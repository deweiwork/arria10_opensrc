-- clk_buffer.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
library clk_buffer_altclkctrl_181;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity clk_buffer is
	port (
		inclk  : in  std_logic := '0'; --  altclkctrl_input.inclk
		outclk : out std_logic         -- altclkctrl_output.outclk
	);
end entity clk_buffer;

architecture rtl of clk_buffer is
	component clk_buffer_altclkctrl_181_4ev4gqi is
		port (
			inclk  : in  std_logic := 'X'; -- inclk
			outclk : out std_logic         -- outclk
		);
	end component clk_buffer_altclkctrl_181_4ev4gqi;

	for altclkctrl_0 : clk_buffer_altclkctrl_181_4ev4gqi
		use entity clk_buffer_altclkctrl_181.clk_buffer_altclkctrl_181_4ev4gqi;
begin

	altclkctrl_0 : component clk_buffer_altclkctrl_181_4ev4gqi
		port map (
			inclk  => inclk,  --  altclkctrl_input.inclk
			outclk => outclk  -- altclkctrl_output.outclk
		);

end architecture rtl; -- of clk_buffer
