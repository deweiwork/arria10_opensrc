// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KPKh8qTKhsaxWJw4oL6mt/XnrqNVb8FoL8urM5z7ZzE6EHQm9kk7QhSgESWbdeHj
jlgqNVogn2ap9ASg53PU94TW6/vWuNspKwgaUSR3bWa+wRNPfiSZcdAsTWpWHDsy
6OU+WLeuIG3X985vBTo+ELhVYpY9+ykKQz45LWmNGKc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2809888)
9SbsSFqHi0z1uNkyFZk1dHFii/TS1Q4DfWI6pjWii4KR7MMXKpgEfo0kDOi8hyRu
gFjU1g0WljfKoEqkP8SN3C4Hgf1VXeC3Q7r3XDBiGtLfyEb/uem3JyJjhwK8klTZ
XJtqG1fBLhQpFtGP0Roc7GSyDjnm27V0ZDOA47eojF7UfvmhaRL3bQynofzh+rwb
9uw49dgPvJS3HxlJ6IEs5swO3iw6AhwmJBZxomQNTnuwZBSmi2WEXNvYIZKMCs+k
aL42akFuNheSOICdbhdoYzZe7+6ixuW0wRewmMBDY8C5dM6nrI4JwqfFBw8ILD5m
qJvMyOt6Frb027xeJvhhdqa02HFGT9Dutoc9yhUONrcDXU4kLOtkgCMBlTPEF8LK
uxumlYn/NGbBbXcauuhzMO2SqMS81fqJd80O6RR9iAUr//VZ8LX6cpYohchMY8g6
m5Fd7nktP18Q42O4WkJ2LjKhk2JnD7rrIG1LG94gHfP6oxr7DBRoW4EjVAwqwJ8T
EFfQj1JbKPeF+UkIOWN1UkSEF/jqVuiBlRYtRToClL1iEgFAIgikenBG+AsmbZ0I
NdGRYR+rgI5EtTmX1tjK10CsAOmim2jDizjn9HIaJNdycfsvy2MIme24UFywtKnr
qE+OEg9QjKiauFFdXyb57ebkuJeZYRf7Vcy7iuISRkNv60MyA2QGpPWMz06ii7gB
YN2QYpJpR83Tg6E0L60VNdddR2TZlG4k7LOsgmUS3LCSVtEKA77MMQQpGuSPV9rs
Z8JEGUf6pKUjjIjkVdvSOSaGaoynsUEbLyuuV3jBvodDOrf2irVNqvOYfhTsSqjC
GOr29B/lxXtI9C24qO4vKwFYDyAB+7yT4JqWP67W5MYrYuKhh7q3xEi7eSWpi+Jt
mAu68M7EpgnepnvAkzClk0qkpGq4+GAajVgGeBd0jWBup3BGMhcF9Y5jYOz0ihxL
N2+blZY13/dTGTL36s1AQwyxmHgWx0HnYr46TjeccuM3BODrr8GijUhN+AO8300H
a2+7Vm6vv/Xb1Ldve/DS2DIsancLRTpa2TSiWo6TFA3tsC+ByTVOsVahklZIEUuR
m4q0zEoeiOl2J9NfqymBGHJRM0nMR4ECM2Mkp9aHRQthPieVG9ndVZIGwOa8cw+o
TA3CoiP6YWpe2tsg5KCF2G2yiE7SKQlWu8JNOgsJDvIdYn5BJkeyBNNOPzlsc3F5
pb/BFHI3vZO1d8rnnWi/FA2Bf4waeST0XST3/XJjnNFIYMgbKHvsa5asHEaSyLM6
Xzu7HugoP+Jc+CsF+mBMPQZ8yRadjjJo530plvByxwHsxrbgzkM5E3qoPwv6ff1g
hC0IQfzJ/PlVtLIk7bQ165RifabXOJnalJxWMUW1XDApy3sVZh0IuarCIGcvu/FV
zyzXhtTTDLjciRgh/suzmR/lt/5Omk9qHG6UeycGE6oEOo5yTejMDiRsEn4cqf7n
SQMjWPhtCpvVAeOE4CplhRcZWLWkm7PfdJtV08+ABN/eJGZBVls9/IVybvNTB/Xf
wi7WZv/LqOgNebEbst/aQsPTQmDsNY+J63qO7A8p+eywX7u9r+M5R0Zfhv1YhxMj
QBj+w7EW+Ck+eztfKs0V/80kZxlG9bniZYEMbjg75viUqJ4bQ6+lpxLqcly0/SV+
oFhjQM8G9oyh9+oP7j4aCrrHfDQXG3zUrnjayNKeLuxwu7FKyoCCw1TdlvfkiAvA
OKgFl8sXHQD0laLN7gZ+R9nHBrsWGY5PlYQHn/428oSZZe8M6h1prraTgVMfi5JH
zc7fRZH6zoU793Lb2froE2lL8HGvMca1uUcAIdnItI9ej1kFXsdmN46mcwMBZz0V
RS2fDGuLjDHYV6jwz1PiaTx3jo5IoHCPu9rDJhPgXSD5WLrYzJHad2kgaX7i9KCQ
3eI5i+YyJCcULg9f1Hi2TUTVymK7I3HGF9KfMoayya9/Ps3PKwAOUDuf4jrMzIAY
es4bReE32DwKmxiPXOa0yEkc7Vf8eOde4cH5QdMdlfcndISzATTNuj7Iy5KCbWpy
vAA2lmIJFXR54MOvcrB6io5oQ3CaNyPCDahu99R9yV4TLtFMXeuzFeFt+rvQiWCj
NeoYiEVYjk5Rkb8k7JnMUFeU37//Ey4kOiHUbWlReSXPrULQ3jK2SGyIvTvIrLV2
2RUEUHHxUgQWWnYhijuI27hsqxunLnEyPhqFifA2cxrVtFpmi01r6jqATKNd7qsa
vLo8hNoB73X7vr8n7D3frazEenDiuVhgiQPmQSqTCjFkuUFcQrPiWxoMdgRhVvBG
O7e+mWITpd8VieBefBzqqC1NF4exTZS75/Fg6f9fZS2TuKGHjuIAreza0Al1sW9o
KJhcBmoTxFQnXRxlK/gyhR/tKGSNsO729Q752HZmu8UVqB+ntqHA7XndQ+9Sp6xL
BANXsR/7UcNtKy5mV9xWRgxcBW7DGbkiFn8uqb45PJYN13hxZIc0NbMmenHGbvrM
zUKNriBa2B3xu2HcWwDZbw86NuktaOgCtuL3Tc+w9UXgBgspZWE3pp8W2U4kJvE5
v1/GUOw3qZrQlFHeIzCkDFSp0VmaN13xZ8gvwExovkBXFIZc8qI+7vxawwyc7OIX
3G3+0zL8RYuluZKDDbh1AJ4Kzkh02liW47a1+O+ALuLVncpea/UWtE4IYTIx5g/x
AkNM4KKWzYxKjAxSROWCFTWII8fdOxJI1JEsRKGqXhbJnFkuiS7cbQfkPe8UKJPx
qLz12vCXHEB9w1ZY93tRSKz16CyY+rOSXFgLx5HR0t1BKBrm6xpxfjiUJIJlvzOD
NV9UBjy3p8LkDcCP7HPol7cr/Kqs+L8qmB17u/prGX7HiOrl+/MXAqzI4mxluK/y
zncBIH1ZQXyPHpu9h/3Mqp0j0mYiS7tfgdsmjKeejgLx0RxeDXlDlYio1PTdchjb
7cJTcLMB5HOq5ycAHmw4TC0fs+EBZIQbC42M7HJgwRvfgfmkdDA5kI8gjfIIhZ/j
XpbY6DCPmJTDgdy4CYsdflk+y8LRxn4g8tcBGWYceXunvfkJS7TbxsWtpeIT/l/l
OoXuvsRl3iuM2BfygBwtGTp6VcPdr/06yPblsZiWZi5q5z5QH55ik024fhEwPBc6
yFcDX7c664oS1d725PpkhqWcnuHiE8y4vQwx0yqhujeGj8B2rvSE3r3cT72HjnN5
lpKz/Q9dsvMGjpHlPI+GVnkgqvLcfzbS0l1CRTNTjX8iGaCvFFpoOk+08SJji3l/
SyO2FY55v/mvgV0GJUU7vhiV/vu25PxNdrBlqcSPXOBII9BQWyPml++erU8orcBO
qcc8mJ/kE/H9xu447pPq+KGxDpC9PpnAVSJoucvWxfAhe0LFBL7KqLFtSpidqg3/
SE8NmaQj4n9Kazk6omrUnBVw4uiByi7RYva4GBfBFeqqPtakDaWlGPDaIE1G49VK
LIrDiM22Cd8nv/IeN51JwQ9p8aWIOLpjEoC4/I+nLBvRA/WxG66SsEAG9nryc7U0
fH095m6dCZ6ROMRVbR5AKfwV1+nUEuB62nAe6E+vqSrYe1oaOvMMmzKmM5LNL52G
yMhZgkur3q7RQQZhmipHnbdX+m6j7/MsHHldvVG0gwAOuJHdUpQ6HiVFWMnHVo5r
bXUPCq52kLelC0LIwAuNcDKQJSyLqp4yN261u1FkdedWFn0D91oHPcsGGRMbsP3Y
kw2stahFmRLSurx6rwY0NLQuv+2vtBwZumCFfWRB5hOKQud9dxpRljg6RZ/B9d5M
uPzTpuDza9CPntn+97WuKHeJnwmIPqKBzpXshExcXYG2Y2hDKGzd8SD/lHLI+/Fx
nS4u5BFzkv2Gzh0IS+LyghhuuPKpMEbYkNfftUpn+2RxYfzHN3fPrQWGLya+UT01
HpB6hGUEFV7JM8/aJVUm9DhklYMWOFQ7S+rxFu34T7a1TiISPYcC/107lYbkZebb
/40ut90mg5WGbQoJEcT6hVu1mqXyEdNkANoTyRLvp+DEn5XYpEhVbQr9u6B758AU
s+JMHMQTXUaV7i+phKDMHpahgXA5LxUYDm9gqgcCdlq8mUOFdb2s8Eia54XqRzIE
ztZN4h59akjezS5oKtxOtNgp7xAGnlsMelWz1VHH7R68Gvz4jkFkAqaUn50SNltf
WKmre+/tVmMVRBtaJ5VTg8sSUMQYfP0ccrhM2KVs22JD1hjfjHjQ8D270WFKlkJI
Bac83uuO+EfiY5sYTnaBih28cvRXMDNXs8jmMxyVQiqzXFy3YxPpLNGtXdcsYN4Z
SFrFcelzRYf6kt/HsVd8cSCjU/57RYy5HpY/Frp+xtrDlPc9V7seO33VgmAUjQy3
CAwyzzNBNAXJQRZQ9x1zK6Sc/S+HQgFtjac93++l4tBhIAzX6r079alscH7mjG/U
TYivST4evlu/xNK53hLU6bws56b2n3+FO2FScMU7whFdeNiwN4U6cefdNBq7Us82
k3WwpVVd43Ls7ylcgw2fHbtxa9U2Is+wAFs3pkl/y85S1nJK9o2EmaJzgLrP0X/k
TAdjhpmbQCLPZqDQFswBU0VVI2KUHcf6bnyJcBAMfH8EhhGghNY1y7gc8d+M9nVu
Zi5OOJ59dkIgvsAmQ+OtLcbmUBUH0/gDbkCfmYzTTORdes9iiCY5XDHqlbbVGE3g
ntCijtbKPKeRP01SNTR0oancxBrkAM/sniR6L8ZvNjfLAyTAFqAoxkBPMOeLOKSo
Ggq1oUAcwJeA4rvZyoja+VTxqUQ4qa2ceKJyebSwyThd2l+3fdniPTOIzEB2s+M8
eNWo3hi7/f87cNNVRVcjUMKJrVD37DuO0jp7HS7ysexNJvy1ixLpBOY17KmFdfoT
t+/u9TLzQX2twm8AUSr2tr0FvXW2DeFeIPK3DhwBT/ryKLHJgUjm0EJlZBlQnojH
WP484F9XIu6xTpVUtfNPWsVDa94pApGsJqncTFD4MI0yuAlANNfbxe7QdEaf1bm6
OeYroHXdtJCuRAo6OUpohcQR+wYh0HWnqJfO51d97CKpRfOaUt+796GAU/46lChv
GJ+LDcqBAlhBBx+ZgF2DNlLZep8o/y2MOU3fOGL46ZXJJebND1S8KOJRbJGh952n
KDyjefxOUzzy6HNqJbLEeZ7tk0kfKVvCt1wbCUsnrATjM+UfFRQK+hZL2s4h/vHY
MxHgyB3/qTHzj8y6zBVmUQXXOU03p9arDwzYsnLimdPK9BZKx6IF8rNcRoKYaPUK
tgms4XdKdpBRaMamtyt90Kl1Xm1a/UCIL2dGVbOjNMYF2i6JK94MZLxjcA3KKy4w
0UbD6/5aMhMMTriKb6fTyqZ1EiI34h4TdCO/eMsdYVBYKYU80vxF42a2cC1Xmw7Y
usumJ2/A5t0wX+IiguOkdP4M+MVSmUHX5FXOa+NmyZ0omKbIc4XrN/fQoKNdukSF
lpEdefUWwC2eudsa/PtRMxx6l3NOTG/CsMxAPxme7Wj22t9zsur2N7JnChM18Gsw
LK0Ws8bvRrTiqbfa1pQEjpCme2tGojVWCX6Ev3IjN9AN8w1ORoJ6H7oRoAF0DYRs
Hfv8mHBGnQLZNhGbTa/LeamDQ1paKaoJOrXVz4K3ItSceD41kzphUJsnBRxIy+0d
+4zedemE7jdYERKn2DKrMBu6NO8s9TqTWz2T0dXrCFiImK6q8N6YdOP0ESJ4JlGK
Bz9cDKf+ekQYzIASDMQCT24vdJi35SRGCFBWV+5tDnMEHq7F0sJN01qJ5K++voXk
jPOnQSR6p7ja+DASWg83tWMQndNFnyGMRXugx4LEHglR+thVNi9Cu+9Oec1fvCwL
baZy9Ct47y9GORW3IAWhaPXmYkOYnj1usUCM9w+uCOhJfd7DhnObr7PB1tTIkXXG
QrEkuV7SkjfiSjC1MgV1tk1HuYAyOyTZx35bz8kZ0uydt5x15K3ZdYlBkl9D/Tx9
qvrch3zt69Wf8eBBp+oMpWBgoxJzh/SZqwW7oQetQW5RghszB0xZReug4j1rKG95
GUFzUs4ajKhmXnWBBSJoBDW+VAlhFuVz6XnmW1mjn2SPyYG2N9w4uy2rKDuCPhIJ
rsvR3G8hiNxmF9G9p50VZhfGEvKrohY6eORUXu0e6vYhJhkQgALJ1y2p/J0cD306
TcWE2VZB/m0clssuyQQYXjZIgkJqAju3W6ueNvpN2ieO38D/uaGOX9JyFUnq9cfs
MARSDBnmY4spfhRIcZstnQEXGz6cXS61RBQUDyHuYbcDeQfTNY8+WPuqBOmjByfW
OSrpPNjotBJ6amHEQIswWDmyhb2lpfaO7rKrXUbDHqoLfaj7b5fanEqVu71OHTfT
yBZOQ7WQsIY951dkInKOdGbdfKSA7+roblO4dYVMC+8RH4J+sgseLZMaLEhj/qyC
wDwsSo83ND2KTOle/T5rqUVq1vE2xTGnXvd0IaG4b/phqN5x0TbcRjxdR5BMV7Ql
unkCcv8kSa/nP91OrD7pquXYYVhdevQcGsXkPEgeQ2eZ0mRnEUQhSADziN3/LIE2
gBMOJ14THGsFVnD/GYg4MuQDozMA7FpOltSHij/O7VrpuRgxgRHJJNkSW1cUwc7w
lQOuTGCc4tNojSRhICpY+XlQriY57lU3wneo9u1U3ylxviLhgmG+BaVfx6zNm0bZ
B6p/225mJpL4agh3TNeQFjvgj0G9hda7xGYY1xbgRJckbWxp7HenjYyctjmAWVPV
qIEfcQ/Wp1MeiYIRTCKY4zd4dEOsw8vyYea7LRS7cxq38oMeNJPdIWUe9TP0BGeb
jNFJ96EwJfHBXCQgX3VZ0xFSttoNTLmDG3yRTO58AtO3ZHOljAGzV7JRLtfD3Pvb
1OpzWYAo0as+MBYA5iOpLt7rSlegiWKfhgeUu2IO9nwfb/2OF6JbQXdl9tJeQetr
rDZUExK1bYrB4jf9F0+xVsncKFSvTj/s9RYSwm4qsn42444K+1cqce6vifZzgJRk
a5me8QSPqwA5JrpprFnBrBZfjNjybG+0VXMeSzzSJtS3+k7vQTOIKphMhAoYLghn
D2/T4SF/U6oAVpFAmZDiJ2jZuBk96CQV/C4de07WPzVQIZ7TbRHdf7cVJRhchlqN
eU4Vife2/A7qqD1NSLd+BmkImLdde1d8yRA5hObKcsXXbJzvwnyaLFPbw1pzE84o
e6JFMMADK+EKWqDAYItlVvy81SBYTggVxjSjRJUTTsvQVvzoC6jNkP1vRIU6suLo
66dU0yxQArGxfbzffioBZWRjMZxf+DNVzIBybafyfIMOYtTzpwN9OED2KiEJzzoX
Ujh1QHS0Hqpp9SFcz7/miFcdsjPpnb/NA+9TC86uhkVt2llfErVOaZMMoqGd2W1t
zH328AHkAfryAIazPYY6/ibjVJggorDvMlaj7bm0GJ9cgH692qsCLuOsljN5Z1od
JYXYYn7tk1oWTGJOQ40R8Ai6UmCWE7uZZ1zuk8aq7ZPVVZTy6R+bFX85xfkqAEPK
GEA5ATTRIr3tPfUTySluMrf2qBSuJuIQ3pWJioTLVW+cfW4p3Uug5M5nSlYK1NFN
ocRmzyU56vUyuyBLI72/E0OYSf5bdENf0WXj1RtwTF8Ig39tN6NZueIUF2q4cyM+
d3oBqwXgjFFutPXChOd2CXV4LNm9nr1ZtHecpS/37bpFk2wMC7DQ7dsYmk5Rlz0h
HjCl+jrD2k3WFoF7C33w7emjuxjosn6YvrvsOwr3e+jSyfcw0utQuARiWT7cdqFm
JnGdyBSxaTpS6GM0IBxyEaEsyZtKn2B/Xrt8jw33a+YbGqZfUGk/N2l+3ZcbfOdw
Hy4YZpW+OhjpDwHbWVB4u8uaaODZzJqQIh+vOZ7dM6gy6zBWRGVWW8t+x49WVkoY
b6K+Kw6EdlsEtL0fLcvP54QmlSslYuTidvCJ4+M67mTOrKWsx//UOwU0jIvhBzFu
gw0zIeWYzSVDkhBhiuoYnhsZqM5U4+1Zoy2/daQd/j0PGLqoZh/V6FUEpS5mVwcc
gGYNQIbK8E4mMIxisYtGABaGLxGcrrdNPLvazXwmz7lhO+qrb7H2SpJucZGY6gJt
95priuHB+cmqaH28EaZfVZy6oHFypbQMG+8iwIO8qzxwqjxAagXcqQzVi5MSyyiD
fPHZftWuQEhQ24wqxn8ePTNdp/7CliZaOQy/ZgWE6G0mvrYf9PnLMcWl+h/YYzPm
hh6k4yPV5mCP3Dg8+FHkXfGLqipj4u8TQKmsRqNfbZ7+gqtDGDTZrfd3+0WE3+dy
2Iahg8sp+QnRGUde4btsnSPeq6RKHfHLfG/aRKqx3fIQrDRRhWt5+kTq1Fi1MMKH
5F09z+PJ8vGyHsj2Spohn7/1kyq8fuoeZmzSZhybHk6rYP+vBpCZK2cIl/wtXgMZ
jhwt9kkKe87LIiTxBsTry9pwXGkEX7JJDTm2AovqiRll/J7KShZPJiFhq1kCHo+F
W0mLkzpLqTDICvXgrmdnpAKKtfC9aMA1xcRPEy9XHElVBaecDJmVwguAtcLofrm3
fPG6+DClKELMdf2EIT10wwakudKICZhb933wOYSn7FwtHuJsjW+B9R9ZmRtzps7Q
IzsNK/qPgYCrVJK5xPXSmMwIf2gouIeIDy6GnPjFAgONmhAW8lww5WbxXsbcaVkx
pMBI2NtsyFLLJ2GpYQwI349OxtkzkVaaY7lxUB7lTgDZEYmpDaOFbWTOz3z0xVB7
eJuGrK3pFEGT7LAcrSxxglfk2CWwYRbEDlqogt0/ODRze5I3wIvJDP0Iqle0gKvZ
0BU1vNKLU3IJWxtzsLeVBXBb2JvT9rkmv4L9ySvWPcSeSjxbdRYcAYPFhkw4yHbM
EK/QfAXpzpOqRYehZw/uHizW3r1mpvi7PQccFCR3CBKDeFGBmb4SjJISn/+eHxfA
KRqRi8BINj7hZSSc+lufEd7+4GCpFseZwJ/eAz9L9jI3Fg2tTCQN/e778N90Jutw
zdq4w9dUkTjKwHNuc3nQ/L/YDDdCrxgNrxB97knLtFHm14d1/6EHM0D4B9D4105g
EevYx8aO9Sm+RaLDpeWPLY0pnc0J8f0oAyNG5/GROwgPVAdVIAiwUhyFAN7cN/Fq
UGV2sl2Dtok4VU6tw7j9w5OT9gszYzHJqEqYcUlZUd3Doz+xP0RVNhOcw7b2NBNz
l1ZQyI7VKlKHspuKEMivQL03/dQXxB5HdEY1qYB/dZ1XMKquRAM5P/Uo4SpgfbBP
rAa8ElipXDd7mf4LtsYrI1jjGwygCCiPRB/Vq6kWuzIC7G2mMUTHRqMCXCFq96xu
Vmq5bVEidVDIZUh/pyycnGgTZvwgJ81IHsr2muCpPiyNo45JMiy0MHGWACfBaiPf
5e2XTywIuIoujwoEt3yrk5U5JubR0VNOHBGkREv/n85JkoSY3wR0eMHjnMSOfKXO
WcUc0cMrxe0WD7srydXSNzpZmcXgxJqposQnB0YmRRg7gpPgK5Qx2mW7PqX8dZbt
892Sr0xIayWGqBQ6lRcUEFiR2gPbjCjcRXrG7ePPGRyHHeflXpGDwKa9nl8mwMXU
bkrKe5yeaZ6jCtiC1uWvARSrj34IzNbCd4wEsW1psSAk7HjMV5b9ZsRpfZxsloGF
INIb0fq9cgVL0pk2L8t6gYPvYHyZgawPxzzKfLhgxG7+F+X1Qq+4J1D09QKrvoZi
WUSU8DdleDE8x/RFOD/5tQYHh4Tp9BFVVqZMbM84h4aoBxIbMvvhNO9jJ2nSplR2
rMnV1wd+jBaD9Spj/LAaylX/Xlce8TGA6w9X6Z04n5J7eQE8H84xhjq/NVUw394x
1yHQLZ79QTnUFyiAb8fHpVnVxVIg1FXqHV4sln50juThB/KGZj9WbOws2pLszdUH
MH4EHvtRWPGYrvwef4SY7Eeqe1XPZ7dZIco3Oq1rq3ETG0VhrtMu+o7szFyvozd5
7xc+h5aPq/He7ILux0UmSJHJDW31hjg1oPp5wyB+Vlvc4SzffOETwWeUXm/rfGXn
HhgOmXwPqX/KP4M9ar9WWLJTlsSFiS5ENAT1vR3LeQ+dGW0K6qfkNVpfc3I8AjwW
XqVhNOWe9Ja40BydbM6X8jaHex/bjomcHDtcrphC/7DPbTDdJjTeHV0xZVawBGi5
7ba2/kdi+kpWNmwukKgp2eyZyc826RPmjie/JgyEKs2mnUNqqq111g7cxkzlpk8P
gq+82q+pGfN90tQu0N6du+C+lO3dZXexPpxis4QR+qqR94ABWJ/GP+N/+YAfrrqB
0gaqcczoCa2KgK0Mb7Erfq/H9dOiJm0tLif5UkO3IitUetY4Ah2J2hJbX9DxJrMK
FoA0xeYh+2eW1G63PBuILwOK/UIL/iCLczr/p+LTynrJ5Vs012pFXt2L3PCL+/9P
Jq+QkWPUnN7+Cn2CvaWixYq5sIGKtEP/tWooDYcpo9c+OSLF9XYlEJHKLeN/m36C
Xdv/vUVIo8XEk8N9D9cc9G538cHXixD1/8QgM3GFhA0g+NgSQ8trvB+D/lkznq/G
E0KDC3utw8ZGk5v/upI3MJtZMo4OAj3wXsmht75GeUQXB89dqdDluUxn4uhTssdh
Au68P3U+jUjFFWG5C8CivhIVT162xvs7jIFMG9f6kmMbgB4VyWlNcdUpqPny0USM
jzhlLU/i5ahzsR4chIXmMwu+Fa/PrkovrTntrrIdzF04ViM4n0JpcDoU9iAvNygJ
LoluRSIp/Y9uMrfvU+3v7lUiBOgqkAMS18op3lB8DSQE/7V9SU8dTQLCnXvbjy0Q
neiy9Z7lkEtnQjRd5WPKWqagmvqux3YJmyXzQyBFeY+lzbFXRQLR+vNEtKIfil36
JShUquH08IjxcYH4A7Yf36RPbY9ckYfiI6udLNtDttCjFoNmuzOFRzaBCQOebCos
e7XPPy0Q1UseM158XRZK+9MViAQP6VthcoOoc0XSTEsreY2V2VRkHxfumBjKHaVP
AeDKjUt2+KnuijJx17/5CWZ/sYXpovTswIysatpfOpYa55cXL14GxKVTSAErlLjH
SVnONJN4KqxAEBXqaLVaGEo/FpuyskqNt4futwhJVcHdEbnbiGS3taYXXeq5Lc9o
sFXWu/q1ot4b051lcIh/vwcYp9YAaXH1IT8tmHjZI6solkhYbmF8qxA62dhGPqbf
qfddLKZHIhuQg07jSdfV5JlTvGj0vcfDDber2EfdeyzlCLgNZ55kknnbLUbvzmkn
hX6fKXEPSPZMdFyyGdUI3dhxT6RszHUhQI6iaLw2UjFUFr9uGfggXIIyLw94yPEZ
Q5gwjqu5Gyay8Mx78s/BPAKCKshqcxhH1JSoUj4kVPLHrABJW8ArOHrZt7g1szWc
2mpG6By1jobMwZpxBAS/qujSEKUMAKSMtxxQKcvdoSVp7n+8C3FY3AUyCXnUGzsK
KCLliFjn4f/f42c45W+lIm3PF3Hgmdg5s1Bt4Jtj8cJCrlzFM2WqPCIFdmI+ivH0
9WbSOsxNZMJJmFoKRvqxIlzxHBSnYrdo0q9RbnGv68d6y6rlcuIxWkE/JGcJPGo5
8rS9Ta3W0rlnQ3odpbs9C+ErRkvONVYVvrjZMTOl+8GG4YPoMP+J5SGibmH4yzWb
+exlNFJ9A97xPu6WW78L+q9L6z7S5L6xxx1nCSw2ARKa0vbY2XRnLFmWzGwl0r9t
tdG7mwqjc0wrJmB4tOeWnaGXghQpOsVsg/A1gMJYYM63KPbwsmMbrMonf7E2wNIN
umndwaeCmkTyjzVmu222fPzAVcfPVj/hqN5f47jU2JkO5Bl9LYDJQnf3QnJQIP74
sGhEWBT2O7magKVHgMBZg8n4Q8LFf+N7aDCDy6KIxLgib0D/phz45Z1mdJ3LIRrn
kFUhEQTJ6z6OsUPEKCqGE5Mwt4hbNg4idcS88R7q01bz6/7oFFZ8nucuJWGLUZHE
osvfbEz3ywi4HKw6LW4V1zSiGbVS4rlMqO187u/ikN23dSZMAJNq0Bwg5ExIbdiT
3PKn25dUGNVSzYEmMUwTdcU6awqpRP7ifGI2NaEmh2mV+cBK8Q0OKhd289xp1rmA
sa4Ng252VLRWHQ8N7Iicp7Sxcf6LoD7logjVl/Ple3BeN7AAqxJ31/Rxv2Q/iuTr
i/x7rpO+1vocnUxVEIvH/o+vrM2/WSsUZ835EegxT5VZxQtIF6TC/JUy/HYYI+VR
WUU2B6GYYoONKxTbXNEvLej+4Kc+tRZr+S+zThZixlgg/XA1rII6xBeGDlIlAKCB
KyzOsCeoGLRBXtAfohNfOnikCgJVAWYFrPyuFhijN0ovz+shKvoCqgxW1ngYA1+S
HTqzGB06jK2+jtOTNzlxH0FUbAhCKs82N6F9KOhCAAkGzYLuTTZ7JlPg2Q/L3epS
U80rxUQUqc9zj7t5tdq9XfanIiIqqEunY1hldYItIctzX7D8YsLfbdsBPl7BzY1P
/iBNRUKgcra3v6jn1Rhz6UT06QpFyQXXwh5rSZLJZiZZABzGDT6SgAWGJIuj1TTX
dS6pGmvhBMGbRUAJsApsxO8PN8NQSoKyPV2ZZlVhjokpP6AzmzwA7/ynZBexHFjX
+nDhvaMB/dfdIJUN3MhRKlmjslyvSDspTWkmBQ6Mp5U6HFOJ85VeJgiyX/TE3poZ
UcRwp8HGge1D1ofB3+aFJxdRyb6iSHSUmgTyEWgAX21u/tKFwqTY2LEJWdPvUBHa
VITjqCoycG911g2FXzcZlOz1In2ErsUYGD/BeKojlUfsmafJ3YiMG2iC6lBmLqXx
qrgNxtl9pLVa8sdOMG4ApHTHQTDVYy9lz6jBiET+tOqZ63hPPz+sPrZdb3KxxqYV
vhVQmyt3pgvWhYHU+EqHA6PIb/ecedOncv64o/rhIIWhT8f8vNJGB8plS/W8byJ4
t/KW5H0/easGRp+PpeLOknbsnt2hDD4usdLfVNoTVYfEHkbMXJpnCdlaNxQ+z9ac
qfAUMTHY+mDfWXHCZx16NPjaH7sSCi/6beJXtr8PlUJj1h0nv1w9ikXRkpr2cTcg
hihsraB0/qalg5QsjP1NqIsbNZDCnMQdyJU7k88TQ4BZy0fhlOBbwE2jE9k3M+lf
JvFUMkpmVEri8MYfuHqmvTDIv7rgGIEUF1otd8xtuVqfdFOHw6SzeaYiBAvYk9YO
ZnbhVPGXK3xk+j8Odof4txOxZ26MYuSY9/B8geEoB+IQs8n8dnaJZWJwt8A+AqTA
HMvf6rTKHXqmsxq8RxvaS3Mp7jDb1flWsufvhQfBKQ7CkLY6CimZAonpTeg8g8H0
12558eQy9dfwTzk5in12w5ky15hwKLLmstXnxFMR5u3xA865Hvke8n5Ncy4V8O37
jw1bq2dVgzB5Umh0lMBeF5dJZU7W7Of2oUEk3CpI19hU3nKiYfpqYc5E6x4up138
R+NtpxqujKmIG2XoT/xtAgk7wbfEogCNqw7YdPUZUyQJWShNaTbWGupDX2e51mva
48Lpu+BMx6Ij7CIN6cRPsK4qHOB3gGFK0iCPZzwnDOZ7REFNA4K9tvOb/PQikiTg
f9Zo2+5bxw7jARMkM/BY/RqdVZMNkxACVQ0rcPEqljyFRo/fubynpw8YdESyHqke
lpyw2n8cgbWDK9SZDzBU8nWDVuXpTj8ktD4Vaw8s4MFxTJ1btbj0rzFjGY5NFwWB
alIsGVr/MdCVaRW+hWkZXW4pTgMq0hKQiSy9az0Ssibs5/aQ+vDF77GN92mJR2+x
ezEAyLokOpHKyTm3gLBbhJD+MnE12Jy79BUsuHPeg/wzBlLIlRx/5WfW5mTyOOVU
k3d+qFsXTR6r9SSWkPFxS3Psan6iJgWj0OT5qDsK7d7mtbUOdj/nYWr2T/uBp06y
QcM5k31mpjqrYqPoqh6b8dCMql0hOILh1CFTbNF7O83I1BXcCfVd1uPRNkYcg63C
jFhwWpHH5wGjC/pSBF+87vagZVGtZ1JouW5jb+lYS9oxSJGRY9m/9OYntY8r6UsY
2h4xvl2sn8oLHudSxSzcAgRIwB7STJ+qo7i6lIaH8dkj5eCkDEhW2zVcsD+f9GL4
lUkvXXWDXqjbjuQgI993OfNDhyqXaJVyHGtQNqJA7GdLuU2cJibEN6Jt0Mj/jZxQ
/vkOE+fOhXN3fW8hXfiP+8CEKInhC+h2IhY39fHvqji/gdXPfYdIY8rddRxZDLt3
WgopvWEyklVRTN7Xoui4jmDIqmmwbhD+Nz4/CSgoRRL0QK44GnfYZbr3FnWHMlZW
05IB1A9zBHg2IWUNXqeXx90QNqRdq5r1YWvVZGE5/YNa3Ec35kHLvAJlsbvxL9Ig
dtAOvw4HOt7RZyqvtkZcdEO790bomoHUcgjuIYDoxUsa+jqWYQeO1fBGTdc7HOFt
wHpHpwyuVrvrjQWlkqLIv/1J3/5IjqFZdUdBDBfvjmUA8/z4OfV+gqELFmRB/3U6
UL92o7Yz517sVX5+BJVqSjfPl6KqQSMgFfibUvK2AG8LT0q6S8Cd39vIogAtgZRD
j8vrWepGZluiYTU5zDnnaOY7eq2HbNuaXRsi5D+FzLbz8c90Hgy5sTgXX1bdWHLY
jnQlnXfFdbETi2KTprf08zpJcWdUqg9qkfAyQL1BT2/ebyCq0O12imeMCR0V2ZXc
fUCMsJwcPoLUkfoSU/JOacIkwshKsIYPKY3cr6UZvpsW8aUndhSMvAtCS94qeDbZ
1okW+nQR7EpUM0BEyNhc+HtDq/cuHSQy35sdgp+KSSq58SIG2/+CgIFTXMutZPLN
FvbK8LGymUWyFkgsLrOyBK0gl4VAlfLtL0JZ6rk3lYARpKERxKpitBM0rAev/ss4
eAqHT8Vx9bpLou+aF02Bf4JTsZaSvI3J3SY6GeDaCvgALs3HFOJDUFnNBKDSaQCO
uoDalHwYT4SydzU5TiFjKh3yLw9krJZIXTqDRnq9+5crx4EhKNbCDHE3oQOvGKwg
Y+GP/MmihCB2SebloYQmmgvynWKRzoh8LxHg44FRU2QisNCJ5Hxuj/RmNhE0lNiF
+GrgUUtaLwjITCAEzN5bfQ+/iLo5EHvtkh4JM0x212blLBuyEGKNI4NBcPj4Tuah
/05YfxxbXNXNNCqocElG0UJi0BbuzWVFNlSSZ027azMNUeYAUCFh4KPIVgwwk/pc
lAdP7ridFOU3y+KD3CZ+a4aXN+iH7Ocw9EI+FGI12tteXdIgKTU5bqrFCDO0u85N
HYmgNWFkSOxpwnp2LEwzGeXsLKnjmiiYqNT7h1WKN+dcs/jt9paVVzWFViOmL4Cc
6ymLQhUU8zgOAbDQD0gBqSEYmp8JOIZwN3sUC4yiSkfk8dFWbic5VOyJ7n8gShqS
vyfyd8xtorWJeYfYXaCFmfyohij3axYFFCsL0cPOAGn4j9nxc1o8z8NaHUSdnBhe
0T7Z1X/v/PJJHjeEJ5jybSbsvgJZPvCKvVLlep9M6VK4k5Cpbfh7tJ8Y8G4tlv9I
sgTB+KzbE2DT8t1lh6Bw/9yJ54Ks/aPheSnzcQQx3XutSlegryanQ44ku4fb0OF0
2zmuKdtSh8JfjT3BBlDLOY/bqOenncY/PkrTJ3S53/ME9PPZdM4n93OmnK8KC4OQ
T4M+0q1TlaDz37GLAzlIAxDF7fN1tLwzqbbmqo4UcRyT3JLfBU32XO49V2ErwL8v
dYgFxTpTH8Bb8bQWH2TazmsIMXOWQKSXmX+UKo3/FN7rgcT+wPfMzxY1lTdlFrzB
QESJnIKaCz+AOWILonQ6IvKw6QEWLst/TbAE6Yv+ezRh5MZY42+pDLkDapq2sATI
TziGvw440J6ZG7O+LIVQetaH5ZqewN2VWo7XW5m+8pKVv0zO6j1P44q/pZG7ELoD
UhyislOvRZTI4SUGHqvgBvOheZN4D6Z7vpjUAonMTzw9q06O0/5avbJ8vcDD2WvD
GugQx4U8fLMAdzqf7qprfvlblbqmWXiWejfPMUT20TCE3F1cgfli26VzhRH/qrj3
sOmv6mmHAjtAP9J97zQ6cBqYYWYV8dA8ZZKe1yV6ag+0j8IAUiatZ5rn/7yGR84B
VjJgERzWmU1gi/ogl9IW4SysFHBRS2OXE3lw1XVvEYX+kOD0n2HQi/5ezuhALRPs
kfE2jfsNIDRfajk+eqB3eco/pkTGYmqUpuPrWKk1Na3bWJmcpYhJhQ7Gy2v87wnR
7CigHl0+8/nXScMu3bpBETlgaNBfbnsZOfOf/nSYnMHBI7DdRl1684khM5Vi+FMB
oUzxZTyRHiDulkn+rfiCUAyyucDKbL/VAy1KP7vVaaykfOYRu9OLnGSecJRtM3jQ
AIXJtNH13pCTd01lSXmyVGDx6P4rkl/PrBKevjNKGFf25Y75+5mpDRva/URoI2+0
5EHlZp6ig6OBLvDMuImUZu/Jx5nzpjl0H3dXM3CwSDxvfe0SZRYORCYy3LWFNmo+
yv4P492kLhE8CFbbOQ8NjJ+2MHWjfI6Y2YYKWhiFGtWCSMAK7CoLKE8gsPqPK8wt
ytZgmr4NunFgV7IPhDgfP0GaLfeBc8KfRSgrthzuObwShGllAeJ6GvXH81KTMZkg
E7VqiJMQXk9EIk9eVCFSDSLFk/zr8sVuOKoeKClSB/01oqS+IOQuFNnaw61LyvNT
05QuNPcLZbM2gFdNBI0PzZzBkUuZo5f33jQJu2dYWJH4yij82Oiv71AX1hjIioeE
KGdIrOYviFEdOy1Bt2UtaHzFTHEhoeicXPKu0d9QE818inC7fBZfKKde0Q/ozzVs
z8CumuoG7UBy4WVn9m4fyohjkMgV6GSgEGWB6aU6ej0IwSdALymSA7RR4cZElab7
JJpgfOjWUywEsfrY27D17+Jrj51Yxfo/E8fQIddd0jRif1028+iKr5Yg5U7o14fm
FoJA/yJxBfiV5SOD4+uG0NfLDzyNyJKrI2Er9237ovH2UpOaXaTryI3FdOlSQYu8
aT8b+EWflBPYAZ5hRavEIjJhLoZ7uHi1mxrwx8bHGMimJk6F5t6hzRG9cm36F/yX
tw+vVsfTqfdCo7jR3SAikPIjZy3OUCEIkVqhXzt48B6kaW263ytbLfmUVmB2azVO
u5u6W5jOyKJuxB40PQ6qLcPrnEvFQNEFI3pqPTDxWh8gVlP9o+O3tqwfH1zeDuqh
4Nq/NKMPSfxKRkIfQ8Mn70uWtzQEaXYCI40xNToU46qqGqFvVTH/TADCBZ3hdff2
9t08AsfX4smN+BnY3s+ifcIISMC8KnpcQ69aPWVY1VuB3hDfHNoQEx+KwSjep4B3
hsoy9lOvWs36o0urRKJ7pCRT3RYJNd0ySZ004flEd7xVh0FGEfKrFo9N126XLS2P
b8rZ/z4rI2m3LxheN/Pa3++QP6uMbnRpDFNKlAxYyRL9PMG8ue3D3dqgX1UBk8D6
kgUroLEo++XisJDiBdtJ07sBN85g43KEIXyJHWyXyjAXPu1e/DYLK5MdFJtVsdwd
dhogPRpwxwO+uLqkYw0e3a0LaKZOi/fWmJMDxwlk5qNTpI3ZG5EcYKDu6udiEwmA
SXHtb7jowq4cpFT6nE1EzTBe2qLpk0K8Whgz3KqRy+550t9x8XFcoxSIYIsYiVka
1+/h45xo0a6WCmUfgFaLilNEJU9A7AOY5AHim8qjao0cXduiEShAKLXoY51HUTE4
xNwg0xwOwL2qqbSaeFk7xq8RHTdBZzBNUpkFoKA3myztQKJkW1vx1GugkqMwhbTY
Piv4F60/kvyI2TCustd+1SLcawl927KTwfnbomhoQIigl2w1x9o26gb8qi17HLKF
vgWRMO2B3R4OYEZHJlgBTe19bLCFiNAG+gBvoJNAqLFedTrjXxqeeOr0u9F9fH55
DwQZqgkvMGdupB1rsXLy7FceV5vAEkKQgFqmWdJskQmFndg0BcxQZNkUqk1Y28Km
H/A+VzPPuT0FEiwgJUAwfa6bxM86KCzK+CaA8GLp9j8ZAm7JR5b+f9NtoOrDXvTG
EsC6eTn+htSBDe17GEcquWDDA4Y0g1vO1iDE3vagYbjirCYPqs+jWQKUCDpw0omN
JteoK4URd6RfWrqPh0XrCP5M+GhsU62rGqOy+gGWUoHidp4ChhXbdN/sFiILCaUr
8JjOIaCZmUn2K+zw/Ct7b7RT85MHqC4KRjEXeypqUM1Qe7W4qVQI/4sjvI5c6+j2
YCUL9IU/nxdEdhrT35IWBP8hCfNIt2hlNLAgZLufI6pp81LKcUF16ejrL+m++Yfp
3Q1t9cw+YqzoXfM8xNURpCnkNgMg4iVQR+4o7H4FM+6AUBt/Oou2BGloo6Ml5iHa
LBBZiJyVJVEhicfTeUhY6UMsMh87Voc/PJq47P4LyX1i72Spmu2KNkLL1YXPD1V6
RK0S5jL/Kr53zU6NvYYZlTMYCGNCz0i4+4Wk0V+YLm6M32cWyShpio8aUB/zhRDI
FvNqbArGojRgbhluEAnWyUpg5SCm2+4SdGXfk9ZWa6XT91qjQrFIz4cJ3OQykPEW
tOX7UNc9uS7BXi8L7TjVcfJ/Ku79Ow8J2m1yJaNbUFnVzLQjUBI560RiZKW3x+yi
KFcUz0wRJLVX1iAxxJJU2+DVynnLOA6XXQBX3a6BzP/VwXc/UQTRQ79jJ82kq0Tb
GXAoxvC//17A+PC13YMlF74t5AU6e0LG4ExYwaReCZnukKovAk9xvYpbVNYlkxtX
THkldoFumuiSC2FquDhuGAciQZ73jWOt0SZVln51OLgErl6sZofBPqqTUR0d25N3
f275YxwZDDO0r+jqqPizcVcKSpzGUT4TFlvLxImwiPsYOd9ocfYfY20nJgV0S4jZ
9H46hjNweDwg9Y0pbbaSBA8xOfijJ3rF+xIMtP2B7qAJnSZIVYqcvPgotX9I/6bB
j9WvyR14S91i9bTZ9r2q7O9o9Oql765BPt9F5XpSE/WcRqaJTf0O0GdGTDnTVgwC
poLN/52ob4SwKNlEvzwi7Xw/wf+L05JxvV9ivkD/J42IQ9XTWekvoKYIffAlAqb9
paDv/3JpLhq+99xSxGkNkxnpOzjx0tP8doOl6ZmtLfShQ+vDcBDrlmv4Ha7UUU7s
J5Dg+kVP02Lli8T111WjpXi+dJZ8tpMfkytrqQJULXhVsblBEeEQK6YfMhqVP4X3
oMiGLJkQw0SpPR+E3e+vBvZT1nc7tMglvgfsDuNR9bTjEDWLzldAz/+M9sZf2XBW
ocHKhsKyu0Cxsjmrr4DyPPUhc60BUyg7edw7Libd0KRLOuh6s5/mBh/Q5bUM8kxC
ydAwQepW5LYhyYYugzCNmowSyixppA4pMxcKKs+zKU1MuylC6GQoZWtBWJ4Xe6Vv
Lj9kbb9DmU+wR0EbevXG6ieUAqYDFLf7EUs0yX8K8LCo72N9mDFM7wZKBPAM/zxW
nEdHcTEN/o/VI0ytzsA12OCyMdhdbVdIZ24dTCUhQNmG/EB0n2xfneDupF2U2cSI
30fRfEvdP8CVAYiihvEhQkroqapemsChx3lXmRTQN1hY0E3l7t8VjoShw8JeB8ek
80FI7t+MLbguCt0AcMSTdvikL1arRP4kuKQVpeFfTjZlp46TkQw0bANBEIWm7imI
CRwXQ+Rjs/V4PR+zGcu5rm2Yv5Gmm+jJk/HKKb0oKKvcUUqTuSNwmMY9qIWv1Nff
nEaxaTKT7jqBBQD+VuYDgSSEbT+nF2EKl8vR2MtTO6CZuGr6vtW+Fbzknxr4+xpl
L/P1vBEwtEj6bYx2TyMe70VBw4C1WZj7fZ6ZuYOzqFMluNRuJPgZORBqzrO3OJhE
w63tELNVUOG8qagqgd5e/HAB1Gni17U2+yD2Sl4jvcZrwtwcqzwNZoaVDg20DY26
jsVXAweuhdyFLOSstRw91+TjXcNiwK3MSqTR80iVNczTXHUnlupJ1M73c2T7rc7v
JWoS2O/x/ptTy5Uy2Tymq6KDhRhRa8FY5fx3PS7usFbPZr1EG0UfmYw67qy/YG5H
Mqkk5yd7W4MfUMP3Mwtyk7ea4ApY2WitYZdofx7hDmdIJd9trDc4PyG01Uw0Ejeg
I19ex8SmDque2FCvjkZU/P3dXYghX69/Tvyk1r9tqsSrj4TehzZo8OUYvF+gk/AC
/ulqG21naTyfN8gzpq/hIuI1l6v8pDtO44TUTMXw6BEWetXdLlntR8LZC5QUmf/1
FbwYG7gDOfqkyfTWaUjK1GYAhaSWNwYYRpGlYXIU6b9BxuKjyctAzUsbVo1ET7UB
RGX+lef0vmnrtMFVydvX5hTwbUPzq0NoS9kDGsAQLbwVMwUKohI3eVc8iUW3Tzpe
sM6DEA8ROseRKb41dFAbjAUN2Z+jB7GAXCRbcnoa9XwOt5+yupG1FKUWwWJ6N0VU
lA6QW6R8Pk5//3kdRNNfc5W7IXm5aOXUTGkD15ptHQlqHW6GIypKfGJ0lnAeBQ9j
88g1XMIeeA8hNCkItigunVPG0c5LbxjMukEJGxxHtY8SAn6Z029BD6vSIZdIY9R4
hyLXkttVWMdeA6pBKQtK8q9JeM1Md3jIWjceYyL1bshL7xdmEH7qAEzovTSCL/Pi
96MlP8ld8Jq8mNCtpSbgZ5HPWEjrIaHcrhnFoQL9OedhfYWtsz+cvTU/pKutT6th
jvddyBNDRhuqFCw+VdxDNwN0Y5Xy8IH7xFCJJsMShxgg3ZzuDGBCGqcfNfqOQDyf
XpMMu74sZBEn1wGUMli01JDiKW56ZsKbkyg8FE8VDRk33OiF1Rt1IJsmNekdPddK
5+SzPcTtOADlVSBuokR9yf8KU5S6JiiBodIiWJuNBcRgM5cdM8eve5k4CDlEfZd5
ZiRipTuxq/Nn81b/Baf2YL4mPZsraP9Fe/NDiqdE3mNe1ksZgYe3WskCrGtsaJBr
ddlbNtvU4iHiOXaXUqP+uI0FbKYbOHDK6NHdIBr3vrmN4drc4hCeZvqU/FP20EUi
B/MFJaLKlaPZ36pqYyY4wMFSHuYFr9VgOnlI9lg+vQ7+2gNkKvSwTOP4vkk/JfH5
udZDBasUQDF99JJhd2qwC4E6t/ZufQUU+zvmM3drOTNUu3ftahi6q/HXmEBKIKTU
ySuePOCA0X8frS4I0Ry9q90ZDnnyRw959+Mgdcp/VZb2JsEiZRTTWt5RIupyfU6x
erNaYgD+ARTeIRW+onj1TLAcbcaFwoAb2FzixlV/WUq6GcZ30n93MJK6koR8tY6g
Qcpzc29tQQlMgztIMhW50D42x1mrBPNE7a0QpohlhNd6D8pZcYJdpb+w4cU9h+fR
SoWP+Bdf2GCW4HHELaQV2BdW9xvccD4MpoMPzCJOfPK7xBxvUt9HmzcFHM5VzqWE
8Mc6wK9Vk0fO5GFvKB1B6JpOSNL9Vaci0DtqujguRDPigLg7cSe9OLR+DWjK6Haq
BqGxJhu73UnjzKqeJ9gYRgPto7+C5m6QW1CzjTWQxaUpU3NiiOcRfSYcAtGO9yJq
7oNkdhvdX6zu4+0CqATQaXwXiEwgji69VDA/q2HsnTexlZo2XabfYG4OQtk0O+nM
bcc5FpcH4KrQzYMLWrDs/nsrZeT/JOAXd0jcfwYiQzTj5imKL3sLFvImhpsD4L9U
BUGNjqk6R77fy4RtMIrfvm/Dju7WxsIe1oV+LEjYPC8yTg6nB1wv+i/ZfG0wvIsU
Tsl/pm/6IwBK7rWhQSSEVXnQCzfpzkeyKj/mLtuB1j0EO/JjN39rxW8dY/CaMxyS
hdDdZbzwouNCC5mHFx7TY7e19rc6cBZjjeLsIdiBvZ1L8Jp4DcrldkrxNnUcnvna
QGzm/Lltk/UEU3R8JAWSkUBWx+v3xYMKZxH7V0u22jJQKQcTcz5/7kMly3Cb8dIR
UVYHmXqQhhYp/N5nGmY6jtlZypP4BUiCeukslbrBPuWeXkwQqfAJ2DrPSyEgBEJJ
glecRMOb4r/hzV8l/VXOK8yC8yVzN4NCp+2YgINOsPpgdit42MKl1/qW8IfPlzSY
W0UOcGJGxZMnPLPwjXwEFOzFryh7JR7EIC2NBJizHbgXYOO+1HXYPkdPPAWPSJNU
/MWpTLh9n3eSBXtc/4MnKlzOphynE4A22YRuUrccDy4nbkompaNFHOLkZqaVN9xy
Fy9oE3Q5C4VL1nqKyTZyr+JPZ/HB+TgX+VPi1SqLrgUWd2W7MYBa0R2TcX6kVbb9
poVUqO2m3zmCvmd+liXEb+5VkV/X14R8Xh687tKQgve3vBp5lDdJ0isV4EB+tssi
nHS8crYYW2eE3ZMAA3kylvyUhA4pTWi7kjcYAN73SBeO3ytp4GL1VPqb88GFfyMf
nY2tdulTdV18q2FJyGy8ODk9kBo6/B/2V3ZXTg8T9eBLD8028SgB8+mdgJYrZUSs
08yqZy46r6tsN8jRq+2DplMkbhAXgdDoS0YF0rfv07AKD0aEXt45EGv/JKaj1qw4
2k4lzSBWwr5uRpiX3dELJN15oRMGMXi4vg4BbGJtBxIf6K4MoIX/Z1PhB5XXfkTg
rzoutDc4XcY4haswYCkkVVjMsehzoF8Ak3uuzzEOxKr2zNmrj6PcnJ7BAGzXS+8f
5t1Tu/Ba2nNKQRipvoxHJwosO6GF4vCTGNnlarPWuwXacQEHWiUsRiBDE11uQ58f
UgLGXtQ3QCtrTv0Y7y6x+QrqQSf2cEPgxrp7ghvE6ibDKbEzt8Z1XcyOVITJzp/n
TXC91hGffvsZbRrzfoxyjyC0vDbcqGXAZV6b0Nrw499MrKZVemwQmdrFLAaf/1Cc
tjuglgSv268JSuU1dNJtITKtmSreIg+YEu1YXzCftbEbPHXotTnT4RoAnrqEgGns
BNfRjKBulb3f21EhJKqnsHP7MSMJDSSsqcdmBC1gulXDhzRRXa5PBtvGkuEa/KcQ
3I5KTluHUTxCfrToHczcBR3rpatcX7DXXp3shwyRAiYHgXJKLgdHKBxUZ18tEvW2
ouMtgUrwnne4jmvIXfysFDTMNIDlUBIbtxUIweWoIm461tzWQRMKbES/1owftDhF
e50aWJ0S5+OBxIA1GqpEPa1AFEYZZ6e6H5v7omAYrDcQAjLjnE+U1GvF+csCrbyt
Or/eYiO5/ilyb2fR2HRD05S9lY32Djrgh2zapUXrwiGYyicaoN33Mywwj1ujAm6e
7YTbybO1m+GgM8ZceZGyWHKdjU4bPPbsHwQdpAKIAXb6ScwLg/0MJYPgL5QsKwHg
42Ze1FBoB2cMT/wUx3uf4PM1dHLcyLwCkqKN78ZjAW0dnTgkaX5nlPL9rhBmGshx
WcosUW9sWgv7Goq8OuCOl6kjTL/8mBPxMxFZjhxvMFuAYWcJS9KewZZKz2l3zEPr
/UxrFvmPNkQrslTz+U8HMXGh8lIHBAPZ+98p7wzVlKM3iPgMf6hFO+c0COhHUG3E
3EfqwGv8MRlhzu5BYaImtlzagpdlOWxdS9F5uzEGBPBd8vJiynGvh0lRIprJxkxx
1Ukre0Wxdm2SfdEZR+9HwS/CZSaDtwJuNvraRIWHp0Dsb6HNrk3Fqf9+tx0HFB2f
7PFSxwLGUN6C8atD6lidXRl7qrADPj45CWoOoMOmXBZaVv6peTIBp6Ag10pAZUec
JJGO4xpumjkNeZW4PM9erkcDm4PLJ9T5qkWlE0MZQUANTa4K1RnQ5bIVtEZpbx87
dUdQdDA1JcajSuV9hbcRyGUxExPGgH5eck5fs4RNf1fP7gjoG9Aq/50Y8+L5tceV
KcbZ716UEvcU+il0LR0DaJXmVXF2/F/fx4StucA+pkYk1aRjn1HtWY0S6UjPf3BM
6UIDb6o04TjF2urrc/G6YkZ6pgyoI46i17WUjA1hShJv0h6PDDhmo1hq3H6dUex1
7frL7syFq6uCu1G+FPzA3G+hAvjD4v2VXe7+dIOox0fWlhzvD8moyp+OaA0RhEiu
B6807RWL/4mdaQV9Dt0WJu8dmu7Rv95QcHSnbCTXvfAIEQ+rUTUzEaRybxF8+kqC
dtcB/nhLAEwKIke3QRkt+C+wDg4e1fCG2GIExcswIu8a4/hm8tV/Ak4dn9S5u1r9
QZrX2SFoIUpsezoSXimLa8JU1dZtZEN9bNDgn4kq/qqbsXjWblT1R8Z7oeXG4VC7
0aXXBOPRn8xXdeFYaXuZJkDActcz3bsP55bCwwUDJL8O1hm4d3qUuvEhCqJFNw0W
gLAeSqUSnSXd3JGPWbMU1FRUFYETcYyScwwK0GIISgQIboyB/4kV2x0dprkXPYYE
siOg6UjuEkVMRofS5Xg11Wu+PuWMKrkN3BUlqT8EPwXH2CLf2OhqRLiMTPEytnwS
ATZagJEOgpBtnsN7Ul8kb52+B23wjlpgtFgI/8w8VaPmL7EGHPdMUDvkIKZ3Jxmd
4lLVGwhJhb3F89mrXQOXFNSh5nSC6LPwn8MmEDlPtvcxvILbkVbDkSfFz8cUcp1P
uL9KEVtYbdrFLEGzoGYQw39oSPTYnlZ+TjpsN3kuGljbHenKNHio/LsWq0Bg2cL/
t67Y4oSoXjkjmtUD7Y9aBbfCvo7VP7hV7+DZMIsXcUTpbkckOyZX5U6CPVlnP54N
WX0AhLLipwkavvtS6XUVfkSMaAvuYflYK4qGhLTbCh/wxFhrScazYZaXk5FKWADI
pwDJwKr1WOK/o0PAd+QHVWgJkfZ2LQup7D3+xZyF+VWxvN73+32Ty3AL6aYEY4G2
/+g3QIujSI/3SSwOo99ZHbHz5VgQ3tU4io2ZJJ0XhhZ3s6GoImTTCPkluqgqbtZp
Zgq8NJ2FibzyIK5IfvYNRb+7NJ9Qd4op5Mx+enliiHuhszpgELbboYCC9buta3Jb
WQGH3o6S79nC0JRio+KLN8jtdiQi3y5r9yIN0+BFNvKSag98eeJgib4PbyU9o2J0
5btnSYsQllwms6X2lGLKpvPofql6MeeegK44wHJjalz4vnS17jd7kFxbMJQDs7GT
fCW/5ldRybR+nd+XiS+UkxcCcVBw6V6+cGYcAEIu4ll/tBPid/6aaVKVF8fC+XNe
0pSDwdI77RBYCxWYo0vknXminB9aBc9+o0/b+RJs2cs3APq9twiRgI6MUMLfAu4/
GWO9srfyZwCjcS27k2nlmxXUoDOdjwJHoP0wWyON7qyO5JuD6B8ZiGY5TbeFfAPv
O670WK+pW99NLvgWg+N2xhLlGLR27VdHKrZDwpio7yN4HwEruxnawPCPGpBWak+Z
PPOrIVfm+TMfmLSWZctbMVkIN/B3IVdX4nwg/Wla9iWuW32DwHCpaTmiO+172ZMz
wSGWzuuy0R96AO5jejHN92eEW5P7xmGYpnMc0y7DZjsowh0wsCLMgSkk0H+1/pc5
UxrWDosdiarxX90iQZJ/rjbOGXuSlmfmzpfJQI0pWDFS/iWdmK+mB9Znzk9jB7oa
AXkMZL2rTYVE/90J2nTVoR/2Rr4A1DvdtF1TZqhsJhyFROfFPMLQdumuxBbV0FfI
oTfrPdZ3ej1ZjuLQkEv1rbxabJ+LY2jNqBur2I6obE2clOR6hObrQ9GflK2oAA+O
PkQPOATNyvNyjcWMXacjtNEkd6u1/q3KHJB82bgn4BueCYV+gD0aadRAwgOQ+DHT
o1YBvKUIra5firRMkNDogpolvexpxTk3Ih3DFX4jER4bzLZyVYZNEHKLM+0AqI5Y
UtjX4tK+D3ah8kz18Ysob3Fw0Tz2c3CDD8sGyAxW2E6BB0Y2qsdPVSn8239AHo1d
j2gE1bzcbe4F0FO6vP8WPShCYzkdzSgLmWcIAB5DevQ+O6bVJabxE5dXFd/ONbIm
B7PhBqTAHBjagZ1H9Pzpy9yqfjmJJFrGUwSObDFCHfjI3+dQbaIK0jU61ZiHVDBH
gQLGemdnMYLdCQBM1laUc9bFOnzOr5aaDuAhUFe4Iao/qW6kolOeGOLCOtGqXNmI
5xt/sr4wF8u9C3jDCNPTDT88Ah88Jn9cPY4ODjp1AluaKmH2jXp6LzzIYq/pQRLH
XrcIRvntCEyGNmx1inD39NewB3Lv3X6S7meF/c0qFhlyvIN8QJmz2BKOOmzKqTEh
q6rXGACIE0xOkii02n635TRB31RolmxdTAgVXODnYEnLpgBYBsn6Z8ljyWqjTNXH
+dcZaxxh8pPxHhSwWlMn9yNL/ppZ3AYcfQXI2qdXlQdVFZ/vcLw3cVEO4gxyMLc1
l1Pn/pNQshw3vciQr3KuXN4DP9UaQ8Ye/DMCeaNrKawbURXKj5ObMTU3sb18sSCS
0itqH0dm7RQ3HUzYjiDLqvL8pjU5Vr6v/3iZCDVNHcE1ckUXYR3k3WZSDQdO+AVH
MA3lBOJgDmbALD/JZLgcnVocnAN8BXJF311vmENrvYZPy4qIjYsqI6ibHV/KCYMp
xKcpXxH9am9AameePUQ1/XfNtP+6RHx9N8+Ajmuvo34fHsNOhdx1XgnOfuKGBlpY
1tzFdc9ImU8R1hT8+OPOqK5z/CwYaZ0PAuhi1d9P8IvAICCArIjOBJunh5lJ1Djr
qcXyEbEKEvBcueBbP+u90+pu72Tqu5RjiRKTJnETl/xaTBWOZ46oP8t7QXWk3u6Z
TnOoXasXcL8EOSLR93zK+9DZLVd7LPiGXuylV5GUO/DmqQ1eZBJ9S3qqVpiYlEDR
MxfKXsXoNVvhTrAm3cx/j1jx+TJBBeMLkYcKUNamx1BwMUoaxSOXrSLTWCQGaVde
JOb2LQVJGqQbTn5oZOE8Qou7V6jntRM6LP/RG1UxnrllyMtZw4xRhsHf3MZzX9Kb
yu5oeHxkH4hwS4M19nOW2ThzHffYPY6Hqa09ze2fqc5EkZhdMnLeyYUBJLUAWI6Y
HXUDg8uP1IBICcRQTANKhjNipUjT2mkH8bXkgTXOhETtQSGK5+qoJBPB+jbxjpDm
K/Ta9HElna/jQ69zaGzdrrdZ9M7kH4wjyDD72DAMmN7xp9Xod7M0jMpKo2sTdbdX
ux4tgw10SZTkzpZ91BU5xklRkgcx1r80nLGT0qJwaULnJx+fpwTwl+1kmAdsHgBM
+px1vucOa4ao6AzAbjzf+trR7UyBw8lDjQH4MVyx4043oqlIDhkLUsbmGMOXuh85
s93J4yof+SkGN++EjHEfXZqYW0Wqq6TwnLAbgHpPdPAXhayoanD8jf0TGm3L7EX7
1kWGd53CDYuoTQm+0Z0558v+IfFhEWO7BzlNuIVzmtnBRrUWAn5KfNcmvpfWMmz8
TOBW2lZfS2gxiy7qwHvMKrqVwh6JX5bXUFWRL98ZEjdmDUxsczJYk0wI1Xt4dg/e
UOtL3M5cxRD0haTJBlmRo4+9B5JgE8rt4Vifj6ADlK9dgPahoxaAZa6MzmfY8ReF
EOjBIq8esZYh5rVbbNSMqzTmfPodNqV6/71JVOg4Do336m0Dck8MczgFTFkk9CKe
JWETriDRSf0u8L1Qg2ccxYq6dYP08ZCTRN6n8zZxwjA9RXhPS/DpsSMP0R8lc67r
XR+TiPM6A/XnkR8eY5NIIdyIWKrMYbx0YCRIQZV9igTU0FUpAydAyWjyv5W7Ze5L
ztvKD0YAIPn4NO6mTarGldJ8yB0MRy6Bw33WCez0SHHNiSl66xle3SSMDSfTTazr
KIOPtlpNKEumNu+zcFwBoqSOBUiyL37OwknMyTQ4QwYBaR1B6fakmhXj+xfoqmTt
KSwrI9vPfKh0cC75Mpioq8DNQLdcdYy/vU13EBL/moS7uHeIQJdZdlRMSKYTaaLF
klAtDVVL+E//Nbg0szWcX1tcRtD7XQtEvw5pa88YPkSPj0rRMBl+sEwdmfxbHSE2
KFxsx1KIgbmFZ94pKEnA++tX4Mir/59VQj/ukZix/vpvL6ogSIAEPviAAQjH255P
MAAgUlc6+32zA1ct560mrnuEl+zxzHk1StPIJo8KB/vejE/hO5VU21iOT8FwZfki
V0oOAVwrwDFSbboevRYGr4/Blf8qK0ShE8ojmksuQolnq52LDjXUDapdPZyG/H+P
l+ODi7Eh3Kz2+vZVSLL421uMaJ75Gsc8hxw+F9oZP3jtKySliddLChGhiqAfAt2t
nNVnuji9mJ3KGI9jJ68nDBTfPeM5AubBNkgOcFsMqnUQUps8epkfNitbUEeHBAST
8g8apHQhiJnNANkhaUYtHG9L8uO0znxbJnwNtXtAX1dtSiAY8FHiIaFtXaDfNSWW
VldHmOMpDSifPP6FQLL7I3YVod2Ui+5D+StZbEoHqXJG12+RAwnBOZSFDDnPz8kI
2FVqNDzBhl46vtLONpk7tlizpCepk2bG3wbn8TblIS1M2uoTFP9zowbs18odg6Ln
ArOheJoOXj70VWIhCk91u2/yyx/Wdm93kAqNItNa18rSAPn0/wrXQE6m09RQGdse
rkzcwi/dNrFMrAvchJxFb19tzlwOTbE5+JQyXhmXE7I5NX8quNe4VlsKP10kF0ZG
5WJ2ixDJN8rj9AqhqdMEIYV80BFJvkVs19hmSCtvHoUwqvUSl93UIFJvAW7uUdc4
jk8WJhqORifwUXTku1Jhq//bpa/lSRb1LhX5s5ApSkf6u12wuqTI6gQ4wdFnSYuX
3j2ySQiNYOmwaatbLijfM1V+SfrHw1R5bmsZvfaIGlpy1BFHQHSokLKXcR4pEXZJ
fQg77X0yVwTMpbSXIYiOYMsEcmELljENlSkdK0O+U8q05HeAStj37aLBYY9SUJUR
lgjb/cfZi+2LTavsdg1t7X4WLtLy9vXgNWZejWwU81mpia7KEAhRkknVb8JLeb5T
Mwmfu+8DpbWrnOMuBZ/iAefuv5meZZTkeN7uzIRC9OjVIi/Geq726dR90O82g9vd
fYup9j25dwTvAPGFSFn+OaNETqOBqoK7ex4ZMiruZDFUVHOsz2O39PJABEI9v1CU
IkGHQmzmHqhh6VysujzKc6o8bvqK+/Ixf56D/9WJl3pqCgJbdK3Wb49b8l41tljE
8vBS8/CzeIuNZ8aEYdjhBeXKNP/sHjYsu4E7B+7ASfXkYGRHyMoLEZYzVHLHrQNH
+Kw0IJy1e9xTvllVHiZaoOu72hd3sQx7UDUI6HuVg02ZcBZl8vGVGefQ2+zAG1YM
9oV4sJjhbm5zmg9e1XKyHLW5PYjViVEXh3WLsaUfYaduJel5MWg4+2wCeYgyQPoM
JmZ7azfOC8l9aAlDe/tbm9V5QNguHmSFpo3y+6LnliMc1tejtdSjuc3fxv1WGs7D
Ipx7S20/DrrROfQVTNHpkxssi3lOphP2ndDJTD1tCt1ZXmIr+yH+lPaXZV3jcyiQ
WVRborOJmlAIuAd7OZwiinyv9LrGp3/r4jtHwli3qsEWrmJGICaYUN1b8PZOGpaF
oD2af7V93ScYPZDPG5pW5CRNqMNKQ0Z3pbTp1tTeiFc6w3dH+bid6wsEFKWZwSJs
9TEOVMkRYHH9bd56hjpAaRWE6UUYmolVsZB8XLgtEFgnz9sAmKdB6sLeAgwYjUUy
zDreTvbx1S1soTVb9sKDAovNlOrYT9GgqPMgGFxdOlJ3iyXWjdqdO/boR8QJgL6e
wIRGZADhjoq62IAwdD4V7nvU4uokjdzJ7Iy2ZQjahzkM184lK/kS9S/1+FAAE2NX
2veZ+An7nQKCl8131HanthlVd6hf5J1QnfOUqVMC6gZN+zOYK0lsa2z6punN4NWz
4yYsFLniF7iMmDkHPKnk+znfpFGhr/aPap26bCtrBJBNRlS+fm1dD9AxlknIU3Zp
NPuKTs+K+tHCNRBBCFJQMsG9oXferq1m030feJLPX7E62X3eATdaWl8avlwK64k6
nUf7d0qJmoLc9BAjK70KOQWb9U/l3Na77GZqHBnKmWcDOUpIMTtS2HSP+AU6dh/s
jiIyrG6iFSYwxhIFljUqBAB+7IHctza4vpGHEnqMeIWzoYfRYHACa3+liAQFL8Jt
lYBRWRF3hHpMELu195aUV8zJ2Q5Z6UEX0fA0ucgNTRxAvjMjZ9a1sErF/m+w2gJC
1FewXQET6A+7JL1kGXTKmAYMEmdHozWGWq/XZeZgLjRgS2ZGJ1yPsyNuhe76udZD
VR2QNOFBKQNFipXsKnDZy9D4CMQyzzzGHxDEJI2pvjJNK5xPji6Lr/9XkQRd62ve
BUXP4w6HXvyRrcC8rJ0WR1B/JoNFxJGeOfjjqACDP6zw2RPqbaTujXoEBkw7zn5k
ot9PvYK1ETS0HgSxefFWz1B7QnOH3gxKZh83qzAsHl46W/QDwU3W06toTPq30qYI
yiYcQIpRaUTbw9jRNEEK48Dr4K/tFy8rtUrE4BvtghpGjc2uTiGV3hDxq5Tp3xyY
la4xPR8aAF5ZHzp8Gg8GXXzXuHHPkHVW5dwLEnmYgHFLO4DOR97wJokKGBOCaSGq
tAZLsXk8k6XmjYhECUzLIc5L1KDK8woE9MJBUyKFNaBvcH0IPYk0lhyjBL7YjSQ9
TiOV9w4yJiEw4KebQZPJKNld3quCEpVS/fKmydabWr1RnHJnBXkFjzBZP7mdKj0V
xVWb9BSURchRvA0FZ2k1gDKT4rxu1mSvWMZ7NWOVeFi1DUrL1OvElPff3CqyzA7u
nNujF7uxbdF8+Am2sZEqri4LLK167QPZkMny3fvKdEmHvbCALfm9rydRmEaDjpiB
rS3Wp8fe6PJQXNdOjr4Ydhv9KwaRJqWdT35xenTGfG/VmmPIKGxxHpO5YiPXqZSg
Zw2jYBbk7yfHdSTw4Wceifw87FNpxFiOsQwtYpBDkI7uhkmx02Ebwt25oNpdsgXS
hhjvjgmcOp0IUbNfVJxA/rTSynX3+WraW5y7SUKD0IS9+XJLdU3KcSJtGWnyIrTY
oI58yxh+hZQQCLfMLou68cJ1JblPGOa0OkprF5flfqrvnPFnmjzusqMAMRmPFBZb
9oh0ym3NGLFS5Q/fAT2y9pvRb6XQfvuVtPrEpNGPpfQy/wRuOpNYBGO6JXX/5CDV
YEspM4JvW18zAyX0veFtlSUSYKGZdWMRo6ZKZRH4vtcDovoswAYOlnDLyD1OrjUi
7Uo1K77l5sKjEWs6kbkwoY7kjAZcVmTyt0z1aqRxkDC93SXrH3sd0obu16iFvOJF
st0fyZl+TpMCRf4NvIXvlBEMSgxajrxcCrMti7kvFmPBAwoa/lU3RZetgUI9kQIH
T0qnjDUQ5uZUUQ40WsFe6UmImyIwp0liGepvDxu9J8ib5Uhc3tLI9oQ9VfI5/kJh
pDppnkQdN6qKiDgH7G/nnc/Vucza5TS3HtENQ3ext/EheGOR3x5sJFLG/ii97uDw
4Apf7PvAiayIT46SI8xYaRRbIHQz7uxR5eAx1pQDwvDICp5XxuCy/KoAQFQXGEjd
jMXQ5U42k4RwluviLJxgHy6Hx/JIYwLAQ7IxxURaZAkNQLLXuYYjQrq9LM3awTOw
KiDvyLvoQsfQZfBH9PKdR3S36S+vIQ2viH57maPiAk8iQeVMSepkw2lBF/ZJWuCN
bscM9AixRYLFo/ChPhUnN8Ugq4DijP5M2C4oW56mQjR1i+Su0B69JMjkYvpCRIY2
R3PU9fTy9Ae/LdiiLfQwkgMMkHA0hTD+V7Ybgb3M69uRzUJu8reVqKqiUgd5+WK3
9qQfthbDOuPvFX32b0SnOwY0c6KC4qebSOo9PXk3vOT8VF9dNRecAuuDLxnV+NEc
f1+U0DhiFBuM85Y2VrHb3pGj2sAjxf5eXDfm8oIuCqLFFRW+bu4WBC9c+QxXuIOM
j3xhZ4qjZ2UPu6Q715OiGmO9R59REql0kdWQecMxFT5MKTlyAlDpVHfKW4DDrdwB
i9J5c+Pe90znXnbjZGjxcyifw3qfSo3Yn/KUfpNsGTR72pEHQzNGt0P6JxrT6vgr
JFxvNBSPO++tsvimbHZFCHiW9jXezI3C5UsS2Ea8Orv4EYVrKzzhiwMMBqcDgAhv
xHE9f30YibBGM63oQIGiSRy9yv/6P9zDJ1GUHD+vdJtrq0rC4CnwfcUcGl5L/0xG
ovnYfqRR9i88DyBvILUaoJHTQoJZxy7p+oiq+wdRIRMAzd9YDOMZYEtcOj6u0mLD
8yR1xAeLY7iNohA5JukThJKeYWt0oT2HHLPdL32ROHjS+lmh2B0HoSdHQwwBEHbW
CeXmYuRMfT1AhXtqGXhuvWjPTUO7N0BgiI0Mct1HzPegojD8Hv1bRi/mykrew84c
DqZTtHk09gv7Q8L6nOZv3kGlDpW1VchUjRUqMy1Q71Xkdxnr8n/1Ty8har0hWcC4
gOuf92KIv6Fbjsq89yh7QsY7JMENaJaDd8Md5mmgoDst9s46G85gnd5XkTSy41UY
cVH6oyetDdMfxdMRpkUPfzyArb4TR2oIpUhubFUMQhMFmyGQ3ZyDyJKcZT7Nt7eQ
fsAAwE8/cYj0SPXN0LykWhT/BEk5COKiRDRWdn8H9aE4npG5FDv8j3BVzWipPA5G
lYMUlDuD94qbvy9m8IjUIxxoXqE3SgFo6HfQV9c5NwLkCDj9KqLREnxdR6Ehyc+4
fcgNSLcirlhuYYZERo2bWRa8tGurhLeyHJRyUJ1MHgBp5ypulx8JYamR6sxPidC2
KjjGNZu8AWR+4VUlscWlek+a9ljyIAXnG2Mm4x5osg7NyLFNPbr1rjXUKjvAOlBS
BAjGm5TMhfiGN6YFvb9wJsgu18qq2xyMC2GNTzbTwXmsM5wudiitqr86Mq5kGA4W
Fmd43q6rS2u0sVx0tAp0Y5Hsckx+oGkFtr5FMTqYXU9BzB/T5MOQpjOtwXmYaLLt
qDsiYRkpmEFCS9rWqu6lvsWWYtB5tJ3XO5/mAnWyeUQiLm7t4+0n7Q/GorkjmYEZ
4ae+G0MYJzwP5M+QjMrJjk6y8v9Rpzv0c9be1wO36wiOuG49k0NHSD53fonPJJ44
hhynAamtW65wC03yQ2JyplYt3IAN7yBU3tEjNatxovxmpSwu56nIjgh5+UXELzGB
wT5zRMLWRBK62mCE27W7c/hw2NJgW2xPGxvR7hjO0mAE/Rq9nv7jGr+UX2vMyYdH
5vijHNngoFw2kv5gScJyi9t1zmkmAyevken0pcuMKWX7kjwRGp1Wpo9s70Cj2DtQ
VHVqcplxgiejkz2sUq18BSM/StZCiFJfPQMWW+CXZPaBxtg9N2dTMkeWaXRExksq
PsexVSBZY9UCmnrO8gWYxbKFobUnTvsn0mqpnqADDFrMXRoLMsqcgxfJ+5uvyWIL
6e+qu9vP2gjMNstGoVLqUUu20nMFguK2vdDewXL3YTnHH+96H/svGJATx7jQ5F3n
uEuMSIT3n/3EDHXewNKjQjqs1wg5itpdIDXJurSJWrWgK7yzVtrWvv514d9x973g
qabxEPTT5956KT6s7Jk1xqngRRm1gKzcPMiQ38K/BpGR124b5ms4AAn+9R2FfE7x
G7ZThT8pz1Dj3lFK9yvDEwJzdr2yL7+uE99EFHCGo1SPHWXC8hQS97zxQyMEsXpi
d9mEl/2CwjoUDvsl39ZC9A994X+lNynUlSuFDziZA/KNdhSIQJz/5gPKCIf+9OZb
impueknwUZS1sXVTi2jv8In3Y2ISBKxFPC3vFLUMki5Izrr0pn5S/yiujcuu8rZJ
/EkoaKZCAaL+3wqC79AcAxuKa2YTM37sehp2Fygb2vnQApISP5A+nKJI2rl7/QBa
EV69EpLYrNO4Du/245t3rcs7FTXSxXnYc40NyF94s4Y1PkyP87mLwIuonaLXWrdh
x7SeRZXu73l1rrO8pSBR2ytCK+QuYWWBd2woNd4g1RcCqsnl/Wv35HqeZeuXPp4W
zFxvvAyZ07m5m1JwLzjIFBS4vDeXt5bhZb91/1zOxy9+7oaWv9Vi1L2lGkDJHto4
ec3Zr0Ep6k5YzNMm6UbJTnRaNgcfzBCUSw/WJLclLtN5sSjGR8mKuilby5QviSZs
fdtlW6rCt9pm0uLUP7IczRKDaDuph7dDg8MpNciLJDeHJBI8AyIFgazWgY2BFlH+
8qfOsGEpPVAhKhEGiRPlH12J+VNDErUZMRsES0jWD+7bNbD7ROM7Ep6IM1/9MKm8
zGJF/i+CKW9g7IFp+jDa+FBxdmrD1BSAEXXL+cRwKw/jWhB3VG4kg3bOWVelyzMH
Iw5+4tcoUzah5HGQv9iL10s7iXLvorlDM5St+a3kj0QgVbXFmItc4WJ5iMxj6bm6
Me8xgkqphqsosglrrH3WhJkIpQ+e92xvp8YR0mUDFwHspVvJg6YibyLeQ8XbjEFj
AAq35ACH3QxFsJRGt79Huqiikv4tleXhU3hfYEG/J1cSV3Z3pRr8RLX965afP+iu
Ma+lmo0/DNugGFYF1z/HH9lMk9DcDQxYpW3sbSCQXDV6r7AfulwCz/iIvFpl0KeJ
QMY+gj7v/kQkAawF50+0J1FZjEGEUvoW4Xv0d6f+dJszSQ5qiFOGkPRc5kDUOFVV
Ir+BeSFlTmmqcjeujE367oWrLHUXg17BBkhJh+Fk4EqFb5X0z0JbEhWus9wZbPxl
XnwDfvtMVf6EudjqoGcn2T65XPDyFxG2axZ2UxLI3M2/5q2YpOsEg8y0ml2lPYSA
xZE99luNBbT5kSuuDIigx/ybgbVCnKIMJE6kbAXDFBQ+qn2s3yGEf2H4lNpnXOvV
58Ue4Pz6qeh7jYhNZOo7a8d2tWwDwWXo+pAEp3Fu2FZiDsK9ucVgSjYS1CYj2Wte
apNYtRFylqEmHCqXoM1/3QpBl5ZVDF9Mgf3xo/hvX5PFO60U2EbXLZri3EjKTWEg
g9DpGId3pi59kNc1dT7bNkhZu+QdnMTJch9RAR0zduPGL+7agv1uP3vwe/UQrZsF
0xPgrvZLffLCtYWQJIpjSLkZnLTUW3I608EMNvz7OH6YAs2Qav3KDs0Bz/yLvEMH
ygFbV5qyrWfbtAIumcOcCrXWDMPx8Sn+AiuJrUFvIQ3l/ZaoHu7Zkqob+haVMih3
HfX9XcLU2AcEHxkpDtp5j5MM6sadTFIr1QJc0NzHBksl1JVkeqZ3aoh1TqcPXFs+
QmiaBzIjBQ7MKRMmgdA31rMLq8yVJcOCV+7bOBShZAANQuqD3XBKeBcaf6a5qh7+
QVQWZwl9Qb6bTghpAJlgJT0S1b6gbz5hC7iXPEazoqs6KtJXgZmb5Z7vXnl6RdZS
YnxEO8F42NoYE1P3V4EApycRX4Rr5GVuXVsg8ic8Gk7C+6O9oMnkyBNl8rgd4OG4
nvNuyIwZdpuXnTJyOL7Zr/K8pxuUh3gbnd5DdBZ5OWlS5eVRGfy1wm3MHuNLVHVl
BxmKhUkh/Xcvr3Aaha9bRW+siGWfxgZxMP/PWwBX18Lt5yv/kC260Op6Ib//g9jC
qp2ECvQB9k8GvrBNay5IqzWWsWgbQ3mukYJUhnWxxlOLWO5XR7UV58CWCzW8WCfd
MXFEAxFURKUCCQJkG26Os/HG79RzMFLQSyy83VdXgjZZoxDEaKBLLGQQKjplrCp0
7XgIe09ohrp28Jwmupa1T/YnzfCg94cALk7c3IYOr4BwSOaID/ijnOrtRIjNO69J
TLEE5diVEwWLT/PtvP8CEKnAFuKWOYBGxQSxLJAY51zqMs0BuvfqMVI9jiABJ3fB
PEVN3IZ/eKfxtI4hl0TE6MHQsC4k9vEh1syR0Ja5oaPkawWBG7YjOepKampT3Bda
g+5AyVT3wm/9j9NlPJv1rzlNSyI6d+hIi8xwKb0IFIWx7rPAJHx9UhXJAe1i6ivF
MCh3f9zQ6XZJ5KCEAr8NfchG5BmGcvdAFwwKBxDGP50OYRuAN91YiuNXtlQOfkvr
I4u90SS+CaJkz8AurRj8bV6SflEqkiZpbm7tT1Ix+JsOJpY9vO3mH0v/pgFRsEbz
GaalJ/uzflPubxFaT0USQd8LTIlCm8zkECvNjHg1zY7a4GFjiswMKXdu/A5ZjMIq
f+P/EWJuYRi3JxHIh1IHZnvoNw5lpqFqtL+YFx8xZQ8rk5c2bYOUKoEDF1aQOs99
MY4gG91dXtxZAOvF/UQ/QlICwLT65eY6QMCNd8elKf2qhkDRe1ptZrXr0kcvvX/L
5j58qWYALtkbnDVhHOxajevFNrVxuiM5iInhq7a2q8M4yDzbpOoi3MGjUJUBYKuO
qlNvUZYuox8fJHfy0fU6J08CRID4ZtRgD2MXOct07WcLsOQldEgXVtrjkSZxpak7
VDsJp3H3MbFntABlNA45y7y01XDWZwQ5IPa9cvILsJODIepckkAkLacQSREFh902
SOY7iWUDYp5a0oy2wEPNCvwFWBun68RDS3PmYUTj9166GELgxijeoHVlYJpLpLul
npFz8gdHuU9xA0UHvCm0Ix24o673dwpaOO+xxNXYJeSqHOheUIO4/9b+nMV0CWAX
WqCd8+XSi293OrHdRGKyXa1ch6fkBK9BcNzEi6XF+5PGGVRhXU7AYh01keqDFJu1
5xBAPm8/5b14ZgKeAwCYAJ8yH2C1Qgbmxwq3CSuuUxX+b7D4hE8ExZ5HWZ6v9SBH
gRh7DYutToDvwIwm5OLbCYmiuZJT5l4sHZP8dKMFWgjdINqXWQ6TtCwpHA9Deo6F
7v6m0/DVbbT6RREGVtTv8LdRXf03qMCf8rtUCvxVE0t0RMUCMfrolec2DZvwACNP
juk0aU04jVgnTQSiPteSGIcujgYqONhiEHCchumBKlpBkLvpt9WikCsYKDEj0jiA
V883lftCHfRPRm6Gj1TbNc7fhG7cz8bb+X1VxM1AX5vl2RD0yLxIF6JiDwP84PB1
9kdTtqEHM2PQvCYJDmOP3Hz7/gAZIl2mSmiiYAqoHtQ4ctmXZsVRus3QyNIMikwo
gEAWncOBotZNVEHPvD+NbILeH5aBCY3L/eyVgaOfa/O25dbTblpe9/SUu5lFccx9
BSyJQBFVOhoUTsKGarAlCSc4Clgw9JY7t9490zodL9jc4aM4aQrAH5DYTUZ9EtVn
8LhFS3DUxObybG1LeDy3zNG+0O7Gi69lBhGwkgafWriJYAIcXich0bjGW4PvL9N8
JekIvRPr6Oc4TNXX5G4ABO2d2S5BKGU4qDpdLGG8O0QQ1h7KOGUdVAoHZJ96Vr2c
ciU6EtGtCTKgW9e4J3W2ozN1zh7B+bN0n17ouVRMkCGAVbMdtDaPLBhYVy9ZcoTq
5YyAX8FywUsQRXiN5wUkMlvZ5tHVOr+TfPcg2m+tqfyNpnDkWRHsL58CXD3nrLme
ubmeBtdZ/vzikpvqVMM7yH/KneqoUoH50fnmdubFZ86sJze1i4P1vLDK+w/IsUoJ
IGAmvviIwWfJqm92lx2HkZxPxnurYcsobbVz8MGJcUtjCPE08k0VB8KArCTjHzk2
WV2CfLMPfP5tJy5djzaFW5ZHPD+7FGeriCOqYwSHfu6TKUEeZCAhDwRHsMA+58KQ
gfxJiaw4L3Azm+zLGef66JyVhIyGZ4whAJVftQrKINvh01m0qH9/Wfu1yLaNZcKw
PGmulTe6c4Vya3gzC5EDwvZQGhdbB8sgRItLxMX1H86q+nVaELwo5yB4Tg1QQ8Qp
Rrrj48mb9gewD/aiuTbaSL7naa9u4jO7gL6qTy/Qg7A+uCfdOd50zjkePQaiUn2c
zlxT/Di0fRY5LpISkayZ2dADGy2Nd1D170b9gcmuIeH9vt5lPLob6Vxw8BeIip47
RGAEgMP619DbtVPlornpppQGCu9yqilEu8EP2fT8bUC/PBwNmYedUUzjfAexY2Ey
A78wuwJJ3eJY9KrZmPovBlqIQGlrQhquAo161FHsL/j8rvdN1/1NBA+yh+gqt7DT
Zg7pJV8RAk84OsK9OMOuEdI1KV6GLAePpXs1Pp0GcWloqne2JowqhssPXJ2uL6iP
fDzFhhH9fR8Dc1/hetgTjw8YU60yUAWl6bVHAfzyULFrm8RjJLXA5gq62TBtV/P9
EqPC3EwNcHG0BzpEvQCcFUwkRpi1nvP9B/NVYhYXp4OkjbL7tO629it7tb8NCWeN
E9LWbiC3eGC40JN3GidO8g7hpoXd/Nae05FRJduryloulfxFpy4HvRGN+aIJeyFl
3+HTrKRlyMgdptZXb/eBejYAcVWGhteyW41z4CDOa5KGQOYXVCMyFUgBghh36R+o
bkeyXG3q4BYyFMcGvwCsHzPr8orcCi7v4G0T8yuqWuRPjnsiB/hH8j/4rB+UsaYH
doxbakXXmbAk+2pZ0D1V8XafXd/KsOsgX/9h2LZOTkpLZRe7+gAn9JQmApRtujYZ
4ISPFK+mWQE6Am50iHMVJucLoN5W9Z9LWXV0ix97ieUpyQlXTqWUkl+NxvppzNNv
dXjcRlgnYSRpqsyYTiaSdlKi/PJbqZp2CC26C61B5M/QCTV+9GY8wnA13NB4CvDg
zq1Ksbr91v7hfybQkh7q+0hWf30vPpDR90JYdEgB6+Jc0PAIMcpO8VgBNYCoLctn
6JpaJsdENx4u3JyRiPGoje6eJS7hs3K2G7zvePAYcDrpTs6svAuTOEECdNRMs/zk
mKXErcU43y4yVYRvtGPd5fiEYFq4qG7VWyiMz5to5wF5kcmhhcK65ol6dJuD6Tli
RI+icxvOiz56TGqtrX0i2K533FHhjvZpxr6bnajs0ZDOVU0o6CF/Qd/EBblirt/9
ooSX1pKwJ8DUzkrJIoPE9LaNdpCBsrN4M1AHOtL2Ag/p6BI19S6mJVsP13j9rUJO
dmbETdFYrkQX35D49JkhgudHSbgYXZUXtxCBkBNy9ZveNlQEIfF7F0S0TgtVVO45
Vd3VougqfTljkZplh79XZU8A1Y/4Fi87w/oKg7gMqaw8NBdwJozDVuBU5OTTaNnP
EUcG6IVebj9+CoY1ZjV/tJXcokgds458uw3mbxeRklaTVUhjj/XTG4gzZLjpLBBb
76JJX6U2tnnn5SV7wVOnMElpYM0LFo8CS6OpvZ3xdFqo7GWUf2QqLlSj3uPlUFHO
JF/savT0z4AgQpOLoc7gQ0ay/pH4kXLyw2BrMSCUO/T8GZcOdeuenmEY3bLw1cTA
0lhSikcgbeRQU/e2PxSYRVf+byAHA2TLibm2AcE/pWjGdU2RpngbjxU1BtO/d048
kkC+fTEH4Fqf2Rl3QLmG75rd6Sp8oI955ranF09dWSXHpxiLMNBCWmWsoWf+9Mnr
XlsuVbTtHA8olgJMKKrmvX+3SWyJd5xdFICaN99O3b2C/9stZjG50htz5tv0JtM6
Qz4v8+8hxInIroeLSKEtelKG8ivrp9ySUfngt37PWQCHwNJrBcaZkRyFaw1ZroIt
jDnamRP7PGm+En3s9rYHEtJn6DtisqDdXcLZDtik0cHwW3pSmzDtv9ivG3y5OG+R
PQh5WpU3c2PhI7hs233Ir0RBxxUxk+QZgzWxrE9/v0Lh2IB19EFYAKOM9HsTJdnc
zpMwk+7YKQ3xPHphpyDqUCTa3aTtp59/1tF/Qqom/WxUBt/iL4/HemPmqGPx1e14
ZusdGAFiCf2MEIsR190bd1RVZMdcgbuwqSgRbOKE9jH39/dMsSYGewhlX3seaZe8
F34Ezt8aE1li4nLhaSgrS8c3rfS3W6ayj6O6ykpCdBUUTPIpUwUlEtpXtgOotCQ+
r+WuFi4dNx+Fx3lvkdxS7XtSO8wwPyDTclnx89xZHTvmO08mRaFP/Agcw+N2sunH
syEaQ2EFn81qRFLwvzDEIbchSEiJNuBnDLVPzB9tDHEHr1Y5zPKlBJI4JoL3XUot
3hkQ0PcEvEZCQsdi6cS7L/Hx+bjR48deo7htDAeP8hRFbDwD+pp3jw5GKo1ySA0J
5gL63LOQ1ongTx9n5vJpOkWBUgiawQhTgLM9Isxin3wFHY9Q2UjmeEDCn/gJVbTC
IotCwwr7+IeZ0Kl6JjidjYlTdY7hZCcsbPPVrbwQiwGI1cp7hvA9eK9Ubuju9/9J
g+dDnxKTU+3HPS/e7a/yrAVTBa4pB3rMvgjdWKuS06Uzt4D0s8GjTP+m/G7NZnae
AC9pFGc4PslQSVJebb+Tz5/wpWPqZwxkPMSbt5PYwe6wXQ9e039FtCmXSfSvCQJn
ncEw6OdBI84C4oXe/pxcQbloQpsC8WsTo+MgCMdQQc3KoYiadtDG4iB6N5/o6a4H
/y+tkC31QpO9/OMRV4mws5j+bW0R7LSo+a7DhvG9GGsJsYNpIvVxItnSBed7/9Sb
+g/LfWUQIU5aWOvQyNm1C7Txj7mU6+FJWwB9cqv7ZREd5LZI07d2QMEGR3n5FzDn
kG5DBqhjFGiBjiyG5NsVQZ3YQ/FJ/N9vCw5uKbrq+n6kLCLIRpbyumibkR+fr00G
FmsETk0or21OSoQQPKrMV1Fi/Slpqpuwk356Uh75uUP4dYB1VUHdEOAp+LEWXAoH
xZw4RS/9g8QdnxdLTC36V2jzix0oV4AYO4jWDvw/2/Lf7zJjBe0I+Wm3sNcRUaGH
C/A5OkmFeNOcCZBoOC5rhoP3FztQGU8AJYH/7YjD3Cp4OkA0RlNblG0SEW5lZR2A
t2Yjtu3OpZZifkJgVrFhTtoY7vsv7SI0KC0UfaVm6Pw83dOU10XjfNTrW+Wyo1Ew
Jd7sN3rtAXhfcib3Epe0xEe8kjR4C1b7lVQLXB1SJjEScpOPCsYVqJaF1HytzRgB
DQn08ZZba/o8jNLvsdrq4vYvGe0zzmVKbRk5sqWsh7F0AB6rf7hY1n9JYSpnuga8
fM23trsx1K2HZ6PgJCSWW5v6qrBjcUndMoXDGDrmu9j3eDUKy8f4qy9c2EYGZxD7
rb/T0LD/qTcy0XZMojoTIzdGNvQYUyOqxnpwmpbNgLgmWhlPHi2vAO4g9ybKbf4J
gy777O9ebmMgmY39OWOTAukXwTJWtesL5xvrvKddxKAvYQvVnQGPWNlc2Lwp1c9o
4KZFvt2dgbuFdxdC3rbE4tsbz0Epsj8CEo2n7D8Av7dbTHfJaH9djFXfTXgFFI/B
eX8v3FGULLpV49rAhUPUUflzYtjPAJvO1UYLn1D1f4+vyW+y/HuahjTf1q00uSP7
NPhjPvBfuNVn/bL+aS0pJzZsU7zwXRDnP/g6+6P4/rYXppju8Hx9qgM8vjCTOjnG
7ag9daniYC3HhM7Io7kWY4jFr3bi+hs2goKOxdSE6FQTNo1rZyRpKZqu1Lr9m6xA
dif1XOt65tdvRzGY2Z8nUhND27/GsB9IcQwmg+L0cjU33qmxLuZC6y0/0Ho0MXAM
uCbQrIA3WD8DOsc7B5dMpdVlH7T/bKTJ5W/d4nWXTXEV5DA/JfmWl55+NRvodd89
BOOx+RT5w2ZS3OkQuroqB1C9+ZrpSRcZl0fu62/h1YDDJuCjYcApNbmmuA/uUsiJ
PiLdvGT9oQUROYnLqRBn2NXpDAw3C/vUE32TYEfZBdiBrvBkwB673S4rQDi7SEpn
7OSosugVnV55V+lc0+bQdz2Xk+UWugkBIau91nFBKf73YQdisXq+Yvho+dPVJW+n
bPM6F6TPMYJFV414RrGGBQDXMc4kuwJvozNgBNWjOMl2YtYElCSR/nWH/Hp9cW8o
V92DVs5xqhWI27AcoZa7XcSgBA9fO+NnjBpIJXaRJp7tJqptzAKD+ZQWoHMvPIsm
5mkenAmkkaftdcq7itWFdEUrxmv6XjQ6p9cXk5uxYqM9wGZksiyIINk3ubBZlU/I
wt+Njulow9c1AAPzXJMbXYpn7d50uqR6I4GGm2rg/w95Kwp+h+y4kJ15uquiTyUT
YKu925ezEdP67v3CLf1MlS+VnjJ3MVu1P+10DanM0dplIcx+p9UG+ksl+1/qNVOW
z/8IhDOTvyryFfC7pBaxUPXCgU0WfqDMPdqdFGsmIT99HVGkRtswfI4xruC0n3wZ
io6aBvTU2hgjtUb2guUHF+GNo69brQUjXAdNnlYtxULSf+IYpwLjPChWWP/zzDyj
awGUuu88H+02ivW5F3S5PDAj8krBYexIMliwEncmEq/nDWwVY0bQcHcbC5EHgjTy
NDh0YvYZgjzVpzNYhl4BSKxNx2C7LJBuMijoZYCmzSE6cU6yBuISdEAc0fYCjG6G
wAUMRIpvtaX6SopnbTaUPCU69OC2Fjo19uez6RdGLHpfGsYGVWm5wSCFjL1ec6NK
kYhngs4nlmoYlfNX7XMkC6SNhZBvupK4eW4RvMLVi7MEAXsB86maQjsjF9decLn9
HkKhI/fUXE55QWIj1e82cQdAw1EzzQOeCEgrwqEeS2gZjtfVDFMFhAH2JJzjRXpW
4XIRAPqgurozcoUv+vTyg0+k8iW9MbuSFi4s/pkUW51OYJ4cHk7hn85LfJCFkDBW
XnA3m44PEbcg4/xPYkJvy3xjnPZRejGbNpQhmhi4GI7qxh6PlyBN7QnUGaNQ2j2i
O29bK8S4JGZJxR7eXXwmboeiy8CrlG3mpoYgU6HpQ2zgGRcmVbaWMDA53JPefggw
h7sT4stZqdcyt4K8DznGuPMrwQZmmkUaYtRDbuX33ryO/9+csNyjaWIUOeiV/CW4
kRIDbbptGVRmkjN9Vr+JyTCDLhobqkrkSynFeUfQIuApb51NRUGFK0q/JXxIOFUi
OvQvcaSaxWyEkHKlIsEnxpKz5CIFNpTl16MI01Lhmd5Q1vR+tMMrPb/HMmf1YD2l
2qFxgFM3QUJmGV9dXJQFOvzucQYt6jZIXWJbcUWLxv5AatA1o678d5SOZk3Mp+7t
ejyJYkcFGbqZekggf9Gd7FEkPDzXpFQePjnY2FwUSojCBYWoq9QCf9AGcA9ZHvYB
iTp63XPx0rkaezVXyTKmHvBEdd65mAEVnW6G+rqw3w8Z6P5ozHA0ywsKO/AZ8ztT
1iN6A1hhipJdmO+JEuUFV8vOSp+g3QSbvH+wzICbupnhGa+Qh0iciz2CnUebFhYC
G1xsTde+G0ZHhynNl6OvYxNU+rcUM6KDi04wvhHT6UbWXa+P/+hvemcm7nVoh3FZ
Rmd26Tc758ljPX97/XBvLkIlEO4XjaGXJMOvjmMZR4+jjlOsx+CE4Wr9G7yw8Ntc
WUlDQ4+dTUe769Fs/j30IgVwgPZZlQ+a4prtVRDewj290jTnk2psYjBmeQV06YLo
SsotyOJwMBjbxiUEgs8Bu+dFiIKpO0je+PYkLJyTqCS90Em3DYVHTMuH63NeMack
U2tQRYMlnb9bT+Hmr6SN+7fm115kUtWfke9NX2HiX0frQxomVGaBh2Tx15miqwaI
JmnLoVoMIA57Bz17qxhfY3bEUNxB9nupucAf7IspXrJeOqASgmLWQG7WLC2oD9MP
TmtnghepeM3GpVp4WdcgxFDc81vKBeJWUNRllSl9dSqNc24wpZSVyRRI7b5rudbW
+nQixPvoyK++bj4I43L98K0+yckWUQkQQshOVmf+TX19zXXGU5fPysMJjlwiSKWw
djSpT+OHcxldp72v/Es64DaZxccng1Z+9Cafgk4WIItTrNeZZnspWXGKFZtGeibA
Tlry45669L0c+TG4I8yIF/DcaTDqQKyiu4IjOlZiJfyzXsrt3B0JxCoM4YD0thbo
A+w0anzLD/AOLKe8yO0EvbQVE8q5yeOUX+gVdD8YaSEQoNr63CEbiAH3vM4FTqSM
6XuH6ZZtsSU2wn9KWA6QHfVbMgOJUIGPcdSOqCZM5xde0cbqpmOmuYTzTLMoXa+V
zWrbUec1tylm3lBSt+vQzf66R+pcQesG1nCQ9CXsP4Ogo9XZuB36IGINzRXLSjix
hwjoe451/QD+zsvQplDGfCgniA3tKlEpAJSX3K2w33PZ1H9Dqg2bmRLCawqzzzoJ
bhBD1scqaSfKV5pSeq8d8tLt2sTVyOat0QM1fMeguH97UJZObTWiwgSQlx3WzpF2
zPlsfEPDWEKTtTaidsoVPp5lZxoT1gBC3PWhbyLvVBmrLLtuIx3axbKBzBjuznmQ
1P0Y4ANcGUyADVLI0CUHOCPt4HchAsl8UEBhHCurVNe4fKmP8NhYpOTBCfjJOF69
yOe5QUo1x8f6JIko5kZAO3t9SXn256NZD5RSbM7eHRoRKWDF5Rfw5yLNGR76DmWT
LYw2aG2xoi7am4z45SfPdTE3XWf/ECqrQKVYByprwmMKeop8nkbq0ADCUpaeWI21
iHNSVyKynyGhadflQbK6iDB45qexqZAg5oZ01XKX6D/OU+fG0e1flbyJ53nn0vM/
e1yT+TKJM6NO/u+QXPDYvo7Wlacubkhlg7PFfYnQNtiKw63n0RFE0IEH8kujFxyd
6vpndbnaZW87Zdtyk4wWNp3Sv9xNwjYDKcvmJYDqcZ9bw051NAk+OU/jVyKU//Ah
f9EKTdvICmIb9t9SnIHMQMHLbYHrUptLs0KYGIttQJD/1jjbykEptO1aEwlU1reZ
r2X83W7dniP40h6/mqDHAdzypTJ0GIg156/tRiZKwAZ+1MxrF/C2xA/+uI2zXXw7
of7bn+510LnIcIz77yLG6/fUjRD9n0QSHKx1fdVtIxA/BorKGCJuwhx81pzVE5rd
rR8AwPHKCFxjV6jdVcmmgzZIfTsvk9MHU4wii13RAH7IIM4WVM6NPa6eGRu2Q1pp
Iao7ijwjoMfW0QhTok10IkMysIFjmBAGQSIzoJPA7+EyKy3+VIR5z/jhwM8oPOuT
4yo9NYjskVlK4WIXcCx07mZTYtrWfobis3sNZuE+eo+oSN9mXP/Qa/raenzxEiSi
oXFMuMJcv7qsl/AMaiRxLwNuFgzh8uaOLEhs8yJy/g7X83hlHP1tFWKPIzCfUpv5
ii8dU+l1Kvw7cwQt93rSvhM4uSs5lv96SafxDtV04MZQvhG+YGD4Le0JWMQhNCdr
0WORkA4fQJI4fSwsSONLhGwumpsr7KtxCVFJy01fiwZsuwGY6g+t1wDw0fROEMjd
seI06Eu92Vg6jIXbnHIXF3huUHov7rnfkW80RxsDsUI8uJH/EByTR2PCEI3FV6bl
9JMHhhRSDjtRihpeRFcoKqe5dQWF2vb1LhyPVb2YRYNXCpsQRQ+Jk5bycaFxoDb2
asAQFtouyQtsIA7Sttvd7vvluXFMD3J3h0wFLRqiPmXAt4Vh2rzXUi8gFddQ35y1
oJj4+Y+gFkgn+8HLRqptDqLn43PMUmHIgTWp8Qd0CJEJYKvvlaXsrUAI4xphPu57
pWLwxAfjjeYjBF5vh8LMIhDyo2wafKGPC6/Atm0P/0yN6f87Te0nLXR5bDIqPc1V
Jo/I2AQNfJkkfbfu82EB59X7nRSw6ri2QBwQW7xGVKBfVYlTmOG+mAKfsSOa5h1W
cGv6yDRll8ZO/NyHakXwdhOKaLNa896asTxi75VcNF6RUiCD/2XE251JVaChBFfR
F/8sqPtBd+lg/p17s3zCxlsYd3SozbuCV38ghpSMDDJ/a8bOnxZIpd8gP7GhquI4
fudZTE/N+feFtuWXIUN1w3Tx2ow3UahEFl08U0yW7YCGrteECmh6o45ecuaBbNBE
QIryIsHwzkp3OJQHAF/H68wq5LgYs6fe4kx0uJ6bavg92cYZuzdDDVLSQh1Ts9Jc
qtEJ9ZuFAfchKgW3K3IvF8UFtU92p+3GouEn/zRyhHQI8+Qqn69k3r6fdWm0Tx2m
0gTPZcgOtqKpYzqvFWxwO+27h9fMYMPB0rQpJpU3Izz2UMWhLmioypy76VotxiVj
cJilFzevq+xDSHLKkWqefjRjRXkSbgY0+3NUBDLHd0cjmyrEHod/dkHze71jYIkO
WXZeCe8OcvLqimoZucxx3Z20aH0/SM/9xZEW6OY4qWxG133sZwUiQ47n7MT/WmfJ
rmrVQjISASm6F/4ktAF+4tqZ0qgZNWqpaCTuzYZXuEz4VdLn+zjSax6Mep6wMzit
0zWqG0SavDf4uyOYXppNlpCMN9fSdFT5M099iFpORv9cQK/hNHw50japZ8FCoEI/
HV/aNuuTRpiSAV8J67C+zBRJN7pSAxgkL5p1nFlCxVJ09IXun24k4o8bslOmVild
EkDuBqT0H94ppjFFB6kqSZKA2uA8Raqba/cIBX+oUOt+GiQIgnLW4sUJcHIBaRwl
Osw55Kxk6I2wMwIYDpAdPFA+aY+kerBVKMNTxQM/RJbcDP19VINMd2+PPind1Wkm
9LwbXymIk2DNobkkZwlIYjbZ4qPnuGr7YMyzh4JxztJLE0lZdKEWRiqVkJhbYWVS
Gk/9eu9GMujIP4USqhJtxrd8BE3FoyKubkDFejC4blMH3CsoCdyStuuo+2/7kPX8
635Hf7jRBk7FztIMV2/dvtW4DPZ0xcY0hWuYLlQkCa1Omvm949cz5hax/bXE/pLc
jEcgsfTHhiEkXZ7Ldo/S3xpWUN7k/bCcDs24eO4DszioWMmcz7xkxhNsmgu+gW2c
SO+8P4RTIP2+9z0FfuRFAV1lNzCAyMi9vJEac8n5OdO58JcNWP0KWCHJjzpcTMsi
lH6uKJqALDxv2wiy8N7152GnACsIOnkLltqoEM+9NlCwKW9qjFPHHmHB3xa5DPzn
suEEW1qhtA+W5cpub3jOlAkAlcMSP3ilJNfDwKwFoTuqUVCfjNx1zZwEMqfJSj+7
dYnqW7JunlrmimM1uqTyHqL9uho5gCRpDWBnAzZpmgWlHxRQiYDtdYrn/oXR5b13
gsg8kk1Pu7eTjlVcp3ZV1Ug0AmIVF4AVTfnM4uZ13MH7/j5Jg6lX7jWAeyP1W6Ds
nb5LtZxP62KsY7OnO1U7J9MYgCSmUyH+06UIUCX1M4dkjO3/yMhmUkhah9F2OJAo
Ixdpgj42reMiL9MywBadcD7Lrz58t0vaeTNVq8G3F8ICIqLoMLW+sjImotqSOjeX
JW41qhbZpnpz4H/vy+63NqdM8N0LbTsiIkXv1KPyCd66D6z0GznbrH7K6+fxIhne
uQ1lAeOhhHMzBSRtF+8oe5afaC25qAKBMWSUukYtiIaXYLQnDg+W4+/fwySXc7mG
hd8QlXFlYvm91aHOcrUUWRBUmk16fqTA75iDw6Wbl2xPEG8t+4ZefMi1TdbiYJF+
lp7VkijgL7neiQrAqZmSikNbh+IHlaiE6FHP43axxLfnZXC3eWc0zAg+1JJMfFML
z52fYhMUZpleCDvB88Zp6DPQ0EJMetCAK5rOm1ytVdXVNPYQQnzkXU3tPuHREZkp
VF4YzIFFrMvno79KuLwYNVzICQuKl3LJLzx6UGkiD+tskT29AmSqGGFqA3CJ4yWu
/qqRZyTAEXGY6cuXtIDAp60u9jnogid8Lrxnte9gVD4I7YJ9J9dD0qZEP9IsHxxN
zgve/PKF5AWXSN89IxeWcWB86GKoaW9Uv0JOpB25eHZQvCXUAORyfgm965EAEQv3
04r66oijkLLsmyb1qj50EMpBDOAJmHT1u5L6SbVY19CWy77Lhiu1vtrI0IbAs0Dl
frYUnxhVoDqPgirolmAd5eH0ggo38tfj77bs1yYwsba2yboiHnUQrLyy/5P3AEOA
BH3O55ylrwIr0wj+HA3R02D3ZJtUUoGs+Mg55SSLxsuTfsQYr8iB1eayF9p8R0Ie
slQbLNW8kk6oyGNulD8ewU77jZa98erTPpuKfaF97uJkvr1zxZSrFLBYYOE1Nlbg
n+4aiydmvvdFvVeH9eUudFpKPCEFp6BkT0ews4aWU/grPLTPyHkv0hdsANGLS0Vr
yFKUkY4eTX9K0LgFMgyU1eDtGW8oLPk+IJjbdXND4VwE+b+e0UrGADKZEIQyY3XT
9KhuzcuFJRO0nfosZKdzA8x3ciSSfYKvjkSUDI4ZdAMZ9YcBFeI8SYSEmErF3iJb
GyBuQOJ1EZo4wlRgZkR73FBvz5Kopha7o+VfGFQAA1F1Zm4E/hujZxlZbRqlSMcN
Lehqn0rfx5kGd8yzznJBfdfaoXW0FPZLzkHZoL0Cz4bBqh1vlo/XO98ZywfgmesH
hp8nOZnzGWYG1PUT9coqFTnvG0yREtyg1RSVNgBakJbC96xbkcCOXyf/u178ITvD
e8TYFAPo4zK7aC4VvnlOy3sjAvynwtp2DXY22DxUYKg477dWIS/H4l1qylehAzRj
61/mYT2KHkKmBLNR7nwWiahyb5fRmzUjA1NOgVS86WuDdQTpnqx2MEGKON8B/tal
cBu5dCCoQ+FcuX6XwgbI6quJ6gs9X/cpoT4rnCmgjJ1BXUnodr+p4nHelXwfYcaH
ZLDKWogOcg/WxkHjLa/tPPhb9rGpzR9YpfRiqhsbmVKAUJNrkYFURXLftsYl/HlG
h2RxGiYrg9QOzosF6M5RICISVGnosrLfVJEH+d4o4ehOuFE7+trVYTYUtBH0/fGM
HMW7JWsdIPJb6ZSA4Dekhau0zuOxKI+hTtH4WYpgQ1L3jn7P954a6pDQ1+cvwYkh
GPYfwmtibnzqP9aaIFqwpLU/ivexQlphgfyP8hBI+nZBoaTNCD7czm9Snzguha47
oPtfNy++348uhzjgKejMq8J1ggD7JKO4JyuTgpoCTF94N2Fxv+EB9AMGfjIbgwUU
xo9RDQAEkL+LsuirnMRVM6jN63KVPpXO5XfznFADCoPAPmELq2CsyKWpbWmZu5l7
EoJ/jDQN6deyW890MQcx2Vjxd+zjisKaMfJxTvECVC/0gT2Pp66FZw/8vmZPOeZl
126pWCKu4kw9KDp58BevtxlYGk4EA4adOr2OY/ibLvPcbEeGM46CeqPslwNSBrBl
/zbB2ZcI5NY9l7Rah4nq7dx9iJGZA3BCwKHytcuT6WKIGBKjD0JZ1OZVaa+ohSFu
HR+tV4tBhui1pqXahHt8GM9x/QhkGFmLENF2Pf5qd0MPxRxp0I43xTFS7mrZKEVg
kk9OoEHz4BHit6cin26ppfNrPaE4uyJeOy0ZAnh+iBQWdCaa+Y6pPWHisECApBXr
xfJsLvhp+HuwvtsKxLpCr/WaFtwUf1WFw37M+Yn05hgZjKVUPK4Lo0Vaz1yWBSUQ
xYlAQXzdG0hVo5ZXKmXJsGtLxl38gVay21nH4o4z1JvoFUjSUvAZAUeyVRlN/vJI
ooKSLBAIy1dR+dunltzmyCtCEUbhOde5hb90KgMrZRIBsrju7CJEjTl/3oGbGl+y
b0qWmIkxY1v6aqku2BPu5ZD3wV7wecxbsPRVswABKcn9Ff6yYK44rgzpPEdx1SJn
CpHjVCugPscM2easoE0JCaPfhl1qkBAGMfPstlPE4LYCF6djuOMWlHzE6au7kO4H
5qqBdnDBm90CZtZkyDAq1iOh6eFb/FfmZPQhMTFlzkgSuAw20oHKqofj2yYqO1e1
LD4vrZsr9gM68heDEk+GlXLEzP/uQ9djtFPALdy+B3hW4SaTT0KGRh2Yzf/8cObb
CCvDy14Jx4jDKHKM4yAPrX4vmnjm6IRzaQ8DkgcLoteAGuZ4JsrJviH0TcjzI/mc
sGWKNFyMEQV3Hf+LKX8bf+P9IdvCPC7jJdjfATPcsFrO+jP0XmM30DkIH+xZr8nH
GwkaYAozGFaUIV3/l3L0FV0xGyhHEMd7xjzx5d84pwBRUh/rC6upVpIFiSC87MZX
uVYOg1nVaWjNdnbZg5IvDOKzNAqRaEKCO5dirNOybQKMVlwguPGNrE8Se434HvbJ
ZhgDt1LzRAi5/brl8bjcmgV+7xOQrVQ67O+nixXnd0rqvPClSOvDT9Bc9fPJx4lU
gmicKvsfuJZYvSfzUmJThYUBWsTiLQy1E5fAQoW2/VxQkTXGZe3vPZAfMeZSTo57
voj3KIzd5GpMIxcQ+eFrGgdyKVh7phKMgNWXt3ONWAAmv7DyoyZszqIX34XcDV5l
k7NwVFEC8Y1erDbmgCFq+EiBym0Liu1Rb40UUtig7lk++sUDUdy0b3Nx9bhw3nM7
YXyKps/bZ6KQE2Vr75ojxlEP+y2gj3dqNll1p+PfqAxY162JSOdQirBs0s6TJRki
SKLG2sQRkPmm0m7VRGkq2t7amn9jPogWwgFKwVUsPPHusJ6uDAUdEyWdzUyxRRUf
A8NYJB8n0sLGVFQwZBKYmqtcJcJgv6xhRmHAaF2Kmacr16mBSoZ0hI0ainsNcmee
mujFHHRUMGVdbeYOeCy4L4Mg88l3ZmFqyaPNS+XfZCchDUXOFZ5EtbXQFxKBs9Sx
9bUpsG59rb0NjUePiVv72jn9RdfygceJBe8gPzdpekeHdeQYL4I3SahXKI8ZvhRN
OHr30rXUzozwjkK2BS/IBbOCClG+3hSVsmYNtf1vwn9uxSGic4cspHbkv0JALfps
rYXlEITRPpX/VE/jSdhU6WlnAgnA9aVvh4TOxS2rGNpJUpbgac7epgQmSg8eYHPO
RavWm5hL+JUrC6kmrq1DtU7ByBegl3FiVP72aui/RPO4Cxgqa0h5udDIBylWa6c8
SYiVccbVfItoAEzdxOArQhZneOY0c6aq4vxOc4LQpeoKLE3mpqOOIYLwXV6mlMuu
9i1qplbBxlme8GuxlXnQPoS01Z04s0OugiiFMdf6AhiL/SXjp5p5NsXqXOZWdaNc
LLBoTp3sOUoRlPu/Mvp4ryNfbvvyZngy2sD8F+3di6FB3LigT57TStIVSppnbj9s
E1ukrIJpmWNNyQpxx+ar2x10Sa26Jj6FUUB1q7Ub/1hvAaMgDs1X+fwnO1rsL01e
EXs3Y+wmcYGISEauPpGmKbjOb/oq2/zqffet3gajzH80as2fmBDjZkMv1rpwkp6f
jvoTxjFXaGicAlC9dbFUAhdTsS38ykbrjn+1SlOXyMrJyCuOc/XFAoTl5VfwxSpZ
dpP5oDsUxoGbGa+Mye1P05zAPD0IpR2GatQF7dRcO9V5DyBad0AzJoGb23oNhJvh
dzEMsBR4UMn5QFBNrjnfWUkX0240skFml4cURC6W1h6cL0iRgI4c7TsxUY9kTWgm
vo1o9+f7iHE4w57yOv8ZfsQ8WE4NjGrvKm+IOo4se9+5d0mwIcjKdYcgZJTt/AVV
FcyoLojJ2ZMapz0BFimnlVht7BDxC+acRITiZYf6jxo1V7iHrCCgalgo4dC9cqLZ
j+ZMTqbjO2gXh55M9d7Y4R9ruYFXxWKAKycR4nIaKM8S6w+mysTnu5rqUIhqosyA
oGSgYRtai1VpB/teqAh6DYD3aKHXCItPzWX5Cz4C2ihY7fL6npcYm90Wcp5007DH
L2Lax06PRglQ1PonXlAhkTfJd3cTWv7OuF9Ft+dQid9o1GElDn5bBiL4mnPxAfW2
JixBsbdWABbxhjKiSlwG4Bdw4907EMuQR508b2VAiqh1M68vhwODiFNOugRn2w8M
bJWozKbfjukeNi4SG7KYlAMUhfup1MKEqFGgIszHqeHXbfc7GnU/360lGkImNHX6
S+1cmhebjHRTLgkZwXs+dX91P8dzFZTSHl7nz/m+gFRsnHlj/Ajawh043g+PhvZN
DySSumQ0cUOV8+jsJ2LyDwDCec6QEIVzZP1iLYbOtVtGWuLUvZbPipM5IDYryQ4D
S+VtmQQU7RI/YCLCn9WTYHRB2XwCxEILBV23QNs4xKfpoc08w1zuUtx07DKUS1Dh
/zMyGtSffpc+aLs26Zbbxy3xqDGv+iyn8oEQJrtxFkZLD6uCGhtYyV52kGnSZc8b
2tuS2/2CsRw7Jv9WYX7i/kzhLzNjvEcKedNnBd2i4UK8rmHmTFOM5lx3VviZbbOB
701QyS8HVHa5QYPZ3OkT2pWVGEPJo6VeguG2KhAosCR3AMeEiBwv4Nk1l/pMsSf4
pN3Ab+7kkbJSeDkemcy626mYTISoQlF55oHXQgPAa8DfzHKHp9p1/ofN3lmFPfTZ
KxkUNTWf+1V97bmoE/be7g5n2F+02gsHv82mib4H8W6zYtRRy1e/clu76zOhPJus
jvMUP915b1NsooUbKpqXOFTVSsFdZMT4wlFdsJP+4FUcib2jUIuTNsyKjMMAbQUx
NcpBGvsIgfyhr1uBRy866/ayi15ZleIFZgrkfX9OiPRpCVE0DdLJnXOgWMkh8wj1
qNpJaCeO3DOMomcMyu9fIfNC0UuerH5G/D42I3NE/vuU9CRdFycFPRXL7KYpL9mz
rYf9Pa1dYEK+ZSZ0RSxiNY95eK/jgjzFdjucg6fxM1KodPk59RYfB3p6C0pxv7QC
gToIyaEtxBdLmimwKGS0Ji4B/AxYb1j5090HfMtJCbRI1+CLvtdU9GUH22EBzMiZ
cmiXmrFK2z4iXXsdF+XWJgluyASvU/Tj/uGd6us2TtIXFIvbBmtoEMGn4PPA4tYG
ki/g6xgf5cb8bnzVS+KcSZ5Nw9iJWDz2a1iVy57wr7eKd2GEnJiwGU8aPbgV/mxk
5PhBSVBSU5PfH08pu35gRLCvqHN0wUFbzUEfo+9CdXNO5HUSxs37rAvWvWnxc3Dw
eeOUKGhu1qGKxpS84cMZpJEtPJfPbAkxa54ik+38tYQmxaoI6mgcLf8wEgvLStPq
6a5D2GkyEc5r6NZCB6SCZP4e5PMAO+XBSgKD7nQiaWT5ERQKDPORV8stjnToCJv6
ppoD9Xq5MbLPux5ngg+TnurUKQiELB0TBY6yXKk9FeUrj3LygkuE93/pdtkD+Q3X
ja27iCiknXwIby6TgD/DiiBIPYqjn8+exRnAo/etB2tpyspPkqJC8SKHLyW2QhH5
3tzfI+0mTxYTr8phvkQjhbG0/G8L06L4NEFmz/Ur9v/rs1OM3g87pAV9HrvF9R/t
IOvUZto/jL0IvDvuSNatSbUbbCiXmDplXebHbd/fybZ9RdCZl4kPgPAJpvmTXLc7
Iex0xiTuCnzGIpw1ftA6Zywg+K/UCHDbjidMyuqrniZO09uqIl9ABYnHEnicScoM
YwQ5FAfIJ0j4YH/LAZO70KJKXtzWGxVnP749y7LQ+oGxPHX+ZlTr8gnx9MqgiIYG
bdoYQ91ibhAJxejXmXdaiL5Vu/1n96SXkRrG2Wf50oJ0pSe6iPWQBPMNjYgvzEUw
hVg7SUDBEh26LLJmXOTbhDPXaXw9pQnB8PtSIRmAG5Wf4saH80a94SJqT77PR3ZC
ZBSjax4yn3TcvZz25gDM8zxIs6Wy83KlpmdtPulpYuTLSshOjq+Aue+p1jRnsk3/
2YHIy5UIy8NT8WqUmsPTcxBstgJNnTO5UXhByviHeT8Pf+tQiPWX7Ng7/sVAcCD9
XFZ1wiU64P6FtBRyY4EIrAtuB5wEGMQ+Fa4b8cLnlV1oXP/NKLYq75JySDwPO3jX
jmA7xv3M9PD/6WJ0XfEb3FpzfRQzgFPj4VT10bVEHMK+T6JhLqcp6QTr0RBD/hNz
yvHjMdOKMl0MFCrrS1lI/L2eR31VJvsaTxs+ZBz6KmYSZxmMj2ta/MZYXAhICP7h
oAcY74KirggWQi2z8GVZAnbOxPK0Y3AxTpEZwzF6BFttLF7di9Av0M2ChQAYDnoT
TtB6vJzJhRq3PRWv2ZSzNiz1V9xRUG8wkQctSgxGlVMEgz7NnD+parAu8P7H5qbf
jHfM/ZRu+9gXIK7WGSyqoytbhk2d+PLBWVUSyfFzgojU3vn0dFrnm0Fedgd/VHMe
YNpih8eajVr4vm3MJl2AtPSh3PCG+/z07te2RJPI5ROuGfqD4agt6u/CxqpWMUZ3
jFX3laPCI6HfY8YGH6o3UlQcCCZ/KfknDKTEsu1GpsrYTOgrTExWc1GGWTBqjHee
fXmtdSnmouoZnZnRnnh1RSCyrdfbA1nXbTIbWJCtBgfmMk0IztplnlyUsSS5ZsIE
uldkAKWcFyD75FI61vRAJB6Uw7mSyfSlTW0/IH+GD4Tlpnn9K8reqryiyOi8bLKZ
dP5/Nq+aqpteFayofB7OVLrAJRT0i8+ZORAYE7+H8xWSHmSf13PvoBY2+eRwK82o
imtB0Q6DfOdzS4xYugNrvI3++nR8ag0gPSJ4BGSQrRoLghIKTU2nwmk8bmPR7i9Q
0ewzJde6UmC8Co+W7aitIh+J829r9LfI8M25s2LIRypXqjfdgKpbTmxe+EFaFm5e
upNIwPw7mgV5NLBitcH+HpP32rGancHJflG31TW2fZ2Bdg4OjYjYeF+S5cfQMZuW
7weC6FCqJcksKlTTCmE8gi+5GHlE8g4mKbkLq84r3K/ZYIdO00J2GzPN9O5vyC4N
Ynkil50SaHLNXixjX/kfnA4InmjPrF217ZIAe2fzf1vyOeFJRH81fq56vQZ/9t3s
gaCXtfxA8t9cOC5tDfXFRK1O+zikU7AAD9eEGahfV164co4eqCc209YVdEkjb3mK
8lvFzHDoOVFEQzSq6Jdv4dDv/Cnic1xUlqGiw7La7CVIX9pZAMrt8ysVuRP/lLxG
oxVP2izfSfUIzyBNTBpcQo+EE3YsISU/uV+Q7MysYYQ85jYW9VC1kL02MEOvFdud
tMSQGeVf8dYEvAS7An3Qmd0g5Wq3U/bfpcZBAxSpaf9XqCNVbyGe+eXw+frQy+HG
GxZ9f3Z1C/gCMSOEyNCK4jhIzsIjM+3Z1L0cfO8FiLH6eW1Zh2C/HXa6hMJzBThY
/EKhnEt4oCw4li8EfEX1+5x+W67AzagkIhNw/UWqAlSkf0fKZsrM79tlFZDhzqi2
frp9xj/ztqznqc8Rzkw7jg3We848Onsgf+RlGx/D2U4nxsT5n3bBvvMF6SCPn5Xq
kSR5VJwRP0TerCuj8B/WlCxa0aDVQdEeovdl44W8NJvqibfrU+r895EsL/LZdHlI
dJBRRgFFbdwzpFWiMj5gtwIpbAN7OnWUkqcut3PPXJ8tV8mZbDDy532OaA+9ev8K
z7VQZnLV56uzCoZrF4L1EX+XU8XD6k6RiobKAenuW81mhBkscgbt0IeVWNFcInjS
yefi1YvrM8JKgbra+fiZnf6F1HOCfbxwBEx029BC0RkLU0+FKfXZFQH6BEuZ9JMj
x6zOEZwqwQcNsYKnpT7EKOYlg2u95vr6c/c2ac9Vr1rbNhArKFjx5oCPz87RHDXt
OEMERvBh9nNEn69Pje0SJLqrM+Xj2bwfbA2iWfmVHxNuvwafRXKipA+JxbSGuLnF
kD6KO/uSsM2k2pckqscNlp3FrkPDay/Yv9k2Hfvqm1ItMf1vhcFYAQvJLj35XEa7
5CkRaD+t374XPQqSVBJ6E23f/amHg7kdvGf8bKyRabaiTEU6PyqwrzMYmyt3B6+m
4bOehY3m1d15OyKK3vgRJji4ReFPG7LRJLXDn2XLvDQyttwoFpcn438LF6aSpFDH
LCLzK5+dL6RWKwJ0Gmh+5BnR3G8XYyIW7RM3XANWaPmMsMAoUoEVwIVhN3UjNM/h
v1JRP51CL7UfjegTao5awrTE8UxeiEVluiVa5jimZJ/czzkIvUgxq97h2D4vPhBx
88uHVwnVt6hreXktkjSkxagkUOfB4hbMQ905raEa9Vb1N0BT6PuYnBl0IMiGbYwH
pNOk+nOEWAKq5EWm5D7R5CYXxKOA/Qa1ZV0GFXvt4lQgVTYpyu6zq1j67utBURsQ
e44LeZEUbktgTBQianNljai3sSc/kPlyp8tRGLgkaFAgCnFhpo4MkbPIfTRY+1hW
UxpQrnv/DDSAm84xeQxPJdVdtyH1tx33tyTOSTOJTupF4mYXh95kkURfz2OH7MVi
52PRU8oe2Rw0bIAzcP0XzgTU0rk8SFSrd3e8LZSkakRGHIeqa6hP/ERZfZ1g/LLG
yZEuzAzAZyp5Hb/kzRc0yoVaVAFp9YSgvmcsmvRan8Kd7YkAOROnkvJHLcAebKIG
pVt7T97vptT66EYrsCKIKDjS0bcPU7wFmmOnW3QSpAOYKdvyxdFKiwN9zwV+uNYR
8pw4M+Sg2Ou1jnHgTcJwELiTRve3Xe8eV86zq2MPzDeIsdyimN9opY20d7onqDjG
f6f7pSTcEXdB1r8tgcep2Gt9mN0lLx9fUPrGgpdwL/FJUul2spHK94ls8rMFv0T6
gSLrB1gLWtVdPcbOUjSnD7x/jCcJ7ew28BEIZAyCbpNv8CawcAu4isx1amKppAHt
P3djAvwte60WrSi6Bx8olumZe4wXP26bVHCz+wNqvV6vSBMl1EPlkewGX/14m4tA
SFMWnGxAthlyRjYHEWOqTm4iSMB3N7az8MYjRlA33BPPhdpMXIC4T6cX29j7phBl
O0biMDz4vddOzaH7UjrpNtSKiQ1ElLFh/RsH0qXW+MPA9pt4CD93lda9ZinP5e4s
21f+ltlpsTshkmDACgpQTSS6VfnYFxj9QqNZCv4YS2GYBGsFwkQtQRUI1fbmF5ZG
PVIGMtsypcK0bl31ycMwvvC9LdHf9jAkP9kXxCtfDLh9fk4UisjGS6BLtZ6NxJcN
Xgovl7yjcFSNcqRBUw4zrjBa4sZ3MC3006rVx6e5Ngfqa7yT2ByEQegRVNxJqFC/
cTok1RV5Lem/kp0LXAUFzydD3hu/tys5+mccinGVxPkbEmLFYCbr58P84Fu5oyUn
xeWEuxyQiZbGX+L4/GVcgPiq+CgcX7F5N0Rz72+t1pCG7zc5rexKpcmDgv2FruKx
jwJ19M6hnHRafG1Snhpoq0esUZ+zj3jPE1klggFnUGm0MJd7mUg8CX2WWu6/BUMM
2JiMt1iNs96N8zURDqKFt2tRO2Zq6FbqOLW9in6wvhRWsklFXbBP9ocAmJz6TFhV
Iga1XTCrl9r3n+505zAMo9tFbe8JgLxHWBGYwvlRxKuMuNcdLvdvOkdfKkBH5Woi
7GbYvWoX3UuynSdnSk+f7H6SHMG7xZ77ufD7xlQje/Af+8kivLuvn4XnZc05IJlf
Uy9q0MXSpeRD+NxcCQirtCV6yCtu1wmc67kXlCo6PaQugmjRKrL66fVkeS5GtHfX
PMU8c5kAvWhJY3xeqXHkF9akD74XWrOQK6Jxh5BBA6EtH2sfy6SRh6cnUbZahwAo
7qXTpbPrWBhWeiprpkWIZ5Me8DObgJMYaYQ3BCAqqC33bWGW9Run/FMurFu6jElH
+FYsT/UdIslHc2CN/lv/2XZfN67vXkoxr9yYcFNweMXZYLikN/Hug3kDHFgPSsay
rbbuck9dCPtPtFNyp50oi/Zxwes587Yl+v74nJtXOHAc+OAQgVaV/suwh4cMHCCW
FR7oOokpS4tI8876Fzm3/w1eZR/QuxWTLm/Vm50C+jg7pYg1j+kMuNtRoDxh4lDL
Kb/LcVR2N47vng7+iSw8ZfS02b8CqxGN87b12UVADI8X3v+PSdNHdwijsr/ktke8
jZx4yWkDwpbXea2FPXD3YxrK6dGQEkmMslZAkUKP2qv0sjv7iU45JnC1dTXxIMVJ
t3Iwjg7rD0UNXAeEC5BkZO3qfuNlMldx4JsHAHCKDEgUawZrx9ZnRDeo1YVSvmGR
VeQQdYaVUQRvNPJEx8nMa6fJREtPtUAh7cYxglU7eYrcCgAZiRc4SUD2frPH7Txj
bWLHvu++ffJYhLOg7twpePJkTC0eL3DfyiOQCCOu03EHIDLDt/j+uZZEjVKx+TrM
M6hSB+r/FsrT9hiqe14CNV+fMLROb3NySeAB1/snulGytQri9d/pSsxHAeYJtPyY
wdqUQos8NGfp+wga2bAqEpIbT7m5Prbt5NmgoRdv2uiNGkHkCOWrqJjYyHB+Igvp
3ConhmRlulKNXNk3zzwhgb5UWXh3nPtt6n2pOceEqmZig3KhmgsLkmZkm+rZ+wxN
E+A62JDQs4XdyToPHtgpkzdhy4KSDbY72FATCfwGuMWDyMeflQ2b2h+jzBGrTPTx
ZWjJhEgrziPwtN55cS59zwNtHvkz+Zq3MLqLhRbWfP2kBwkbRGtNT8sYrbELuzyl
p/NRGZ1S5HuCoi9LOiH8mTSSaMNJCZoRt2bIukqWfTegr1NcI3zY0+r+xViKnRyi
0iSoupS1sNK36oe6yV61QxQJSt20DUioygpCla82Ttoyv4wOgJ7f0XfshDUQLc7W
XguW5S7IyRpz1B2oSu7CX0lWE8TnoeZ85Fh2NUaKVi8H8xhQe6C1yiu859LrEfgJ
+gIzyClVoD/UWbuB0tFHt63+c/SPBBroS1ROUGoZCKg+UYuC2Vlt3+B73I36JvDC
7nugNofWG/GySt8yDD88kDK+5u3Ty7MNCc5xHjytzx+1IAVIllJn1/voiQ02e85Y
jF6yEZS5nUrBKqqHRMx6Ytc5EhmPkOsfjiAUcTuYrmL2F7+xfHHfptXdwUldUPAw
Vo6xXtM9wz73jPQ0Zhb8QX25WloBDCyQuJgpOnDFIpjSKYPRjMnz4rr3A3kOW24l
10fffslN4WCahX8I191slXDjJncurubXdOQ38aH2q4YcN+s1vS6tXPmeTPzL8SBS
ED4gAxTQoD96mFgDkTWL56fcrHRFX1ShjWKFMWRmeZGMezVLo6QfRd+/2rhyHZm6
fuiyuk0yBJhcwvmcfGx8ApL5IDtzMRQE7m3iF7uZi6axjZKrCeprwHXBH0crUjAh
1lSh6qB3gmI9zMiZ+ndPrP8pfYLTPUEdZtD55+RH3pi1GpeKaLz/2X/fQougj1ng
lsve2/V7i6olP9t+kmom+Izcjj++VgmMejXAMeJqSguHYfOfUXxXvpdoLIetWSHR
Z+hs0sS2dJRf3Ov+5Yl+OX+K+DAjZ+sKL9AwD7QoTo5twf+v008y/RK935CvAUrf
6wgXpgaMWc17dE6OmoFs1Ba1Oo/kou0awVKPt8E7kl++BxiXAaZpb5HfPyHCZNXK
GyyMsyCGguZ/4h0DqZHzrK8CXNSzAmRim36r0Dvmf2o0n3jruEP+HynYZzvDio/d
Oya4nRouJL9Jt4GpXo5CfFaGCO8G1RIYS9YqaV+sUqhqyU6IDrPUZnuUM/4kIBni
1OpYY31kYNnEMYwVsJQOzocR0TOB29mrIgEg0vxgBVaSeG/iwUMrUnTm5sBv00HA
DTS0jUBlO3nO2az+3OebfKXRCzf7D/l7hjrd93oK1JGWEijkoDccHQ50Q7E1zRAC
qmwMvYj4Mz/QbuvbwMnTYdvGyy/IYYiOphZjUGQTJbpS84GkEdkOA8Zr3QPKUnlj
OzM4Gg5QwdpIiEgeT2jx8ESTFsF6YBjYQqDFtBFJNbJahWovYU9ncya2ej+eUvP+
F0Tm2Gr5m74IH2Y91HSzDyl7rbAk2ypr3qFCuF1OWw459p6t3LMosgLSSxYyedGT
LI3/mup/XgNb0Y9WPrI1e3hHhz/CgMNFudXeHcbaJB9hXTFy0OXKViroccW7qqXY
upZmUexZxJ0YJ4VHxsRXbSpYbWvJZZYmTI1WrHiGlss45jp8bg1cYUlIZJuMyr00
YQDTlhx8CPk7FLlJrH4sQPxW86TBA+wy7uyDjBgPK1Vea9hKWE8Cx28TsfoVEPF4
4Sx/mYADTpleSIyqtF2+vBNs82RiL/WO3uriEH90FDlXvNwVLTkeoD66JQHUJHQt
yFyb5gOSGx0kt9fDzq5xn/yZNjA46NPvj0Q4TD92REbnee0uXqqA4u0J7I1CDjHk
bmR9+MZlDWMVybG4p2MhbUQyJ774v7Xn2x/MDlGARG0PHiiJd+dR+aT7exF5C83/
gkT//R+EuVCje803oCjSV0zWATu/yE6f95bC93sXYqDdn9j4MO8w7iQlVHwnPFZ8
9Qw7jc+kQyu8+/dGOpxLIPW+ipXlo8UWY8YhYmIjwApzupstlBeLrjsEITZwRovX
u3saxaSf4lNPPUApsHdftYA1TkTpzJViYhGH2TUx8+MsXgIplk0kz4MFlkVSq6hR
CJFOhT/6RYbVz5F50EpdjP9SePWb5krucWuYX9ktvZmZs505irvmYIn7jooKnBa5
9/hcICrCtD3vM8XCd6B2zvA3UTRmMOHmAjK7P0N/OsSCAKwe/iX2yeRs9u1nf1NQ
QcrurIeuyggkODDYSHoO1nj221tC2mMb7dcnJaHvCrA2t9bawGyb/zkDBAqmEgtv
TcLrFk2SApp+sv9i5SuDIKM2NGb7153jnsT04bBx6EOkMIJ7Z4WoqoQ1154JzCPB
BZCKGO/5MLR0JSMr82fiHh54xPST2C1rkju1mbmAoXXRIIBb62HC+s7HUzJCgeSe
3VazdrsPrjsx6Tscx0/jN3K7p1nzdEER6vbLmfCfrEo3I0KTqKlIZqreG6XCDq/i
8J6ly/A87c3gL5W7vN+/k77Ynh3vCCV5zPbUrlXlYmh2EhOI+wDnYKOAVrXUsXeq
t3hf/ZROogptVkbizOJOtplKcCFOCD6Ndk0EkIvT7/NLBjlArjq0oUS3+soWtB8K
R/cI0c1ttjV9us9zLnJjUCl9Wgvf+EkBRPRmkTG3Lr3QI5Wc16EdmTum+SNXekm8
t/xGejUDck1eY3J+Ch9VrKVpfzGVbQSHNuM+pL8ARsBobJc6BbfBWgtCAR5NViW2
v9iqpJp30tWvqEDQF/PZEXE9Hl16A9mIhNa1prhRoVkHS9frG9N9XFQxPh9X3HGo
bZRN42MNqkx43zU8d/PyYQZt/akJl017PJXdbkNzTJrt1tGaRPEgXCVjgXco2u2P
soondymwNBwXHiCeP9QzipUiMDk0M6euhPN1PZFgf1utHjOcJeVPTOC4WsRLz8kZ
5HL7EneNxgB9E4ac0OL0Zth6lchXo7vUQMoCwb14VdweONs3gZuOnUWsXo2sWoyf
TEbkbd7UpAQC1GOAEBCyOilPqUPoYdnR8jF2XNCs3fp8dtvtI01FBRhOO9UTi006
O2KM+MKSj0667fLyaFmgm6I263jaipFXmlN1P3nfCBvAb3LW3hDgobybosOZcxKU
lAvybg5I1xFqgWQ+ODmZv5rb/cc5Ga6WMrcfFL3SgJZuJ+RC4488xlQCLdzt7kU6
V54hdXUccX3tsp1M7lq0U5BpwkGIMeIE8nXM8meW1wm9/Bz7R7XsoHk7JTy7LM8R
iJazsONL0jyVawwAV/SSkvnOw7W0q0OzDuRfKAaFZR/0wQmNZqZw3lw8aBPFmzw+
HRyrYR/fdEsuQsjNnDSTeaMfUDOJfUXAuyESkRQanS7EVIt6x5jcgFaNTqHy8zNn
0RVRFSMRioA9VVrCFEUAhJqoX6N6eHsl6CU60cDsajDfQz8S9blFKVAcxZa4QKlM
C/iuujXepWYPxEUKStRfBz1xG4kAHWvm7jtr3m2hproRwafP2qjTOb/fuOeFaEB0
sFTuBVMYjizaKfpiyTYZ3z1FLuUPl+A0oiVelb2+ramT1ZG5s1BElTRoNA84q5Pv
kFX/VbsUpv8MoA6DDsXZOZuKrJAoL4GMlVhKqUbjc+l+BZUpGCPNcLoLhlgCpl3D
4/NeX8m3jBibRBvSKe0AZK0epxgJDQYTBV5c76w4nalo6zV0yDfTvASac6xmMK0e
9vTFfcD8wAReI1pcX8bOrL4+W49gsMmCL6QQoGw+r90CZ6sl8S7YrEp62+p5TRpp
OFJ1Bh0ycqXgR0tX5kEzQVtXzHcTB1cqIp+IIE6Nxqp4iRIM/Pq3/c1z6CWDl1ls
1oPYi2sCx5UCX7B6Fd4BZDQvb7+JutyiU3Sq8PVoB+FtBiifaP5q2S75erY4YatR
niiudh4c15Nbpw4KInvq94gFy5QcoNIjkTSKDMqENlbEuU3lw+lz/2XfYtTN7WhW
ivd5jQflEjxT9M1ZubSfsrBosnvrsu0vPbtcZG5pfGs50yoGN2EsmidtAjDn4K3h
j9pMpRX0JftkoZ2fiYrgaSdHrcsccBWAWTtujz226Lx+8WgcxvWna5ju5b6P0okU
W+Spe1RCe08As01ba82rd39yV+E0rgLVojpsFv6VuFvmv1C88We2P7tvSWhvImzT
SVXE5+d2Ct/CBuV7NRz2mc17ooAVMujqbjrorlbhSFvk24cW4qYOcjufiPlZetKJ
BrWYwtVoIjc2HE/sB8uNkLpHVPaeAQJe1mReDDlO5hUQCXbKwy5iW7ZPKlemKdNI
58iwNmNwyC3t68sJFud3UOA60vOZMjPAQLnI6lfTFczFt+1R588Iojb2nmX/nDZk
eCn8IaTkswPjFk+z6JSS6G2V4Fz3vMBN+3kBskoW9RDvebuUU6Y3Ibk42ozlxvUd
U/VY5mZHHXmc7frvHa24PNrvGLXuney/AdhIZaTbof0zJDU/Irg05p94UMqDOweE
4C4ArHMvSU+dBeGbnm7Q1mG3PIXBLf4l/euoTZ+Oa/7RFAa3DbcWgB4BTD26k6N5
ZIb6yUDAWcjQyt1SsaBb1vt5JsZkt+yeZJagIp8JwxQEpiuTC6eb7mUiMedX3ywz
Qcq7IVXeNXX87LY2QsPSp7PTrQYzzO/ctsTzfov5RuxVdU6dTHUCMhmSyuPeVL8L
J64B1fTxas345EMVxzBxLFQFaDGMtmcStYL8VCMNqM7j+tQADu8vvDP9Vjv4Xwc4
XAEmQAao0XYwGAbWpl3fxcQVNtvgdTVwxtg39AmTjoJ7uuOa4I/JVBRm238g3KRu
RLBGFNHnZ0RWkl8niQoXEL88GT9GEzPpXUQPbmTni9UHQnaPn64LVlmJDsyimTer
mq+Xs3YQTknhzyO0rfRbC1xuTX3Xfcn6swWuzJTtqn6HdzoDg6as9NbF5ZJeYL2q
PJUpTSD3nIaC/feWPTp+S0jLFrCp0jUtHATbsUod8ejOSUa4306MVgCoryn2KQ2I
BJJUrgJHk68VnojozKlaZIJmRzX70C+lu2xaYV3faGm0myIdES4LTfnHOM6dA4u5
1Zn+2dXXOnkmYht9aY/EUUPhHqqTj6t8I9lLQsmRljqyvbk/i6xeDO8/pPX5q17c
O0DvALh0gTSvGegsCpqlH8SDHgOs/HqZXN62fTqmUUzDC0YUrLJRoSOHKFHon7Pl
qck6W1DA1b+hAUdsf8wlEombdX+3CJlaxAmOFak0IrFFlXQv8FohHGv9iPJ3NmLY
CfydsgyUCmpyJZo1n1W3+UnqkcSwcorG9IUvgCfKPLxjBOwe3pGAp9NmefNkI5eV
PFHxcCK/L5kbEXvUNGfZ/uSJCEbqzmyGzf8nw8SZOFCexzoKoAKHxCmJZ9ARhqmd
DYGaytnhrZ6jjOdre7YfL3lnzAC0irKvf+4u2SdN3Lo0q9bsXfZ5yVngRgcTlTh3
m0hC8h4kak8DkTjJDIJDEUD58sRVLfPC29Kw0gGJwVdKMu/T4jSeTT8uVh7KuuTR
yZ/ohAUf9VhWeARnN2eor00F9j071YammjglVTPPEDLwkUQgsaNNvra/3JT3RrHv
6ra2ZHdpSq2Mfw2/gV6ICEqMTQpFsQOGMHj2u7p8fhErO8BS33dSU1kkWixgn6z1
4518WED3ji5R4v+41pARKAvwbjZiQJQfUFiF0AJzRQmn0HDwHYEPLMB3TUF/bIYW
h0BynmslE3k1WRvXkrTCNQ7ZCtwTb8c25h7rDZkvXCMOZS+xS86x70DWspTF/VHj
KCqA4JwSF3EqXkqSAWM4EgqobtPpO/H7YLuTKU+cIU2imwCGpRPDFO0srCm4AqHO
Z5cnhU5qSHO4W2joPtMxV/9F+JPonsX7wLHemnhQyN6rkvE4pp7VdqsLItSoYU+3
CQsi/U+iZbrtvJjLVMBRdNpCnczE+o4K2EADlKMUgFi8E4qOTlbKmIujTJiUccAA
PNDG5jrGGGYg9wmHr/Kyxdq0Q2ozOMMRhPuBOG8o7asE+kB1bqABD+FNB19J7cSM
3vEGFOOjFRtxqgJ3g4PgikrPorttAXWZlJ4diWmv27RiZ/RXGuT0t+5Ev28NpjMj
XLE39lcI3+yeBtpsLU5L1Y1rrRw2dVmuzh1zs4wNsGAcknq3/TgwgFu1erBK5n6W
M4NZnNGskmBWLp0a8JpMcGYhY+HlwOPYy6rvasUEPGX5uBFZwDbovOqK1NJ0rWEZ
QSe+Qv34pBgRssXE/Q1kvooQwlN353BGtm4EEb4u/d/hHiHKjWJz81LU7qN/abYv
Yq/scErj4qe0x80Vh2aSiDCNwCqNy14TZb2aGvyfMevGgkZmoo3zTT86tvSL9dlM
tm2T67cuqDO4uVx5zxyHCjQy5w44+3Ttwist8i+dDaNLMLVF2A/cNa+Q5DBfRcg+
OEsIDW8srvqDQ7db0mGqOoWsUB3FJL/Kggm1P01kgj6tmTxjowh7TWRNbPeAiycu
NVim7r6BjIt3tBnri899Ds227+euWum7k+z4grVa1XE0Z4nKc6IpVbDHbBN2fo9Y
MGeYa+FPGWN72TzS2Bq7qDhAkYfRVbw9eJ36HKjaHhBf02WR34N4qj1zdwPVhfBe
v7mijAyx2XnY8n6Ihv4xK+o2E5aL6V8EZIaF5wx39JhYF0JYQForATesB8F0OFW+
jE7taw7QFp2UmVmA7ydqe3/al8G3oaY3JDrPQtTm+HbXjhmnIwTX49zHF1KscWZ2
cU8/HSpil+ev4QXPciWRLtpMWl0MLznwTw2aincjnFMyxPd5XjEEkK8CWqr+Q0xR
DDeMm4JAQI9RnwdWzGVQaUifHJY7aeYSEKxN8OTQ0ymbvSaA7IcUl/8QNGD1W6ud
jDhHCysbvjjXMyrBvDMSUVzVXyQfa4ro0E947FWy0iNB4rwZrTWuWUZB00Wqvb1P
x++h0wTxotrdqCp+8WBJJiY83HTg42PBHVfFKXvp5bnblZoP8xod4hrB2bGHmdU4
diWQKyD3U0G8u18bhIm2n5UIh/YCWNUD4oer6RY0JEUNLw25jDyAUMxLKD8JYHy9
MjW7/AKpQ+u5tcY4yOUSiaJvmlRE19JllUYNeuPdYiZwvWsXM6a6wY1OnmXRT2u3
VpHGEsNriJJM1iLjv1upnh1tawA0W+PWILYUDbNaPHKWTqKl/2mfCS31GUZzXQSr
Va2vTH6KR8d5D60upXrJpnpXuxfzDhYV0AnRuC+h9d8gZ/1A0QeFekAqTLCicalp
SYqNpPqTev0+gqsnPjVutXlooQiENZY+2xMZwHYR7AUOb13rpVVPbVXyIaeQMAZi
bpA18t5DxgEe68sCPF2+Wy62qJz3hUKtOvPtN2GxsVA5fqgXotX9dKRasegK7ZBD
rOqABRtgv6bASBXvFtVvZ6SKF7fs5/FMEN4gWvRidtqHkZsaVxA76Vu9BlCcfra7
bS9X25jgVCLRFE6CYZQ5NdsD/83ecA18ejbhVSilf8eP2dNutlc3Z5KNx/RC5C7r
LJPsrYOB5Y4HkuDal1VN3zGw/DDVdEUEDUcgyPdMkJ6+weoN2QC3ojVuKsGNJHxq
ZQR838ItHeieO8nXy38HMs+U3tbM+jQ+JXDNh3Yhh23KyxdVdUdEDage5ZXlqGG+
80w5m6wmi+r+HJ955xc4SQ+sbZYgcR2ZyYattV8I8u082L68XAtSVCqmQkw9aiGF
/dZB7kUlQlrJSYYB79XzDKVIS6JmntS8Sb/hIkzc+9rv5C8yMS6MVan2GxNLc/Oi
uDHnCLbEwzp19ZLeRqtCwqTEPqXvrNy+7I0DOuAWJDvtZPvkH3eZ/oBlEtL+zoE8
RrCJnl9fGz+A7kw4Vust8w7UJnDovBjgyTuYF994Ao5EKsp06a28bUILFBPJfKZh
yaW3t5Nz791Kne3Z6Gl9AjJWB1i+0RbxXHj/t8eEBYUUn3BZq2D6Cd29yP6vgYcM
UeguZXxfWZ6DuB+YpQZNJzIIw7OUigz1evD+pRavXZhWbvcaETfbkJiJD/UVXsRs
s0tmwIr8WdnUaD6g9yKQZ+8sejNEifOK5JM9wn+IKWP1f832EqdxMa+TDcAZq5UN
hhB+dRkFzVR5ZM9mAKBquCabtvNvlzN5Xzg3KTUkPSTz0E4OpdHB3zVp+vtIx2u7
KUH4decHyKlnAOh+XPa8Vn1Knt4h/FvAyMDtu8yoqCQ84IBzfHtzco4lh7BZUdkr
w5yLgy6bCB3df7waHkdEm4oTn33Ss3rLjXlUalnWDaQk8kxjXF4DsbKeSCgn+kyd
LabvQvmQwygM0d8zrAHHToAb25CDJ1uOV6O5kaS+jEXW5Y5MK78mxbqF55D/9IvH
t4hQC7BsC1Cae/vWD6rITNSTW4jDH1KcB/21DVbJCbZxJ0p/Vt8ScJl1K8HdGXVg
zksHPSFBBLUgbC2kXGKsilNZUrp5+NoEXtZ8DK64Qr8bTkMX4I1UP+yZnY/GX6ci
nuery1nacxAQHSNkf4EUZPMe4dERH709QfIiELYfkVz2aUkbbb1MJl7nPVmecSoE
+BCFUZHYjgdOvKMtNaJ+SP2sK33GqOdGepu2B8bJH+8p0x3wddFF10YHCH3kd35Z
sbmYe+WvD8q9SPshFHL6MzbkKbWB+Gb6zqpvNuhSLbdd7HLJuD1aChlrKXglExAb
Pzmj7ZovvUatz7NbsW6/tyxdUKeufL/UbS2CSVOiM/YEodRD8MQTuHe3BTEKpdx5
P0137XbaNlQjlbss18dler6rPjrQxCVyqdU1gBVkShknflQIR8Rs73ULv9sm04VT
cPuYP/X09ijt8FQLBygL7qLk2yJTtDUi9tcOt+fyKE7g5rFFJTtuiC7+6bMZVF5M
anL11oj0PjxS/4GVlMdAWWC4I9AtSv+wnJP+qJWAQjg+QU0sSEjgX0NGlM3jHn9M
2NMpZ7al0rNdmh2S1kNTVttHSp5relCsj5ExrJEQc0D/JMPkuwB2J9UQtOkdXuB+
3Z0Yq5XO2DyMc+6weeKKMi995B2JioyzjuIJJtjXWvmPfu4zAQk6SshOo9DLV5/J
Hw18zDneFRgHn7Hd8cBXqwrbRZQ2FpsvW5+Fn75yOmZ/hmNFvga/6OuIXnIIGRjx
7v6dbFC8TfA3py47JjS7uq8SqrqKzguOjSqb2XbSYDKBMTzE86/43lApBI3ZjVMG
ImzJzZXDtWdKkRK5MADKXIm6lcW4qvYFUtDn/3foRIMGw0VFoMTQI0skrW6f3a88
H6flYzcz7YFNmgdzyEcMyRTIUWfcAhIWochncBHmDfJ5hGuEL8FDL5oFpRJJc9ZC
mRX7lCoh7SKv+/3yZiY6YZ/I5BqHP2B2MgwE+N7rSCHpi6oAmkW4vaahUWYD+Pvw
oEpB+6AOXG3MzoRMLK1cDNaC2BM2dK+UoEZaTMlZPr1KxiiO4ubOVwd+TeoRkNSb
aXepkF2tvtqWAPzWJPzO8cRK7+fGFC6t3anjx4ZmFjX4p34C7/BPXK/Bea2ZZrWx
IlaUFYZ7hQN3BYCHh7nIJWH4kHAvumHQk4ByiEuJmQQ/KXa+SQ2zcLbGtPg/RmnK
ZRNGpWxqtShwp4TJjn130ueWBbmBujsFMTTMRdslj+WKvgswCL8srl8uC3hY1zh/
nPqAyEpvVZjWYz9s4yHCYW5+fVKq498JUkSteXC/YfU9DVQxbn/sxwNyGc04ODLi
D9pMazWIWWmyyitq4zg/OWC2j+exgpYdbT8+CnELEQ/ShDaP1NlY/1lpZiAJ1GzB
VkEhLSiPIqw+YR7DIEIcQxTIR+VGJ007UHfG96OJVwbulW48lGn5YCKsS9iXtPbf
HeppVH+Q6+IFJp8NlwSBt58wFq7daQBcCUMo7s9g99r41STBMx15sNPOCvANTT2E
pyJdiRa7Dl9eIxi6AQ9E26HhT3PubeeJC9T3itVxi2xcU+b0I5k7tCQVewCS1w/p
kDG0CU6mWQeKhey4nQ1fDXl8gm23zb0yjchaB+/SoUMSfb/y82lgbS1AKixcV+m+
Q6McKKJ/q/yASWN6s4RPHBsKTmrHoHvje9k4/5byJZPVEFjbl0WmZ/W+E/RdQ89j
NdjqjNvh1cJmsSRMG6sUg6FapxrGwJgHXEA8UsbOtEDHXIvHXwBv1pLRrNlh3vM+
U2hVXqECHQybwOCyEOdPFbNp/vU8HJhIij4iKAw1QFjNCaciNWRl0PmVFHRWwFuS
nLrtDGTsR1iibl5rWYXmYsHGqxs8kvb/cqhXQzpyS/V20bLOCsbKkN4bjYq7cYTH
oDjH/YEpWtyD5ah4U3vsd+4bZE9ywxll+68klnzg7tEi5rKzqX4NrYM0A8coCho3
5ehBy5eN1nf8rAyF9Hi3pYiFnH1oWUbv0c6DWFXPuM/J35jNDPMa397x3aryKGW3
JlYlgTj9JTm5/9hoYehQoiJ+meHRzf/M28Mcz3yPf489CrkqhJ0fn+oUFFi5SMII
0LVcFnNe7jfGJdBDnTgXRXva+JOiMey3kw/DLKEoYhL3m713CvAMZyQgwJ7zzdeU
d1rZBkyuOEx+ptJt7+JPBd+47DSdxmx50/29R64BvXz6JCOjEoTSFoHAXRicN9br
ctum9MN9SapBhE9lj+MikJsW6jXokSEnGLRJZgE7Y6RFuPx9mU6w7BoTMI4I/8xv
93HGLaiu9PIUKYcZ6mU0Ve6FlcFh02w4NWH42KEfwynJMOD/pck2KkEz2e2XjoVc
qOcHti25woKfq0eeCpwqImymlanTjzcwqLGCA/79wMKFaOsv6uCNYbKRevn0MpKU
D0yyBG2cL6usgvISm5FJ99kwqOWsRQ0tqQ/0GvvMrd3X4QDT3vJTND7NuucpuQX/
xTZ1HSOyyR4v/3t6cAmbCanKjgW3YH32na5+IQurbqS8h49y0XubPjF8o/wqqdj9
tRwZfZGCf2wlDt4G7AEXR16dgNs486QdXxOKNwMzMtjztzD7XEzLbG5WCSkfGDrL
MFK4WL/ielZFIoEDERx07SXkDaMhfm4QKAxvy864qAT1wE/Zk4+TSqhM+/OT9dme
45KatRjEIuRV/AFjkZs6CrZ/5Dc4dLmqj+xJsCr7o9u6Ghe4xYizGo4SRuKLLMND
h/Pq+NVupL+ioqB5XNi6eaHf8d6AUFINtZyFZTPFsKj+Ufd1w5R/YePScR8a1S2p
HZnBzLZkl+uG8qcetj3b0W2Xd2EpgMVyzGIrjG9XzUv7oeh2FCBA1uzPhtJdI7RL
KSSXpb5Gwo/3alT9GE0U10wQKwUH365MPS1GU3PHQCCwj8ioEBqYaTTczyZrKDM4
H9f8w3gZZaMkzIs76EJqlILJ5dLiTGBhLdlNRRjn4tdpZuUnOKbJAEM9RxLoKdSQ
nTrwYflyIoVH71H5IWzDi0HUhroThSP3TSYWENx8ebRYazThzTvuFLt86JCEUnlc
K+Or5dIeQVCm+4S2X1Hrc/OnnfSpwDrt31OosCXCG/DbF5BK5qo0r7nCkGaf/mNG
gYXrTHjvzCemDD6XK3NI2ER052wicNOHpX2lsZDcPMJm7H/VVCw4rpPZnQYrttgB
cWQPMNhSA1TKwRrdhbIjlnYEJE7AtSXnYOM757ATZ2k1XAO851NQ5a81xn31+mkK
ytE1FAJ/zbgB1d/f8z7HaDJ4j6jZzPXS7juvTsCEPUbzgZI93BK3L0ZOCaWGXJQo
42EkuOAgVclTRl0hLfZAacJA8fILi+YrPxe+m8+nHIQ2tbtzjFZAyReaQ1R69pH6
ex08vWsrtPtLu2+XYzPvWnA8DO+Zz2D7HetMu2yvqrtWUyT3y6gs9oia8cuKNZQs
S4p3vCiWQavvSPjzJtV6r6ninQsWdZvsr2DFBbwp98RuUqNE5t/F0B4Rfjnd3uNh
+LTT37LmfK+UNc6nE4R6+K4boXpmJNYnzcws5VGcLUoqdUYo6FA5/F5nNDH4XsDn
aw4d7TTFaXE0XzPdPS4dOJY26klYSaww6ac8OI4Ow0mF058nf7lU8yonJvumQb8I
4HWL2G9Ty3AkpD4IGeFUX1du2XSjR/EmxV+LAweA6Y53HI4GFHqxGbsrzsHnqld5
wjMqRLNw43aYzK85TBOgfqI7tWF+C6GuzjmWkMLfMC35ygfQ5l+SfgKMbDWAQdcB
2vWwjKtLsj88TqDreIxt+z+K9O9vZMDx+7HRY5U0TGZWFCVnSHNDP/9sxMuvFdAc
Obv1rjuuGLZjAsu3+AcpSqRcF9X3xgiptfegaC6wiYYnnuUh6Ojl6YPgug+TMJFh
5x3Fu28Ohf6oK12G7svXy+7h3G+KuMoZfN1Q3dOXy2Sver39nJ5SW0LnkcQ66wQH
8rVTQ50dBpbqKQ6BZzqGgiTe6ffbqxX96loQtist3UF6DA3OCbJ7eAVurQiMlKk1
LJk3BGLsBtrV6L7dKCEJtd0TTS3S5r8hP8xoGyE4RMNKDE+kw0u8K8PDEDZCxmck
JUxKBZwBHzd/jPzIEgS4qIDbJICqg415B7j4e7quN++B8U5qXTCQ5mzkWW8oke9s
lxvtxcgJqzGP7yl3honi9ECdgpn9nbl6g+fkhnI0Z6KNGpfevDXjcfATzVhy4Huz
JZu1zZTZ7Jn1ah/sXH7fXfcCDvhbvjB+OZwurkUuBIw9VPnHQXD2QY/P29P4E0n3
8EnpWts4AHkk5FjqnU3K4tZ4D3TwGPs5RKEddM2YwYRSUPk2MjVTddzbTpfGIiuC
3tg73lByUc8I01FdeIaxsmWC/Z7ohysgVTBy/Wnf5enDRB9LKAdtTIksKVdNyEAD
uNof7bc/VBT8t/Jjeu0cK8XXtqpjY41qGSog8IX7qdMkifCXu0t4SeIrt0mTKsI/
ew5M4KToEqhnark7WI1kEo0ZMrfWS2yYC9QYKbSgGWLMo6q96Yf308QcSg5uQs0n
ia4JdU92qPSuowM2/iz2DgaiwW/QknrKfT5YCHaCklALuk7hVD9vIG0bsCvwCfJW
gkArGNE5zisIN5sbSI4vV33tHop7ycViBepREdNTh0/vfcFTRtUDk9nf4bsSEscF
kQkn0qwkVBERtRsjMTMUZ/9QPj2yIXJ+Ssu+fBx1iysH2x5tv9KIwOmZxCp37pZk
Mk+Bo0F/rQeAaxoyfKJg3hKAWprAj8z48SsjdkaZKhHRw1Luyz96TTpAN/GjSR3i
nT/GhqWAC53bU+rKJD1chwytC8dajMV6/asxfFgy1zxX/AxunTtFUo+anTJ7ZrJt
GVU2XPjHvL8g5qgPOqQ2d9obEcu8JIopGPe9MDeqfj1ATu4Q9mHcRYmwMRDVW7/w
I347JMnYrWLPrQPdPp70pzYLiVgVevasWWio9HiD/FNzDFdYI4wuOkSJ9bGUjKY+
kkhswdJfs3NmwLFE8sSIsd4uo5VthQ6c7YXfIiEUjD/HlcB5mJr2yt4Hj7hghk3H
ig3qL8orIha4R9Km1EebY1vYEl/rSMYyPso809vcpmzZe0eqQrx+I1+HfkMI7HxY
P6WM3+Ga425AIH6JDLBC7ygu0aRtGxKp7Faa2wpqpg4GfVlXRgpWoCgJhY767A+c
bgqJqw4RJc3oxcvXBlIyjKkF2uGRDVu0HSR244hhoYiJNr4BRd2gWHE7wd4flA4x
lrnDOXcJ+TpGjFcCx4FQMiWQ6Z8NGFi0gG4MUhT0V6Y9fdb24Hg7lvgKhAacgU5A
lhsRs1XIoxHwJPSXAl7j0R38fKXyrBxwCZqUhRehonMxQFdfzy7tM0ZlUNCIURpo
Kivtkfx2InyvuhkFMJGqijSDIb8Nv+1zZRNQ2+lvIvFNNSX76IwNyMMH7whwRbn1
3/UhQNjt678KIO2pvaan+xcedhGC/TAlryCno6CJH0mXFJXmZ2uMx2Oa2vKUm5fG
q07f08ABgvpm3cqfFVCksR2GUczRntu7JEhGim2KpNb2+UCtlr7L19s1+rTM/XdG
hFGdU3TUpgKCWfmg+MVXNcbo9SINxx6/GWYeeMSg7e+GC/bYAvkJB8NrPyx3FPhd
wrFjFfaGRnZNXCdUharXHuJjGVAxC2jvxc9KahOMHZk9f6j++c++5O0C/vTkf4Hv
JPMlg8LY2enKy+K1zlDe3AHhe48sgDsIq3kkIolrwJd7dfxNTUNYBjNc2GbBFSQ4
7HB2xXSzCCH5NFBKw+WCOdja2imGhvlVXhEY1G32lS0qUTUIgH7Wpl+AcmEEurgs
JNrArVOC7J9aRgfhVnFx11gF3fPT6DvAEGYf2dWJn/0Efx53UqKy5FuUowJHZpQD
UbeR3PjRbhh0qv22kzpgETr2QAx3zyZyIsfbmfkmwfCL8jqR8PHQoaYuUAzd9zZa
BaLAtbUioM/MO8ZmHq4KrOdAt9I7y2weYnhjl58uQ2EcSV3xTdirJxPgHdpRk6tW
E9n9d5vVIViSf49zoiIVBhCSdxAqRKpeNxQgGN9yeTSU5v67EBhPDFggNu1OB8JO
b/V737YVkvUQIbEXH2VnFjT6WdXyQ/l/iyipl8R9ELoqMIoK2uHKYTR3kl0uZufc
LJlYwNPdQzpbK0mf6ugKlyoU/mzDnMHbjf/AsDS5woczQE+Hbzd3yV+8hG1Nuym8
BnAI46R/gpCrnSj1r02zB7KZhIkSAndeldBv4tfRwjgEfcGftNXtOzwdPBpJ5V4t
YHr95HWD0fi28F2SIHRJhju+BJh35RfFeSc2wX7t7NPZwlkvilV6VURntPN4msee
ckWQTvNTjFoyHCecLZoWi8nST31j0V1HPhOfJ0lbPNDG6DAapFKra9SkC9RR5Q/N
hrRi0k+f0oMoObaHfBmQn8NPcIJsgLcNFHTKny8+HLZHL/F4vsqrdEiRLca8A+KI
nviU5S0dg64+FewUSJirbm0w9nCnzyejPr7j9qK1f1i9ChR2l0lHOg12zamaEF8E
9HFrUGfo5EjbVUQbW+79jwrb5GJNHI+FplFTbacC8c32KFtHlTL9150KUSSpoDp+
bvCy2vLUK/AHMoveT9fwsY93kXy/tQrb5wMBLDN0SB1BMrZYG+PRWCtSi0tJXbWi
t1kKCVIfFMHMLzNQ05SEnrH7NJTAvJVLUwmdWKBM76r4CIfWy42MmoQp4iAnKweL
ZL3esC1AkWX66ICxj/Ef1/OyW4NEG9+lLq6Nb35d2D17moD+mJqJj8P1qM2xqgXq
DdMNyPF+u6uaoxEgc2RO7qydzfhfaxpCvBu0X3kD39y66w/WKmos6PIop9qjAW3l
b8F4H7SDUWKD+pa17A6CH+z+OiXVI9kGnx6C3tJJ88WRXiGXry7DWaKQXFmIu/Qd
XsxZYObPcqPkyXRi82ULclJvHU4J3A1emDyCZu0b8ycnD08ew2al6XAe7kgUyV2f
0pKENFeVw2exCpQEYCpIbkmoQ3dZ+80vYr4VVV/0THpmdwsfdvzLdgKzlqdiJncV
UxiokRp33Fg3yaYZehf0O4xzLIhP+rtq1bUEb6/Ggv84ei08ALEpgx2SLGyXpNUd
XPmwIvZFULrwu3QBGfzMVqTJ7mT2EXTOKAM87Wq/68NaGrpyWv/l+Yym4o9LTFrI
XwjPfObEDsRsLv9kqbfWvYVA0sAwO1afGc+hkW56h5kuiJKtx+dFLPDtAT7VoEtY
t6l37DKeItajFG/wEapTv/nhEAswdgpznNYoM4XKcVutWpBaNBUc6L2q25cecwe9
KrZfFPjYwgwWeq663gKUn6aKbdbBK155P2aCUjKu+kE0Q8COT1C+auEM2yX5uGzQ
eqY2Gcqe9PbRx0+OMZEJr2LHkjxsgsaTcwO8sw+7oCQ6qpIGEEOKawBH28ln+h9d
QePXJxXI2cyn/PSyv6q2Ctq1S8Y1bw89kkkEgEe+DzFJHzFkctFKg2sOcQ1yEcGY
qu/stYi7+C45v4erqRU+cHTIy8lWKwl5oQWSsqJdkhqi4ucJXLeAqLctUD7ufsVx
OS35TX757AKAQk390zsjrPC17/fpFF0GYGr8UOugQXpWToVj8seO/mRU8B8yjwS/
plpNqDqJ00dKJUAcIVukPMLB/X0fE2nsX/EFwBnGmldloPAxXHTl5BsRQQXjtt56
PPi1U0pHeRSE9WPm/eneKJyvDnfx685PpogYtwvi8UCEbXVdGsAYOOXpr6w2Gc3F
xtY4bgijZDenixZLVB4Rw5X4BJmMS5MErgnDkNy09WFb5BKQz/UJjI5KdpIfm/yi
D6ZHlqFFM51RTPllOfvh3b+a3bLWm0+BKAjw5vAxk/3XDqcTrQfoZ+fYfIT+dsMi
hrfciI6dcApq6hLMwUFY1tEZQVgbDDufqt6jfBRJueCOTMGOul8RL9ibYyV9dp3O
D2KxDWXkW/e9aM67T9NlhavFV83m0jkQv6CK0n4r+KDPsOXEVBmIgx4oD+x1qs0r
E5t5mGtzxup9VYq/YFK39pBewWMYMQvIjfA8dd6WjYXW5///7KTnYToSGv6SGM1I
PAhEuL26B+18Dry0AYPhGE15kKOxz32BzK9hKisepN/TkP8kgGS9MzTboEpovKwS
x0nKEV8StUdwcnCvMVtegaUWoLK1rdSYhE+0u7CQXWCyfqilFqphYyU/LptCH0/6
vm+Yv5LwWC/qr3K2+UyocKvFY+K39sIO+is77URWmPBE+2q+TBIOYazj4xuX/8Y2
BIbcm167T08pB2tVdKqRVKaGez3o3eny+dakaH5btiPE7d/uq4Qi2St4180z2+TU
vmoXlfYV3lHLREx26EMQet9KGgYmF1+okb92vyIhRd9A5ETjOobVikc8MxdH+tMH
z5hvDhvMQTdMv4UrgaZfd54zZHECHnWljK6UdyK/VN/RIAy6mgrMji6HYpfVzWz2
MQ2/3zZIHPTC+mpzwmzWq1hJ8CSNcRYd3yn9TWqM/uOomKSbOX3TQw00julGb0Fx
Ardm231Mg4LESeQJFebghuaJYCKj5hIV5rbuWHBPi3UCutbUaqqfpaAtZcSLeSj2
aFR1H4K9bltBOlVGLh4SsKL86+FTc+SnfqsxY04gUy50b4z4pLKeCNLDElgSnf5I
VASCBJhht34AfG5A0PTDwSLQnf7RYGCiQZhSt8rQZaMfKANyKO7qpK4GNrG91QlX
wK4PLwOUjO0HqM+A6CQH+VatiZB+QxFWO8madCCh9lPuVJvUDyOMTuaqEKD0plno
u1hqhb00M+j8/xPXUuHrTCzf71xbmTkmRWIrdQg4/yk5UcY2WFEJgGDo6xSasDDn
jYfU96x3NX6CgA2f09tKmiJWU6YE6tBHtBk77stBsiaOFZK7/ujdvVpKduRDZbJ/
2eH+oIBvNpEtB+ZcYwj/fvBCgFTm1j/tn4XaOTKX2bJhGpEcZLV3XJxMReffk94q
3Y6tDk53gQtV5TKuANXZcFAl5L6snymq6A6ZBAt1tnZEf+HyDe3V+PTQ3H1bcqVf
8O16SiBFTga0Fk7jr6bpwbt84D3VqU6aaVF9cf8Lu82l8JAxuwiVka4LGlMNAnIq
yDCIfyZ4sBK9bF/oQ6F41Lhvh4FCCf8uCwoYqCXwmAPFuSutxNfNsqkbfjHHo9DQ
CAL4A+WJhzgEC/ZXp9HLToOBjVavGhuguXDz4thL96GNLcRPPhnBSz5lWFfkuUuz
irwlRa0Yrk0YVShd0N/yMzMlexcyVxb4A4BC6o0MFMfAMuszFWP4WaSpc1lK6H0A
adGLJLlRzX/wNXnqvcFvdFu7Y3t9Xwa49cJWeWVjCmOTeBHXawiI54A/A0dO4qdi
mLdpgQnuEQL3meMtNjkjGAHxE0XYMT7XWR6qfCVNCDkTyvysAKicF4Rhs3FGa3Ku
Tu4qlGxeCd/TGdBktY7e5j6PqxZIuwAsiJny0oHSnXCeROMScp2xg4WFOgK6tFnK
tiA40JQUsAsCnlCmz9EQCx4c3gINWNPgcDoGOBDzCvpfvttD87+R15NPwsxPMSVF
4BWwqXxtb3YnB7EdWuyxyFPUZFEd3lyJLVBQz1FrUrB2fhYh5WFSmQtj442r88xt
O7yqPtuvzOAUy/2o+n2CfB3IozC3cN+EG3rBMezaKE7eRAHHOMPNX5SKZ7wubC8D
NLvHYmzR1KPA+e6b5fzn07Nu+yd6N84B0kDZXDcthLBBnTMfprZby7I0RuBsh+aI
T5ozHeFOK3/pu2MlgR0ESB2o8H6iL8XUwyKv547s9Jvv/3CLX8jnctJFALbwpgTv
nDIbM62ZRmZP/V438RZAODkecEFuMvMD5gdo9f0t6tRylPNxAWM8YRjx6MrSs88A
N995QuiYz8K53gglXlkhOmyPgMe9Mxe66zCS7/zVWLGf1aiZ+T5m5Plbm487tpE7
2FHevEJ58BDTX91jtkQJb9+R6qiLF2tIvXPdLI/gwAi05qVzTC5NaKicqUiWn+vZ
KutGilIjWxszm9YVnUux6SYG1aG8wGe0hiPvg3u0Nw1bBuqctW6gHSiAsSTbWS5R
jLq8mUEs+R8jpvZOfWYzsYCfjuHSvvAbFHeDzVFJPe/FmCQTmztuzlopkRG2Qfyv
FNrumDoJLcxjBbK41BVyALIusi7Sp+a5QAk8KJ4jwgoLb/GsoSFra9TldsKGwSAc
xiMVA840I893RLgCXYbc/R+sgdF2d18IRHqmVZkipGltBvZk5xp2otFlPW5JqaPe
qt3svJB1Z8Xd1yHdFfA4+3C4sogVVjURDhomkaKz3KOk1AI0sqSP0hbdzjeiR8Hh
f2N3+c+fRtnSnn0Aa69huNJORj6ax7XULaRf+cR2oT01fItQjz/xG97sl0tFQNPQ
ptN54P3q/3pCDGmpIobIj0VRGOhBQ3RWyPdH6pCIFS+morXHRui1FDmzuQDapycZ
j8Achy2oFGy4wanlR8KirJps3DVIUlExjs01pF0O0WEgCg6aUfYNugg1uFsrAalL
ebPsU4ywQ1T1pcY55r0atSWD+7SA3cGlqS59HngcTUE466wFH3smbhNriXcOL25F
orayMi9/gD++lirWfTWihwF+sQeTydsnhs7GhpMz+hqzBnspSyimzlpc6T4iF90o
N1A4G291oHuNHBNwiCNu2xrpY9LyszXIoPg2LUFuNWY4Lgr3X1P719zfKiQtFp6T
h2qdQzWocr7puiu3z7zEo3AJryZYGkFrvbtn6IPznB4uBdsjyW1rhHFKCgCyEkNY
mOtY9s69LVB3LCaIdoc3z3NaTMbmDFfsHxHj/In+ap/FS7UQ4A8ZeMo8/zm/zNYN
8e9Usx/duMMaaQFk4d1A/ZML4xYOfuipmHpwjWSJEE8ikWP33zkjz4UzdFCT6qIT
RE4Q0QgqGEWXpd3s6sBOa6DR/xsBqtseXX+EBQgkwC+56S33n4VxM46tHR6E3eFG
j55HN/5Vz6ZG5mfOUY6uSoiTv4KErE80BfKJq8PufJeAGaYIptfR/upDdhk4rkpm
CPA0/zX2MY0sP6AXPZ3TE1pA+7lO9ozNRhA7PyPjsHKBnAop0szkwCzfAe0/YE/W
rQPQ3HzL4ltHLdym2QFKc0WBa4AlYF0rVYTCgmBSDc8v0LK+aG+L2z/Tcs5D9DaE
pUrqBYLluY2EdTH/IA86BhHmQSqG40Hgopfu6O18qgCkSjWiKeZMZD92d5I1bOIs
fmAcPJK1iQdu6m2gqxnumrQmnY3U1ttEBM+TkNCAmfXiGKJkgHgLbzM/Pu9WV3QZ
GNGIsjdKWt9Gc+IGOatw6NPW/BQjJKvPLr0OZeJFbkpQzrmHZomNO8Pu/Ki1+4Rq
tAjieyWTyTSR11VugwiMYRIxQdqsJO9INt14igio4Wd2a7qEmJmfskeGUNeTxkub
7ZyUmX0et2V9eZUpewSmvtwFiaHKUB6P2sV810Y/esEB2XM7teEbnIE5vMh+v/gD
DvMqYNvCBdf0v/rUjhFl6kah/bhUkZ1GiOTrETbM8Vp0PCmk8rZw9pVJ/4tz1YGU
8YwD06i6DuSwTBPsRdC0ROirgO9l3q/4b3EcDrBPxX40qA0A+1JhvWFkgwl8WhaG
43x8UUlWBca1oqJ76V/mNKdkQdeLj9pwckd38ahk8YokKQ3eqXQrCrYJ6N4SgLUK
QmsJxEnm3MJElkObCT4j6LHfH5Fd31ld1wIjR+mPqoyuMAYQpb963Par+W5WMxZJ
QwsG8GUpu82+kCUvBjv6wCsucrc/twmSNo60enFFLDyLBkPDuOd+XFVZ3qI2dRdn
xunijQxBLbad1G0g4WnVD9NoEFplXensBMFAlYl+VSlk9ozQ5x4A2pe2infZHV/b
dk8wh80maa5zH7ChWOZBjV/2COBNAKxkMWk8K8oAihTMjvW0Y/6jpmoWDGSy3uEK
lvAhXw3ng3iccujC/NjuUQ/ixQlFKnMtf+QH9owyrJ1oa+dvUWs68ZnvhAaJE7vj
/oQjNEtnOD2jrIyZQUs4VKuh76+cEnexzcvY49izsgeXdnxznBdGlUb5/+APiFYt
b+up0AggA3OI9rW+xvAPDAn+WYl3DN0geWaMSolMV/S9z+3U0+zi6yFWeg20Lm6M
OGTivnzyv/JHO1WFPEBL0oZn5CtdJGH75QPc+/jZGiMnupXPgGLrAPH0k8A1C61H
0BzE9QS5U7xhRWo8PhQg3DOdJ0pmVH1+31kOyXV4U+eQU5kSBV8rVXWRQIRcFQlP
+0L8GbBKX8UuwWIg5i8FeL8cHbkLYVLu5MMUt9MNiYG5eVl4uoOYKnYX4vlCPZR6
UoA2ni0wu4ZG+xS4Pk3gLQzvQL1C8uShEzlyhMc+ZTLLFLRGXy148anyqwbBZjKR
qzvBJP/WIsehUtxpVsugLc0rcNP4TXVOx0QRHMnQBhAVhP+E7r7OzyrfCATLBBq2
xdPvDjDOMyxKTc0psSdEnELUBeW2EjtDsKP/sEORnmyC65UUO+io5DbyK2Ts5AA6
Y+3K31ujZkxtzetb4YW/v8GrJubFofa9n5pUXCodpdoXi+NeQYv0t/oY2jDKeHET
+nCdBZ5IUlpHuZiNW1LGPFESWReoBf/UAWodxq1VlA3bVcPE+DpnKLEBvvqBkgZU
BEFohQ3UxrcEkjvfst8itUo7x5H7jP9fNxBScGvUudgEe9EjeMPGvGo/57ax/I5W
fbMUxID21j+1FqxoSC4yGwEcDM/RjQbJmCvtx6SqUQ2N85/yrRFfHI1HZSCnbFa8
ev+lLX8qeJEI/eRA3tauY1t1q+gZfxq/GDSJn2InDEH4PTb4Ni4NCY3M25AOeLVs
IkAqAG6sA0M6/HtBHAY3QTBF6rPTAY4BS54knE16rpUN2Rfs29ctxKU1EKPMleI8
Wl/wCdJoqsWE/gYr0QYviUFP4mPK2Zwz02D0QCHl1oBGOPsFGhm1gyXV7fYBaAmg
UOkXr8DlKDmHsX39jyHujmz/npdHECwHC/BctJ9JVxJAc7kBYxhiLAUbleIeoESC
q5J/m6471fAjspOJzuBnpBpNzF6IOwBO9My5rnZ5e7J9o/cxxmWsU79JGZ6lYbGC
rtywWn1s2nKh1a3phC50QAnvCYMtAGICJspfZXUKwNcpqLRCBBQBVfQAlt0aBeAn
tdEU8IxVujD3149zfRi8Pc8sJ00kThxCUHh4k8fgzKx7gB5jzLFFtPBRfRgM6eje
bT7C23DUXQ+Bt8IXep7zEEwaqxgx7An57YquVrXlbeXcto2i0TsEz/Ox1gPafVVE
bwCeMzD9grfctAM+d5M/tG2CebFBd/BBQ4n6pDMKbjq3nTVA5Q06EFopQBqzyTkM
VWaFUV/ojHO/KCvRpA4pNy5T7MH29t0Cl1TMUyRN39KaNPND4ooGrHKtyfmBqQaE
Lty2bUjDLASKT2ux7eAFpT46KZgcud90QJYTdKbjFWTwfT1lPc6MsXigBFYjp9ui
bvUjZx3UKcpt+m6heDMe2ODnLbjEz5T2SGQNwWDRy5FXmyhYFlvpOt/8H6e/IH7/
IU4LSD3yfjW8KEIyChFMHXzoPjdxoT3HR+s9l8tNx+x7sCMTKD8cwHdZ+xLBf4dw
SjkNB2DXdg/ZlH2w+PM0O9nKPgiEDz5QLCr3i7CyhDSPOHYD6p9qva5iQNkCV490
G7NL3Oh3mgV8KXy+t1IN9NQCTWeFS2UHtr6If3yi5eduwxP+uXt50tj7ES1gABWR
xSCMF9I0jSalhytY4ThZWnEd7UjmsSC5zIWXU+g/gfDr9Ok/oCYlTRXh8m/BkAgO
/gSEzxq7Qd++6mIiSDsdpTeGN8XJHjcCPL6J0SdFz9Ipn59CerWRpO8j/gRinJAI
Sf9eN2rwEO8mLvNIkiEaM+h23DpBwrU2PYWz7Msft52WqkbZUMHaH9I4Oq5L2rcX
zsexCHWXkmxCwhBZzYs88JB2nyGbu+awcjrDljeiL65gFaDM4rQM924kNQKPzJuF
5fwv1tnJ9NaBvFrpXBFzcFXZaEYfVTqtSjJ6ZVFHlcNVuOfhXErriQHD4MY7Zv1u
QkKqFfeNvn/bsGBk5PwmcSwGm9Vdf69buq4Zoxcr0J8wlGAl3QEFHx7bCr5u3Jid
PsHw+LvsXs+30JKYzjR+am3psy4E0Gfp1e0Jp2KeD67YiITmYgzKkXyIZFZ7XXEU
L1qaciqjnZHzfr0NGtoyrXLLWU+Xk9R6EpQL1muV6LLoaAciyM+tM1EwQar7aDFc
VcIWX1km64YX/KFBSZpmLXjhsiLI90kny3ywX+8nOqYiybuxDDZgo37EwYoLHlBh
WdNSuSGmQoe/kYuVijoVqsq5QutkKauG7XOkWiKyxXkfVIy6pIF+z2rc3hBqC0gZ
Z1SpG3XRO4K8KDVvcAOII09SYYEQRVmp9AQ0l64dCJxiUpQh72yQkGz0n2sAAc6X
/BknmmzNPkYLPtnV46Q+e6qF9FXhwc0JnjdP6P3LwTmC6izd+//Vsu4ru9OO+3xY
NMJm1xfdZrvtMtydkflu0+2f0NkuiQ/VUjfIHIB4v1wc+b2Q9CX5Y0KWDrfh7WZo
KcgOb1ubyuz5HNiBfluh/q+Z1yYs77cjEd/k0S7UHwf85lSrbWBbuA1bv8AlT4i3
LDQxnZd76JBuruyIOLCOqaQO5BlzCQwvINLPsgZ//+dK+jypLB0BpHg+s1xracGj
XEv83juX6XogMBvgqmWyb19Stfh57y9dOtuUNGYW7X2Z2fohEnqBuULsW+hXAT/G
ryhq8JRY4HniTjFaznJgGuw188o4nPnjEmzTl2scsYvCTAtlO/ox9mRrRNoapZrU
ZOKfVOvdp5AcJ71FCw/Ic9JJxf+O0yjePPGc4JkhXrknBzJEh4YmYjo6gpl0EP+E
C1x58HTU/rqoq80lFRbR2CXDyik4iPj9o3Vek4dlcgteOH4yZQYl2ONPDVgXtM+E
RpSG4tixtuJ+6Y26P5LqspaFFzRJmDpAki95cJN3DEpFP2HToVD0Hrdb4NT1HnqB
wJz3sk31XtsY1jOWScKlQs+fQnBmQbMdYoty5GkJggP5MskbeZUNyOqowr8GfkZ1
yfg2B18nVeY72atEPOa77nh0fqf8zsmJHYsUHr3jzMBzpWJW/qSqZITCY9e1LcI9
4Ye0nwWQ1xdih2y4k7zh4qM+QaCtkDasf9zb9yOMj5THtOpAbz60jiQqNKlmWaZA
aJ5HmYiFlc2EaZMI568S6Ruev2wJKsOAz8GMYzzrM8LR8wmBtWm243/IXNBzek9H
hhveMGoN3CGBJ0ZMyeXNqgU6lcq0h9oqPgnRkhKphqJhlQ+fEOWBsPoEJ0TNuNwR
PzX8SAniIQtFo8YXfp6JthjVlPmEiExVoniqc4IS7BGVkPEdZZTgnfy7xY+nEKSU
BtWkGj0eMndWpaMFNpbfTzdxLHRTaDpE8lgNlAc5lmmvnzYIkQTCgFyKo2YK1lJU
2CiaH7j/QE+bqggOB5Puiooiy5Hg4pw7uFUE43IQEFa7Ne33OEGnCjgoOVoNg5+v
q1XFZWjV7EwuiOCU1CWIBjCN/wi3WLomKsfsLTppvV3LezRmh5xFvW99vOI98hXF
J5Jp2580FXAKuPQP2Cvs8Fep++Exbyd9PcxxxQaNphB/lP2vFFQWpS2SRW1QMFAQ
M6nuQ+EYrePcWS748LVwNi7mQsRAPNDF/1oSQhiVgH2DqXLySLTcOleIQgVhn85Z
m4iXKm6XKrvYYszEurkFxcRi7D8n6tk3Uj6q9hnVvQ7vC4yEWk+49T8JU4LIp5uZ
oNZaTG6zJaJVkc7HYkQyvqlXqRB8VXeb2ghEXfMcdZ6ZwzNIvtjGcTEaQQenea8G
eiT62/dP61yoR8oPE9FnzUbKwCSF/n/7tKfAAykrs7YqnEwKqz90JOZIJU/CVdkH
f+UzXRXIlXeFg+dGNY2WEdQDrhLtfg0o7sLuepswU16GgmzXJP1nRwb3sAsfjj2l
NZdkiBowyPgTt+lnW53aA44O1UfcONkLMF1nZHTV2y/zOlSIephqvJqf/g7E7v0M
RaB+Fg1Sfo+zzxu72v4hlsuD37dbTKyZPXejVZlDl5LmiVi0iJiI2Wx1zPqAzaTf
nw8KgrA5vCuKJAIq6n8Dg+2MjIdIluGB7og2LFgzzeUrY4B8GwR1C7QtmrknWg+n
1dVC/OCoA7qmJJTziGfW/sYgcbXX44lRwfAaeO5lyTT5CYpFio26WKcnoEJxsXtt
+hF9GwBynAI7FvTL7dvimkQ/xbKoT81p3LYgwenmKFJ9N0t8uLZ/TdgdV+4t3KrZ
wPr/qgwwORGw2H14Nr+Gm386g9xjgI1+dx5BmKuwe/W/yBuK7qJYitha4ctf6oee
lNFGwutoZq0pz/TrHkV1+VCQ6B24ebuJzLHAfxABNdxb9xjLqGq6XC3nQeFNBpWU
p1EmBY2uyv2PCwn3G9z5mtfmNRdy+iwMktnh++Us6Tcu4Uf72QH/DlZGagcqeXEL
2yqiKJbNRrjUiBjfniQYiSPH7MYyCcT22w45L+PUBYfxBQHf2g+dDWkMj8ga/ztk
Wx4YhA3HdkqHWpaRWgEC5m2EEIPHSNWcDv2YRYQH32L9nT2z5ngT6mIYYINhAK0t
3nsoM08u6CbcTOdit3Y3OlgEZnf7iV9zoct68gsMpY+fus0d2MmT+naRznVEjpKU
M0CJydn19Iv20ohdf0FZTmS5c7oGVQvL1wmoTI9I9B32oaUBlD0KMKNKfAXyV6v7
CJTl2N8Y0aAlD1h15p9ko9s5axponS+jienxsBjpaQMOanYgMAbAEudQpo4AfFIj
zTF3dzkd7YUSeMKIkmuYAbzGNpwmXY/SFZ6/J23D7LN660eyBCBXyRVPP2lJdw94
gZ4Xk3pr1d7YCetjWPShIUXVd//V1P8v5GhQMTjCFg1aPHZvHUxSVExOX/EPKKfW
enV22KNV+skTxKIsgTJNvhUy2G4dV89SUuOPZuJOCxO6PcLFKrQPds08zJzl+1C/
iOu3jXnu9Sia6OfSOfCVLt9eQc8uwbUlqBw6kRSyMUMwvae74BbAtqb3NV62Z6wk
UTgw/qTcCQHsWS3RCMfcgCG45jUJW+GoOm624sg0at6AMcr89+u1WFobIdySMnYS
eUI/AhJfv4FPd3A9P+FRQ/NMuTKxQ2nIZ4PYalxh69f0eHGDZinLgXaZrPG/l7JZ
pr5WTpEhIvlMKGvFtJUpKHWnNPdTR1lmFVVqSkrUXRCL+/yDJ6viz5JoRt/3FLB5
Oyf45VLW9MkgMmKfxm3qsKW4lRfuTZ0AQRJAIE1JEi+BFP7cCqvSIl2FEXW2DCo9
SjM7+yxqZAZlsueFfSN+hXcsZ4qnvOhTw1nKr/Zh5zhMVHzFgfT45J1491xKPtON
ZcXkw9sCvp15Ls63bFtqshhbVN0ZZ37Ro9qZyjPplPBduCth9EgCO8Vr1MNi8ttK
ACy9x3Ir2Mkoj8xfmkCJq+BR90NMVcck+LmLBTc+zTi0xVWbLeQ9pTme+XJtIAER
VAXmp6g8UzY8HBaG1ZhcABql/Zq1ue/0QK3zbZlAW7JkpyFusSAjJRSspctMvKVn
5ZKfY1N5ZyRElK/p7tkGWqmCVSTpjRrxWLXRUpDNhJwinAXmFWIcBnPg+yHKq3xX
s8OkUTLhqRSGAF+5eNLr8VZEqkcprvW58m7p7Z8UJ61M2z4iwOvk5BKb6lEYCRK4
fUlgkheewStnbI2RD7ng8mhfK6wZT406+vsHhL08+aBi+SgOuiRwfX70LEZFRLqA
01jbtS7mnbVf14pRWOGhMH3mJuicOsc3FsEjRnpJQ3Ow3wA6GpduDbfFP18qwd2x
+IPm3zaIU9M6UmVKfwrccdf6ECJ8JlCAiwmcqnD8YN4+PptYo30bDn2dHjTlMGrj
R6J+s1x9yT8dgRvbYSHpL/5SoFiSohz1/NDsoyF69iaza8SnP1pqNH7RygIcfbBi
ZMet4k0t8EqYZyTPoFN5vDIBoNWb+9V+jqBxPt9zRCkO1RKNp8UQ6ExsPiKdKWV7
a9/9UOkwhcozZUIoH3RnWAFmAb5MNRQDlY8NqDjM4RY7J7ukhFOv6TGJZyZwy2/k
lUCnNpTNPOXG0btr9YCrPLseKyW+pkbY/X2PvqIdk52I6DJF/SAB5QgrX3w43+rj
tz+37I/0ihQcycJDLRmz9TCIPMy8ytzmqpG7LU4HceLJGTCpi6VYv7XIhY7pC6LU
UtBiou2hBkKFFujVnvsPyAbJsY0r1IcSfkyM/NVYDXch5fCdWVkoyokYtZVUBqp3
f412tyONgCgn9HxKMM9iGltO18Ho7fvMYCQLPnb5TCS6vn8LP/xk0PwtYnAIRJaw
IdI4YaHjo58DUASS20Pz2Dy/Fz6e1jDLOajHRQKAOjGdr+bdqKnuMpegEdEcXxxK
4V5Rt+CK24XhaDU6qqOazbCk9DJeaHlZJcyyjmVIV4uv2jmx8rpkTLi/3NfaO+/V
lV0hgcD+lpmjuAEXz1fMioLjWEtsr+h4eo8Yqvhwc8CtiIUa9bjhy7/6nKf1rQXM
3fHFVrX9zb0jJnxPWZANJdhHIVfR8KFDs645odHffWsfcIKkCUgioXTxg4F7fizy
IfQ3MRXUoaCWRZYfRu9a0422HnPQBYsBb2SJwW6wgSB6ZHQ1aNdAknI91pWz5lYP
CywKYXPgkW+Kz3WXLni4EI7VeH/ffKDxrhA9WanD5jp1Ba22LN2pDamzP4IWwwF2
rO/MoKz8QHLMdxTsGBUKunkvyB9UDQJ3L0yoJ1xHKpo8iszbKVyDkoHSoYn30nG3
sbj6LV33dHbSe9Aaq21EEih8kd7CbveXWbdiMtoQOvszZIhtGDV/2J4TwZBBVX5a
zEGTuWs7N+mDG96dIdMcN2wdF3RDKy7Qe4KvuSGKmbCTnDgY/if0Te/hMiRZTTs4
tgR36q46bEjj+tZkKGc3/dIcVDQdW+dVG+Mfg0jubLY5G6chqJa5awmKB/0xV2Zq
7om87PggsRGJg/dXQIEpCpl+2ludiyomVx0oRiIiA8pNTdHU0WVem6di7rGAV2wy
n1638kSvT+ujaa3uULfWcK7InzJnhCd8lMZSBFF82PdCjKcWMR0NukCrAjbGpxez
eJvvGY0DdPe/79+0L7x+wd2C95jb/cqhl4bKiKg4OY5fDfOAzENW1fDyQTyInzZt
R3UmFel/PVyLCyl0GRTNm20OfaoqCOOaZLnJtEUg2Vu7baGbIXI1TeddaYQVbg6q
kTvFr60DOxkpwkHEw4hNL/IIS4VNvPbLkJo9QtS1GIk7l2ih77t7llJjP2OVmn2r
q95o5kJuwWsWE14a+K+L5yZzjf4yYHMEfWMWawzIDUVWV91kXZms5Es2WGY0bgF4
w9A74wQDDhXeJZdRhfy5m2Mofj5ICjUAbjm84VhIJTjMzgQ/e+w99MJpGCDvJpDc
NMAKBHfYVvgVymE/jYNG63TZsN5Z9qK7DCWGzKwwgmuW4dXBpkBG45NSdcCHQ1Rp
xMNioIqgipc1kQJbZU48jKO21x14L3sv7ovQrzzY4+rAL2wZQ4iXFmAvRtSG0qnl
r9eLK6Lb7gUYWGz/pIBim1xXahh1w/I/x7gnH+5r6ygkBAkNoU3uGZTKXtPdRobC
8avlKyLzzarwpbkmrNgl3NxFZ+3KzIAll0L3C2H+mBPKn91edxhj/xC70CGvnSRb
1UgFKju4TvCYv76osAxNTeT0k3Q8kfCR6ajBU90xBLQUKZ7119s7VZZEpwJj2Fv2
O/jyBLtoAltLo6NI9FDq7fxHH7gtXEGlg+jGiKfuZqPWU+JWbR7Aki+ZZmtcnbB0
1XsJacFFYrKQYFwMVgHXAFxAhbAMVtQL7FpAQg9GGJDJjgq3xvkKRmUgEgQ1EfR/
1umUuokiUAGT1KpxTBQuw7c5xYlwD3fNUVIy2DQof30Wrq1JACPTMzZYg6QjOJ9c
I4DKFV57EOWHJNk4foCo8di7Ncx2qTrvp3/u4Ak1+0uC6+0jlb2A/yEDlg0XDJUy
eJPBIOVkHX2OP+KYw1n/KluwpJtwmAhwBcC4jeK4g7rH0/5kZxBFnrWkJEazKEH4
64QvFLYtSiWsNGnuSpGe3LqVzVIcNRce0WDBBzvll1TURAXC253nB+j3FjIFzGQC
hDrtjSrI/SKgnclOEJ9RogkqZPgxBTYTu8POdxymlKypbZwdQA2TXJOLr913e+EJ
ZZ7dYHgP2JihwFzwQcWGLSvaVWc/xhQObCzAJpc4XNHTsq6XKKFPQRnB43+CmBCS
2W3F/Vc2oztFVRJIbWiNZ5+sxzpTMadU4pLlwgMxQdhthqK6zmKZ6G4QVXgAVfgZ
T7AkKMG6XIHWgFhEf10Lp4tzhwv0slWwOl0if+jwwCrO7nLeFfOctUipNKWrtmmT
+OkDodcA9BqBxG7hHe+z9ERdfifWsXzr/47W6VnneHMZdEUeDJwO6cCqbTpl4y5/
oefH0FNLz+7ZtqvrFbXy/4N9cImJkX3cNG4V386SJo+PZz1iID8/Fpg9pjMkSpkT
ISs4wUgWvqADE961ojH8d0JhGG8ZD/QmOQMoryh3d8BVn9xPGObajBQX4ZB8pv4c
z4/HRwtPM0FHKGhmw4qCMDYfl+laCAJpvVT464+qq7bj9sDhru3ydcYBOrvRXvJ8
aRmb3DPMdc2396o/8SzoMtiIrafHweYhrKfBjTqv1ec7ZRzTPaBYqsOHlR0ta8Ag
wmAPEkhRjljaHME1wO2HZWK1/yGIRTwZMYuQdgp/dlJEY/XhJNUW8ZzVzTnc6LuZ
k8d0A4CSSN5lYMWssnuhzMHmMeH8SYUs0yTfTXxTqLZStxresskmJK3nFWGpCtuP
g/+cSqjl+eb0UExteSYqkwRlhwrMwJFQl9YLhzR5fR5I57tt5qXRmr558rYJcX3J
pp5aDGdxbbIFwEVmWjy4eAAaTZvNfhcrAf33TSgTil30768BJbMoHxjXV5ftNvhY
QtMU3F8dM8ZOAu4DSpXzi/ibv+Yw40aUMObvOXh1t0m0KhlsEJ7pPZ5Ddk/0kz3c
POARrpurpdCZ69vc0IUcQ4vDIBQfLVoH0LyZeQTJafIrNNT0pFhR4+3LMqC6NF5O
a1LqWXgJsqCJeXxbig0RD91MXswJ38gZvoI2DPdgHdLrwK0tqO0twLZkyPSxgxuv
FF0O7sCVAcQBlfsisnWUmo9KqpUV+UskiAVMbDjF2zf/dOGtTTnqjBjcnB6CKfl7
td6cR4Wsb8JxE3h+KJEtlOLUnV8hOTnq5KOptuvPacrChxcuBDJ3ZowPkeVqnLXb
3xpOhsluIyWYk4nXS78+66oWVhrmiQX7IJtt1evaKl6yJUNq7jPBIdmazLb+BCPt
o+qbiXJ8xjWsqSoMoaFomm2cq+k7pBFaY11Vi9djjBy3r+m7TGGSTXhQDLvqXuXg
Q/hQlSUWZuMwHha6J9vHsrftOWQz0hAvQrGaVsUVUxX9WjLjzPk4vjVkvOZaZWBx
tz3YfyLCcAttNTBeRBvQ4vU1JvkXJ9N6Jo9tyl3/UePrWwpmARcBjdOuWLvi4W/z
hj0+e7vlf1gxBuQ36L12sExiJenCBLbl/3E6/qe65dvhEbhksc+LtQLpL9qkSztL
t7dkaYsyDY/uD8yxGBq0Wq+4eyFb9mlrQrnCgQWO7gt3xYSyj/fb1ywm5IcvSXLy
NJhNAkcHZt0fnyv5Y8QIPDMwHq1Y7hA2i0WJ8U8MqbreoPmA2IMopDe5euqifKXD
EX7K0aJ5HityGhTpnlFrZ5sZGatbK6GGVpXlKeUWyJBJ3VFLeW/fiGP8RaUu/uzN
8lGnaa5xd4t8Ah5xEa9hDCDeek3qqT41hzVThFJg8xsl/F0aYVNcKYI7ems9GdjM
r5G6Cd0RYl8yrDgbAdvjekv3/K7vHA4XTkIHnQSMeuEOSjDopILhaclPGUH7vkXq
6rGlJfMDdfqsREjkxNshWiJHCMsI+NZsifaEdoWBgf0zJNuRGuxIpIAbIQkze7hA
XwilDWtn3gGinaC9mere03koYXTjZzsxtH7Qji059L7LkWRkh5Mm79x556gKoyAf
kCu4hfu9RZ/C/J51I6ErWXyi+/jHXo7sE7kBiiYn+MDRHS9Ifk9+8jY0NiIKv/du
8FAkpgoAjuaID/QvFRWlkncbu798X5yaMf/NJFDrNLJm7dWIHqyCWaJiZD7s/SqH
AmjA2b3pRuDemhhdJ6FwoNNDG4qtA9rw5ciZT3BvZ5T0nwfK+pLk4H2V210l0tRK
Fxg6VX11tbQESVdxMagoQXPQY1iPso7kk05p4DktyS4qV7aejiCVMrrMTKmp3JeH
4KIOGS4ZVtR+MMVoBzrfhadbIRSRwx+oLweB7yZbikQck7sXlEISZaJlpfLDbHqB
86+mGSnJYxIEET0dpYW1TgUFAQnjuF0sFwh38c62Ukmc/AQiL4VIoiCypIJ8/LpD
bUZs2I6i4hFFoRUrRf0tSUwcl+AmjI+ztMm15kHk+sBVtvpR1EfRkOLvSjZWPrZ0
394jMx4bPifEzcqwwOUepyyKOZyMQXThjN4uu3TzPhNINPbDaBMZi6Vo9vasa7im
P3XwbUviofkqcFQV5NV5RH7A3gtUyc6j4h8H3MhvpoMP1RpbiuAWuFhfWG3P7k/G
YDwExkcgz+do46Dkll6vD1DfOMt4D+I+sCRTbujDqb4umLA9zcOdoUxeTCBaMGS2
d8ubdR1y7kfB1Jxo0oFhfrnz0i2jknM0g5uc+DOQ27GGdRAzbN2nIU01Gwaj1hxR
iXs6xzNqAKpUWmQ+zp/vHfbMz0xSAr1rOFkAEZetg37WaQxBj663BsURw5be03Yj
HMjbrX8SS8mFo6+p5YjqMmRjaNxkg5BqhDIq5ofGzJ1zequY5joWoKM1LI6Hsvx/
8V5UkmXD79rj3Xyziv2RdcfHAL9pDB9bIRLD+LcpJxM6Kr7d5muyzn8EjxEvd5NI
AjUhrxuhB6PXwOwvDwxf9WTqDMwLuO+dA3tJCaj+ZEuYkDSVO0iDR/+3JfAzVh5I
/G3+2E9/+XaoYn5Z711FHRtRFFYlTegRrDN4eWEJCieVwSZS7sgOsEMwLLZtX61H
K9epxdNpTfQOzhUaSaRx6N8C8YlwXmmF4eS7l+1LJ4qps4fEsWxZoSRZ5Z37CKZn
BTrL44tYkUDQ0/LnL64b580gElVyoxDgvixNMC1e3SxBoSI6czdSBWLaIaQE5Ij0
zC6lS7PBc42GUxgB85OdsO+/fm36ew2C3Ms5a870p6mw0LMmnPedkPQOkmR+xXa+
BwHb57GcepDoZsNGgvP6IdFs0iOp3UbtrGJYwKdbk6oipF5c3kdJ7OITfeU4pGdr
HADC2UrRNraLq4nx5JedKxnY0F9MHAmUbpPDwsbM8aQHEIUNO2KVNRXsPRpXxGi/
/krsG153x52aghwLEYX5SZaAttvtLbAKAgATejk3N9tMMW8h5xfXqKqv+vokp3To
OilGB8nkBiYVOH12lslRi/YNtUc/YhdncPqe2Nv/YKx4EqFhgGkE5bsOoxJB+7ai
bmPqkMhdrwISpQBqXY2qIu+HnaG9QfA+N6IIhb26rN4uKQwtcnS+MhY7tfUE4Qxd
Xny3VtPIASNfGCXC+HIFbFPizZuToJa5gka2zsaTccmK6LJw3kGrKOQxjpJZtfCR
sB0o+JSrj1UgmtvNaIBhYErygWq9f7AlvSajxP47sfes2Fm2OVAMfHaZKXtMWPuo
e5h/9a+BV4DWalM0GROiZKwLghRFKmIu69PPe79GVOFp+Ciotz+137RyOHr/pck7
aOBvFiTieRK7iB3C5Uc4etHtT+wszDPWlIIPy8ZkBejhsyDlvMZAMysPidHYtRjv
W0jsR0buyK0BP9NEzdzbTzgIP04wCP6R5r6Ikjh1NySSp7Jnf8eJ/ZS3b4ckPMvF
C7bDjmN7Nytm3F9Eja9//MtdB52d6l8zo6+42t900gBDiyYUqO4e2C+jF5tDiFMz
rIU2esPtybbuzeONFkGP2u8BQn3U/NDGG0vVlwlihRrTs76QVJ5qoYGQXfZO6AL0
2AbNioN+jya6ACgAdYJnoeukiRmyQ5rUT/fxHp2fxYg2GjWzyc+npAFnXKlgcvX5
jsvOYDokVUV2Lua2gUp5rXtCNoQM/ep30E32Icl2c404GhC1uAl2u/rnKGBA97CY
uDODbjpicBeucnD1uDj+3tBlFJDyH9MPsIzEaE6XI1Fn63YhwQS6VuCD7g2cRP1J
qLCK9N8SQqXbcbci0rxcjFpLUm3WCM4uu/H2IDVkWlXabHcOOfekpcARyA5BUt3F
pKQIYY8gWv8SSGpuEWYfgY+Jy18guXebgzKMklw86B4uD/wLggA5oBq1kmFU3VBh
b00o4eTE/Cmde/4F5Dt394fWTu2n/fBjGYHYv2ugPRtNyyb/R/MhiijGwR9rKml4
gS1M1yBqGPLHKnoTf7uiNcgwAUeqghw4GmLBMKab5h2Eg5bqUDNBmwdaKI6Fvyno
KtcSuvCCma6EkWioOVi1He2Ty8v1zQJiO6PLHRIcbN8VMINxI0QoBHShJLV6PJQy
0d0+cX268BuyblssXSohu/Hh31AWePBJUm2cfoLT2FVhfRQ54reisckewPP8HL5+
D/WM7QFF5ul2uXRDZ0T2oty/2ZLMLwf8E6Tvf3z2t4KZaMeSNR/E5F+5Dw31ZZC2
09CVUXkSpnmZ/bcXUBW+j7xs9rUzdfndJbR0TUhOhE69VQ4GEA4rgFm1YNP0rwJ6
g8+B18eg645z2UdeF7MXEbQ0OclY+tIUsBqsp/ef6Mfmk3Dittn6TZj5F06ar4qG
jUiXcsiQnAj83SRIB0g/8qy4TRtoUS950yxQ6s0xX4cgOSxgmjdmXxNStwKaS1P6
S9bCgZKi+hMZQVw0jcGcbJL5+3ILe5ks+NKFuEQrAvNjeDVOeyqiGuqgEUILH3id
jFsl2bvLyeIFEPAGap0+dMd9Ijs6q96Ftts0kBT48vu8b0OJNFqYy6k1c2vdZ21T
cKRQBhAMIryFNDPOfDhdiyASQ6NDNzWCR512CjNrQvBw0PSnQk5xldXyQ0Ff1Ng+
0+tQp+1muePjMV3EMYefa6+j6gXi0hrDD0yuSbpRPSCPJCebpeQKDVS0NpRo0CfU
GZmd2FNzYmBTf0mtWg00XZMSLE13WYSas9eq/PydYBz9YcRd6XSZ9qhqZ3FZRHta
EvSIpaG4Wy4p2Jb2SP21g1bJIX9qd4dwMJttLwWP4deV1fmLNDKcgmu/qdObUyZ2
GOxKph1WHwauv/SEIivCHXv38lCFPW1lqYyp3dzfobi/td2eFEI0PXvfymeQvU5I
L5XbF7SygzO2Clg/6eUq8Jtv6cXjPrUVmwZObpkjWgsBsY8P5tfbXjb5zBBUOwj7
YrFQTQ4dXRBthGzIUkpAiDLOKfyHFcYo4XcuqpQEfe4EOsBZJlFmbOPO1YMUjOjn
sEfcyg2PYtNCkjOwbjLlg7FIA6W/bLg0uGZziSkUFQ7hBymozps3OqnE/6Tf/qd5
kQXPYu36Tbu09U6tJl9SZg/vk6nLbWUfeQcxDDkcTPiedzxsZYQtzO43UdCOXLoy
UlhlTSFI3j0B1ZCuRqCuAE8Wt6B5HN8e27I0vI3JpTYNFoYnVTDSVF6aD89FP1/h
hEQKTic9M9VpRJXKFqisqh7EuOsD895tG+RBaIN4VgNDYZhHOLIdn+7dJj6ibMs6
LRAHEMiAKYdN6K1gaqo3ts6k8w1ppvWuTzLsoYitKLOWdntbVt7Ehlf4pfImh/Kn
uha5INveQ0vK6bVxTLxLr3C2vothsbhYKgEI8/lkTRTSwXa3h+U3p4BOPZ9cf6Pb
yXlQxczDJM7J96d4h6R/K8forNzaqe31EAyLN2/QkJbmBq736JBHj9AOQ/RuAeL3
qEMhzkCtNESPX+QKrHWgwJ2XZdJTfmhjPD1W5pWS9mgadEmowpBIqWHoFWLHoUMS
hJAFcsUoH2EIhI3QqVk4ZIm+kI4iPy/zpYtAn0CgvUbWm1x0AgBurtALHC6Ks9gi
ulSxzsQd0KWaTkDm2dD6op/oD6C0x8f4AlknL0OEJQvhmC0hc7vp82nS399SS2cM
S8QUR3ARab+YpsePhjTz0KIdBw+0aZFKchkKxFT3QPVQj/Zp1y38b82tL09t3OeN
r8JKxIOMIYUiPY0UvbQUUlUoVpAqNBYtbLFNxkgqs3ahu6RSjFeKd7Yo6qPKoSDl
ZSmDq7Rsy4tgVpGj40KuYYbam28uP+iAZIJevy4lWovp4AZzRolk5w2FBk1o3s+7
9NUrZwThzWwS6fy3hrsAKcDbd5wVYKjrW67eHcoynzbhtKEVCIaUq0vv2JVAJhgB
ZKj2eqcj6M4bTLB81bsL7AjCKTHlHhSYOcEN80rno6qzTLNt5h94FNunC96cDEfF
MpMwtn1wMnM0saYDfKUB7a9ooCgJ2O2u7JFhzXQJ0QrhU/dHRgGy2r8dFlFcoFEd
o9DWnh3HJAdtuva1QBeXi1nmaoP4GhnKEyfIBL6/OKpr5Bb2ZhMnln2oye4HnWOL
hqzwfXy3M50ZidNZpGZvby4ExCbHZofh1QGfWqnrTKC8OuPH/CzHZ+6NipHG+ft3
M8uTbRtPcluZsfHECBMpqUDUAu9UW3SwjbL9f8urJVhV11eX9kXSJFQFTO5B8w+H
jvYa41VYdtbUykTUQyW4mvR8RCayCALpa9plb9TDVnk7zgpcqsFvGqbndfFY7nAo
a0r+WpV4bvJneXb8Y8JRTYVyNz4J1Df2rH/FTvwTgIsnhlkzBSnPWa3nFYyl2RLW
WqWQ0BLDoPy8Jsbv2wTbUOng6a06ir2HhOV/306JSgpFqbxmisUHfOINR7xGcvNP
f4+QN9UuM/fP3EmY8U8tI2CmXuFxHYSGptmjMTuqNx6J/i68eEQ5MP/SPSZhYvFW
G6yitXIfx/g7gQQ40AIXgPq8+RLYuwL62B3oZ0xouzMYISH4tcvOnl51aq+l5izn
ldkVAGP46hXF9lG+WRv1oUNqK8cEokOq2lqprGYtXFDoZ9M32jrzTs6rBnRezV0h
NW4KcHNMdji5NsLE2Rqoo2i0DB7tNF2dgAXLXABI0EQqI4QXCZRZdqt6nXXm8SJG
oaaJI/kCSC+0mkSXRHeCkUYdGku4+T8wg/QbPh7Ka6K0b36cmqdHRWnTOWVrCYwU
pwzAYUEzsQW/CS2ewEBQGE5slUwDE3p/aNugpfvrEAwONpw3vA4REFQjlhNPpPHw
dcQK2pL6eHMhdBnon0oqA6tZOJGq9rF4Qa1Feibz7TA93IiZMKk0qMna7F+ECaao
gzf+yMxWWHC2FGckrQVyRBkFsG32/jFM/iMvREhP+Ln0Igd7B3xCZmeFp0hyTpQE
5daHVwJe1IadVWITyp2edzIUF415wMvEX6VbFsKltRKiQlwaTvD+Vx0Ok8/NU3Nk
UDkBX8ejo6GWTYFr48YlztcjwMKVRW5stwk/cLMBWbnQXO+/65TFUjCq/moSOhP3
sl9OewStgYfsPeyoUDZD2LT+TM9kNPue8MTI/3GlBbqlgC1WxoS2VEcRKROsu5VK
Pdqfu+FgPBKK5vZxxk4fY84Bnx4zumR2tp1Q9xJuVl49sa8xaQljiJmezZSBgs0y
l8RDgre7qmjQQp+nu8Esc/Xw7kw/mdRYGZOgyTugfXxfJdDKgDkBpEWrf0LIkzUV
Mn4YKxJ0UBC8bj6hJbS8NaXmyUU9gg6R9fP3G7Ncq3QcfW0Vyq9qfpwb+EzUofRL
4qvR9jyJIE0vGTc2CRxTC94P1vkYZLzHQRAywLZCstXhwMsdsY0GQpRI1sPMtDlz
jfnUzzdnMUApo+D1ia2crJABtO+/B57gOLeK0WTLn5/je+9ybwgvFFxL+WlG9WDo
uTeUsP3QdTOkh1fv5BpfdzFZFbumqjuvzoYbClW/CzrCo2IwuGAc2+sugwZYZLY7
NZnC+WWCv+QO33H3IEya2Z47LgN/fCYYlQUrGJtjOPooSfEiLt8gjhcguXf7Bkx7
TsXiyYo5LuormIgPfstyhakWI01BFeJ0ljZNlM+04FQeNBrVLxU/fK7V8Gq0FXZ7
s+hjSREiAhVCySJse8N+PI3k0q4r/ZEwluGtkdxeIa7haz84VcfpnL19i1StSPuR
SPfkx2x8MwL9+KrguKz3Pkdyj8PwiFwt3HGRkhfDjdvRzV/iaA/4w+I2BnRt2qz0
fhN3ZrokbLRonOzbvzkEvwKhI3991IZ9NPw8EjxkBy3yrZyFQMYpYCXmosLDIRWd
20zLBt/lPjRGmYc7Elq/pzvUdcXDPNTonjSGHmQsc2cPpl4k/iqTKAO1ZvDnj5r4
r8vgHfVJM/gWfwgNnfCy8mIzLmBhc3XEodRLA516EJrA+rv49dPeSyo6ZaQ9dmzx
HJMiJGKx9acum/RBaKYgiFDGWDa5GYm9bkNzhBThZ5pG7s/XRRpMXldFM4V3FFEf
kYfHpoeJxkur37tUuSK7hfIq0AdrmJSZSGA2dMXTfqRINdenW3m5L2nOElj+D08A
QhiT+C/12eTFIQ7NiuJ7Up8ya0FRr6jfFbAwF2ULJdpChXF529NZ77f1yjAOe1sf
EZycrVtcddkee8BQhS4vx4D0GW6kopl0FAjx27rs/kiuiLPDw6MZolZMHhv9l9tq
yQSKBw87kK1k07BETfvqgJ0+5OizA3oBun5FEFuaF0HLeuuHuwv9vW6V0rtvxng/
sRtDr4sC5LfdYj2O63kN1Uvrh5n5lI1Gi9tlKBr6kSmoWcpbpnDIEhp39E3GqmyB
8Q+CvvaXuv7Rzmumr+cSpjaG0jJlpZQKIqGKRjWd50BDpy9p/vy1YnCEmAY+lje/
To9oRw8+fUdf88hhVSmuINIbYhhWsM0xmMqaszFMefXsEyzxTYIbPqnjxjbSouz+
0XLjbHeyJZBfPMA/ntBUc2vYo+cOtbbRBr40z0n6oyLIFeB/o/Q/VPfqsNQbvA2N
1wFRpG8Nk7CyukjT4MS7NlLPB0ZK8B+UYxFicoydWhz5xbkhBf8Q9GBv2s1zr1fY
COkl9vRyfJbVEuDhNGwWaz/N2qFZ5FxtYtZsdE91nfL+0wyeJ8h1x658AjO3G+XJ
80YeT5YJOgGDURePdgprMNAtN1y08ojI4IAaT6uZ1J9c7y7SP3fLamI0u8+0NoEO
iwkdRnDULZFodSe8ZRo9P349ABU15Ugszjm1HXUJe88BkvX2frxKm5A7MeY//PIV
YH/jxjdkYbMFj9A1ks7p9wCoVzTZXtfXhM7S6+9Ki6ghTNC39hlQYHIVmXn/SDtB
vmQuiMra8YXv/I5FyvgZBkU3H/xagZWUcSgP6ffyI6vobKAJreLUq4n6m/lWf1xf
7iGVMjvGE4/yLh/3dF5n9o+VAPmMzSg1oe0jukkPHqJll7sB9NMiROsMfZtCr5fn
8bqeAzKzcI5muy86r/YDfp8u+2PKrPknjLS8n+KDoQc07sk8VkFXes7gEtEKfyyN
ke1a52PYeM/sSdYa7FxCU76DgmgXcb2ZLfXztDvaceqvRmpcBD6c/sBSpfRSTfYA
Pg2see0o08eXpULXVZOVGVCeauKmNp6ACC9hJvNDY8oQLxGm7lzXmMPPiSrWDxkV
v/vrVVMU4Jcl8FlQyC82Mvo0ZWKxquuSBZYCewrfAb4Y5pv2koDrlMpZIqX++kjI
csC+8Nc54X8CldufQjWt3pTQzp9y90ZhpWNzBOdWzUT/VOenE2BQiM/la5rxpiR+
d+6AbK5I9NFlEvYwCItGmg+4Kl3UIYq4khDap12h92rxT2KZ2CBTWTfYryZ83rKv
OypLzpTeN+mCQGVfAL0VE7BVpbeJtjnn0cCZGaZqGr/+0ewCN9zzqKY1WPzU5W5e
3jAafWeb8oWqsPeQXjqqfeZax7YlCSb6zOyeqYeYuXtJMMYiHawWpaxZ590zrdZ4
eN5j84DSCqmut+drmCAdr8TOI58+QR5K7eqzIkPDyK4fOlGHiyB/CoBvgBubCLFp
JllDzs3gPum96PvA3/G53mkWd8Ta5qNlWwiTrEEP+jYKWeQBUDOgT483T+QkgdCv
BSZPYuy092DwNwF5UX8w04NVYci2sC4hL8lPZONSuFyB24VpaqI4cxaMM/BzESoq
Z4Bj+jhIS0nArV/JpKjVggkdz5B7NvuttO2r+flt81IdMeWYpFFFJ5ZRNSQJLxZ/
lsZj/Eqi8AKVAwTA3tP2aMFOQLnnfmoyQqmk0TqW2YGjmOSx+/DvS7h4hfdgqQ8G
+9QKIE6VmVqZw8xGAfHOR4pdTudiqJVlxjoHKPPMbjuUCaXmC+N7RRcXjjhrbyWq
4LYAFfjpCx90ixCiGoES4BaVTKOg+BhuDD+lFCIy0uYsLObS/9uZ02levocm7K4C
ymLuc2g9UQcXwjUaNo5Oc1aEEjSYn1qscOB3Dx4LZpAg1oEWRAnYRVbLpJZIcQNx
V8ulEtyW+isamHkQYO8PeI9gP395fxVH3KG3v2LDtMlSEUZEPMPLUV49G4IfrDIg
KNeUtJVaRZ1YflVzdmehy5qfB4EXPVtaEytI1DK88/18FOXrImHMILtxgRiN0hcO
kVSDHQVGxp7b3JFYug9iotzy+Mr+yFzm93SDBACI4toWz8rcO0VLpfxS7x/06lvA
HteuNlwV89+XUyVVVZivr04ftE8rcorakOJDUBUCqYr7WNxueEbeWaXAHi5TJvqa
wWcoedBi4uMF2IPdAmVBjSRH5YFViarx8g3lKqR6QceZVE+/IkW2lacUKDO+PGBI
RgVpezMFG7IYaB0A7OBaPuJyCiF+8mlc/7+j5Xdvkf9Q7raIStWpe4v5mzwq6xzp
1r4XvNstGUkyq2tp9JCf2Zf9pUCkfZ93Ahpi2qFiI56PkM48oVS6mWLyXsBgr/mA
W4uJ4alyiiE2Xlomd7ACsBajhnFP4Pr8NT/Yc6tjbSHdBOBPsb6qqSZ9piK1+Hdb
e8mCW99TMibxb/xbiANBKENZ/XuXpqbxL5FkvRaLaMzB/oQjAg1dTMwhw8uBXaBt
mGzMegJELdmXsep0e5dsQG719kYTqPTbII3eOg+LuLC1G8gNMqyN1gLDWz2w1rmg
uVY59ZCbGK+1DYCkNr33UVJC6bNXk8C7HM12kVM+jjsC96nJabot1ryEJ8nrwWrP
m3oh+sNFUMYXawyQX4XPs3y5fW8e8lj4Mxkxlt4hm+kOpJAp2l66+8dIC7mEsVmr
y7LqR1t8/B8N33DVamUDET+K1eHMN3q7EcnjaSNmL7D4IMianF7xkyQF7lYOVM8w
ktbsCFIRoFu287zQZKcg0lSQiLLrcJRmHJ/SEzuKRgkG54DDB2dzvopT4UXwIy9b
rSwe85W7hDXVsvTXi98KfKyz3gabdxVb1o4/e+0jRWkHMHh7AI6vsIwjc0oQj/LQ
yRrn0YnjTsd6Tegdv8Z9EU0eret1obc8Nmj2oKftUYFtF4vA7MpubjZFiKxGEAYH
5YAxzndtFEMhQ3FAEcGaM6XAjchScQe16SBDLqHJdWl0jQGdp/6O33YIH/+uxqUj
HayUVPj7ZyP1uTeYd66VIkavbQI8luCHGZQt43erbUbld/nqky1aFuZt5D5OEas9
ORpSsjH2jXI1TUe5+d+h4UkwMGT+AUjfCF7r8UCBYe99mXjO3iv/yzuM7TfZtvO1
Vd3e+N25d6dqI4bIcT0A2vzSjoGYD7Npg/q+1cVxbGpH8/Rs5B7sq8l3FotTwg8r
hZc2ZTDSwNmNT2A8jlPzGGegh3FlZY483JytypfYgF22Ev5dk56xu1x3wy/qGfhC
Whe70nHtmp4llUYjqQ6PznVouRdd85Hhkw9taFYUhZL4KmRVtu/AH4WTI46DHL5S
JuNvYVRktcE4XE2uE+x3Q836IwJpXLt/uITwZRntVqTs6/N9Ia5/gX+JdRuEYJY5
znf5/7Kuz3TuQgwheny5LqFNWUnRVmke20+p6F89N3GHHdnTNGF8wFdfacnlTxi0
mOT1qf0AraNiFVwdNbuEIKbLnK6JIgHHcNoawF42TXuM0Qyt45rtlXXlREvtZKZh
FoOFpGQFFFjLncVWgXJL/xxhbqis7Le5PwdvyXgubo7zgmsIPY4NW2hUdLffsHid
UV6B9KqmjY6guE7Wiy6Th/lYXh2R6mETgXCOcpKMHjfayqEnkCdwE2JXtvVCyEwc
gjBLozUiUwHQbsVj0xsZw33d4sccKQ3kweGihy8CwCcWC3rKsAHOKHqfTrqz1JOd
LYO40kqdEC0YPDDcEQ61yzMMN/GeeK6k3Ec9jvARTvJn37S2zY7w0qsEWbHVtpO9
wavYzJmzXmrLm6wac2NGB6Z4Qawc9HZSAGm2yg8AHCMJK6o6j8z7i4QkVpsbfoVV
NGM+exZmjNrUTSlxFVh0Eg86540MC6FB4lM9UXNelBXUG8WoOqRL5SYpXqwc0Wv7
hdImyNHVITTbivPvq0q/Mh9WaX3FsPSiJU/2+FZ2Rdud7iN/O1EmT0YZIO3Z9m4c
8KdEdmCfHbOoLW62lJ/H6LrFNUQyVknYIB3cgATStuqSR1lSg4LVQRHbe3zorGDp
vBOBuxJixJHumyDbJTM5sazODOlqkzNGKYc1gTtVHY3qjzoJYd4q++yn+pFCDPN9
9IkuGpdMBRruTeff1Ma9ZTwK9YuIEsBA1Pk4Rugo1X5W3D1DneOLjw2x/cmqemOt
TzFHqao+E5t3rKaKtYkpNMBBCIU2KM4PcyL1tt+2Yke0A/UNm6jKkoYpm+dMfkL1
CzqZgCWYO69CeJhSPAy6W0FOPansN0Yk+J+eI6ZsGyQ6vwwklwbrEDkTVttXVSQk
H+nnoo5xp4mZuAum05hiK5zhyir+NAZ0BeYBk7DY41QHQWp9ailxilf6slLRlgP7
DjoiZQ1uJ+18GXeNpcu22HHTmxCsdIk1rnUIJuDNPqGAJt4i7S06LtOnasq4/T7y
zQniHcScuEQDvSA1A+EMdjoKL93XqwDurA39gc6MBW+ICIurdIsKOqC9NCflQNOq
W4uZ/xoFrTXpqQNmi777elTgsqVwhrvZBFwIgohxD5pYfVS58BpjUOV8mDBX7gXw
KjnUw1lrPfbu5//bqVMX750vLeO+YE7U0uRssF8JOOXi14mEneHg2/c+eu967lBv
gxkIWMIPnAgBslbnQmaD3Bcv5tAfpmcwrakzYaQxl3w+Tbz7HJvyBuuJ6+2vmYit
ojoFjsgndJfTv0AD0oLaaNPhVacHyrJAGCdAWPEaIMsHd5Mpr0OaQ859QdAMG2hg
yD6O7J55+eIgS85LlGG+3sfWT1WwcltI75Ptn4VieKPkmfFd/shFlizFfgpzd4Hg
ol9eEIquirlABAc7arSv2fbyE73MqSmxheHNUctXy64wZ6edu4zVBdkCefCzDb57
Vt1w1EjYzM9hc7nVn9kjYgg9KJXXnL//IQ0XCaG/W5DmETydouJMAjEBORasYllL
ZplLCGADedgRLFnXkusaNX3AyPstY989dTIE972Om/Ab9slvcVCB49XS8EHgsg//
dPpGspECKuDr3z1ypj0wGeFc4XJdxuhpm5xq1SHiwgTN/fgXILbetYvNC9kaQkOh
6FqFgicynB2hrFLOpB63mtSkjpaBG1S1qFZOaEF/raFvNGwMkdDw8al2tWngJFmx
FqKU5RH10yP4eN19YNrfbpmdaAE0ap71Gm589iDaQO1uptLqTnYn7elpt9uov5/V
Ts5b/20035NhUuQiIhBNJsuMx/6LAh2nFx4KDCTfgfS5USom++8A1bk1mqedkZgP
RtfuEsBRD5ATBaCcYO60VNJ4ZhOPDP3A5FF7mkCTSyjHWTkA4FMwP1LT1qms/8+D
EOjEg4Du5kfoiVFabNMWr/nUifpLghO76O3T9PLiYyoX+ZpT6XgURwGwO1Uh3U37
PxDjmE6oG86LJ+RKGTKuqzIMsPyJ4xRwfos6EfDYAF29sJjG9SWfj1bgVtm4A04m
o6Q9ms5jzUWaHSUBqu8bK/ba/RFsNPxkMfokqf2BIaMbPVVldxGSXPBoDgpok6Ag
WfSHmEwduBoVAnvaAsDNZcQ7c66O9DmS7IXrA2u6vX7TflLxej8JGl5gNwOEX/X0
8AhkqgQt4i5AEYsTxK/2OXs1vCdu8/Ab8SKEdpJ291hnsLhBNzyOvAdoai0h1Ejq
+jLrCG6sLJIwcwI34MaLGI+m/fK3R9IZsiNiiUb5to4zR5ORwlqft5UhNqZHAcgM
U9JoQy9W6fgXNjTqAH5Gi1QidajLQEuA0eTLNMveYq9gHkpLgLV/SvjlFJLupWFM
u5cvmMa5iNg+7uaWCSt/bfj5awtKdhS367rG05gZNg4Wuc3YhJucI/5dhJxEkzPl
XvfWo/Dih3roRoUSnWrKnGvgCNoFTkXHjaVQIohMgXUYEP/dx2+gmDeCjttTZBm1
dZBiI95NUNWGIf3OIuKpdqQqGyUoNC+gwooKCSMBUCw9AQ3/gAHNpvnC4ADrBFnS
cX73Fp9EOl9saKegqp3SeM/ERRwBEmK3zJNwFL3ssTcpkk/44qhc9Ba8gSWX0l45
oVxEVb5F6f3T2vaW3U96S+n1a+u8VcmhUOKvKECCy1Rq3QwG735c649zQdOCsVOa
6DQm9nNL7oSq1TwGy/5PNgIsY9PS9UnOltzu1c7nEt6KnCVGPzNbXPbYsOHwXjs3
qchEmV22P5LRFcCMvTozCqdsVKKAK+o98eJuuVSskeABaLCkYoCBycxnzQhA56pJ
vSLyjRpPljgSiPez7atrpI4sdpoX6Muf+jdm0s/6kPcyXfMLeb9+8ztcGL9mGBqs
k322WIPiBHz85MQT6rQ1fznLl3efuR0O4d4yaqJYm4oNTP6wbScaoC6bcj424+Ko
vC9oPj0LuYG8W9CVhU56luKYNzDJHPIlCsoWq2DlirO8c1dS/QtHJAcNTQCmkXCn
jcx2GRZbE0uWgirxqoICOOSAN6mOjQ9eLNA9d45yw0Pn9F9rUDn+4ikbUqnHB5mU
QJjjfvvkEmDjY1M4Ea2tUNij6LyZP8B+Gf+NneCIcNrwb36U51+fwSmFOmvw9Crh
wrR/SjirRDo0RAXoHfBTN1JzeOjg3YpKItIl7cuo53uE61b4QP2Q4zPkw/Gh1e3z
cf+cflxOJV5wuuV6MMHbZkp7xm40+Qba8CBvkR55As3OSyuVAR94eRKZYoAQ0tdt
JDCCFJixPCsK32JZnVSKWUF00tB4FslwvzjynOcdnpak/mTSK5+tNzIiE1wzAt4a
OCHwMconlJKPDNo9N0/QYflXOtv4kL5crg7AC0VDfR/ICVUAFG06UpHr1JRqvvFf
gy58Qr8JjC+WPwXBHfgGSAsKipMOuAFc/MaYEe2LjIqkk11shYyx3Fq3G/mLuCWi
PquVJsvrN/ttvDMJuwFvyTEC1cvF7qZeG+MFEacPMyxavl24uVip/DNiOR6SdwXu
DBznjBiHwwXkpaQ8KyvecZN1t/IuyOr6DxeRqO8NU90c0+aaDtdIKVx8BuMbuEoR
Hq5aaKvUkwnadHlyQp80yHt+j01wYQgxyI6rnqgHw2pBuaFqB2IHuq7TTt9+N7DN
DwQKm1EPrVOHAuwbGXhACYojUgnerN0ttTXJNRbccyMQUdQSVAuhq+9f7+50ShTI
gVf3zKSWCH+aKa1PrlTA1yCIl5xxkDcRpuxsV78J2IHPpzQvvmqTeqK/0+znR6o+
BBrmrALYIByX+1VUsUwRGd3uuNnyA4sPcPhjc4cgQJTwZO0Fk8Ifse+HMEfO9A0N
kcX9y4Hm74TV2zAPQ7my2Pxwk3G1GUYqyG2T0KwasVeBBYauBAJglkTRrwylYbJ6
XR8NByeZZ6sR8yQKKA+SXgooAj1NCDWXstzTWLxa3e6YH4Mh05DOPctG2c7qfxfV
7c4BGd9wUdoNetNUypc267u88nX+J0wJIXMG1hxuZVgCAI8MDDbWJGmKeCuDUKJq
QpRmi2MjyHG7FyR4joWXn70Xz4JwKA8Qcv13v211OWDC2Eexz07Wk/EfrPxHjpZu
foiT7jAi43IJ47VmtT0Fs7JXOP3o4Lct4211wPVyxXhCYMN8sy20JfkzdfTVv4uF
OoJtPJd4QO+FxTqnVsb9lNLpFWkFuzNGKrOTCYl3o6UY+D1DW3rf9FmL5zjRsdHX
8XajwgFrmUzrLDa9QNF/zek/A7Q/e6+PWccGtxlAI2cIotUhhwfGup5EuDoTie3A
yB9CCUZNsUon/XrfJ7e+7QNeTxfAVebs/ZTAvxDggPMcWWC/FbxzJyYgH4MWldzh
JqMoWIJhPd9iDeMqPi0Jdj8H/wbzHdZ9X7QQaAYG32v/LcW4P+OP8B4ETak5lfxK
ugPJ+RFu7med3MkuVr7MH+Ovi/ilB/RoZmHoy4axzjxr3mp76DcffVllH4M2Llmr
JnLlat3hweSQKYDiWnjS8nlh7EtyH6a6XSwc5Co3gE61RrU4lUUKMmgcvUmNX07w
aBPxNguF6blTr4zI5Hdn1GmiEi1neaQ614Gn1KNxKOO5RncAQF+4lS0XhVSCqGRj
xvHTSl8Yc9yFjAMFnUJNTFFljsYutxF7ESdAdnRoy/Fm4RFpyYVoYwV4P+lXWBOR
/9qg7obTc/wCLDigQf47fstzCRGU+4NzVoobSAor2RMeXE90imY3hQRxv3gCJojl
SD3HJOagbVolQKodLsFFQ5Wsvu28bz2f83gf1BxQMnUeKTSZIqOAKmpxmwPUxw7e
5dMPv+2Py2Gw0jzASH9n97UQGR5ts7/6R31DMazkAm3HZoO/JYaaoJd4d67Djv4S
b8qP1/qmHGiexaxv60KbUBRmsWuFO1TusJngOcILalIDJAnP+OIqrcDX6vd3fqp9
WFVcWWYoDWCtYQtQgsa85oaf6pMOPE6RZ+oRrsn3EWB2orvNMFBBxIlZHLwL4vy3
AOU6ypCjYBsl3Mkr5XHhAKFATqsSUoYmgEPiEJXEvPosgC3zLLncsuIGKLzHjjZJ
VcWjf82wdNrfj7iFStfk/ArzDt7cCu11PgY7QDkWUp6xJLCegT0UZawPRdXmKggn
26ebyRgcnKNm8583c7ZY95h3R/c9OlpwQNkH6E5+Mqh0FVBO/6u6l7hG7ZAZeLNN
ePekKzv/6p4oVnBilEWsyVJ+iS13FBScEJvojNOkFfR1RV8+OBZyQquB892sZvVY
CDD5BsUAwGFQ1eratQqlKaIEcginULXP/lix7GiyOiTQzyolePuV1ZlWLjGB0c9u
qqsLg6hqk+8ajw7WvxM9RZxpNdVPxnOVD9qReQ1hYv/O9t7REAhHuw4tXhHxZnp9
n1UdTieg6H9DgOXVVgoqmLWj5Pe3nXV/Lfi9ykBFGWRcEEaIPLJ2koOVeMYarW7j
Rc1uBK21rF5xLhpV7CUVymxebUvtsIMvUdrWHVQdRUb0QZps6rhLBp/skR71vdJ3
ot5xrinvvbjT744Ze1z/W0NoN6bzG5OlWu8W2YLLrzuvVrpBrXFA6K06dePcnwJx
DA4kxhZTCcB9XbcGqiNAtzxHgySr9BmuimOESrZ0sS6VPO+R9+MMQLvNber6BN7X
G+LeG7MW2iBdpGOJTP8bBXCueXRByCBCO4zbaDEnLpxXWYwZEV4XAHhG7rBx57wi
ZnAJYGoyU3+Y8tu19eaRIIYGIhuluF11C4rTKyyxsRk57nPy+HbU9+UMJpgOLy8r
3CSV0cMBJyNeBEZ4oIZyeGEOnZb1xW3XhxIt5uh7zoPLFcmy+yMqHa2mLl4edDIq
WI0iIdozhUni83nnHW9ceywxdLIZXXspzdMJtVr/ereyBRC7h8fJJl1BF2QC3dz9
SHXfzVL8A4aXzj0CM28AXVY3x4DE6Mxx6A1ijCGU2R2qy2HBHLLdiYoxs7QHDgUw
TEF4FNWtWR2docGIWgbUOqjElHOvZeHhHC8ClqHc9/jPaOiQTzxTNwaH9+3lp0SN
+aqEApalOnEFjAMzK1lEJHbSXNDAke5/kzbOFJvc3DHvfBd9aOWBaG75lx819rkP
J/Lok7MofQDdFMCUIeUVYPbd0GsroO/N1qpNFmQEIjlcHP+oGtgfbyhiFpozJyhU
Jokbpbjiif/wvoVEiyTQXsTDyklwL/Ma7Wshyce6T3P9M+deu/gDUT1HhhWSJoCO
NyWGPdWi1IZUpgDmSoWdZFd/yCHDtkL7/pUZOYTZtWZwJNaLhvpcK+DNuZKmR2UX
TrLfHJyya3vGmFTkrHrkLkBq+3gJlLAHmSTCLXj4mqFJG1eiN7knK4NbVrfwC8mu
ocmHfHpALifYmyYpaC3YkdIoSB24oyhMJpMpDh8aSzrnIWaBAbpjn54s/Mq/xyEY
uEPwXDrHEdJWMGMYLOKhPYtlJ71Iq7Oh1K2rx/kcmboDm5GxvIpMSkFzufqbt2ny
jf/tE2y1JqtTOY3Lmq6Ns98lblz8ENai41RqW0KoJs7Va7+5knZB2TBKkWeAueFM
ozlRCunqQ/7xhUmrWvy8+KqeHv41s/D2K3Do7M++ogueFzbVKm5LwnVppwhgkBBR
s5vodKoGucBTqcELfoiJLZVn/7e+ipSHXX5ZJeZ1RwZE2EE/nr2oe/WrfhsAC884
3kndJ5vl6XXgyXf3rNWr6N68XCf6iNjyLDjG0I68Uf/EOmeI/A29RyWR7yPF/jeX
wdAI3/enR8hhyJ2EdGqLUQLXcL01RV4LlRy1G+4V4DHNWNtjx1jn80M2ZSOW+NYg
SLcoX78vCHJan+R+49B5J5RxZZpmvwc+VAwrJx6VASIuuDOCEcq81rAFRpFVBhdu
VOw6UZOWeHiMAJ3sF2xsscR0El6118Z7MLCNxxMv6PO4JwSmFMseGXzlGM4B9lpD
crCsu+eyQ604ppfuP4BXiskxN+f22KOeowZblri5lzLX0vJyVnLKqPs3Oq6qo43M
wihOAbkyCnOk2OKwJPh9C4p8eP6mGHGb0HEzEE4Ytt+jON50gIXAs2hpYnC08Vp3
0CnrZa6fx8wRdEIyoGOpjucey7pDLXau8iUZmYfPzVFhNIgy653hTH2JEIWTAXTa
WEqLP52mXe8IeBNA6ons4btHL6PmxrzOQSIHv9VPm07c49GkOkt5Md4du3a0vNPC
03OVtC2WJGdhtfkxw6rSmZpknZt9IkzBhBJdobGrh1l5JprC2DgBIDXB/FMZ3nlD
We3j9r/I1H3BvIde6os0LTDiYB2h2C4ZZi8tZYxlFn1ZaFrXDvq1PieS0AnxysGm
yezRMmr2mhmT6Gimd+sebESfw3HfBZjYRXHdYDDnXSOMqm1Iva+lOyzY/FX8q0mW
eI6kG+uCJ4Cur4N0Y9ZuGcuyfSi2UKR7qT00PV7JLyet5Z0toGvm2/wAN0Ol1Ld4
P14oxxxieun+kmG+S8KmCjo/0lk431glUdrAi1mSF2M3ShSmcUhcP8hxxBHK+NBW
27sOl4PVIMzNX2zaWwLc2wJ0OvwksL/rYmpC/ao7Y+2bUXJWagXJ/3ZR2CqjZZgO
Lj0VN83sKifFwsmG1g33Lh5t+XviGrmayuf0Gjr7kQXXchBO9tO7ZtJa40GGlCEL
9xEU1qp9juu0kADMVQr7lCbGO96b52prJiV0X1q83tArjeHGkcog8UADgHPqy2i5
PBfM0rJjHuT8aAiqqdMD8HfSHs/SFRpnuWwxXY7djewU4omNaXZCtGCWiEtB2coP
ch1emmjx0VK52cv59n8w/qsXkUig0x84JE/lSoYi0L1/YUC2t5JJns82SwpbQMrH
cOfDCpcsrmeyrJShBdlz42DSzRuwbrUMO13Hu8UsUMISuQB791nxySwJldDBPzk5
SwZl0MRxVki3p4KZQDykzT+r4yHLp7SDApRd8Z+qDDcGm4LLHWn8kkK6Zs5jQ9jU
kyanqbIshOB1Qdd86TnQ+3ukhLqs0/HxDfwybBkRJMxCO9vfSGhMMf/jYPVcKwcm
XNSX5S1f7QJ5f3LXTpkqJZP9XuRpwSx9/vWUVq/vuNqaUS1BHBgT3ZRuva8qgh2v
IdndRgtDuE20gAzaOgbivXTbOT31EQnB2Ik0JGTufNWS5VxSdhIg7iX0Ya1jQMEY
U35V1r44951e2TW6BS2dYISHE1e7nEOVoalwQfOT84m1enPskU3FpxGpghIXBYap
uI/mLx3VXKJ9AyEN21jEV7m7MZx/8Ti+VQ3EsL8CeiEUuh+gkEq7y8D5Mit6gX3r
Pn8jGADbG1594eeREu2eGKS9eRq5f1Mfqd8JuaLcsAzKaCz4SnLZeaFPXE8RZDmK
6mZiHgGlphEKJQ+PBuQcmNfShv5DzqB3coseU1UFv6M9KMEIeZ5hJ1KeEO7wtNIT
s1cWU5+9NGEETdvZYcDz6vpBpFn+ubs5EmBF/Z0NEsVCeKL+kxjhK4TeSRyj8ilE
aJSp/Bu2pxET7Ta7KwleO35XbL9O5eb18L1e5oAVYY5UbI8ZhmdEcmT3BGfd7ETE
Nx4fUkLeWzHr2SBaAc89YgaltT/hzEDaGG0AMiPMyjiaChjnH0pBHDI5ixbCFVm5
Yjve4376KUOX+cuVPIfcz2Mad2EwNoYU2b24u24L7UvwDYFY6AxaBJqWDQvcQna/
paWjGBJ24IfCR3U7shuN/fugbOY74tEHVGCl5vKZHxUdNMESKsLq6pyv0/QowlRX
qZKtBe9bemVz8p0ZPpvEBmY46zDH24pK51zP4jGcTmMHUBpjXbxKN+HH8HuFalTe
oabQX03jWFEtLW4sNdY3IZ0VrJJDvllCefc8TyL3PyJ7tRrxJUiYskNrBBrL3m25
6kXbcjNU6i7RnhbvmMS/vl4/Lzz3wlDc0NZYhs8eUpu5Fc1UWEkMjg9RezDSN+ri
KAbEaT6AaLZHw5GYljcdSnN7+Qdp6ob756LWMmRNwBh3+kHM5ykJ3XvaEAwG9Oi/
YICwAIgjHvCpBhLa7oNkqDSJyt6X0QF23Xa4XCq9SAQ0GQ46ttWghmmNUxzt2buj
QPoE09gLcRoSSw/Ih3+oPTF+msHSJLgsURB/lfur1yWyi1o4teNoHbIUOpSFClVJ
VpbtdldRqzusxKt06296Cl8AAA6iafAgAwpc49NyDLqv5VagwQ/ithSQtNjBTo0L
cTr9i/LvcRdH2mNrXwZl1/lwsqtc4Dw9FmD36w2qv8AwSLzenq9dD2p+9uirk96w
Z5kG7NU1OHsIHcBB+BfeaYh8lSOx1MqjQc9JPPgLBiOo41OhnLDjOxwaJ1+f7vdh
aRlzABI6BVdv9TB3IU2+oM1dQsw0uagthlo34PAvMf0f7Ur6WJ1GeruJa5DoPGhd
Xbz0gCE5mBUtNetmS2S43yfAW7ZPc7tKtvsHEvDxB2o6dvXHDjFv8P3Fju3oeKNu
614CWp1W6fDvKXshDhAXjXu4OrJssGmFrQav4jkZ0JSPox7LANIe35LNdfVqPhYg
y5MnoIUqN9dm9aBXiLMr0KsqViTrUilVehNiWwzL9LPza5MrgCq9NG53IMqoQNny
xdO/0MLFCBr+7K45+RfBuGLTxSKCI4WLsK7dNUq9omMbyQbXZ1rTpMEv7/HngEvq
HQQO0L5JPri+kLKYiTlOtYg54EjLhfVi0w+0tHPrWxv1ZL5t63s49Ttk15RdHR7F
vAhv75KaXy/GpdsA5Nkr7Y632S0YwfztaOFLr4CZ6DhX49ZzE8yGdHm7bLFjyMm+
i3BCYmC/V6lX6xhxsOTKkxKBuRednQa+MQqnMwUJg+F8aWCASVQK7tIiJkc3pH8G
mccfIrrZy3RlOd8Wkh39CE5J7YFWKZyhn0UE4nnSGucsAMkuXH9Zv9fy95K+4oU8
RwobFT9uNPQA/xAr43Ph+lIKDgxTgR2DJ/PoKn52t4lJoiNlnxrd7pcOhDNR3Hcm
vPgLbdOnOuINrlbUntdBZF+zYAuXO457OSV/ADtyHo3Gy1aU3dSeDsmXu9JxTLHr
ov8fDvScgUj1KSCt/ik4tsf4/EUFTsAKdUMUVesrqC5CqT5gKYEE5cSg0iy7+4Y0
B30W1OKrjF4pLFzdVUb68GZfO27wC7gc9OiOskZoRDY/gqBbvK3kpznSgg9xhaPo
uWisPhQTB+vfSkqrt2OYPXDPIKEVyztzfXgdQoREJk9ipQ9ntKNICwzncf39LlL6
yKD8bjjr+QJa6jZx73m9FM31sGJb/eOkqn/MlnPDAKyvjjLhjbiwRipPOKqMzhLe
mBXv1vuIfQiqjRXz97O351+UzwQmaUSNzy/T+O5LA9T23uKUGsIkbRM3huv/LpHC
aeso0hQdYjn7cQjqq42pm6i12jbQG6s8DLBzMbn8F+x0/emZSUr5zfNizZfjOuQf
MtGVlnCr20ijxn7OTjFeZfBaAD7jXmDLukAdTLpMRX9QECaKhm23GU70s4KsWsrz
KsALWNCIVJP6BXbMwowIkv32O4FtqRZdORzhZjvsjb7UY1u2x6DGvsTUQcI5BxGp
yH8PiUngN0qVP8SebV5tHgvkQxicQj4a8+Gj7oSa4Waj10kRl04IY/guCUE9CMaQ
5oGRVlE62my1fqNR02H4nSMHaGX8w4V12ylnaw/2EzMzeN383aj+Fngz9GlfshyA
OJk3+d+cuvmrxgT5rEAATMH/hNCiby3V0R+pfAc00S0snl1B4Eb6IkPGMWZZVogX
W7zVqNihtxGMCVwonlhesOMpE47hHy7U81qcz23zVZTogj05Lc8jHOpHG0esEinH
//i7H6re+iM0mgssZfdC6L5F6+suoRx2lqaF4gzVwtTt31JxYWmELo8St5hHfsDI
zfa1XcW8K0skhdxdlE4VS0Ui9OxQKGFv2uFA2RiQSUEg/+I+VCU1XbeoPrKbP2NW
ZB9I/53FFJXiJUiDa5HZgtmENTFzuHYLdZqM6HHFFWLHwO2j6/AWdi8LZpUgR8SR
MidURb6bur/V9i3F814gLXTwuQK7JMV5vcY34mRq8MJJx2Gpvmc6xw+ejkKZajbW
Cb04bef6qCw9VXHQ/umToduQwLZ46aywTShZKihioerY24Me3mWS2ziJwet/fAHl
rT0VEgHMCPROtAzsH9fnsXdOoUUZnfhp8p4OEmcazK1Le+FEPK2t2Fcba2Bfq0PI
pyuviCderQHKv7fPBAM/qWJzfGNnmqrZ3EenjS8sg5r96LQrLWbhhN8Ca7ypkZ9M
u3kCdoHLB93ACeFLEwrD2khKPuDeKxuTjJysUxHWIH7wbZ52FJZAeJjpVtmOQ7Y4
n0ZNJSQEe+E87VQGY7nB+dmFxxaJke+rHr5VeWipH0s7CnrJe5JeHnPv06W8K8kO
V9itpIrIb6HzTEWuQw0ucmqW+8u0mUKv7RNQOwJ/iFzAJsEHZyIxc1zgmxbXqQ7t
kuM2yAavdS2JhEQIypmmisxYTiwj8qhrplhjLlAqqu7Z4HtElgxgcT0GhngLy+Jr
J/xLLqdBmBkT2+CvXglwcDBvZQiQ5Hm92tdh54YX/sVWtmAfllIEk+4y1Px3Ovzd
RRU2Qpb9T5enD0tjbtBqZdZQod1oC+ZGItCDuXpZkcoF9rp7wRhq7kaoQxqHdsul
n4XOMbb7pTv5X/pjxtsu39bFeO7Jsn2pzic8HUeM9C/bUtdrVYyf/tK5JCsQzvpq
V2ayCUrGv9Zza4nLpSkk8gQkD+Oeyd0n6hSU8xwtWacqHX9yWRTgp/Wz70tWluHN
9BylYQKeqDbmlCpNfQoE0+fiAHJimnxU+F20RSjyjX+IzchCty5aae/vWqESfnaD
hnGJ+SPU17D9UASFeJgquhH0AxYO1i20bR82hMbsUhYTc38Xp0wTXOrOMa1j4f9G
aIgI6JxIXeRqUEEci/LcGLXZXrP65GmETgoSJwreqVyYW6XM4jvbjW7M0czc/PQ3
eLcejFaG5AGtgzdvcSeE9SHykaj2KNRJSaum6w2ZcXi37rHr8nXXlVlfu3AHnqzZ
jj/C8nrQCLzW7CprZlpiM6jOiCkMPGiwfXpHJ908MWdbmZELtfTUVewyRZLUQD65
x17mMEaKlpj3pgajEFt4yBI8UKYJwwaP/1320yS2T8t2WnIuBbfyU4pcwGs4YW+Y
nS7/L6lul3c/ly6BJ+nehDD6/gaSZMD9h4boE8J0d1HMl0999M0GZTg/OKf7lFCv
cqD1NNUxXJqotxlw0plqweBUTJ7lKiQCehahUp3S9EmHk4oLdx94ab95a0idXNsj
PzeDqKVEYg538fJoC2fUMBDnrSMV33xs1Z8csst/UDXAFDfTTc9Xgv3LLeE7DJgV
kxoYuT2FALCrgKGNOHgX2bH4U2T+rLHysL8R+16sJQB6B1Ufy1V0Ln8gZB2OUqf8
SUj+Oz0w+6b6lSHxG+qPlIqynsk6cU+uv8Xaa2bgXJWkViCDK97v+9Y4lKQPr16o
5Ku1fzkoo5u1o1PJJfx/cMoIhWg9f3jVDTuDXYGGwQZk9LC7iK9oM8VFWTdwwNIQ
CNOo9ELLB3LKl+RR3VchCDZQA8RHIxWgSjSsKH7YFi6Ff01FLdudEmiA56J1yYsv
T6rKq2C7CmnbnuTtGMOdCmdDx/9Y7BOtX2hvnwmnlRtEKjqQ4+jfzLxmgv6V7COe
txnQ0j1TuZ6/jq/Yzmd+0VZarEvHjCUcvm4xeorlvQwkB0sbQ35Gjx6kWOmHiNae
8vk71xlEHXNWbbZlYN8qq7JuF72yCWmEGnTHPlYiaRv9W2py3U4YBeTzmH7N8h41
uLhhZAQIeX1bxN2uSwu29j46l5d9H3dLQafNVyDjigBTxSStGV9WnNg78FMyHk7R
doKyhFTeAGgKCcp7KGOIyijZvMK8gBT4P3IxmEgPb6k0hnRdCs3o/INLz7096Wd+
XC49Vc863fGEtsKEJpr+FeTwSqTiGa6RUsXrZSV0Q5wsLYbtuXRTI0KsgL1UbnT7
lpYOR6sYGWHKCsWmR7Q3wpE0q2VNC4alfzy3RDIm8CZkmXeXNi7uZeLhVM0B+9f1
ZF4Go+2kTOFgWQlFu0S7muuxoVBRSmh6BV5hd8nm7gjY6DvGNqeODpsFbIF9N1gp
wXElkn+PEjzbPFv6Vg7/vjtQV6pKSpPwINPuwAdn9lwasgXjxCjC9J87n9WTtskP
gMda2yEK4wOQAkQtGJHvzv4rd37x16wlh0B2Mgr9C7xnOC8sHb2Q7fxLqFYs3jP8
8F33mmtM+PPCFC5fun7TobOg5Txu5EmatPD/hEeYA3LRLlzZyrEODm+BLgMB/jw4
P5UtiAZcZnXDpSw5ExlvqWK/ISyhb42fo85x8kK2vFVxaG97Qt72kxiVEnX5kYi7
KIskkuGoZqIG3cfLgM12vfkSA8WQZuzIdNzE+PZHFgHQUAcqDfSUtwXL4mFB9fuo
A+T+89qnPNONJTVJTBGVdEpC2qQ10CABk9qIGTqzh8dKbz0wr3HQSDwkvgcTd+tf
iskO4vYWwJIrIEX3b7e24/t6ynB4CaGzDjcjwE6HaOI/9ZMyNS8fkxGL3IEYF3A7
8YG66/WyySK2Y1KdmeWxsg4cThU94qfo+rv7A9rYzh4v8TVRFoR46H6vpO9P7JdM
qWuM0dh+ZMCknAB2eF9RJ4Ko9gXNoVMk/RMyu6IRARFiCo05ABHWF7/0+UOYW2jQ
Jjh5cWwpgPZOIjMH5XB/81xL0vU7RLVeA7ARTjiS8ws3EXXnRAGCbV8INqcUrpuh
a7AnHDC7OeElP+wOTuATob0T62OBVgF6b24fkJiool1kGq+Jl8zmqbdCi/OGrFyF
5RlkqeTwBcKSm9ypMCkxP722ZkDTaMyI1z3lszjzLt2as/B2mn0QmGxj2yoULvi/
AFIcC4p8s+4NIL+AjW1VsMjizIEZefm537L9NOMAGUiAN4PqR383l3VYAvPx6Wsx
1gd9RC5FMVO6vuGRH2wVjUNcrAVTo78ykrKcEYaiFx9DM2e6Mcl9aLGDjAgCS2/K
FohG9f5p+N9FHKfmbAAEFEFFXmYtZth0gC1QA5ZT6WqB0K1OPh2QmdkjfrybVKTX
dZvJhB/o7IisMzRN9zMTaXVDi9Xwi9TrkFlLu+VPbQnT8V7mATAAP3Rza9BhRWSA
3n3RFrAFyr9y8xy+Coip5ptrHJEzu1Dx9J/eLhr9Amn8/sX/pMIehFiScMiGxsh6
peUskXWRGua5va/8hKSIjZajZVZ2FUwm8GJfBBzKe4Vrc5BUdi4H0KbYzd9IH7LA
Yk1f0KekctWWJEyd850ucXg0WgN2DAi51VR1hI1t0mP1A6B1PQjSuqnLCM8mYZeu
d6oEz+elDwN31Q2dmxV0ovpJNgG3yJUS9488IvxB8pZBoaBPgCXK8wxmEpmbk1VA
bizO+zk1Cs4fdc9y7hwSzSF8yFBTU+e1WnXc389CMpYVfrO0mbGnVv3BoCcSb9VT
EVB9oH7eyyH4tUIdVSwEXbWcYaUuobx6XEO9g9ghQ3SKCfJ1iRIrCfSE4V87zCKP
uF9rf2QfsQzmA71aQIWJiGNtjJHL0JTl9WrQBj4FXd5v5lcU6Frosjc30VG6ulOU
x1oQFzVdP8olz4o4yM0gUovheueK/gk2mxOr93c77FWnnaP9kKSw5gRFvMoUGJaG
sh3lL48Et6UUtXlwAqu6MoU0EwP4Bt2OX/Qcst0Kp39Y5OGdlHd6eyUvmV1r91qy
9ZfGW6Vb8Io09Il9ARYdOJV/RjS8Q529Pw3HN/aG+8fVmg/WqhLzpBHffaTAPkmQ
aKgf4bpMCJVAryKSEJMEO4sWxgEm8jRZj+Ns8//1NNVedpdy0ytzH3zFrsfpEXks
nam8uuIEkpC/f/ZJGPjPXCiTCVBSfDAhTbYURYo3qlQPr3jQ+yfZ/CqLpoEF3/u2
pqXZ/QDWBRmOclzrjUBHhP+fwCyQQQMReCfps4eXMttaOpHOmjueGiU+kullvsOE
eXiymyXVTvXB94QP5awO9m6kbe9k+2PnqZVxgHiy6CBpKT3YXftaS89O7F5WpEBh
0fNlV399GsNkXfWaVa/ZXoMsXS6GgGww9cFjRaBjmj4WNDZ/cnFeaKKaq4+YvT5a
vA9A6UoiXfLPlT9a29heOwd3tf0v/zFGxDaSK564A5ydawbms00jUQ2dVhKkVUKo
godiC4ZVqJ6olcI3C8Di2uZZhkTIsniPFtDgNgb0BTChKD07dyaoNv4BlpJRq/eV
OfsNGJc1jyinnx/G146alrHoKD0IXrhuDkdQfL8BNLdV2FYBnSarCiRYvH3G1b35
4Nn9hszhr2zO1kbU8zhJz78D8BTleK+GhHCRg2J4+8sSHUkcx6d2TKRbhs/yAuDG
dodjIL0YGPUIpcckGstRELWG1rAg6jqlXc9f/0+Bhfmu0vwZiiAVrFOPc+QOOjHA
+55lydse5AUH/iDdh4dkff7T2Ad2jO3qQDkJIs9WdWeBX+zcdiXcSq68KQfR9dLY
CVn+N49X5ojzwKzGsCFdHx5Ko97dNkyCQaz6g292l/raz4ncBdeVo/RJdjPMprIw
5/bRwcL5Nyi1q3+bhuQznWeE38fpmBvc5ceNtAFHOufwtE7A+16HL5lrx+UGLbAe
thoylV0XpRNnxC2MN8P++fADXfcaUlUVDnGNCMRweOCOU5UxdpESMVhNBiYu5B6l
0T6Qod2A0biT20fYOfKfObwgU+sptlU0FlCtPlQHLymMYXEkJIMsybn1QT8+oJEc
FmQEu6qms59AmEa9PAzPXVToZTT8u/ut1o7vwVo9xbf/3qqoif3GgQA3ehgyLagr
wwNI5usGqLgw3O21ya0OkjkIno+xn5t+XsxFwhCUep9ffqTjpgal2ijshfxui/ps
oym0WVmTC2Pd+Izm72NEjGIEVqC3ZWaOGI7DLyUNDj2mfHv37Xc2Pmx8j+9InyDX
CgZOTOSPxXvT9Hk9sHdyKAVlEyiljmObQ4jN9RjTA6BSjPeUswrrLMpuSlRJHihN
Quwl5xMZ1dL55MPgbcKZqo2t7NjmToIpH969nN74iJtRTd0uL95GG93E7U9i3TdX
cLTBxZM/8ersR8H1qSmT3LpQhK2s671DSMgWE96D61QrCT3cjUzzi2M722ncu/Z7
6bYGG2APh2NBtnpo41zZDefCjvuq1JDkA6TNzNlXf3sIf1dIGcINyQumEkB6TWd1
e7xCetm4Ndsr/S6XqIDIZWlIAMGM9ly0ONU9QIXE0gKofml0OyVkGPOrs5MNyQkF
HrScru2TyRIWHtST4tZLt5D85skdt8epQjVQ25fGdgDEDjNVUMmP6E1R0oCNLUc/
DBR1Zam34/P7B8xD6LGk+3DbOEp1jBTf0vO167/Gh6eZJn2l0w0EReDFDBPWJMtN
fOHfKtKvWlLS+HYHNtWssyNf3/taNMLNmrV0Dv/AQTKHY8vXKU1bbs0b8oPpPkxN
cnKXR+unPDaZEUMw+oqDXyIlQbPSPFCIJbaUCui7WSAHKHgswThm0wqz0OohCVbi
0eEONRypGB4X70U8p41fOfCQXdO6xVykIUbuhbFAWq6pvGLz8olTFkc+9FOm/Y+J
k6QyYjL3hYncIKXyX3R5RyGe0Na7y4t1YFHAMFgEaWafwdeppzWABu4eMbkpYSLg
ZnsDxquXClYQiBBKNH3QvNyGK8dpZPauogzk5AsTL10TvyFfdM8NVVuy7q1A2AuS
0fVPEwTXKhsDzl3sWqWAjl1DeJ0rCQzNxtRM+OzOwRqpowsIiMuXbjWBYzhnfzt1
dWrarAckMRiF+m0TVNSga4CdbDkRMKZnU2PR+7335Xc6L6Fb9c3vSKbd5j26aFnU
cX5zgnRk5tw8eZdlK9YzjUQuQH6a7lX/Qo2BUH4eLep/yr0HjQwLKQBZhCrz3mu4
EkXVDudsh3zywfc1Pvey+vn4wXVWeehbs6K1sCvIqQlFv7zJ4qbuM5vveaZbYfbF
TtpCz75psEF6QgCFlT9tBwo7yD3EFQ25gWD8ziPbcABgiaQbXYWwWbEk2a7DaM97
ZvoMjqMnIqkv1946G5BuljaLIzdayWKRed+3e0sNIK+JwW38aj/VM0uUAmh5X8Sg
t3tDw558SwNDUp8qTXKJD5IMogevqQVigdcj3esybnOre5SnKmvfrXmE2IJlyx2q
wFJ1Pe0Mv70IaM1w19oVqvuooyjYVuVC6oADDml7CtjoMaZwL7xtE8eIK4K2kGsz
jyirlX9f5fLSeK6ixmO6irDy+ESmwVwqIaGWJ7MflVkcI5qy45eHO0n6i2/n/QAL
cHQAfyZCNc/2NDYv19eoDQh+c8PNFvrUD+tB9b7SlpeRMxXN2YiYW+gAdDwc60Mr
Y5N2oxVMB4DoxlypTFQx1gNS08DVnkksV1kBEYbkFYfvcV0v+LaBdLct4oquHo2J
bIt2eNl7C9+OQsssMC1tWKVeZe6zHMFp8kVFKco++Z4uV8uaUsjFaudnf5oSKBZ5
UCs6o5K/W68j447qLXxcy7yTqob92PF5AHQBPH8R3j70n5TKoOZ3qNnMmx0o6npD
W7GQz/lHG7JGCa0CxESnAWhXRKg8yZpZ98hJyCkcy1CY68aokbnrwykG0+dlzA1z
r/lvEDuG52NXv2hkTYb/YnyDYBYoR4aTPthp3NRjbkfE5lcbU3YCsKPHJe/ppQYt
kWLbOesZ0T4ktYbNGOCnyBPnWBJikI/LOCubU4PndaGN78ezGW6aFrF66lKrMEl1
hmOKJ2eBbGGrm6PFZuP0+oEVwcmXt+hBeG+SJ2jPkaxzdmgQK1zJFeRNjzpn0/yC
e3iKf6tKhKsI43PogRFiKajKNBrp3/YslLJJHMIMUA4jK7vzlv8cfHm+d0VxOdat
7FrFBZ7aXxQcKnIiaPOZMpY9PzseFCr4o6NHc66ezH7pm4wEMQfO0aCvITj79sjl
ym4OeVvvr1unQZ8fxki+gg77B4lhnezBCLNMjDhLW9g0KhZyz1l2Vd8l4F4GqkA9
IDOemkZeO2Y12njyk1laAFDRvoxT78bOemsuHNLdRoepos9fd5Q/rOW0KNu1GVBW
Uu/4NDUX/D59bjn2Kz1vWFpyTHdFUjW0Xj3VNQmGH3PxhE2DAuAAd10FarmMaFIW
ncTMg5EFBN8WvTNekGt3ZHNKoEbk7xPIL2XGF8cbJ6XBbTXzX5NvA7PrNDoPQDqA
kqTBQA1y5UqfiK60uRmX70io3x0u3rGlSwSHz6qF3jgajHmsnXy151dStD1NU1ri
3ZUzT8OQCKD37h4GjP3dpdeWXkN+aITN8ULvHg9gBpN5vnVv23PJV58ULsDP3P2Y
6RBT7uz6PaNBFKanIRqEUL/V8BCc0U+A0IpHFugy3RZcM+9MThAuBmH30gwgYWpk
E31r7Wc+9USlwPEdbLUeKcjOs5fuDvwwnKelYkAkmbgndwZTMjTV7aUygkFeWiHD
uawdIHJle5/SKS25s0ILEZZF2KvBhXD3+ZI4yte4bpJ5Ena/1CSEoQtT3d3l2OYP
jDyg7sdF6ggF/1/PJ+2GUpuHTvl6PlcyqWu45P7mGIuw5QqIW+VoT/wyG1ehtgva
kB6J0oC0Yd0AKlqnI/21A+hltOedJqDKqipcGnjNZJCFdQa4qGuEyjEOpECuu566
I3mZb4o/nyPMiOGd4E/5qSTCCc/JGcPP9J/Y7T2hJMQ223wRtljIs5FZSXQcNtl5
0c8DwljESxvaB0SoQWOFoFCWxKJdNDYLLDZE7o9d0wz9u77w4BFjEXre4GXU7rKJ
OU2QeTHt+L3+zoo0gVeJ0S6hrzmCO+5jcZGpvqqXPaxnvd06eRItPl40Bmqopm91
wRTNzCWuB4DQVS/l39EVMy1bwEE9M0LcFLp/FmavCQrKs97uJ9BNWy0WnP/PYd3a
jgMirBfK/NNmnS86GAIyXgaAjbLDNS5xECmTVSzt+TcTV5ZeTtmpoivu5RwGLz36
N/I0xRmWyF0zqomQRsJ/Bbyg04zuX49qpWHCIpIuKdPs9wIBlg5XW0iZQeRPZ5U2
dNiZJe4GG4DaSNdmScqdhgiC0QMu1ySSsG37K1rZmaNSnQXyu/fIiIbHLkG0zuXb
VEKtpgzZyApA47vVPDX2knL4eoPeB6YmHDhrcKSBUfnnFWqHVh1Ik2rziQ2aUH6r
Z1A9nn8pnUnKXYIfrLZ1dqcZcjSzed976QpJ/QfAGKtHBXYAwRSCUfU9e/ftcw12
TNcXSlknX6JueI6u6drlH9LlI6V4Ql+WzRvJzNwSaJT9TaznbujnCDOsd90ImD3f
Ddd0c3V/9Kp8aLXOETishdcvNa+uzcMlbzkl5xcbxtF8W9iZX4UzOWq85mMMK2KW
PDC80DrtAQb2woxBDIBMEj4RChIq3H0T/dBui/fyvBJ2dwaMIl/Qe9sG2hIr+rF7
IDF7XKzWqRPC/J6D6VPIfHjILrPNOtlO3r+mkKwHAUITkcuiJkhBwLGcDp42mhtQ
UGMbZV3u2onhA8s104p/n0FDUUgWTRvCmgKFL7tyL2jXLgyj+wTzptViGpOWqIpq
X/6v7q7Q0DbrUopggbyeEmgd2pLyYZiC+lzfoF99aJjUgzCMQEHXz3EvjCwz76oQ
0b1Ku4aDvF/hn96ovxQPjkKZyWSapbg/guKq8hbBzjb1ZSNSOXIl7/FPcrZ8tugp
5j+uXbsaY0Oyq3SHetM9tsIfb7MCWSTwfE1vnV0XkDU66m0OmR8sOA+a542EHz/H
Ox1UzwZm7AczIRZokmHecCeLN5FtVFu9b10xdUSNOtj0sgk4zpO0kHvipzRxqSI4
lW2A+sOz4hNrsm3sqLFPT1lRvYTiV5FnLdqq+G/rbEdxs07kXfigsTEG2KRRofP7
qJctUOVp+fiATO/s6GG1gTjtxt6ZvWwcpXBnJju3ihtESewyLNEiBMxDpQX7xjas
LKP+H5N/H1dniA18eGcm7waickxNzfTRhuJKlkYCqHrYy0PmwjKxhQdTOC49H0Xe
h9rfSkFqewkwYXuRESJqv5ox+TlQy/bL+3Y9y8PoK3C13Uuz4z3HsB21HCjUkpv5
sxkMZ866RzjKA6X8CIH+3UW1tHrQdi/7dIyQHJIJyxX7m0NSbLn2wgSXaXLZTHJl
dL63tRsmx8NC2FSnHV5ls++8JOFR8jbi9I4Vtv2Sg6F84uhzhSWtVjLELn4dVhdA
Vk3l6qbA933+h+k2vdfyjAOrbl5w558SR0GrNz7CGnSrvWb8h0xHFwWkB9WkdWOm
K7mVrmFFxpzyYxUS9XnRDwxJFRnjpNJx3Vl0g0CdQwhlugwp+KLw+lDZ1/brHFav
XTnBYozWSXpuwYN3Y5D5czesKo07+w2TeFKC/sCsc9ZB805Foi5DLepJsAJdasWs
J5WxraK2n+QJOQcMoVBDcPxMw80krhEgtMaTCZDGX0ZwWE01HIVp1J0ZErTCMoec
t7o5NkRnDkaq8oL2RLssx8pxa4mLMyK84c72d8djr647Ycd6ybmt5iXO+mZgBJnx
YcNPnjFg3NO+IT0/1vce83xt0i1FNlLwIomRxz0xxfGDydyuRdb+E0Uq4zXcmb+Z
8ZiVWLXVnXYM7INw8uV9ySrGy7tAgYBCc91LocQE7rImAsGTEAP+xZR6oBgEC5IE
y5b+6KNBIbO2x/ifmg2nKiHjf3ruTRGidgTAaHIENjMZKmg5ljkAx0QgCAGiJ/QJ
1prg/Jsu5pBqj0LaZ1fSzgZCqPi0DBaQfRUVX6J1Hqv7i8Y/EjjiT3RrpxcbjHaH
xv2WuIV1KK30TvpJuI6HZlMDVULULN9+wwzypC1gxWtqaKmsq7l9jZ/k29lUji7v
LrwpGiGN+leww775VgU+4Ens1C+78Q8sbv4wqKu17w/WRoMGSZYwxIromwuZ808d
91+GoUWOXddmjY/QzMC+/ySd7WNGGU6dqJABPA/Adr+UjcNs4WNqOP0lc3im0wIx
l9OGquMzZFqCuV3+4RP7ABy1g/Mo1ByyYLbwBql8BZ/fXvWAnZqGY9aBIdyCH2fq
27H5EWSJiW9YAmN5uY3oDyMcm8EwNYnS8Hq9qIjKl89mYpQH0GXcamaHrTaHmP0y
2HjeXbVPGzYMHZHcTJjo/ZDii9qQlNU+mCdDcZqPrKh6bED/EucVOA+bZB845TCO
NE50NMkFZr8q7TFS7II95k8rB+NEXvOYcy/XZbbZWOm2r9LBtGQp4SLsbouI2IRG
0fCtuOi3IwztVj+EShgyZXWhby1qxERw84eih5kY4MEal0elFWUjVzSfC3gssYz0
yHPR+hHGy0QDT6zg0UPqXq9VxUJLFh+hSjZbFj/9O3yZb4q/oRMnozLCf+illLY/
hc4cthNXXPDixZDqUR6NYh2NHIXLrDKUV9r7CzNmC5OUV+AtZhf/ZJK2+b923os1
4yT0QE15jhJf3BgKJegBOvXHXqPn01YUNO1OQI+jDZDotkd4myAm+ff/fETFtj5h
gFwPFXvFViP44ddS8QOV3Q8xQrkhzyoBz0T/bGF91BsTfyCdQ+o1umWO/qiWMhpT
lc5Sqdz7wKxdLTnIVszXbXzPOzk6eXane00P8MzRqBl+daz8pQaFHJlIq2QGrP7V
iE2kBs+BX3gfO+fRIDFwnuxkt+VogSe8O9lSygilWlG4AVMfrxNl7dBDXL/geLyI
rwXSmfTX/tk1N0FoS8zicJLBlG+lm2xs7tMteayExoDUC9HXVLYwbdgFktAj8c0k
Y9R+mRG+6dfY1idFUjHLb0fQME+XtFng98YJQgjZ5VUC9N8L7V6B+8HaRJKknzL0
zHpYdF5/AEHUi939OWvtQY0V+xFGG+p2O5v/UaH7VPHGuotyZzB4br1tY86cc91f
FVGHwhxT/jqVdz7xSKRgmWBxQ7J9w6W3YyXx3TGFcblzGp64fFqcnCPV0/6le4q5
wWJ+GD+RymLESG5JCrwAGCFdPSkM2eFqvHIgOVPzcSVyxql59a4w33LuQn0WPTRP
Od1G3A8FwWw5LrLgXDBbhL6hUZguvSPLMbpwjyetXY8g6YbqJ421I3gpErWIHuxN
V2b5iW9dInAhBpKD8Nn+k7a4LQaBmY7fOuUwU96b2xAfesrSP8rUoh5Gr9QDIGMq
nC7A9SnJfjTGEQws6JhQWcAYfJ1h19hL06kTTPeUJpc76DyFInZpRvO/46/wJ1zH
y/w5MZLmH1ZlxLvSXpKqkFCl3AMak3OoNmg8CzcJNGd4S/1mk4u9zCaM1X8KheI9
0AecF4u5fvnDsQvmP0g0V+s6vv7ePiod6DW2sXOufigEgmdcJWcs8YyndWFqpe/z
zJsWef/stMwJ50kBKelJy1hZo4LoLcY42cOD1qx8Hburq/M4zQvWCWam1qLFV+TI
Volh27NYAwfPzEUC8DD+O9b4IWvvA73zX08y+OW1FY1BuPnPps95W5akaMquFkCy
dfcTdPmPvyQSQL/E/qMm9HoTHgUa/GqCHNFHDXP8ImhKc9vNeL7er4Go1MXiKliJ
MUOGewA6y/QVhjxqJ0CdsCT54LTK7fGSPDh3HL5SlwXYzrvEOlEf1rMA+WeSQ4Li
19Wdimg540UUWMILtrb4X6P6JgA4bTGUYBCmF5j5erotdfWWfR8Tw2WhCttwclH0
5gPg2FdNzDEHOuFZpu4LWrBPnCzeWeHbFQJ5BbSfbbUF3IlsGsifnKoMS/iUwboF
t3yztDvjPNn+li232FWoFh0DfC80RJOr9dxTjeZjRGeRfrDsciFY/RucHYoL75lz
GoFObn5+Xbgo3DuBWGusWuOcziSG2h6nFHQwZ/Wb6J2xzVJxtuo/8wuTe9dVKyyt
gocsVf1hfpmiWvcTqE+rXXC+ouv1z75Gptb11oOvlLEZ1h9+hENkxPrPult+xr0n
iUYDOf55PN90aWBWpSkB3w4Bd2Cf33C/d620WXYBvDcDSN9zk3hxpAeo26cSu6XA
MfJF+qr0D0UoO4njHVYBzW/YE8OMfvrrJnjdH+WS+WcRGkW78ppU98Aoxdi4N9nP
/QVV0RuSey+Vtz8R/iZ4BuuV3H6v+21L0O5h8+QR4/HxJ0nJy1Hxru4pnnrZKgXa
pAicCAf3odxmE40n8A5G2FtxBNk32R7PVexj/lQX5CKG9U3jjthkaDpN0FLrYuLo
annXy/90/DYrcW0SA+WBX8k4uSoYmeorj9iNL18pbEuMFQ7lfXMwaFemdqdp4SH7
TqZyfp37otyvboDtDYGVilZU0bsNzRYMPaBH1Gava5GGCFI24Xw8MOtXCYVSmmGk
+czTNmMDflDjwvfyuiBmcIuN22Zt+FjN7tvE5Fum5cpgPRLywe6uG8HvjgdXsiVu
qrAglRolaU/GlkRCKhcWIQwVURGBNpb85KH5N7+6b21QBjzsmYEfZgB13rO35pwZ
gmLCOn/ptetzLrc83UKPzIIL2j9BHOdudhAm0Qf66bMf8YlJ0gU60pr9XVxTmuTv
iIASvtI0bSoqJeWeB0hxjRyKnKf7F7B8lc7GrMeG5YJ6jKbsYCWPmBhotWkJr5yy
UQcnTeLQe5ckbeWVtugLoNWWoUqzi63dfCXYSkn0gYYXfhrS+h2QcrfiiIpm6zbP
4cG3bYYnWjTmpb74X4QHoS3pnv8dAiO0/KW5J27voX0pHpQW3vqP/rBltX15qgRA
Vzza/NBYRnwVzwsAkOi9IjCVdl/bv4nLnLdS7nBIvKYLyvaDGL2+Jk1d1lfi6ORU
40muwtE/x0HsnSN4LnqUHE1MaP9LpCeXoSsg7lPWRe9eROAaOpkxz0jlnGz2MtCU
vsQzO+ayjtmTSiaOt57yj7yXZ9+Qf9rPzRfpsdkSs7sZzI7vEKkJ0Erw5FLrwKKr
8sZyq5jqC8fqjXXN/0pec23tqjfi03p1Ilysd3EFwY8aQ0heSQH/4eGrEZzoxIbB
lyfb7MgEEbph2c1EUYioXUU0WF5xTLmLzTnBoGZ8uv9XnRQYcwIuTdOSkPdEjxkQ
Q7hSInV7fsoIcFQ2aRnwqjDvVmPWc6UBQDaVjtyaCHmqFp/gHcXv9qKDyPxwGuGx
y5AbMIbc3EU6QSCyQ00/+K4PDqaBw71sWZig+bU8NJpHUtcki7OW++C6HP9outl/
zIWrtjOUm+JI1HClB/iVhb3NPDGfBLVREYnOW+pm4aDCkLzNACI9rDW33Gh0G0mX
PR+NUpbh/XjX7X6VnYG5GgF+lI/bEh3fwu/B9YbnLNVGNAyQUWtqgmbTZCH9Hhxu
CH7PCCceDfDT4AOrHGa/d54eYNG4+7OWQNG4vBHPdhlUK93+9EZUFbliuCq2hALo
wavr5nGSfhpFdFs91XZWpe1gOfTZ7T61IW99WCrk3P3WdB++BQfKVV7fZhyuETzU
Yb/HerizG2VXLS1B4byIL2OglFZHpTyBpVDlT8gFmpnJ5NnvUVLPt2hwTD23JlAF
qDV/yoLcNlI6cuS6kOjdhCD3q0VSYZPnxHSft61QxmnuXEU3hWugPlIk6LFh7LLf
F0E3L7+dykSKpf/TcmZ5Xc/P79+LkFabHPX1FUhbXoGw3XKW92hsWJoXMQW2Q+Hb
7BIAl32QCpWs/xmlp8QTTKNJucVHbGba5u1dSOx0hILLOV+j5ACaU7aBW12NRyZj
vvZrkytZ4cT7d0KqfMWKv5joXeEszJEbSXuiIA4cp8gx4dydQFGIohez10lzKDcT
91qNdaQoSMQdmfWbdbpap0412ceZpAx0Cr7VNLxgYuC7r8Oso9pXsCXBPKPNaOu8
ORN1NJYN4azZSQ0QqwqLORrx6/i1WN98c4DSNJItuSX395b9pyUMp+RV5/98kJMp
JgGonBc6/Fu7E5QjiH1K57gDzOVKX/x+StFODlmw7yZx6dsHQdcvCm9JW5m7JXz6
9hGrOcRwpAZ+Qf00zsXLajJ5naTL7Du/CExyRWxv3bk4Yy76HWjIfnpki4nTJHBQ
lD3Kjipl0tq/0XsFE0/y2O8rAbUsKpCJO+cO9hwJ/TNLeFxNNPm6IxEDNl8vxSiI
xHNcu4X2mT+uiS3lb8RuXPyf5GogjU/OQhrNtRmIQcMHIp3aJG7TxyqvfvZB4Rb5
xhZcRIkSw7JcvAH59fDR3fKA2Kk78FUOKaMmryotb1hAsyqXnkwyLjTPID6VgogT
DRvNN4A81XPdPICMHfjg8TEHn46oKooIkH7ON0u946erGmLgGbFWUyJRxB4OIr31
ggVbo+lbYGV11jvq9WULgUOM5l1m/Gdl4quePEwMRLZAcDt9wA+a2zpwBHoVIMio
F3bybHIMYBwF77695oWXvOWX9X1lVkY7zDaNsqSl7I8wY5OUbm0hagPZhrhlWPti
LJxfo0R3ZTM+YfPh3zzqjVjmOPQMili52XgcBr31n6BLl6gHytJOepSdmjJQD5LK
/Muw7tCAqhKmdy3hLNVar/8I20qfmHWRmpG2QsuSZ4HhSRoOIh+r9fRJCLOG/pLI
QxH33FN0FGl6mirbrrGOKoWWRRzQ8I1w4l+BGfho9tHMcSc3k/ZdUN8wg4MZfu34
dfZtDZC6f7rzY1/LOMoQf7feKWXVKOfAUdkxQJGlm70Ap+W9QF+Y8S6KwjKCluPs
LzqxFTXu+K+8rjQo/9teAZpM8X3+FGTuT7a1gkgALNdNiM1evIlwjEvjr546cKs8
X3Wt8yxrVRB47gJ0lg36QQGZlAEfg6IviwtNguquDdZSuDkmSluwF5aGh2S5DJvV
anLR3b1rreZKtvm2fgIdMiyNfsiXcSbIKe5uO83Co40KjaGsV1nbAtFBsVz+qVcE
uCxK/1ptQZquIGtpm8SCR6RERlnJGwXKODMVMC6oQD3HyGv4Xhd6IJOm7kZoUjb5
1HI3Wh/A2c3shnXKGRwY/pEYXlxBDbmBv/Lm38yeOeuOvS5im7eC4UHAiunHM1Vf
BqIJkCYsBNMeU/FJcvdTc5WvaFKym21Gh+yMhzoZ/4cD8icm7kB+9M7wMZvf0v7t
CZT0KW/J90Cn0dk2kuhBJ09CzNUldPH22v1aMmQK/jPuNkskpKSFhIOeRF3ZyLIz
hljIdPKcQeotAZeWq1F+rTcDCHY6s4fHS1Q6gnrjkHcPm8FdHDluqStyLziK3ubZ
7EdEB1wFSg5C2RjIYSMq09gQ/v/7RmdS2v//uE49iZi4VCQxi1Jl+IQlfyU5bLrq
xGX7b/RhO3pbtVQw5Jxlw8Fu3uORgexLUYIfwkd6xzhnd4+jAE1J4SauRuFlUJGR
qlocH31Sn9edX9UkrL7WsNtHy/qOF2cI2lCmC0a5Hl7EXh5tv+Fi4Dx7orbltRNj
mgYxMGF2dZZim86fVZEfAVl84PBMtf8acFgNGoo8IYplwTVZksQr4GGhePWRqaAi
vHly8GdK11+Ma5jUKEsZuFpPYroNPElZ8QxgqW9vdbv/wlEpTR8Nfi4PEBf1Jd9k
HKcNvtfwdpGbSIWbn0tfICnEZt37cruTAFDlfzPDHFH+qHgLXLJsFftz73HjgJRb
C6PyzQ2/+xHu0TalKewJWnIrGJ6LEl4utBFTqney/8um1HBdTPd1kPW6+lfgcdHa
1UQnRIV68TETDQBa0naeD7/snUN5ad6Fauy3T5QxrHLe43MRGAt5WZniAG2SLSL/
JathyDjAuS3lg8te1ePwTAHZJbVgCoQv1G+Dq7FUv7SeTUM6dr+U00l0x4nsCf2y
5NcjRRRbxKMrmx4rempn1yCR28UiKLQvP60LnUW7Z+y2VviKPbaU3/YMUnjhOXGl
VR4XmUlutM9iu3sF04exKwTw8uKDSoiGmayS4yGQ6MMAmmT537qQMjDLdGKfPAo/
F7Cn4m5GgQtID4XwP7hwVMLIHhKj1s1Viozp40O+GQDQ/Nv5Ie4iCTRBZAWQhLGo
l53rdshvsV47imn5ouS34p0t9/gq6Rvc1oABfyvq/etGbRwYXvrKnC74TTOvW5VP
ipkApQkkiR5+29IpE6T/Xi62tiHcN0cul7NNxx37EL5f4Q9hFbktLIe5gCQMnRXk
J9UJzEL4db0WfHA0E1R4XOnLmpr8mSW2AC6bKvatbsFEzcuHi0MlWOS5abK2aEk8
E78W+szI3jC/TmgA/q3JCbAXLD0ogeM3bncGPgmeZJTXm/vUa66uL3v28yZlxBM4
5l5hY9F42jwMr2JZ9k6wv6WgTxv5h0+eiqYY3omgHLHDDbyfq64YTG8KKGQmhWLi
iHJOsLlq8hj6L3MrjyXSGyZ+oAAfs/8y0dQQUILcJQOX8F1LYoWb+BnHIEuDbjLR
Da6q97lvm196J+U0zim8wMdgzvunxBAvnLCZ1irP4aase7UlAoGXLlR19OyMiDJX
cm/net0BFkZXjUcKWXHp7xzb/nmBpBYn40dcWL0zU77COZT9S9WYNy4KH3GeCtXO
ndKCgnZKdN2HcmQY5esNqykg3QJft+B+50XPXyjKkK4Z8/UuA4rN+jBMahYk9bs4
B8IoWIW7Xyi+Tohq/B2Yw20tiADdtNhCxVy6E1O3W7ne0qRzd8TmIEkBiISkSJFU
Ojpesx77EHd3xJ/MklfoXk56NnwYdK56eT9d4dP2n2RiYaLqHMspNW99KzYZbDuv
T0HPMA58bW+mgzrmbcmVkLxszin4B2eX8hVM3iYGcKqIlpOu0G3EtVQtZt2jBaWQ
M6MUeloxRI+6b6y6wWcn7qdLel52gVgJUQIxRGHJqUOfkPq+0F6vkx9sBbMI/VVV
W0UrS+z2GwGEXxUgTkhroyG9a0v3M1gXxJWdnKhRDezZTKPbLQUODGFSphS6bvMK
F4PYIMfuSRQgM23k9I2JaL6Qd3Xxx5/wAWgHhAy1/8zhdqsXEnKgzMi07KX5qTDd
BiXLaUW6KU6DuHASzgmSHazARluCBcIKui9JbkcDcIQ49bO2zLTXmwoCV3fVD6C+
csStB/JRJmUOLQ5iTsfXOXTJJuoOSaW0Ca5SuwWWm7AXm5iuR3tRsa0YQ1OCK1Sv
e8soVIlz13LdYhD3LsoHsVZJsV0Um2pjioitTIW8W9P+yW/Vf6jVxuNLiNUkxdeZ
QNIOCHUj2N1li/v2p1laQDK66cHC4jXuLZtBwjvI3n3iH8QfWYNZCw+tooSuYTtE
oIL0OadYzojyXO4W0MPCj+Ko7mgsBA0Ysd6jsQ0OixHklZnQLF1wKXyJcDl5rciR
KEh20AnZSX5eaVPWR+qnHzQIiBv6WdDLIA1aIEEKUEQV5acWduHtv3ky+RSmS5J9
AHlOloSs3i6UveHE2MiTxuZvvfrGXSRyoLLm5MeyTXGWzaudDLsxXJhmC+QDWasu
yJ9VXsLkikahBufGMKAfE7lkAmV93v8SZOQSgA3BBwNWmlgEju6pBeMZSK8Tg5/z
gPb70uSepzJ/5pPGWWhrM4qWUT/w4WEHLRACJ2V10nt3nMoMzF7kfasaRc5WN0lC
otQM6dbly+J+kDyqLk8Ug1mQOdh/Tw7ZxP9OUk4fB2Ov+F4oU+W03aC9cJCHQ4HX
O87akYNcReK0yLse1PjaohfjHUFfn5IPDgIPfiHhTeEPHj+l6dZvbXF1a7Ff+0lX
WopylLMFM4q2DjY1ev+M6cnHeamaOFwTyY5o6x1SeVB0iTodT+97r26cZLesWTMp
t2uPHarOwhk5mOqqClbjntyIdcytM9yBC+y8ynj53KzihDTg2TfzLx4M99KoN95J
etoPZILOyVew5mQP5f1H+keZB88pBIKY5mc93V0NDHniAQFKgasKwrGisFcTO0m7
JkppQ/YGuhA74y/OGlVSBUg4VYPCAYXaVxRna8RVIg6tcAwJyVkmeWd0CsQGm21+
TxnrmzkdTEzrAHqG6DAVa4ZsU5W+NdcDSBmBaJ7myc0U7H0N45GHWNHmhh1Gao9z
mNADVcxXp48HL6P2MkieJr4C2g8ZrgD+bAWwdUIMzYyotHvrAYAMHj/q8FKn0O9j
XyYjpBfycAUe15xIBrlagjEOKrz7GVHEnHD0VgNzYx2Opf0FRNW1Pb0QiAHV3jjB
H4qMge27MX7mE6+BcuEEOFe5ZQDY4ZMKzi9IRH2RU/fqv2xhFuoYQcMP3oKLIImX
LXpNPfWoLe9DhK22BvbsSdXltlZ2AtERGfhWYe0PZt5310f0ZsUZuesndqSOXELu
jfjrf3A1cs2Pn8fNH4CavPDNf7YEuE0AKfthDE8R1V4k9quTx+t2ui2d5E4TCQUl
Ti6VsGi6+31NJEvQFyFUFUCJu1VmFShS8eLZFU3Ql1UKxc7veBt2dnX9o6PkIunS
zZ0xcV1nWenjVr8t+IhFBlSEqeWHpRbqRKggKqJ/Jp4NF0wq5PEjrntcRETZ9ybl
Hdhs7Nt1/ca3eySVqeWKc9OIZDVfTj7SgeDirFxqlLT4FYIYOww9PxCMCayhqUj8
6BxnFxbLzIKniGHELHz/5/O6PipcvHzOzM4GPkxv6OhfGuYUg/D8dsV43J9VhcqW
E8LOotikMjJ/3S0ZPAlUUC0tXwx5fy0rjXIJ++YJT8TpRlbD5eOffMqQFmbqIxIA
IAr/KF4eUYHXoidmcxD4sppzHaIgDL2YilPyHVXbp4ndIlUUxhs2I8Ar7Ev1O1hh
M93auj/Bx5aip8Hfn4DOmjIIjqHfcBs76O11MvKkR2aRV3masKJXBpCl8TfRQQAv
GvtCmwJAbIox9cHmjjPNL5HNC4DLdJCY9FlUe2zaVWACnCR9oMJ3xapG5cjrWna5
ZMB7yZwGVW7RRPi9vqFc1B+Opxi5wLS1C39xVWv3vTDkr1Nll/3Kc9pSrLVloW00
0DYghnXddbkuL4n+7EmCQyzbCU21HpLgQeicQlVG2Ezvo2u4J25kBgK4kSJvPivh
L4XQ1kyNGgdf3okrsfxqU2YdVzvZ5+V11y3AzZG6MsW/ADu9TgDGjTqWdOhSYS5X
+vEU90YcEZFRNHXXza9mdnYrWnAhaTHmDX0c8RNvtZXhI3rhNhRhz5CUTjVtotFj
+UmKAxfLIbxFGtuOKhb/gsIZpxE+otF7JQCNGGBTjONShq9b6vsxvnJkP+1cNHsR
ATLT5dwi0xeGjYAhX2xj1WdXOOa+xpvIYlW+/KdaddsGtd2cxUQC8X20vbEo1BKd
grWVTmyJQdZPN+GdeB7LzpVFn5tnd859FVK+h6Pt75p6vfyiUWDtlkWL1DQPbc7D
XPHnrEtTVY2So3zPiM8lj7aAZiBaI7bQUucR3W2dQWna5lwOMFBAmLGBEjxUA2BQ
WJSAiEyWUBqxTWLjDVHC4OlziHVIT/JVunvQHe0P0XUN9QRqJOUp9oFQ4SCRaKeh
uTm0VJwuTzfAZ7CQx8rHmbE5EbNrty+LTKd3e3Jio1rUeKyVN64VvTCjRX+9FUTq
bEvHaGzhZezi3mTvx4cQ9P8S2w8uZegWcthRCy8vwcYV9/Vclzn4cZLQNCJUucmr
HX+FuaDivKhxZl2DRCC2geEKlC/RqWEz00yAbT+Bs4IqX8S+dCsVyVmZgWfFzT0D
ZfJhbzzc26c1ehpUDUgjJvOJ5bGUY6iU20xZAT9qeo5MtkZkG4WDh4k3caWJ/f5q
MyF9hKCG/vyX/UHyvuRfaRiKqSeIGBKNM8PzFVRuvdK+O2r8WfLGE7klx5LgA8HI
VKCa91XC645Gixuuu1cMxsDkQcz8uH3SCcg5Yrb7ursV0yLUs/nEqW+xcnLSlLJR
jIP8f+dbztmuGQRMMIAEt5GRsLuno0YXlMiKgRlBNUhCSvlMqKHShxHPo0F8fiCs
Q7mIrL1/EovE5/TipSXCX6coHBrZc/OAmRCOorTymVLdlH33mIHRjtPAfc8Ws+jE
ndzCJkFsMnMzDJ7vrOhDzaKH5woQE7cn8fELWJbtdeySVAIQHuiIoRSHjHnMv3ne
gRqtMsLsNqZOX2eZalVHcijOkac/4/T00HuEryWiivwIV0KQNOqNpVg0En5II0UC
N4g/g3SbGzkWaEg1nM5e7LsSCFTsGz8fzhOjaOWkCBcsqVd+N1abtt0tfmBZlqMX
zigsAD14tCZC96t/SFlMYBaMj5PiQG2CLkn+807knbPbTIE2UdKh8L8M+1dr/zuD
nZGqdrixNdK/wrk/Tlnju7x0fi9DslCMQDXBGzcxl/lcAZGDrekplFFJphbhKwkV
SxOJaFOI7BR53bzrmu9EOrd1JF62Skc/O+UBS8Y5yyM5DyZEHKSD1AChImm5HJmm
v8d4gvOkP7OXP7g3/HtN0RzlCKiZkd6dqymoCqJme4mUL3nNi0CJB7Fy/yQUbgGn
pMhx277rxycy2uzPt0jlNPSx1sqv/+315SQSjrSmMFlLRdSyBI/8VdK+GlXqNjt9
GWOU11SMhk0W+7QnkLpdeK0GXGryjojEBQO0Lpy4LpGXmNAyZPCINXvTqPUzfwYs
nGFluzRunLDjMSbPcunZ/bE/GCRuRi00zsY28T2vdD1AYaUGkVOjS+zyvpSYK+aA
m4NfOj7YoTVjVTXCZkwDsIHiNigBV8t8t5HtXmEJT5xRuplYaI8kzi2RkXVWiioh
G7JWprSvwxC5HrO/U5dKfuYcPG2Kz9pszBmJ25Ga3St5uvxaHxLpInT3ShOSiGRY
cbtudPA9PRwLzaLuE2AazIm/Mmvr15zL2UDFrOOwnOfsSsSqNxhj56Ytn2SnF3fu
/xZ64Rq0Tk6PSjTXK9T3pXj8D9JGLvZqlYIkRU/AZnSQJEh4mOgZmSi8AwfUBC8h
Y1uyk6H7KPurhXTj7/IFHmMioUNcejhGKaqy33wnVPCGz36Qid8DcKh5I/DaOCyr
qsAwfFBGjzv1sldaS4ZHPTiQoEapHTJcpQFCdju5HRBPwWesiI8bP8jCjhbTWDl9
Qr9Q4gRuKriSo0NKK56fvw3kLGG4iiFvC4nwNrzXh/ecmrc/dcGnii9Z0Ug3td1p
HAg8+sNjSx5DuIwEHrL3a9RNNdqfcpy0e0Rc01vztYRUdPNZN2/fuiIbnK39tZ1l
oSt7/K+aAtxbWn2Z2vJYCJVV5jd3y5F3+r14aukNBts0GKByoHG/rGDmkQJVBhf4
qQI7OADNkjjXRcZhuSoBtTjMAVCxlhoYgmGn8PpMe6oDdWtzP9RNogm1/9zSHbfO
6TwMGRlGFvYKvPv/Z3LO/R3qJ/TFCiMF3n83GOUjx4zYv4Y8g0CqHXR8M8FRnuqo
QF//bNRFsOptyrXSfTTnCXm5MH+Ulatw4fzabwIzx2HXqQHlDeXNnqdKaibgwcYd
OCFP8QNSjzFKih+G6CGviKjP/7R/LijfmPDDti3qY8zSobJ2TXm3WxoJUQ1AqFmN
wcXfaHgU+FYKhgj4uG4pY12Nklzb+NExfcIOAatO20qaaAfTb6jLY2AfOyIlRmf+
5of+epy3ZMWPizWFqmHuQS+HGCYPFXfKzBWgJzhbg/Ok0avPH3/aHOcTJzYM6srj
qdHZf3mPx1lwByKS6gVreJcFGeDKikw4dDfaeYoBt5sCipRiAXszuF6ng02bA7Hq
bfPM9UsYZYwXNtzhvf0bPUJhBArQAaLQOjnfbKG5hZZDdmVxKZ7Oc/GrzmgNxHxD
IwlVnh74YncQfoJlvjonAcHHjvlEtZswXcqWkXgipIXlbkiUaj/cYQgGn8zwklL4
mQaKyVkAADDO0V8eJw6rMSipH9cK0L2QMJMqZrY65HowmFPaTgGFAvGSfAf+L6+7
qPabBWVYUTtxQsWoBvgboQ/j0kovARTT+yWwGeCxWqIYPEKD204Ii+DEzrrNEHnM
DDENSkNkztcyWEikcmqQOLVEcPUyk51M6QXfzcaFQnWOGENjp67/Y71ZKswqB/G5
4fKVJ9PWQ7vk8dqwhe5BiTLd1mbJfixU+PTNrtWmI5hvO0cNl5gjAorf+aiM286Z
d0omwjAG6QulyZZSB2f7yGqe86sZZd3ktQObdnn/T5+CLO1/QgmD8LjmoO7bCEQh
bBD6xVHx1s5nmMu/YwLDTuSRcPE06wdxZyJHiVX7ptXGBNdclxomeK4B87cJrc3b
8sq+xR/s+g+FBtMoFFA81DgXC3U9v/DEDr7h7LY+4485fpE+i2vyne9jAv6/2wKN
pUTFlggVxxQxcm6SVapZZISHR4ks/pH9N3OnN8EFeR48KcOO8nIwflb3KnRPbpnN
alriOwm29aHPc8jdPEmQssHChZGaXEYcaFkgZt0RRfEDQ/YlgP0sbNFTbUj5YRGK
1FOCTychKWEZ6CxYOt9W6FOfsc+KUI6BGwmWGx1+kBg3LZVj6Aj2d4bk7NWmOul7
QzGdGP/1zM/jTP/2Ln4asrvoBHiIdKHJ3JZD7X+hBiGwkE/xGqqhMxO+bkI4inTR
g1m0NcNT88W1ljdKYFaqQiD/Iigp9hi3YyvmG3n5MGuf8ijXOXR4nJchV6D3/O1B
z8pg3AfAXVz4eIb8H97h95PQ0iwXnUz5YE6YdzndwHjuw209PL5nAitGJ06mfMJr
k/uCONeSLsbsJKTL1I0SYUNrTFT5KaiwXDIzqavPRBcI8HcE7GOeU5BbGCTITTye
VKQjcWCVzFB6aQlG6qMmfsjezDjx52pHQr61GFWtkzlcpllUor2BY1hjS+KtAZrO
9QiWHfuDeqO1C7h0ZmG2Mbp3Ht2rSUMmylLMErbi/j2tRqBHBZG78J/lhu/PQMlP
Fomv93Q8/rJGdfOmu6HUN0wHQDqGQp4rNvxUV88F2J5fqDQS4SjWJx+U7yzmpUoH
NrclA8DtodlhZ5GBUVuGnOUF2jSIr9IIhASBl+u5Lt2Of32HaAE4SOoPFQjZjV9+
yewtam5jNGQ2c3KctvKg7VTkv7fqAZc2ved/H/CFpvRdhhOZ9i3j+V4EcgZkJJ6D
/oGtMcRwsPExUrxAU5pS4eFVhWRuXUoXLOHxB0XzfqFKbv/gWkBD+3pMkr39NJ3c
R7t21nFb2/VNternmICrk/NVa7Gbr3cmQIUI3fhRDhy9kcDUyrzOCOwpGzAtMJhk
EbJ3D4Uh6BIvrqX2z4pPv3LJr2K5b7rKye5HMBDMgN3jLXEY+psZDFBq22ZgpRD+
ZgcegLPdosdSfZzU37Ik6R0IhCQIoz6pKt0R8/jsxG08PVSlH53ZsJgv7z/KmJPz
VqwrMo98N8EG40KtMigGjKuWJ6Lm98jx8rZVBOML8P3CfGe1zioToU7nKk5XYicu
GsLkVK3eQiIzT2L9+zlMx3ILGLSdtcwjOEkD9vykOgZNUQgkStiP7+rBC8SfzJJh
k1lkO9KgOGMHUo11t887qaufKq3HuVmn7+0LXLXzO2oJ5rfEV3XE/njKcbP/8Z2d
hvaNVrrsJJKyFBTmkdQ7/9BJ+WUWi671GkpdLMrBDhsSuu5ydTXojjUjv/U3RIuh
vmbTuioxPOOLmR6A582oZIlG983fqerq+gsUlWHpatAQmYuJ+gbvMAJm/oAqw+y+
mixcbBottnnwyYsU1NRA6ujZyuJeQTz/HD+1V0IWf4HVD+WaKwXYS8o/DXYsqEoF
qBQfdVa3rd9Ff6Rn0PVF3GwM1/mjx5zDa0m8QIOY1n/IzYQfBK5TDQWzY3enbzKF
rYWuX/WVyDkE/RsG1sIhk0KiQA025GKsJY34FXDzd16tuV817ILMl22rRzTuojqv
b+DSOKodIvdPJn32d0pNuNXaZy4Mk7i+6nQ9PyxCe/WbxpOAJJxUyo6QLp0bumBv
BQjhEiOtGttksRLXUteftLWVWevHucyAKZEW1t1XF1uDXvMplTqzcnc6B6cBSz3Z
cNQBHfNpnucHjFobFWzbimcMECyFxN02wfCf+X0TD9DDsWPVgdvYz0Ma0z9s0q2c
MnB+5GPVkKqbWOGGx4rsmY2ZUM/uhKqRzd4tyE8NE2GFuHcvWjHJUlJPuOjW4iKJ
5Fez4l/KOmUorXS6UjOruU7egxd2tt96EpDaAZrYMqZgmOOvQaGRNf58Zz1Ff9mX
eX3oVh3a24EoBz+XSpGg4IxL5CkH7JzztyfO5oAreD3Dk2GL6zQ8cuHDDbo8oQnP
bjpB9sxr9lXCpVuXrZTdhELpVZW/khJtrdIpZJYNCigkROwSDzUKS0TCb9JMnuuO
MBLPN/tIYiRsh9fJDXzgMNtFLqKxlJCE496qUyCIOR9gZb2ERYu2Gzk9ZvMKkz1o
lsPu18YtVpdUPhBZize2jHnUlBP2vKNjgQyrbxGReGUm1K4bGoswXSTIr7cCI44V
Yj0O1tpC164GMNRhFtEMTZH8ENAH7mKFSX5x1ETd/kIsQwwmoJpez1kstmUg2Xxg
bgJvGFXUIJJAM7ejU431FzFLw2PDhVtqDm8vBUnBW05Tpj+ktn7XpQbrzoyL7qoZ
Y3IogKRyVvPC2xeNH6hKwwkQBsRP/dZOfdj026AIW+ZR/xbowOrDNwSa+KgdGrxH
lobMEXR/6hLZ26zsBYpJd3oqsc3qSQV6Eji5RV7uAIuavbBLprb4wRdpYtygvS9P
crQkmRyi5hrCDG4uQzniI33HOo7ZBEINiQEG/9XSz8FuSk9AERPHGb6AwHjK3NhM
lIDIiFolupcuonohBX+NmgRK8INe8kax7ViHWl3sMdZ7sJSgsZySR2onOIrQjWOH
nZoGNDrCg9NnBxdzgywEpmwrtopL0tJBL3r/rays8LsT2DlDCiRRCjwSEorvcf8T
+RgxO5+TLjpQ+gLXZ3BQbeKyMIgg9wsj5VYggnxvQrC+hU6r9ldBMODrTOEDm44N
AhYw3LqbXSXJkm3K51P5/CTxcH791fHvUWFYXr4yRaQ5kbosv6mXlobqZj0LpQRq
RFABtUwUZoD3SLOENB1qK2bhUFoLMzuKxrPHehOH1K6yQRdwuBmgqJ5daNjSdPjn
q090J/Y6FiT6tvsL0LPysNzOUceWUR84XUgTe5Q2e5VAYCvLNk6eeCxV3IGmbR8H
orDfzWmNyRYwfJmbE/WJXjY3BTA1JWJ4++nDSINB5yPnz0XGSorVsw9pcdffjqvB
49ffYhCHB72ujaIpfhumwqXTeQSEQ8colvGhx9soTJ2rBZhQ/C3uyWhTw6DpWuhK
7AM9Jg28dobZgdTxtfQ1FrNwS5yxF0L8NJFARU8PuRZ/s3DsO2Tz8iqKtZydPIhe
PXaJNnNUFq2uUymnkiF+x2qS5skHA5QrTAozDpd9HuVy7wHetps2hCR6OteKY2dN
UAPguJWlj5zfaSDgW36TXy5buvM37cHLh0yD9e/U+sMCVcm+a8As82MsBqzO+glK
hMqMQ3DsQNCPqW8HAl/myFiENz0KpF6TUeP0tG4n3xxkYzV5l2Y86PLdpw1sav/u
N4maguNk64naIeEy4YuPus220o1J0Y/aUJ6Q/0HrxM1tx05YNwGK1utv+ZaMM3p6
qjHIzzaRKjLFKPjMUaWWrSfZzpJePR63rBzcOSiUg9CnMw1Tml4hTQUvJRqaiqFY
zjWsmbrgnl7lF7+e6qn1fBES3e/+o8+ftxeFbgWHgG0+RCtk7Jy86HVZ5l2F9Son
qbn3gMNlTRWZO5YCWysnjnb8WfxAwUe68uqQftdeJ/CLnf7lNJ4SF8OgKlSD4l/8
wkSskzp6rr3iFSOedQxkrp/v27ov/BPaDvi5+1tgjfgVClpKfAIeMzgwkKxj+WbU
VFxcqtFLr/RbUEVxMN3IOi0znBrSJLbQAn0AZmF5TNaUf2roszW4gm59lf98gr9g
RRhhdsaryrICGFp+Vu6xr2Z6nudPh8lvmtyKqxUlyFMjdHaFeuM14otB+m9jILF9
2RXslWgndu25ukXbOSu17xyA9fsVgwDoxxKLBoqlm172ug/2bs05JZ5g0ehooqh7
Ns3gTk0BBkSmn5pEtAuFO13n11199fqhbPAr4p4pl4CiQSsud5ivhnNze34YZeGe
IT6n14SGhFdAkTer/R6iv3vSpJAKwIsywjdsndxfEO4eKoOFlprNI2O2Jkg8Q1bR
8qTuVE7zGHg5EzuSm1AROJLuFpAGi79wwlpy0tXrGCWP7xda/D630L232kOYMnfs
nsNhRZYA8RtDdmm2NMzlH1ZoQEjDPvPIwfK4ej1LQdZQnKhf5/0O1lw7eCZHZ9PU
zRy1K4dpCt1ao18O2Gb5S99Z14t+P98A2ay63CpdQngPZY7tb9ilSj92TqmVIhoE
OphfLc5kVuuncFJ2PswVNB1QGS6PwJQ51fA+IfhK4Znk7YJp0UhYx3POh4t8KysD
/o6DRbhW3N39OqodpOnZHL739vZkWtq1TBdz1jnkD5m3Va7CiSB7ZYaONk7mjWbV
7i8KnwhNLZIjSmYw875ToIi3zW8VuhsN6d7q4qNvpYPM8erLTsQabXbXm4TNgLSq
Y9+qQcc87nk+tqS/RIgbyxuvwPyseLN+B2FQrUM+dcpEiOYx1vv+QsLLHsFb3/Y/
dxfj6m7Jridv/ukCjme2pXGC4hy976tRxDEQ99/pEWrjhz6/goxIj6OgViqOueX6
NJmdBoOgJdLTDas2qsnFaLPHMaO5a13Q0dJLbmuHTzjEo1KZKN69Ql8ymbQoIMMY
K0besgU1OL+gZAGZpF/szMFwHhdI2ghHUcTlCg83UInm+Vnqh2b5HqvtsVLWd5MK
l0nfONDpmrurT/BYNDRKlZ1ZhyRbB/M0VWZ2b+XOe78bahu8ydU9PEIHbtE0mpj7
LHXZpfa13HO34stRKhtrfq9OBr5ddqvbY70w221KFe/7vp82xoY2ncoFzRer38Jm
4kyJcYJtYRYWtlWPz/Mgw8YMX7vKoVBYPgrUd+7hGfQDwldXw0gWPR6jn2qAEFF7
uI8e+VriZsROTipN9b+mJUvnqf8t+8Uf17Cp98B6sLOxZjO+raWrLk9FZWa2ZWhY
5kqqrAN7nOw0QLzpfgNVP9my+7+OP/ak2FwcUFcvjyZWLbaJfoKUKTqQojx2SIoX
ZKI8LK7yJZ/J3W7S9+xl26DGCQr8bCBoJY5NI4HgExMTWZTcoFiEMMxNZ8IrlSR1
xISaby10uqW6wP09UBFjW6hdp4KANHSnW9bbdNPjPCZNCdBaIez+U6cfdOWLye+u
tK76EiOb/VEGfXxIcLTDE/zMuAW/ZpGdg3qJO3P3JdddzIhhfTBHUmIeH5HAkIDS
+DifKI3xYo1AZlAJVPiHYj+oUI1o6/yIL5NqAce3ORPDNyv+3IOXeoKwSKZOqFe3
qWC/d8S/skk+TiZdDDn1qKByFHUbbWPYialVZe5baLvipJ8O8MjN7RYLMFymU/59
5GwbIvHNmEX6IZcuqVn53ydwrh1dLcpXxKI1Dpw1lyINCRL0LlAgDYkQg+7VzY5K
5Ltlorgn0rpQjc9pWjydrwRkbxQ3kv4nOrxBuXvCmZYfuNHovnc5B4QQ7aJ5b2Gy
b2sDBW326W0IptdikBc6c7+/hBolBJpVIaFFsNb8VPyqyEKCexFI+dR3s6nU/JOY
LHf5CD+Z8ZfAKPQ1tE6ITz+eznRVmPwR2jK86yIPLC32uzALDotcMe8fJe7fIMAv
gCNPlOAExXtjPOBVHEF0WQkFg9xVNHIo+ZC6VoT6XtnfWqsqUuLogBgvobJHcLaj
6B+zL4+tZhdTh3YMiPZrHZfI8ZgLwyFzPywjF0k++ikuKYusSEkORUQLfyhfSpn5
gozml54EGl3VKYONPZmi4Wor3KHIN31VpETWY73G8Ab6ZlZiQV0NYJ0utFdKlNgL
Ik6oeTh+MHvfWoEoRqYVVj+8Buij73QeSVTkXKnQUN13Tmtn1ugICdgRIn7vqJ4E
5AgcC2Ch0Qj4kD15I885xiRzEPuJfHMK/X8GI+IJLKGxd0ZhSapsnitGW4/QabXI
1GeBIBU5N5GQyZDuOxT5fBS0K5WzcAgx+Mzqdm5vXIZZbA9VZmIZ/n00HyM3MyDu
mEpXlUZhhObe6ihN9U4wOv7ZsYc1jam+oqwcl7AOngf0pFSg5Bmxrf6dgV4sJkRP
36gDztmsqyXZmLMkzMAWilIYuFpVdQWRyZMAtl3y8q/2DgJGxK16LEq9giezSGl5
VWHgvai9uXldAocRom6Xmy6CMbcbUod+v+3lzsNd7sGOOoTslvbvuQfiCJuX41ph
xD0e6qtLPvzJaTyYzaEyK+iRCnQS0o6DikW64CmpnNpTrge1ypPHCUxOaeQpoPH6
Eyd8ZZpUb41ivS36UapbFk3dzYRW7quqbJ+e9iWel6aC8UXl0SxEiGHTBUKCzWuI
SnRanOpJfDL5yEQTaYMQ71/g0K31yJe+WQRB+eNyUiT/uJHa66sfvS7LtYhy3u6I
FmiSB3V15XK7KPMXvAubXEwGObuNOWqx2VBC5M0EZT5TF0S0rRZo1xQVtyGpzwq9
xLlj6V9wK3kRsPMoPWuhdVazCrQw3Tt//87y4SYT5jtya+h1SJNUX00N8RoYs8tc
H4TLITb2ViZAU+UwNShT4kxBIbLGJX+s+oACSqqx0SKiLVbnOtnOePPTsrSKU+QY
d05Mz9iDPx2xLO8pAyDKdzrJ58cufUdadXLH5Sks1Dz5FIwxp2Lfru1T984QUAmW
ekMFnIbMidgkT0vz9K2fFpUpWAvQRPgPW/gr+BTZy8FzIraS66waT+o5GG1Z74eH
p6oQh9rBHzuc7X4poa3CyYTb4AKUMU7f3qIUNk9ounGuBU72JT3dljDQFIUza3W0
FBUA2oRITbjfpQXAJ9XmDBgRHgR3Ifg1k7xSqT+saoeJNAjST1Y2lK8ER+19M/Fh
1HedMCJ7RatOqfz4Wzcci2ZDH/E2D18c2HoECRd28YLBEofAF0oo4hLjJgwHqnPG
gegl4onCtjPnGx/QpJEp4bG6+RmXmpSrElYU8YNL4OxzYvMj9P+OMQZx6qUaFKh0
Qgl5eYdbZhM1oHkxV191B/oUo7TMlIoLduV564rOxohERFAPq7+UE1hwSHopGNjo
FsFYqJXVM1N/vMfeznFrb6Fu0aFSh7yTJCjnkm9Ib2w2j0TO7JFCH+SM+UHbgRA+
ud8KzAaC14s+S6816mVQ3hSDRW/XFft+qFDPIdfxVHYTuzvD1je2iac37XSe7QJH
N7GkE8GrBOxEBwfMXcqc1+vNL1aAKIiii8mNw5d3wypsiQ/K+UsTs4ozuoUu1w3W
B1DdII6pj4I66WPgUoO46oIIJTUDnTCYU9qcqXTXSZTlcl5ry+soIOzHOE8tFgDn
p7rKqufZF0IDLP5HqEw5ja+6nDwZKUuZnDaBDiqJ2XXGZO0iTvxq4z0BjBF3w+cy
57WnTEK9caQIahn9CEQu6YK9+fmDKyW3TMo83MPU4TA6dRSjwCT/jX46wkf99Czs
owkLTHvjneny1la292PONMQQr3W805A2dtisGTNvKCvFOEcPsPGT00foMp7Ro6xW
5jT1itzIoKTOyS2WL6iQBK5ohIlAWr4FvNn7jYqlmsMNWl31+uiGNLjawHUpOOPk
p0O6yBkIInuSYtmAs6e0gq+j2hKboRBtEBNRWlEma8cazccA8cMG0bxa6eRYixhl
BUi/uzzkSTR2S0JECF5p14F5bxyZtBc19YHgH0FDxsfp+TPwOuZv/dkxjkvJKQzD
Zs+4WRsqLJOYKTZbGWVZzH1Yso6mqz9R0JNgXcULAr31FXa033HxxMZlybKoIYCy
baXoplzYpZVaCPMyos9H/vuYuO1Vd4Di4GrVyakoYdd72E+S5TDK8aw6wdfmzvGW
xutmBpdtBMEAeirRrRlKVZ6Od8tI/eA9lcVcmCmBSO5Sx5qxw8NsST9sAc7J6nC7
k5RMJYzKUK2xC7jaIKADQSocIDAevScmivPGMsZCgkSMzjCRH7Q5IdKzg8gdujZ1
M7PCGtBaw8dyx6QtSq6wT1Dk4kwKIUSvNJpUnt7Yafp1D8J29/M0ChzmUk3qJPay
1+cuZ6MVjVN4R5CMcIH3AJv3DUq6ya28vgUNxwvtQDAggk9CpHZDQk33wTGkJZR0
GlwOe6kiOis2FMmzjKtg1zOFOtRQSPVdKucjp2NmdWv4hWdvJ/kMajBHe5hXdmmm
YD2MSjEExS2qExB3Qhv2dbCeq+bWDu/XGiZJ0pr/lL+Zgho0t2f5GKiKKx+1h4xz
S/42RvVbaRrTeFIqFY8m+YOqnz+ehbO3ELsReGGPMNA2xb76OWdL5Emmd0SBAFET
NoanNWK7gKYQ1nKfI3SElWLiF2ib3ZQxBtIs3JCjyGPozl+i13gU9cgK80rjHl5P
mmBL8B0AoB3th7/9xQMG1lDLSe+tGIxnIqyH0J7KmI2NMXxmmjasYsYSzb6Xlsm1
4P8b4aK/IauxGBUohn/WbUbV+71tHV18TjU7JeRGIw+v+9wZXw7/6m0jC7OL8E04
9fXlH+AhFRM9d2+b3hWb34xKcDrDnyt5MZ/CTa6SxHAJN9T1/JaEZQKSQKipwL7R
rGLY1sp1QaliLpf3g5K6HiIL48IS9Ttwz1Xfynj3R7Lo9r923UMkKxKU9/nFcjBg
tqojlBgTsvfuEJc+ZcW47gxPb8V2+HmXOQbiBD1BeYPH43bO0tGel4bWK5dFio7+
u7nVH9hncBNME+9Fb5yjbMLIP0ifNsm2YZ1SCraEQyYM/kYaR0CBqPdlh0mwIWmK
5vkWyIBheVLae7iCl3+cQPqHZ1leQyjGbhR6D1z3kmNB2HbG5itMn2t38YJE01W7
hFVGVem7cvwiSebpsNHxLsYoFCg/NgoUX7+m3tkK2ste4RPeUqgKxhQJ77Yx+eeh
qMxqe3MJco97nH3MbWWqMlQ6ihy8E7RagtJE5gr246910ffDCLRX6eo7zvGVb0Wy
Y6N3T9ItnMNcwWNWM2IPWhptrxV7srh1r4W1saJKXuoI6FehWV2dB3CXgUpwuViO
P50HRbryEiKosaJ/akz2Dk+rr6vg7pzPsvzbwc6Vv//r8V1R0zMXryfQ7ZO2HbQ9
yi4Y+87Xox63Ju0Pnk8qKfXdx7B1PwoEbeBduRfajW34vt/TjHdjRi/f884H/ONm
RYEgG013YJY837arFAsp9NwaVA4lq1S2bLLCrd+ItoEyCSQNpRA+J8q0lfN/jcK7
rxXRJ2FYETW/qdCx326boKE1Gjtfj/CtmeRSpM/MU9FFep+5AKwfs0hHb7pcKArv
1l3xywqCqXQXJyCOcfu+Wt/8CkghYvUdKOpPou1iY9TUtu7NkGYghM899aNX7wIy
fC5N093Bz23KH4wd4y/4tuILNMvObqA2YwwqEyZ+Z2QbEW9/ql4yQbxbKIkHJIh6
ynCInasET7k7ykzi889tE45u/nR1f9zniF/3elfrxWQw3kxgHRVGPZxl3fXP15wJ
qhVQpODi+cYvl/9kVyqSTfQBKyJ/CZ9LKrqgdDVXl4MK95oWi1NuvydoVPzgFrbY
WSGhaKxL/ulgvcIbnrbRh32dq/x+SsAmnmwwbU6IIZjQF8kSB1rlyYrVhyve/6+i
Ha+QJMC/zWxZUfl0m9aej1tXEpuMHo87hZpciVvJS7LcZu38OOcuiqpQuMyNlH8d
RDmUKWD/ituaEhTqGPjMjD1fkDg4WlnVgAWPMA3Iy8A3NAyRWWEadm+mPZstYuHb
YvCoPtiLKYGsCLCIzk/DnC0MPMucRGra+R99Zk7wB0t1xVrC4U16sSCjiJt7ej9F
bk6OTM2l8kInyRAtxUeCblW14fnkT/bcm/91nI3of0kgzd1GPvy/nw4q/hRst/aM
4H373pJLJ5JSHrVJAOsXarkkN5MnQ35UEI6Wk7vYzgYVLkx538FzxS1pbuzWBSY4
SDVnuUIr1Ofeloi6j4GKa6vXVFLKlF0jhQriEE2M3eVM8Q1Wb3TXM6RcBnVVEH4S
+6rKErpushiKMxWZ75e2dAVYItX7B3y7j3/O6T+Ue2cFP8VM3w8w0rzelgTBLG8r
G7SXakzAvdZdqgwOuoInvQxjGpPbFW1MZXb0d6oAVVQ8GtvyAftyjOkpeT4kJSMw
03OBggfy47tBHUPklGiIidCDLvboJDYNZ3Otpc6G/X2doliIeqbv68HgnBXPgHuB
LxbdjtxetBI9tFSJjDJ0RpEKj9dwVIORnFi0HzmgytbI6x964Q9UI1mZ7blRotdQ
gXRZnxm8pWnrXPcg0Z85w6SdfBc6IxKQiTEEodYKEVGnVhOe9SUTAMZEP5BrRhoG
6jR27NzTD2govlbeJphSgoYHWVxLGs3aCEEtbv87iulvrS6qBwBJUa7tCybspvaD
mJ13VUwtuRDRGmtf7vO+UlQAsCoDa2jtA8FNjngfB3L1ROS/JBDR4gHhhkWz7nhM
sQrj369OB3Y/HyTpLNya9MdxmIxKKmmG5YOsS8p8/LqRK6RA0m7VowU8aAH0r0de
LePIfe3DwysgtMapNQhOLYya6FVZ6V3lipOvjd3zFlhiS8IVbbkc2NLQVUHPPGdH
HrQCy2C8pLgdDtVQIeJ83FdX9Gozo/7nLtbctoDNrhNdDiQmcx0hGHrhStGnGaGE
G6i+Pp/x0/i1d9h30OO+GvBSGHerhMTb6GQDJDY7TGVLj6+CXukJ/w3HKihzQ5Z+
/VwGbW1TAHRMijhdqzCNjEE9S+T8hE+ed2XOppMHVYPKgKa62k5Bods2HNoxk6Iy
ww93a3I9VWBu8w1emIHn4fldGTsBwBg0xAHtN5qyA9JVYFM1rqpOE1/SjNDVAqfo
1DzbGO501azoUZbDH40GogNh9Z1DstcezLbC9VbYnZw4FYgesu/w+fLjuiG40EhQ
tsDtmsCnzOnhpxB3xiswNB6SkOt1yOGQjLlHVH4eSKnmojBfV1yqvjkYkXgutr5O
NhrcathTKm8YZkfdJ6jo+DNSb0X7PbiZzRQ2QvKK1tuc1FCzt60NpY2WSrZZxwJf
c+dLaRabw4MdVwQekEUoFVxBdCUbM3DqIGUK2IygNSXKgQZOA2NeO1itpxr0gBF+
/MkJspDewIhAf930x1EMqsDUhvNtrT41ipqNnf0sFz9rGWZT2thuq9OJXfLjmmnk
KAak7+m7ZXwSlopBvXOf9ywYBCxWdkjdN6j0WAkv1fXIwSUmGROnQp2wBTUKIoN1
K7pKZQv5PFW7qjYHrG2+UQ08iHXmJMDxiHrIFs8TGaW3fKL12fcOvxWfNn/8euDe
ssBP/1xfkpsFuaBHVf55Jc5yvbiJdRjwrcmlOObz9ZvI/4n2pBeZ0STtBsBsX11u
8eYwPoT4wzBxOHq+UUsIG+Wn2HBsAOF2sO8YZS6HX1g7fU0jtIiOr5leMpcS8Rwr
yhyFqWmjTpbLipaHsASDCSDbOSAkVefGACBEUB2UGLXgWgCZGGHdkw7+DXSxDX3q
aXdsiymS4pxrvrsAPGJGVaVs3F+xWPwI0WmoFTISJ5VUUresWJxdPsgrXKaL+vIN
EeNf5ysPZ3LeDs0HBp6yF+d4RhLhZ/OxJcvMj+K/PQ6Mx5wA9tyJDDImp7+hHMVv
pJ5HcQRY8YLkWZXaZau74AkGl/ln5NC1rJyA7saqukZEuKjrITt/nKDe3Twbh+Hm
k5zTQjUWpp1xOwwsCHY6n0F6G8VdRpZEYUDxfHZm3ZUX69zhEvRFW3Q2v6vcXo/6
yLV6Kio13jnxjbJ66ax22V+Twul3VvP1Pl5gLKQw7UwtxU9qp8a/u+mko0BEVrEG
hytFs0fwanWR/hPkaSax9LEXQDGRIVBJfwgRuRs0uPO1OnftVGH4zbsOs6XGR0WL
8jpU+c3iHJyfYfcpvF7h1M4vVFdvM78YIJNkdcN5MRfK4g4t4gDhg3c1b5b/GxtC
T2XC4Q5eF3r2kZaK8mf48Lhjb32nTvWIlK1o5Nz/fCzCOo0lHdVSDFwJ+PcnRdRK
F8Tb251cw5keYm3gxaoOQCdPm+lPcF1zKZBCLE+UdT2nR3UBkW8IWwWGQ4j9SiSe
tGR6icebNHQv8gMCtZ5kMs3WLbFwn4kflt8sXfuWAGg3Cx8zW/x9rz/s+cEp+5JS
5nSPVWBfIDzNmMk0rGLjZhkUoon3iQfWhz2YwUF1Que7QMhQRrMV7/ymnn5AQKQQ
+mRI2qkqy4IrEZGhO2WIsSpd/veU0kge0vWdrprRhI6ceOoLBcnwsB8DHUgU4c3O
ihJ9pAjLeQ33Waz1fuoeOpxHdUVFtzEJbXHa68SlGRBRNk0dIt8IYGVUDZFfSQL/
h4aLsxeHeMMjQhh5Y2JR7BxpQbLY3QnOfMTJTR03pv5VdXRQqsb1DS+cH+BYOgUa
f0Hpi1I61a1GyHjxH13y7kpnp5NGHHDULCMAMxEE5F3LS2+ws56n2JaBHqbFz1sY
drjtjEsP2tlv/RhBXJm3UKLI0p6cXc1Bt8zmedK+TbSvYLpTqg/udVNqlP39weDf
3wRZtotBhLrQAG+xv/PL6/OqD3uNuRsZjAq5iMxQhxvV5Ty+Bt963iT1MoJtWQyp
lN+Cs70fAS5Y8ph0XwQT2dh2+CzZ0M9vx9/LKT0REIk3vr1uZmzAitwBp5DtUcVP
pxjOmBzhT7ThklTENzAORtVwpZIVQ1KvgQpvCcL2SthrzI/g0ioP1VYXJlegy6Ey
3QdtFHV+l0eKr2wchqjcm1L9tq6vrF4tETBp1xJxkiTTfViA1383/9lJUs+SrNMD
DA++r4xFQWR647Q3FFT9fZBtniPrinF+EeBE+wSUte6g+dT4Ciyv5T/ywKcdpLvy
Muaxn8pkGU+3r6h853Up1Cxfzj6xZL/c+XrN4oBISaDBIa40BC7GnNrKnlWb2S2t
KISeEut5QGBBQCnYYVtwC40IVmCbYBY9Df7dJPbXiNFzzmwB4lzAudIY8u7sAiJx
MV3qU4o/T6bnFcAY5+yKLWdloQES/VPbGv82EIfmjYG0m52bZJJqHnJS1QBa3Kvt
B1xKC0Ya8RWpueOlewcDa8hqy54LHpzfoEUV1ZuHsHIZWVh5CD2DGzoCb7Fr97nv
jVLBwsyU7nLYDtqsT3zzJQ7/WoB8EMoqEOF+EMJOS8a3CrqZsQO1J1sikTf0SPeJ
m78Mr7UVumlC6vVizryQi0tk09KuJCXrDzPyI/amBqKtzCFswGn5iWDDhsjvw0yM
7oJ2eaDgQZZb8tTqYQnDkKz9L79OEVk0SPx7InmBgJ+XXlfvmfTSfpqVRxB6erPY
qpfV4Mk1RzbSM1rjAueuMCAWp9PqIQt9sGHDlIBeKWmRtDOntZg5piVAsx+doW8d
Fwfqp7cw3Wc3SBsQ+Dd8YnLjiMm1RMSI0J/+cj10RyqYBMKdQeLV1bZOEzh5yC66
R4I7oeBTY/5Ut9VX47d4ujndl5iDja6BykEBebtXKmmA9Fy3KFYiyGP6X11uyH9O
ugLjZzz6wrqFVFKosiryfkCxJ1gM2md1Qrh2CytWguHBrdae7G2+yt8rzXAinIHD
zm/k20JElhCWf/XdOa8O4t9D5eSii7rfH20B0Pp6byEbQmy/hMa3UB6IEA9D4eUJ
yWrZSVSu9rYYqW7BHk5IpOSa3Hup2LURgiJOmiPcgW7Coz/Kx5cqkz+diUtmj++W
j8Uhxa9kYU9A2wXATYyK4p2anPLwiedal9xd91NNbnhvX1wC43o+WWp5zPKW4x2f
vlezqDG3B00GSOQxr7ZFd98j9AsdpPoDjH2vcFRAwdC022sKvlRLUq4y6+ewPSva
M7L6BdJFIfm9QAv9COtSrSEKK4Mt+aPGSnHX46tjttxYz8dgJ93X0BfBY952ztPt
R3lU1c/dLFJpRMaUDYGs6GT08z5lN+bDRwV9UCcXZtkqSccyVZ+Dphg8Yb0TgemL
Ez/c+2hIAgrB3nHVoHqtMdQ4DouTZJTxr4hZ1buIoMRv6+b7mXe1Bwa8cJUnIyCf
I5MVi3hir1V0dxX7/gpNE4Mk9OD8xCvzY2dZGK8l4DFKuyjA5JQmwnDBIl1hvbXu
Th+BK55LCx2Xf29yv7PfOJJap4CcKWRc4L5hqRJnKbLUTJSRvrcAvvetx8fx0qMG
QB9k5TT5xBze35autfP7FDs2JRt6awD0nZ/iYoprWPIzIWOeTfV3WHgsSd5K9DrJ
W5CQ1mJLtKWNI8OaG0A3lZZWXu7q4Jy91cDfTUqDXqoY0589AAmxjee1cfXtHjMV
EGYfLGeogMenHXMbYbeMZGSdER1FQduz6K27NApVpDFUesylb5I6wrUWaKTombaS
Or7YU0rfwpv+I4uSG96hndQUfZKQqCT51acotlLDfcCBlLy6cm8h+1mAlqI1/5mk
ggVbWgZfmifWiK2GO2Y9vuG+3e5OgQM2CfCnwyyZnvwc8nLEPTiID2hx5Bpy82CF
HRdKwXn7Rto/EJEkzvKGqYlcvJJLmO2bcPl9YtmWNhXLdkAL+zkiHuoMDkdGeFlS
leGXBDkfn1/8A/yobIrDG5pB6mSXj2iJ3aBzZYls4M0Y89WQAfRSXJYMB9WFk1H6
IAgDOqoAa7uRDcFEgt9+pda5TKbqw6lkVMBPBhwO8gVJz0TYsB4SkflGzQh2z2Jj
hI0vQwoWOTtLNdbqcHt1JmeqIQn1L3OnlrzQSfCl7RrQcYKw0NgfMavjJJhGNzKf
T6bEcYOoQxmKXLRWRE8OqfiEHeUZGZKlgSUT+owjCN1TOS3u+KMyr2FilJzEO6va
iu1YWBaU7ALtILuTUysHaNvSfcR3gF6TNcq/Ns1nLKhKaCRUMhBOZkp5yUlnyvVE
/ItRb/yMbGC0Yu892frewDzJGW0DdtqHh4B+1oXT28xfgblGZh/1GVVH2OqqMgHq
jVi6mD+YjumPfuhy6V+z+S8i0/zhr1FDdOUYF2uXFSPFOUEZPIEXeNFfPUYpJ44w
v4CFy4OiqChwM5nJI7ngW5Ezi6AmzMG1FIBShSKqI/Y+Hrqqhu9tHb+khKg91nJ1
en95FUPgds2EThPhCgoYtX7/rET4WDUdj5oossOrSqz6b8nUDnKebVXvyhZnd19t
Qm0uz7ohHtPj+2Hmk5w2aEN+mS2tqgYWTEEYdrrT7ShiPgN0Z5G+fxI0rhLycIOE
mjizhV+/VMA7zyKVpeFirov7NO5EmalbzlYWEnfgioglHqFJMAdOjdK61mlMSA7c
+4DLt4cTmHH7dTVvMmFWNjZlust+twkWf5BLJhnW48xkEfkyilI2i4/aS5kJpmeC
NNigYqDndL813CTB42rmWKNxBm9JP9tg828LiZk8gHrEx+/jxJsxfMHdRkS3+GtC
TP6WivkD9lVAjphkII5NtDqrAfSTX9Fei94WF8qpjzjnfEUGrGYKm2tplDdVCgzH
xjtFyLr17ClDowjPaVcpCc3vPIoSj3o7XDW7nHBp5KSqG4NIDfI46R2ksfwmdrUS
mWx4zuerSUATfnlzYY1zcll1cox//KpWsmF9g4Ada8t1bU0LD00PGXhxHeKU8+0y
X8HlM24pGEfvDY7RqUThd1rDXkQMF44q2jmFLxvyFfRfuyxRf2wA6HwME/JKB4QO
nAvE332M5LdTKnUqxU8kgTOOhBYspJ+FQE8QgKBel2qiYfEPshXZi1QLUtu0Omsl
AVMTidp5bANzmWcl6r0TOoeOIKgzLUK5Vhg45pO8bVMGc3ugdiumfqFwC/K2QcuT
XdYA7aPETDz3z6DHAdvS/1KlEJ65ol96u0f1RKya+QcM6ZirHhc0hORsT9CXaST7
BfFoVcV+D7nmedk/0YG1T77/5vXGpx+LDB4nwiUgTgQM1wiBwWh5No1AraAfBac6
MaSi7t9RfkacZxgejFsxXQZRj1WWxV/YgNRHibEKnyA0VnDk18aYIab4PTy335iC
rifBJCGLADR4X29Ngskq1nwwL865azRj5g0aDOazyslXzvW2vGDrWudWFDJbQuhO
ZCpHcSBwxDyj3HxuFT5pbqDAvSZcE/BO2XQmnMH7+LmqN4Rbmrvy0jHtMB9GL22+
ZZkzsDjQVu6J2trhXWt1q3pcdlw0XN3Tt4Woc53e0JGKs4J6JMCkIXHU2gzirXM3
woHAbhskTQaaTlT3Xnh77JYfh198Oh+QW7qSGfmj3+AmU1zs9DgQsccWD5a/axKG
j4Jctgdh0aArt0uOSMOqP0iGkZ9zUSGVGlBDC+ta+lso/TX8GUozREPLciR9EjBk
yjt8TbCJnygZi7QliZBK156JjqqSB52L8gwf3E+77DN1Oyk2+Nk8RT3xuDKalxQY
ufmtYPUt73DjnDpKdY6x+UPkzxa55iaszXvXua7eRdNKjpML8UVejCK9Dpl2xKOr
EZJSfz/Evr3aXvWPT6E3bPquNeee8el0RNRFcBgB/uu/McrVUbFEr28V1Fs8VcyF
03nSQDoX9D3y7HcHWM1HUtEiWBC31Ppf6KYIFMPxBoW3NLdp0hw67hFC2R9sOa/Y
5Auwnb2EVGYp/w//kUqrzxJdnqXjuUwabtkY9SRsSQ5qqzLmsS7SZwG2aLqGWvFk
0/eCuuKdzbRA/BLQyW5yMkiX8InqBpbkKN9Y2WwXG/rGSVfwM8S3ZQD/N/M2notE
4jtPITg99rJkmfZ/YELStiXigAUt0ERad6MCboLrEietipNYmq7fSK5kkxOK2U6C
J0dHSF573N1/fXYi8aGYPwDA+ESgNxfwT1zVMkI1VaQlEruIf4jHhcP5XgrmcGZM
hoQj8Zk47KIvH/9MqzPW1VO/p9sHn0nI7D4GtoEGsyhRRPPGJM6FMfd5lSlDMTsk
XJ7xNVoCAwICqQ0xbyC8KerCMMnLny9XWkI5AavSGgWtTbRtkCFXYJEkBBvEeGKv
f6v3n86TmlzvzCOt99vj/jiGJQpgcyfJX75j2/PFQjG70CbDMU4+b3wr+BMTLlte
h9j/lOzz/42EwWs3xxbCfRh9A2BgCEvb8yoJep+fL+zIYpmLt/qiGaLn/3sMcuxd
Za7gGKCE3Pp5NY/OK4/zU5sz22BuLd5ZfwgJHg0afGSVpnOyE0/AoVdywLXagKBs
4lojn+h+8/AGmeo2p7cACPHzd+EcESp92/0GtNW+N9yFIlf2TqozfSQuqx8/msCj
ce8rPftaHXwE3z3uZFrIHBJmtkaIbCKv4bUhY7Bgi0gFTiMl5BpJkjNCA88IUYir
gMwOEqfSFKas+Qs0pmBCmDlcVDjcmPSWK2zdrDgYVdi5j9xN/bPqYgr9xfz7dFWV
fJPNSwYI+pEyaabzKwYYLavArvL2UTlZsqrgWk/tpS7TcoiM0n3X66G79sCxeuRh
r3pzeV+YVqpy+/AbhIJE/JlIq6UyNBdSduiw1cAdHYi/6Dwq0Z1XfwW9lEoLcUQf
/7ZM8o62BOVPFJXS7J/2bVpYXewxKeYZt+7W3TJ2dg0H1x+W2lowKuo/mKZXF6qo
GcWsUzhmdlzpiuhe7OYo/cy6MGamg9S1OcAXQZ6WBApZuv85Fax2JKYbaXu/1MaN
N/qlgN5FearHHVOlWqSky1MRTfE7OMVOXXcktH6EJKLOcabMmo9eaRWzdIXFZxNn
NAK+KrplAMdkZzbcNM8W3mxRM5N+c5kbeN5uXgnBKTBVnrkfZB7sRpP67WqBJ0h7
Gz/opoCC2s0vhW1LAWl+ly5dQrhdWII5GMgGoATUTnBVYFEFIHh7EghGAcJ14n8t
zIRenayJaKLVkNTpj53l+QUa7q7DKzCk9J+tmtrt25bbTl9l5ZIVZMQbqJWcl5cz
yUIEGvU2Y3jTN+QMPQOKSPS1NfvSqWeIjEHjE2KWGShVL9HZ8eKHFGsZQPTVE/b/
yc5WE0qXEzCeI0gPz/w5SSuV/NIRhSiUUzRVtv//+SI2FQXlpbc5uBtBiWLRTZe5
CoIVMqtMv3yQ1b4GD1Io1Q5pIU1yquBgdPTMI/jEBS2xO9zfAAkAjJZIsB8rEhj9
jnop9P6/J3weVXNmm0z3l81F+PLGt+JAA1rBmjMpqK2TgzBg5w6hxDFsj/zLfhE0
7z4bfyY46megncHy/fr1tQ1fP+7UI0DN7DNb2SHIOTUyRnH6YBw8Oifl1zmpykL5
axznEtx3ejUvxDw10dB2aUv7gTNsrYY4fiGXZLkNG9SN4f/kqDsnzhah/2DeIu5h
4dEXdV2uANZBSbjt6mxBmkRm6h+1E1V1fxf9ac+4VdH1tEhHRBljBr1B677va4CH
oc7d84vMfWiruFXFsrJJ3LHSaO2pges006ZM1Bv2j2ozaIFMIvNjYxtbepbIcBsh
xZnEs02HDJqZ1bvA0fumrNDfU7lvebT7RD031VPWQR5vE8kWini6DulBesJxueMn
ZZNYWB+IsGxKRvbwYAINCtixnCTmGtQ+LMtr+Wt3CPVyslJzmNbgobYAwa5mygly
iJ+bd9JK+seOF4lb+kWRPNeXfTbJbaOVOGGYvWu8wFwe5r3dp3TjBA+Ut1yumqjN
hijJW04JGdLijrYKFWaMvrgoZHcntHu6XV2CUcOIIplUC9GdcM65mGbezDQLDG+j
tmeq98t1CSjwRWOS6rauDy0EF5ktaIqlHgAhzCikt2affYJF0oi4qimt7zVzK56r
6/8qarKOBhCEcd013BEc7NghSYmC0EbjWP4iNrNsb1nAx1At+JD826Xbp97+bJPo
6+Kh35HQh2cfH61omphSzIg2d2yGVUkXCnq8jMxUsttFHAWl9H9PaCUraXxuwTZa
bWMtHtV+gIGnhZ1YpFGTIVfgcLuljPVYjviw+v41Brah28g1LFbJC3Y6U6b+diNJ
Vi7lsoxiEm6ThKnICqZhmrIKqZissVdiGNWxfaAa9xk/XZrohV2aEcIDDfkj80V2
87YjeZRrqegEfX6qJ47Hrjeo4/1zN6f559SoZyMdf0EGMFs0I7K42Iv1NxJ5lnCJ
9Ii9TnDvMs37cva1TTxE7m94W6NClJMOX4ANfPSga5NOIxubxR1gYMWmoT+mGN2A
wtISnslBRBJqFyPkjaFRx+loJGzyuNanRoCTNJv5hmjACuaXmZqGGYWCtf2KWTzk
xQxP+A1K1mQ9EXhkjYAFbsRkdcZiCUcwxzQXKjCoJs//jfxtnSugfvwZuw0w1V7v
O7xo2VyAlxDwJbWHVMIGf6WNYOnFG1M/b8KjBJnpipiNAvRFA7d8hLbtEDqFQMGC
4QJb6fTQtSuwWOUKUIiyeZ33IN4BxuLbJlv3ACh9lGksNJhZDQj/d0jzjlQ9DjBg
y5+UEHFBEBfa8x8Jjcuolsyml188lZTdykKcdp6fGUITEeqCfW9C4pwNKROfHwlG
7bFQ8SKwrDhJbmD+JLRpQjLZ6+ST/YcwnALaOC1PCEpN0FkFOMoVay3b7371Fx/y
aexrkaD5WTQYtZkAy4P8aCfgwbYIscbXC6r0UcVODIOh+9vPeu8/d4TU+ODRUDPu
+2zju6L6blnzfM879ATs0n7JdhtGghpfS2Eg9x0Vy+gI+cjGeG6rjOQatU0VWdSu
aZjhlzPMfy/w1CvMuftG16J6G+UG+4sPaF+Wy9/ea4ElhqYZQb9tZ13jRSJnUJqD
+BtRegDPjbCOTtTRJoyuwp/isBOGVnI8oieQ4oKXh4/RnY92Ed7b059XaIonlBNL
yDluGEbJxUoU6nTGZh3DTqyauB7UrZhhUladtUggJptDAgm42uxz+hX3GIYGrb6G
vPuiv7276e1qgpYqwn0PiT2rjlQUtpj+sF8/2dx6F7nEj7u8741o9pfcHsGr8UNq
D/NKVxqBaBmHZ24dIZBLJz9wcTmw77KP1dmG7uxUcw9S777ngQTKJqyLtJU3AYAx
ENGS1y4E5JwmB5whs0e0JAm52MpAB3yhdH+ITTHYWV6Fnrpi7tcUYuO1+xcneF8h
itpvuQIRK8Z2gv6zG1MgNQ/oGFPt7VYOdfksN/EVAzFH+z5t6Y0avHdj9+HNFafu
k0uGf/Dnci5DMrnJ+viVvOndHJujeMKctkcNNyUx04jeQWHBLCj23adh4uoOlQoL
UJ7XbHDZfjNzzUIAyf8CYgS8dd7/Xphi7iufNcIooejk2gGn9wSMUdrkqAQlNsFw
uSN22t63rSnzqvYCBSYKtb1AYOG2vr6+DcpUV621+IIDqhRii/ZwccZl2P8uHhD+
tVPXM53uj6MDY4HpMe9lpTcX+DvlFeqYsrIRrpmD8j5B/zu9xlepO6yDxgz0OGTC
pJWNpeTF48BtxUAat/qxISxasOeJWsk+HNkitpKkLG/ZbHP5Jmp+xT38uhUdUSNw
jUEVat+h16LDB4qppCUZqF2QPc2et0+J4+IKWyJ0oCkoZZ2ZKwDXMY7B67yBWcyl
bnFy0h1KPrfzKDeidBAvVpXWsJTRAvNhygv1llSYkFuii6ghoblfsjnvcYqGdQJN
hZiQSkUcnTRSuv/iinnd0AkzVmb6K9foumTv3BatDDmNdUblqruiFVad1AiXwQ8T
rXNup7MwWrtyWeolhluIEcMKkKwF3fepBAJAWnwcUM4VIyG/rj7d56NYzHQykJUv
cu3zxN85ssy+RdnSzKAIdlSObE/L/qBDOeuvvMENjcAas7S8FSno5gmWFwAOsmA5
qNpnObiDCJC9lcrjAj059xD6ZDME0gz+emBJMdg0E9O1K6O+jWAQbPTMQ6VI0S0J
mczdxKeTjBApPHQx7T2sv1G+1m0LWUxKL2AF0GDmHJnHkN7QORkbR77M90EuIkcU
bRSQd0gftOxbHhXEUSKgHjTFjmdd73DSmLpvWTsMCHf6jC4wvF5gl7FpSVHyAE2P
1KBthYpOlq0VHneDy13Xx45Jh365z7BxOEyLU6ixhwfYBeu7jXg21WjkpDdj5w+A
ZROGc4exrcILZukNylw1ppC/jEQ6h5hpgjuyvKGo8oXqUrxM1soQf5h3UEeFWeb/
mOxA03mZN4GqYlddmgDSN8ZmRL24bFKlJS6uXroBJYaFdXkQ1RLqcoj7HDLMUt5p
qTsuBfQZVLpj5BerfxFlcwD0Jg4KVfvlK6rpqag5Wcb8Sk7AgcjLmHktEI+s1HeL
XaKO0Iut59eMkea2d6F4b7c4hWVn1VQiAgV3nlL/BK3po4fWC7UtYAjU9CRhWpCz
0AvHyI2kdYpt/zBvl322+vJUJkNutB5+BEZ0pAFs8SM5RpgdqJv6gA5r6EFWor1W
foCORXNk0KataZEInGX0FQRdL+z8PrIIyK4m+c+/I1pBxKm0I4HN0/4VtonsmcRe
6w26m+4DFkeHU6wo9p2Z8gvUhMnhZpA8GwmNDrNLcyAuwF3iYVImxxaPtx9c8xSw
toXSkj0yeukC2BCW2aTEbuNCZ+FmaLxeNRUofnPtZHkqNBFjcv90nV1gyb/dlB1G
XG/Dwc3uRzvMBYV3gD9+flAmy6QqU2m1bXEaIzqfiP2pDxlVwHqHUszjojvRVNfk
b4XUF/MWWG3ultrAhr9+mIUwyo6m/+hOyk5z0wbVCnb+5OmAR2f0Ksokt0FjF3Mz
sfPB/q0uSE9wszWB/k0ZLyMkK/TsuX88wbc7etiVhw86ekbRjF2+2kaGdQriZ69H
6O5zw8/PsAc8OlOA4Ohj2r9UEX9IM6lf/5q/cs9bKZ5JGiXuikvI6sTZEw3i7PNf
EtLbyhQPLBvgCF+qVpu3AdPJnkSHMPnecf7vX5OtyjY3LIVP3B6UU6VoKaiRPiTR
HL0fxd/osI3VWmAnv8h+i+gzF2VU2UkEfEdfKPeczVSt3QTEh3b0rx1dIPVNd7rs
Qjiud2kDDB1K+Er52/S2UQMdOOQUvgH1fRd/mCXKA8FoX/k+oIaZfnZ0YTHNNzG4
/S1e7DbtC8udBNionyqFtQhcEHgKgoZwBM8HUzVkHMdTXFVABqUVQ1wd8Xf5NpLo
Iq1Ra1xK0rH6i1dP6iMrRExBwo8jajzQGTPXytUqstSF2xZZ87hTQbIDjppltPYQ
2q+fs0EYPYE/d/IqkRbtMaMoEnbElvYpndYxhp5PtbFnBM4EH/QkQnulFn1fZmpg
cbLu+zqhd58F9hbWMfvA6pmJHPecoxQwh+qoB15kq8f8ZU6bCshm4+li0yLNy3fZ
iUzDQhxi0gNIjmz8sOaVHYRrnoLVn2pfLNGU9EJTdSyttXsdJ6Xtc73T7drQ+PIc
hefGCcB06FkXN0EcEWN3jYrAUTYc297BknqwrAvjooOGZIDtEdOurWSZOYngA4Fv
civ7zEDr9ZPuILWNG3Ev0Up10r4ZzolXVVBceuXBLkUcofooz7ruBF7bC/lnmQuk
subz7EGTlhL1p36Qw1BiHj74DK4vy/sJlx0CGyy3sjvqyFqsFB0jZyaCQqfiHPj5
1aB6bW9/ofyah0HaYVnWCTAl6LnpOUaL+Jw1CbbqzQPmdHRWooefRj01Kv2F+ivc
9p49J2nrptOTpxpoATkfrnNkpz966iAoz9wiaqBr6T3yEEgOeob3Lhrd2c6XPXdy
3aFDBF5JLJh96ydfLjhqBsPEHUnj2XpxKVerPRQ5mrpgK7MNqmFwwK8Z/1PwBIu3
usxGcfgxES9UEgWorxWeOq/cpYlvbV4FP9hYTHS72eJnIGUP3EFaIxpwWDqcKWxN
6VrPDVWxiKzZ08A8RiH49BNZ1m+QBYacdYj7GazqLpdQDF4e5Azh41Aj4Pl2os2/
6J3megGme7PkiOnfmEYKYM7QhnUE7Ww3EC95iVPx2khyhififSUJOfDzbae0Bfmk
jKKyg16uSyfVSE8AN1LaJVZ00WTPhs/3UCPCS9bx9FDxKpeNrp5/D8pfwdiroWUp
2Wz9uCmHtfLaN00SypMW6CWLt6h+StR7fDmNWpXUqoYLrGIeG8ydVmDH2vF4u0x9
cDXd0e9nobvPoXoj881QkYYdbqHRGxH7twfSNzR/lI7LVXE14kDrbXi9OMben7W6
g+AhShFwsKrg07/8GJUlDvuqQcAp+Tip+SCy6vmU59a+U7d8bOKwGIkpYFqjWB+h
tvOWaD5IkfxgWmyM6NRWFcSbuoMgvJqVYHAiGnwzeKQ/4kgkO5DDTt71EIZi8lKo
IJ+Io7CQBAUmVGD1uaoIXKh9XpI6AZWR1e5AWF51qkxsFVgvi2vj1D2/dIf45I0J
pHp2Q0dC7wxSMyioWPYkkBYnq6UCiQrS2lXQfeiFzLST6wnCrBbdW5sKFCm0rTRn
sAejtkioJxwHdHYMkiNl60SOA7jDwtEqyoLwOx7heHdT0/h2pQE7meII7jO4inD9
8tJudGJau6XaxiZecorixeivMOhvl0FQ1O9c2/ZVUvFVWXTZyT9LBjjLC5Ujxemz
Njb+21BO8xwPBoiXGlQFqkAVzfAh8sbpJw7jAHpJam6I+G4HC/WrEga+65itsVwR
gZUvDz5QIdnY9sdwUQ/ScD19AdVh2C1oW/pm5a/pRFUT253f47uqeq5TIUv2DP0x
IiQZnlraPIgzAUCthWZK6YwX/5ky/y0ABHZ8Ggeai/mwfUezq5bnd0j0WKHyiMMN
q4xRDoR2Pjy7bqoOokVTYlr+oLpHEgBFETuHUntG1SRopKhjD+SvFjNT3Knr5s16
ksq4BveklwoBiC/YBPD5m+gVWcg2MUZvWp8XmO6FK0MPZSXxTAPfPiM38Rs6xevP
dbqbHuDxXkG/q8hxlYeCAgznwE+GpMrQP+dyVlBS8d81ktk6sDHg4qtQBDvGOrp0
exx9TrSKx8+/dcFxza0ke4sgWlesMDD/gkMdBZNiYKSuHHfANwldqqxNrIA+TfXd
gjOjjXRnVQDHnSvk88uuPsMJSyde2x5Hg+DHbnCW9hDvJ99XhvACoOMNBq/jQ9zt
8WqK0r6imnMCHOaDeOMJT/Ag592MUlKH2Rdmj+UgD4k2vmlEVzf7dV6fgbWlRadt
zO19DbXSWiwbYvQwvPdac+R0A4Pm5yl7zU5FzAzGzvc9v0MNtknis6RGShyZrfGz
nqRwOgnqGL9B4asXzSDKzSDrtt3XjF2qWLA1wJnPhbi0kaFwcB1s7LWD5xSQdoQc
lxvdaP3VHYPaTYWWJnbCmCLTxgkp3N3Kvu+Fc4zk5mu1MWDqOT3/NKURLGE4u7WR
ugsVQS5HqO25J2bk7hMoYx7/kT+TVa5XbbwPwYrF9lqw0X0Jp67BADvRd0w/ibNV
+AElLiaBbUfehaU3h6xME+gFdrIbQbwJ2LzlSopZPqx9p/FOcY0jrdslhU829+Ba
mH8bJ7dUvpoXSmavt6nklQ8GVzqu95+paOHhEPCwZp6vvRtVZcP04F8+zWBznUq7
38OXRN1zqvDGxnNxbUlIg9gwYNcN8ctHX+c4ZMNMNAxkaSXa4Ss+UCi3tPoluUko
QtQFsjeBVCc09SxpyKhsZTdu1qeLdz8VGZEBsjoVprpeabIerwderQT6YEi8IaJo
bdF9iOoz3E0RsebE6oQZQEXXo9PiHkmISmMgyA0ZsipUujhQvWq6ecTjfznjxmaL
xJ8YcoJXFf4jqaj2+wdSD6UGTXDxNC0uV5w3+gs4U9pcH6RphMMs4RVXtCVIUFHz
XZDwB1mhex0/Ffq3C4NMgokvbxkG0+UXKxCD8D6AfTbSor0jg3QA9GcMEx3kzqQU
mztIegXR7WUhh1VylYN9wfGbJGhFQuSOSer2Gbj2b8tymNvdRFnhm6k4AUujxo/C
yHi+slfDxZGAcI6nhT+ajW5jYf47Ot/bGV+R2iKHpMPnK5y65O/cFTj2Q2hJozub
l3gWdudHc07zhAaLxgFNhzTBDGJKDp4ycXrRWa93UNB93Mo6Hy6V5kbYoJsuGiad
31yIfSih9Stn66hQq2rkR1ZrW5AxMciN74tNRi7E+aw/0MWGAKqEPztQtqwOaz7c
xVGB9uoM97r8srbcuJT8r8b1Il+NMFlqa40d4dfiBnkbHT6LYh0oHv+16q5TgmOs
OxtkrLNGlUjtM7CSyqK5fZ64hQiN05MCs75GCqXzOB4avy88POFO53s0R/d1De8U
qotOEzhUFdnV8EDIPsPyAehZBYnH+0Z6Z0PDU2P1EvU8VtxSZEfLFP9NQQfG6UJD
fYdsamZutGHsr0kg5XnKuLZeRr8TrIGKNgwc/w3/7pi/ad2eTf23GnywNTHcobNH
HhkowKjoZFHpoJchN0vtlYRj2ZDjYPBs50FmNdcylqZ8YG8sPODAQwLPlyZzwnA5
yaCWeQVYp/AujIaRkf3UlZYQqFTbZ2Td6vsz84Jgqp2LoEQuo4K1Hm+4QJMNCD7I
myZPGY1y8HBQHIrUTP8HtrIu9nCgQ+oOMVi56tsyfXS1UZ2rbGyHq5gkIerHgIgd
NvmObZaZz364bLh6nz+JQBiTnTwhYc6vjh1i/wUqf5bQ2+Pq8SsAU5FoeFxbuTOV
gY0JQbO4qK4ZnFW7FHypvbPGPhbKn7HXBVY5F0xGDnwhfNFmBBpbFwBCc9WFK4R3
alhkPgeVFCBMGdAChN2cKq/qn3oXoQKQ9w2krlY9mjogSVoY9F1FbvIu44+KQygj
7HUsL+5ubiHZJxhk6jHaST4rglLtVpHsW/SbXCI4PB/ONUgABKTTQFozUM4i8xu2
zMVtSsy0gBLWLiNFj+lzuKlPiCY4dIXnnmPuJRKNyQFQQ5ksE6WhTmkNLdgPH8Mr
EdSYENU9wAh8AEYc8m2B5JVofXt65swX6lPkhI9ukuJB5fyYXL8zxOYTD918+euF
k7Z+O/M4mlQPOZKY5O50KZ9cmbzC+szY6E1w36LxdIfmu51A+2qoLv0XJYRLjQEv
Q+9ClCxfHNAZaaklD14iW5DJT8CbgV57DjkrAaPtQpgx25QVv0mxDdWyzchKQBcq
yy8fT9YYzhDrUdEYJNvxW1OIFFLLjIK3sYrSZjE9uLsFaxcDVz+ez1pCZcrW5wc+
HK6w6iLoedTBOb7D78Of38KmyS/GLFaPQGq6UGTghFEucGjYLs0m7UEGSZWkc2A6
2YnFNiVi/ZfFAsO8kUxOYAE4T0EGFZBwR4noIoTlid35VS7oABE84rK7qbWwxulL
ptOxKINyHPFArfsXes2ueZ5w0mMhk+4ZYKX3VFKFgDkoYABmlXGRm0yuhuuKlVRl
8tRnYlbAz78df8290niIFRx07TyUaHVzcgXOkavFUqMzIecD4D1ZQro+/H4voqqN
F9SOlmiPoxN2vQrrrc1EJ8fJTEfrwVFcSi6DtGv0es+gBp05isB4uhJb8PtzlXwQ
JEhal470Gpb730Vgu6X6UzxybjZI/i8d7QFLM76mBlWgFcR4snnpbEsvAu7TCpC9
0gLWk77Ps3fc14Z9HidZ21nig9g6MBTzNPjrBrj+1pFWeSx7tXLwLxJRE16VGub3
TMHziK63iSieZjqfiE1dV6RWcsQCbLdX9ezgVcaLg95sLlc3VVhm5fhU2/2d5KMJ
TnmTUa8q5n1DOlabNCG9Ybx2Agohbc8BeYO47e7x+hoSBPi8YGLLADnGZAWrKsVH
vrsBFhIFcYBQC+lSGpjko5/VE8US/5d5vD/Do9+n/W96m60mmtMmzKqU2DcfGJAC
+G++j/UwuXxtRtisNzfrDVfW6i0AUgnuupyy3Xg9pt4bjAd6xBFcWzhbOp7Q+GCe
EW9rZeap4mlWIfyVsaGwidomfF8kxUvmpgBtTO/czjfD17VvmMBp/2Z5R3upEy/P
Oqpt7UnGe/q7oRHjg+DRu5syRWywdLmUK6xgPbScM1ye6ZTO6+bqvlj4oJYk/pgl
dxKsLuU8cDLazapVzV4IT4PF8cJbJi6/WYn3pICrEE0nW1jwFrSYzP+IFhfANScg
AnO7NgMuVdGbU51hTCVJoqwv8/B2npcq+ayFnxyMH71oItEKyFxIx2+/OjnZ5iaW
g9KoRd6GLbBCje0Xkw50P1rKPcKllBa7naiU73x9rIzNc0mslmG4DkI+RW+wCZVH
nyG/mIFPQYaPAb2fRqBWQsvWOD9BuBN6mvEY+Np3dso5BhmLd3Wh/otuP8n4If+I
IjxfEKpbeqg4O7wpe+qaZyGvhsgXF+i5z8zhLzS/IhGYXi2uYwhnmcT/9gCFohtb
OoxofW/t3uOum5etqu9csFQN71itKlXrThJc8qnNC7yVgF6GLpUIurPlY7d5S2H0
rfK+QehGJSLzoFeZpRns52pIgVgdWPSQGjHxEz4zP5NgF8drLzrHv+6cdUOFBRRE
73RHwZ5FKb4f7T9sBMVKwf92dTwK2b7Juza/YorUp1Kug3yLjnEA5q/P8Z/xtOYB
GKppXP/aH755X+hVj1aErpl0FgHdBgaUN+HVoR/i30QITi1l4BfSV37PenfJH7kY
8J0CMuKyurQex9fVR18sBoMynkLap2Dw3jebOgwInVyUEWJtqoxbf/VNdgB/3gHM
Q6mZk/9UE2OY2I0FXhZkGPKT69eruk7xGm+By3d4wxnfkVoPvB1ay8SPnkkzYju6
i1UERCqMFKjzS9z3ppWypNc75pVhylwiYbXtlCIPGdeMzwOtkWKF4w8jy9PM3Rgt
SkabDtyn/F2KLI1D3TOb6qed1kYznN54Q98pEZ4MbhxvZgT/TQ7xtRLzGQcWT9Cs
ZkFKtkX5ul3orDeJrACYrlcvmakm6x4nngrMxS1yzGvpeYiitTecpka21vhwFoq5
AS8BNtbnfC/To8Xo6fZx4uRgyUyNSa2v8zkdzZ2NFV+ogwJzNBB1c8oGe76gCnLe
y7HVw8i7c1WhMsZ+C5cV3fgKEEJRPWctd0ilgAjLuumwsY4uoMrHla4q/RLm4+Le
WxjKcZFmD7GONOei9VOv048Pv62j4smqbdlCqQuP697Z6AHRW7lmovHEK8ISZvPW
1gQlQMwXtLQ8/NTLhdVQ4sAvLhSqKXbzCZvRLt3aoLi4Yb5UJxTUNzOEotIrbIEe
cgv6x4yzf4o3MWSR3KMU++6jKgXVuxAI59XcFkuziZYhDpMYvvqhrZNlD6WHRgJM
CfgDkVpvs77ECWPDuFsZIXZo7z1ksLulLN+G4pug7qiXm8QSyNLJY8Ji4jQGDBy0
6K9BriE/UyM1ja8P2KZUiDAalD579h0MuGlY6dQ9kgW/dwHyhkPsV5pROD5zhrD9
iL8Q0I6kaE8IOXDM1lVaH3DwrYi9067A7il8Rwc8bsfvBJVTdGNxzR1pC/q9tLCO
5dcDqqATLdur/VLu3r13GkzzBqX3FDSgKqA32c7RCQzLJrM8eqoFo31ZDAgmQwba
uYMYKNdOBN1Pm0CJTela4fQgGGZ3DkM6/w84z/WbJm39nTl+oSsZSTm+HFhdfk0U
NchET6V5ojpvCgc6t40YqPg8391ykjP8ES0KY1EpI9SAz40N2hRnC4c8EehbDX7+
ieTpet/woQH8Voi5VSOOX8QF3aclbrnJ1OIHGOpa5ZOslDmJv+gbXhkiOefzSSre
xftMLAwF6lP8anpFR/BbNNUIpc4hdkbL/miHRUVUHRR47CKtdeQ1YuNXAHwC5Qai
W7EPVZSnAsv3pvi3AtnBR15jMec9AQEbK7awoGohyQLx60dahxiQSCgXk2hhX8HS
uW9Y9wm9r1Cd43BF9LFUf4A7FlnRlnfiDUmT8jYbvmahFXM6dy2O5qQY1WDBsjVM
xoWO44TNSOe5ahNuLk2YMpHIljwlbyx9IzlS4pAf3ucXVrOyp7vwKN4XVayQzmya
sq8gHW1b0nt0WJXXvIpVHDrDr0zpkFXDbI4ige+sVaan0xhPXGbFhCdr9Ri2KFyX
DAa6wZoz60RJE66k74FaaYxs2BvnOAFgT/K9HF4loZ2aBKdwxZlEBpkXh8rHYjMc
qwtasMh7CIKNM/WaBzqeaNM/T4Vs0QCyy7lVmBPIARIHdXLnyqywLCLVKSou3POy
ujjZcg2I8U7Dkisi1Wvhb2fsgP3D6JZdIydHayDDikmjztKJckHIs6MC/Cb+p3vs
qTxZ0q88b5mnD9DfxjKKtcW3US4iSFGA3BsqzZiAxFkKsdsWqRFN6fSo6f9wXWoU
fXrxRq9IfNwUgCg/hcGTtHs4KWJKZ0gMG8dfzlTxT64VPJXOwvW8nLzPdPYUdefO
VTi1AnV5vJ4e+apq/zQ5JbeL+Pyn2owEp7QJjG0bFFGMlBM4k3y8MjZRrO4DPiFV
4Si+iovHgAO8oL18PhuU6XYUCsZk7jJ/xmxv6O1/E2GoNH0QgAHvCw5Zsp0AqLX0
1U6x2LXd7RR7zBlj3lBhhhABEXCP6IKg/L3PcHF6ShcgDvaBGeBlOFHaaqmP57nM
H0ayiXmiVbXfSnA16jWm79J38N9lX1jATIbjTrjF/FhsMJKsg2xjEOfr8SZNuhON
vLDP4QDuaZzMkcCwLTnQ36LzJS5pr/N2WMfwHIxeeJMCDkGrI5WKHVzrntuuzVuA
F6Q3CmJCRM8SQX6BtyJvZmoLPWUdyRyeq+8EG2d/miAL82ssdOPa2HFRFVcS+BAS
8UUqUfhqLj6DPEkfiSLUpFEJMt2Ul9ScuYwdw/lfCBDSspAKRlPWvpFxvKVwltvN
uTamyoc0N26HyYYmz04QBxZpRqShPvgjHUxruRfHA++qOlt5AJSpJZeNDBbIwjz+
kyHZhmi6p7j9+0+vmjJreixy/h8iJLNQT+6YP0yAwRBBdeuucEB/u/oiPfhRjMti
Xd6pPecPwZJWd897JMfcoHDu4MbueOjM3ZvwCLNKviQNS7HIloMebkTt+DZT8tCz
hL27bu8Bpjg4/ctxdP1Xb3jYe5Afd9ttlF7aPEAs2wwCJPFHFteQwZq6Kc5gRhje
QPrFq//9mJrpSJeTBR0Y2L/zyPNB+UKprkieRVxa6rjy2mk49q6xs39swImE3Ntp
tRQBAehixcwmgz+e7fdHgld2ulXsObTx3azj+lLw0NEa/sq2VWywDLfjulx2VHRp
3HzHsu0vrI5U5eEQ6P3xWk0PCemDWxBf5KF7QtALg4dkfCUnATd9m3Fiqosffsab
ANNwfloICkjIQPIjelKsDNqhtOu3x8/kQKojPqlstLueebcYr0/P0K0xJBYeTVKB
chNZ7N8t0vEVjl/rdmNyanTIYh8hGAFJDormZTRV0HPFL4EJd7jTqXYuidcKQwxB
wjRhjlL9mi4cueD6+gonASOiwQsW6A4EKbnhuuQn55P12pALbqs/dY+JWIUqiYcA
3BfZm1nl7xCe5w/xo+/aBDRdEOv6zruw3epX7GEABX3ox9zT66S/DjZsls6fE73r
ieHBmBGTYVr1rxCDdNCoDgm5obb9K1S3HxGMIQTQZplrwgVsNLyuLYbA39YphJKg
18tNemPvl2NSrmW99rwxikTq70IpvCvCEs8vCh91IXamdV6W/4tUgH0CR252U2mp
A6krWX3ZZs7dzwZGT6zLSwjqTPTVIhjbQl1DIYe88aN8WBGuHtHuGW1dlsSdMUDS
9qqwROy9OkqVzzaCGRbso2s6N83SQeFrM/P9Ahmbg9mdpj3tCXOB9sWxEhxi8nKc
q3GKeW0PeoOGNYSwK0u2RY+eljtqhW8syI//uVrC2lkk7/UR1KmgwBlyhSv1F1rb
M1wl0uHsFj08S1BNBxOSeCA7a1nAxuO/J+4Lx0sio4ZDLhCnVO3zj5W1RZ5Vkarz
BscM7BeSdUq45GhYvm9aKCZwpUmnITWIBovD5Aas/SVujxAkvaU7fOIzbzeB4Ii8
nltBdFpQfyAgZcWbXwLvdFTPsbtVEHohGS5sJBtc5PKZeYXVplDtZ6LAUmFpqDUn
sW5rOX0NaPE8rL9+WCoF+fZyp3NHAMScxQ3FjqFu7KNm5qP+LZWyjZWSltNydd7N
APcTHAh/0MM7MCUuxg6dX3SC0AoTM/e3O4dhdAJzUTEYhF39UEzz92iikZqx8z6F
Ius9bU0Ye7mIqGwN/DYf094viItU0WF0MVfj+80Ghkyh/jSIA27DcZAFDwjHUXDh
OzzD6yCn/Y3CSIy/pPGvCkJJltYFTuTPazUuUn57A9dDkQtfLXjdlGk2Qir+90+d
LoZTKTvSorKimtjt6dWPHx837gycAXEiG2eXSK+iHx23Vv+Ikm0ef2psCine/ueK
AiigIs9rFvEjLzRTZ3iLOWJrl7qY6FAnz8e91Fjq7SWNfX9zmfGZbN16e+4XGwdB
WujpTwFqnqKgIkU3yjDk2KG84IuNl8oAKKNGYM92bTaLXAv5OhNNv0S9ypuS5910
oGgNYkFuqAEoxa4J/3ZYktNVwaAl6NdaBB+TFqupwoP9BK2ehLbojNPvPFNgEyn5
wWnDs8Y6sgsrZi53g+Yeb2eziHWGn98h3ciAHkRAwJqfsCUGcZeVmYNvqa4NuPUM
VfVRLLKzsn7B6h8ZFT0PdzdMW4LmJOFfrx2fGQkpQZkaCsNS78Fh8SLxM1qmS+Uh
pSEeR5zQZzxBXPZg6rFkEc+D+RI92nPpmQKAg8Ez+y1/9WJTK8yykLWDp68VrB0c
nG/YMQEkIk/UW4VtuJDP9paG0tXMK7U2jf/grifYGTOg8g/jQawJUh5HyCi+TwtX
bZXEa/jd55TdVtMjWD26KhMQtQD4Tb59rhPQqt0WVif8C8OiLjrN8Z1/8tMPPPsn
zQVRPZHfRFE2k/+11T/IUts0d+gTWtwNFXybrmDWT2YaJZQBQaddAeDB6CA2oLdd
hbooL6iya73LivGe6mVpkousknukUcYV9MGxujoNOgm8pKwZWMMtsjUiGCPkKunf
+eQJ7Wobr79wVN0wW3z3aI+AYRdapS72+ZVUgt1iCg8G0DirOxX0O4Xujl2nOkX+
HuNTkQd/KCO0I7Ex40SH6gVWIIR+bTBJN+m2IlDIY4709YqxCj10yxnadopcrRmI
YjbeRJ2uBHK4fpDrggrI+pjtnkt/4CjVqOaxYRTJrrnKZYsjncCvUz7+JstEwdbN
VCPRkvzvX4mL3nFN3UwT9LchNgcFucmFHUEJDU5uqgiH95U/H4ifyEPT1Qy+vz9k
/6YNtIhIJmcEYmTFS+gkG41zun4d3/DElYhPLMYTTTHrjJoOCTt+83Mr/TM/CFof
vdPLYFrc9mig5TaZl+IUDr5UNHzHrexpSTKi6y2ZPJRWFT60W652gPkufVxt8rxO
0RIcFC0tQawku7SRSk/p9w0q9Xn+710upR7IlbcMDN5ba0gPjszCqqB2U1LfBd1U
D2zBemqWmTAv5ePmo7DfN4vmZCdbtsedL9/x9Y2430q9MChG8SrHz5TxRK1GEzwG
fy4+sOpL8UqIOUEigBKrXGFAyjbqwiLwXm32iSghx3aVn3J79/tzPWxlAcwC8BmF
34qay66e8jLi/f26GDFQEuRj88OUdeRTrDaqXVmH55f2Ytww1BeMRwTYoy4oLOkJ
UHgfQ97mgH/dmsJ5/j4zVjANMTr5ab+SX/Mm/9PSlIc/XEIH9GMNP2uHCj1T9dNm
sgYsO/dqILdAV6mSDqRSmsNHUg5MHegfTk4KhZRDzmjvuOz8EiGDV+uJouUNovsY
7378p4ueGvz4d3EjgpiKC291qfZzp8riqk1G2/AjXytHzILyquxUmDgGFN8E0FOZ
ePoyeBtE2x3mcUhAjAt9Ax0PhpnyC35/Wc+Nyel0Sn0f45iO++zXhrslqiZvvT9H
8uNSyVrjlxvOjwhuvQb2K9Zn2gL+0qGGt+kbJi/LKleilUJOvkOkr4uPYtpAGgZ5
i0i2tYcm777F8/9zW/bQlSt2ULldvEhdwAw6Goz375B4Eqg92Yno0fRIGR5eAt8J
5FlW/cJgefmAFYtGRaNLAAfIWAFn+s4k4SY3C/keG3QRcf97tJaBuADoxP3sBAFX
l7OpmM43MaQrnqQ+KjOICY5YNUKUkIHhPSjucgCxOt0VwTx+vIxlP7HHH38emSbF
MmuGvMarXBzlYE4tx18pDlBerAk7bfsAN09o+4p6eF1cMBBPiHU/MljNy8hoDixg
UcM2h+HzBWLqYa1z9dW3ZlWBbRGCXCjeXFT+vsYvsEfLdsFGr2Wc8OMTijD6C3P1
wd8eyK8CsGoJ6HOeOQI9MDICKU7ZWAVWVoUMX2nTEyAxSoIkTAG4xeVAhpBtejMC
fdM1DZxjLq9qBzPQCoTCAgMqkl0gBlemBLinQhLVRFOpVH4Tm3iM1sMrOIXgJYSR
3CtLs8JxxnCvHO9bpOygJzw/a1/wMnUSYaqWsWbAekhaw+zNGPw/flujcu/Lcsf3
btXA9VYOXy79imn2PidYP20j0/vowUThHtB4xErwPdrhRQs4zmuHBE2bLH7Vahv9
95bn9FklnD9MMS0Jsf7qZnFZa9NhKLolN7ip9R+F1l9JXsWPhGM+cq5VEBBfTX/S
WJBhsNEsGEDjctTw5wb2FNWyHchSOPjAMf1bSbpCh0Pqiwny58Iii4/k56kXekBR
vWVCIFBZhZmM9Xc5an54iBs1vIdjNSX9jowerE5tSmJ7aUDLRmtUUiKtm+wb7k28
UfpvSx9RGqt990EOCeSvPXIaL3IyVV4PVKvsHGwhR4mnbex2TAQb1r/MSAF9H5Ka
IzxNkhhfm2Ry26w7g1BpWV6002YWiZVq80c0JuYqUMG5yjovtGOl9AcBt3HiTQjC
wxQujg2XwX0HX3f0i/7pgGzsXQ3QQeIgN7SBYMHU+zkCPzGuKBVqk+U7iIxCUdTR
gZDFNHWODgW1JQE4AQWD2GwK1OI7z72XAKfuBxyo56YXF4EXVR+048IY3CbvBVF7
7m9V5dkgmTB2a1T5Mlg+AjX32gVQSh0JKkMQtISG1QSZ4R5I577OwYwEw7za72T/
6zmi2tYQhnnu6yqdxv0MaKQ7ulKgSaPKUJdjgmi3AVw9aCYOaZBO85wjuqP4tyGG
R0uvxqyOYHwsQZOeilVpLfXN2hHu+liFnRuJYVoGlrhoBCC3QL0EMdHlIyd63Mqx
EhWJSHJ4jDSVK8uF6d2CQ/16zTFZ3ALsn1WS2EkKHoUX8bvJsNeyTUX/vBN1w6pQ
K2N780Q+kvBNSlLIjL2HiRUfvZQqoou5gACKkZYqmcuEuOooqtjuFlDHTO/ygauf
ihfLS/ufV+8L7T3FDda+GCdXJiROiejLSUaxy+my7FGBs8e2UFjM/r2pEQknAneh
/Y0gYUWcth7CuB7zaM5Oz0QdlwIJmp0FYiKu6K55NrPPgx9sLHwNKNH/ZgDs72Vo
1q0WRCZoG9afWaR6VbyQcfNW0vVu91yjOxNIGduO0DHBAGCihd3frLMn9L7oiO9s
UhmTd2MYHjvVVqMyII4PkVd1g2t6sqVmfdHlPatZcUijFUVMGCAFI/qLGl2WAVB8
L7ufdwEtdvfbH13kFB4ui+0g67r9G1R77DwxE6pq8hZSTuwcLIDcmexV5rgpepfz
vhYnYDl+n3GybUyJX68s96h6STb0nEwS9Wm2EE4f7x0+XYYJNxH29duw+wYg8K4C
HH6jzIBamwobni26z9s6pZUXWP1T6kfDlnSUig7bPh+f6xyrU88u989BsKtA1QDg
sm8W7iKvbOpo9ovG4CHCpP1E+dlDsG/ggfU23SAMjl9yyA0qRMPlPzStSZvNUjDQ
E6DByqJvQheqknVHrtdI5J4moOIluVom4eW0C52Or/L2sNexzlzvosAOy9b9c6FF
X38c03isvbfLbndhUBmawWJFnqfTbCKHIIeMtOjY7z38eoVpaQ6axqYuxf43CETP
FmoCKlZpWtR2ovhARqmhfu3kN0rcw+1JYdw2YENkzo1Yf16yZdjmUt63wXkEzu5V
YDoH7cSy0t2xxvOh1ZDXr8HjyOmYvKVNidS4pzZR6GDlSOWOLoDrHl+glO8jaeDE
sLzowRC8b5bLXg/4ULETXPKhNxz1bTmO7t+vJeYY/t8+8+lMIbWha/QSb4vm7sPC
AVda3z9Z8adUsIS4ea+dTBFkbxawLJUZBE+/rg+mNpRwQ/I5VnJbcDorHhgdUHiq
rABgXqBh1rZswTBWVwlJERDDVunEpzrrrI19qtWG5rlD14BmwOvTk+qN2Ww4N++L
tuwYF2BjzWR7f9RjKtB0YpYiIB3lffWNqcDkuKsLL2NoTJ3y1qQeJ6fza4X0gjuJ
ZfRIlKTfYl+ietbrX/jZOy4758+IjIOXrH8SIpO3Pk4cLUevV+UcHifjKnmX6L4w
8JGpPhxia7Pyt2lDDFwmnMyHcY00EIhMnxQuwzCdXU6gx5wAmOb/Cnc9WX9VqbX4
N1eKxcJz/Ylu+WfPiqQAuZv/h89gJNlwCTQ8Ad6rCFjzajn8tlhd3F72IFHwSdkq
wnGHwBQoN3xxv1RxXaB8wd8uyyYcb2h/teZqmRezYus+nFKQiSv8SLtYZQe9N2lq
IKM2dtZkGv1g086a7brzsvhnQU8Ril8sdFAWQmk3X2KxGF/UNKXcP3vrm5BWMrAp
xCpblDDgrAGvxHJG3ot8eDTt0prMECFVFonxItELGpLFXp/RjQ7zIt3MkEFfpkDf
EUdHGy8Qz0vcasPqpMaYob2Om+jMuOh6h5KRIfVfYSYYnO7NNFKp91xt+6MVlyqI
mHOHwet32zu6qub/7MT7zQ1DwucutE6rac6qp0BDSS1kkmtyUlp+EiwL+Rh6bryp
k06gw19nQ8ebvCMDjsiHUrX7GBWrdRr3ry3k7EyrewbUJecNiAr3ZNjBw1oC+hzu
U6A4xLi/r8qIW2azBl+LEtn3bDwL6Hi3+pMB1uQk2jMDS/+PXBKfLAnoafcHhPjG
RYWgBDSNcIp7z1kT9l3KB+BCqMUoLA/3z9JL6mOepctUZ+4WNcWuBCGB0fIs44CI
hPucDgGD49UE5SjZ1ACD4vWOTzHNF6CM4h35ShHtvNembo+oge26RdM5SewsbdVr
hhERjBIXaJZtYtwyIM9xhWFAPSrl6OIjUgWd3Y6WcGsic21T7JPQ8SaG7yxdN5ba
mPijowCZ8XPmF2SU+Cm3Vp79qNdBQHM9jPD2ksiVcuyONTOdpID/hGV9C9XoNMqG
oNguScMh4z+k0R3ltZj3btNCD/eGFG00BWKn4aFRo+TSKAalD0lRQUdA2p7fDDlR
orlM+gJ6nl1HyAM4xoBf31DprXTHJfZjJqBGJwZ3rKUUcmrrqgFgJKqJAtjuN9+7
7ajQ/n3nMd5Qz2qhLhdB9Yq5p49FZ+hlmC/mlu+BR3jpwF2QcqITZfW90GgEESGv
VZTJl6AGQH6bhqqN/KrzAANHyJITMjcKOWHPLnsc2b80bCo3hgphYY0o+7N5CJqK
J4ZJ4Y3ZdLrvymUhcGPsVgKEtJCIdMP3WranxvyYkKeT5TTz1b01njgfHnliaO1V
+EfOzmC+DXgXrdCXbNzkT90voAQQ09nBEgW51Fard36OzN+86qv2ISz9G+uDJK5v
QSi64Dz2z4jTknFjzeUFiMrUW6n2/LWXNFJwj0L7LBclcirKzDULwEgKsZwVb3Cq
ZaT4ujMqRoOqQgoMarFDw/YcdJ8MBibJcdv8oy85u8Fu9+jlD+za5kNyDYX06tTc
CZwcI2RHUHrBR1jm0XSOAF9ZiR6uCny+BXTSnSJ1ofrNReq7bU5rASmR65KKUYUV
8TnRXQdgQg//P7QdGpMSxg+VW7hjQWMwADSBmreWjojv/khqle7eIpoXmB2Y8a63
pBtyqdJJ/nin3fylsjniTy6MHt4a45uhAY8/kfulhl+yq94G/jZgFv3xxpYkMpVZ
Z2rT1+DRxU3YRpwqnsyQSMB7IHjI3uYj69gsq9tdDZ7S8FmeCQ0ebhDb7jMB0hWp
ivT6u+E2IBXV/yG9p/T8d/T4urD+NOStNeOogvvMx0wjADF59+3pq75aXwc8AKLL
sRyjHNPz17HQCMWscbnd/0HoYLEJ+H/E2EOiXbboOb4FWRCShYdZDlHUlWDrsz3h
SpNe43g4wCOOzY6gGJ893k9Jhvz7Ow1fIa041bRir/1YG+hxvz8K40fPrD0e4wtQ
Q/xQExvwOpnnBXYeXC0uKzkj4kQkIkaEiLtcAHF0Kd6M4aFtZt5n8hmPUFXSl5R6
CFnI9ifwfqVVijQ/f2H1LKZNS8YYAvK+M4+8urgt0p+RYviWrWLcUtFw3+cLWaSP
Mv8davYr01SFubXAZhWgDyExana80wAF3MopZW5crukFG5UeW8NHMpPp104vSqHy
pZjAgJN5VcUFVpkY1agvlm6t9HuLtAe48t/HohP63+3nFzjOGM55u71D16Owc1dm
0di+bVbL/LHxKs/buZSoZix4ELsJwbkJwhD+1YQzVl401ifEzHh3ofKaD7scIcyn
APvVpk2uQAi2pE36pr3xzffUbnCggYY/eGPQ3NI+LNVduRNJeivO5l/nlcV6thMY
rEAGSfUozivvtMJUWIgI03lFNAtWKDRAtzA5RkwYEIGiBC0TdsVjefeZbkJg4YFL
CEE/RPp5++eFmzKb3prPVQPXPqN3KQzpFlPvRgNIDKMP4e2YJKxAej8S6ngysXWV
Kn3/tToVrHeImBkkdyv7vVCxRS1XxY58uzS7Ztkuyj1qLbbd94Z3JewkXc7g/2CE
3bkEXGaqkC0BgpuxBc5xzw19EoprJuEOiNhL7r2rYyZ/bm2s0OlAOPfyjiJ1Qdd9
odyn4K9U/bgw3iP688ouwcSbaw/DTCzwn1ZSB6beFTzhZo6Wunt9H3ZKfPWc4lxc
eFoaHs1kTG/EapnFyAKY2ZN2arP+5HEHn+v6vk8Z+rFYSioTkWb7D7/6l5CMYVjo
P3o+JwcK1FFhUrXG+iAattCCcLz3vIDvAwCVDYGWVCRalhpusc/dB69et3K73JL3
EsU7xycSgnt6sQ7xiJix+1f6tQOWWgBZbGLWgKU8Fu4sz95ZqN9fwMAcRN13Ymmu
RoScGoFwKNPRykrubaJf+KtBRABfaKY7CVrtI5KTXuE6kOhKLl7nnIilCWWoK8tg
EbhMq6V+NRcaxcH/mQYr81setyGLh2btK25MVhWwiFGFUAgekuhqoDy91CNV9QaG
6aw6t+68iypIIY79HshwNbkE8j8uV1SNsZ2yqbvQ9RHcs2qtONzPC9gZ64zhveb3
Yz+lmF4OxYsRMkhQ/V+vWSbYpA0/1Z32cYq2ISdL0Ox+KNrOR9t6JKpB6o9Yo6jx
2IklB3SXDHplp4BX1owuwW0wHYoAfitIIRx2kKk5m4iyjyM3AdxfIGP92R82+FQQ
b9ERmvW4lrx6PBhWIwMN+JNVrhrfq6zdvDv79Cb4fPoxnXQQyl03yKoR+h51BvHv
LZCeyBNh+fDfFTd/Smdlb81d06Z8CnvmyR1mftdMgYuR4amvNMZUNvWSUTx+77Dl
YRc9lFD2ERQWzJdn5HcSz1EdLLCdiYYC2468HAuQ7VoDzyNxTwgOZ8m07hpTawO2
LGXsO5RUjCUnqOLKwj0j6WfADv8O+2fU+JDF39nAYJxT3JVa8Sdg9kRMnvGsN5bS
kU5ClvsSgmhRo4JlAUxoSTmkqFDrHQxP8N/9H6Z7jf/2Fx+2rzCR834W1z/Rum9G
/7SDLafc9qaZD1ZY0edqqnasH1M57dpCpHf4nNpBf6C1q0wsF5lF8kujgT50dzRT
4GRtkF/ErNlPCC0mfojisaOXW8vqrkuxNGYMTWGOq2cXcqX1wXfe+7rAD+v9UbGe
MZVVEfk9IdwsGYIN0ly3E54wOIcwLDE7j4dxsJlpkLf/wpTsMOqmKg0C5Qqk9oTq
fg5qZ/ZDfshdjP3bjAUCiNIiv2zFlctMTvoSi3o5wc4wxhFFD+nxK2HdTW3MEtgp
XqpWVu4CM1QYgmaaMaXkutc9h3EnQ+V+w/A0ctaWOFeyzjy+r8LMkLSyvR4sdMNa
OzUDxzpvsYYppwkMCFuVEVwehMYbSxihnLvIQj6qS17tnlp8Z9bpl0KjDOwHrhMo
9nKDZzhWUCO6VJVL6FUyabDtgw1JHLr1ZSmOqQpIlFYjdzGcb/jvTNTmipaX5II3
U0DE7Ad7HfNZdedlHSjHMV/zezGHXIbMAiEpNOEZyinooUxMDZhDCaCCbvC4PYBv
0znRk59wKek3cz6Di0gT6utcOmU53XmyCIKWelBAxHZCyoVPBv8yTx+q82F4ZZPP
kPF2nqShbfKGQ7nMLsy2yl+4SmyFlbBW5Bhp0dIZ+B82y54eNWtlApuPoGZtCg2N
NI8EnnU2SgZ97uut/RZz92WlbiAI4B/LltjG6bWMFzLaFT6v5RyLHfEYmLURHorO
EpurIA/da+c8EJIHEIansvYDT0+Stszd2pkvEZu8iDqByX5H3E0zPZ9oBBeHHJZ+
MnHisDZ5sRwIOLEnJAO+DWmzrPhWACffxlybJIc+eWKlOxi/RuKD3cxRPWVSDGeD
//dqX2OqsC2/E/tKlfbUfKatNaz1sdjhisN6qGwqu3PIAO4HhxHWuExdMTpnB9my
/1S/8Z2Nr0mB+MKBqmBLC8wLa5XCyoweoVHg44XYdGSS+uW+aVVap8+U5yrIj6F3
hAjkTwB8dQ1AOcq9njDa32rh5ZAKZl0Dbr2DfBtsx9kj9JKyNAg+6eNgWwwxvm27
KZWAt2I1VQb6Pw2XfR1/sWjlSan2hrIUnGt6Gyr8+ew6GBK4c16ewdf6ygRDiLBf
VagGlBW5zmXY/dlaLLLZpZEu7t5U5T+2bc+2Pa81Dyz7Yg1FS+CvHj/e64glRazU
SQljrR0z9mC7YauBCxoSr9RpQmOOqxMEo6bcjXpKcDp9Am8oaOeqFlCyGR0UIqaX
r2/G/4ob7vJb85se3wZtarI4UkCyw+ubVoq3FwLs51CiCYcOJuGmFRoEVxCEh2v2
UH3Ce5sLzVZBIZywh1E3nT1IiM5vThrAgIwksx3aa4r4fJp6NiCHhzPTpS5DNIUr
FFX5tFrHx8DuNRb7Cl93ZoJ9NatLxU4F8VMm+Ns40iqbJX1I4S2KAhHiHzWTyxKK
8SExnIBXNDISQQ5/jHoellLizEVf5qGhxO8ScbLLuKIltpZoaq7R1V73kQ5Xg7IV
swPkRfJU40AluczhD9OMLiiK52KSOH43VqiBQux1BtrTfoASD0jCuM/PK9JNvdYZ
NeFO5a2JXosMoR2iF00wptcaXYikmzfnBVABm3mkRkAFNDLoEwssDzNjU8qXBuea
BEWJhtn+lbgNjIZJodCcV8GqyDtHvcr5aKq9XAll0kNgcCRp5QSNIajNccRwZR7w
VrHQjAA8rFrGdBGiPHHf/3jEZKv3N+TgFdsqhqDQNohAlBNgRAaHvfwuS8CqpNRZ
MKq6AbK8irk41H7T4Fv7LDRYZwn6pm+ytQm1Ggytelodxpbh7yMtpFq578o313+t
ewo3hPEPXOX5T0wjQkMmp4Ob4dbGmr+mWz+Oz1IdGgNNWKtySH1Av+YNQvaukjqw
wya4Ai/YTKOEFAOWPvkm+XG4DNlt5m+K8/ZZkwQsxQIaItCcjOhimF6y5pcUGmzg
MDhjDWb8MWyeOySGA0ouFqzs0ZHp4gn2CgOqwhADUvU3x0gxZqeuoU4PL2afWmsz
SNI1OJOvu/7IL/Pz7tHR4v/nFeN+BPG8dpH+ylaVHAK3t31J9tpxl1jq32lNBRRi
ZC2Iq6WDmECRmaPi7f7eC5SUtxJUyooAVU/t1NSts14B6q8fqH4Nvt5c1/CF5d4O
qcDMoCy8H0I3bXSZzLgI6zF1oggI8s2vJG/x+4leWpYtIE/javzB4JxN21ci4f0b
Ujti6HUnUWTYINkmg5x/wHimDHpZiAvYovcL6ZymkBZwEZG8ifxsf29JfaKxw8iP
s0n9ooQYcgPmUeRR4ls0SOcsAfD+fzUNQzWZufufswDNCyms8DjL5GYJZWTXOvMq
4OPAyzQpJ38yCbnljAlhjEcnRkU0cCsIn5xIJY+/wln0ajmWV5pK74hHLtr0xMMB
oc22kpQL/INTW7tJB06AhPfTiivYUNywj6QK+sgQl6nGY31ZV/vIv1hH3s61YXTG
A8kwY5k/Wr048CGCRPwITEwk6LZYX8cy4LN6r9r+0M9yoiVIK34PFVKf1euCTV24
d2Qt2FXgwb03x9/I2m9fQXmAdL8zMci0EN6QG4OizQuBcI9nKMwleBDO3xOoZggA
OKBJUDw9mbBp2LiScCtfgSND+rHBJFklL5LXmJ0hJ9f3E9neE4BQb06I1aQ0Rax+
f4ol6JL2anh8jFaLujVgd6nMfxRy0h50lsw4woMIp1g7H9hOoEMgTxn5sZVOJyuj
WIXeUGztSFOlrU9xtmNpJi4SE+dsPe4GFGVHSf+64fsk+mqdZIoOIxLnP7H8nVNy
BVlV9dCe3ULZWsI5EY1VmGVXzzl6+05V6nyv68sxdN/SPbxpYzQVQRJEyg/yOMmS
Id1pO+xzzZF6sUHjP2aSKn8n2va9FVuUOFO5QjzgLB0SFk/6SQLgXvjU6SqJfYuX
k/mVjpVIklaaq5Tf2WJTmBFy6p1NxkMs7DtCm24mtMayQM0zEjEuuVecxdzrltfG
VKsHbHr29qn8bnqixFgzWHLUdxgd2XTMgdFrYGPbYNiTO/p+ODv2zkBcA0tgqysu
C18ZkC99Krr96XD6RJf60KENDZIxRFcO04GFrlkNzJwWI+o7j3vHONN8PsAK5D+l
mhdlTuQ0lZBiEVKpHCOt3r5ooojnut/DvoUd9S87LTLyOBxnEG//UMuFjHH0ZO59
8K36RVEB9HBfEiXWVRMpDd+bDT8hPj/s+DMxbTbTbBAKjnwUd5/f5YiC00lO1nLI
z7MEQo1S0GN52NxUwa7wlJ18wN4vEY9zeUJCIB7j0Mgk04wwuAZ/wEIT5pHfvw3x
yOkdwumYy8CRkZWrjAWWO3B3OeHdCK4CdliyyToEkyq0OlGo2xpbR38Wd7fv4opi
zh/sJX+FP2Wk2Lq2/uaRLIsH9f/yiLSr1dp4uAws30lkgpPdL+KgVfqPC4ZWVgTA
XYLCrj9ZPXne2+qCrvkFZdyxEpmbAWxcOdV6qALhON6Yma3BO4vz/Ezr43w7EBdy
DmVs5Qrvzh8aliWUcXFA8v51n5JyeNV4IxXQYgWxKLU/OTvIuDmr8v8HXeG2XCDP
lyfLOUyqQZezaKcDEA+hISuLk5U+wNlqd0JkV/cMWZ4B+U4O4UVfGGZsbuSw0hWI
p8YOK2Ldfugnms4oJwxKAnz7zM3TBl8l2tN99JKHgk67JUQJINjxbBrP+/DZk9tO
dq4CoSuDhqMeFQJ1QjJyIcwnFY0hlZc6byKel9Maih0EvAHbps9y7wMsTeE/tgqf
xb5760X8cO1jx4J50mBxsWZhtAHsTaYTUbDW9N/E0KTL+QAxk6CkVPph4I2YjC9+
I71BtTV3MER4OXunvLi1vnzcPkpWXaYH8FSGS9ap8h2aPK9AzMzUxlXQux6eBlCz
GooL0eeW7yHe/3y0j5Gmg9T78YXTPk9ja9VMbgxnslpyOe7Tku4SA4tV6F/HBmOv
1OEcvY5uRE1CTzIu8tQw7ECi7T95obiYa4vJiJ6qzduXi6OUCJbTtaQgdPqC1AGW
MLR44zKY2AJHJSAdmb+OVLAeF3jUU0H39zjizm0ZeRYg4gqKLK9wGdoS37cYLAS6
GBZYAxJw6CBowY3IiucpTbP28/GH+XPYspTFdtTKAx4bpX0ihOyQoCOHLcEYvL9I
o620fVcPEAjQtKBwcnq5OLbQV8+uD1EqMuu1CvWeck5N+p3bXdjrW9RMdx75Olyr
bEGjrWJhZrUPi3pwIwDX7F4NqsvrAJRTohMDqCtVb317ppJQJUK2amvot6zBRM91
TQysE62r5DzHY/uHQDKvk+hRE5BdKpMNvbyGrVODw/p9O/EO8os9C6YW0D+Kvz6X
DJ/c6ih19fEGDcCnLHnIFe2YeXkdVNBk+iLdqDN8MBTwsA53mhMHnDJxunVbFB+g
8PXahfS3VVkYsIS8zY50V40w4hKCeQwj+rs0PRRnFUpP/vp5KWk99LoRwrazyYnv
BUaNhXOA0E1DW4NPdVbKUItUeBL+FZuWkBg1vyTN5BLQI0jgzp9ddGzuUaQqh4kC
79h2/6TCKP+oGg971Hy920Ovp5WL7DTkdWDuEKsNgb44ZL2rnwY7lN7R3HHbjx8k
f+ybzEAJts3HvmH5Yjg3JDbbK6cT8JWy88Y7sC9z4T7hm2K4hP9k5NLgLVROmH7x
oJ6KMaB3feYkKS8WCJFrzhi484c6McV9sFEwf9jLr/eEM1LsIm9DFAiEtOA30JKD
LdZ1MY9Vjug8+dREBmE3+pz2ItjtlAN6VTfCW227PFWVOkTgySyFor4uvOp+V/zd
sA4K/s9vDFeHznrazB0Pnq2Yf40Zj5ZM2JeDAV3TPG0IYqrxtKDd/9lzPTvREYBW
fogqQHaLv+3JHLkHBtnEbbPuIJ90qexf7cg/VY6cZ7bFj0RF8VZDHljLJUHCFhpv
2O3t6HwSWANEs+WyGiQQYZlBx1oE5SOJcKCM/kOb43GVAl0BJAWgHs3HSUSTkF4X
UGdC5fTcEYa+hGjPn4YYcZLlcnnpledVw1Lqb7i7MTj7f5k76Wc77fYSigLosGVX
Bx2VcgL0O/mTyzrse0gZBZrqZweYy9N3y5SmJ/tcYakBc+zQUG3opn8BT4MQBpAZ
ei4L6TLBjlY2n6EdDdysohASbuUv2Yotpyoynw1B3mZGsF8jJUa+o5PtovqbfQbp
PdK/bMvgK5oGbeH80G5Vgr+nXD3v04C3/7dOTGBQGOC53voRpaYp7joEPYh9Su0e
gefejo7mMdvVpBtJ2PmDkwfBS+/ekuuTiHvWd6vNYoaIZOr69noPQnqW2gg/esth
zAjuCNKNDl045beMCfaYU4pvcA/oNRTS7FGzVwjQFOi7KrQ45IERL8+BjKqQs81C
SqAGuTisZ+ZrJW+/zREg6tG4pTW7dRT2zIr5cPJWvjem4KkMIR+oDnhkp8CVQqSd
4j7WWNBMKA8nIhlaBfqYhzoRFeBuChr6acocx6l2FD5mNj4PqdkM4kpL2hIaU6za
op2xC6jjcE+qbLuvtISYZ02PtpZVcixfsFCPygiQ6e60lVIyeNWtAQxpSQA1o6rA
psi9LnC9oEEhjC0RTw/iU9yaAJjzNZxw96TkAxXXFe7ClxwFVxRNjT/iDfutDbnK
OmLyveh/PlYXmvQMXKfgZLyb1xG7ECUMVx9lP9pdUfzJ4I2qaXukfWGc5Gb7Ovrp
ttCMEhqmMxc4VqA/Nr2APefIZoD2bu9LuiCLMksU77FynXy453lwDbvMsVzGdaYY
ioNIN8sSiff/jbD6ZjYEn9K4bEP+BQO2Tzk0yXhkFZvUFNXm80AjuJUU2jznBYgG
p5DQ+jSKblU2aqBFfgETVKoIlUVhimfiSW08SCrMXHJUCAAbfDpksrLD2rVh1ytQ
W9BhhY8EXyqzKuv3KABrJ3++cHgUMcAV7V8b58opUXpI+rkREIwePKNVst3L6hD6
M9uVToZeWuC50Fp240WtPvRzr+Nfzvz5Byi91nivkxh524jSdiYzkdm7coQgb+Ji
BMZAw9CbgTiebZvGpds7BO8zBrbfWi6jcqfnfh0ithfvq21wySIsveutxwISfEjO
ICC8jcc3v6JYN0NuCn8DBjDVIAcHKlcVyh3qsD43hYxDwgRMheG9QvS/KnvavTP7
WOPW9Sk+Ext42O3Y51luI9HNbXpwYtmwIWWZdavSHLCrmLUnTsV1FY0cngRz2qlM
Mug4+/Q2CAmiTlAshxa3t2g6uE8jBp+pWmSQ3ppoLL5kPSoAOUHam9asCRo9C548
CRuowZ2awuaEaihj9w+Np3uMTCCM9Y+MIbEr/WApgHD4rwOcgBoA6AnNl9WPmIow
faQ9HJQjuiiDRExz0LMzQ8ZY1aalhEluuTVR85kspz6YHDFWHX7Zu1G4u/FD7SUY
vZ6Yvsm9FT2d5W5NqRGC8Ulhyao4K1oIc9J/fjYkPXpbSPKwgml6gH4o2FsxXQoS
DTbw7VnQp/sasm4L0IzWE4trXmgsKgtvElwFYxjpXd64W1gtsqNbS+m5/nSFab/i
L/+qDp/kt3XgjwDz7Jl8jzXxmERdomnaC+KjFqHyse3wetaevpJ8KWlOlCWJQMba
KU/xN5R4lgXvI5NTly6+HGo8plTmP3voWxRl8cGeB5xNCIm3bYWGb3Eo34vH3yYb
8MMSP8EQuYzherhsJkh9W0o4z/ggfecdQFwT1bMwPsrx8LqQzcOf2/9L+Px2Z6NK
a1ufegThKrg0nw24vTUJSIZHFNWT5170qRdSMMTgsFp7ciYc/3ev6d6QkypKqFz2
jbjahBwa/9XU6d4NEA4DWJJ+N50D4B3wyRSL8Q4weW79UpDAmpzvb3MbQ+w/1a/e
WJoVNL8Oay+761uV65C4sp0WlMcY4yEiRupyv/CQDphu3w60s+bgOc9quzCwBb66
Mnl2FXPy7W6rh95PE0mUjuGRB7pbHkryOG4fX6UzHJBG/CanzaPsZJr6grMVasf7
X/o/Vla20cCXSHj15sNA9oX2X4JabQzv2xqNqODiq2CWwM7QTV3+tzTvXwGNSNTH
THA8gotq48HBJO0whpRhyF2gcjMqSs6cIFlHPtMJ4v5doosKA6wq1aZwUqRm/lEq
xkc4kjSNn6OvnLv5XGKALQOAaF/cLlMQ+xWEcLkhBoklYV7ybqhpdfB/HU3knh97
e9jrmpADKGtXc5sXFpYOHVfHLoygOo183g8AagX+nWqQe/71tTtHpEl3AURuit5j
VVqsxSoAx1ZjicHVNr2lGR5AYJwzKNIRVLOHxf+fM19jhJUVhDGjHEiRxkq2NIPT
slapg7EfXsNm6Lgyb7xaD4HxwwX5ZCB3cZTUW6sPkLm+irIZih0hFWod4ee7k0IR
i7cJQMgqycdYJufGk3HYQMKQdsKfeUq7uJo2KAHX+mYKn1YhFUV/rVSAMwVUpFsA
4uOIvcox9SrJWF1XNH3BQXcLmCpK31IHiO8eFZmatcMrg2y06hmLnLz2naZHT5NL
1zgg+4U6HGml1RAZXJgX/nvZyvazMY/0QTOmTpzD3JqoYxE14UWkSS5jso7+7T2t
Y1W5/L1xS6nL7g+rrKfnoTsEkieLxZZW80eAYMSZVfK/wcSkCdOcCDEwTYvgmXDm
/W67JLWqmOAJpj9Q0UrlaaZs33w+qvZdtifGXLzt1S0MYJCPPnZK6UjzqvffWL7H
N5d6UxhISy+q+SUtVfLeOA8MltgE0wMcG+lcj0hY5gnLXDTUYSIg2Htke85cCHzD
Dkjpg0BwPNr0WstNK+uo+BtBW9yWafcIxXizjcxRZgQMBewQoPRpCUrhLJusMaiL
vTNDv6hw6r4OiiCvPJckmNs8LXgUtdqd/nhru29Oty/ATI8Uf77AaqQQ3g6lnFUd
b8X5+NXCX0OidDyWklv/7ena8AJjzM8aKgA60p9eV0c0LhVRpDLq4Grr2B7kN8aZ
fqSxtrxPpGGBESxf1eef9awmCuHuFwynCjSV9heGEECGau2inHg7H0PsIj7i+/Gx
DZC66YUwf+nYKkzhSJOUNKxOKrpwnhu1Ary50C//1CkfvVIZbBaZ5HigvghX0wms
ybJXIKqUN7kE8WU48EZJX24bfb0hO+zD7TljRMWSIRpjRrqMR/gusDVQF62d2dSC
OlOK7JM8d5HJJWJSAClRQyxR4obxP91ffg2Hn0lOlauxe83ZgxJeDyafQx9XJb6n
E6qKR6pLCKptVMt0L+hFhAZuvlpx4yVwNEq0KVbOVROIBGL1uUbNirtN04E2WUCY
Z91OOYQq9HLocXAjx7jqN9lCXk4VEGeESOVDTfhodDzp4bsyr5siIU23o4G982Rr
9tsRnMV0KSPPg1JqHh+GyRDtKtznzlkfCEuyxNGqFX3pE7XOR/KCzNMNFKb3hVqj
L4HiCYeV7/psrm+fxBImTetZrSKGWsBGuqYYhSVCrHKLWM6zA9AejwDRF5eEjgpS
1bVUqHqZpjvEHCmIAUBnbvodyd0WReH25Gxe59wLEa1xcdRmd054KH/jPhaUZnVH
avmcfyW7ksszaWFhpZDbskcoQQ8RVaTU/xzh7WVWQy6hJL+D81UPHL6kBHDCIIC4
kK2YhiyZWu7KwTHHCby0SGp+I/ky+pZq7QNiQmQsnK0nIGQYFYHKWLtfMBVAZh3p
vvi4Q83luQRnSiP4eHu/W0apIEIUT36DJLSXlaYAJYqmNQrphijEyQ9STgmZNNTd
xhHdaVHLmxuNE+lG3HXwpxN9vc1s06FnDsY/XtXouQTU2V9BeCLaEYcsCp4SxTCE
hipQ1cMRZBzqUYwZ3smTzDbIpGuldUL+7T97HxJHchDtOpwvtdVGe2XspYiyz1lb
5+XziXBVFItnr7FkWLHuWjXimUiMHBo9MV7W/kK530SE2Si6vlf7NTOYzZzMIVX5
E34Trj/+eWW4xuIX+fNtoD74fRZHz4RqsB9jr59ikagviAHLO6uoZb55cnaO8MsN
ONxDczX972fj5TJT7p1+F1Bkdw4dc4G1iPKj8vL91yX54q73RPv/9v/5H6NaTw7q
eGHrNKIo/9wHopAM5V6ZOWFSosIrhRmlOhXCXpFakxmvn1rKmFQih24pA/L7zaNS
QJmHjySrhMvgvauGa/xhCsP/z0oBDqtyLLQR5cUvq/zzvywa24YyUEc4DrahWLUg
FhMlMvwiph+AtR06VZHKn8EqdO342NlsTnHyJprcE3gKr/Dhx05GjzyQNYG98NYK
rxpFkrW2C8WmzEF+RWHx7QiMmOnU15+L5zYw/YuOrfsteW45Zt6QMxR+GvKNpDnx
cloG34nFq/uaq+yYU3Wz+bNVKp4vWOo306fCeKLaPx/xYCqPIxGoBladGnkL4A7A
V1fcL2rK4q+n1lGO/XfzUKI1Jubj0jC0u7++DrWepkhJ3Vv3pff8bB8qplrE3dIk
r8sdRMmpMuXAC5AZAbZjBtykOSmYCDv65RGImjRce2+8S7d7xnZGQ9caQAVHQCYH
OVoVjZRBQA6U27ch8lsZj0BA1e6qZT5+Dfi6S97IBLFeisXw555PMzny8uKVrS+g
lhNQ6E+9srj7p5jDoi/H8FLZWSvBm4BBQHkNhPm+zE45dOl0Dq7Cfm79tpSz2QHU
FcXFhG51ZfWrcfyJv0otbV1IMrsZCkoGBR2bSRjT2lTZc6lL1AHgVFqx/81c9KwJ
4ZHaBm11slYMBpGzFm/cOIyTfNR6P7GZ1789Jxa5WLY8//eiRJrPsDstrmCncJsN
4QPm6PAosm6yUUgReVpYQe8SYstc/oWSMuTsFJfkel6y/9n19I/bdd640jb4ndyW
1lJ+gwRY5A6NiE/sB7nNU6IshVQviyqrICGbrI9Lc9zWWHNEQ0DE1+NzvjwuYM1d
va8d8e4CUh25zq816TezA+KHEG13bDj1y88jf0w4jxPby77op1B8ErzGT+Kfj9iX
8eVUh63IWmstPc87CoiGMGXHP6OQfDdBdK59SC1uGowsc8yozcCWT4atSoyD5msp
I9rQORQUZgryArP57KEWrwj2pRJrxehvcOt7RQ5V4F1JcYo8iIiOdeowrjzBK8NA
Tzvy+cNG9InOwyvrG2HcgevKfAnbj+jdCP0l3gUrECvMSRZWcnH56RdnQeJYAB3g
5IFGuzWQtIxLLwos1m8wnz2nqAF2WN9IIzdMQHTjOMiJsmfQfXD+0Y/iqd8Aw2T/
GEEWOTy5VgmvJ+lCrjxVSDLdUxGgj3WVzkxIe+qNGzNKaoUqNGYxNwi3qCNORLVw
jPFaCmw9darJ1crNh/Th83zFBsZmmvIHuIpotpnIMhu+4R7oYjQOXU314SRUMeyw
XSKZoYb+x5wkvbQ0kwMbi8o4rtie2MEoNBLxiWS29RWCm4oLtl8D0BfzBuYZ7nhJ
TMSpL6Dd6PWM05Yphn+Jr7GKaLz23JYHli+pWqoA5Ogq/WeUFj20ghLtuYIQBISr
xWtWbOJxcMdPpf+YNih2qtp5XT0WImEmNIllnkyqNXceGs99ycHtV9ooP5tQrzWx
8Z39XKsEpHi00LVIO05be3NPZbTWCAv/FdvFWLKLWuvvw7X9jFZo8rV3B+52BCOV
3Qu5TFh9jNKaJi/NTb8K970pb0VZqSBQEk3wcFaAOLbbAEOCv6KOnbDKxwPpI3DK
DsuftspQY0BI70DHBw1/ZkDCe8cpP162SfniM/DP2vyOUqBnK18Sv02qk3E09moR
Kgyl7KQCwbBlyFd/4yNRgxSuuZB+LNSsadUGkVvvjQyMiGsoQcRiIIcLxn561aNA
CdR42hQ3BkAocVmf3Ff7xK1GakSp3+v5EfRCrreaR9e8b/Kc22X9B8dxYjPD6NdC
MT0HJ3MOUIhF1W7DGyX9VpEAsi//uo/bI7jsfAtlmDePQEFv7M3/05mk1XrX/zYy
QCK8/wClSRkAJ/c8HxFng8vhLMpT7NpZK+dVeu57WpurweVDd3MeqjlQkG1IH4aF
qMqQYS68jLlscCve04yr8uT+2J9Hc5lfTt0wlyfGcRLFOWZ+dw3viL4p18S/2gmU
xtfNnGiHklGFhhUegaP7EoNYVwV33ZNCflr9AmNK9ynSl0xRe7YHIGPJ850xPN29
PINn/iz+T/0A17y1HhvONltw0XyYS+to9urUY1ZT1jAzvmZq8rUFHxmGxWmlkDvv
VcIo9YCGSJhz30SEdRXS7yq50MbO6JEL0OoTSHHQlgQbAvXBk8aafaclpqFmEIMa
68kPTdDvEj+yYBVgB+KdreW4sQkan0K4Uk041+oXiaV9CEnVcC0aOCwiDsB+9Obc
7d8lryv/+XFdij/sAp7m6YYahbmDiLyzDnrNTYYgMEfDp9kfIiUON+AEdV2LcsDs
cqqiM+q3gJY+3TxpPQ4Y1jSANziFzr+IMtLUG3RvwoRuxVGSZjEo59X41uu0hyeu
WZwvJRwQf/73fxiI+voQpwanzDNtEuGNFA8vdTb0PYh6gVLdmsq4dqd9lQ5Vde6y
GcLTxkPH1ZKcsi49ribKIEHzbFnxeGxoqkzPV366irM9/8kqwYHI9RDm88QWDHRb
iGM4Ge6Uyq8/15bCIZn/1ck1cPKlDtNE9Ne0vt/WBCofWml7p93Af5dm7hic7pHN
ztWYlx5lRctxp8EhMoPgANuhjhb2vh0nHlLf+rvwrXhgqfquVIAuxl1Wv6U8vssa
nehdSHMQNqo5Zmyp6HwwZ4yGV74s9PetDkGHzUgyI02wMD7eZNmIN57Z26usceSC
yWAl57+lgeczywVVVV/SsxZy1bcX3XxddPpakJ2/AvFHbG4FWconFCngNmr9TCpf
ekdQV+9VRsv7Zialt2Vh6yZJb34vadJRyp97yBkxWZBGoZMqobzaGW1xLlphsFrs
y12aqdLHlJnG+yoTIQMckFSfKhvSTXxG7t3Ck9z8WJw+Dm5vQGQOqOMUWDCD+/3I
EhZWqNh4NP7VYyL6NGfTPcVLImRgcY0hlnpekO86dca1f/NddQtUPzQwyUGT8d3T
mXD7UCJARk6THzcRrVEscbohbBETnr+4vSYDEAB+LsfwuFADc5beSFzpw2TD1dYU
OpLjCtIbxzrFXNYYGiRgc/Pye4Qda5OXaaCNYxgIICQ8O9ORX4at1B81zmUBcAx6
n+XvgffR5gVzP5S0m0dKLGevGoAhHApCn3Lkn5Ol+5DG6psI/nH8VmIfYZlLe+x2
RMbVOq428jXOauxnULtohJgn2YmsIQYpMEhStklp4DsdOneqV6nQ1eQrMXiAHXde
3vNcCv9LWna8xWVXc3traT57ayi4XsegjfTQ0+p4fGSs/9+BUtCRZq2IemiYRfGo
+PHTVI8h9iCScnpg7Q7mSNWbgdqpgOvjO2CWtzAeWsxKgnn49YmbUxEX9hMA2jiF
GTk6FdyMEyxLX/xp51XV4kM/Qa4uDpkzVTHhgNj2+Zky5093XKWZD/cmhbt6+bBm
89l1KbApoZJM6GChtBBjl1iSVPTZBZs8TuH1+IwjNF2UnZJsI5Blh7MutMslW0je
Bnbe/9enEeYMGbaIAfDC37IngwhWrE5elwbZpN1ebnpVjSfbeNfmFijgBL0o35SL
iCvgjlmjjK3C9r6DwN7ir9+AM28SgwOyykNSJidCwCMTdUnYM8DZnleBd0aZCwc+
JS6DxxEyWyuUd7kDYUM2mMCYNyAFMPd5FbaO2YOBUhWd9zCQi4i8OWCQWPu+h52q
TJcfBTj/KZKU5KyZaIfWnuft3dFk34P+G8sFzPK+45eqBkZng31glfFXtnPBbcg+
wkTXsCZLRwP87o64XCuyLvWNqEd9WxKW3iQcepUPoiECLTZ1fqEZ3fEY+znTbuut
IolLDvQSgRyqwq5rSWOagwSBYUdIwFs9TL2n9qNKW1EGZoPsE6IjNRdBWcJOddKa
giFr2hxN4RU2om7t7ODQYfq1WbigZSHNB571JweK5TecsGGjjnnWxfJ5w7HooKlP
GaL1xncDyUZfDCakuRXIDkqw5FGBOjIwK/7ARIHuGnIiKGCtpOOvzIZ1HmgBnLd7
Ftm57Ad9GhY5VA84LmM+Kv77s6ZTqN5wXEATBY2bI6fAu1ge51Bzk+WHHE5ulF56
nJFO/GyFcxxXZs+Ko/hkcfoJ5aRta1zIYACqMMfhNajfp21pFQ0ZsyWhGpkCYgNW
24wTs1opy6JRbh4m67SfeCbgdnulNBYYufXLoUJSKKfhbLq0FYPfZNhOiu+cvsdm
3RAIa63Dny1/ERhMfzTVY73CurtJ/8B8BQiOvvQCytNy0+Aj1SBHuPR39OstrOWx
y6XLP3oBqu9K/agWs3jXQoUFzgc+Echu64RigOplKzrL+JFVbpZw/6pOU45fopzj
V2iiu6UHMw6ocINwSBGDndwx/2FggTQ93IGABRTqVn8EzJWgDrOZrP8Zb4bMGiuQ
3Z+DrdCU3dM2QODo1udS+auaL2Iu8FXMP5P+w6mnm1kyq5YIekbBPVg+n2UrXgcl
imPthk+7jIU5E99Kvui02gv0xR34NXEiTLp65jkeWdFzsKPw5l50kQIIt3qwNqFd
mvKNDxyJ7u6erPQvsm69iTGzgor8g6MEpMoYAKimhl9dunW+x2iSqPeMazIPE2cT
4uu5EH61gPkFslYB82xPOZ5MLpmk0BKCwDQ3TghA6z8z20XFUx7sfKNV3N1OFQVw
sbWNQ2WfU9doHHUlwV2tlfcxo1Cp3JWX8PW/EX2+T4rD6Xz+wrC2hMeJccHHT5NZ
/eyNfNjwLTC4Giu5LIHsywPLch6/E+drCC3FfYaH5+3vj0hdfAOlYIzvwcoNis3X
ymPGaULevEc8vu4JP7k7KUf2a4Auphv4YhsXabmxWPrc6txLNZbyk2qAYU7yZZ/b
a3Jr7iOrrTo5ji+IV99nIGo8Yd3QX+Xdpf+1gl9iAMy7yo+llpNe20Z70GuGkWam
32SKs8Nyo0mtUdOg/0qqssuwVGKZ7lQbqqgFcwEtF+fXvylGbbDE8Kw+GjIvNRkJ
nWhrVfnS6RHdLQy+fo1dJ3TYjfTA+bWzFYDZe2+MJToQ8MnFcwey3U0cdf6+MOc1
r94U4CLn+zO1q2t44gabFCBGbcmvd3gPFpTvC8wGkQ6tegl6UizC/ccmYXBxgv2P
Ec3rsj7tLtOAf3ElFH3l6smdt7IyX5SFX9z6K1XGawtToQUEvM2qy4A+f0ia06TY
OEDg1BDxqKAR6j0hULbSRaGeOBfMNvshU6E9aqTDG1fWy5R1kGbRlEEuMH78F2vL
vGp0IP0Sooel+RiG119c/FLg2GrdLaQD+gtOLELnaBnM/ryfVaGIIkKvJ9prgVYi
DjJbjNyg8OBRHZn1cnV7Rph/CYuwX3AL5vWl1Mq32MYWBHhBAObpIKPE31YlE6GE
KGUMJvQsIWGvRqMka9A0KsTYDv46YzqjfWCL36JlngD3Se47dx9CidjN9dKXhOeq
8y3XQwdAF1sWuuuIyUU+EwWLdm/tcunlv/PPX8zaDkl2zYDNxNvo97IgBl5Et0zO
eV25z0j00hVenuGK17pENggLsJhuDjee0WgVjY9IKpWKtL516jG2oV3WpG5OnFNu
KxCW2Fw3UeRhMJOldp4DZDsc54NmW7E42rOpHzKar0UZNrtZmpR/SwFGVHAlAGZP
cLM5vMeZ9kHyKxX0t/DkC7/Tr7oCBUwodeN/OqTquwYa81UkUzIVkiAZ6ezmoP+Y
8SCkMIVC116fsLdg2Bhs0TjL+Or25KMf5vuxw3rrSDSENb2AQU1FRTDjCwMeGnc4
XMc4pYfiVbf8R29hwaGevrWGc2VVR3f2Hh4dSOPxFymGXOp6+md6jNQw+RkqTUpI
YBdFK8ejDNbGztGuMb3YDRL1Z0R/mJ+1Iu5SWv1Ci2r0e8DzQwlZX4BEQ81JvAMs
6rb1b7R5k+xt205JBYWE4SuKokmiCFbU1r7BXtWCoADRlbnnyiYogQcKabfY1yQk
meX4sTWLeuwGWs5GzkYIn5PPhP8nXzyu4fgu0lb3IcJY48FIyYATWiSQUzw0G4U+
dOf7fXZvWJvxxowiH8FMfv17Dr7QIiz/ZXMjv3xv1bfZN8UWQZcgl1LeYF+eZUUR
rSBh6ZeW31B3OcE+TmjM4aoESCnYt62eiXdZ594dAcAyLMLnBIQS3o5n8fRowaQ9
d6qdMFqvkAsVxRYgdWqcb2S1GC1VvqUlzmC2qr7eLHFo/nmgETlaEwnfUgsZ/WJH
EA4ZDF+kYh/pGQh62u9cU5vvpY3K5AIwQbla3nYqmI1SpDqxohXCfsqlOE/gOYSs
Khj1f3ClQV5HbTBjJOf5bGOCU1ubO3bWcthLvYA9CdNWoNAH920VSLQxloudSyZG
sM4s780M6/5Zn9mVMyC+GDp2d6Mlo5MPvGPyR45jAuX22xkgTqMr3GvD5YbJi0VN
us7dDazFoCM1DyAn2OiehT8Oa+f9xNjwa0B5Jf63PHXPmSYdMppgej/D8izMiYGQ
bZaKllBCh0plY9rptSr6JmUS14ddKQaRzemNLf+qHZhh2wDJC4lowhLdG/KywX8n
X9RlL6KL3TfHKRiwnGARv9qykgM36Lq0z7obfD0t2ZJXOuIQz8cnQGtJpkpPc1Ko
UhRyJLzV87XTcK53SfMExTPZBMMcvQFpZc0DbflizXmK7vrax+J3AuWWGdqLAvKM
GfnE5FKKR5MlPbrz6ZlNW1NVzQk2WBgUmMT0zDK3fc4ZjVfiTVWsBuYLGoIHceY+
o6ZtxsZnVU43OS1D0jYOtSXID2EVDgAA/VRR2Rq6xihph8ssHUalz4TD8+rPTq/u
wAsPUMZFI1yOataNIITBnOJ9I+dSua4JjAZIDUQ5AlRDN1wQEQyEi4eSXkiaoT8Y
JgjUMbjw294d7/1obsYTsjz6qTBpyV62C8G159MjkCSHexnS+0/SBY6WUFFUR5Up
HON6waIQ104cVRooUru4Vm/zW52jB9529xYUOo2IBcX0VVk1yV4Pm6oZCGgbg/xK
iw9iav1NOoY4wO6Iw1o5x3CIuEzMT7vuG4vRuh4Cciaecn6OL870vbUbqFc2d5DY
WIHmLlxcT0L7mYGiX9N3kRB3ndXYYBjpLEtNKkbNUcG9qonE6mcF28ZlgaDfha7y
Ha3DPfrbRgyUEA0elAIoBTNHGm8N2OV+s9HoTm1gkw6aSmR6zjrjVVMYoD33AvCF
Hp/E7kwAjQOPtkmVj9vj2W+g5vs2LWfCwM+b3MSrLe04cV+KdrlXpXEMB//Qnkye
lJokQGiuNcPOX97ULr7zawOGOb0KxXz4s9znQjEc41QzI+23DWLaQYWuf9PwtXoM
IstQQCSbLivpSQtzOePNqkruiXHEO9WyDO7YWLfDcm2IKkvWxt9oZXYSvypHlFWD
FcF4OEceB9dVGrX94N39jeCatxx7FH0+dE4bfP4RwdgRcnW8dJ5qfO/X2mFVsAJZ
NmmeXqHQ9Won0j1B+HttYA/69d0nxWcGxnWk3QyoZ64H37AIvxQfjqDa2LLRqovX
ZEDARS4WzgH8W3cYzA0ifHsEzvjfmfW7UZHPdZj0k3/yKRmSdB113hgQ+N450d5x
pOfzNZ8sktEwDnbb3f3oWN5ZA4ooOP6zTujXjHJhcxmYQrzOi6coHTTng2J6dY2m
444YmXToD6Wmw40BwzR/o0H/TgGXUFnK+WMPSgf7Xf4oMmA+hqBj5FKySWiUgODG
ti6IYFSKTq2dDb+AAZ+BSgOFCFk4d0XACxHS7BfpjqLoXLU1AVG4Vi2GwIaunL8I
99ZER6vEKNejEivvaA5jau4v7ZWiO3wVIh7UxgrOyJzdyAjeDExG3Wmi9z5+JnCv
OW7e2ahHRae3ThqDfGXSH2bRN8mnaNH6F+NVTq8PWI/zZ3wyvn1wOntMxP648U12
fOPqwu1HdaI5FlrQY3sqI0ircGzyJ1WUYvPOlYj8P9WXERZPdTRfnPldBO4DzQ+8
fZF8nFTTCqP969iyzXoeiaLb8hoeklsQJfHBYZw5BjQJhgsZm8k3KGY9wNcMgyEN
L+vlUwXMcKDC5HGex6PcWYkWtbSg19xMcoyU3FLCQk/jNmedtl8h8trzUnJHCQQW
MckvYIiNLRx4jwJE3MGWsjl/EspecvAqvYSv/sJktq8BqIx0LufVCcA3r8D/doWS
UJs6DUU0Swh6pw8X/NkfoXYZ79yE+e/9BdUzGtge2UcqwAaEogSYhkz/sCrIURL9
aXdJ4plvtaYrXksGM3rTB70kH1/EI2pZ1WvBxA4cQ/mlE0dLS7eb9J1puz9/tLmS
oNvi9teXtTaB7OAZeNS/XgbJ0O5VOyjsBdFrCjk7llkvHrMYIika4q+8bLvsOV98
8bTdmIvJQezz++23wmttcTqJQHmL/kwJusUnhS3lO7jITH98hTgXbYGzSuDd14Ai
91nLWdttpKor0U7G61ql75CELm/aJm+6gvmqRUXqGGwBeeYJIHmKYoYr/5CjzW6S
66Z+W7DhyLCSV8KP2eDp/KygYspMBQ8tB7agYHr2PsxBH+DTf30Uv13PY8lW/N+a
N5mHM06kvEeD0KMYSgNTsieexD3+0Lu7sAplDUqRv0GTxIz7m1xw9gRyPeFqrKM7
1PTlGF421P1eL9VZ4bMqTaNM2CKN/oXMyLtx0vrhewByX8QYqrH9w0Ff+X2fU6Vq
anwP+v91/BVFVopir63og6zi+quQc0CfhpCWMokuhu0JYtaqu4yNJU0C1Vi5ePr1
MWIiZTaC73p2cCDbnyfFTK0P9YzEJZv2HtcKpdnwy3BmyNnHUOGsNsueGR3qpUdu
BLY0cKWceFWUMVsJ64heEHHe+7pZ6NPNse6K8jFArnNhI6i4TEvzQOAypECr24gE
oCqdGdULSn8B0xR9KXUmigOdxjFkFDkiJdHLjKDWvGyOdb9Yp1jMbrLkvaefpeTb
nxkVjycqgIPutqKYhbTM11Ij0gnRnbwCP6hbBpLLrbwh9yKoaPBEKdCRnhSuqzbY
DCKUlZ+tXDLTjHzjH6jFuwyLl2tOuC+prWPyXG7fUd7SYHdCahqN+7/98Oh23jUV
0Zfat0dxowLZyECfJL0CDq4d4cXCb93Vrq5peaoOFG4tNDyH6VFVOpLZpqJRYYEH
yECcUsLwYXWfXUirfGtWeBJia+LVCcxc1PoiJRDHwbiRWC9up2BfnZqrJTEoluIE
U2oI3qorM/tlyt+Gu+L5tmx3qdyjBk4fQlVWK1azY/+KhW4BS4sYBSL6RRZQcsyw
/uh/2ZTvGT2JqyCmshLoTyHk7cGcoFsev2asfjKIKFWE5cILfrYOrUGfYxUiVUgH
BEOhRtbfbtDs4kKDChZ7XdvEsZ0Ig+dgixUBB2D/Jm4qiXPYtFdJ0p3TBF6i4PyE
bazO3nhz4Mi4lEA8oAW7Z5PCyaaNA5NB4YnjKQ/Sj9VapXTtwkb+aImVgfAYxlC+
68U9eET/2PXhoYf7v8tUKC6mTiAiTX1mAZbK/ZFoPM+LJpcuAS3sTAm2ophru/tx
1apMMP/nqgLK2kH4/lnlrHHcADz/DEdZiO3x/rrxhgyJgIuRIueJ0v9as+XT0LUL
L6jUe03shfnijRecGquzYpbaHZisKDJW5xqAWkMNdayJmqef2ne8mlDCL7+lWlm9
Qd6WZ2nkxLfMKlRhId5jaMm/wnK3dNC2UitJuQomXVeh6oXAtR4mEtygnFsZiGtt
igxwW9/zngH/6ZNAZPTwtEkKuailA8mz3IIV7E/Ju7UPUtagre+TiXKRb2f21O1/
zs3YKtX9aeQxX788u7Jbu+A3mX63m0vfNxIYribQCwKHj7c0dmfi0cYV2/m3XQpb
cpWvTrKjNMbdNL2N9oejGqWn1a/iaGs/NRH+qgNXUDbaBN2FAXGV5C+WZhPmDirk
tKTXmoz2v77WUHKyXodpZFbbhZ+SyxKXUBbudqE8NFTn0BCLgOM48Lqnlx8T5sPK
8lqDjHqIJNEGDGjRzeacE6hUCGfNYl0wKkygWbcFBtTwKbxtYKvWs0jA0j8+xCmq
7dnt32omfE7dgVU26YOpabydsvVOogI6p7H/b3iwsAM9THblCq0NrJY19HRLky8h
+knoKCVwLql44NYVgWnSbvai6vWE1buA/g2TBq1wR2eTTkTBWs497nr6hTs8pJo1
c94L0sfTsoqCx9HUPPHnn12YyBZDH9iZRNajVYf3M45jtkw8LGBqAKr7f0QXegUM
+4kIzZ3MgR9ZTxfm+ZAl0EEeFTkx2USTsejYj92eO9jQDZsZlTtz0m5cCWzgfAfC
f4LmYf2iTY+igFx66sXwLzGR+if2PXXvbChwEw30Ok52NdzpgRXlhHzqTLGzres3
82O22dnC56RftvBztcp25IiCM3A8/6iXL+ZRvoKpYrDBoOFWBCJrsUJDNJPn1mt3
kUoIrovMn9X5YTkFnCHQqW2qtMDfejx+YhgYuJbCLdZwqRU/hEXEgAqvzYTOXjJ0
JP8ma2TkSyj5tS7kDUm5CQ7lcEZFWuVTfZDhSEOTwd3I5qqGqOGxs4Y96qOHm2fO
Fkoy0JWHWlU/BBu5MpVk5bmesp7fMD+57fj1qvA+g+gnS+YCpp9bP3dtjWUoSrA2
kE0UvROeCNFNkcSUZtYYIpOhmXEVdl/v2w3jXBqBY9ViPSoUXIOjZsUVw9BdaDBh
Ld5u1eEsn8yNZ7lgUXezLIM52jqVvnoR8zNBBILZeRW0JENUeqqO0ueoC684FKLZ
1zGI/2KIAFTlNNzSjSC6x6ky1m9Cyvml1R6mrgcEarlNaV/bkWqIg0GHeZJ6U6+H
CIren0JPCpd4Sm0Jdsv+A4DERPnzQbE7c3fioQ34WUd66oBFjHVVRzvgYJwTNMcf
SxQ8nexRduNbwLTOB8cQSIqHDe68u721E/g+dA1Wa3f721rZus8snpVgISmbIDZT
lUT6mcWnsI2LDetOB0bkDGHKagniKxOkbuHPzzJ/rkQAEJEW4aoYEhcaegd8RT5m
WYOdsTaTFxHwc0HJqnQFJSmppMJ8dCo10AEOGRChLoGnlQdIxLp0sSD4r9DIau7x
nvG5wm2tGYWC+zuWNzOlc5HOd/ZspNMD8Qyb+DQtnVvs0jEnwzAqtI9XUUBZ9P7j
edZ0JZA3WbqfDGZzVQKKF5zDRfLdrKLV9MSVKcfguCwkxQv60r8KVmXnIPy6A4HD
AYKTtF7e7qB5Tb2pqQrNY3HymTbm68BUY6aay1pRvsGM1jwG7nOk1nv7G6TQIgWu
rrFCUcmtKYa+jOjC1U3v5prfCO++qgIDCccAghVMT2mRF3Jo5VpbZV0OfWMW83uE
dsAWVeWNU1CiqTIciZCir6htF+MhM4yyWdBKkT11gU+oY/+ffdl7VPnkiBLPML/b
+fWx21B51BHyRwJTe0gH7XbBsM9HrCvufW3BNxfl0D2oDHaxhEhXYvUBRD+x+NNW
OVXdDqWgdSNsmCr4m6I3m59+pFdWZxMyYnlEn54Xyqnnbtjdnrv8VshZSTjYWnTv
pT2CmajIR5I4bX4og7I0b9w+3DyHnCWtTTI2r98w00N8sRxnKZOP4Md8bUSD/b13
w1KZ5378wvwDkBPBUwcyl7QWXZN9eK/y7jIPJU0jj068B7fYUhvNFTGZ7K++ofsJ
Y6kxfBlkVwDuvuxN9ySVIXxTQ7oKNltA0VuEgSupPEcE6xJuo+hQPatWQf26Wbtd
Vvf0WuMnPM/tOVgKnwTlK1zAzpanfbRK3N/rd51TtVhsK6SRwmb85bn3ujx534lT
V/NFbAZL6ziDwxslFaMoEpDSgIdEWZmdHIo0QQOYifabXzhGjoBwUCDrIevDZBI8
yw40e+CNMMe+qSVOWwBanD8jW72CgKYJE9jhq8nbIl69W7qN4Dj4S/HreyOGMtgA
Al7BJLi9x6LQ3gED5lQLBRsrFXqNxr4kMwn6DqOC3F9QovTNqds+ea5ZvaSQXw7Z
TZvxrpADZzFQ7C9X4THpHyXzKIpr93lMeh/HpMEEv1Y+O/mmdEVexPWyeVLKFIVI
aqLvo9g126e/CR9awWBubwDYu4myHsD4KYi+R/+vMNLfP6YNMapAMBprvDe3JKSY
nCJgpqnEX5f3FVyAxJ1xGMxEuwkYbgS295uFmsPwJlkafwV4Fcy1DqygIjnnqI00
Ql2WZgTLP9uKl7NNT8xNSpOYZc3mKIG5+fZOMA1Kg82OXZArHm7vbOv7K86dTSBd
h3FufX6j4MN/7R9fsDwaBhxrBZNudN+9q6WcOz7It5jZCKX2qjltY7e+1qIhF2Db
nbZ+uXPjSRBumN7dND5yC0yeFPwQ8eFwMjCJ1y4T9bFb+CH5EgP0y6r63zKwwDj0
Wm7u03KU0kTVNwxtswChulR2Iea/4BGY46AsM0BYvDwMII/JzhYAZPGOjnnn+2FU
jNYPhxeXDF8FThGFMh6yVl/4t1AktcteK2vWHtccyNvbCe/kVjuIZivGnVY3Y4Q+
FQRmnju6rYvOQnz+x2aguKgNv4nerGQFqHFADKfrpNHMGeIYZFKU9qR1b7zoA0v0
Tm3js5j0gUBqHcynve8l6L0Aj11OsqdJcC0BK/AI4WkM5CuY+xBxlYzAud7aSipI
qpnvpEIBQl9nG3DGqkiWM0kH4re6FXCLsltEuAiz5OsiPCmXbPluVhExMx5m6wOz
lPeoNs4VIehCxcHsDnOV2LLtN0/0iv6QRYw5+l8Yg0ASgFAfhicqH5apO/Mbodxs
ys66LgJF1xKUdGiJ02zk18q3WQstqPeUUm32BxkvkAfK9F08eTqJhZGGXiiUroJW
OUjxkYahq6cQO4tlcY2xIvhAt0LUOYv6epZdW/mi7MShGKN8KC15O0LMB1OmUMHH
cHKPQv9K0DuhA6Ps66/WNhrZh53I4PSP/PPGTv+rL3J6cXrdyCJ6UTYyuYhcMK28
+z2BtppmzsKmZSQOlbEY2folwnDU9XEhtP/ZKOuIcUTAri6SX8o1irUddL0Hz+i8
+3gwwhlVnpCftNaCxH0Ryb2EKGEwB+mTsy+Jnu/qgo/6beX0WVHNPVQ3XmXX0ezm
ALLFBVcbdlTjJAknldPT7QQCIyxSNGLMGTKJtRPfwIjAk2tfg8qV8DSNlEg+7r0J
Y9Lhg1cjRlbw3YYd1jPXroXeQ+zTm8xjOHLWNWBDkIGtWumstO49px8IGixNfzcX
NPXm5EO3Re3PZhOCBpuTDbruehmtqmJJCJvon9kQu8BxJwKahiBhHO//4iFR7+dv
RB36BjL7HsHXDmXujXN4dAl0TIGMMHHjX2/hxoNVrngdAvl0tR+aZxjnb9gVmz1c
BbIqpLcQ5Qc0mhKn0fAyI+Pm6ZPoo1xvcC4Qttb0hkuJr7gJmJSWNIi6xN7TSYBZ
2MPN1YzG43bi6dvDNWxKDlarRAp9cpqTlApDFTS3iSle3wjFrBGrfmA2nwQvKtuf
NuYSLFQQdI3PKipYFu9pZbIyrFzmHifWJBzt3LVNWUbE+2PmC3Rwt27QyJi0ocF9
Nh2rlZmAQr3YWdJMlopYDV+suQbzCRg7tNppIDDoa15YckfagugOUQi7atZQVXm5
idr9+ySRdPuLF6seffwpRgdJdzc+ssARmnKHPeh27wGl11mqC7En71VoHSTqlWwQ
e+YAiDJnlr31Y6IeZi1f4442snGjtVz+GAO2HtLffG+uz+Zhwd+29yjpoKsI6SnR
6M4SF3oEEzrs5h99jrO5AW/0Q00zZ2iTEbiwg2AmGeFg7kqqgPidnVl7Edh+fwRS
PX/m7oV+Rg+6MObArLfXePuS/qHR7vlMMOgnYMByCdl+1w4NuWUqB6lk2aWrqVpR
1RQY/zbw5lMlsIPhnN2IQIh02Levv8iGr7e/CLTdzoVip7lzOe+9/dzn8ALPXRQR
obxGX2bAeK7ana9VFqqL7QvQ6U8PFCXRVUgdsmZfBuZOHLHClvouOcJxosMRqGQw
Pf3nqPvqze9fwEISPmY2yGZIxHVVC+cLLLJirVhYAk0wLn2TGMdKRyAIhYKQICNS
0mBK8KTCuUyULOARWBCSHnJpgGF5oNrM1UPs0N5I097xrAGQzK64fuq6KHvLMCVP
xhxHX/3SMw8IQxjdUhicfmtX2kLByr7+s4OPaGD+fmexKVmN2/9YamAUceLoARsz
5K+TSraDbUH9t8wFRdMWhvf3zMGUchi0+QY41WllIpmyCUPyIqFTBQ8jVjvRkfbz
FRgmksVwChMEkS95n2TMzgDhaXF80XKJ8SvNc+WlfRQTAPWKjpl5UGMELUYDm0xS
KCMDfVXLdhwlU4uoJSkir+HoYlQX3KBC7UiPWMoCIsZWZPkvgvTbDqtBTH4HV8N3
J7ap85sIBoEGVYcX/Ybr5xVylMSuaBI1ETGmxkHlLHQWyKoMDzPvXdqUmfOapxWN
P53o/KY9zE/+yezzyogNR4GwK7CDaqr5mzuxtlOhcUbCcxAr1lRRIF/kx93OLaz4
363zfkXaXUUtzc7mA7XFA+nwfs3rTyXMtBQcNZe8SM2eUtU0CGNjkz/jmDaJ3QXx
ZlpoFGCzNnA8ulxUBAnVddxx1BdaPS2ekiFV6/9Il6eqHctUrwhgcZ/n+ks1t0Wx
N02KRkZRPzN3AODwOjZtfjspb0lT24/ZRk5TZzn5Ivjik74dfxdAs5AeHyUCb+Uk
sHXstNyPL7W83NMLEhv44xkEXPXj9869+eP6NDi3ALsfA+zIa5cX6/8JY1xHekPl
Pus50cMaE4eOm/0coCdx7lNhVlNuQ8ehLiv8leS/FZA13Ngt/JVWVxL45UyWbBy9
XaPPIIi9B8BiUvqp0X38P++bNfDuXxPOd8VJNuNbN0N70irEcmuPCP7Ey+X6iF6T
7AhXcE1hxy9pZaFAusiruySH9NsHUdbMW0JSn7agvRapfgdnHhqCmBY+F9K/zSdB
vLJsIkZFCcyTKB5Ujx5gR4unPbHvrukgR+w3XncjoshzFMf7uuyv5rbODMuXXyl/
xNHjrl2GgA4/22VqZCW8hhTI7ih08Vgt04mcKcDYvgOuDqbP0RxpVXAa1cWjTCGO
XKXPP5G4EVLiMui3gcInA/ezZkOcQrEp9Dv2xFfmvLpLJD2oMotRhhqf4y1rJXSw
/NrEpd8v+KAFgrvlEiT2Vx19K/Yehxdhr/8ZJBDGDBti07L1SX5Veuh6B7Jy3b63
KF1kIu9fegM1miWr9AB4C1YSqvHriQSXExBguQqMLEn6x5WaHe8OUATGdlRQJqwa
SV8isHsb9ZHG8V33PIraQodkdaN0zJZ5b9VTGhww/mmVi689hJo5FVWJ7qu9v1im
FUHMRT242KHXfb31467OKy9kzSfO0uw1ow1e+kZAyyGn0H1aBxwWVF9gR9yhkt8n
y58wQIF4wbaDux6fHCxrRDpZgmyrxPTUbc2TK5HOaXVW2ALx6zmdcCuklzCg766d
E+CWLYQSZzlDu+fUKCox7mze7+g4L5Lpg+X2UHqVZKzpoucZVyymFi8/J9T4TM3Z
JeBsSyreQnDxYhSDQ3GPHtq+155/tuf7Pu3aPOw1DRSiZlpKo6bCLt341qTxb0a2
oSCUepxywfPIXMb6bfoAPaPiXbpBcRqd0j5HXZ83SVkcbmYV4Y9C2OOJbG1bVf6k
UyXn9ftmZfy35JRE2bF8ketPfQtIJTt2Vn0r6Au8YkpHqE85bbIn41qVRoOlC3R1
z0q1J31c6g/I/UzbEA8uc8Uvx2ZKhn6mA5rGwszOCJ6r6k2DMwdrDrlt4LHl7cfJ
JKFAJWs13vHtXxiaQzj1uuAwinAo3lzftAAwyXygDDPUgWJQjCi8QzB7s2EAVcRO
3LKp2N6J1z3FRTako0W5hKKXcCeh/r4tedawxO3Skb66E+t0mmzMUvmG1hj75BPG
fIPIwxhWLXYRfwWZ5tN5s+qExkxaJ/hIqFjM/PazEpgv/EYrCOLcIgYq4iAxokEV
pq309/SnHehRY1I6G4pFK9HKE9FuE7x06xeUxqonNVNotI57B/eaFkSS04LME2nQ
KUhxE2ya674oefulM3jWAUdgC/q523FgC5M3MuEnxgua4Jc968mVyWAiAoEuNFyI
8L9wfixiL6/+NHc8hp4fgfF9yRuvPC2avhmIrnqEsw33MsB+UshSboykp7l4WBk6
0KTjBHPqdXFQbQaW8Jy6OGP1YHHm5GvjVW19LD2DcVp4E8dMz/l/rrZroxxgMp2c
WPPucFUmsGPJpkctwDpF7df/5YNuWLTs0kjXM5v9HkfMEC4olzvaWPjg0F7SDscE
EX/9r63mWomIGM0nnvz60Esv8DtPjP46IfaSMFQH4zxmS8GT1bT5WwvhGNtklB06
b4U0kkhVRLA5KpAffk+e59hV0ZIrz9TeVK6q+ave/mvY2A1VbZhoHTUmzWBDT7UO
jhHn5swe23d3MRgOiAnu6AGqDATN8/LKHzuO0rM4TLo+DL5jN78e3zanE61c/hpQ
oMmuMwTaUyTVKqdiOHvSDEbXATKRV0XLOz+VzCb4rghAsqUlcI19KcmncL2g6NRT
tRZ5JSa/L+lvUQd9kQLDdEAcvgJJ9Ghm6113fKvrjVgJcoIHTYe/Xep9SK7Rm5M+
7zBky3bdNXcXy2DY6zIXP3P4ffX4tyua58gVuy2864TLwzYQkwCzzZ8V6ebOlKTz
IbPg6vDmV6+vF0AyxaZxtzfrKj+kV9Iynn0VNTx9A9Jpeh80I88zzg2orjjK7LLE
juBgvuAGD+BhZF9angNHrn9wQ0S1UMei/y+WgkZPTmvxy1SkNoJXBhx9wpKY6JB8
2uzuOB+q8B7NbWAKopvqppCqiVTkhohCKkGbQ15WmXxjO3+soaw7nvixHlgUiwyY
v1d2mAcZ3ofgfIogWjF6u0SNjJVzgw7i1UZ13+wOSERs8MOm/JmWr53raiQbo6dN
UG5I7SgKkTqtxSZV9dx/QH260OMgGiG5NoaD//obB5nJ6Usa5M5KkHkjBq/1SI+W
0HvMkm44rVunr2L/URlu8Zbt0Xk+IqidLUekK7cePjVzQbwl6MpAjSCFoLExV4QG
wOy4RYul8OvNk9S09svuTs2ihjDuJAH7p/efGKnnTJTKxJSrz9noAmwy0V/MuFwX
u9aMD2bwrokfwZw/hLBULR1W5uuCKgVdpgk3Mc3GjR9vO35YSqcpwg67yQZGrSNr
8aYFLQgIs9QGpRs5zh7T13oMUzCRzwjmJ92Bq0PSm6miQNJk9mGDeCtpIlQtdd96
cIxmoiPFiPbfA/jTeQ0Jg9Zd7ujQ2koeWERaAS+rfKhrVTB3zWU2NQOjkoqKWh8Y
f7IGoMdNFRm9g6OMrtg5K2jevvAbyBSt63i11DkVV2IJBmEDPn0W2SwUHnYCdUmK
H28GvUG82DZ+3zAaE3msyf0KqeE6RZg0zAR981lWF21BtTAfLkebaS7F8FvHHkqv
27n2/wr3ZY9wegyyqQbhVvmzZPbFEtdvDjPhS6LTGiASczNYBcK+lMwvudkPWLrd
54AtSU5Hpet904qZQBZwWlKpSnrqe1C9JgRE5tpvEquHNr9L/4cu110GThd1SnNi
CAVjI+kwR/SvWGCrapEkEYFC5WsuyXDZEMHlqyRAirdw5R7bNw7JB0/o2pvbFhH8
MEu+LjniZWRJ5TcQprVUfBh20bEq56XwRrCibDYJFJzwv6Wo1oB9DnNwbPX62MRd
f5HJe+zwrFR6odMMBh8lEnwzusCV4mig2AyJ0iOW4YRoWgjSY1+VOf8JpZ3vbjMl
dUy9wTxP8mlUwKm8Twy3QMO0z8M0CwH59ewyXCSnKsJ42sOcuiupzOoiWGPHi1CU
WHxUAQYj53P6VEAVmrc3+gSy35Tzl1v431LcTFewkpe+fSQjHiImqw4tl3Vsa1+5
hUt3fkEfZeKrNFbEveg4IenreQbumvGhb5nwc8xfx7OktWwU12NR2Eo9dv3XUFGW
g8oz84RvQrNOS5otjpLUNiBhqqRJDit00KCUGVXxmP5AP4olCuxIAev0gyReFmPn
xdFA9eaUj+KpPyswWBe9rDXu8TWzjeqtA0zLXbGDYE8dRz90k7ZxN9b1AUaFmQNe
44mcKRO1Tzl5RDm36coRWCJqtHu94f+z+4c85PCx6myLtIk+bx49d/CUQPLZH223
hJRGdTdcsfwaT/lRZkmBzU0p1E2IzzVwFEG/27HOaW7TfM7JoUJVZYocn6cRhzAH
5kbxoURzO3tyefa1SVtfeOeR4iwI/36Y5esMQvSz5OZFydiGFDI9SmIiGD2Ogr2V
pla01dDwaNxRNG3/y1WNMQePzzMdaPgiCKZgBYZppBPlV4NuZvpWgOOu3C01oz+B
v4C9qYAHy1ztkCwZTPNc5H5mp4i4UEbrqOkuPKGrEdrNyg295gCieDknS3IJLDvh
IUo4+1kX5DuplDNUL3LmGvVVbbISnkEp2Vy+1MIh4+FPWFLX9KV+4vxQx1bQ6XKb
pr1o2952mERXTOr4lRmGO3pk55Lmqsw9hw5MMwcw7/+eWt5oOWfeij11TcL6zLJj
lMOc/HFBDheQFHiXBzu2vXpO0nuz3s/K0QcSUio6m7bc6djCoNeQG4+xpJQNNgtX
IaakBcW/5JXW55RalNVU9BF1gJHgFM5XU9DHkFFfHkWR06gfncw8QwJNh2lipxcX
J9ycKYfFyS3fDG9knTke6xnfLG05S3ARLJhKywYIif+eB+NPKoG2srOJwEJDXBAB
sOmEe8xOQ0ZAq+6H9d7/ALpQqv7pDRe0YKoX25e8YUFE7nWudrydMKPRXj40mPWd
3z0+0T/E+VNKe61NRJ1lECYi9kgAYHKog4bbvSCQ2bhaCWjMaMHHg996IzOMU0G4
WTB7GvAq+IjkVSmOdAp1wWrNAZnYlkMXqOICaKiF/eRyo5NhHcgTa37LteYXW2dK
INN9ioMYraS4c+ScVlr+fnyB0w5TjScH/U8tO5KaKjU76ffjF+BDzRGkEsthLuo0
zB9iLESHAIBiNKDC5oVjhMGmoKcAnjWajUW7YpnbXQYxQBf9O0ORf4Y6lGS8tpsD
79O8b7L8knlU1dEEXNZ5GpuglPxq4m8Lk+pXjFysVRVN8KSBeGJ/eOlpK2RQ9U6U
ti265IVOai9Nvz3udJ9BuK2ws2uxDCGi72ehCQCq0mvNNfj9Bs6DCCNNqfXItR/P
7oIAaGW9jkgzuSRmu8oMs3iGuPjUW9XDml8t2H8ibjDKE3to1focUHimUu+WQ/fJ
Fk3wzdLr4b2D+radbYj6A/tElCitBWa4fr4v3iuWKvI6kJb5mEgj8DEVWfrknB9h
tZA/fLohkUkxDnhyPqN1duHbtcrod2nJPOTzS0TU47dF0gNFsOjUUy1+MSWAczcb
NxwfxYGpSHC3HgXEL4633qxm2lIuvLQYgaet+VWeWeFsxhKfGGqEaUfUomI1V8AP
zID7hsx7KuCMzKnxmWwQxfw+Cxd3QDQsahTd2UHs8GiVRwiaRgzqRj+QkIxWiEKW
E4JM0NVVulU36sfiQWT7Dd/Kb1HkwYq7HW0o55ePt/59vZXIrufcKQfjeSpCBVVJ
j4YY6IAICXWlUvTfM3UzvKHsBdK+lho+wnVdH9bS8M6gZ796a80rM5XUEUBhMNmo
EywmJ3wOmxtvx+NPFdesLzW18qLSsU7duKe5S7qAJmNW8yXP54Sx3I8Y4vJbpT+7
OdGQNFqJaBpclO8sQ+khSjeQ8AQ5mczasDl0vbakL28WzHVUv+FsfqHl4IR5q0ER
M6ddiA3unMjl6AKTKcY654oLS4D0Sv8bN78VOvvtXFYANxP6aD49f7layFhXgoRt
/RYEyiaFypR0nDjMNs64DTkKklKpvq128i+z6XemC2/gA3ygmn+LFmNjG12ufzif
qkH006IFqxA1hiL0uTP0Aivf3TBgYplRRKM2wWKpn+I6LvZrS8RcfCZzZa8EQ+e3
WURuV80QLYtot94cnNpQuPTTVWnTfP1w77d31I6XQdptyGbOR09VDZ8LzB8XgtbM
mTDAeBoCj4b9MgCcZC88IxIMVyQUnR8alJTIztfaaaUhOfl/3fnar2FhQEpOYQVX
7Bi461SRFTbtc80WcDxFl0q6HKzVOTCd2cD/UvJO4ZmJHqbbriTH68eQJPPRCD/L
0AM19hbMqeVkqQ7YfbKr6kuJAHg0PzxaveLvUs2tt6N79At9CqbSSwoouBgexN9+
nL9AWXkMMjcJWQJPu8CCPoYil7iNg+P4gdTJEbqKgQVfywQWlHSP4sJWLnmcPpZ2
ktXZDDBciSJO8X25Y6+eXsQKvWP/jqUrL7uCWZY5zK92eiNPeIs8rmnPh/prR3VU
fD19vISX/tAClcp7+/szjtZB9/7fb1MBxitf7RRJUtm6hW1uELWpsVFtGzrfgSP3
zGir+8uj6Gxli7dT7Yvtr+GzFD3cutF8Ztd7CInV7PG1RdbeaKpNftuVLrIsCQzd
DNEdkRfDpYXYvg+fc9nFaDxKvbN4565rHzfvvq+ItWKeFxU0vLfX3X62rcrTfz4i
nCORq4pXr6iaEKoYb/A+xi6txyPy+S8OUCDE9QSBYwBdihvPQZGku7XLTO9h/miC
OkgOix50zAlyWO+tKPl3R/ucuZxSaa51DG4MqhLcyhl2fj/wnKmfFBzHRJoS+55D
hvoFrJNTCAeZuhDRifoSO9fQZudIMJuU4PveL+vhpak6FQHTSnWXhoRhYBLnBzDz
x4oxPyWPh7h97RWCz8hozl5eHk2l3O5vzU2z4Czy2S/oydzZa6aeG79k2+5tJqkz
148Rz86ivKcVXYTppDloFZg4ZRNEBARQYjh1JAG0vkpKiLTYqsVGZB2lv5MNTvdX
1IjX/gVJQSb9YP/jfOyZFpBl701PvIB/EDCYZkiVMknDeowonOhXQmbFDGfZtI/p
oia46q+ZcOu/tg53N7w/61EQmGEqWNIMO9lKvK0ZLYBGRA89U9wvb0OytkB7ijw7
zQaJhPZf93O6hKffiiqDk6sryh/EQzHZRQNTLTGu8NVq9WQMcjWtjzBbgoXH75zd
oRkTRlyIZYZveDs0Iq4ErzLtbTz5eZwnUQVhNEFMIkT/nZrZrz6UhBi7D1xr+fyP
2JC6J1bp3867MHGK7QUnDMN8WQ36EtF8aqUtFFUan/71AushClftB2POHFpjvU5i
x93bteh148nZbnglGlKMcsWJUeNjh3XMnDO8oU6eA/7C3jQiExNZhTiQCXr8V0zl
20OwVdOq87AZhZQFn8woU+4PYlDOmo8BDDiFTJnCcWhSHBrhip+kN42udRnABarP
oNDktmULBVrXpsd8omIbtGn+zoHj59eNbi8LRzEBuVU4JJtZs0t1QkS1HdCiSCTD
eC4rmQ6Hr3MwHsP52rZnOFSjUnXFjMcg4nM7W1WKSw/jRukiYHG/ate3+Gi1leys
EPxB0OBiKtnRC8xCoYG7sGwA7di3+QoJtn+Dciik1zXO54m/PJmgj9NQsijKh2Y7
fsq8r0xwX3oAyPp8aRhkz68hX45XINQP8EkE7OLtkAbOvRcuE2IwPWVfXu/JRxJt
IVjmSwWZdh3KhUrnD6xMRYt/3aQt3prWEZJfx2p9D9AGOrJxZiEepitEKe4EWd70
6Tb0tICA97MByD9G0CjH3JRgPjzXv3xdqewMTQo1KhQj0vYlsbclcLU7vvf6kdFr
xGRl7EFZbKdIU77LvY1wJhdI4PszMVpJlp7gnaxTBU6MnXygt/Fb/c+6XNcYsF/r
u5g+NlwdAduIk2tzbKXMhng+TkSbmR3Ic9S55hDODlbapQ4M0FDaERHodQO+RiTo
AJf7MdiHERLQr3/+6xWIKUJCu4c1WAATvcMsiq2ZAWqr3IXcGeT90sqEDCnW7kAD
ITFvP1HYYctoeaBH1hSZpzMFvztoKWsjNuJBdKROVjLFSsG9vwX1jab8EPob/t53
j4YQOo0GjiZGrkLFfABw7vezFlPgh5FCkiV/gNyn/qgPrMjI2bzxaQ40LCv3KJ3v
+iHtONF6cHkGfhKQE1Ru20t70n+WsYo9RqmR/FOyuiF14jOyzhi6fOyCwj4UY6Fk
POQPTN/+lICGF/CWzredo48HJ9dT3WaOIvYcJSvHCFT2m4XnRETrt0ufteHbMmvy
RVZ8HC9IGBAchamNdAXB/t++cJ7xo+14o1EgYJUmdbYnzIGQoV5EDelTnqkVGNG9
/cgJfW6uE2+NBuLgSr4z8PBDALUtoJ8Rr9lCa1Z4YRFd2nxsNAhUISug33A2aV2O
VKLovIeGN/ODej2rmtIcfZXnDd+tlcXAY9nGjprvrNY4vwZg82rHgGqXEbD5vlBN
e3QRop/EK9JATctJS5tqKROb5Rg+GBntCEQmw01YOH+c/FlYz8ezSqSqaYb1cfLP
hh9l0qvqohamsZGmMYCExHRde4Rg0TZwTPyFwGIBqdH8o/t9UYlDLuULP25Wasto
FMjFU499kzhwS2fTL56c2sQOkPQMViRtnFPJbuZi6ZTnFFD7HUzm71yhuzdVA35Z
7ehswvNalI/e6EhU4qHCao8tZEgN1ViksjQXc1RkITxhNhfYQTZq0Oe3QSvjTDLf
YfRXA80xP/GtASnA89nQb0sCeIIPYeRbQixg2VLAf1jPwcXr9BI4bwMNOnQZt/UR
GriQPoGIlgin/SBiYtAyW1QoDY25/ZuPuNCRGcV4olt7BG275gUUH7jFlNXUOOqI
B50iByWUCV+N1vUOODIvZzEXr7Zjq2flyeSTEvNlqpMQ8HjySsi++s4dnte/BOfi
JIxqV4/0LnqyeRKz2aeUNBvH/SIvFxwYtQecl5jPq3FRZZMNLbpdCbqlG2NeUWra
jwR7JHk4tUiwkah54Bp1WKayQ6rx4Cw8QnCZzVxqa2MUVQ/E7b/hck0f3Bj2r/vm
XMI+w5zJ/XNlZsHjcThUz0kc5Z16g6ckR5YYNYytuNVUKYBaOERYl2Y933izyYXP
+p4I3KEpYebNVR/UYy+pUy5aGuUp50eibqlMVGPtIcj0WWb6fw+ZpXkTnbH+27z8
nqObAcfUqnL2cRsSAWwtAryWTZLD4cR11Fgq3hdpuLN59tyzP2JIF/hiYq3q8aZ7
SJjSuJUKPrS8WOZ6OPb4EXZ+pmlq+SvC/a4cuRqsrJPT6l+kfBCfaMgPCs9SkeKd
FGJbmE/OiY83rtF/0bEqD2RYqf9WokXHf1q7+4/CL0AgbEFS7D1MgdiY1YqqokNa
86z31aSmiFG4P3SqxAJCRJk7Urd72Ph9EQnnBWMWSMFBDVLrZsqyoRWoxVcRX8ZB
6zk1g2Cetl1dsDe4FDibWMNz4HFjKj4Ah6HPhLIb4O+wo3NW+QOzgEYAiwkqcXXk
2mXP29kGTElAoHYNVT+bzJCL+GO+TnIaLCp9L1Z3uOYEQPDwVgjU6F407KWvfVoq
iypT/aNqtRP4cU1c7+9JYNdi5MO2fCFmDnXYL53tDcuq1riW4+Db5G30Bkhqupt2
f9maF609PjC+nczgeA90Sjn7H39jwV+hOKHYKVBzdEL4ROmVI/4+a7WgYjuav0Cy
tD0glZrb8LinXGPsHT5PhvZlm41/5Yk8jL1hVmVzrG27ol4bE3i5cciAWQG/5roy
R65KXEE/RyHpkCekuSmELNpKH+UciSes5AwjFnAAovv7e/TEQ0Mo08O4hLy9Q1T2
JDHqS/oCHn8wCdQEVc4h+Gj21y+S77BLXwYDZlA6ruf/Vc/q99GmsvobTUVjln1p
pObIil17+siF8kBYeJP4LfCC37HChokunERiL/nFqZ65IGVXwxWwUghSQQEjBzZY
chXWyPAVSDTuugzc2KQPK4cdvQM9R4rzedk74SD/mYXs3NE5Gx7CjYpNk9XO1TEa
qf5Gy1XZuLKYslr2zgxUW8+kbj2zVHxwEpOoHtfEvUx+7MLO7msOG1TUGnZnEGOH
w6mvKA2LcNplR64N+So8glYSm193zxSzs/r11nznJKxy7fvB9pIDiECIi3X4AlFP
SEI7TYFs+kz0Upt9cj+eV+r7JbXWeUPuubiDuuAxCWt3qxSJFyKeRZmlZYu17MEq
wkhHIvxGsBlCZwSJrHUdmR+1ewdjxuutvEq+rDzVJ2BUTk/ntI3wJzMU/7ZUso+C
VzzZyIxjOmOC3wPdXAHfF6or//S6Z0DrnsyLb7PeoiXuj3OuMLcgPH/nw3LcMwSR
vbV+qf96GaT7r7i/fB1iSgX+xKOwH7036rj+w3JNxVd19Cg80oWnoJo02vjrNbIE
eD0vTYoM3YH7m6r5drpsb4Gh3XdpaMw3dk3Qllfc8ZBIsBpTSH2HGa4SU5vUTa9w
JjRx7jZ5TmwOmyxofOiulGorP1u5I1xOJOlwebA2T7PyMj8ZYT84CUIaMnKWb2zb
X5xXz3AjOBffYtcGSGdq6h0KSl3dMnSJ7tkWqWlutVBFLkAUmbdNzN58Y/n+kpeU
M86M3zEQhXJDadRPFzp3WUhIt7n4ZOUX+st1fn/9urG9UdGpezd/6jpBYSDeuUHY
oYdZYc+YYs73VzD1WzVbpMAVPljzQaD/asX354XeT0KDhZJGZWPmisnVc0EhF4Dd
6W5zKgjLpqFKn4aDX7mIjRCs/YRgcs1x1ANTEwu6EBjicrx18Mf+zvFhqv6Yz1Tk
WA8FGRNUqYS66gCyR34RfeGxiiArWbCytB6VN+C9qJUvot6AKL33u2gYSuvDpVr0
/4Jj4hTxQ/7UgDrnQF25lO5MllBRs2ga4mgjBb+3a4SiMoVD/hCbOYEMuYl2Tl1p
9Ek/SJBWmIbCHLEpB+5yFCxhaVucuPs1uRcoamsVNWKm/nvjT5qtP99UQTVWG29o
HUMWfU4Nf1mUvUGrxRE6pmIBFFeB2pQHZwX5b8eZ4BfDN2qelUwQPdCM5UvOR9/Y
jbcEfhammkpp7Ar2K/vaKX+b5KRFkApIq38KyIZboilPbGCp1BletfC21+1mA+xj
NdBJ3KoZFcJVX15IfvqaE9wFNyXVi/p6CIeGLpZsHSQVEaGbJmMl5hujOnV4okoo
eJhdhWAgxQKctLS8jYA3Bj7Inf7bBQp6GZNOpD80I2Ij1IZCgyXZSBzYtyl9XKRs
adrHSZfdNZiW+8vd5Ll2MXHbpw2vW6o2ak9TNvYGSKD87WyfE1Wdmxre1Tks+4lr
d0X0a9kPe/k1T785eaEyhH/3M4sYMpPmMYHfLRQd+IUkq4XHMA0exHXdFU9uixwv
Y4hnynjSwu9a6D06pmA+Hab/Apu8uWn8tY5Z4J5OtKnS3rWm/bIwKl9po95jUqLD
WaAiwQ0CTlwcjFYnmcwGso2PSbKKhmxdkUbg+bZBHjyukesl9HwJ0nRH99yAOoU3
Ld5D2cRzbhGd6JBkpLqZAXiJOo4Vnzddy99lcKfH57GZQubinbzSYDZ+B5hq9sbU
ts8/pCHLvYsQEM+UJlHv0GN97hRMOZh51BIbS7uZZqRfeOWYgy79Bra1VMcUO/d1
tpSJDruu7XeyP8CKovYR+Dr7mU54bH3/jn4f2yT5TABuCJXbiPk27tQJw8cP3v0e
JKgOt9kU48EtZFkuHmYe7VLbjsTKr2WhnCgxNt+ghd/sp/ulHow0jhbDIB2ZxOq0
cl4QNKlkL3TYDMrp9SDSvGF4+X/nko90NiD73InRztINBEQ5EmLxl1ZOCE0qLM1L
BUat8PYLbDHPkb5jNyIB7xKnokOggFx4d/uKwTD24Z0TdIvc5zshfx5GrpwrInT5
t+1eRL1lDgSl138o50jH3WcWS2ntXGsIQIusf0AlZ6c3Q2w5sV+ktcMcwNP7hgaG
05lvd0jP4GtR0NQdTXToE/0cRQwnd2PGev0rVhoX3NXF25FlpQh2jsJY90Dm60fs
Ho8Ra0fILNTeWEno0HKeQ5j9PFg1SiA69Y570ClVRmQG/nEz7ly/G9AEFFy111+C
hPbhLfGJ8bnJJm0dsvXEjlKdZx8qJoBZnm95SGnF2iaRjMR7rzQ0BdOrkedhgBg3
KWdYEdTehMa7WByHBT56QMDmqEH6Dhin3azuy7hQH/i76CGPJ8ryo550cc/ee7/E
0ti2ih6NASq7UWF8+aUAost77CbsYceCLzauvo2UPDRRwh2OCJ6fVqQ2EjbW7Skd
6FdpYZTEKgyl11fdCOIJl0iJV1hZRxWLDI7TW8WyFY4/0hr3odcDQ6Hu/I13LhqQ
TSPd+FURhD1w7EL7SE/eviZx2HCVmAFXU2rVSzfp0QYzPxyTTnkbcyyd62MIHUw0
4SLPDY1f8KJ9GIKdtNsHHRzIrsiz9lcPUXhkz+nm6eW6l3FFVeGPEVA9OGiPgqAi
hytldLsWxwGof/Dsp4Cdh3nPhZ78Sq0fzqx/Vt2jp5rPAXHtApDiwHMw18ZsipJC
XVkOWDstYEPjnBfiLaG1KRM9Wf9IGjYMxUDG7rhXPFfLXZLYgsa8c4ZYfuuJW2Nb
mdcSZUyau42Z6f5JLpgzpF1gI+S7txcRVyAXGZ2cQbSMEKJDrD2UzLD19A/KrQBN
qcS1daZ880jqyuMuh38Sf5faJ3RBm62+udR6OdyvHw+3Qx2qgjbPHrGLLjBhQkaN
UYay09PNWcVxahZhybYIe+/pxlODCEbFBrgX5Vb8wS38DPsqXjPzuaFN5ijXlzDq
0082wqbQSmcvTVtwaAzHT4MOuUtLam0wMzAtLr/HTNdxmBZ6fHGfx0BSeOBpfm4K
4HBaTIKpyXnPRmRYdF/u0uvRYnW4OwNVZfuTrnQw15Ua9o8eehga5slPpEOX9sgi
8igB3KhQDk5xjffmApBDFYED93XEy8cQjpugvMc29tkBsdK3/C8nrhvunX7xdiP3
eXU8t2Uji1i7s3KAkSBqUydvGC1pA+ZKrWrZbHuhS+Wug9TJ8c5z2fT3hzrYvtjC
1HFbcSQF2JEO7gFQKS4ercRHki3vdWZTNGWG8gX/f8OHTfQFNtb0yAkVkZrU1ReM
S0u5biHudu22Q82G7jI+WSpTkN5M3U/3Xw9FOkLBqj89LdSK5utwsiMeadIhkuls
XKpGVP6H1I9rA1AaZWz0ukhhghwJJUsQGYM4E5/xwpa596LHqUdsKBSAJfJ3qjKX
YbKyKC4PCJRf9zOHahqB7w/2/1Wjy3IwscFw4yq0683usJvfMlsbAz/ogepSw9V+
PcMAOcNbFEzWDgkD7RzFH8WiNoQQzrqWVuSU/SWBUWEoejGZCh6CqD/+vyeyOtOr
eBeeHyzaVy13H/uxqetNokQzfxlYk600Y/0U8y03VWP6vZvEpJ10FDBnfEMj5ucn
Ro3l9jtMr22WOCXUEAFaScI53mt4P6+UzE7vA4mFw7MDyFOZWaepjRCwW7UPeCjJ
pPKiEFLF7apwvwLFfYDYUgl/yq77s4wzkzh7w+yCwHNzfLUb9djXj3PnWGVx7KEm
r2QT7h7GVI2/y48r+pCP1gtmCvivnKk3q9bo47drC61/XSr1bRee65DrxZRdg9Kc
DE1br+1naFoUyIutsoFdI/Og8n5FU6+DqnU9U6JkBB2IX+PeNmuaJphryEyNCs1K
i2zRI3Q9eTFS7MyKjsHF1xh+R3Qsh+lIHIcOHYf5cOMiSwHZF9WFj9mAIXUodMuV
h3Sb9yCvXFmI9mMc+gJ79fGqbtYmcXAIpAAMGiOBgLkEU9fq76wsoME+WMysQolm
Wzh02htjwgnsESgrHZK5RWxf+C20oFDVZyc1hSotOX7/2tem7Gyp1ytm0HgZUL97
b7llHn8myldRJTSFkI6bvoDdF2jiJKRIstbisVVBrO/o6SBUYMtwjDqX4gJ0lp5k
e0E3/moMcxIqB8F/9cSjuldZykSd1s43JGnPjBdHQ+PdgnwPtClL+u/9fyiftHia
zmnJNfw23UPlQPJkzOejKZAeed/UY9e3zq6cT2xTb1aq0+X0buI82EFzhonNapak
H28W/2U6eYnnmLfXS8sI4wPt4K1VVckqHv7bL8D0paTrB9B1Va0ljd6vcV3/PcMD
328miMdZWnZIkKuzJir19+TJG+FkakyHa9LM6y3S93kWr4atl5f+ojCMH//0MHWO
HkfX9hawDRMlECIlgUmROfWCqPRtPV3Z5zVwWDWIbVH0VnlzCm2RzEs2Zm7edQnT
dOKF6SP1f+GckBA3LMLyrkoO1IBDe9wifIVvM8K87qekmLccQj/TQkDpHuPSdXo+
7wOxvPTDrF2dGmqfqa0S35Web4ZTwXojPqjO/L5y7ksV9eTg86SXUQRWd1xUELRk
8ZR/5lapQ+dlIIdtxnKnyGysclk69vohFzWnMeo3ZOu+T50siMI44e0jPEUUnKqs
BvtKMqRxLRiNASBuhQhs+9isMn2UAWQ0RgXD1XdUWUyaaTOJcS3jYnQy8av5NFmI
mCvAS8JUL5Az+p4I0DuVy4Rq4s4zieh9YTfWg2CY4CZ6Wb3lczCgwZppCIZWQsYW
1eMt7VDfMtP94Puu0uxoupDt8JFMXveT4MD4t6i2FCMZxyJVojjRiZ8HrllZoyyf
PahOwRChGrkQYinWyupAM8k5IAuyF/pCKNds1niUoHm8gpdJc8ll04tDu9GbFTrt
kUlW2c8ObI57tgEr008UsiSPrnPcoi9UnVDldah6nnN4878ryM14zi3Igt35+O2g
8aQAyHcc/ayXU3B+D7c0hk4CKVdWYZmrzQqMM6sjuVKcxFLhutqKo5iGrktwfq1M
eZtLG40mZw3ND2F8iHFhQQ/yfE4p2kiuJy9mZyOhEXw3ieufoieBkZwCoOJ6yr6H
V/5qHAvFlWm8ySxyb8/6ceD4x7PIBmpqZGLR2tOUn0bM5JmB56z9vwg08TxS3l1f
J1nd73YyyS/IjdEFZgKNRx9BFC2yOjSB6LoM7YznqCSshWab43cTJRqTHYDIc1qL
zPg8JXhKcnqRAl1jleGEvDk2tTdlZRh+x8taDP6ta4svygZbWztLkkOtvHzs3vzE
TW0pxJcHFza6+9ggaJJAtnKZ3vrJnli9KmGozJfP3E/R7/jbR9RAbi3+OWqBsJdx
yAkQSNicDKg9ZV6XsoT3KfBQbAThqOeS4Dq2op5CkBYXuey02ixbNflk8Om8ArRK
mi20pcjLyVszFiCkd0EfPpv4gY9nO+iwl6MU7BE123BKqSnkIfogqMdieEy56S6O
2t0ZKjD0mXPjMaBvhYPC443rq+c3HFkM1KYflkyVelTPkd3A76zFxJ9xapFCR981
McfvSbGZL+Rwq6Vk98gpq7gc9RIcKlG+nJnPjcdCq+fHTW+8WPm1oKN1gaf537Zf
pNdeDG8/DTa7aCq4e69QmXIXaeD/1qHphV9ObzIxvc1v9xHobKqF8WOpIgCuBWOq
GwTtSAO9KU/BNqIE0pVDnrWogvWBtTMmvgGismgTWDKA2h3m7WEVxximBk/+7js9
KmRsFwBrSqAieu8JzpT6ELF/7x39mMS+nejXd53FKGIne8JAD+/gnaTMWNoKcuXn
0CNbX53+wFiE8fWfafQ46dFwIkTlL7oyPGPFZ0lfqAjzg04HEwDL3BMHTWZsu4pf
pnBCilI2BDI1nmrKmZ8T1NKzPRewbzLnzx66+U1WPu1YY29Tdp3wVLvUx7xe6vYT
JukIcqfxfSBymMP+hsjX3Kr5oAQAYj7sZyXUroqLnzXEmM5nevr0z2T7O6nndgK6
+gts7lW6LuUID7GOQ8O8/jLJKXae8G6/9QAj/H3IWyP4xalV/kEgzml3nMYsHc+R
QwQcCQ11skg2yjR2UEmSH0TmBSg6bfSJs5ElyBO6tGB7mFoOo+79NYCkHLBViq0Y
mqHCEn9qoiFwGeWPKXHPpb5At6V5PNOooGIAzXqpdaS8AWjZgaZBFNvEGjBERSn2
37ZytnC7eXvopwH/FiDMb5eM6vwfC3FpZ1NnS9nI03I/OX/X7A0prA0a/JBOmfvI
d/AI3sPJ4rRBmYQcyMZDQ6VaGVOn+tODBLFztfu/jDTfSxI3Fo82Gvv7cHoHv01u
I9dBjfu0X4V4PmruXZwJAkbObRaeFm9A/NAOuekdOwG+NYnCMlfPhIVStxm8Ltwl
PJs4DB62ETsGyMSNBTPARWxNlFg1k6lo7aJiiKfBScRVp4oLkGxqYgiSA+ND9dKg
Jlilri8W7c3k0v6eRpBGfHSGCaUMD+/w3SSNh9fJXv2YDw3WJCYqOq/8MmGwdm/Y
XHMnbw5vm/LgL5mJTDqreYziS06og+MIGlIG6mVe82UDFQtuE3/To6dufo5i/WQn
Sp4bIpqHGSsDFMqfUW16WW7rjkbnNT9Dc4Hb0hEJtjPIfNswjysF6SGUG9ikXhR/
bCcGW09YvhZwm+o5437MqGiR85Av4B5VaB7r3ZYgI4Mgkqkhp3j+RwXckb7bKpCw
qsTjjPgTN8/svbtapNNCjywcPsDdLg7q3FMHrljOmABS+NwjUehSi3bMzKRkmUm7
Z6QFIPFSXSVTQgNGAmwo6oXSWUYKLeQyyal2bxi4IUBAhgo6E8YxxzBXOp0zR9o8
n54uMeI0YkxNupmKxzc+RSn7JjGpi35LKp8x5McI5uzzMXJE8ca2kzow9PtpEAjO
vGbJCZB3F65A5AkTb/dreIwEBDpRqpP6IBoCekBN3nZVhuUeSw8f9qbh0UfBTt7t
5VtAp1YQvec9Rm1T+B7AByIeyiLltRdLEPsdWslXoH7JK3aamYo5UgSSylHeSRnU
qYEnyH52n2DKRlbyRk9gH5ppgPEyhKP/eoK228xpGAApYQAA7O9uEfzUSOUrtK06
KNsQbPBtma0O4HaXdZXecz43BT7PfwMzJTC13xQLomSnnsbEdHZY/ZsZuYRu6L0w
+cNrbNJO6B/MzzccvJyZyYeK+O1XwzZm85X0scL6B5QoukChWkA5RzfWhLFZsnwP
yFJPAb8x1oh4xG8dZ7HrfvRjWNyl5hD2gyJ1ssBMNKceXGj7EWIhL0PPpcwmJP7z
BRrL4zRLh/0ALNQkFEnKTYtxFvYSXqceKRGaKtz8TU9XV+3sUQzmURUUcg/6dV9Y
JXc0ZthitA3NUjjbZJGjhRKgEmvI9Hs8PLEBsA6av7wXMUW1IjwEcH1du9cHvSMK
fizJD7xvub83lvgNieMS+3+rDVwW0IHqpM+ZUx/u0LpItdcxutJy3YeKB/FCmivS
aMGP5z67rmWtdbx9p1ieSUIrjA37B0sE57Ez7ZKalRE3Urn945RLdGSyavp2Hsn4
F6TdezosCA6PIvFgLfUUaMZKToEIM+zNc6I0E/mjsU6BeV6l0Q1XL1sdRw/ObS5u
DNkzepdfRTCnifB7+X69Rw5NEvmRoi99aT8FKpogK0pmIDEo5TvXB85kD7QlUW+H
gv5A/ZC28VZs7XUHeZ2BVaXd+/hdpZoGnKW6bgsWnTz9ZM4VCYhwyGsHpdtl12vh
NHf+cSLoOH9Sd2whmDj6qiCUWM2pw1scjgeSmltG4LIPzAFZmTVaVjz2SW8P1WlC
RSgDc1SZ2tjw2kUyVxnu90JWGr9twKrcNu3j4/mt4yqvBiCO83uuwwEpcetJoMFC
fVjKr85uoKql9MpbDckZxnwzsV1Avs8AXVsQPT0ohaS6ICCbSD1LQpux+YuEvNOM
iJW5w6ybbwv6iSW13uCG/RCXPWapZL9eJSNxYMwgp58Wo12nYEP7OOPiKOk4Frun
NQkp3MAIgi+fkIWCJUForkQgnD0C9z7czR8kx+CWo0ckmZP2pmBxndpifKeh67DB
T4GM//MR4aD9BrmgE+gOv0pjNplWvcvbRPAHdJVnOP90F7VvFfCbNrho1ZxEXXup
KA1HYmeOblXIRV8eXbvOlx5/wICqbNtK2ayO8JFD/x7/kYIWCl78YR/ErrwdzvGa
rFnEp3eVwvswxO38vTLepsrBwMYWXgQML3PfHYoCvcRjNw7DEZlzr886/u/SXfqd
YHDk1ccJx/ssT7Ofn/B2VC75EJ0ATcrVV0XIjk+fgaF7b/YTq2WKUimZLQP0iTzF
HQK20sE+bqx1pWZtc6WRT2V0TDezq4Y3bXdoXwchFdFWgmur+wxMl/uyN2ujDEMq
iiD8zankXp7aUu998VzkBulxnwDiw8Ct16Danc9ZBSg740WKLfVo9sSyZan7TBPs
HabEIQYJTvM1vN3FsH7WD1MXOeDGm9SHcGmVg/i+xrYGEUfhXT0A0bgpsArJ6iKd
mAqZYQzNZdXAY7Xkg508y5TuV4K2grg4JR72VB/6/VvfPnXg/AJ6BZ4B3dr99uYX
wplcsF66X49DlF30aFqG0fy2jcifsK4I7XWcWwfXYxoF/6mHePojmflP2AbNoD5m
m84UADl0abXPIKD3zUYwAAgQKeJPeDicOYH/H/cfBMmvTFwWb/4C6RF/u2y1c/AX
zDko6KMrmKMWGObFR8i53G5U5QtnD24y22rjo4gJjxeqMTT0xQ5URn0UMQGXZdQP
/XtYKKTQbm2dpty4goZkl4WU3JsRkgZsEIWgm0Z9G58arb1dMug834ANGeajHdKh
ObCIRXDDmnnr9SR5ycmeIncKtDOLmyn9mFapHQ9I5WFKX2UwaYv9Kh98HDLupk3C
HdrE4eFIUVXm8oyY+8IJQTr+6u0UR5GY3MlSHDrF2jJG0+x13C5v3JmuBEIbZIFh
L6EDBXKEoJFvOQfckhD5cAZYu70WseSBLvHGNT+CV1P/GNaTxJfFHcLP2+BQ2cuI
hAp7IuqAl5jBPOV6Swb4S73pg3sBRrpWRypPpA0oCw1ieE3dDCJuLaVR1Vo9dAfg
Axi4N0YkwZYzBOTXHLYBd4I3duNeC0GKdLrHJADoBqiVncvKqiBxWa5qlvQ764hN
pTTdZzWWwd3YfrU8OTKDFNO1P1slzlqjJpY2RwMCYVu08XKpGMQOKHg5oMtQVq4u
jAT5poj1n36GoZVnX7ytU1CWd85+4phHuLB4P23tUCx+XQo9950mcX4WpwxWHjx6
maTiWPFyYiKjPsnRcSjirMae7kYXs+0ZmwgBG5QnpncrAE98fB6YiJLufBBl0NKn
AnxxqKta1UuD4HjlAxunBH6nZgr4Le7r+4VS1+uHrSQL2/QzSx18gkjx/cujSM8M
rCdILzi6m3DF6tG5rpTZVhmSHrJMP4iKGpDtVnkMNeVx0Ie4rLWDwvXMNAqvBcdj
QByZrt0yy1+B6LXRcSUVlgzwTlLPWzYibRmSXDaQ9DfGtEsYcVegz6stVwe/jlzF
iYe/zG2dfkO7+wj29KOVsSao3L2n359AR61raK/vI231bT4BsyoZuYt3dSxtPO7m
JwoQYQ8WA07Ilfqc+qMk8HkrwkzvFf6MOjQ6RmJtwsEgnTVSlxYJI4REW86hjR2Y
uUkU7BMAMT2iLHWATYp4ggPNTcnletfq5k+F5u8OCIvhue/Twx5up4+yZu4z5+oi
rbrTthRfHM8uILlLVweM5yyj9oID2su6PEIbvX0u8Wv1mS4fQr4W3aWDE0MfTv5h
sJGWZv99ltVkocA6JkO1sGREHt5/OE1OR14Zk9MxsVtxiyp+r+O6P/HJ6241SMQs
zIHOC2ns0YCoBJVkfyKDPqKVyNbd8pwGEZmL1oQz8J/WQpauGJjdJhu6LUOPvVSS
GZML+zM269ZyYLpdexnNhkcU5JktWRzIcdcOt+137toop7MXP3g0D698JvWaNiiJ
DKm8Z3ZU5Cfh+6ejq7D+1Dh33tqvoEomnZFQy54Cg/2OIkxZDdqkD/bACgIz1M0z
3VgP1kk+nktRZLqPJrlYctO97Gn7XLonAR+bLhhxCVjhgcNCbrodf02YUy8BRkMG
WivqvG2aHryJ/I5G87TtPvRBgQPCvpBNEhB4YilSasvOZenb+ZRKh2BrJx7vl8H3
1avlJJNUtAc70J5f6k1+mD/SD4FizpWuIuDHnVWrCJQ1cM3HjvAAoskDkB5ObhFo
s33hDS8nCWcJs3yRYRaIaTHmi3yZmAAXShma2Qmegra5cwh3aV3fqh88BCmzGspG
aGL1hwVT1NDR+19LKmL8HJMxrSizvgdPyj32vTPwhE151qna5ZbyG06qrTUMnNVG
0PguXhYvajLHiYAI2WqwwzEABSrFpt1Iq23h0oCJDhzsHDVx1k2U1wgQQAoaIi+1
cV0Exd15CH7O8eq4AdkuIyVCQfeROyMq5vpzkqeL94X/1hCdaalFgHjyiqR42YYY
2FjZ78PBlQbyc0L6uMj8tKri6Nf3w/uA9AsPNQNzAUE3BVW1PdtK+OEySrjQUaL2
Ns1U3HoU9I9wj5Ul77rjOugJyXzUs1oGezPB7v1ov+nVIuOowJajjcZOWiNf8wlH
6RfXVqbNMb6ndX8JRKcvxEPWy270QnVrOVPBBCH2BaGsvOjhrbPaho1rqp0l7wvv
d8bFoHJP9cNQ0+ZGOigyt9yJqNJvNkmzo21scCsE6NmXLrcgCX0omY2zy2/VkPSk
RLtXgmCmAqOyRXz/tNy715gL1KKpZ4rtHesdyDCddBIQMy/WYQCHlM/x+fKFjIFT
zTOSGh+WcnDGQrgX8k8EzPOuKx1XDSKrwOVVsFwFg75kox9/g+bfx3nBGCFHLdGH
XyYWh4FS17H8WUs8MUXeJ+VdRQt/M8v2M4cd3f32sOK1OV2XvccaHTxolA7yVoED
z5Ls57rtu5fQa3cm+IeBiBoIUhNmrvJ0Q+yfLLwWu/wMDaNr6RJkXxAGLEREw9B7
wvMG3kjx9mIQpzMPfBEFV+/m+e5ApqNGTwdUHOL67at4txMq33uwcsZu3RNpUmoK
uxwABiJDzlEq+/vll4pcrL4e+a6k7Gu9LeVRk/QsCg0/YNtUqMXsZX+nyc2TVWBx
fWSK9E+C3Md5O+rcQkQ5hk32z+f8OaQZbuU6UEdBoHR1FJ7tnivMuio3hWCCH3S4
P8lMfxl0pSlnJJqjWccBAlkIYbRz1FniFFInzQLJRypw4+Dg0XX71ZW9pzTD7jhb
igYvQkvq3/PVpxVH3oYrJKpBCCO73yV/x0oiidIlGgKXV4omQVsZ2uU6i1RXzTHK
ZXWNtWmUfUz/5YNkXkzACB58jckvUil5ldndTHthsuIzRNILnh//vLYjVRRTsTv2
A10AIbX6/TA01Mx4SerHMZQYnj11mTR2rXlEVfkOt9vy7DdsMPULvtYXdD/nb6zw
ld0LJxW3NvbBSlDM5gNCZ4XKc8a14WZAiiLmP3pQ//X0922UHau2qLnxP7I3B/EM
/z+BpXimOd0kbzQ8jZZiDfzdFJeaXx6UGe1kyLqupX0d3tumKY/2exMmW0QB30mV
+OFGidOjZT6j6YzvF8TXJVXLp1FIgf5tKys6TO35FDKxDta3yERDQjh+NSoP0VNv
SOTqjT6Ss3a95PxDLLTbBGjUxWcR1D+uu8GMdJQC48+/ekOyKV1yAoYetqEJjTYC
mT1CKs2z+olNFnflw3kilz2y8JAnuhBQIWcJ6ApTuS3GtFLLlU5RXppDp6U8WWNj
ITRPeXhVTRETyyxtBLC9wPlekh5zBMRPOH71yEIm9qmNYD5K1y80IaN8bhduCA2w
++upihoyjCEa9+hWpSes4ksQrFmNtRPjOyUYToUGgzSsmKt11JcVW/ajzYiCSVZP
TzG5nzXp/r+LBFD+DyV4Iqa93T4FwLcIO2VfKFjH0/MNKcLjUmV39mKL9eBWDhQ+
ppiMYoNTlK11SQDYsSJj7Kor3NvzYhtaVXK66dVwsssofGEx3gv/7guQIR+HlNfO
DRIf+PtyQfBw5/BxmL60PCxaZj8PG1L7XdFGTF85QT6jyyQ4iqbf4vKRNTJBCAEt
/ejg8juc60ui28OMhJKVaKX5v+dk9Fo194tF0RG60cTLjwxwxRsZH5D0VAxbi2hf
aHJs5t7YOrW9YQRXbbUaw3puLGVnSjAdYOW2beOgEanD6FkKf2bQp8wVzHHwOFEL
/pYQxBUK7xiYXzP7ulg1zPFK7SmtBnisEWDcQr4gdxBretuubkwFA/Qk8jm5Ck8k
P0Zgc1DSZeSukaCyB4XuAFQbIww0KvHUZIUF1F+PylhjEDAf21+n/hVCPhSwazKB
yMllaLJWwtSA7QV53ocUlWX9MYWd4pySDZcR3MYKxq8RSuUd+H9lYCVZAZZKtUSE
GOzbqkEaQRnFD+RfqHOwvqY0J2+ACc+Oesm526QWhg9TsTlrdz709I664ypRBzUX
YJuXUg/0OchIqRzG7MX4+YyZ2w+LaH2RX3GSjInQVSa+Hh7MNDW+kN9HWBQXG2l5
9o7bXg+7VfkRfp/QTjtl6+d6f/Y94X8+qVdJxTNnS5bbGood0hDCVRn3qTj5i6X+
1FQKbp3GsYCmh8jeYGUa3PbfvVu341lPwA3KFkEclUK3ep2Xk+a3Xf41/cFzPRSn
M3Aj77bBjYMRMN1/IZ03FcCXlbVQmpQB7u0uyZkH8O7MsOfeTP3yeEHb+KBzKbyp
R+yhCfJenQU6nPi1wGMu3XvBSuUkNHdShPnL5tjCp2/Q5rchYDx1AyG7VA9jctOo
i/PyL6PyuedsYB+cVBZWQfHTWTBHeFlqBGIjBWN1tz3XBCz1JR5Ja3bOYN0yadfP
wM1O+qyNVTf+OI1G8U1FJFvqZmZzN5JIzbSNlbIvlFb2Lyu2/Bo/qKidphxlVQKM
b4yW39s3tie3GSB7PBoW5qpv4Cnv14fMb2Sk4gbSlA9RQL1ecy4AlsxRKSFPFZJJ
4pplATdUAf7csAJn1I0r+kzDFl+zWTuldovB2y/+t30b/0GRUcgM3+9/jDENV7/h
MOHr79i4Tp8jf+WK/diRC+gakzTfgK/KIN/4bguw47CfseZs50QKYNq7ew9oxZVq
xKQdBMGq7fH4OK/1vaftLl3dlErnwPK45zv4R47pWDDn6h5r4HdQxkFR41L6lt0X
006esMjOYCFnibfSGNmci8CKoBYHC2MGB4fNO/KpaAHR/t9fjm/CwId/hyWXN0Ou
bIQjSj/D7ch1lYTbxMa79YPgUTDKCz8pXHBshcjktvtdV5vTMV/+mkUY8CKLBlaz
6Ok3HvF1rX3RLsxL9AiJmJFuTyEnrq8tt9kIF08VJbgoKFhnKSCT+MN3Sf5wX8mT
/3r3hBA3wSi7usS0o2l+Xg7Y9JCBOnxtUWlf9PesIyztayMmiMX9T+zk1HHy9jg8
y50gYCJIfAkksuTWeGUnJcpLwqrimJO79dhizM9Z5u7WcrQe8Vkg6l/yrgk9Cj2T
xEreNnXdWPkFJ/W/SXtFqecjQH73N6r8ZR++2dQDC0FYRdoWLkR25yElFREHPMvd
q1VggDa/FfEhZRISTQLovyfm4nez3iIPGkIboqw/fllu6ymru9KOFQ6Z/g56XhOO
pI4iX/ti41cFQTt5FaXxZEQ/48B6Bm7uxrGFOHJFPzVMK4WMO/GCBKKLH9F/Duqg
5YyeZyB3dAOiXGGfEJZZ5XaG8FXIIMT9ijFAScFnCTd2xSSzF+8wKod5Ri6qcFgK
+oHAsUcLdv2YQUHH+Q2MM6FqfxRdPpmpF1ZyesqNNlke1DUMKQ3HM2wAWZsReDGa
diy9PdVw+4GS6PQsbyW4onJKD/pp8r4iBQgAacp5h2RcBpHUZFTLu+9v/t+fDa92
6IBNV5yfjxfeWW771oKGycus3WJLnlPhiVdXDvfItSYhp4KaSUFX9JAToRu5QLWk
mf69se/gTMFy5BKuMaaSCqbwnhBLQy1NXXjiPDH7xPrePvmXnBPXO1fKmBlz6VXb
6zQPkDAYRYIBKI4mVSt6b1IVWuErlG3mJSP7e5WB2uH4jOQhmtJWj3PZpmQnE5MH
Cv+NVTeViT/6eDcR017naB+m9NO/7OIXnObpwfGXO3kSwE0eb/cxabRiixnT+a7V
DAKTglcvMtsQsZl3RAdn+UoUI/dRP7RHbywFT74riYySIP45sb2eFLi50pgZlxiM
tBwuX6yVsVG8CcKxinZXy8dzPfAeEt6KQ8QtRjbG3ZK0qnt9ccDc5i3KuS7M4Ahv
L+wMElgWHVEbntH4wYAxr1cHdxpT7HRPrCBnyHssRpBJ/dQQojVgmcRk512LF4Nf
cpmye/6iYaJWkUzl6wFwvtPfvs1RPIX4iLAHZTkZuIzI1qpJ/CO+vVOmA7BjTC+k
QuqZmPkbw3OqCMeXcZc7ztYqzhdsBtc38VhRoZ1/4jm2+iwlaUo/LRlh4mVKdUmC
Oc2bZO4v9D8QhryKGRZoR3Bo8Qmn8FdJxbUym5niuY24QgWpnFt9aPhVwksMGB0/
K6nGuUDBA0eAa25joj8tDNEC9vxBihwcmIJsY7Ojosn8uOHxGnXJg8eoauGgxT3l
Jzs8kAQZ5jb1k91XwHKf8x1BkMxWAvu0ylnVHYRqSRUui2PECKt89zf3eltverUP
ZfvRE6c2IP7sHOFfuhGmwTSZXUl1xzxdB2Q6hoILQ/GI6VyJOEGF13dNvNy40pzn
VAMG543kAVPY5e7xrJm58T4/zbpBRKYDj0Jza5bbubmkgwAeB5gUEW6a+7vDkI/S
Rv6UJSQwpqg1GhHeYWrlQD6CAF0+MX1M8tEab85LI8idTqI/ei8/nN3V81wJqzB3
83V/A+FBOijNRS8VtRNnRoGqditMlUlbxzuhcIt5vST+Ul2aTLN2RDb4iBFOaaxO
lJVsnslTP+Obt54L0caIPVlRuXbpNOhvAogIxNBwmAP/f06+xWSkG7NFLPTJSSk7
HyNaj/ypy5lo/bRpyTahD6NYutaVZum69tJvj+cfKd6/g+h7LOxAvWuLoMLCTKYv
UMIyuSZVoi4+b5Su/6iCPDecbIGJAih62j9aTEFaUt4yZdDIdNfQiC8lxDGq5G7U
KA7upj2N9iV2l8UjTkf7iu+JAev3FUygvUi2Qd70MI8ohLuY7z2467FNV3VLu++T
wPUfcCDZ+yakIetl7DVkCLu6NGXR2uolAc6Nfcjooq8GEGHzCDSJHYwVwr32yO8x
18Rjvlbni83MZxEqUSQiUm+KfEuSbYjIJUy6vAJcsX7H43pOsVs3g/SeSg8ndbW+
kwZIUbzk0T6GS81yda00IxZj40sl8eX73Mfw4u15WtHq6mhXPF2tYIQyFFS4bSL6
1wgDlNSfIlrr8g2Bfd9se84roz1iLtlsbyBxxEBNtkKOf2VQHusMzwXzDxqBUXim
7TMB7IWM8iZBYms3KTCn+DyMygezjLO6pGxooWiTO/pj4lNDHpaBKdaWecJOzKSc
YqpRU6Wr+Elfrt+oA5GCrcC/XuIMSBeAiyMU3nL4wAU9t+3hUx37MnJFA/Iu0Kab
JvrMnl15IHdLjGNLlo2RU782zslO6LvaetEMsh0XiQC6AAY/SghzABRqkYFZnbZW
7LU1bhbssKxCjQwR5LJXcaCpWvDa1xocxd5FyB9Cdqm0Qii1xoVBuiQNK4AZVv+w
kUr6GBPyxRz1aPp7JQ08OpBUCNl/9NiorcxQBeacCxgIkuqbbiFMtbnqhbhRDbMU
9e0p6Gy95jmSWy+dQ0InD9mdxoxyX4jENsHqlUii7M5Cu89wuNviZSOapimgdyL1
i3DLldOweSdqu7xhaBk5vO3N4Ia74izDSMW/QT2kLNCcibG777VwIdDT59i8D8/h
qmdtasSvKjDsD3z2w13nZGC/AEKUExCveFCgPYP4gYvixzWNcfD7xou6xJTqHuqg
RtTS7a9UzahZ6ALEIvM3G0tLJfUMTqa8KR/T+obJFWRUna6j781RIuwfStNjuooT
1I1v76r1oJV4houFNmf8jNre/WjUYYmvfNIBZ2SkNIIs1iCm8NUh+AeP+spPM0uW
inRHFXBEdigIHXhMfp9tqxgCn1AKy+HCPP2UHTxzLbuamu9jE5bEDcTaoy+GTMRl
OmLI0SfdVjqmzG+Kq58eCr8KHAcodxbDwM4AtLhoo9U5nGnPfGFRsBlHiHgWNNwr
kVplM2LJGeh5+0psk2/446jKBpsQW4c8tOFxcAjFcw0iPVlOSYysA9iF9v4fEDtm
rG/YgipXg4+yAoqL2/wZMCtvSPkUjGB1HP6Vxf1QIk3igtvyKNn2GpCl5rz4I/Rc
VVj6ZADH53b8AwTDsaU37C9XMTvZ4Ry+Gh9lWzVtss3u/36B3wzcsR4/QxeWm7MW
olpdKnMTaog/Q5MZN23Ok2vqC9AepKyugmBIbVLcVotdY8ZfU3fTIpcWxexMgCcP
G1LbHxnJlhHd6KvOTAPgB3GAnzIGFIYw6j1bQZxNxMouQSCdd6LF3/vrnApQkwFx
DnB8gVU87FSV+baO6Z1wayQBW58VIDGBAoSH1pvI47fSVgJId0nlav93QYQlQB6F
WokPRmV6UCWuXH8jpHxXVrRRShiKfVf2g/TefUDfIXt1bTGCnvCFosS1phxvruPK
t2IzNMWCJZvqIwsUl1wsAcpDBtu3YNq6Bh4T0Vuq90sZJwVUrjkbes9lIo11+b7f
+AxxCVoVFWbpajIhh3xNhaPrSljEL00Aq6FqpYMtR1N+FTuAiIpce+gKjQ+7xhSR
7F1pfAHZ07y9ullY/Ui3uL4g4X7WzipWbcDXwVVgmh2MXib2EAWNrS6MTgA4/IUH
C+xu7D5sItvUBNXDRJF3dFimFVTpK93TglBc81NQRKToi7zIjhsVn+cL+XGbtiOL
eNLy+m2w5Owu7QD3eNTVHkpZvmUqSvNNiwKH47XIeHDrmS1gyuXs5CJmKIDK/ogw
rqBriIZbsFLYoaZh1HkCNxumstWabwAgYTVIRUSR9hNAsBM8m1ZNHs+MaSMAFPpz
7Nvo0FJ1BAl7Dd+RqOQ8yxPUk8EMx7i9ziFLw3Yqh1hWkCYBbCtl1MsbccuDBbRv
4rwkTt8UXYtK3gY67oc7cfOaAOIhZmggoz1VJZ3h4ESMJLWX4ny1gyjWD5m3gzKh
8+Jl4HZ8HJNMJYIlqLLuMEvHcoWtH+zadZLhlR4MgvNXR6FrXMbRrFpWlLuT358I
gSwKOKAX445u1nQVMfdrRQq0IAK4T3J+cGSquaZXXKFtLElK9ojIGSZLiZyPntQx
MaY+YkYDC5H8npL+LhT56x+jLaj3C3I16TRZO7Q9k574wOuzYMif/My50tFbFfHD
0ZF6datO6jdf8QAe3GctD8uDM+lZ+Wnqqq1JisoJEHs7NCMHKRjg4vDN4R9tXg1G
lbdnILBR8qlPCpY/R8XBpCTJROgZXC1bdYnBJecEhmdSBXkCkd089ehC/NLMEb1w
TAFZdxIGLMy8MFHKcGqyxtPbnZ8vi1nXzNoz84ju3zj+9hWyNd0mfYG4Zrsat0ur
lagdvGyJKtfuao3o6l02QOMlCQy+NVUIfVRc2R0gxdaI1OZ8p07XHMlR9mJ5PCcr
jlQ5W/WXA7k8f20YRavkKFu8xodDu99/y4sU7puLgPlcmSNJ6henXNwVueuIJSUH
y9F5Be1P6ahLBQZGkeQoMqSCO2V2WzDVtHllCt9vj+JE41wB5ob+eoByWAx9H257
2zrK2zghpaIfCDZNd7m8veTKqsSn9y+wDCh1OTqGWr8qqziiKaT9EmsexDFakWDq
MXAk0foTW+EoHJ0llmBsy1/9BteoSppYLljBfc2/O3JdVxFUk++WnC3f/ynh8mGL
i/sTc4FfkFF6a0Str76iVMFseLMuoS6DWvuKIf1zbGCq0YIcCyqS+YsJTWCqXI9M
+iOE2uq0IrK7f0Cq5QgDXN102rm+IUTxv7QeQu+T0tF2pfV7Xx+4ge0f6pMklOCZ
7y2BG7Q1yGbHhkVVWCD6WZIrDNLtp34YusBDMLpFpyeYq+dAsgKn03isCRIJ3WVZ
uNLKPw04SUlhIr/OC47f0XO/pO1ZuYjj0TyNk0hcLOFgIBhKEQUntiEqfC6dYQPz
4OsTB2ssLGeTAfVBEdionKo0ZnRUCLgJwrHwEmhozjOc6SYKIfLDQlI/lRRqrJk8
H/hxYHgIzptDwjhXIMneroIKooB8Yq+KOzA9p/4x33FaF4ZizjoecL8hIVj5qoHK
RbzHnN/G7K5jnB8qXmIH0DMvfgL7BONR3sO/JV+H9PRjwXtsYKEpLorLcsRMQx2q
Q4oFuz/fBJeXfgNqeVVh3wCQgSbRJQn1lVaWK/B2/ycwJEUwoGBTY7n6J5Ls3sPm
HIxd66KGDnxJSqGDSJB2rjKU+xOd5NCY64Ws6JRNus2NOjWkAH6qr+xExQXz1Uvg
0u2PVMjLq2zDk9mJHxpGCDUp8UAi7VjNG0nbDRRpefq0sUJPukiXWlGAw4YhDwKh
6uftAdDKMXFL8jK+mGk9kFinB/T1xn88o0fMGyT7r4Ua4FvGr2R7woBOJmJ/9Z0w
uz3AJueB+s0TnvWgSk1EFfphTvXpwxyk1D2gu4Mj5EzNf0jbsEg19yDR36DfxDRB
uyOA94MGoIkZdvEVbHa2S1Y06IgOwFHaJZG1hGufoM+9WpmBXGvWr0LYLFqfEvxv
7ai1BcF3r76R3yYkXb8oAoqvec9yama4br5AvEdns5YumEP3vZ/u+vDarA5Yrri4
SermpSWR0hgl1tqaMti69VEFhToplg3GHqMJYOLqVPjpQ/K1am8ji441AeLlz4YA
cRzZBYQb3UeUqAcKmwZOoQAZDOLFu1EzmQh8UyPzgSafBbANIKbmhgnJubAfleSM
xbKRhIWjh0fLySPd9z76xMYdg5MmR0T2HULTX5qqMreIX5iwz4KU1IHWcPiMzrmm
5Cobagaf55/yVKXpWdtacD1IttloxmKVAoDL8RsK8Nnpp3N4DjDcO4yNt6GL3Uy7
5hWzb3Yh213xDddMzkcyHdVNeBchSNvhdJ2zBWWpnGh2ndX+WIk6Sa8uyd9nlX63
g3dxPsiSzhzQP5m1T+osWXY1ArhDjgLqy8yUL7VbknCcIfgPxLEyOc4t6dghISRM
ByxGA93npdlbpnPtmLYmoCJ3x76SkZ+ZGBPB9/SiZ3e2SBGO9H5UcKLg0Nq3i0uH
YIE8rUS8YQ5bY2SK4PjucDpG9l14z40rpsryhQC6PgecRRLuAclyhEfFd6HKLcJU
d0sSa1jMB3rILoJAQ1zWGOPHwD6riTgl9qA4sRBA5LcMh1cz1hFQB+f2hgCAq4UV
ro38ZdfV8tNGeyIdnj7FQ04x4rdoXR1DGrJ2xo7FaJgLjfCMyLl+b9u5YpAZpbOW
RR/tnh4vlduavuOWvB26vEuYwAvCS9xLUtZXmtuqV5ksFi9/88+xMRY5tBbs0tNm
vQLgWQuGuN96oP6KfMWTX5oD4xQu1CMVkGtSMwDl6xaf3KtOYBEL7xz2+bPNAO9S
uGQZCM4Rc/xlgIHjY84GltHss8izks+EBCuQp4n3Qxco+/GgrpOPiXCBoQ28aigd
B9rKwsXj8xZxfulCO9QuUdml5ocO9VNBTRIZuCELvmSC3EVlLY90hHGafCctrLqn
5F/OapRYQWisquNnec4K/vnboHGsrMVQ3yzmz8hmT9KfXJv8UULXPVqECKA8aKn8
gPYxpBdnV1A7TcilNjV2/EzMxmGrwIC92YI2vQNDnZF1B/wPTxeen/J/HaiW6k+Z
fO3s8LyRZvDAoLTViUQ9wXBuX2XOYLPMUsoxcnkRHdf699na0DaFtsBRVFFMRh4M
wgiX0UZYMcjQYq5XxZEZlWthLePh0C1jayRixJCDa7QFCIbWGdVYCvdQS/1nKpoA
628m9gNC7zhGw+mq6TjAfKMYBKr1U1Y3AWnm4nYgTBVar8JrC9Va7fSpXsiy+NhZ
RoINhP3ySvxmbRQ3wODX5GVAWHOF1TpiuoeoEn4SpzzczOjaIjCz6VLwOTEQHkYD
vKL7pwx632puYQezmsbnZB+a1lNtHzo2dyrlfpliUVFEKzAl6iK3SnGGmpEbKN3k
NPfkIZp6mTsSj2sSEtK8G/+wxXXltmmPCU7NYS8YLI52T1spi3397k8TQyNGOpgw
z4xWONj9AeXbYtofMz+ibstHmhulDbkdfGT8gO9Wny9txEW3vfI0J/gW6ce77YOI
VWOiqGR7ThaGxRyq1f5OoyIygvDh2v4DmW6nAJEoN1GcwgbkwL/BCwEwc137/I/i
bOCaHlXtTQ0/pdLynFqzoIGOq3zjsG4x7Z5hxwqNV24smSFbW/6Fu4rFAJ6oLoXU
oQdrKywuiLRNqpWgTR1lMXaf36LP9i7tEA4VLivH+gblVz7B9irrHGZMxaUc5A4Z
8Q5yk8fNEl4zh+DLD3+FbPYQTkDwBxMGtanP1upvYu3psqUL3pvkzoy9tfQMFCRU
LmZrELayQSlmfhK7ei9W2UTMzgZSC3lrfW3dVmzPSnwWVamvaFV5tCniCBimdJQY
JNZxsqGzZ0FjPylPu8xDPjkHWfNyFQlDcPvccjAEckekGpNiy5pP0Ul1BbrLL8Cl
6VSHQ2t/+szWWDdE1Zz6NOcAaXj5R8n/oWHWXUQR4auCKoCIyL/pUGHjpc7B57m7
lwGqYm4xVL+UpmEysTeDCNs4P90oPoZWb+Lc6USoetWcBHC2ZazSIaBwRrnRB3VW
gnKvWZhyEkogM+tiPV7vVGMkYdZa9r9QCehdvecQvZMR8ymyEA3q+ZBanrT+7GE9
UU3OaTrKaSWhgdXJOMhbQNGdnCNtzNutApDOhgt1jWxLkkYftbRd+yJVqbamjaeC
qqyMacNSH2ZpRukTUu7QYbUXk+mdoVcZPvHsQNwH1YobkLwBgnPL1TebnGtuoMsi
TAZ0zFH0GWGkJwGYIML92fymOi5n1r/442PBqqNTHCRdbrnkx+uRCIeOZOWbbo65
cjA1LrLusHgb8nkWllKyl7wVzf5+c3xp3T6zNUK16m3F9yZvhiLd4WJRE6Y9ZarG
QTvSNhKRzXh8Mnvw77jWLR+X+bxT5M4JIgknzMiJAMmm1vGoaNINCIl7FmW//owB
Br+eCchR2Ckin+gPvJ/Kp74i99FsT0jjbB35qP4DWTRmgfKpKmto1vXyJdMjfNhv
amTE1piQuVGHxIE3MF5HvXSCZXU80Ax8i7KcbXZp8RF01J+gbjfAWo9e6XxTDDeo
IVTveHTQDM6YAqXKgmDcOKcJUCAc3lgFhViU3h7WzdvLQbDmLbv3y2PLVH9YWZ7X
udGdACMrhd5KRy1W6o8uHVe53I7XE57Tyr0pTqwUDTOD7+RYgwYeylEivt5yIr9J
cdqdR/4K8EoWpI+P9hpKFGYBj+MgLzB10B2p8zvdpR/vWaqMCci6npZ/s3pjUL8u
KA4euNZNQ+BeoH2mHu+VgjlpqbN965Sf9fAUfxcdQUHtqHcWWUcBv+e+rT2aHdhv
5fUkPopHjSxm4p8KiRQs9HZo26XFkyqhMb4APp3zT4QfPgEfCkFut5VeWcicq6jP
y75iBpKZU4CxOHbR8+dxjHznzTaxZt0ESYKURYt/2HVXYNSXuJn6yqFrgC20fz02
HSrOFQgiunEWBJ85GhfZQIOPZIVMTtTUepbOd3VkJqkUSFl0jzMG5kDV6jkIrwGe
jJtGNTECh1GMQkfYUamTKKGVW6GAzVnNs/80lwVSq2J16qCzqfAkAvVuo88K3qLs
RaupQXC4n4P6p4U5U+oy+ISXaWY6GKaFkQ2W53zhH4NhD5ij+z8x7UbyvdpfMljF
mTy5hsjduibrCyEzUtzLrURpRfJnGA+mfehjxOMT84VbyrEbL6MhoN2Yl42f5Hs6
7z9csHMe0GHAbO1NgRdJsoag9fvhaDJP2DIC9E/ipIGfnHv0N4TxI6apQFBzmKFJ
7d8GD9DwQMy+XNJpaY1dnKCRQ7GhpdbJoGJqM4D/f89tVUhMRvd1lRTKe47nC1DH
w/Qi3/RLPdbi4p7nZBU2sc8j8dHTZ+Ytq33C9pBvB5jKaMqUh1qQDyTW/K/omu+C
OT4kmzcBZkPpPk7L5xbprLdxbsz4u7zALU2AqcbwqTGBH9qQHFe+ZfVOj1aMhIpv
COESKAGS1CV1TxZHb9+j+hpsJlJmWIPgCLQFNQHyGhHkYuaEqrvG1eIt7o2ZBbTe
EJlpl72ZAFHofS+1g7J2lnpA9MRlIEtH0JSlLv/Yrcv/q4BjGfnFhfn6wWfNnm/a
iQj0AYKjIIMbL6yyUgx6QVr+J2rLM7/u87llE8lE6eoobPnyr0ReZQw7Hag0hC/c
08wLgg/57YwfBxG+b2QOtBCU6c1SzKEAO2bGTncj7enibUHRXt3cckYL5vOox84c
BhKkJaZcxSY23wNmZjb1v3BWzqg1xOSCVs5KUGOAaUA4ZlyCzvAfRUucNrspo+nF
H6lLoS0uqE589nr8PzH0HSYpOMRiDFH/rwFyYR0WDoeSo30nVSY4R1M6aOPGr3ou
6l1XTz3XkQgTs+KlVJmsEy/FhLOd/sPItRMToeJZvEZEfXQ2jYibAKPiHFNz+DC9
YQWZoEXi1K9tgi1SHB1MDm7e/oIauzur3zKG3kP9nVVq6Y+mIwGleMNNiuLPD/8k
XUDZ5kosLcb8y2GB0nzVy2+jvkum0ZHp1STEblAozleZt3W+SReWXX0zHgglExMD
wJKRPso+DYVbYy42PqdR4myCQIycJ3PX1B6/zpEh6ngFGsgzHlyIbVEPR+RfMqYC
0d0VzSAxjCSh/T1AeqAZ4wwa9y3RO1XKTjsFfJtyb66AvjMTgJxbSz2KvngsGAAb
7zm0tNh1yQ0M9PR0AuzlzJtvuN9TVQEa40uzjicJvBY768dBd9PCYEhhQzQKaH6h
Hi0siMbNRnZJn2s30h9kyaefk2U0Y25cbTqbCXUP4aJoVLkfGHBIzPa9NfiFaSLE
L0Rb8UCZl7+5ZvH4qEoiKihYBA2/lBg31GY2V1IErxgnZdqGPBTN2JvnTbV0N9O0
Zey2bBHonsgsORTd2GjvSUg+3qEBBMn25aIPT9i9lwaKQtVQ2pKwiSgdcBiVq/Do
W1yxf8hnyYUC2u448vYEdyBy7FNt0XYP5U5WciW6ZBjweC9z5XFOjco06rRnW6IG
1q9vAHK9u2d28PxUyegCPfkUlYlvuGNabObALccHhGjqWG9hRM8oIv5UMrTaor7z
WuyI1lsMF6qn0XUHeOvhEiwZnXO4BlwupVaQfkOv7TDmZhefSMaKDCVnOw++k7ox
V0vafMXiFPWGbsQ6ptrFGsVtBDoaawqxHIdtvYvJ8xubuTKUL9ZxAE/Sw6qvJScf
ZLFNZHAMOcAW5bpyDMzLAKw9+jtBX6nV8dDlnZAsCtOwN/BLlc6ifwRjQNxEdKYl
pFekHe3Dg9gUfjagUIDYNpgIuJA62cPS0eXWSXIKzrSOUvyWNhBL8ATMXQDbuIUY
7gUSUfPUagKpxguSzVCvukSBYIjg0n+Szb0xyAB6sPo4UxVlOPzNbtZfA14rJFHM
fcsAi8Uk9uEy/m+btqa4MweggCWXPkjqv48zrl3TdxZeTF4WprQBo1uTcYDf65Xb
hDqGkH7InRXx9uAVWdZcke9oi7RJX0QNI8D87+zqYby4SHnheuZx6OA73xwLNy5s
pL1mLLKVSGrJGBz0EuXh3DnodfYZxaCLkDAXHGWF6NOByIB7Lv2j5QsmBq8DzZNl
08VwjpOP7WhTDyAqMDMRZz8B9VBMpRNOKGekbH99HLccUsfvQZNDH4z/GFS9djxe
zw0A8tsANUqfzenrmBA6D45nfJvJF6FnPIJKqfcIxsMoSLKp4Wcr6nSJAjgR/ijw
C0ARwPGhM9P5KJ0vkjWVdwxqHM08CaTQVtNABuOqdVtB1gxAAgkEC/xTuKFPQHOV
B1+U/RQJ1vg0Lg+jdxNMxktRZHiV0L8yfC7Bth8yoos2lPmCS7tNMRFEMy9p3Nvt
LBLOZsraYmQBy0PCdUUYxrZ8Nd+Nw3GohqQ7ohZ13+mVmsrJZNEtf992HbHrYAPx
O7e6EkKzN72ertEA9MFuBMs8ht/R4MmtdRwzEAymoTemFhFpm5l3oDBrSkfg1UXh
aeMG8cCzToGbYL0pog8tO4ZO13rnM6uTOxCHSBvT4fbykZQw/zTSPnbmItF51zeB
1BZWz+uTkfArhnhG4gk62/hseZjCRpPa0JAWuf5Hcy4rcF91AILGznn65VB0qdmA
sNXi449uQUIUXKiYpo28fdbWYiIUFOxpfDOtuGc0/fCE5OIlIaFFbi+nhKBtaWmS
FD42uGhQIjZiYUK2FYPWg0Ze1+RuIz/du5qsxKwkBpjOVymFOPSoej5bvtZ2jYAE
w94YV/3yXR/2atm5E3jWeu6WoAu4rK7IpI89iCMCCfkH8zim8oisLPp0WZd0C3jt
ak+HGFVJp32hI21tuJX1ep1PfF+1W04BlwpgW6XVGJkdr5i5moFXBeyP3T1YhfPP
WP6QMVUquXl8EA0kz4Fc5iYMHVRdgZoRDfnB1adVsQq7pfwLLSEaA4UWHZQreryA
C2mkc6To2LZ351l5wOmrK8D7WeUU+v+UY14N3dpZJfVFcA+8yZbOEcxOfzscVvkw
RnlI2xlfuPVbfESQQtobSQke0AjCHJiLr7wCPaFBGXUnoJpjg8HozLxGs0wF4A4o
aXJ579NsY3mFSruXn9iMTb46dzZOM67mUSE/BuzMCw3i/auTcmCoGWTvD/cGGH7h
zWq2IhYYhyq8SBzfcWA3n5K/ZI1mnypkekggloRYwN80KW6ILO9NeHhazaUjG6kq
eq7vEOPUXESSny/hF3c1So31H+Rc56ACMe/M7jIlApbCi0NlzleduPFTUoern4qi
S/nQNc/K6OatmFE+B2D0nhHgTrr8mbsD4TOR5ngL3BwIdFJeKGpwXicgY/8J/z9X
8NS53XETgfc5UDL+0kuvA+eA1JimDfCGUMzMzilEh3T8mpfbFJDlc47WwXhpIcn7
y2rfZF3xHXDiIs0KgK0AHFbqV3YemlfHIW1az+urPFbe68tIRm1G8hxXulu1pwpG
iwzx1WGvnydkTd+Lm5l6TsJTUj5y0mP15wbp/9q7chfJkAj6/eYYi2D0NDu0IcMt
trHgJTcBZ7qGvF2OI6ppe7VLJfU1qZ1XccHMiUXV9rC8Sgd0A8iQhcc4b1V3yVvT
rs9aZ9bjJ41HgzyRwPIRpdUHFG/GxFJrK3ThdEVSexcVvd36Ff1y9nXT0jWNdDFr
ViX5j9Kr8YGv/a5eKekBRdVRLGtmri25Zz5kjjX0XJM+YG9keoeu6A+UXttU1QZO
2Lt/lKIbDLZrFq7HrfTU1srbG/BaweCsdjEWDbyYiBotqxgca+mIVGC+ByGodr6+
Zt4uX/kJ09Y9QJnhBl1SN01TBx4Ae649/uwOcXjMx1wfqd6a7lSA1YoS6fKBSdub
7iveJ3vtdfHvWCnh/ct9YkDxnW4vohp0i+ogmGqOT2Z3tiesCWtQMXNSsx57Z4M2
lwQhrnhDS25hG56nKRJ71AP3l9JevJJUKdq+M9iwZiFa6ZGMAJOGr6NVoPhkvaS2
Jeqgra9RbXw/CpmLrZUFYjqoQcTLlrtGkr/Ng+62da5tM41xF9c/vJo8LykTUuDh
spG0AEGrqVqtJn9D0GSki+ekRym2WHNDayojJaCNB3ZiLvEaaCqut/jREyAh+gsD
SMpPNPEWZx57cZA5EciWO0xAzE84MqikrLxEcfDvDZVyfBjblSCcqtwTDRMVnbib
nhXKD1CeOl6WXlQ8TvVQu9aq7A/OGW8PhpbmWwbvoR6/ciBvpij6fCeKpBix96yb
GrkeSV9oOiVynDmSswH4cfa45caYWwhJ3kqXoFCNd89Tds53LmFXXAd9H1KbBfwd
SYXGy7O/tJuTJGubpGsFVBXyoo+UjKMbtYIFucVdoj6KgDMh3EbrTjppvHasyfSz
ohPFc7msNbZboveG6kPyyfhihSucHspNxQgztj5m/5+GMJ+kLxXulNZ/TKwg9518
h6zueXGvOWWUUNrJzDCKPs2OJcE8O5xf19KjVUBW+V6jwDJTMyTJcbCd9VN6OoIf
7ohBGb+f8bHCSSygKGOkImD6GTi0fKMSiyDSdPVGiZl6fF3J18hMCkAMmul3exO9
3kMfxjyXV7pgdPSE6xtfefcDiglulF+t2E6jBMdziUCFtWxh3UmELFd1wcx6fclU
taLdJi+PI4XLF78zUq2NyT4ULTu58fATLPOvF7TIfFHrp5IWI3/SXMiLQ44M6SVz
FC7PbAtOMCr6AmXRgshBh83mHeVwTYMQuv768XOtzV6Bm/nE+hjPDGxkqSUJtHeV
htAzt7aFXaArAR7KkE4O5QnMRAR2ONXxD/pik3Ubqqz0FT049be7qFJTQqfkXjuG
Rblat+0tkKOJYg+QQJy5ffIjHuMdtUHbPmsMwQkXqMFERTR7JoAe5ZfLh1ICae9H
hkc9iNZQHOO0ET02dGUgSwShJ9h/4RMoQVEPKTp3D3il+5+YKvB4oNQTDBEOqUsM
i2qrwqsg8M08CHqvUfR0Age+GfauEMhdLDXq4/Seo6OLdso8/20Q/gzijXvxBzxf
SHZsM1HvnCJSfYcaSz9F4bvZELCgqhOphLeT29GOQXa1X9ke6Xved7WM/UMUMHLp
TytuxamkZjJei4NmPzYBcoUMn3+rIICNGkJaKQKd0GjjqyUJABC0Rxwnm/gvJwYY
16c4ihLLasO1r6GykvAqbE4ziGuJA25xOxYJNpSKGeLVVVncW4qLhmTuQXj742wo
LDymakDGpg1nnssjcmHly/qHlxsIZ763a+O6HK3Awf1KOmJEB7OMHSUOWQOCzf3c
sr9FOPWQw1YvHW0GHS0hZFf6AXhAnOTvLQv7XGRrMJ/L4hDqO2mJTUdSkyjaJTKq
SzHUIAEZqr2AT3ser1ZyzvK0tGfIoYaLbd9rTiLAfp/7PJ+Fn7hxP8iwXSVHBnfM
ahZGSCWFAacqvXIbDTN88lbvxEHugUpD32RVZmpOQ1LkdlN8HO47NQjDaQXwdGIi
MA2KxWrKoRQ9SOD0yzR8Urw8qXOPyRp5awcFUFB/EragUsCsyEU/eSnwkesK5hr4
rNUwTw7hRw7E7alCiJOoe97bONNYhYNSMmbFz4huap7m6C7+xQlw6UDHUci6lb5Z
NpEwXNMNPvY8ldpxObhzslotorJjnFsbDhnQb3ROiNarq3825chX1a3yetqKLfKP
t+6lG0pQc8xIUlLou3/zH07GJkm29SOTzyLziGvcuJIxDaaYS2+VQZhRzV50svI8
UB+T5kiiZBT/ZMo48FYuwh5C0IxnS2BCGwjzSt5qCCYnTCFUxKWfIko/4HDl+ACF
Yq0XNQwLG11bT0w8AIjaz/y7VBshzX7zDDHetuf6UH76VHOvYXVEpacfRlazaF10
gXM5jkRnDScOveTxcyWxRTehWKFNWPtyYkII8amMprGpDuZPvyeUaR3ldPErUbd7
hqcb3uKJErHH2jSurvFNKjYLfe+FImJqy/O6berahIJf1qSDZXU3c3cprJxfw2O8
aCUgm6H8f6+v6qkJ/2Kk3zauR2xpuq3uw/DdurVOR0nsPNXuClPF3zWbwPY6jeTY
J86qz9hILbUIxprlaNhU/MPsoFXjL4Mwljxzfsa+X7dRMPrbUxyPv/CLUX4PILaM
PDElEKzQv0g9PHtsjkloVZyOEujPNapr7XR2ZrTPccGcQxvBQQ+clNysi1xSn0DJ
IZJH++XtZB/1bQk86pbjSpt5xs43OeL3v5oMwDq+SPzCQOANKCHGRQJmwG6tJ4wT
iZ+eeK0GSPKRpCmDOsK2uedHS5XBD14uCFBd6bD61sZvZ3sY8B9Y12aLSkoI4yAF
sjK41Jfh9Nn5XEruPKEujqNljZERdkiX9YeAhsk5t9p+hS2bAFz22AkMvkDraEfN
buabUJqHBe453w52IC3FD8O17IWJycS38qN+9RefROS9mKm6lsllcojHTHD2oxEg
DOPHnUhYez1ivXI3xXZXJpUqNBfcQ5kX9ccM3ScpA0bOyyrXNxSNegJ4y69s8iru
crqHRpBh+IpLOAm8SSreugeC3+tWNeCh4w0KmjbmUNGDy9RlUwhaCmruysh7747r
p2p6mBJps6tkLcRQFGUaeT3lJ/eRxWxsNdWAeJpWf1aUfzzJctRIlFhnHkDNs1kv
oC5cxK8XDuRAqD15S7QZU1kb2PUat+fahGYlo+MzKtwMLe+GguQXwMvlDGabSDSY
BiNFoOwp44kQxaqqrxjTCxr/fzsADLvZltdgd9pHguzoJsgTjWqEUI4gWwjip9ec
9svjsfWu2Nzw2dpKnczA8lWawDQHF7c6mYb3NL6MsKeEHa0TcGHyxjuckeV/AUVd
YP5/Xf32X5ODlyATi/b6ynvw90wBY2BRUEbl/yrpN6qJFE6u4Jg9/gm2n7UpwHc9
xwktpwWI9jc5JA61SmVBf6w5ZdE5rs9jyHbnWOlk9IBAsavK2KHCne+OLdoDolzs
lU5s50llPxfIkeZbDJROvngZQjX/uTL4rXImDJ76jAhbqeqv9lYIO7uDVKl2/dqD
ny2k1x67Vi5oETrJCzjCDl9bfWNk7wIp3lwe5Q9yN9vjnDscEfHw3HuwH3W6L87o
quM/SlT8Jv+lC5X1ymmVnVPOQGYc8+qUnbxMpZ7RlVMYma3EZvRbUiwYD6IMR0w8
HkLyBtYv2npw0wKKtyUC2ffnU124xMpuI5g8YnSlCEEk+Hpzrm0xZ9oX7bScdgjb
PFrB1nes5uHnM6jyDTtuhNHVZ/8xMMbKVl0Mf8DY9RElKcuwo3nFKKamTv2+3gIk
ha4v/hjn6iY8sP5nLP2f7is5ohauoKmF7Rcb7zcbrawKv67kJ5TgImFE66ojHn7j
iW03MlHscgO5Hn6/IGETnKfBqgo6lWWGnsf7qwboWlXip4PQcGafEkAvU/N1SNMy
qGBKtQkNaMQrtKBVdGVkhPkHjMd8IQlzP82Snv33Ph8+rbDH11/bqA1LSeJh0HO0
Ti+0m/DpDk90EXrSB9RnRr9+e5znPuPBOhCoe4krASLao2OHBoGlFer+DbgFVIeD
lMV3XeOcqU/m58xuw7WonUr3vu0timzcNNPkgH/fwb+nbts1GX61/fIALgF7d3nj
EnIkLkst7ViGO1li2a/M23Woyj4a3ScGgJyVxmxHLKG03q2cpx66TEPoaq+guLvC
sc+TIIztmxwYoo1UdlTzo76hU54gj6LVajbJS6Itwo3GlFbclzoMJaMgPTMKZKEX
lPWiVYCO2c+Pr1WuHBpPgt5GfQQnn/XPjiSoB1nuGTWB9+3jFPdIiLmNZO3RgmJd
jcdwyllXyqRo7ojE8PSy7Ry8wms/QpROHdGM1nZKhSbpGELvNDlJJx6rub0HFrlF
Xqq5uE5MAaHsGOKNKmrK1gmLFAiboWj8RohPE5W7OYp1pNz9zy8009xviR0tY+0L
AI8PHrx2jMbEaYhItplDmxUX3ZrTDLRyY4jsOR7GmIjR8DbP4GZZsGiouYg2mRR9
5K80hoEOa7JHJhUL3vKUSYETLznEjYhFzJssp5XkXeoWNM3RNucwGLdwaIC4ah0q
mfPZ4ySIlrkyQDnars5l4O9jJBXoQD0wNsVPzcN+i1hbgT1OpuvjsAZVaRuP0v04
L5Hkmm58/Ow7EjORE+MeQK3QKPz5aTPzzsyq9NBS03SyKv0b2N/ZZBxEU2RFsTxp
7iG+GlEopP4BZ17E0DLFIhYYIts3eUbMfYqipzr/2e4k5b8s93dQhANmAO04iEJA
2XBGNjDHXRkiEt6CgEYPvYLcXVR0EFCuH7F+9C7C+dk9FQfKe7a3EV+NIRhpB0A/
u+DmV1BSXsmoTy1c+Fl9J4S0YN8hIzccqlRGL9ox+zatImoX1K9Lxh68o4oiJMew
I+e6uf8IdytAODBcawNAwp/tF4yry1fxWL4Erto0IsJP2yWP0XB6TBWLsvHCSPzV
lRarV6gvQaMiIRFpQwwBJoRIUnK5Olt7QSRQo4oN/J6QP37O6rLbxqSsuUpxox1R
VclHRS2lbBliRMDyLQtXZHQJk4SXsIqFvKnWV3lOuWhH25m75Lz88e0yNvEmWDTX
IGugOgOA483XcKoBUtr26zC9jLCtquZHNDw+yzkn624gaT623P5W2OA3ltqwQHJS
3Hr5yQ24e+8yZA2YOmQkx6t3502PFecWhZBRmJzgT2Y7gkGZxwVZXoMWDMPxgA6m
nvZNnrA73MJZFfn7a7qbrjLuFtvY6Xo6FAv7n4rxtxfh2FNjZ4wnAqWWgJLPDM7w
XklCZnC0kQMK0YZW2/ixagpTJ6IO8k9MYjcJtH3GhE7mcvD0uEKcfDF03snghQfH
8YJwkHb8heONqF/r8kFT8QbIPmzCUdFG4/dTO1vyqILnKMD18LrMLl+nEIk8FE60
264Igyj5VVVOJOuEwJp+lGD7rycz68vcOVPUgCRCbI5rB4D5RxhK54P1JfaaO9gz
prVPMjMLLrCkga9B08kGlHE0g1Irl5E4ipIjpr6L5J333zMMakBVeyPu/DABuFWA
oqMEXUAXfIsC8jRsi4rJ+Fca1JLoA4xPcY4Mi35KrGdghpimGyO0oMK9OLgjMmhh
qViLuwSZbw8WHomEZVYSbemgWvpBG8FGQpnSUZFyYNZue/A+khNJ5vFk5VBaF1H/
DaGOGNDXNlK/l3GupI2ClPg8P7Y1nkoZ81s5kGgqJ9yy7k6WpU9zG2zf5UFbN8lu
sEKwn9Ta59ajAwZ43+2fqBGnPSaut01+PfQUAsLmw87jwrVmQU0Nw+PIC59oHjNT
w30whMtEqsr5uqDScVUtGVm3UdjopqdGc5+qqLuADntuZn4kpTNbWtUoM9H+Eaia
3AOR8rjjHYYe43lWeOPnuXLBal7pmD5IkJTw4+bhvmzDXuxiiqycQQ0Vfcl+Po4O
fws/KBsN3uyGOXvhVQ2Hvgls0qfyK86vWvmxXip7DhM2BDl9J4XF1i+y7rKT+on7
5PiTphv5xMXc+rzVZvvCYlASSS0M+IEXIHWLyY2AgPJr9GoxmcnWNkEwrm3pTY0f
RUpHyK0VRWd+KC8r/zqf0utUjM6m66HDMdEdLEZTTghONehpK8H2Uew+thhfuiuN
VGRlQ/IEbpkKilak3yFy0Ut9rFBvHdhf2maxJtyrtOmTJA2v+ji8mybPEjiZDfJM
wRMh4p8bztKA82B/bSuu+3rIe5FA3691/NEPhYTdf7Z//CeC4C8pSu4kpUE/+veg
0dh4TFeMDmekjBM3bKs2Rcos+z2zfRioc+/UmIytYPvbTBrpzPsHIXaUGrEDvyTt
isomEaVNGQQsrY11p2imtKp1SqRg2mH39d3vGObdukKjdqqY4L3k2afsHdDLZlUu
KWOMm5qiYkGhgS9Fr6jV1LFYEQyLRckgqV8E9KIxtgdM2yUCGfVn4qK1EzzAxWDM
As8BKhn4qS5Gduw3m5Ys1RGjkIdQI/KAi9E/wlfQam3eegVC1yomOg++YjVmvZZN
gxOM8Ffy/1XlAAZrGo8vRn3AbwBWZG3VpjNZVi2SO7URJWkyG6JR3J4wgrhP9040
2quBskPzxvUEbI9hOjWqyfQ1H02uDXe0GlrLG4clJ8VJAvni0htBJaq2d9w2ni2c
hQ4Z53Og5kD1IqJMIxdGROBC9Rm2UrjbkT8CAD26/AOO1/SYCiiFhnjkJakhXY/5
LhJJdWpYUCBGm2OmydNjv4NZXG2pWljbjzVqc0286ovYL1T5arLKmxXEu4CdnqS/
2kiYO17cj9HFhZkxRbQ+LFOvTkMs08FA/fw3yGL/JhC9fPHdwGlnhOmw11GMOpMK
Zudk3JEfC9KshgoHd2j8b73AhFnZl/GgjngaIdVJGrnSdRyuwUSob+jBim7RzCpO
GIt2ZVl2HH/d1Ia+H+ZZgnK1QP/GUpA34PKOnQAt7uqghgjYue6/NJd3y20N7TKJ
wY7HiiJ9FlMA9chZg2mMKwFUah3jY0VV/ASfSbtL0sPVLcmJmlwMRfFC+MxuhI2O
vupSLLcnjpvU5uO5rjA3x5u1bfrj3wWZC5r0DIjAZQdvc76ACf9g9yPoM4t2Dq3I
4PZx9q6kKcw+e2vsh/qePwfzpAo1FGTq9zDmeee859TiyzVeq+kzCE4fsW/9yv4x
5utBIOhw0WZbK1GnAtXsd+BFvmh4U+PJ2Ex16HaMjtK3NpAspUWnMpoGl4v1LLSS
vpUNB8idyFfrnSK0Vi71WNDi+CMz+Ytp9Yh3aR4Y+YeRLnyzu9MQ203qeO3OR4RF
jLkeWjG6jaDmAXXx+q9Io4CdIFYYcgzzraLkrpDyx8AGCt3rYAFQE1AywtwpoeD5
7oEEXzqvzGUAvHQBB84CYQXegPG4OqQqzsbdTI+4bNWeUe5imExEx3cqU+8xCxCB
YcJ4CLiTvvFzztMzsd5kc2i0OGJ75xXSzUb4C7YMBf6xtKea67c3kFAJjnclzJiq
ou1iXemz1duPVz9wlrdTaEWU3AZWnpNerDPqzwPOPyh8TAJNZQaPscmriONonzK5
xcL0gPn298hIOyb2zMn9HxdfqYARuzVoM3ANSd/HKM7NMOE6aZp9Vwg4DvskjlkE
7l3t3c4ReVWwNfiiQTvTxfVocQyuRsKvVGUibSDRyDfFk2/NWnyvDtLan4efVa87
fW6Ii8hgyzdpAMT656deTv5QZluV05J6gOHjBKeUedyWoeykWlTPE7brCySUEgdv
iG+1mfWFvG1wdgq5vly/GIwG0XQYjLz++cwThpP9ibnNER/i76ow8nZJTRMceMaY
/5EFOmWItNbJUZ3kHtMyF3nvByEAikCTlcQ2IEipOoHhTbc9YLfNOJfu0J06T6mu
BtRlHyDYYcgDXUbKR0IaPwIWxEuG9WtSVErQDp0U7Fjx/9yEto0/vLbytsjcmYA/
6POqhjB9YW7f4/6jvfyR76Dy0eBLl/qU1bI+tqHXEf3ZkCHAFkvWPzjb363pVPE/
A4KW+dDXQpOvD/rT/9X1b4dMWJ0XZzsRevFYMmDkQalPznxwpW5ajC4ZwwAVShrp
fA2oTLr2zQpethttGP4j5DvYTma4099BFWnixU+YKcXka0hQjqiL+MbNlPGmFs21
Vtw/glHxWqcVNda04R1eJ1iV68tBeejy/2fx5eam4AOeVsslTiyiSYXgsVRQ3Fyq
VlwqJkhu9iGR6Boa6bHQO6eMidI+k3UMoOF8vsFAjBUsLE1h9j3A8yFb9XOJ/cxF
JQnEcU0LhXs54r2tlhgNyqOb4IolWLzefkCG9LqcksLxyIvY6jjUbwlHPeO+u2ev
U1Thp7VROR2Wo88m6e/DllYpjDx09ZBNQw0W2idrnQlsDm2wyioryCHhIGPoW/kt
6Frba4hlh1iTsWyOeDjxMOMpYY5iuolD2SpDNHYToKMkqglrdKfKKypc0Oji1f1d
vMEu6PRXzq69rNV8Ib263yrvsq226xAPne/fBAdXh8JKDBsjnKo/UiiNn8urU+76
c/AE3OnVf8J06shfS50p4kjWfuj2hXO062ISWxymf4dDlaF+1WjNbM20xeB0F/iu
qj4bB+Uwrkt5WO0CzyQS3zwc3gjwOLn0H1EkTWXTLB3lNd2SlI2fi0qPzxBPmdlX
BPMFrcCMOqH+fqjJ3a1nyF1EvxU0qkGZlhA70URDOYDimVigNMn8wgjXwTVK96Jx
pQT5L+555kUv6PmORAanieFSaqNRMMLe9ZL0o6rQdZc53doKpVB/CxtK3s+WgTSe
1CIcICM/bfvxIJRQ+pHj9qRR8dJMrrZla/HABd0D124F5YqVCTIoZ60QO1iZaWTA
WRuQKkzbu49tjjk4/3bpVzlZmskZqTPMA2/v/HwpH0QY9aQyQgqYImOmo8vID90U
joo2AKs7JhsbF9NqYqjG/NJEz0xsbMqZVOx+bmPa54tnJ01CuIBVLoNN+8DrpoYj
5JkNIb703NQi+kQ55KvCge6qITth9Y57aPYBUeIarI+7JGS8E4W9yHga3PH5f2Kp
L6Wzqm9EmoOzXzJrqconhfuZr9yUGA9Ic/+Mjih8cO4PIV0NKn60Xde4BAk13bv7
8KRMpFN8L23/D8/OclOBHz1YWKrGsn0X5Z/J726m5Q+vTEVbYhBIo7N3cYJwOZQj
Y2d55+o5zRHPrZ43Le1xI4WuHwt25MENSgBLLKNbUlV61WGY/ozkDeGh+hyRINUL
VThH8iNuytg4I2uvvmj/kj4kkzTShtzKDRLeKk74g6I++kDGVYBH8netpsKQDkQz
45ktKWtbVISYW89uHcswBpRSAEorrEKn1FB0sLPxljbi/msHVEG+TiozUfo2e7E1
rf1NZE6DQIrmg3qujaVnuNpFrJ8jl5Tkp24ADiya0YtOaYNQmnOVkkrXosgxUZGh
kTFQolr5EsW64sVQa7nkviSYFl3VFetAGXWNN4XNM9rqR9j0lDiG7pg/ZDxBSRds
APzsTBlgNnRDNsh3YSLXA+Buk9KwQftpFz+7vDaekYl0soQIhBvc1YYQQgaSV8xe
2D9bbGwrc296Qc8QXKeHHZTGv3Laz2YaRYroWIzv1Jl9t7IYbYw32tulLiDcWhfD
yeQP4w7BXjbuouzxkGm4BTnZoPJHUI5YIhoabS7MLEr9Rn+qeU2jKqrnEs7CGdHq
xSPYRqmCLadtizvp6ltp54LyhYlCL7rfv46LaR0auHOqW0dinanhRbXgG9c5aW+A
di1eRfusR4IV4BNxu/EnRCTannD1SftSNecjSoHBQLPor98lAPYHVvRi8HluJQcy
+rPgaTVpxgYZYi6TcGDc06Y+Tu7qzVDD7vp9kbqQMTilC0mbHQ/2DzFbkX/5X4v7
r1htw4BsNqiufw9Hykrs6uOIpuHQWJ+n8xHsxZal+HUV9ZRlr6eh5vgtVe8xu7PP
ZFPVp35kX9D/lLICrb6X2lLfs5PuRaq4i6UdHMyOZ+dKbChK/wJyCF+okrZ/fa7e
X8BuIDakb2EmTUBl4P2j0EHb4oiz/AjcA9RM8T/HpJZrews2RiqE34BTNWPRKKmB
77/r77YTraxDha0+8AbbW1xSnaO9UeTfaUxdQUvNVCffehBpZtVqAbiTu8SIWXKb
1Vvh/VLiJwTBZSoj300lF2Vf4fHMV1NBbeOfoq7TrJ0RIhnzpMPsqAvF1l18mmy/
8hFVHqsA2kqi0OvUfRdPzXH1MsbwZVc+IaH7c85jmEvgGdYAJpeFQVifOZE/L0w6
NsajUIjadY7YdSOZlOzw7LAIAKLTLO0rN0sqsrCs6BzzZfxKzTUx2+U1oFHd2KYf
Ub6buoW0saFIszG0aIB/TM5QpUkX+iEruzH/1CpDb0qHFA2TCmKbGUPhkft1L/qw
noSfgct5RMR36grEccgtCmVQt8+Cia50EvfYMuperV30grF3EOuM5ZdSK1Hg7HpB
7Kb66zf54IE6SX6chHpcDdL5/7w5XtG5YMO2O/zyQmiKHX3rw9HfxmPF7eOe7c6Y
OoKg97Ff0rKZgLxuj3DzSNy//vcFAPXtAbxs7S7S5SGNWIu88IN71eujldbOXYuw
1mA5HNcTRlXOFzJbxe5ywbB5V+pzf8Krn6VLrb5fQ90lEGtWtIxRD05fydULWr8k
215CApUdsxshY/h0EKB5yjLKTussQDa5AuFUlViTLqNQGPUEQpVpTvUIuIB7rru+
j3Y2s0BdG0kCszj0Vs/eT1hZC6kGnQ3bsEKRUIylm85GFk2/PrO095IxAlr/cuQE
iMIZeOhkR5jNqHNKGYUc+BDUreddJF7GFcg4UH36meX7umOIY11uA5db8jOCgw6O
6OUZL7B2I3a9v8lmYTdRQsec+NRiZIbkP5QQdgOsxyOHuApwQ0Ebz5C+lLKoocQ3
oJ+XZi410RxQ/L8QfiiKXsAd6Kews1ray0R2KSefgklabtb6nhuxgLzj08cvRehX
WUot2MwAOp1MowsmMvzOikdfj51tvnuw7fIj+1Ak4T1WZjJ/fTNKAvnfgixQ5qNz
26hLIrv29OyFhrmZBIGOQgFhESMO9Z9oayf0jVMC9jeDFWOQGs7+tSBUfdxWYUhI
SrEyFXA0wQWfpAaJutM0ZXAt0WcNZPyKvkuzCLrT3tWAkZorDVrLBhsWhIVLuD4k
ZeVt+Cp/ykDxVqkkktC9PIK86fvCAa3G7jSDjdb8+EIrL4BdcfgUixsN3IuXfu+p
QsvM51AJOs6HHfBhx70HVIodAzn+foQH+onANHAS6Tzo7iUyfZbPgEnijcn8VJVt
SnS3OuxRYYKipHOLY3kVK5BmNJFhHTNNGZefeOV9x1ExNNajPQaKsIITFECFAZC0
05tWMCPYQh0gwX40R/RkWoUEQnnoiook+zQpblH393DbX2q13ncOERPzP6jdABIZ
rIp6GzQu7zy6d/W7rtH7EkUu9qQ62skzJkHlKU6N9VndAu1rnASavMiW2KLwJ03K
zAzQe0yj803maJfx8cqJbVb/jLEGJAZkJjGNidkOeCm2Ap6eCbqW8xFcJ3ZQ4v9b
XfQ28NqeMd9t6/gTVV1J8MSCYrsF+fY2gOQkVHFx2UKMK/KiRcseBBZxIhgLtPJI
ktzaxPVQ1nSVEArCVe2t10SIggbj8IjJ1I1zUO1uDYmB71xT2puTsK1MRHMlzKJT
7ZPd9HVgpum5amFkgGOCytH0sLZQtEOdofaTCQLD2kZiAfzhOMrIAvwD6S8uN+My
XZ9pfC4hkMjStsyoI4ynOgCBGZxwuWVwo7oda5FkSQckcg8tUa+z8nwMx5NaeV2X
TGXI7B1TNx4AJfIeRckqNZgsJ/RO1+cIbg/dukeZkrAvgE/4EXhGke7JIfi75EoP
8m0U5VbZML0N2a0jUQibXzHbtIsGZrLm6KpWLYjPBfj7wHLXVHFRhSU0S0/1XaSd
u7RoJBWJF1nO8FvZES33DaU2vBvtLoP7+CYykJlP9anU35o/65XQ+wNxXbjzeQ1S
U4dACa1dd9BHtpsVmle9iTkkVVMxlX4vH6KA3KwHm6ANPbUFpBGEUXVVZ8v0pc7l
ZAX/iMT/tIZosevEaNrRMXX6XFL25DM3Jn6BLq3HvodY1b94scbDkh6gi/bwoX2J
8HMmW78aTaMU5/XQDbZRCp/5jL9FjVmxvNb1WmTsKvk1T1m1mM1110qciiYVdzGH
DsrpK6wh0yRJGChLaRWp4OhSRfXwwRnWqZ7zk/l6k28b4r+lyavPmga5n0YRzUqx
3nGrkSva8VzDdar6q/8ErYr+kqeRPj20YKxXOlrWRgAXxHm7MVlb0yo1UPA7r/vd
FepTZHEcv/NHMheXzUzLDLpyFkHawchlWSc4sJOqWfZ0xOmuT6ozr9NxA/8gHU63
MF2N7PI4Qgrnr+JgFB01sT0RQlDz9Hvebi3i6vPXmm9yVyTljq5fOsdquDDvO5Po
nQjHF8PlFlUC8xc5OlrRT98oDe/W1/RiUIGDMZLcEgXBYZZVLQ1Cor9AeTQDF4gP
vdKBw0GbEcMQAPNV6RSilZbBXh+HasRJ5unyI+X569DpKaCttd5i2TQNLPprr4U7
DXOITTPPfTydYMAZY1ytHXuJNsnxoLD6pw3NT68NTj4aG8knGxwCpVhGbmiReZpM
rIvg2ZKnZZMK0p8kfq0e/RIKjM6Ps8HxrMjciy/WP0CWVKLkz0Ywpnaa01FxYcjQ
a+isJRmChHCDUlr5vd7cR9GXeoSMJMIOSyEaM15baB5Kri9N6hOEHIQ6tkCFc9LE
OFjXyvzuSdPeaO1yB7UikK1Ijt2t5sNWQ8MI/WMYIktqb4c6E6MUxYkLU5WOihyq
KESUSxCxp16t+CMFCowldL2EIUKPDbGd/BehMTRW5wjHxnp9aWTFilkW5hsivIgC
qGJ0XbeYPrf1khykKSN6M1GRUwudcXGLXJtE1nf5gm1tS9AKhLthhmFAtrS8cHz4
3LxeP7jHh4lqQfO8n/f+qeKqerKkzUejUbcR6e23D/Gy0bruN0cjcg+3xeTX1amP
/ppQlHV2lu/hcB36izxeAwTCKUEmC48BxAKwJmxSOPA1UrJsKO3aP56prj/heCN7
m3Uf1r1dchdrFwKsS5fAAFE2rsLqb46ZKbABDz+4gGIXBkbow/Pai7qSLen9UaeB
/DTZkDfZ5IIGK8WYftg93v+pTrbUo3BC+jx7p7ZupCbA9VyKeR23E0CRN9iDpCUq
qczjRrG3tAJBhuryphlElk3tnm6fyhYjIJvuL/Y88wohCADBPMCziuDAGrT2tBUQ
DOw31fpK1FDbAiOZYF42EPBau+kGEOnHICwkPZx1+QqR4HVQgQ3zXR/QEnchjSNI
N3hOWfROZR2VaJyOBzjH/81TFccJPT1zNKOfTW8i7Fvld0n2Q0HgeXcxvzn51Lmz
THidVMAB8ZMEqDzmwRkitT3SOrjl8iVIdROuNQdEyDeJVmjg5QOVE0BytGQ0LeJq
qkTathmVaIaZUHYXjGdBxbWcpP0ZA+J23X+UvyN+4yc8jeZhrwnVMC6IgyZuqMrT
TQEN6vkhPBLY3qNETKLEALejuQefEfM4Ei2BVEcwEzKbtoyBwRpeepmiSrlWVXqJ
tL7B74ydc4HZLMg3gWmME32oJWC+64VQq1eWvsKTNzvhhVXXRhlz2bXqEKsJph7U
D92gGOfkaMV2kKgeuJap9NB4v2EIcnHv0XXCgZd4eSPPCqRwU7mIjiKxZdLCe/oq
o+in54s4DuAhdFbOmpRh5eFK5DUMSgyM9DZfZcb2BAKkLLsbn4XJWJaBAB4Hj8ft
R7KKCBwlFnO/ORelWb3Rdoqvx8aaBRVswR9Sw5GjPAVSCoiz8sNwvhrWt0zq1c3m
fUu/HcXI0887CTSQBPf2XTk8npeNd51XgwN4mYFjJBeqOl+GPv28PmUD0TnnWrdm
UDV3+qaE3c1mI/Rk6Wa8V7wMAtXXBKAn/5BMwleditIxS0LC4zhNNGCkwXPyqWhz
L3AOJ+LJ63+q5TQuknIoiiUuCRN9PRiuyY5Bc8rlfePUbZlzXHLVn7ppQhChBaDw
K86YBYM1BN2KMGI9Cx/+wikQtlMAjnwuftmXB5WeeaM3ie90SHEeaH/HT3X3KvGA
X9Js3I2yL0VZ6AhkQVLoRRAmIwRdr1UXKQEYrjMQ7RggM0yLEYZmIyxwts3g7pyz
lGEKLIEoHDhhmwh3Hng7exPFxCykT4lXMuDlaNnwIFXo06DPda63BXrpQtR6Ncx5
ZqP48XbscTlAEepuk/IMYoWSIlz2Unam35sVQE4CzKPFN03yvnExytOYTj9/QRWT
1s53IeLsgSQdzlRAWtYaqMc3uAhKR7OENBBvHYo0h7CXKvcJ+3kK+A/Kylysif0d
cDW6jeH+UpOrdCIeU+QRbvPPjQ12s4NhpKECWB04QONZ/I1UYXp98dbUCiW5RHiU
Zbavtr+/RwRODqFhc/f39fMjhJBWTRfoDGGhMUjsQR59qNqXrZ9c9s8YkLOng1H9
1VJhSKf4l5U5bUh5+9RMZxPtEaoyNiYmutMukZf8EFHossAKz36Ix6xRzXwbPydc
POFqYaJPIp5k4uhMSSQ0nOz7YxIlNH0ymAzv+fQioHWSym0TjkOT07lTAaLJvDIY
hzJXJwqCz0pRaERntmH+D9e1OswJJrczXy40I39jajBcpWx0OvlgsyS702p3tzLb
duf/M1QMnxLUsowugeckVbSpi3E07g8wpyqkp/1979C60BhSWQ/aHet2cLHMLWbo
V0FcVm3DJpdxVgLMJQf40Pb5pu5JUxWVo+LRu6aTMcLYqq20eUIxpTaUQcgPQV33
t+y48LuN5Yxr2kFUn9/3cWSvB8MaZex4Yu2NvEOGqNyFupWvROJi+WcsRGWMsNMm
Is5DlCeIPg9fCCp9e2pmYgXGoLITtj22R4kUNcn7eLV/EeoEB8OVONopqtyZ0n8j
vVdEStnfEdGcTBWJFiDfBHAAChs7f1V4+/tvTbwV2g/x808Viia7n5JRIoHYTkrk
3GTyPs7AxdGfDegs9UGy14fVnV0AOYFYVzq8c4NugIZYR/K1zrY5r7dxyDkCIn3Y
KwGZciFHzuaaxI7fzyxwN1gPqEmxIrdBThq0HKylNJFvemHZ9kC83kVi2PBgsq3T
XU2gTVEljI0wfqZVuLEfF05PA1EMmo1ZZZ8Rwu1D5MCz8aV/R8ozH6wlapyYmtHJ
VGYa8yxWHklOYMI+kd2AXkwHgOo/aJZnRSI+IIHExwCOtQgUj0Dt7LaHxqun9YPM
BJgdqO8R3pLPDECY+/c11waYznWqwDPpooS9+6UO3woeLkLdlH0sEEUn1mRo9FXp
mkMl6sIzpzgvnBMj2qJhL4/VHyZDuWBxeEzT/U3xE8fRwbjloim8aCLb8e0SgoKI
Y3/Yl65qtrNX6xqB1ihSeqYOiH1ooLcDtaRsrK6yt9UswZsDQJ8Y/MIyAu+Zimj8
YT7SvOaIQczuKkF1yeLfo3pEGcgCy00i+knccgfPYYB6Pwl/sQ6cwmAjMp79ex3R
xbdLHVk9XJGL1th3CAF8ekAgieINB7pMRJ4FNRtcrK5QzJC01rmESwL1TTwlxiHw
RW9rZkKDArjjyh+VZNVmSMKPFv9iTptNFe4DQ54+4zJfqStjP4kg10vXcewKlued
3Lh8num4p6EMPJz7/i/+MHStrmrdPxzPdV71w/7UxZTyw+nAbwBoliwldSz//FBA
8ac2TYw8bfLH2OjJuk9R/O2d+1ZhZ/jDpwEZfEFpY3wXkssxbt8rLRuoeHvbtxoK
PQ7+eClUn/SLMTrz9NCPgmD7QFloaYcqnIl/hCin81jMm7HaTstIibdrDeFvhi9Y
g0uUX49v0KQtvPfHNTivLBKurM6Z8QprCA05jBX3en7tTGovcSCeO2p6LdN+WQDr
pBbuofCPn4ZAm0d9o+Fyqx3DH7AQIapT/IZgtuxyxqcE3HqR7CSXhXBKMCx0c7gI
REvTI06n7e3ykolBWZHdCyAFvhJt6rsTr8Kgda8Ut0TzHaRTPJhj2ed4EMxsMd9U
a6cGbotUoat5MXbou+4LJZS9j6deA+EENHDZcUDr0bPT6D3e/MwFqDoxt1Dsaa/Q
gyKfBkDXH6Z+qT4O3lHdp+FOMdkCob/zu787t/m2HtFC3S8whnbIi4KeMbjfcUtZ
ju3ARfL8ky6rsdwGXS1g8d+Ly1DxWsfYRJc+mvzqMHCoSZEyPUJyAjKi+Od/L+ds
epT14vQyiOLWzAWtCws7mZKUbmS8k8iYM5BVrDZqkmVnE5Eh9zGYlEB2a5L/M/9B
wgWEk+7EpKvSrdVqCX/djzW/xz3R2jXheqrAKGL+LW7H5eq+hbfl3d+1brbp8mwv
VR95vw3FgJpVD1RCD+xrMo9yoM7DT+IbbaM9APGKBdH0tw5v9920LGp8jl4fnTWP
T0wxhnRrw+h8BO+2fqSktiCCiCfWduPZpkUKsbvbgmb8RC/dmoPd6VyR+X+IQw4k
9HKFVf1iS0P6cTmqY6YWDRTmf+ZLpyLXQ1KNNLnS1TLO8pexh9PvncqaXZHrv6CA
JprBJr7zwPqsmXVNob2yb6ooSIFwC95aFOFhVT2PmHaksMQNW8WfIjK/tQqFAwFB
7X9xXwdm8Pk1mshYfcmtE+TwpPyrpSbPPGC/4LdB5cxjc87LGLCKx1maMAkuLSkT
f0oYT5T/jXLYrEkCxFI0tcBx7Gq8XbWA/sfiRPa7rDu+HRsJHUJbJ9/f8Z3tIo+x
hjgF+DMyKKL5WVziXUNRYCGQKJJyGwqVrU/nGaH7pPLlGQlW2UgQ/GCjYTy/Z2QM
XRhxQORATlFey4kuroX3LXWchdmIIO2264sY6zGEhVXdTPzBRIdCJvn3atr/CO07
DmcbmmuDw7cHDxzhcS+bm7zJA4toTHp8ekuMx5BrV2GmQctxUwzZF8t6OksCdggr
FwyDlo+UuvCnzZLfLsrSZn/Heii9gCWsiWkCN+T1NDjHlYdcA9jHYj2aa1swrE3S
Bcl/onMpFi4NRKTGHqDGo6edIAq7NfvwVtEFP2L+3UFP3jwDJ89LZeQ+e3VMwYkX
ZY2I9+S/5zum3sUnq4WtmYaz0sHdwXaqy07IOgiao+vQf8RdiT6kl7L79P4B6xgK
z0LNW1Lph0gi8faULvXWBj4HDkE2yjs4trzMj57Enfl2M57zPxkH9OwP/5Zhp7Ub
dMoBtS8NccepUIxFEEs9zbabnW3bd3Z2gthwPcATU+SvXCDQ1O8R62BX5ML/K1qT
Wm4QqTyu/ziJPdK8MTzcp5J+M9GxqccX1O27XnWEjfsneLWym2IBVqYyXoJMhrRb
oIsHWdC0Blypfyl4AHhVK/bJhkbQaBLv69ye+NpplwrRNmaw3ipvoHt2LgzHZrWL
28dwD18VhWrIb2pDTuzH+D9A5mMYIupZtcjxvs2UzWrqlqf3l5lrOj+35NyHKa7W
CZZhKlD1XSo8LzPwYmWxJ6+1PQfspb8RoLVQO/fssNsx8Rmw2TyWz4MI8qXg5zHl
zgWscnmwzZjxvaiHPKp5FvpNPKZ1MSYL0lIla6dJfff3ovThYNyJg9R56ZHbXNXJ
nCzg/29EBheoOBg2aBYmLQ3JorBTpAzPOXCyCazpadUqyJXszIzQgR/H3NxNaHOn
CAa+BdylNUraxZerUFmXugcbNdZvQbRPvZR8J1IzPguePYQ0fm5sYMAD0QSiVdGU
MqkL9i3JwTjx2cs/4orQoNcDeAdeY17YicKy4YobprW7PTF210NucElu/Y7Cd0Q4
PJeQbGC5GYj3rgmxvzVgoFsHan7QQnFe+E4DBAug9bPYU0kuxjSGrv6FE3a/Wk9H
gkQ5IcIyeo9H8YWcZNjunTFJ2lOIJ6rHOk2kIPIZeqFDjS7EL8o9Crx/VJg5XBly
YH9iRoplEVHPVIxcJ/VD6rXcYziLgriOkgdv28vpa8YOgVFGsAs/4QexzoJAwKfl
t8InGBNIEzLD275h7ml6yTnDhtVuauAWEouZugjiCePB98DgcIbg5bfHtbNzHMzw
M8+q9ulZXHkOlWaaJkBSWvGjBhO0srcq+BQZcgEKz4zlZgKDfRipCgmCBC3n2XPN
3qae071FcKPT8MumSBd6NBRDGB0Gn7gc6wGHWElWzBdU/VcXhAKVp6IMiKGZMVY8
Ncja0Y3bI+8TZnqikfFelX7flBAdPbrUjrRiBku2rRuS/M3HD/MHULJdWI+cwx4A
asrahHA9REgfa+kWmR4im7azTsP4ddDmgH43cm3FUMAZJrI/ZY5fxF2gNKmrEeyp
5xKjEeWCaw32Gdn7ZMOLyznrrKyHW5S85cr5oTwxqnkOUlIigZ8eoTAO6SgV66mG
kDcCDv7u0VIbq/jWaEah6nV+oooBohgghjOnD5DncOFBGoLyprDPorgM1ujOv0DH
YEJaeWUxnFBOkuTNFT+bML/l1G4pSUcY91QCrdffCUyB3lX3SaqyoILvF57d+g6w
KHieVwxsSY8jCBqdJQm81ulLFBMJJibbH4+CZwPLx8b7xou3NjdSs9kOGwzOLROH
czT+gzaF/10KjKXt6QNbGMxysEdyG20ulnHAOO05QoGlKv6BR9aZ4kH1tvUV1yc8
hnSLFWl1GyiFx+kn9ceq05JfJ3HzubZuRq46rUVq4cplcGf6ZyQ5DKRfCbsjZpiV
j79y4SOmgiVEBqQY85t61UMp7WR9gf9XJ6L+mcK8qmus3shel4ae5C8ksvRvjECH
bw6lbVMkPX0TGQc76gQnQLNdSwRM3NK251uVP0RWQlS5+IK+Vqi+/bVU2SSGZNho
gkI6rzpnoXlYjG5zOqNLt7E7Jn2Cl7q7uTiua2gQH3ev1e7vSitMMMTgdp7l41jM
po7zmD0jzXz9Tkwq0ViCMnIyKWFcEq4qRSHoLGxczJIcifdhqAIUL6o+NR9GaKOp
uolFNaMVtwzgNFCS7EcP+1ZkdgF3txNJBIyQY1RvITzksK30O3ceNXb46neFNy+7
2DMGFO2MYpNRNEo+aEwLCWhyUOLk6L7R+9cF0F2KLwcpEfq3HYgZ1xpJc+JkEJRH
j/1pr3MpRZ6EgZdAOQkjHzQCMvVwYzTZ2hIA8F6lcc3REUZKGqChFb5WSLP802Mo
c6wX4D2pP62Ne/R4Yia0QVIjJZpmLlkcqDzSLzm3sMWhIrQqI0ipf6iplI00uUZG
HW3j8RTzVLl9iY5noMT1i4g3Ssfb7f32a1Xn37kezMpEj8dFfe4Y41G+iwlGk97c
joo3kmcVtK2/b5lxkKyZg4VGNz+e+NKJk2/k168IaAcfoSVMHzKPrvrRdwFb2w2S
w18874LXirxallvHO+iPczD2LtEBicJY98hbLJjj9LS+GDbbT27eAw4fcin9TKqB
Xm1+wKAIB6qVB3kvT/F1mdLnkWxz7cZ7QElIxdoDv4w3AGdv7z+RrGMrthx8lkJZ
F3t3nJejnGON5mPd//E+OV4WE+6yOA4IL4bGRSQImjV83hhL6XxYOH0SRbRDUNec
gYKwINoigK4nsqHTQmdSjQ2IJ4MAjuwm1iaxs8KgfwCuOzQ+j5RAP5cV1QFNFKsp
D31kwLt4LNzjwBRNOx5wgKPmTHn/cCsvpJG0763dva5ydmB+LO2S3qOk4kn/50YB
2doJvdpxJZtY/FdVMd9rbKZpw+wAw2oy7D48jHsLm8vlz6010f/L7V0gI4bZr5/N
7cvAmqvNhFmDRXzaS+Jy0kWovWR9l3GbWOjfTbP/IXQZVMjJ42l3LcPEkB2odGSZ
4268G+tQInObW6ESpWFwxpewhQssq1x9CnCEOCj8iUUCBEws6d01QVLls2C/XNo0
BCfAwOiBPUwus4JXARsSpHEBZ2YYwJg2BAvL+96/i+eVio3nEROq7EVVHIay3Pj+
mNYKHQ6IbRqQI5MpQIKLz1wJoHrN1xstOulGlNoO1HMmx7FZG2nEEoh36ZOHg6iK
khjj03EUDu6HKzZ5YkSKqs4B7b+iZOjN1gmaunZYthnUwNoxarfXsKYe1cR6KuNF
gCvjYD/kAaFz/z1FRDJcM22BTPn/MhA2EdB63af8GUDG/GnWhJY1MzHndRbftbF8
+6FjhqLOFinWw4vu/an19ZAtVOVGHcY2hui2OQ1r9Jndp0z7JNOfVmh9OvHzrcfG
BoIOrnvd34Eq0Lf+zkbZHYw4rDzZJzgMY/+ZN8HxP1mymJ4sG85iZPbbAmiCzRij
xHR1T4+x5sqdiEetmEA0LpUVACwJ/2ZmKrtB7R8e//fFGgOG3X0R+LeIAZOxd/lZ
q/6IG3jiVcCxofApPl5SK8lClLTk5Wwt7FpBO9MLwNImiu4C+JKcKXrsmTjA45nH
sVuNDH6adR8yNtvTvQulahT03PBLAVtaBTF3XY3LgX0IbUzDqswrE48jClzjSE8o
cYLrXIxG9ZcZCzycXvkLDLeArNTvLFMiKou4CpDBVLiDrTd57M3rzzdWFkWuQcLR
d4VklJpsX9utyngvH91BT2GB0wsP+tYkVbkGgoat7urmqLdVNeh7weK+Pd0/UjeD
ixJPdB/OLOFFZ2/l95iTt82DjLBz9DM5g1isDHhESU0D2iLPHIYsK75vQ06vVxP7
5MjG0VMRlJ0i3czCLzwejTSnfCGSxH9oarAjw3E7P/ZbAAq22wqL7JvsW5zOxiEy
zbvEmDheAI6yBY8/TvYZK3c7Ob57s9r5jyea5GONfg0v9E+fPH/LKTFQfjRC4WWF
k5e7C+Lf1BRRfv4WPIA9BRXbm/NSb5oGgPlWJW4uL3qDxIAiS5Ng2HVJgl3bGXlP
Cl1wSksZDaP7MHzdC4meiLCGjunru1mqTmN7P0E8mcTwCkQY6EcidXf4uSVJpEWb
9RUFob4SjnU+3iBvutEtdNgq/KkuXkK384wL1YRxH5+RaLTi26d7wsnWzNWhF5FR
f1LOcqI92+e7XPqYTIWYWTvAXK74G30raH+lHrQgrlM9JOxhaevxwdoax9rNQ7hl
LpK6A/0GWKDZOMc7VmBvmQoZSluTCbD7MCyX5ITvyD7Ld8iwvpbtTt6DsAQ42y+U
M7XLH5thPIGuN0IMoKQeI0DC3hJr+rkxPuBojV6+PHG2T77tMLAbQ3PFZybGEeJ1
BCtNwRq7aVHWy6jVR/+d09FOB1o8WOFGfUAiGW4wqahW5VyK0/PGyly+L/UC5YiM
oo859S9kkaBq4FFSLIicWrWEMoVRksfNWv6wgM6ERTC5eabE9rgQhsddo0C/vxCu
6j5P7jgVP0pt9zsWSV3BA5HR2fTLLSFhK9UTfawuIrQmwS4DDe8XeLQB61RCwSt/
QOxK1XN1zccbWtcgk8RaKRJRKcoh82Y9zpCO7KcPu2vCvOCBZs5yTM+1Y3yLr46O
yqBSh6yKB/2+65/zPpvgPqgafmf7KRF7sUTtPvCw8od46nRexZVTO29VpntNTG7q
QUyM7vaHOsxwlokGctdSsBT47F99EV1dr0AWf4vxfHJlmr4vY3+GpMsU9WgG9FJV
++4h5M7nPC2EkrVe6rCPueZZhNPfgAZJzzDrMw1LjyxyeYCL0G97HIrJ5CbPDTCe
uwFPWV5rzYbSdsosQsg7UVvLuFL/V9tT1CZqDt2Kef0XiM8fguaBoHFsmlKIaN6D
h43Dtk4vlTDskDS7VtvdcD4BMqMK8H85ogKqGDupgL9uFDxGn+PjO6aGUXLVYrtJ
86LEf9AJPyvf/TYTbIP9q2JPGlCzhNUWfmHZ8wk+VFGjtk7yHFdFYiV7Ip18CbOO
AJKSZDTpEw7vJ0qZ9wmhJaprnqFPSGyOuUINYk8sXocXFk2U1a2mtZZYg+EBmZJy
Ky4/GlKbxJRuEqrC9a6RGBAuFA3nv+C+C9VbMJyPzRGQI5EJfK4T5lJR7p53A5RC
pjEFRrbITy7vHSV2sJPls0RBFXRrr0N7REeZ+M7Z6/oZZSrc0UHB4s7G6W7b9b+b
B1uTWzZO7LxE6AFKOgswkKE4cJWQiSfXZQUIP33S59BzqmfW8YbB1VEGi5pcRaRS
Iczzml8FGYBHAoOGtzvPEU+FUfdL1idunph3AAzcwhWnfiSP4lZxWTbSqEQ4M23Y
7mKN8tk5RR8Ecu1Ert7M4KiUK4ub00fkz/41oMK6OdrhRX4QYAsEbL3x+LKLl91y
JXQzhwWdLF0GGfh2ZLVB41wb6IS14uRjC/o4hIbeTlbE9cZ5Izm59TJPT/Dk0GKv
OWjbmhkbIBX/wE9cf5iPXjBSIX5axXH9Mv7F7XlDj/m3N5Fw6l7y9hmVexNg/S7/
47GkFvBtv2oaBuSgGor4BZGQfhPshrD+4G7tZwCHJBCb0L+Tr3t10z0lYNZ6fd17
GCzO1qvENDAIGNwvQrWSJQXptVo0izT6BualZ3eOveJsdl3Vkge95MsTtY2BTdf3
nbk9Dx1gr2sj2c5AkXEdxyVxcD3LK8IRgCneT+wFt/4+Cwrme9XZ+lH1UxN/Sott
MdpN5nTEwQF3MXt8Z2eC6Ko9SpI4v85vZ72EYa9pxAZNn5qO3a+Paw5iRWFZagYq
+TtVwCHFDfm4bFHFwtdv39jxyvF4I7++gMdVmLQwkq1M9QilscsiaCeM5j8QLPrw
a9Eu8kDp84Dw405QkE5TzmQwT2x81nQocLY9vHRbu+8SVorGVTktGZ1lOu93HmH2
Fj/gEuH7GhAgiJ/nffS8JzLTo+dXPHDGWUTinzGrDW6mO9CMfGLSAmh7YHYBlOeu
aVKY6a1laR5rV3dLVfD9B0skpvYa9GmQqfJiozhrxF3VMxcU5FqzGo3qPsKbCOCd
ckOpQNuBKw62cuN7mYorQCauTJaZc8R1Tnj2P2d97sc08Llmr4eqahMkdwszcJ1+
bqNVj6fp2Xu+f1KKtuPwexhNYssQ9LTNLD4h5rpMGvTlcdpB11ZJYWcB9SZXTO13
sXppVuy5oY5FCWRgSzOU3/GbPOjydaG0MC0JnlaVlVOIYOjbXDtvc6TVNY3vo6jY
/oYjvxkh4Rv5d6VrsqCyT3N/SWnDiLYe6ChnFJR+TGKJ0PyhbLFPVT+fogWx2yYh
m1zvgcm73pXGc509TMdTLk9tXXj97tgL4W5QsxJsVPqz/d7SG0mn2gJKALzJ2QP/
gcsc1Y+JWFGEqkSdaxMFLGc2ktagvQBIYLjFMblHbmFkIzruxfg/wnpTo/u5ZXDd
6PWHXh8wpQbhQNzM5TTcpxXMNYDxHknxwYRuvYF64gOjRAPrjzxzxrvX+gCiUMFt
hN0eoPoRpwGg2ZgBjy6FawYXBlrB3PWpWI+0WNmDerFSPOigLoamUf0JQpj3UYIX
tsEuh8i/1zMwVGQxIHTIF1XExXEmN5v6aNGziePzAYJlLEJYds4rF0dEbQKTvCQi
kiyFPxeo3cKWet9TxFcqFut1V3+e0PHDvlMx5apVPs/O0vWkLqlYV0HPq6l1rjqB
mmHvcImy1AAMuQY3XnPD8wXMxoVF0qi+9x8NnVOLN5RVDMRmKH74xcfn7WATKlf8
CfPtf+8DK5qntCuqo3uafD0DKEoV9wdGDdScavusy9/UeCKdx+L49PQKNMFDf/mq
9ZO0kGEw5zXZjRjyGsv8D3HFWOviaNPgyVgOoED5W9ZtoE6RQzkz1ZR6m/jKmjzr
T9Lo9ynG4zGPZsbNkjJTK6vHIV4gF2pwLutkfsGYZ+ZwZkhenHqPRnfZvxv9cMc/
qTvFsEQW2XcroAPtgQrzgu5PY4d+NvZ41Vw1dpbwBebvoIEvH6YLCOH/yvAUPlFU
bKZzgpwXstaOo6zdrCgA3Lp2Hpo3d4XMlwWWaA0xy+XRJ1KVLixTJgYDlOJQhY+p
R0Y8AbYs7Qlt08rx4Y6vbu/JfOrc33yE4G6kTH2jhK9/Dvb6LKETfV1pZFErbMLU
f2Vu0g0PPcBiq4A3UlBlkkjP571et9Ew4bEX1jeWiRpCLcBr6rRj7U/mA97qupmv
AfDIJDY8e9G2pM5R9VebFkV47CScmxOleIAlutnxDbqSr9+Vby33FgjhZNLtQWkC
kjRN5U1Zh0m5SnUhu4CSED7gYHFvFd+H6YrATmt8eaBPGS6Gur9RugyPQOkBKZjm
mYfxfpn/DKfv6FMxg/Eg/UX4N1dbYBOEvSVRHMaKXfnelXHYP/5u/BXUCknwJNMd
ItIAPLgUumNC6fB4Xx4h119izlvktKKahNt7HxdZvOevISXkcFPKq1VjoeC8sFS0
4dmTf3mxD1NyXs+YIIdFS/HfKJJpVhs5dJ+kFrvnMmZatBkRx+XBUo7gkfYiCMaZ
evZ7BheEuYB9WYJgCcOAM3cay/MWxADb3C1qgePS5UpfP5EhCl1YwxtvBqHR3oRZ
mMkrAw2C/FQKjwI2OuT+F5mFELJImy7n5FVptClnqSwvGvQbPtOZYMZOOMEqxitz
+KU4qrwOLUJhDeqXMIbaGbykfMSlmiPASKzoit+HdX/+I2N0qV4ZVqJJkZM0hcEc
91EE+3qtQY56kv5jcWNgYw0Uv4O2ym4qFwdfztg+Uy7AygDLz/8GGlhuYSL3tM/I
scO+BD7XIzidj37NvA8nTi5S0yYMDAtrVQheTl+oNNMRYogJCPhpz9NuktREigfL
r8aAhsbeOggMSwhTSdyfwjF6SGO0yiL3lESfn9Pq3o1OR3pBzArnT0BTV2PN1f1p
DhRPRRsn1JHyv3OwUctT9o8L9u6orMCejoQn6dGz/D+Ha1QNwzCBmRzLMPanjNls
aIUZi9cFugwMtZXm+2n/9q6AQheKJReeW970xKCOOZGwbcJ4bHLhINzdsW96XqBX
CoD/JoRGNcHxW5Jz2noFB6LoP4Pw5og3i3Tu3L6Tbn7tce3QYGa3m/4oTffRdyXo
yWXnisjqK/QY3pXUo8rT993UqoqLffYElJ4pKAwP93Q88yLuHyk29+CDo5H9waA9
EYF/ADyjLdKbW/sZWB9CM7BJonNWxjxcVh/UwEXg+M554YtYRsXNVQn00xh4DcF8
twK9nID2NLm2Kassxaz6L2cWPfK06irW8h6D5FDegX0ANmnQeZk1z0coxPRlIXEe
KAf/LOJR1v/GDDtoCn2TtGIhvQ6/gY4HlQvYLbqUKD4+DfY3RlzI/KO21m7AKb+h
5cl8i2pMSap27TkhzDaPRMLFa11wXgY3UJluEYR9Yjn9RoXE4m94Kw0JZY9sXCB/
k2u4wO4MGz9B8tvyUMJ6fnnSyQ8LfGhxzA8s+kqYrn0gu9pd9tofeDfd/G+quB64
d5wFntannB8jJloMCGwDZFhOTK3fBwhir3yMHfwOVg9CJxTDbOS4iZTu13aQLk7M
uBfUKg4g6Q6dZhQoMFrvWk2SWDFQHHbC8szmlqLXGt8MrKy1VFKheO1aFYn0ThuN
fPiFhupQQcC0FXKJ4JffjltcoZmAlClTL+o43cAHtlFOXQeFk2cx4eHZwNqGi7Bn
kjMAphGYBlUfEPPkwakFluDRw39J3RZr4RtO8oBPRAmBd4ZWGc91ZdMwwVs9QPez
R/X2LgJQglptBGcU9qoTSVL42ZQEadQfyF3DGF61LB5WxJFBHpTBbwB0MAIX5971
xLOtZ6CP9pkRW3x9EjluxhwwElWC5DPHSOWMRwDNQPVPl88ymkxOCBR8hfAG8kLK
N7Mtbwb24p5F9fh5Jeq10AUSnjsem8kEbwflFHtD69VV24nMbevoScVT+InFUNYy
Ciq7hw6Q2ygmoaLJuC9tMeQrPx+UFmLpjE7JRZSuKOG5YIaHNfhkiZ9h2UUFb0HC
8PpKiFogOU9Gq7TExPHg1SAxBXTBP6uCs+wla1BzECDRw7UQlznZKaZ3XhK55g5T
65LhPMsrOGlckp0img0BBF+kFdTAhrz2gw/O2tcPdCKzXdU5ZNmAqX2NTxrqz+O/
+9Kz1Vr5g3JGBEHYPCrXil9IVx100sUy4Rz7W4kGQl9evcate4DpyanthsmVOcLT
g88ENUVRQPhRDBr6UTlcvNoQRHK7wBQ+MGbDRthasZNYFcUehNvwBYv8yjZ5zzZq
0bqoXqYd2lD4iSFW6plnZ+VGRzzxSG/uTnD5kfacRZA+tCbO+eYobiyTaXmyk6y5
lTyQOxqqe/L27PYi7gT9AZ/2qtgeEXgnrJbq4VWzuodMXek2w81z74OqlrPmuCqk
1LGllCI7f1ohxtG6yMQmhGHRxLbyZdrW1djRr8zVs0ryK+u+OdSY5+FNT5+SZGP6
jCDF4xr2XSAWSfgClG0jtrY3kKUVGcOHwZ17ZcUiPmQ0M7kiF3VVElCIlN3vtIrp
bMK1bTl/naX6imldRxhT/VO/e2iygwKEqEuoF0bLP5z8AdfUQxjab6L/kSQ+rrAp
729+effTqo+3s+qIBldfqBB4pGRRB+m9GpRQoa+aJ8NYS/K7auqbOwmFBbMu7+Y9
ykMH0xV7tHNuibFGtLRfD/mMZvXyRx4gXKOs9V4uDl/Zwnnw+hZBxeA5/bvIf7/S
El7tEa6KmoD0TxnA4lznb/IoxCMa/1cb4/cECYtzNyyaC1qx/U2TvFY3UUvTsBHr
RnA5PxAG+eTDTjXgU9U8ekf6OkxWdo8DepQs9bdMUGiz5BFHFvXIWuC9GtXkswiJ
s5ePi73eVmJ8RhlAEu0OShzpJzzOP440pzZKUO9HjhtmCO5MK5a7yI4mRQTGyq5h
zQXTJwV90aZip/+8F30HbiPw/64lrzr8Bxw+qGCtKGACQxA2F/6yWSskSrBvcZUU
owZ7pKvUUxWVnb8Xk991GNS2Zh5tG7bOMF0QkMs8cCp7p1YNs+VoBPFsfA9Cm/UI
DXf6uDyBzRw9tPh1nAcJE7lDQ36MlBtwD0PF9gKcRRlF1WyOOvIPEL5dMcnoNHJT
wAOM8xReUWbj8kzAeJ8v/vh9eh2btPY9uGC3EW1m27fdFb5czbiKNxSA41PPsi5W
8K5i40D8ROqqS0u9sPkdboLlCq4QyqCIPOOg1k6yZgmHN+ycOMc2TGpZkLiHsCDy
umPx9ypQ+ffN/IZUtotOmEv2My7uQhk4zpk5H2t2dnaEx+Lfei/Y/YkmsCEd/sFU
vxZBtE+YWjyj532piKxPrEq+B+3FdLYkUZpAjUi8m0BVDOdcZywXuglqXq6jnFuq
6NdvWaRyPEUvonPofSqoqCPFBdHHl0ohTDoirQpWB5Dj0Ky+bwT9Ht0zv8oiu/1d
75Vp4vJi0yHnhp2cam9ryiecszyZR2vqqMdygSI1x9/sERqy9Twu1g9fzPHchC4f
fS7k11z4Hn6Dl077stC4YM5XQdj1dxRGUY4sFFYQyt7h/6VOKXDy5WFGUKdBqBf6
ILDc7zQ8KNu31pk4j4hEIFS4Z9ld8ttpnlM6OstZKg2eiimxqEAJcVtCy93Ss6qb
fAuR8lVquM4oJtxIfXyMjLub6jFO/939ESnXe56Vu/FeKrxHoKLuIpL0nwdCKbY8
MulunYh7rhhmm5Sqw2Qc4GnprkoqqYSooiTgLyy03+xtqHvqpgfRT4lIU2y3BvE7
sUrQjILZSMg7wc6LBKTAh0ibhw6aSxmMXgALwg/I6dx2Dm4cvWoFuM2/PtIy92Pb
NmzK4c/+reDlEcIAY/6CdVHtcCzwS5UA/fcnq467LWhR1eIse6lw7gRG9e4htGgW
cdKsKd9mpJe899lIM7g3hkWzfRT44p3SKKOSPXM6qba3llqkxME87Ac0MoFzGfGU
QN+9Pt1H6WuOJmxZwNzuLOWOAAVrT3UO8TpPckjdD8qjbcL9gZd8NN4UXQpBgCgf
OG3xOtF5oipG7b/mVbH7oY4gE7V7IDpC9vBwq9NCnC/To86LpYbamRMYpRkkxAW0
gMiqvntRmS3K+RjJb0JaDZijG8H8rf7ZJ97qETb0jnpFU0qOp+NrKV/zkFhhKI0D
JyxiWQASKuVhgCWPWD6jHcHxj1yJF4xvtorbxffX/97G2YRSiocu+vQ9zqgibiyF
zUt3ZHSBHq3nLvh2oYJgeT63qHDpMFSGPeQUam0lHNMr+D1qrCD6fH+Nx60F9eRB
3IIeGt4Xoh+pivkLXYm8pDzeCvKfwtEYXdUBhfGu4wf1ZSa+EyCKJwke/vlvUsqW
7odNX84Ucf6wPJPTfSLerRYENc102a+Begpp2WjaLgtfyKCQdTcd0/PWGgS2djs/
iE1eW+k8kliGJqkDVEIR79yHR8+7qbqK6wRifyrUhR0+vvOK1VA/3qu9XJIdMFyK
y75nrsAG5+R3R5PrbCcbYa5AP5kfzEOGlOXabvqds+YyMYcAi7kmsoQXTgtMUAgs
OYHyK5zZdC0w7pH7INzuPECa5WGsaVOz0zC9ABr2ER6VIPkXqOBfEsSYAHxibBtZ
xSFe3/I6W9RAG3ScJrhgABugV7WaFJWIB1K68QNDuSkxSAJ6OANE8V533Nk33GS5
lKMClFzSYtjhzvB92nyCLO60MSjK9eRF56FBlnfXXupYFjpWgtXLvd6shJ9NiSSf
hsUyuaxxC42U54Y47r3KZKf1DURWAN0oMo5uS7nYP5OfGdFgKmMKkj2H3SvlYv0T
UZEP11fa/7uzso92paXBUYkTT/WNuspqeZsTc/Wy4y00hEnNYXJb0kZZZCdzTQzP
6tqtZtmd482W6TXhEF93GAv3uPoxzmrTGATiD94xWiroQOp15Se4MxPHJ2qG7Dtx
B00WhNPAvWMa2GcCzxbzWHa5VdtayTeeT0d3DuDpp5oUbbzOUvKfD68NPc3+r1M6
yH3nbU6WFEhO8beUmrModOey/JFijlEdn99MgbLvrnr/wtm5dOsJ+Pi1Cz8XyoYD
wd0eFyJgah4k1QedBVtOGf7hu2rGyWmL/ftRyQpzIUKpwhpaI/T6KYDu+/NykfuJ
/fJqO/QJW6K8ktK50QSqbDrGQQUcp9parC1vBOVCl+ZBKlC36/0v5AzQjdwW9TCj
sPiXFkKsluZfFUn7FK7fQ0Zf9jGIi5UESqOm8QXls5I7DXLepcryiqP4HHqEurSs
bwmXdQRepQ3S3gmzg32hv0ZFaH5iaRnhQb6b/w0FyKTeKo6Xr7vGmVj+d0pzXhQ5
mv/ZJjNiXH0R5M825u4h3AD4EbUmkayeUUjoChsmidGby1u6EDdwJsFKu31Az51w
LX6dHTj/1xzbeIYBXvkF7N6ukzKzbDU/rLyeeykk9/3cdl0URiWd+IMHY1mLbe7h
dkRDGRDHTNwz0b6BkwuSE0TlB9/WwqYlpO4CE8BnvpMrGnapB7B5ntwN7NsI78sh
KH5SG2L7na4IctW2x/UHVNBtvuVP4gDdyqylDlF0lhQr0oa8Y5aY3JS+WUa05U5y
WN5o/OTWUwRqsyDUdpEr52kEGyv1QZCjIM8WIQFli8zIjEWASQo5A+rRCshDfKz1
9Qk0JlSR+VsH/qPvZdU+TfYtV1PS/fen/uFvoHkqVN1fdOvZm3dhWJKSkQVxoVTS
stxs1VYJ/cKbKHAT3oLXkSciKnA7cku+9wda5o17NBAUjVKa0lYpkYXc3YL7GUdR
10Tdc31hjt938Ii/YUNvMsjkwyGQbU1kmp5eqZ7tdQzBL046pTpsmYEBM7hMsIHs
/Nf2ZoMATuUEjh1E0YQhwGsioJCzJ1sqqZ8ocdn1lApX0Tw91wemS2htXXgVbomW
KI6LYRoKQBW7kDxW4t0Cc51foLxFIWNX+IJLQNNOZ58/QH11iuew+z5Bdn//XZjK
lCuZvMAy9HKhCp9dCwrQ8d9tOEumLnisE1iVm9ua/ilMvrwAAsEP0vW/5Ms1YJsC
WLbhCO6eUjx72UinnjkH18cm6s3M7HNo//yjSMK1WZX25BCNj9RfIiA+JynzJ0EP
o3KezJFB38gKwQIVwv8OGPdU0qs52PBk+/HCU/SxtNulQy3Z33TmDTH+k9qfSxfk
FUfLZA6w2wHVTT9JSsIh0pdMT+zYUYN/wXqoSv8BXhzR1HSq64YAyLQwyenuhf4n
Bdp/4gRbXd2hAdx/BDgMXDdzvNaXc/xcb3uHmPA8A75ADLgKNAvEAuaphbjQNePV
zLPYtue83MIUDHSF1lFViPACpMkMyHQeoJslr0FvDVz58mEbe6Os7zVi0YRIOO7L
Omn3S0hfZGi8X8Y7tVJp40jf8VOE4neVh27sFj/1mCB8laYcls5XPJBIO/nDjL6R
UFa2PM46uy4YEqeJOMy38qaRDdno6wHPFNtEcBG1rba9K3AkXIPaqhur8KhrSBdG
qd4yrlqLM3MHv4Yip51EkIHrJXCaY8ODgLNtRuTM356zASKcNvBXvygIUnPBpiLc
CxKoU9RQTtWH+J2doQUXTEBTvyu40l1zH0t5zXPf+I8SBLpmrEZKhMZ4v9nlOk0o
SVLBBgFU5aqX78Fu8z3hH5qeLHVjeQQjjiVzNkzG9NcJK+fxRr+ow4Fh1E4aOpIf
NBeMsdhpf1zzr+FZv/9OuW9+HvdDf4vOEWxWgiOmfGJh+uNgLib+WiINygi2RQP1
JmAKiU+n8lvlOPjJZ32Sre7u4Q4TBBboL+qCyGA4bQpYSSe9zHkGIMfAY1v/nf3u
pfnNpKACjGtcSmgM4pDYjRkp01R3KQxLgBE9tk9JALRx3yPqQTioFdhDO2DN+PBA
mzYnQlhhgAoRVailI6YVOHgI1kc1xsqJ/5W9Ug8mqclvjOKL/NpRsv5PvCQ/NiHB
2Ko1xEcgOzEoe86hATJKg9dNNHU6DuDAx+pG1ivXxRf7m9fNDyK5bmP+v4k9Jq4a
KcMysRarGwl6xwq6P6hl2nGWi5uDCBbv+bYtQ72nj8B47YngBr13z0a3kcnBhFIN
avd83mqxl8ChjF+brHgtuqyUlIatFekKOX57wLqPRw1agdjeVneUPFQ/1XSVDH7u
Rc/MLbyDpK6iHH6A8JKnwsqyH3IkrpBeTpUEAl8EJ7QA5ljh/hxzcei7cTokKd8k
6RPbJSZHoU2SjmkXl8UQxkzirsL+n6bBL9pn+A37rtKHag2v9OeditIjkREU4xQy
J8X9nSlGxHreZcQUQC8NS8LfbxUvg37Pa/Uix9i44tsHGQ/w556sh0rQQt2S5ok5
2H6MfeA4TgEj6FgqsWUJ+8z3kIHENIYWSlmQCDGMFArqUPGx/CpEeIZ7BQx8P5Qz
nBb4l26G31EsjXiIPgMzEP9PbEfU34eXkF8waqfeMj4R4MMSt3zyo/iF6X1MyfKP
X+nhX62N2VMmODEiXsrF+F01npIZKLCGMjeRKbkR7Y2uGq3xh24xeMILGImMdVat
54bQFsbkfuANHviQkuDSj2F0zIlqP/5evUnyZO31Y8vuTWE4lIVaCI4O3xhxUj6W
bt9TzF4D2gnr/gVGVew+FdcPQWYf15JCndJBVpAxj8NrokQh4YbRdIwVuhw6tB5S
Zzq0vV1T9Iht0+i2Niw6SiG7nrMt9kE3MmU5aIZuMGJLo2L+8df/H/vqefz5pfkX
fWGaDs/BsGj8xTeM2DRUxCrLz+2Sxj1Rrdl+VtV1dRFwmo6vIZ22QIMgVHD6bzz6
7LC5yQMgvVi355drRhQLwjUcG8wAyjunr5BTpwhDKU0epQ/7SjeN8gELx5yrikjY
BfDHlOIOE4xhheIar2rETPYpYK5b5knlQaLuZ8ZlZNw9uP/H3mzoO/0+Pp51GgeD
7CQAdYQSH4A2L+tAP3tQyMkBEICmdY6xM3KfPwrXr9MTLs52vNBfHIs19g4kGSMf
n++BSpGfrO7oIzWP3jnpEDhqGTh8Y/7mXoKNOoS2/pbID2Q9/WEYa2YWq9RrY1fN
opWSPyEe4JFObUij/jRnSbKKIH0O9rxwCTTJft3PLijFqz/wwTf+Fbb36BYcGJ7H
ldZ83fP7I5c0ZL1sOkQbAINW6+w3k6KFXV7EzCpG9d6pY2dxJFSgTx0qzsEep+67
TjItaHF5VSOj+dPPNVefkg9T6Rsmme+1R0WAftSbhpbr0iNcPfJ0G5zBQO8UrHQ6
8IrZZE9zlEzYpb5YlvY3ycXrH8y3X44FEVRdyTD9ZAU7JV8he8uUWis7dz9QWon+
FAK/4WSsJmHIVZ67nkmwDvQ0K7esXQl/SyMkWKJku/t0frxAWnbapL1fDexKRcoE
8d2bbNeXL2NvY/81gEvSBwf/NYFOZru7SXTxGMZjpc9j6L/Dib5VUVmcy0sIeWpm
7rRelaVAdO1hKXuEC+FoMOVA23LkDiG3LENf5Q6oBu4FQQXj1Xm7udEI2dv2MPbX
erK1fUYzrJ8a8AnUBWCWAEOO9xyiFzhg0guiEvHNT/ZMzxcjUTIp9m+TBXy/7LPx
ErJWKXB1vutV98psZOQ41AhkgEjAHBorbbt/e/UMTxGU782aApkl0MM4OoAGSxyv
jKseilF/jYwIrxROi++GfNnyqYbiYpYn2gUtyiTsvN7lyoWO7wAwWk1NBIGXlErG
Mi5qwytS7YUrMMSlQyclbo5bDlo10iRXYJgyUzDR18uTccgbGliOMsFIGFtElZT1
TvMfB+bx8BdXCzpWFlB26ufzPIzYHulJe1twrTSuWcE3Px0LhFjH39H4ptQt4Pas
5L/H5VU3gRTJqihiTRvZDWc9TXOHWRu/mLbsSJA8gurl+Yt2ZP+wxvWh9A6/eHjj
cmebIBwTCZ1nafSLzTUheViUcq1Sw7ZFkEqRtsKjtLjaH1wWU3A6BgNWDM21h2iH
x71XqTNO/ZTPg8vUFwqnLTiULG9NXo/jkq0vxk2SDTHb8p6vycXNE39JKdnqASIL
Xe+NcAiIxFEjfF/9g26gECRoMyO+ujlJUZpJqDTr8pb19gCWTFahkxV/tgbzyX+B
qhRSmSBPAw8owJa3AGMYnW3dHyFPzOJPPd8XtHEESnCrCk+AsQxH9u+3gFT66Kra
f31HJVVAnjym8gFuIjik5eaGDsQU2RUxuLB9H4IT+akmtGcm6F0oPilR0MRaR5sa
LFKefJUf2OIAp9e3knrlSeKAQUqt7ldrCR9JlAZMcREmkuxLdq4LueEEVo9/xXFM
7WY5eUP66sDuJ7jN4d/EDeohat5szfnmdsSQgnpzGdCZIbJC8ofiLt4dSSEw0/N9
OJXn2+X0HBNT2RZnROokppZlvouecsbI3dCJL6fSf9kBUdqf3TmouISldaKC18yk
6ko1kP5grmzz9CjdDrGc/zafJEqEONTVqVpbW3R5kg8hTgpy/vLrVZ/3Xx3fPrws
TIGRSfeKU/wdYpzSwmsGk1+8M/yi21spAm0ySaHGH5LZ+bHs6YrtUoD25OWpWxk2
YKd5oHgFSDlECCERXt+fAeBvpTFi9Q67ARt+VminujIZ6pgAOwJiPU4r22Q2XIzN
IqTEP7xPM3nU+3AaGQVmP7VA+JpTVwmMFBhsB4u8KrcpjYbwzNjnOKqpWcrrhRCA
BuUt1J3wW2qhbyKiqwYk6FB+PXGdhWmO+DnwPDr0+drGiIuQKMb9xXL9sAFOWcew
e8gIAPFlan2NtFf2HS3YSgLps4oudcZZ73zMOSZpLZX9cRN1ZtDPnjJzLbSl8Tn8
PfCaBah5BDFiBrwpM2Z8IO7wTVI58BgGKXAOK23jqzU0dHO+Fs/enx+zkXLlA+0A
Em15N8UkeeHCspNTk8UwIM0erRp0jwPh8mwfl1obKSyZguFvm3V1EcP2Flgv1o82
bF7D5fhLnIP1hJ+5+TidbL5HivMz5CJTS5Xztq0r8wg/RSvDQDQKp1sPvxhptnc/
dl3CWLblH72tsJLKIsgba+xR1xu2UbsLClyBK3uS25lonDioLdGMCRyIhc04+zlc
MoAAvPe6WuETtEFkOtsKKeJ0z6RpwVgTizSsJi0mFKedyJv3uWHcsXuEBzt4zd6W
gUOKXRhd9LP8BiYWskHS3WNoFfgS3g1y4Y93j0yEapWQUd60SEEQ05mqXQKX0GXC
yc2/uauadn2GvS/1EBbuDTkVJt0wZ0txQpSqWzVxJea8mAsSe5IN52xcbyH2dvsf
d/4Qt85w0PpLHdawN2LnFRySa4UqbpomOMbhQ2NB4K2oG0m7wl/e0RXOJ5GPgPG+
A8HOckKPP4ctUJRLDuH9brcMgZovY/3Ap9ULiNiZ/fZ2ZoGgqpaVB1bRNQWORISF
bmG6Rl6q5o6GMEC8TvMLiznpLjSoB86sNuIyYogWBN7CFx8yhSty5Ril0b/M37uD
qR74+8VhkYA/kLNtWruTGiNj+USN4ApuaGxud/UU4U5fwUGDvWyZLsK275CIWVV4
lMJ7e4VA+gorzcrt1yELG6Y5RTSdbabAmusHnrxWILUdQeFJ/ZvYBJJuy3Pfjj0o
s9CNp6LvOmQWAUM5l6MB+rCgaoyf4s3YmDa9qCfFB9SSfybn55so3Bou7UG0NYRB
AyY7hdUuH4gg6gZSJ8M4Wc4oEmQzNmaJP3fmdCY4u0sRX1n7ew6d2jPtr+wnJIUb
0c0wCJJtwvkoJFYqjjMc9TptYsurtcUPhJZjOvErQAFvI0mb5TQ0gIlTdKkkXmMD
ov18wEVqaGKqvgMs7w7jLtFgFwROIOPuKRFQlN6GlrDMIbKUhGyI3B25CmOFe4M7
Yrd3GS0FulqDCreTwOegt6nQnVo2I7HvPLT557fPrOdrU7/5OOwzI1BtXoOWf8Dg
3McjuEmoXLdlpeBPrn14fqUQ0c0po0Qx+Iy5tHT1m5JWBGuM18BETAArDoEoYMG1
hJC4xHdaZfS4Vb+sRtksUHOvxD4Rpf0l/1xqroW4gP6HsgoMiZ5fdyGrix/JkX5X
ZHF+zD53JmesjJ+F1er2ktgqK0NEa2D9QuvXi4NFCB0FlylbKWkUHa1cYz35PDr4
f0bAoW8DQp94Z+jQG2gFsnldtAzPa5KrEQlhkWZ0wrLzFYc7X5ZeCbrLGb9LeIyN
yyfmJrzfOhJK3yf+66sWuZNNmtdQJmON7s/T/NR4JTlMwbPHwiPq9/tAl/Ch/j6Z
S+Navi5GBljbSJTvTM0BNxiqzXqz39Chw7kc7SD30o6qL4IE/VaN/m9PgxUrOcG5
kfHMaAkBb5ewHq6FG+M6iXc3gB1Fb19niEDh8Ybby9XJzig/BFxNhnrJL1wT/FsD
u2e1qBFu3phPET4IdGVzDCfDG9rp8Mdc3R+WXbFZSI919i46Yuhh1LBl5/7PRvQ5
s1ZO1j6z3umZfHNUrM02kZSOx3zJR5hXAAoar6gIENDeFmeaOeIpmpza5fZVYd6v
4mSUqtzr+VYQOYNOB/98hbNon31vvErvdMZZbMnJhpQSVn1sGiH1NYXWtgXcr314
p6R9BmpLhnNM0WbSM4SmZSRiAUJ4vRX1lyh8VHBk7RwhD5is0GyEIyUvTyaRDoxw
0c0vwEE0Ozt52U7C8l/XPBADVR9QFZ7d3SiulARgrT6Y5an/EE6Er4mSRlkYHuCm
j2b/AJEBhrOAXkOWummeKppTJFzaG4S6UYkpPmPxUiqWgo6LzWxpGd8+PJyksISV
fDGyRj4whLzTXdeCeV5tt/K0FqXe7FHWtquYsgc67ec89cP7CaHjsUL33+aIukW1
Y6G8CHqWUOXJirH4Zh3PbQ0LHx2aVTK8SuiZJTk1lV/B2bESg6Py+TBYu1b6/DeS
tHF0K6EfJC9kgjOQAtRUbOaBzrEbL4XAdkqBIoUrqKwb5S5y0nC00goUdwSTGops
flyqGrHtSPC0yHnx/llE/MRmgu6IPgLOiUA1qn2xaOocMJql82A7RBo+RnmeUq5C
0UqyrcNm5LfDJNMcV/lZZh1KY0ncMMqTbNKSf9mAYrs4aUTUw6F9KjBHXkU2Mn1J
feiI2xSQnhR6G1BhVWBq5w5dIQmPbYXFqlVdQhaJqo4KmQwIBWWVTHaE4ChVCm2J
IKZTGuy5Lo/vtyYvyJs8Op75Zg/P8k3P82Ts1/loHR+AzN32EarrCAYqJXceXbnV
fgoqZij8ZDo8F3PRrEylNsZgFiaAi1yj73HuKSIqVqh5/n3MzCuMdQk8AVKtQROm
BKpxn3ngP8Fj6Dcj2DOw/Fs6tAUetgaMIKLsz2BDLVGXO4vVARJ2aDuaDnRnlnLO
Fnss0dHymr9QA7D1T5YOCVf4ZulO1yIHCh/mMFyvJL7yQ6rNW7B4iZ26SOTEAKXE
mRg7biHZb5F//1/YhGyeSWpjzfylfQW6mNaPWZXjEP6zccuSaezb+lvgiMkG4Z6s
NFHWs4/lOGSQmwhioctkdyj3nt1RsZKNSlxGHqB2q9YTghG3OWswAnpO/lR8eu3U
ycijJQKJDM/XDDoL6TIOBvFjfJPPZG5tjWwRcLv/ILnOPdXOdzIw+sKdWf8F1sb4
I/L0hCDQybKeFj+TLkG6/DRiYHKgemESEKHaMFBoOZKXtm7P58EMMtQHYiWkSqlh
Yq6FPvIeqliu8GWB+qlk2RjSYeQAgs2HSrPF9HF+1f+azOZ591HzP6l4z3FVGVoN
2tAjyKqf1/9u82LBzAIQe7Zm5hXFmKyvGUGyKYLCbCa4zx+67Arjt5tCkmjIRvLy
EtJIhhi1WdLHglSfc/eFa3+/Pb7AXN3utMg5LqbfpdSK1Y1zfVVIXvrZ5SaqMrgi
n1Le5WoZJyaMaLWZDl0AgThcI/d2RUumDx1ygBaEY2V/gIzf3V5YzK/xg/C4nTmT
MR9ozXc4lvsNVrJ4haMccV/Q+XmPMzLtrNZAA8juTC5QyNxzsZyUp8LE+M2jwNpJ
O275l7CqxJKVKUCyCWBhdAgrcRBdz9deuIP+8bW8yqyLMTEvvgXs1nrF7BDQ+3fx
mCs4G9XGUzyW8BRE3lkd8cjSyh9uBcM0xgZbtV5LGE2kwN09HSNUMWgEsEMdCAf5
1pPVvDUVXdYqEH1P48zKLgeBwJpmInJS7q+0DtSoin8a4wWvndrlFCo4XsWYv7Ta
qW9sRdQbmsSXcMsjcABJvgpnrRbQUopGolSdfKme+qA/jfVc3O9ZHRjyFY6fK+5v
zF4+zEdryz7fJVOF1flBmD2Qnd494aRjx7xYB/WWRptwXaCejeozXYk5FrTymTaM
lGMt1YGdmd5vjqEjqmeddnrIfz+IzMPnoP74Q70vcw/HvgZLm3rP+N7kbdpomy8L
0/xd23ZC40IwCybQVICBeJjGlml6CbN+Y+p6h9/vet2hplnHwqFR8dB8ZNgc7uIG
4akpv0/bGbBCLkDLxgY8yfvy+9NKnqjR7gmHOjDhZWY64Mxw6M4ID4g2oxyFv19m
mdyIlp1547SdCNLSo6wHVjK3qU85gypgO/SjJZvX4f6TOUyVc4yA9tT6PG9e0NVY
aEZRPsXTab5XGyUFz/0zjQyd1Hofbp13J14f9ou+g1Bs3Uo9mzT4EeugUkq/gTGs
FgjcOGypxN63X8jlIGhLWUxkjfITv5zP5Uj+FY7iCSJSxJ6q8z0W1oVjGbMaTh5l
4UCRvJu1ddJWUU+tfgC2Z6rGm907+a6FPh+nwUnbnwUIRfcXAGQCqybxLV5b+FG5
82dTcfS9Y72iXdxM7sTNge0UFPN0ojnBTrO6zgiOxA3k3jNrkTyyZdWBGp+I7hIh
2Z/pOxR02oifVRALKLKzZdyZ4LbawNWTOWtjZavCMLMTanWk7PtZP9gv+6hkmSBu
cE1BqKJGxdBGLEivkWMKOyQsdMgekHknfeOlHSSAg7FvwnCHGpbRI21EqpCiB2Aj
coIGuDShjk+kghSvA/+s0ipT5uTYJ6b2pxjMOOBHitpsk3UHpkG/VAvyJZQrdfAW
iRRRlrenFzeny2LzInW6cdbonG37r663Cr+C57a620AUECAqC5mVM1QCkBGEvnbL
GdxLVUt9VJbg1W/nldEEE9gcjnT+0w+m3ROnWcNe/gUtWcZnJ87X6+cF/iwjJUWQ
HrKrkVExwRI06crurjlO1Mqa44jqWm65HMfQDrwe/URAhiJ5PxqtInuyF5Ac8SZN
bbgvwEWhpr7tbunT0kxezFTmGmLTP+Z9nlu97Nlj/wA46b+vo2c6RCklLCfGYb2R
i5p2CaQVLWmB8JU90gll6ppNFQDmz2uR5bmSjSyIAUV0t4ktlpRkqNJgEK5MX4oq
TXrXVmu2PCkA9d9++BAHvgpVicIxPsOk74C+gFFoLloSADFnMdR95cGrnYSDUOeF
LblZ2tCzmR61uXm+pM1XkTrHNSIc4xpy8Pi39HtowhrLjBFVgkHbXN02uAWz3J8f
3SytKAaUl7dq3WjyBx1Dyz/kLRpdI9uCLzY7joGiT4ThzVbklp39A1SZyMaRywI+
uDaCw0R226TNyKmw59Ocu+cvbMNYyePomm+nVx7EsPJ6GvdwVW56otlJ0KPtZ+kS
tGhNUYsgC+pOlkAf2c9qjw8wi3QyE3hSpWtNB0g73DpCh6TSFYlDD/4vLp3DNVeg
gydPYfLAMWAUWJsEknOvADullzPTyir3bqwoLMK3xVPC1/+D+E8WeKms24Zl0yLM
on1G9G5qaic3ItFy3hMCJ8aqQAqNoJ5QmtQ015OsF9ClyCFBNKOqqRp745U6AYl7
T1W8KwBxY3cyDBjRdR20/2vB2P6sG43n9vURtnBZlEI9Jx752Sdeu2aMePJV7iQN
I/A2Pl9Cm23xjiSIO6V7cDVRW3K4vIse8jCesztfVSmjV/MxAilrVwf/ahmN34se
t+w1PiBMSNuNj9PqgkjwWYAyOwfSTQUOF6GiO+rf9f8w+ev0V1CkMcDSus56T5mA
4/eNA6YPLe3u+rwKAJ7dyKy2htzAsOkFlfEvqu1ovthNQ83W4XDkZUXzuenpBkMJ
1ihFASmtOPYcETDhclOJb/yu6jIEpj4hXdD1cjiSu4lH5V6w+I0GQY9qqGPTbT2F
aAOUg+KvKCX4DBBXeuZbbH/aNW7v7/NEAPL1iGViB22eMUvq4lLiaBG9bdBTRTVD
qWTlnvgmIV54SJJU3e7cwKR8Jpwk1A27m5p2Sal8/JfmLaMFyf+PKTsXh5qrRLd1
I1f1kfcCaB5FYLKIigCqO+BZNIHlHTGjbqfMtmL5S2xOtWTlm5s0g4xoPEAz8DhZ
sk2S27uZGZAOHSHkWThLvlh6OHKJXBsNkwQ5qnbmyOX2oQglLHHxdGAtOPDXUCmn
RcnzwryhK6Q5ScdRaX8AFM6sixUAJiqHy8cPJK03rCMezGsWHuS4i02XGqtFNWci
FsMafK+W8klKymA8KcDSFQ1KAWdnlSjsBsXOrc/EfYg3EANgz+46B4uoiJmVz6fM
NcHMLN0hNmQVryEu3c1eSFxUMs1WaYD0P/5snIG1YRzcdGA+UaFP2ai7bV2Xkh84
hebOUMK/Ep+A9AbzzFCA1Y2cuM2lZT2KRr+EcU5xCo6t6dw/3SsQktDVR2G0w+jN
/gQOa+zU8GfNOqFD2d84Ev5B2HnMPGvYrdr8rjRifqhmhJBVvztPIQd2Ex1l1Zbg
ZIPucIeXcZOTl0etMBLkQ2NdffiqB2S92iQ6PptlS4AGj5C7e8j+8dON/lsUk3+Q
JW9QZoiu35IAi6F04KupNY3PQzU1QVaAliqqmVNrwbp8wvdIoehV83Xj//tTZ5H9
n7v7bySU7MJOS8033P/hnlXrMYwOm06wh8XvipELfzg1STRM4k2BM8Va//nyt6Hn
CiaixaiuIbAL/DV4hjXHXuHFSEER+g0jHkG51aV5EWIgYVyZjUYYfxK0q0S4tC5m
vmnbE4lphLP16VyptaVJKChtuk3+iF3g49mKy3sADrwXhImd/QSEdcW7JOcJ0x2n
crjEKnIfO4MFIlBYmsV9d4qF9CAYAngpWQnXCuwvOuksVYj5V5yAKTm8Zchw1K2e
b18n/fnaCYB/xsIFqW1kce0/NQXjJJfAz2DZh0kxSRfe9jGgGdpxAjw3RVMkvo0b
cuOGzCLLv0vAxADHKr67+ctfiHuP47WiVIkCH8ukNpoRE2n3wGClDfAzLcLT+2fX
Ak1lU/zegdWlBQcUwKoLxzG0zg3TuPDxLiSsTcNa3EYuWw4MUV+to87TxI1F+S74
Vto9++K29E5O91KM0cFnpXogC0eOMug5l4KHnRnIC62Jzw5vbYOabLIt15y+Rkhy
6MSSa3VE4DIelFa+ex55qYNylOIXZo/VJfeKuklxZYGVineUt5tRteALDrS24ssE
u7IE3JtBR3ew6tFL0TRYA7PtB5fxSFvBrqMvnZHtrTLcxD5MBf6c31u0ZfSYPCe+
UFWnq/ZyFArZLrg5yPPuMKsaqKg+oyOMnzWR1p/7qBIdnickL/0HV0HHHYDzp++e
NPbKOOZOGUeJWh53Le9x0zDk/0qSLfA90pF7AIhmzl2WSSvVLPz2Il5AUOfsmWXY
DnDom2j3Nj39ftN9Q1rQ4i4tP1rNJUPbWeiZFhY13Ikiw7DbONg0++yvnsi8tdGy
5PoY2/pNHKEoHYCgZsJfUkAv1iXidjrLryBtPjuDLRfXFa4H2neC7ObuQvMMnVS3
LUgg5GFbvOrTm8ceO0IDxGcO/+6mu+VXwnwJjSbr55r4XDMDeWMBV5m2GhwFtWYS
cmNHLQ4n6Cf04g0AjguruGddb2kbk+JGbem+ah/NTO0F2npqvhyG4+QOYpFaCI7T
Ypz8EuweM0HlNEkoChrgz9RTVsHoDuiTmlBbwLcLcytox8F8RuuGi/m2nkiqfc4h
tXZmaIrcZfeqKxqX1V+0hZKm0PXOgV4cCFf5hWVpUjn+6tfP29D+0vvn6MgbsG/W
pXGd3F+X6fyKX2MjVlWFZv6Vb6nGb/2XhwFxSWn79XWwlwrC49v+LpGQ/RB5QaM3
ELlzbl5hkVRUvS2osQYda9LD7eA0OOA3MIcu0woybha/FXJaa2JtnL3iMecvT196
pqmAg3iueFTefznWgP1Ge+O81NbNdGqx6Al5E4f2Zo8Qg1TGkmfVZkY5EeBdZzCT
XQ9NbdLiZzL5QMiGn+VL9PO8/lGT1MK+XqE+QrwNOPgg0i5Fuh08ISC8d6/d1fpO
IP9Njenlgc4iRgYLcz2Vff5umT7jLiz4N9To/mTXg37nIpP99eRjym1oBbneeBLQ
ihZlNOXMyJMvM+9gWCRiWhCoDF/9nEwi1h2+VLp7Pi7TmJQ+b/M6aNxKiHJ4ivFG
IG5WzEN1+W4o1zUvUq4Z4ZrQhUjcw5F4lFmdzKU4Zzk1NBIetLevxMERdh/088Kr
44LyF+OqvKrd3x0ddYuIovNwbDT5GvEqL8bN2KRrRNeeGpmcMdLTfTkxsZD11N93
GJdk9QNaOPimEeIfsDOnpiFYQKnRzOM81ECWe7h0icXvaElopEqXxvrPSmTB7SxQ
XG55TYE6HzG76KFhK1imz1uUFDLN1cIda3C/1mcnz7XijIbjXXbtG+c6Lv15i7BE
PZAeM86GMGdkO+DlM/NzcIbCbEwZm9PTM1mavkFBlbphdS5N8Mrd5zufNhuKAQjd
CrqZWcj3TPq83HSywafGdDlqdfBF+8otG7sX+u18IlulRIff+qMJHBC2PFASJErV
Y4Fd1CmPKj5H98KAi9+mumqbplEv+FBqgyinm38WMRNlLxXAlr4OUOeRRCmcxrKp
W63TLpPEpXZVrgTqFHXp8h0/2chMpfiF/XHWTkFJXZgARkA8gsqLbkG8EM93XvKx
OpEM4qdYbYZJYuG3FUQo0Ag4xt4Kz1AsMREof1x8nepuQDdap2yBAjrGYL5g3mC2
Rt3BeIK32BkWlze0qHvAOasuwSHZGhQaDz1z0/2ToXtcsjC/pcUvIwN0D+6VVDx1
/ezNup82nlTR0DbKO7fSyhHeQcjOmW0FRpge9oATrfrGtQr4gDxunhMtNbuZtWSB
FzTJEMWGlEJGpWYDznsijHyN9arH286AI4kge94kvrqkgWJApZE6LtMLM9kmDb/h
Srt34yc8NYTYEJIGXCd7Eqh3OFjp6sQgQ/7fR65wPCBxzx63L5czS5gOA1Q8e/jp
edtiQk+PofaRzaO4DYbWCSUeCBiX9Q9hJwu7SV7f3Txj3OzcNBm8O9LYIaPRWwy9
pFNKQsbbGFA1xi0vUmXhdHL+cnPtfkoGFilCRrLvxdDxatzkR6BtIXAJREI9elXF
yj/ZSf5nmEAolNde5vbrOAmKi7SQ6lknVkcUGx9Jq8T5syLByTMsrFUBJ/nybvem
Ee1VPKmi7MNcaHsQQCU9i5ywBiklLdNoWYYKy+5w595V+FoGZYFaCJ3kPoUApAel
7CGU3wO7AeB/Nwo+q69ikXNtzhUgw31EoO2YHjq6dHPwyNf+CS1mumfLIXQS8vJY
RDpKKAp24RjYjAS/Q6KQJR/iLtDJ+wadd7SC5Ua6LE7oCRWHtCo3CiFYmMxbeFsv
kqtYwxB5tgoxgisZtCLqY+cNMWA2wXoOXbyS65eu2fYaWaKeSMXnDxSLT8gCXF8o
9vZulpYW56WwYF+32b+Xt0Vh83TwfrhVDkAuLil2mzd9/plPPjq7GTeAJQ7cSonn
oyLzw8MQZfEqAZ97gDDGDOf9c1fXjopkTCIqQSEn2SL7xJRryX757o5X3LY7BTXK
GU3PtlYyuRu4mwNwlqHVsWzqu8Nxd2rAMiDRuQSuviFn4q5WxKMz7eyBYInsUBwJ
lHrJw1t1Ye6TsIqFAeBnErCEDnp5bXFwWBsq+SaVuk4E6In6/pRLdmXjOtoGwhFk
aimQM2+qqehb4+XMO66QOO2s0pjXyfR6kWfDu/xCCp0s03nfI5Oo+lPpTeXucnkM
NcVHhSB4wS3Vhy6o2LhW1GeEu471JqeDLc2Zx+KBwa6uO8mqQsRV4uu4KZbBIaSK
UNkRiPnMgn0ybJ/0tYnCZtGyJ30JDeHvxrDXm7PBI1axkRWvif1QKBVBeTxBNog0
QMpb0L4J2+OAsxN6ejbp5CY/Q4wgm0V4fTvL5w0AOqhs3gGnxBN+ys+gCjp8Uetv
dCU3Nr4gGs+dLMpGBsN2otrQs9TeuTAHoynJVBl+0rAuAQDfULKF9mNCVZQvSv2l
X3ue6UWNEp97qL3sE7vRUc/cUB595lPFkdcS+gpO2p6n0ZRYCEqMIsePLyxC6Qee
fSIoNMleIRPggz+kC6cTsmfAuolkwG91cUQ2UcRdO/th8lNPpIltTRjkNE6Pnp+d
w6evk7JydGWA4PfQjSLljH//wTClbGBxHiyd/2jEjwbpO3RRSgo64OkPXFF47Vi4
ZV0bWVbh+efkxE0eE5d0D9qWtlflXsR/wNFYapw6jpuRBrWknk6hPJKB5HCJbQCm
XfJ/Zdmi6K6vllh2LdOUUETXmwj6Mz2cvy4KrU8P991DqSpXUBqhE3Mo6aHwkgcX
iz8pIsvaGZEnG2mcuiODe7D/1E+wrejYyXHjKdzdOhQ4F5ffv6uxszgf/RvmfIKy
oZ9wI5eLIMX3cK73JPEeZYwJ+aWY29+xOxV7ePBaIyQ3RACjhS7/zCjFZ/2qyFNZ
OuGNv+oPQVtXMbjDQ79R/T8neXPqgIZLx8QWmfZMzPWE+gqhlxjHoBRyU0UvNmFo
Bxxus/V9lLBVAoscmmKdj/M3eKX4SHZxup2nst0Wv5me7AhMJR/dQ2mcxBnCB5Jd
Zc59NODjhiRDbtBPTfffdColR7V3pu0GwiC4XnAxOLx0yozZWMXXe/V8oUhSWD8q
vx9ouNRAt/JwRpNMb1cy1kgJAEnJB36F8xriCfmcZPGsxOrh7I7oW6HzgypbNj/8
4LhZkMSXnaN0LHvStQoB5LAb4nwpQXKNKZAgXTFISr7cHQPmNjsr0PIE9AbwFgkZ
Iy5Ejz2hsBCouqkRGEpx4vL18LzsM5Mpq1OHCrpB/EO9aItTG/6TYHYvvy8mUBqy
FprKr/zSj85Zq/QZRvB9Pw3Pu/DP1veCJ6w0WTiUbTm0gjso7ILQZG7bAFOYZB39
8M/FPFto3Lwv5tSvEw/KGkTqFkad8KlXkTmMH2oHf4ux8sZkzd7pFa79WJpYpnoF
4uZRPNoj7camt+esmA1AmrNRF2N+0t6GJjRVUWD16uYZzLqddIht0N9Kl5u/Cc/R
UFqNaYGoEvKGz/hHOkYAZ1636QP1IP4mtvXIkmYN+yiZCoi+pl6WbfyjeqoDTN+F
enhRtaZT687396cOjnhy7nHXC2FKNysN3B7/qxfjhnITbWFvFGVW3CG/vdoi8/vk
lMUw8qchfS5fDyOdACl5ncUfVzzfcCiFgh5AZ2lVoZnHqhmJYMXfVOitcjeGUC51
Ec3Cq2O00uiGC9aOlZ1WO/fF/HqYAIdeW8Yr8o94iDlnQBjGY5WteQnL0Dd73pzH
EThg95VVAw0NkkpvN4xPwLuqGjhrrfB2maPy6aYMQNLYkfZhrsoe0aZdnPdKTr5T
GiMSTu0rZHstdme/4xsuJC9KPZYc8dw0+8MFndcU6p9bJWV0WRmM3WXD6TIcrC/m
jzGqz/kHzCOHDW+jWotrVzaNcPK3iliNiRZk20KT4i1FCqoSN1IDcWF8LBJCFc+M
xM6lScJ0lMJX4xRWrGiVNhWBBqLGFVx31S4zwXESbmFl0pcu8fiCc3DbQZF6XABf
emk+3HwpsadLD2sgSEykk5Q12jepmt7ofvu/L0e7OBq18u7QeADMZRLZggGV9dk6
y7+IdCWCHz8KWXbP4Oghf1tCKCxGEfRvXmDR/iZFakfxdbiukFWDYcMlH7EZwJb2
CuhldpkPypfJgYA9n/1W0HBlLoX3OLvePA41gGhZqLWEwNmSNNcIyvycghzRLOkO
7lHi6SMxfeI0X3XmzD52T4nGAm448bI0c++5LiN+cT1VcZ1vTqAv+b6RFYeEtIO+
lpjP2CvFztfncyrd4ELeSjoZ6tsulsSoFtfwYum7mxzFYnWZW8bqUGGqhKAtZtwv
tuq9O1WTU12TwDWWgtTNbmp0Da50/pIclryL6iHFXs0CFRLX3D5s1lZ71fwD05Sl
XorkasmYHOmgRuLjFJpDxkf2sSoc/MdzSI3HvzVch4+E3y1Dh9M9IOh5XXztJgCh
FBCmffZdzTtpj7fVCl4ruuQG2gxKxep7K3xrvKMARb4UfVX1dyX3aYucHRvss4d8
uzphn9xMDc4yrTn5C9WzhnSCOujETsMPbu53M74NypChCQ027aA7txpYgjWBSods
ftIsiw0fgZQvv06zuNT4bzjUOMWKk5Q4iof5y+fu/zFbHA+lMAC8KyAlVPAlhIQ3
VI2xA5BUOCKyzx2eeyg1SAQPjrqWELT3kaCwJUa0A+HAWYZkgndfnf5B/eiQpf7C
XE2yT9BMaNGKSo1x3Sds8wnpSlDMuIJqAWVWIjJwBZiEmbp/OgAT6s/dZ+8J2bud
8LAEwTask+3LdLGO4DzviLUH0t3RO616TWtc/ScCzGSjKPhQ4aic+EPjUE1GDMlR
90KjzFDUZpKktppr/FO6C6/fRmlZczWT/mmnR13eFxyHthKmHhl53Ys3HlS/l579
FoJ87EJR7TqBbsJriH67uWEEicuS5vjtzueDxWjSdq1V727HmwCdAkSkaH3kiHMc
TKI/HqTd8sgb0SYdA0q9InA+5Fkx6zukwiwt5iWZ+4BRpQwLQl5y8JmsQ9rOuflr
iWwY5njz+MRvAG1bHxialB0CVf9LuR5Bf9UcbdUdI4VPTLt2MlTUHXnkR8mQuJYq
NYiO420CxiLpQ+1LlSEFfmQ1WsdOsS+39UtMz3YvgsWwk3ticYZoN4bOFTm7k2/f
1phlSwHHdMxI/o+votr6YPKaRnUq1JSLqFP1G6kR75y0/RNYwhU5NU4wTUT1SAsm
skFnodxF58UhawbAhEf9CugPwlc6OxF3N0x8vRxUPJuLv1Swyem2df5d8pima/n8
vZtF/K4hg8FSdTbo90c8Xy3aulVQO+29ejMbkltQ3pzFgCE+zK34zBqB9t/avHxr
i5Uk/MEXhFywbie8vwGQSZIrnwqd/S+/YnoiRAVwXw/zugQOeuxtL+HUFAb2Uxy7
kh+RhrjOdRKvg4yMQf65HSvP+81vPQXh0l+gcA5i0/02aNL1/Xi3F30/DV72A29f
uaONvPjLF+OxQISo+akgiB/fr8+SxbEqeG4l+jR+837QBxHEMHx2tHfD3SsTI+As
YLM3nhIrU+mr3SQcroSKpAVXI70Qf5giD/6IP3jp4IyNrMkhxTpOG/VFvj3OWHZm
wwD3Stpuc+3yrww76jtKZJjuBjKf41fJiJUD9b5Wb54b/c7ziDXSJy/cQ6RBNxvW
9PF7pEpfhvVL8MEdh6JTko54L+Gjnk/HQV8otBFhjp1BjMlJ4pa6u67Ll+quWux2
3LhPgcBl00u7obI7Ia0Hs+7yTu+2wD7eHXp57/5RqykJGpnqUBNaAvNQCp0pmv0A
on3yZ0tdWsfOgqugdUOWwPrXJAMpl53QyrjqqVElngo/eSF8NBk22fCpOu1T0yXP
YPvx3/X8N8SFHwG9l8s5RpwfAhRn29ZwseVY6vGm71nhnVxhB0Thk0AyFzvx0Lw2
oJLPjq8BFX6wYna+z/v0J9VByBmqErzqPaTaLa5QnK1rzw5+3LPVSVVa4ONwnkD5
YHU59y/vcAaVii0AoFSbLAwNYhVLIzcDzZQKGTqd/Rsc4mAoUMtswjmsTdAer7HZ
ppNLoC7PQ6fYhrNq1WdZzfSrW9Uy7iYpfNSKov/FtAJNPdpx4sosgP9PWIEgd+Rk
TlVA8S8TzYAvt3MwIo7TlwO9s2SYr+BMAG05/dBWOwjwtz287duwCuKEuYpkg5Sd
5wr//94MtfYhSROhH+UJY8qGgiXHrwpsinAoSjOvX2nOjZpfS8i0uvKWxcrtzqWa
QP+N6WQqf/Rc1J0zDWbaZNULZpU1BMoEDRVPnl3eYBM7swOXHPTY5yw/wurHTkPI
5lVT18IQNy0uFrTu0+vjo8AxH/YvCOfpIA68CGE1EG1oPkj/Adjl3STr8EHETNcK
loGWl6zs19e1JmWbXoQ1Hb24eLDYXfFIVLJ83c2iwyLO0WW1tYB9+YhpTTx0/m94
YIX5MGVbwjyTNEwBvumlPXXqava4BL9z3Ms63VmKDUdBrOiPdvGwINtok7Z77cVm
DwjyjNE4SoRGbD9dAre9aYvw0bVjR4H2L9u5QV/tZUS0BX2tJDKFhptkvKL4AQFD
2XSMpm1SUzneRn7dH9KdVAJR3o21OGX0BixRjweztYDlnyW0Q0sS5/P0J13Wbnq7
dzf9s4e6obxktDL579a6HbjyMnusIeCfkLyIHOpaRPC66Qfc/5y0Tl9LNBLpGhBs
hp9kE8uoMlOXKEKzIww5NSPNDEUmJG4F3lY9yhcajBF5vt1GFroGYDZ71T28dK2N
OS+kd0JZlwI95xl1/991nL75Ea6RIjGKp2E/e1Km42sRnzwAJLUoHZksoX0bpJKv
CQC3rxdFco5TGeh1n12vNInQwAyM4FNcFDCG2Lx3dovPPUfE1z9Z7E+3cHQixVk9
KVQNxAHJepspRTW4Maul42s7ca1e//6I0OErEWFxyXGSybERzScLDWONlFG3//Q3
LGsMiT9VN0nucTzdHTVqCjBx7e8hPHUqVo/30J4kq/9t/ptqym3MeOGsB0mU4ZgJ
utuILK69h+xd3E8h3A/QEZaNe/IMTIYsvOHxo9rGFxmCrU3S62CdWdeaYtPs4iJF
mga5lM9AG3H9sAuNgQ7R2J0QdeA3/+rhpTXY9razrLbQkytqHQ+w2dezjq+F9E1G
sAGOAnlDNUdJQ1ExNK37vpvxKhSBzS58mwYZIJ00ZXgVNIekN2nuaQ+PGOTlLUAf
PGv8DideqAM74UWx13BJBPPdkdkf9i90ulruhmARfuwUxf/Ak/4pX6uTYGmj/gsn
Q8QT8h1KmJcWTscrh9zGFgTQ1mBlbIwkYFOpgOD524r1ltohgv8MNQ6qLGULyoLQ
Q5r4VMdaC9FRZAU3wN3S56MuPBfvJScIM/VQvvflxAN8GYRVKDeWhZZuySJcGnW5
J885mRr4/7/v3jGGFzaiIO07hNRnqPv90MSNM/fxzJJ2LI5my6dkmHFSqEj4tQqp
iZAVt6oR/c5yLr+i0xaxzimKU2FlUKWsopbAyP1T+7HTmDKsMKu2P1Zw/2F5gPMy
LcV/A2g0nsp24F3iZA1JflAMKIWDm61qbI6P3d1n9XOF1z5uWgFuibpvR/T+HBOZ
XGB0L9Epc/+8LJfS55vUdeQUWtAgzbsuS0MYakB2V2rjyuiBh+Dp+aylwRboYXv1
JzlC6ZJ3LCGn/o1mkBtXba7PP6dxWgA2ln14hxwwmsjdr5qSUXpRxrSm1RsVSvLd
lSNc+kVn381rSic/Mrz5vXNIdnLHPb1odnbEE8+Q0BSkB0fA9y7/e6ns49zILRnl
oVLwIovbdjrV1IYt0bV7A0vYWP92d1PwI1S4k0EjKezqTBEguBcAeoSQjPMU/kBY
3vkBOeXIKdtWRAeC4/bBvGb+m3UUxMVIri2mjuZTRFYTs+91xSW5j+OXMmqn2eBu
9fjSCyinprMHrUN0biV7Qo1Kla+nr+BHoAqE4BGHK/8r6nbQTzZ4TzejjW16ZA7k
w0dh8XoeGaBqbq8EJYlIvDLg27/ZQgaU5AuUnoClGNXhS1vK03WsX4sAGWo/beoK
Tbnc9FqCLbJGVnBf3ktqEO9yxjQYXbnF7MCfv851ouOYWcatZhEVkkHrNukhJwLF
ntcGZiGREA1TMG5M/7ozmddm546M1Dlge9KAupJtePOFL0icM8anlHYm+eN5qoc4
xMwQjyQx6ZaLjHAjJ1BcFsZnL5TgCh5cJVTW/XHdLvHExAmui50U5F9zp09ET4U2
G4F4b75cookuho5zHzmMuOdqUVeyN5hwCppEb+yJTRdFC+7e76BH+pmuttCsaSML
cIALcPtZvbgZn1qynzcMONwPizkzHJGyE4iHZJFUccNaLgqljYrUzdiJsINeTblW
WRY/uWNwytLuMJ4S+6FqQZcP4HwBHGgJF+wRwIla0yB1DKcw890AF8OwQrxvJHWj
ErDZ+vaxTb+8DZVrDmG5BCv/L978NLtIlPkr9Voep77IYCOF9ItpuwKbJCv6wM4e
kWGsam7ndQXKiCW/AAPL+mV1GTDipsWeU8sUaxT2hGrZOPRfJcJlkG6PoNDZOQ9K
wPXeYHbsOUDSIYjuL6UVm5QIQwNUzzRRAk6pQdKmBzKOnTTmikph5Mb0SckVnjh4
0fY1qVAyPc1VNjaIGBWBHQoxsmfgA27lIi+4rAazBBeMDEERLfLp89PFt0Zh9oxI
0jej7fkLDBeO96tJOFvsepd1BSlbzuib45eAHfZNp/AXs1f88J6x9hZSxjfGSbhn
xFPxfbfoAZbVBd9BBs1WL29Xc0jKpZGJFb0r9/rUZhsmA/tBSSnyGyVmjx8eSAe6
U7gtNX0l/Et5SGVjcxlv6qduMblmwAcJvmKOVJvG3WKJY5TxU42vX8SV0WJzAH8b
/biZq3XoPTYKfVz3aCIUDs51We0QFdYE8GRMZ+dktOcyvajyL1yPy3H/h1+oLl9T
bJ61Zr6ncDzpTlbwOy7ALfHwJvuj58iKWNKAe99CjmJ0mA76WqgqsEuwFdH4KDed
9nYIiprL3xS7greZquxjDJ4evY8uoeB/QkvF1T8p3HIWf7ciUF3dXLG6abkqgrYv
hGNrjy8BEMc7jeGiOFOKCc9AVKpxWiUDYYGZaObcB8YlG6MhwQn2OQnfrXAHux01
oxVlm2u78uOf/JzBklTDIYAjXTIB7lt1n4W8TCNV6+TvaLn5o3Xz/tIW84UFf+AR
1u8MngIoIPTxmpJ4lyQQTZCzCjqy8fWWmxI/Su2TRe921nM06jSM655sV+kXNUg1
PMROaaiYoMOLXWkIFSt4N4IbQqYxURMrzH46HlgmoMYbenS7UcAZqqezFfzLDVB4
XOaTqFQjFHX4oTaeywBJnGo5NLTCmSm1iOFwWe7j+wKpxqhGHMwM7oY/y7/wOEX4
6JktOTxJXuZzmXtuWvBm5ezqZI4E3AF44ed2Dj8iHj2LR0laTWKN+s62SHrr7kRK
MVothVMpGx2rmcYs9MSaRZsF2RORSfGr9nnvr5Pb+8GV01SEqUo0PQVp8SFOcpLJ
D7x8nCi0huWUu/Zq3ltk7pUd1RAuJpwHMvdWI1nskvvgLk8Ar3JAqd91jTI4Pk4Y
MsUs0ZOsuSpg07gcrD5pmcyrfGrI6qU6VWrDD1xkgxVCzaVJt5ttI0TzYUNq7EDZ
Kte3OOlrK9EIDtuqvBXercQX25UZsAtC+IlN+j5/FljMWzzkJUbGSB/Qy5SzAov0
6dLZS7UPOYJWZuL8AyciSnl+IsZ3Tx1aSAavlQ+A7t4Z1nsvYJOPtPIv0hlz4x+B
Ymx8dixD+P5AFS62m4sAreG59cbpkPVezKAyhnGz66Ben93CfjT9uru/2rIBBdxZ
NB0kwutmIp90Moujggd0uC1BIz9BUdlqgoh3xSU28OdmvGyXFGC6C9YCoZnzGtYw
c+3nOW3rvkM3eYNkV7Wp6hOQSG3JNT/uaZ970x9OiVOaMpnJxVXmMfsEbHp7ItVA
ws1HbnoY507Ev07IAXRFUP3xVD/D1E04PoXQr3kxwki2ANu/XPsQek44N1Zw4l+E
257pcXFqb8yOF8riUsJOuCUrb0iPCviqV3/JVAb1Rb2VEXxQEQOeC8GRYSsayGzM
EMaIT29PuNGkD2YU5hakBVLZ9l1oco3T1Fdz9nHq8aFSaKtcQlLYXLIiCO5LolU1
DW5MLWCKEjDSiQFVO0pguFXhhTBR8lWHobcyKAwZyV+5VpqxEGfJ/aFIxbHRQ5Cs
ow9965HWdpGv7juCUyq3i3UVQa8D+tFtvrijqQOR8TpSAe3Kbztr0OLKDi2cTEBi
2QvYBkXOtb06aDjLvgQ1LR9/8lutmYR2B0S1VSAXbcgHpmPpGA8r9m9JvUXBVDuA
trZyio61B5k+jreujIOjd0SSGA+FxGZAnw2HvxAYIvyL6Oy5IsMJkzOPQKi0c396
7eK3pcoEQDEgsKa78p39XGdRSDgVX1/wuzRfKa+hClK85nqrErQpdaiRS1gRgdu0
5lldZyd08PJC4Au6/zNwr5O/ac1G2TNLx+hj4p1xcD/BIbTZLEUNLjaCsXBlZC4N
/5YR6D4TqQRkY6jlQVGNgTsjHN9C47ImCzgVB+vF47PHnT2VftBZTvZr5MccWlg0
qbRc3Po5a7siBkwnRSDuLaJzBrgh0tEcQqhQbXejnb1Jb7KUHoxcKgaC1u0JbnX9
DubiRfH390k1+RtFOzoimxhGg9hrvz66cUSIPxYrIl6uHt10cnBPhAC66BnD4BNX
jy9y0h25UkkWviGR4/XHSVHoqTgUzW7/dHEomUMsAMp8SKoC7/2Apwnq53sNySab
E7I6exZzMTIlNj+ChkK35xBZgJDK95qI0dDGIxqfeiZwgaGIT/b6USuMe2Ex/o5m
TSBePHTTyWvbACotb/27JpED3P3CWN3RZubebhCkYXkhqU3KIfBLFCnbuEFLeEkG
PEQofkPS9HqRz87kZzgTVsYJ6nbQUTou8vYa3cUcftfnOeHu1G7uWS9yAO3ewL/5
q77q4+25DDVFN689TllZ4nuAkvkISedKiMfptUuTOYN5q6J5tFvumpEznftpcZg9
S9LOvYZs98arpKMHxjHroaDlpYz9ZIx8GqQN+5XVotjLXzu4J8kWWi8bFDSwcw3d
gd21dzVhMpzigtr0XgHhfApyqrm/VqRvJW6by4U2TWylBwZJeJOLJ7wMqWcsonJL
xHL4/TA0chJ12GYmacr5E2xGQSZOMTZY3kxNHtl/0F8ULhTxuH346DsJuv5RxWQJ
L5SoowjRqKEYMoEeceoUI2G8A6Ljnvc+vX0h7rrITYM92q1Pmb2oMbb8xU20Lwt7
kXrboBfDez8aijWjnh4YRlBMFTodLcXOooBwv4mmouGI6Y+sUtrWxvOxKXGxfpbd
8XkySW7yDNg9t/MpZpRTnRqsaOuHj2FDRUrXNW/VwziugoFQXDKL4pBBXe4dCZbJ
QZ9FRC3KBf6DqT/NRJYgtwsYkoMlsp8I6QHDszLFyLzLo32FyixR5e6gbuHuN00a
jMNleaeehbgR93qi8SYRYnRgMvvvPvt/AkBkhFiYiqS5ilnRyfrUaXZqf45X5Lkx
YYFIflR49hXH4jwmibqCl/vqo6rTvtwpsuJNpQEHvX9fM3aKxT4Dy/bq5PThJGib
L1Q8bvS9WPK3C7NGfa1uOdhWTg8jXTo2v2n91hTj4hn2QgHA+b5rjaKLYaMGB1Hi
kssILngXFTWuklrUscrOW6lHSOCR49fuchoY108C8Rls5J3b9rMs0DfWM6zgf/C0
PEPCeFx6gXNdmXLpvqVGRo++4KBKYXTu1SFdPHNlh7tzXup6T3t/UejYFqvF5mEz
vGjogj8aOeibT0Da+K6/KY/VmvVJUu/zdPAQkrALS6Wpd8uOXVDdX3uyzQKM1o50
svrE3V4PHDTaZf/o6wFuYDUmzhkvmCoOS77E6oc3UJ6/AJSen67W/qKfqO1/6VB0
KamjeDrt3O4m3UxPI0BhAPVMdCH5jUZJAaXZxaT8XTZxKfd/mrzGoxjBxvqYN3z7
2Bx069fP4U44q+4QTYLKAaYk0a8FYqEag+hQSmC8BqtupBSaWd4eRdLJs7StR05V
q6WjfsL9cMXpIQc+mxwrmxBCd/OBEvvCubfwDUNI4UL8CmCy2EYIpTLUXyaSC25t
0HV+u8wzyAMepz9Q5+OvyYZUjnPS2m+Msfld33mnPLM2uXAxCY56vn50cst45bVm
QlFoyLFHqB9v6Szwj2XgkkSTFQd0hijDV1ufZPKm/ftpVdpv9vz7s6nAdvAW/QZj
RLkb3ZOj6CWjr4YFgbFQ9L0616lqfG9QSTZrlGizXAC990QwROdX0eYHNHahGDSh
F1wLaG/ysvqucQUaVLZa4lHUV6gePcmqiXXxhgSy/ZahOMOUqTwh9gS/HhE2SaSk
l04UNH15EIW8o5aoeq6TPgFCQ7T3u3LlJMVMAt3B1y8/VEjAKVs0XmwifLJDYyEM
C3bHCx7E8ipH8qu8oJXChK57qO9rLOEEcYlwfPWxLOEvIl3f+bmmHRgeFCs/zTuA
HlxICRxJoAtgoPklIpdABU4phr+mVYhdAohBxf/SyFT32WOO7f63RRqrP5puS94O
OzT8nA/lGCP/iyrWqv42TgWducQ1VafZg51b6GM8nXnNQv4IGiHZUtUnL02KbEFH
tbJtk61bcwmtVa4gtndhXF6x09PZQdX3TfgNaTCl21ipyYGw93M380ihQukgcyBr
mH/yI4Uy0Psf/jmweoUTrHgbo+l/08jt5My/AuhVqnk8AhaCjUDNXaioVneYh5/Q
yJYP9BYldw4dZWwXCn9xJHxE2LyWW47qqV8Lwofnhjk7Y/j1Fh2AGEteWmtnS1XS
j1iBokfoPgk2paiLqbSQq0o14bFFi/B9uuJKAGFn/j71lDItqJ8TohbGmBH20N0s
j1zizW8KICRzOSg5j1SSSwij56q3xV/2qxfGVDmySYroiMX0BX5B5/Ql03AA2Rtp
K10cFaZhgUJuWze2zoI+vjtvC81+2ccgx4JZ4rktxl4rqHRJVTrI87FLLAckCSjq
nsCT+RuH4cts/KKRPV+kp8XgaMxpH21Rh2BN6GmOvdhyisVqk846SKNJWelczCMr
9CiwoLnhtoq2L94G8k1xShefa+c//i1D4kjtL80ljvIIvZAGJwze+TMb3vuO79XX
Im/ofEVSpfW25+ub7FMY72nzyY8/JFCrxAWZkFAmmo86nYTwzKvia12zBfOivJXb
v/KgyVf9l7uJFDCzSzkdeZc2h2fCNsAGdT1BWWla0gX5fROXrKWsv3tzsauPDEVN
9TGzovHWZq8ziy3xZ3dq2zZuLp0ywGNRvxdySc1e58bAQBQBt1c0yV0fLCms8cY9
w8WIYo73tdjZBdgfP1yDJXrIX0+ueoU86QllhoHW+4EnhMxoxP9tf4IBgNaO+PuL
KSQm6OOEBoJNd4tbWn1FR9aSQW44Bm/PsVS9lgDuomMvkDVZO3aOet6siB4iMujC
FtLisFG5HYzPrGaLm/oworOFnQOxp2siQtTDcfaJjZpNf9DFI/wuJUk2witUq+KX
6tYX61MwLNqg4h9kdLY3X869LZSS3SFGCR7V4W48ZRCBzIRixdEef91KcFG3qXT8
C1mazgpOLHERMj9zjByNxZODg8WWZPM1UngYiQstTqN7gJ0kRaFqQ5+nHLrO/xG2
PBAbkl/2BroSHwFC0hVFS3vHkdasp7Oa/fE7sK6K4e0g+9Ki1SOJkTz8blM3xwip
7ZPllYXXSEas9V7uxrdkivK+4ksz+hWzF6avtUwo8kmkZVJrsh/wDAxItgw5GdtM
Qf2rIoB3XDhsriACR6ALo3itKR6GcmXau7XbYX0UbbxUX9AiCdXksU9x+9dWSMKB
FnzBePrMl4HgnaodgQot0dPVXWf2omNaHtPAUKeF6X3XXnuymA1sOjxeR2Whe8Cg
N1NsBPVvkc5Ysarpewm+5Skn/9tstg9okHGtXa3hCaFCbS0i8rVw1mptxjbK/WBi
kuRcsAxUw3L31YyXvPKqlhVzY8scFLfatvDrVVB8QEJ00RRnXUy0oJcG23VGb/vT
WDujDK7rtSHdI/H4a++2eW0IaOcV67hmtP6V+MtmyM8xSPow6VT0ZI34QWc3y87N
Wb+EA8lmSGd7n6tpHG7hyNvSRMXtIWiu89ZzThFcUT8eCTkWxOwWbns96MB5i3NV
2DmVVub3r8b2qAT5ei4m09FqQJy/vZupt9m4KouQjXC9XCVhhWKDd9WL8uWR74Ph
XU1cu/wOX9LMcAjssnBEhYptwThk+2JkSfavFkConmiEXckPvBopKhA5XMgFFZ9v
oXE3y1svo3X96rFG3L0aMuuV8nrWj5LJZSnvlE2NWglya9s0IfsZcEjUeI2bRsnC
gey5cw2ENLhKGtE7sLWtxXDxkKdj1W2BDhy3cGXq6WYsbd33gNDXtTwXTuf/5fU/
InrOjHxundjGl126RluJkZVLan6PvbJ7ootBBake+unOC6OCeWLvWXAz3Zd/R3Uv
pxSaR9UV3mkCcNBz/1DVQGwZj5bJPjbMo/nUaZYCurcQ//WyG46ZpWin3jv2DRp8
JSj8zUUo00zRxt5napIbXP5lqSwKVA54BJNXKY5Y7WXCM7qkH8werXuQaF8w/Zyq
vnfUx949J0UVSlPzsO/0J+oFrD83DbF1MCu1MF+9g97JE1kL2+hc5FPxlSKWAZKE
YbuFjA7xR7RDs2RGCtvcKwKYa2XbmmX9FWXHVgOTRVmNdsG/mMEqUU6AVnzH48vS
ojoNerxVT4JDjGmea8IOGnS/eoeZTO3Hvs/KU42GeABOwdpbAUYqcD3mUyp2aWEu
A9X17XGDxcqxh+4rSiccEdzwmUSm+CvGl8ZuO4O/4FoJtbWqzE554eyA62LId0hr
Ix3uHiJ5HT+1pQUieSrh8d5dMXwwbHlUV4tdHbu36GOHd4wfwFln5/IFhPC0Pss4
7m6cTbqgUab8WDXGtasQHLfYTeCgXTtd2f8OYV6t0jpoCqRCXyFbJxt3YRph9FQ5
OpevtzeL4LViPQ8h82oVyrHeyJOqLalNOBYyuLdAQ4skLR0RZ8zf4Pv6GDbjVIiJ
+PKORjWl/Qa+pc21cdT+zYM0NDjQuc2P07tggbTMufACe8vqDFLsY3SFist9F1dH
dZYvjvY3FVI2tHRV7frueVALLT96qCLKIK/zeQrqc4sZW1NXBNiwABZ8bOJGMudP
DYHT9KVSdl6pHkgRMWPiU7m9YG1xRhJY9mQ55nxikiT0shTQZzKWu1d5Gw/hGegP
ZCUCkRZCXeB6JrxfLj9CNfx/wYtMsHHyvYXsDXRsEEFO6AsZMa3ICQ1qCvcCc412
55h8cVVQlr376rEbrUp1MppQkCYWgzGoh6uH3q3E0GKGPnTthgElZz5v4cW4Er0v
esQYaFgXR97QNUWNDekYsQBKe50UtxHUR9L8q+lgMpWlb377Tvy1uO/Xpf3LOMzN
KhR5ufiU99hyx55A/L+dJ8G2EWz19LehYFGLdyXmVyEtR0v1IhJ75XoHBU7A0uiy
F71yoYUDwoxbYlkkxCwYkKEBIBDy5xdFyCvH+DdiFa2XrAo8Fr46XQ45+L4XlX0H
z9SL8zinQvtoyugpqTMcPzT2qpNI89oFfgK30ePawjBsmoxPOnQuvtmZAswsYbH7
adoUsQAZd+c8HHO2IjTvDzCoWH4OKMsX5RbolXmRRswf0nZuL0RfnJtF0vZ4N7gd
1YhmPtRKB0hxJcoqaknNAbPPYolqUuftwl1H1E6+4OI+mWPCHUUFX1zKTBx8jvJ+
Q/YUmz28XQqZdLlO/aVEywj2a8Pw2iPTahL/6VGfcQs3I/wykR8ksMwalNxhI/RB
ngE42qyPRSJ+f/+JM04X1S0yXyAOVF271lQ0VJz+9tmpd7K8LgAWjCkD94yZgujY
QXYoSnUTtNfcCm+HL+/VkAu7VorY54YVWGPiBt5hzt5sSqAtkmLWBbvfQTDNbhqX
5rUUkRsBclyoRN3UJMn94hyKLs3uHYYqj2kgLBC6bDSeZWmUSIiOMs8NH/QmZEjY
0KIMdJgGsM73XtsCzqyhT2wxZlKBXQvOb4fg7tpt37Ky8doHiobthmduj2Y65kqv
uHOgun0A2J9S5Q6FlzIdsZasczChND5MXDTY8byT71Fo/2N+J7u4401+w4wCbdDn
FXjFDx0SRRHCbtAI04d6PiMUoEg0GFZpwUqM6MFktQ9lOYl3rmu7kZ7i6A8U2hcw
bgytbBT33f7XYBc9XaAQsWkiG3hBd5NsZ0oqubkseiut6P/O2rhh36Wxf6CaXqmq
vh4lCqhBVubkr3odRMAUqGcRBRcVLu5XsTsviEA4x+uyM0h/nL2cHAkiUCP+XE5O
/JJ4fPpIaslx//5Bg/2GgsgnBXAthJ5Mj693etqQb4L9p4tSPQYXG/QrcXhLNw6n
HP++FZ3MppqDy5pagJQb5Oj7436f7zSwP+QSV/wRElK3KXH2ToKLyTpwwN5Y33gb
dOrLEtTZ6qOuSafXWAP7MYElg7X6Bk9tJEGGg8dtYAUdKimN4IOnYqn0L0AlpBkX
7vskgkWi/TrZ+99cJGvZCl5U83UZfCYsL3btqL9fa+84GjugmSqkm+fFwoEXe7Fq
bygnNaT6k/SYBALEuFW2Rpjz1lo3kjYfUkkkh6N/a2hIectHqrpl7EA3IqAswCJL
x4zq+y/tpNiwo2hcPgzQVm6PY/jLL2da14oHwuJDK4dlTWDUIEF7PrwcPXok2FKr
9DkHDEQiycF6bD4vqs3G6r9SgAjybNmdXPjB2xiGVqZFZM1R3n/9f/3kV99mJqfb
u6mTjnx526PyDtIrsFINX/gaUyJRwW9wQFTLiuCkB9TxQm6UGTrknk055QZEKDWS
DXWFX+wFjeKDKn5noErf+eSHAOB3MWEVelorkJRAwz8DerhD22wgXw/7VtqgCn9p
s24jrymcWrgblQ6DGMS5FawD2CzofOA4KNsPHH+SKKXuHrw8hu7YNhlIcVqja/Wv
Bx09BKA6pQxETVyTjmg2U3sX9IZZvPTpvQ5XBhC7kMGpunNeOYr/Wx0oj2VIlLvL
ZQvghgNdhY9DhxDEAuF+l2lzZ45RDX6ho8XM2vm5h6U2BSiX17WXSVp2+ul0zU/j
GNSllso+WuCJIC0dU4lQKveN5JBMUPyJCMKizdPZOnzvT/A/mpmWs2X2tw0b1tjL
nFsxG9v1MLtdgWGZhqtiHBWDn0bTG8gb95kZiRVYtmQl0EYIaIAEF+xje3f5OB07
LNLK7hwpbvMQGjMiDMbXI1UtzQ0iqn5cauzyRnVqdtRZ4T9V+4DtDAS68pL5TKmn
Th5WA6mzZPiVUiMEgqnaO1x5OQpSnGfoLuMN0lYCh7d1nPIYrsu/OkSX8rce9w8h
z2w0M0sgabMPQrsDIfvbgyhFHiWf+cb9O+1rzxcStuu6VnXxGYXHjdCDRqtKLVzx
26FaiGXlH/8+TfJebXDoLlu6L1bVSxTfW+q9x6flZ4CdVl4bRi9dNisT6S5q09wq
zqjh9dUAtuAh/2E+gIgNqsqeuA6d06OOpnjHKG+yoCQ1BuRJ3MtvKDhcnojIyqKd
iPE9HL5EbyWmrS/dNeLC9ueinsnyGhOyb106tB0GTdvMNvt33bTvS/BnS267lTpF
NBwRPvKdxWuFkbolURvTI3hMIlyqcpQvdUAehNiMExoDkSPkSt8u662ugHTPvb9y
OO5anrEQHpck75T7kTYE2XPJdipaEwVpV9sBGlgIPurZN206+gwj2zJrZFscPBFk
Ua8fvyOl13RwcG5Hx636XWhPEg9hxHLW3futsEQHwXSKPGtRXG0CyG+I5lpae/Gg
zmxOwsfgH6JdBkRRmLySPgleBl3p7R99zeyGImzQPIdMZayUaLjN/oYWx74E/yHz
gcAPNGnYP62xzy1d98Lat3We69/NrP1xe9njMx5KXixbaMd+Wb+u+9sQmN46+4cr
AE7dOeOyTKxKdY5H0MO0fYvlMa/VRY676WywWXs9cdpTTCdMnMdgVLfp72cTeceW
rLK6RlEDWVbeCU8uxk89zgPhACjK7xuJhEueX6Mlk/Bfv0n5wgmAz2WmWIQkSwUl
QVgAFzhg4nTUNLbbhDMsd5Y810gi/0ONcDagItrju9tG6JVoVifAKS56MzbpoDIK
e1g35MxY3t+arIEaHBDCNA/n4bd5srkid/QbBxpor4cYfulJBDJoU8W9DBelKKjJ
rIIfqMjHn5MzzCoUjHxiEv/Zq2/9zgoea3Y01a9OWfe78XX7d0rpDLvBBEnFNO6r
/8AdIQQEFn4pNSml34FC6MDaWr+QFxxhSg9frwtD0Rqas4r0S1BQl+B7f1Qq2qlQ
QfH1X7ygRQA0Xf4XtvqFT1E9h+noLlpP0pbH/EtHCGz220m39sFT4skngA8mLrn7
a6wVyKVT4p9Y6/QIceEID9ETEjwfOWz/IrByRecf/gryLyjWepwXerHAsb+0tWQQ
Tn6gpYKactwVaOGtb6bREqigwz1ii3ksIqq2X6sLxmqfNkLKZEVqIYmJdgOI3s21
773ylEzoyeNzZJrNoW3vZvduuH/mdIxLBVAkCjvT9pTL/0O3RojbCNS36lPNswDn
dfBYjVrN7DVTIv/q8D/Vzh7+xO2CoT9qq1DNaB0Xbs2xbQy+FR8JaNVJ33NjyIpi
weRHDkxl/z5buQ58gPw1Kw6KV11Lk6LRr+EwlsmLkNDlMP6+8BMBlcIntI2og08r
wPoa6raSWhAa6qD0A/NpZgtJtp/wWroJxtBZ1ueZpriWbCLv2izUphLG+Pn5/oTQ
wWf2JTZ2EVPd/CRFy70Uy5AW0VJex53G0rYSiFnC+UzX8YDVxJeNhUJYr5g8E0ml
m6xNRfFGjByBBfsz/W+KRRCstjR75Txm26Qfja0lyAdaP4kB9dF78kx8xf4QCRme
DdNvZfGn0mZ0H79bp7f5+NFwlOU5JSQD28zIoPm0Ez5YppCOHkyCvJOOP7ocDqzP
CXzb7VYwG8PFoc8yRcvsTcqCHZxVJnEa8b28vYB4hT5bbitIXqWkd8us/eW4amro
DHdMMW6GGlgSHVL+7yb51iOGD55G6d91BoNUji0JOodJJs9DQKvVdcOoPzNIu9aE
NaJD8JhwPAaQfxusBcCDhmgOapTOigUMRk6bQfs177jwU5EKAei/qm6uZNSE1LTs
fKGWKVT7HNPQu1tgst1h/i8n+3ExDfJu+XDz4qCungbjAyuWnkyhp/0Sz7Ob6DKh
zoUOcQtd6k1SxO59Gbi6YVamRgZ16gLdUQo6zpqA1cXShNy5dLGon7Eq5NmFu+tA
mOY2b5hCCzGt8rFMYXejGgydwJ6NLiFMF50K8BUb9sOwSCTz9Kyy/wS8szwnsSkL
Vi00nk+BSZvAydRePPx+5l9pLl5sZb0BRHaEDJI/oqlLVWmYruBKLVlEzNDoilwL
wZ0Z7aN9J5XguNOlj+JOGl4OG97VP7qt/xP2ruoRivqMo0E5rmhmW13v7h+5pknY
Vu/Vt59xhZfZWThaoJaDe/43gNhiaYCUnzYpJvHJVRDrBwkfwUzt3oB6GdLBZwrD
dr8xSiLplC9dbdUUKO3agiW8WxjAFZYB9CzgWWFLHtJ0ggm/So6Gw80IijLV+8F/
Qt0NlyTBnMkU2AFnErcRmEh46O+15NPly9HV3ej7KX+GpM/f8thHu5MRCpXS4xK3
mOHUBKVfBZOp3+5+uH9hbNVwkdV4VbO77tin5fdDm2q65ADOX2WEUs7/pfoo3h2m
C/rZYMObJSWRlfo8DiTFGTV2bj9KR5tYQIe/XT0CwOLkhobjeBHu5bnYzwFoNP6S
WFmAXMK4sbr0SMPG7dWeVMK4Clvvf8BaW4ND9Ch6lVZh4IC1l0y1t06Zv8WXVHsY
BBrI1JZXyH+ZNiUmBuIJSBFe8+CPMs1VqENJNwkXDSB9gN5CE1FDJFUwEvjUvppa
JKCNcrUod2aebOvyP4F5SAucpqrPv+1VChskauNtMS58/6IHEH9xykud58ymCwhh
CPJHNVWFV2iZz0VIarWU4rmk2G3DT0fNU/fDp0nRqg/SkQz7mwqyiQPOrIB+HHOq
Rr124LbLV2KJ9Yxxim00GubB4k4xOc5RoWNWeqeTvamHtSlQxIIsLS/sG+jLMkrW
t4wAIEHFDi4SxkMOQa/8dGEqC4PCaW+XyiAF+NBFMQaEYFMsAXizuYkoA0AvHl50
ZrCzW/lxeMMJD9JRWYC055+dnEUJJr/ZTF3obf78dKE2MkQpd1UZ6LPk7EH0ehTt
+U9VE/s9j+OJUFCNQz3QE9/Dpg6STFNqSUCiCUyRraI1RiRaZCm+lk/oxDtW4Vpu
joEdwDnGZ2XcPMSUiv4uny3N4qWFkvcRUiC2UN0Jx7HR4+PsIUOYO9Oz4iYjDepb
iE10PnBlqdutTnJqIF8HwpYYAGvC4qO/DHZuF/bl4rvfOQsrPva6tkn7qPJfrBqy
MqzcbsOHm7BYXZ97XIWkFlcpfgVZe17o2n5BlBqQBysG+A7Vpxw1V8E4/jB3gCH3
CNH5Z5QkQpbBt7MGdoLHHzpYTWS3jANqxdq2ueFZuxKuIVdqMDmLUABlZvlwzHY5
WNJA+Tsf9KLXEUWBhwSZnvxyoyGCUOLFyZjgowmR3Z8ymEUNUIAvBi3LbZ+USO7L
qhKcsYqHxwdflvXg7jNF8L0b3q9vrGCmfxEKBaTAVGbqwf9SnC4uadZwUgpyeIFt
+OJkg5JBrVcb6htKWYh8IeiDoCLOK7nrFBj2Y82vafWQMUeEOQjnfrvBNkGmx9Xb
yReQiTCU1s1LajVIQsNmfNn3690aQYzWHI7rrlivuYr8x/6xw9k3/+ZA12KXmqyM
v0crINbuSAQgFBU9vaP2p/dpBTN+gDCaJp5Xx8iE8lmOtUYsknZheaDSuZRgqahq
eyCUZgKzwthyswbC0cj2YxsJd3jFf/f7YDuhnQp1qoPNk7cjQohpLmSnr6K20nGa
6/kZKsV0J54T1x2/cMMYFlO5O6cpXI15gqBsnh6J8ZRDus8YALK7ztFatvPUyk3I
37gr0d54sTLvCW95tx6bHDTNnGMOx/jLCyYCEQvBkpg0LueXkePtYqQHWtbE7BSG
FE4j/u2Lu7c1WrcpWXcBuUwBNPXkZ/IlFkwyoTl/ukO21xrkzEwnzQ1XwlO3US8b
Mcxb2GCYou4lO49MeY2PqyX+ypkr0Aq1Xg/A3RRxN8gi/87aNelPtQz/8Nql6NAg
xkHcrkkG5y7aw150/JlBUKmdeefCfYdil+8ku+NAd0S1tz5qWMvtxZoBw+2i/Jkr
mzBixkrDcYAkeqGz92UYtPGJjlRPKuTcnOKYYKUk66gSJ5A1ra83IOs4CMno0gv3
2zadrqaMhdMxFaxN3cyjOtpVYtHUQ7xP+J55oB9aOCCab737tKLAlNuMWLE07UtH
5d8P/o/HgYpcOV4iA0tLGxi9bOdlt4FCCHfXZGqiJd5SAFgjskCImKHl8MxRuaN4
dAaa0YYBC1OAVIWal6i6CLutD7JeGcMVGciDp/QlrPM6YfdJ5SnnjplNf8AZYS+0
Z3dz3JoWL5vXqJPQckAJekNk5JcrrYVQ8IgJ8LNwoZcNr8npwpoViBrNA9AlcOi8
ldUyGPakpIBmq45ZflXMyxnH905LK58s7+fuWHH2D8xGttmd/RyulprmNJI1Y6/7
StaI7fmvNeAbbLRZrBjCDw3JuNRAgnlAh2xBzOgWMcAbN/yO/5MwSymeSQLoKH7N
/6mC2KVZYCLeflhb/SOzKIW2js/6Bfrgr6zSzx7RDAJkwmKLgN8prHyXw08mCgjK
5A+Wz+HArKcEpf2T3v2PwikFgwxVMIXEQOEKAuvz7BuJYMKhNU0yH2liEeYlPKLw
SebEYctmxf+2K2Ce1ZVxHuA8KBLKpIj8cMbinCb18ytE+Mn5bI4Ccc+sN2DO6HY8
Bs1ydwNo32DW59nrCz/yjThJydhCy97D/zbtMYVCahnInOGlhC7sXwe4o3TZEFfi
9p1W6AccaxQuE6hVnFsIGcU7sU6hHo31pvRyil0kyKLEz8KtiZ3viVw5s57XYT8n
QQO6iaXpBZ3cz8eVS/HicuaY6j66JEZ72Cm36G5uB1UXbMA1kxIhF/Vuy/ianSwO
B7rCOiDEFSvtpiJB1BE42Fb2ioqNrLwzftaGIyQA/nsvxPUUv6eTsT1tqrXEL8wG
RUMqN+ZcbRFBMoKPPL0Qe1uJAihqKo6z/H5sL+6rQrk8DH+KNCq3IE48ygXvKfiu
8ECiEAcxIY1OV6kQ/hWzDFDcviRhASvMtTnL9c1XiK+LVIqMMFnBsHZNzZzZjkpO
BOd109FpHo1cDIcMsjWpidYWzVUV+rz5LPou5C+F16eBDzdWiGXc+6SAMaupH5dJ
H4rBSB2ia78HdPMmrCg6nUrQltolMTdpHS/i0XPjVu+8jBFh6IVBJ+mg05wAGFT6
v6GV64kNofsQRFVuYvUcBOpQPH0ZoMCwQ987R55QndOuCKZwu7tZdh1s8U1/Zu9H
EKJagqMZpdyxy6G+sHL4QtTP5AXjznFTfaB2VXusvieMwlxyNX4YRAJQGgsQVaa0
XiHKfxe+qWf4JMmfO27xmvHfZtdugJgkpxcIMH/BbnwLetbrKBl37IzuOId4gjB3
BK9dNXzpQf1hwkdIOR69ijcdCVIeBw8QnqEcjb4GHOwY4/WBwu1FXE8UVsJzPVGK
3ODOgP+6zMvXMcVxKBv2F6I4VY3+XpjsN4p73HFxZ9FrmY3cZ040x+r0Ako4MrFm
SW47PdHJSKcgUIH1ktrD7nn7JVR07hXtyDCJhjQ3uevG4GTTIERUD2xcnIS1O2XM
7k2HoTZVz7XNgd4SkeWzhaSwTff8vSSbBPd2fSxfU8fHv3bTRCJoqvXQe0iHMvS4
qNrxDKWO9CFFFvO7lIHTvegQ0KWTgPiVoedan1RxQOiE1V3Auf3zENlYG5o9gdF2
Wbm0fEEHoXFFUTFmZdPbjXzRuNDOMuMyp2cp3wbly6GGdRPyZArGPjadduX8MMAQ
qhl5x1RZFaNQmzyec9zgKqbMCEP83rLG6f86tINkjajabmDSxMm85fMyBw/OyKlp
60Y7/usB9cMc6e4qSyb0u55IWOjoaqPQAGd1OdE8iVuoy1oZrffd3NcNL3zFzuNs
O4dy24HhZf/fnLO2nShi3H/f/ndMMv8sb6Cd7Me2IQJAuH+GWcQHxArdMfhYQENh
TJIN5hWin4tA9BLfXdSmOn2CD4MNRH0o2Nw/lT+oBiFsHJglbxkAR6XEwkerCC4o
pvYAqJTpSj8B/ZL43ril8lf+EcXWYGT4KdDLPy2wlsfIpNlTeuu/ZZBOcGmNZYcT
3pGy/hpvbSaUOy5MmZnZtBCcNZcu5T0UuW0O6jHgf6HVaB7ks0mytBhK3pifWRq+
8wrzkI6z7MPXdftNbrBIHWWWNxnJR5ZysqfV5vcNq9FIDdLEqYdOzWxgcV0mamkX
8mR5duCZqgfFh0vfhZxW8GddDX8O7cHpD+UQyTc4/1YMuJh8h9v/7x8ZELMWBA/M
eRaZxZKyjHo14snOE+vKCsdHPlQy9MPGqlS53Yi6jsnIvmPnfspeNEHAv+NBYPkI
MRwT1z0PfrzuPn1g0tMwVOEowSPwNjqnD8PuahkiUaac+324kN7Ji9dCC1U/7eSR
2pW/WmWnXV8mdaHnYZ6LePXfCWRc1dnWsZq/J8vWW7pq8yIstrBMOqGe43horXEI
3wRNTzS4IXq9vSc8p3ix8RDTVHYLt/1cBFNTFeOCFynl+1hPL2lllOCB8/DGjyTV
5y5uq83aX5gkyT+/143Y0vB5kXbojWjhDCq8wD9gpWi0W9S5Osvzum7YHOQTeun+
TEylsVVNNOahYXnNgVcbBY/c0d7+lJiQ3nPEAb8i16U0/pNCB78LwvHHSFbygz6C
DL6XMV6WuCwpyXC1EjjHOV64Vp+dw5EJIICG2Z5yEtcno1zrLGZEi9KG63yZfJH/
Dv6ipDHIoPWW1EW5qRu8vBZGvoDSjU4RrQsDVxfdWNCpt6PcBcMiavRHXZLoctxG
jSij7ZRJ3TMQdJ/DfHq9PadkciRtQv/iElNSmh95+8dIL6bgkT2Sydh1JOEm6N4V
uW4qV/xNWE1SUwkFIeUOgd86/qNob27fzqYeEIVhjva9lK3Xvatmd6EZy4bbrMTt
3usfa59RYGl5SEnctdOxTxK2mIWqsYLynCwGD18wVz4JHs3oMBK7eZm4P8c4O4Go
tGFG+LvBm9zsVCCVrWuyw7PGOxS+LaIdTaanMuUQcOv2DE1KvBJTukfyygwvcELB
/g2JZkwjUEt82siuECoAMTOvwzUr4LbSoKnPSI+/QcVcZ0iIsCiWQAAKSUeNLe19
n4Ru3VkiAsowMjTyU8un+74Idx9lgXSF/+SB1iLJgJGahB8BMGFqA6np0BGIDopF
VeOBX+mg9MQHzwFyykMfzAwGDYJ3C9VZgNxV1+8WTo8R5das6PYWvy/dTtisbtYt
HX+c6eMxYdhtUTf4edo8HfBqApW2ZAH4WxtKuFexwc45fTv5p5i25lCNRp4ItIt5
k+KfYFNui+XYEJZJ3ZwP+8OtYToAh+61FKKOZigltPT9JfLu//IxZmBNbNfbruVh
EHESN5aqEwAebHn2XwZWJ1Or/UwlWl8jtHWpxSryw3fMxp5PWK8JDb6KLmKT/fX+
s9ZOk6cr3lPxO94s4XuaTIYrR56J2EKW0MBnhnKvEjKGwH2qc4TS+7QhAwNSsfgZ
QgANgR3ExSeN2h6zjlwt5K01LSpokf/TAuFTJAqepZ3bdiWJL5253EROcqfPEWDy
CreL/MjvQkpkJ5QjMoDTM8xJWFPLEPskTX+TC1MtCa/NVy5wJEOPcDjSdwUt/YnW
i0Iw5cMsQRhAbLXLQI38uZ0itQQ6eRlACIZRDkYGdx+lq//pkmipHyPUyKO5xPlo
oAGb5QOP5tWYEthA3Hf4Ms7T69m2XRG3kYlmRAiBGev9XzMRj8qxU8X/k00Lgt8M
3FdGP9bu+orv5YoATiOCaIN4OuKJI5ijFa1wVEmj8QcjSeac7CcLwiYlVIia1hDF
yItKzMfqZXssbAecgOMvDwRzMSt3HPJKrgQ6XvdEvuP7D20e2cd3KPNY4KNZ9ylv
9eOZJo/lMYwglr2vO1OgKkWmRF6WdDyUyi/TPMEage4m0yLZ7MEageqTTeQ1HE36
Gi+EiXhEiDcIIeQy2poMn96c48IDJUdz4f5layZPv2VT+UpWujNGHkJeaJVEVk4B
z/Y0rBJr372lvVrcFYOyw1pLms+WI2Jtbg5vxSo2wFo7RaOWWhWOW2Y+L24LHqkU
Rf2L1y+QSEZziOEsMccgf9HRBF+g98/bHzuxE1qUUQE+zqlo3xhjFhOeBhVbovmu
R1A1S1vpCB3u7UB26JpXXwZ3IfatfrNTWYE/Zg6eNQLsUq8wdrU5ASjrAJYpt3k8
NqLVTB7CokWztTLkzSi0ngL09gPJghpeTzO9W+e+Majz0h3KfXKW7sM1GnpJdFy9
XFEAnuWDE/92BJOYHtzDn6imrxvJd+e4wauvrJ5vGCL9QQ9VuzMWRrxnEe2rpOFQ
3h8VsNhOCyNxmW23sINVp6algXkf2hfOTd9E/dLE/+eVfi5s1TZWB7tls8NJq5X5
EQymWIWaZqYJe9QOPONl5zHi02gWq0uTJdd21caTMKKVkW81Paet49+Rsx0adR8i
ueTTifyJ1lS6xp2nv4Krknx5P/IO80T9TOu37PlYc5CsF5VmPvglfUuBPzHKf/fw
qaSBgXMAVipEsOgYwSpZQDW/QlvBd1M8pQpcFeQ/Wz6YH1SIIUxtTlXDMxMp7hX6
lf9gvajiy5BDNKnTqYeCGR17mjP9hA5xnpgzUiihz3tFhEaBU/6ZcrBSqdR+3347
GF+4Zlk/OM7ztVxZfC7sMjZEC1IZkUnvPLFh4j/1UtGdgAf1lEmVAPrNv6h3r+sW
yCaKTK/SGGQt72SfFz/j2O9IoZ6NQkEuY8hvDlI8i1qadVnDfLaFYdGwB10Y6XY/
g9HzOGA36hHutB3LWJrfGAjpVutpjl/yBgLBpZLnAHBZVLqVto+nogrfhL+hfaEj
K8loqMP2bTE/smhbFcchADSPcSBy+FxnAzpfBVuyOc/xpStyIL0Bgb1tjaI3SZGH
Ffa4eArvpHwofe0rTnxyOdEbbzLKsiSrECSNY6OWIwEENO90TGozij/DNdAe+no3
rZLIz0BjHq+hSiSSFRU9buwdzpaPGqL4BsaZ9q+evQnJh+vLPjOnIlIyqGFFMYC8
zDUX7uBEdN6F9UKYdQYeB0UiWxsmcgn9h5qhiMj43gc2o+zt8hwsX9R7qPENPfBU
TuQfLC1Tc0J7Jk4B315AMQ28s8IgaxLv2eX0A7HKDE+SK5df93ZLHg6DCpsTqZ+E
Ndkb/tc2dd6jnLtuKjV3RQU+NNQ42IJdQ0hIb0BnzlIQcLEKrGn3eHVXy4UNLONr
0926Bklpv29myAS7mtWBZoouAmc9lg//sg0ZfRGlLzrZm7uwU9jd51l8YshUsiMx
2oToHzbqU2+Ip02uvExRsixefpYm+mbj6AYNuzenfgnrJPWc2EzIzOguD90vJFNG
ZdfyR7FJ4DMrXgidBwGeU45S39Us/4vYcjtZt8Q2ku0bRxcsCAgqenJrtDzMGvap
YvHgoINt3D0XJeOkZgSorzVvGgLml63NsuiMMFORDz/7rYZxtKioS6Zskm0D5FfK
qKlzx5DIRSnfRAfbcp8a/FLdnAKh71TeVQ9R/d7hcMiDDXjBfX1eT7OjOUkWa+rb
PPbeDirwmwkX/ZQRAMyUBZfjcJp5pxOoHbwiEH9HIkMWOG0QgZG2zDeGaP5Xis1+
UkfokTub+OF6QLaap+AYa5dsMhldkgJPAjg3Bf9wXkXUZI8PZtQQ/7+V1Ob6rVb3
gkMgqLDdT13K2P+Wp6daT9fB4UsNoRR7bLFW4JerZGyAwK28Loj3zQPljhgOpfv7
cxg0QWjedmMjJbbr8Bdg3GuAAEn8RBzHg0Bgk4bK16QelN8Z340N2awL0P6afQ9Y
YAu9fs3RaeEo8xBKjINNXWgSRn27KiJhBu/LkYl6wMYkhZhVQpFVoYBdMGYVsdfU
X2/6VMxIW1sAp9gMbyHdoIpdPKPI9sxB37plUsLquJF++g5HkVxNmBHs2EzIt4Gu
wyhmzoWqNCuNskOqxY2O3cp2ClP4hrQNEZuwF5KgCPo3dJ8r828ancGRGB+LctFB
x2QvNGwQOAY4n3j7HICIQYuSXGovEZfn9QIigkxTqt/jvC1fJcGjN9ou6em44FK2
LyPr9vYQ8GoB06THg1yXPuER1RWLaEkyf7rXDM4mTNxREekuYBP8O3Cz+stkJKrX
81wwWe0ab7DO33jyiMoFrPq9QMkKDZrTIzdvqGpHHeYZPu55hzhukrJRgvWQarRy
YtG5g+88/6R2FWgCx4WI27NiGOKJBzXp3KQQI3ohoyPQiP0rC6Pv7/qfL7/rDMTb
DGUVLx6BGW5vkVRbpqu5/nxaNuzMzRTd8J+4zYUFCjUt5DGvjZEiSJ0iXmdl1mK/
Mfp0OXSotfMLotRXk1L0ZDgwhY4kwIwAVtes8W4u47xGTTPUXvQ3uOo5uHCP7RbV
Ic6HMC1Lrlx2Fs336KaxTvtDcic6WSC0VYIoNs5suCNTm/WNMQ4DFUujrPIWCp2S
Ifnbyc0eRYVj0HAu+CB53325h3tj08Z0OlKxMGPE1gFFWLJYOSOm+FvdGXC4f2dJ
lbDlzvW0itJaRrrOqfVUYnxz9HKQMepACjEAn+2KhsBeQiN9YDLmZlNLKRyKZ3YQ
bNSLkEG4L9c9Z7EDsLlBd/CipyLNrnJnk/AKu9ol/n6dPozo5ZmwMG5L5ed91c9e
H9zF1oLnQZ0AnlwiNPT8H4FOCV/2KMUPx46WrXjawa0/cnmEGRppUVNczjUBL65N
PFnassGaB6Uaes+rW6tS1jWrAPMw1myxqDjLKh7ZzLdmwOn6RjIis5MBanFq9xwo
wYrPI7/DYgeTg9K4oGbkt5pifEcq89rQ6dhSnaIc6VUlNLbl4k9tkFYGQ0CkfA1o
eFPLOCq/gwGNU44V+LE8hDhZqlDjilIOSD5panGLqshGD/fuvaQihUFjGBs7RO9I
xqNOh2Jy+wqTsSxwxy+iVJ/NwqXbywClD6XHLtsrSVBBZNH4IO/4sqLkZHZsRKQX
BN4SKvzL1tUwZ55ye2/A89UA+eF4GYPLo9yNWKewPFC79XIgDQY+YppctoliqL7Q
OD8mK/duEYrZT8GoiU5YKNORp4yWgrFF4Pj69Zte3nBKKDooWYY5OpVlU5rceFES
qKO8oieXw6VGZz8N4TFUvtJPEPWL2Qig2RDg5MddkiyIbm/cYZPCFzfJ/mvTfNsy
eF4dN64KKqeJBzo9Fu4WVw4clIbC/YtIrn4UWxrmdk7R6fduMYwXMnPrX3l1PL/n
OAW8PzaMT8RIr0IgQ3pMPTA8xT/HpdYs89Zrl9rcqfVZ7g4y3ggzAuzG1whfW5y3
hR8wKosWwnF/OoPVHNFZFpbK4AVH9Nm3VleB+pXN81+GYd+A/tcFeeWX6LiepGRr
xMr0NTcTOUcJHAkuDXMw/8ZY9mUQYltISz8JPLsx/d3zY9yaTiV7i8sLDTNT0SbF
E7vmQe2AHj2Bu+yKO8Te+pN61Af0yp8shitlBR+Yvv1gPd+c//cJ1e8vTQu1oBMm
QEmE92Sd95K6NTVeF3frNGfO9YkZiMtFO8bGjd7DlJQjfo+YzHHCZ+1ffeTTFHit
N7p0vrk5ExSYjJA1UgpJeaylF/LWTTdfU6ZuoS4B99/EoTFnhPuQOAEWO4/5xW5w
UiY3mY3Af5puCSM0IWNRUzTTSlhk5lbVQ2zShNAfrJWS8u/yVmJ5f5pJsQnxxSfi
vYxePjhAP8OdC77rqsKwMxb4h4DsyPGNrMIM4lp3S3oi5oCMnOoiMsHguy2D96GO
chzWMA/NcaZ+M2x31gGYVRjx+aAfHFBpv05nAUbat7yob5rO//2s+wC9iBj92mV+
9RQpb9fx8oI2/9E/tHupw3HsScjuS/4O20uUOfEpwkJAcifSOQoNq/0yg65HqYuw
ZKrUtirmAYFL0s7pB4HJmhFVlQXZuGfAZmBkrqQZuDqxK2inzT+Y2tr8WJdCC/dY
fom2MO2wpSX7PdGWW9CpKg7liW0q+4EfQrXHekvMPKwjo0CXr4o7raseeY90OHXE
toUoylJ9gOfQH/t6hg5PTa47aOpiPKujvyvZDqo/yqMlEV156aTOe9s6dfSi5sZd
qF+hTSeWIsIncuYs/uCOn2M7MQfx1E4aPrefmuJSCl2dC1XTLfY+dPQYcH+u/hG+
U/9z3tGNUz+ueR5zKgXfxbHQLtpGMQ3XiOF0pgKgqRNz65tSglTMyqTlZtnUBCac
PuBzgeST+sTsrhIODBDNCMxIDcJd7pieX6oH6lMyQEK6XIGFTKzBVoGoZDf2h0+E
r9lppyy1DFZwjh9ABi5C7UJObB+9Ij7NjPQTMAjDU9KuXv7dx1xsQXvt0NIHatJl
U+T4evAZ4C2hx098Bgpn/mnSp8ZV3eE1VPlnhp5Gkvy/vFOCWrm3lJunwRNhblJS
wKvs4O3hWe1agh0zysN9K1RZvvzvdj7qJbfMHO1SEVKT780PjOF/G2fSiCk7qexG
lqXidMhP+BuYK+h1RMbOiOVu2DzvBqpcZFCOYZEMwxH8B50OBJ78q14FPcrB4pJH
J5FdqGMbpjmmZkQzCLKhQ34n0Z0LjlkFTtly/nu8l0Rc/n7jlrNPdfhhOFTsm4/i
UjRZ5MsMyncl5F3/Vx4unwdlH61Y/DRlOPEb4JINtGJjdjM0tfjeSqjnJ0OXCwHg
rGU7lLVzi/9OEThPdPcQzHJNvIqU+hgQAxUBgUr+dcW8DVDhPjdnhmxk0iydDE7K
bHR4uiJ3V1fAIAnHLTmFW7f57PUNDxE6n2mjv2lFIwSwfY/hiYwHrhubzlQsNoOJ
wXkdU5Q10nqmKboKZGTluCRKm/+kukkfYXs7YmKGiVQ3150uVZhRTuZ0vFIco1U8
babi0pv182umIkk5dbmsiNNcg5G9FQ2hdhmMRartuMIbBhxg/rgBJ6hbDOfZBnST
EeOyRMM1+GwjD6WHF4oQL2hhYjCiuXMjTfHFfVRYxHeLNlA4/LujIqsSscey8DCE
TAzS81LyBBscbNErBQ9mCz48546l+IvMlMWea/glX6knWUrYYMVjZR+msAcisjrk
fF47NTetCi+ogXXq6wuoWFc17gWMiH50rwWlAMfRD9uMmfr96TIiLwYvv2gSfngr
GeaENNkFKjl48sjHU95yTNI7gIx15a9zKHRmFTd/TK5+d/NVAYIlck+zn4vw8Tx9
Bwce9ucC1sLA54OL+jXqFBbxMcY0jHmMZ9CF7an3p6k+A/neia6CDHQDUWV0LzLq
/qkGKKE7UijlxcOhp5PKaYSeg5DWBSkoOytaHZmaSyRRt+3hAyRpWTzGtMl2m7Qp
aobXFMK5Vu0qdcnc2KNKERLJGlHEHxOJ8b0BYX3N3LtaNtdjM6fuYLbASdkTTBqI
a6IPUwZQuVWP4KSt6U0G9bgUDhSGWQCW6FwtsBOx8PdK1uzsq7RowUdEy/k4NWjY
gdwf75xcXbXfy+CjZ1QxVC7ACujHXikcbttvcBhqR5IFu5G+KohXuBG+wa/wQoJV
qocT3iYyf3XVTM+vhEY9bMX2tOlMgWdkNNETDI8HyJMeia7LU8+EtPlkebInYb/q
oDOl29xwWCtmNIjwCWnITNr/us36Uqmywz4qEu3b0YYwf8po/rbrLnrjjiwWwX2R
5T+lweiqwxBWUOaEJkFrZPzLwpmjy2lF6+3mh6+rzSazhZYUUdRLpj3VttNNu6/l
OXRD5awTp22dKa2YqIeLkscl2yKfbxJWTPRAzBgghIXrKY/S1H13ADfhAjUzbTd0
f22F6BNQmtva1u1B18zSw201kGHDWEJh5qdp3jK6KBEoNo0bnwcYhbYR88H4wZ3g
2gpbceBKBiWGVRyiPjodHUBtmq7BHLil6DwT6SF2irr2qwFhYFuY4lh5tcJMdwf7
/x33gFkSRO4Jsp/VRH8Wfg+YCIJQsWynOlVu1v6mo4/NyHv351jYoLL96uiC/bZZ
ub/fEzfazjJLHuOIkcInCqcCa2YTjLQtjSUmIkF64vcNEIjCeuEoCL2LLrhf5EBU
DASNHJfkWdTATCKHL618YurnJyF1q2zs1sNOuu7T4lV40EMIxutioWouWZfqvQKb
qkzkHgDfOUsJBE4CPVMMbEGswAEcPoe72xthKZ2/6rapmkKiSZtTUUjRSBJu822N
af/gOmQ9h12v6uHFbmfuPdVZlPv50SuvAiNchu2M4QVDQ0rPWYwP8Q/wqnSDQnvu
MmriZ5jLGLQteNafBoEMvczLRk2mvWniWkFGF3p+VvVtFMHpOOeOpheIwBjfQ/zc
vLNLpX8svHKAoE+sfxjCot5Iwl4GSYtYg/LjtEZpgLFOA83eAehCL/i/4b6Fe502
Bnz3hkrHhOYslnBkCXWoD4H5hVxwE+DlgXaonXX4WuvlyXsFRyxA4p2hrA7s/JDK
AyYKfK0Y9gRFCAgCgEm32YUGncAJq0W4utN+d9AfD7RTPAVXMRD9O9YMxYjAL50b
Z8kBSro5hYanA2QeiVqWBzxVOtn5fc7l029qBiqbzzTtCqfPAp4aXzkMidy3Uw6D
vtMXgH6zwQvnIdOZnUQPQwDmScrzoUp6cYmNjTglpvtM2czn/N7J8HAmp82wZgi6
IUfPwyLeyXpf+OVZuiKbgCfKl5/AnT1W85UC1KLo4ms4kczQ2Pn6c0flmkkrvqzu
QNDr2dat4AgppiRtZEmR8pHc+cdzk+ErAMb0k1SMY5gWz7yEBGoFaADhU/6YX4tC
xDtXOLPMuqcfTh1Tu0Dw3j/h0HTC+PSWhIu077RvY3X7nJkezE5um0ho4fGWKvhC
9Hwaw6t4Y7c4CUpz4Q/NXkxeBGmJPIKw1PUBDHpGow9jBeJn7sISi9Znq0N6PtVr
h+snglN5HbFoeO3fscM2Kud6aobLaamPJ8SnXxVx9rMjpXBQLky4ZRxH7zkIBzDx
PfHIEiouNScnLFEwNzEC7TdIRbrdnp0VGmRPPPOmhYdbHzogIvPZBFF4z8QadBpl
Rl0h4OyvYf/NNXS1b6iN7Whmk9+YOJa+7XVl9OpQc3ZOptmUK6aTlu8bPy+41GNS
H0q5vnVmdZjGOZzveks7VNKGYe9Ml++PPTJn4IzAbSTDXq6V3561fxOvsesB80ZZ
w43Apdhb4oqcVq21sQ6mfWDxj6pozLc8pGbYxvYAzNzKozlQUISmwzwv0pQL/VBP
BGGOUdO2h/Bi31IicDwnz54xnhw4avK1HIsjW1afhsZ1/LVAH7U/390Mw/3uHrvZ
s/c1dgx0jGgULLlb/Gbdz9lToUEWNnQdv8S1PMiUYos9/S5IzTJjcAnkMMsHO+iY
DCVknc7B99CJWdwxBm0Gn00saS7nD7YXGb6DtW42FdIUVQvMA+s2/wEbeSL4rsB1
00i5gSKodLk7aZqFfrsqBRvP+1soJJ5BVRKS9jVOt6T2i3r6XI1WqIbhv1P9bV8R
hR4QntwbZ8gQ1/vm24XKkbXF47FdLAiI63Zeko7JdsRlnMkuYFXAP5mLVyxbikiE
V0yJYiDkomvXTSnBB7yGK8LRN3l6QLOiI6fwXtZb+y7Me3EJTxRWB/7vRHPa5U3+
L/+psXxVjdgw3pWK1tb4T93ghJWozrTVZfxac3L0HVPVfSdZo4LBGOXHBzAshUd3
DGwTpfTaS+7EsLFoXnDwsQb2wTXSLA4nOc0AzF1wHpyzzxvR/FDqAsOsFeQBhJ6q
y6A3AJ45Bd6rM7KN4vvMf7mvv+mG+jYbYU1VPdKFA1OyEHsyH7vzfkUfahUnySJA
0TO75iA6/ISvNh0I3hYzTKnIkaaksGMSCRrkQ924c468IS5+8UObuHTK4m9OE4b1
HW7hwOPemO7XA+eE24RBMycPOy7maz5A37+p0T2fbvGyHeiWD75qWmpz88w1aQOj
TcYUn2ucd0InZ48e4lNrtzx5SE4zab6S97m6tnp26+5uWSGH2OwGrM+7b4RTppKD
c8TCxmGyedqAijRr1P1nzf+8EqTUIGyizKWV4VuJJoPZCt0F0MS+escF5MGSNNwO
cxfYQmPzR2dW+RyrYyyY7T+dzUB0eW8tW327ls40dMfuxIcAtX0FY5T7gUzgnlsL
blIbX6tDgnRUVzcSe4wlffhyjc6z5UpAwg4Sfc0Q/6zZ4lFXmaa+1LBOkiwk92Qf
bVSg7n4LmYLUVjjgBI2XjK3aAx2LqqMXUuOA4B08351iRtE1njtjMUlpvsPJ6Xez
ygsuU2BfuM0h4HQlh/3LRrmYgULvZmpt8/GdYR4769IZPk53Sy26Enmr8p734IVI
WpQEbhAAUYTEKhkdNgsH7qmA91Kbf60hjFl8DR2rU63OAoiVgwiNNH9ntnzdgamw
1dvkqIBV/AuT8tSuyfaznWb9h+SoMNVzf2EcYkItQLz7lkIIit2sCD+XwcroxEav
OUfMRmSkRf2gm94W49b01k6Eo/l7/oIlNwOehuNVo1JYrINFRNrs/WpJtp84gnkm
tOGQde+arg6flNdDwi+e7CKaBoBeF3Ilr657DccTth6JIStbuxGMdel7bhqUDe2d
nvuaSPJ3e8lyXFNK1ZuEfK0HBez8v0ey7sPXrQ6MqpeXVvcTRqruTv6BEYUF+TEo
JjCUpJq3NbZsLnLBe3CfipsaMtpUJFBcleXhY/7R8Obw8XjcLQ9YCE+FNxLyld7q
zTZ3V4RLZE53zRBmHcy/WOonDxfrPMq8bsP/S9IBVxZk4AmJheJO99YBfbK1lQN2
C1zHxnvHZ98rEQQ8GtHYu3XKpHjT/tyhA0LMn/rH+CbnD32HeLKnlu5/uIl7RZBE
JhgGHQdhVxoSeKiizuM4eFrdbJMVXlPFg3CTR7NVOKHdtjGMh7R1n+YqL6+fEdX9
KgmqJgD/zNde17/cbtwHTmUbHso0wCUaHF1wGJ1d0nKViBbwmpXMimMXpgdHg/DT
7XLnzzsHpzEdfU0WrPbQLJP7Zji4+PLwP18FLRayvZ9QusMBHbJtVpBYbB3izpmo
t6T6GwF06ipKdFOeD9L2ckuTWSNJgQdEcWrHOnd9eE66N3FWaJ9mvMSSQO7Ppzso
5okvCpv4jj/k9ptjCdgSInxPxDpddyNPyFkpGPPhjfM5xR3IFXgVoQFl1gsPtlWH
liSh0ZDTLNOdPF6Gc6AJkGqPvfmTg6QOXnrnLFqyG1sQ+WxET9J3FKrjE5tpiDD9
iUenrdT7+X3fZPD9vcSVwveOrPBeixmqJnOOkC42oqllD4s1dCQJ3B5/D9Cc6nDr
dselYL3nvjZF6YKUvk1eF2LhTwfJJTJPvbZ9afWeHTTEH4JYZXIJr98j/WuSfccZ
iKiF3K3T405AxNKFlvbV2ZAiSQwBWERCMb9u0hX3AGE7f5nSn04TCMk4thVx6fhh
gs4Ib/Pkqb7LxjQlV7N39uqIwENVvXMqkheWrTiMB4iFXKUl0zwbj+ByuiPwX1lD
DiUjQgsogtY3DLpSfvEheRkuYfHuImuYuF/iWkO7B9pH0VvDCKDlBqgFbZt5xvJ3
4uF9TDJcV8yliIUWslary0ug9M29z4kf5+mRCHrPzuAf+6mFgxoFrvrdykN45dam
/vJ7RO3OWhT/RKpBrOeux6cHjpPEyO5uPcxWqOqRj838829HRsUfDO9RSu58ScyI
aCVoEx/tkZv00ATLrKB2GAeDgywdg9qSLommpPxYllUA+o9jWk2GVYFUFuWan8H6
m/1dA5eHIs9zLdQNlLZibM8iEupEdM3XKIvPPnNm0twF/hAhc+kMqmQEfL326mpc
sStBAoyS+1JJ5ciCEsL4rfTN1DPrHwLqvxrktdakW9t8J1YTYjWAxoKinxaIoNpe
Mm2Wlxu46ggNS67AOHQltndOU37iGFAxPfzzG0ejrBK/09DQB7L6euwmCkaHnxkh
SnCRT22042p0JFMeKk65hxQIVRibBsjlRvfjUMUkQCzC2ozaVj5C9ccjSAwI+mB2
eVqAVMQ3XjMrnFesIGeGIAQIffQ5H+nTBc/I+K2jvwJM5/jUIOXKVjMKgRpEDgOB
3SsH+2A/oiY4puqherr48mhTaPbQw0cRR2GHwCJWAdFvrKfF8S1E7VC6PratLHyZ
N+Z8p0V84x23SH4WojqCUyKPvahXDt67pm7NEo3wLIcX7taNGNr5jQtXEOQn/YCp
/YR25M54NVAgiQ3qpzhlh4iXz3M/Iv+761wjxrzStTP+8MiknZ6eVuKPjKwefOt1
qj1IcF3r5/7t4L2P66P/TmalmDDsLfBRcO/NlLxJJoEQ3OmFzXOiFh72QML2RykT
8IYF2od+ABLDRPOvZNeKn6gCKWq4zBLlVNYh/jCb72oJxVQLOheChWTf/iy5/pp9
D3WZJ5Z2wEu1iinCyYM0qhra0F3RRnGE16kF9BjraZXD3X9Cspq7JyVzF/Nlh+BV
6RmRILAOlQPP1TUzc+z/ePc6akEaNrBQ/iCgkfekIKH2Tqs61knX+eA3xRO5ES9D
SyXxGZgvnbgkY6zNFkyMsGjfcXO/+qRyiAsVG60090kRmAfqx96xRaB91v2nIBv6
YSNRY5heSMnU7sYUDj5bfDpcCsr2kFOSdRBFpUyAAOC5sDi2QH8CKYdGpvhpBhfm
zqkDtyNSiT67V7UDAG0mAUkRTD5oqP+SvlcWkRVvZP082+tjApzBLCuIzDS4SOg4
tUZyev8GaCmmv+muiCM0nCfErGhI3KyUq3PLmMNfd74F7yOD8v0/P2pyA05fvniB
uVYDCClIy0sCKTMgxu/t5CAl+wjFpWYtxhtHrKeRdYIDXReOehkqs3uIuB8YXUTI
clQeD+nQDSQIENAIG5cbP9/jIkpJlYGvufb4OxiE6qpnV+8Hfjs1ykfbbTL7c2Jq
JT2VYf7G2IrlRB3mkHH7ns6x46VDTbuGYTtp2hVDFeOWKtky9yy8wc6enDWUOyfe
dLbFG83eQw3T9ZBamGN3jO79OIOdM1S44c0AGGnKs0cGXkBZiITuFg/W0okLy4cA
BdOOrKxSw7Whc6CuU39WKKQMaNBs+a0kBeBm+i6UFOO1poObLYKD6V/6zD6eXEG2
YJbxecuclWGwJREQpBbCPmyblUvghT+DJ/N38mqe7f1smYGfq8RJ+UmZNFBX/Zb8
ytFOhcsB1LJqZ0v/GpyWcqq8zLnBNoyn4371JevevVcmc1/5DNDNdjqz5WbD0L6W
W7tvupG6VVmq+MMgou6ZPuhqy5OfrCr1b7Jf186mBjQWHZQr3H+MjM2NTyw07xsy
/IEKAh7CUK1gXmhIPGQx4cJoXN5kGx5zJV4PfTpKNisiE1cBxbesIWc/7KcGxKZX
jQpUJXkbld2dhKTWG8uV9cj07g4wCufEqYfku1+qNtJjA7ZxEqp5viYhBENmkOGU
Jim6l+NO5+e4MoW9yK3c1XqHGD4rGvPm1GyqVFurXiCJPFE9o7FRlGUhJvNPZkW/
tey6v+8Sr+/HnaztTMU66u6kV5tkZ18Hw+PiVx0SEiol45vuasgPVCM52FlWM8r8
LadhB7/XZWizd4MFNMaIxKG0LnpxqynbNBkV024yCBK9vekV4a9/hVKtIKCahgQC
+Ykxpwz0YIXPTt3VWnJKhpxrpEP2Yf/unWCZL6wDeDm4yc5/fL1IJXllwdCd5qRy
PG8rtvnDhxaelWqQu3M1PvOmfDLSj3CUxKa+gHaEMGVZ0+NxBxGaYf06wvZxrnF2
mLmeR3Ne7o23VN6utKBj/uqjXfNeFR2APZrbPsWwrmA7FL2RpTKZOYIUjf+OmUJ2
OhqiqICNvuDEm6Gxp7aK0fuJlwNiCDdQ6vrTw8Was/NSJN9fWMUA0iS+KDFcO3a2
/8TT0CDjL3/Ayp4CgMJThxsYiZikvl4UYQxd4tchX1WjEchrSnDM5NjLiLGVStG4
8FcCbTQSmkekzkZVBJjfKQJPMR4C7vvj4zL3zBlpcM5CV+fi3EwDa1dplWUMRmuG
LwpY9BawZ7AI3Rrw/+qesaJCvTRkFuSOrQZBsmvd1BEhsqaIlvY2lZpo0he12dxY
wxJaO/VXN7ApTw8uZulEEw//6xaKUvL4bk6hrv0zgEP8OM1wkST1BbGI5ngIeS4B
t6jIHaDwLqtFABZrmvl+0zpYEg0YOkCPUwj/coZVxaOtUeQSve0Uf0ZMRbLG9OiV
CAQPURaNJoZcDfw6uB+oTnwhOTTK1b9VjQqf4RmEDiElv2R61QYXjU+RIgVUclm5
kPdw06a360fWv0HCyEMezgYQ2LK7blETVk6qNN5OCCntkSXbALzk7+6sk2xmMDx2
JaNo60Sb+0XHgwQ5mSJZ1ryRWSTPtHHSv6OLrUxxilE91WwV33GXh6dfJNNuZi80
i4h9x+La5czzc9TXIdlD8R7NQhU6jkhHHwqovgEMTWpkma159mcH61iA63F4q6d4
O1es61tvg3o3EvLacTaI9MH4GHm86sKaA+BInlNrifx060EmLl9lF0gE15dVAW7t
/PAVJhz3/YtEioxqw5EEKXyQVR4meVQ1mJpqNcVNrUxz3ooHKWSjh6NuLJgGiC2s
59fbTX4EyEwOdffJfZkJomtVC/zHKWrcsERN1Q/tF3X8BntsWEtDP73TdLNzS9Rt
HgJNaFb/XWcSEB8HuoqQB6AGPKnHf0+DBPmxqSuH7B+nj+BJzDUCX7YiYaCEevhZ
zAU5KqfYa+4xfNIMmlXjMMnm7bBGoUf6AE9V+LzrIbYG4jEK5V77b0rVKmTpMI+D
TXOvqJ7wORVVUIdrOH66LkZFCZahduModEmM48IrtA7vkhbFbj8h1JqwUgbzAJnN
9IL1R4MCg6qSAdB22TQ6y6usc/RcCy0U7ZEVEjUG/moj7HjfD8pgjq3lHekZL5VC
jsD70OTHxzO762UbC+jVTgNXSluqE0ZJO4DGeA3yih7a0NHZxoHxnaS1qcYL//ii
H0ilQns0vtXk7Mjngm99NouY5whXpYtIxqseODsMqDNykyFC9kXvmNwvjm/nSFXE
LArzlXhpph0A6KHBR7VD1bdx4T1zbIO0wJD/yXBApweqwfHiH6SsmK++ZJWVQtRg
7z+kH2WWN/HLmYch/7dlxOv+YO9tiXNvnWsRXvrNMn3f6ua3+hq80QzOFtdH5/Je
BlWIKLPGARHAG+3vKeVRn8u+c4IDB2wxxH8jrX7hKaoSsXXn8VMpBQnRyijQiOMp
PHHf0BwRmcVxzJwvMn8bST4+Sv9ru45PyJpHv2mqxS8RCOAeCKmKqhyJftU/2AWF
upoMOzVd91DWLbUHlarBiePM5GzzvQAy/dZCBQF4tj5pXHAi8svoJBS37tmnikQQ
kWi1vYNU/8WKcpQhN3GyAJRuKDDZ5wQb/m1DR1ea90vxlD9EmHwxfe67TgiJfWMs
N3YOX1ZOuCIbzlSn+AVFA6JmipxwbH+GVcpL3XNuI5GFgvkR7uPVKIobz3mi3nq5
SwaSI77Wi725dnKxmvBjm1O8H4rPygecj1UVPBBLWmTdxqBBJCUM3Xs7fNmSkayS
Qly32PwGq+fae20B/jOxMS+ldWOyrf1xOFTKWlA11rGy2nC7cC+6aBFK3GfeginO
iXkjJOQCnsZ7kUGU4CGSS1EOg9keDi9sDosT1lW+HBGvxOFoID6q9YflEEjEoKPA
BDUR7xq/MWTrfTWVJP4O+yVlHZxcqqg4i1eJI1sjaIfSukPyX6CXTHwSUvvyc/QT
Ie814kV3zLhCHbSMi1P+xQx8cr6chwf1ge7d5EwqavSTE0cZIm4wink/0g215jCQ
zAvPzII7p5c0rxvxBcmtFt7K1w+P336c6Y7974WNutnc8C+yMkX//xSHKBzyBqMf
6UkpFlGUm65io08BGpNkl+2u9iW8WvpYRI1rFpH6Ppb5HBUQ4muyv5Rq5nfhjvhl
w0XrVGrsolWVilnMbnO+UNAbb8h38QTdsocZ0l1erDp1JIM4K0DJ1M93oCv9coWi
78apIVv7n6lv3OIK815Xpvna7lvaghnlzmQpxDmNuLzwds08h0zyisEgdHSGDa5a
mGotCfbrkQZ8lwZAK0r9vKw2OhQbPF5zlT7V5D823Bz597dROPIZ5FUdGlIUPJvG
yTkJEGYZT3PR8r6IQQCtuJPQTCROVfhYtnJxsB8Z2T8oG1MpmzfO6ZZ6rRpVWO8h
NCWwf7aSYLzw9pfJMyfjouBimDnAul6kShmQanvAFv2/6S1Sks4SkPeSlF4M+29D
j7PUQ7I6kVK+YT1z6GKfkFye3+lYSAJdUPOBm1JZPvvjL9/06HTewcofhxCLEn3+
5+9oaGW4Zsv4Z2GKMlam+WENJnuk8n4FYEqtzIx8eIQulKI0/7E80fZf0SqT8L22
FluS/BLjQSogK32sL2hCA0YgOYK6m4oTu2v5YT2g07kktUpRuNIhh3Bmgd9yrAiy
tRq7QbdurjSLnLokDIzh1EGKI2/TWsXlaomigVwEmona+2lU8SGc7AWlvSWI8tDX
TkDS329J6SdNr4OTv03vjryGIagC/GImFobG0rJ+rKnHr5U56k24I6ycwRXn9Jg5
SBYKqnkJpN+A0DVAuuZxiIinwn36+4Zj6GZScVkHonJWXlRpNdrBJka5WIMebA9Q
nr3/ZPm004osU0kVLUVTLG4PKmrvwPYPWjxrqQqOxtmmJkVWlsILUdl0/FnPkRUs
TJyeGt/7Ow/FHGC+THRScjZQw68+Av4qje8TJokF+NbfeR7Mug/Vd7gm5Rcb/i5Y
Y64P5WOBvUOaK61CE0ZJZxG+TjkX95YcguPp6jmADSbpCpl+4LlnnhIudiLh41B6
y7b1bu6le7AOklsVN6hOXfeARsdpeALjv74SKuORzHIrfRqW0PoD6b5+Nl9z5Ciy
bEHS8EFiUPlWbLH9zmxZWQMA82NxW4E/fnt4lTahqCUq9Mr5yB65tGSch5jX8wqO
/PXwcRYqfuWnECvAJ1tejk1IOqP4td7CbivO+AoB0IAeObsvZ5k1y5/oAITqIBBO
VGpmVGZsoh72E68IdZuppv91w0jZfCTx2+8DUbjgdL0Hwn+hpvwMZc+KA/rO5EST
3wL9V7Y6p8A8Nhtz1U+0X9pu9NE5dn+iC8zgeVjvZBPJFPPPDNFfn9xoQkzhxCCK
MJ6qPjU3FE/dPt5ehfzDnJMoCk/2hOzsilzsqs4RWf6Yn/0KdkC2UNSRzSNNqR5A
3luimbA6c5BVyaTx1/ztSH8CCpnuUhs5d/ldjLpCk9t6IQBKTDJ2XIkpOBBpiCtK
wc5ml/Z2vdIT4/7qhS+vgR5o+5Fa1TQa5oWBHy5FmeHMxB/hRTvXnUdMpRLIDJII
jl3Tce1TcRIqmxh8NzRVu2dPhSwFqyY1u82QH7yy/FsF6OpsWW95Yh4wYBLwK/vk
yt1lQk6GZRA3Vhi3CKsRiuj5Qf/3dbv8OCh1w08gXK0R1+/kj24t8YO/0Sn7Bypv
rwCMWeNO+kjbfCX8EYjYpVRG6B0jimlLc1pmegSrHLql3ewEYoEa+kRQtapaO+8f
0T2f+XH6sxi2q67NscFYyZBJaWUXEoMq9vCM8kvA8dh8CjwnYoBcoGqCgFp7ez0B
/48le9TAFgg8Xqt3LeAaRx9UtqVTScFNFFaZp/7MvLMB9mQGYY74Htfdt3SgyWPU
VcB1uRcpNHihGbvVG+ZEl6W3YpUvwQ5na+UfEbMvx+1Dazlr/IHGzVwm6KQ3TRSV
e4/fn37lW58TtNH7BQNs+GfgVj9FIIYiBVWgfifvXy+xvEBg0GKy/NL84/BvkRSp
tJZdGkBRxPbY/rdfi06PXT1xAlAI5knIsB6KvGl+qsaSDmvUuv2iRw8gtCirQ4Sh
4qni+yQ/g8RyPCQRGz/5xLj5wLc6biyzSjjnQJJQzTY0mG7mrR55o/xZlriPb37s
AiwNvmNzxqDFYdaXdSBBOHAue2+hCbsyD9KBYn4AL+OAHhfc/zV1fZlpU+5NIRIp
pUI3SCnzhX72QxkwIO/qcYltseZpr6KYPl6+vg9+C2FUaZNT95i6kxL/2p4OqV1O
fJwhLVHiv4NiYqZoWqrt8+ngWTtppESDnxKPHOPCnWByR4U3Pk4aciF4Vu3amCpN
UijaG2TvlmW0MitQR1W9d54AcOwqwH1uFkNV+Wx7zRo0lYkedHkjpGmUUWtbFwMJ
IaiuLJ3fEaiah60SoinFpS1dHOSkr7ubZOcY/Pc5WEtdecNzM/HFT7emWk6m9EXx
tB5uaokUue9Tsx3a329Ks5W1wIk7oxTZV7ndxWGhYRNWlvYDIliSvn9W1bcovUkg
XirvGMUvYVrtC6GhwpmiD39DN2HoH2B50tBwupg7Y5HOsMfesbGFe76anupgn3Eq
t/oVV+68CLoShU0DrfPxKbcmfCz7wrDHOSfgSfs+6AU9ZIvY6/YZXU2YV//X/+BC
P9t7+P/l6hSnj2jHA6s35rSlQcmvYE6ReXVON4Pzj54miJZghqZdoJclFXmCX6Lj
GsHRGuEcJxFlHR/pqwzTlEtZmYA3555aaVn2JghKByDpUNiVxlZBNgpLZ7BNjJWi
4L1H0kYkrJnHSL2/8xeFLV52PWEFpdCkfMrFEfQPqwYmkmL7y+D+Z3/dROmRgQe3
qjOa6KzHlGZd4y5smf4vkNErfPbEfNgn2kMWidOeJ5Uhpi6BfJiSjSwsH7w5XWE+
F4Hs7xlKTw2aGZWxBZNGgt2Ld8qzsG+91pm0wyV6igeDzJS4Cc6915KloAVKPDzm
T4wy1EmzkYqVbyeY970nhkqJxJVUM+13go8JipglZFpE6YoSaPl6NWuiRIEBOXB5
XAoaRk/rrF5pGFX9c3Bmy8MytNzCmTiTN22H0B9taT+T8uyNMOyj1/OGZDke+uc1
NDZb2fBMRtQgbDdFvLGcmt5J8WWIGZ+R5vUkBBfs9A4t3TdeRz1xZ7UQefPSTjhC
JWJQmRWbKpInkdwOgIGV/nw5Vl9VkGsBHxdwm+zeGZSIv+k6mAkhMp+nAc5jFC5W
FaJ3tFv4LEnBRg/yRsw6wZ5Lkp756deuo1pklZzbInNER38/haJ51TR1qei5+r0F
wG45Cv87JBHP4hl7DwQPCqUX73fNkHYZygH1dYHn91WSQMjhDawJbC7/tibtHMwO
78eZKCIVlBck8Cc3AeHtiArfMuJ0ADVkHH2lDZuIo+abtV2DgBL3ZLLd4FMyUxX4
KwRPiESBQPhICMZUZakzJDdGMt5WEvra7EPGQMRB0GUVNQotaS2fOjWPIfeOGxD/
UlbNFzAXYCIC3VKYEqzkLiJbhlpPqNb8BfYxu//8Ol/A/vlK+FudHtv+I6iKxqE5
cBP2ZivdISzfGqhEul3rb5OddYClRZvaXBN2NW6rMwOAIdp00hhMDYXQ53Ott9Ps
qSWj6Kq1BtYOCQ2gaNuNFWpIFbc41V8n4gAm4+L6BE4wYCPftFRXm2aid5pxQOrs
TLX9e5XBhO/XCkiEiqq2ABjraYa0Y/tFM69M4mwvfIBdfGFZlqHQzHofBPVoka3u
SsoYKZz7OZwdsZZb7po2o1K2mgMwLSCVfEzmzVc2h8+/8ZFgLYE2MUFxpEH1kJig
a0kbw4/0M/tm+mOVci0WtvYsi+rF67F6dRO+aLOqS/OySI+Omqkl2rXj4885pHZD
iLmkx9N0DQbnXjH3iJFDp1+F0IZwuzkBJefOtHKM3neLQs6nX/R7z6z5NNwPO/bh
swq5diDXanOdIgDhHJMcFqNmNVX2MfU4F4w5q28YbiQ1dnEykQhc7osb2EFnUuED
1d9AzeWRHbYVfKOlMz3nJPEGwdlGFl3GozopzB73AZiGJS19ogfzPxSJlue/iIsu
ZyA9WCyeXbQXZl5pF49w3Rl2fbd2kqcp8gNSBqu7O+KX02Hc8xmYHR9mNK56St8Z
tmMb3XZ9D9uEs1tzpiugJ8R3QjvOhie2J+rEDCO1ATKHWCyMT8wVlumekxGf9fo/
EX5jKtyUPU7oqnFS9vOorRG0LxHvLTS2IZG8Gf/C6V9NQYZbAydWmtfe0KHzcoSc
S7GGyyFbCd90AODirimvnDfIUfj5q4m/n2PbXVtnvO+U9UdG9jFaBS6YB5D9UJCW
6SWOpuwiATZgZ1bp29A0fGKR/PzESfSSCk8lW/MQw6MLF4p/E5yJJzfJ94BrZfac
k7CmC7Rs7NBJIER/8yURfc7o8mOfDjD5/DvzkLYMP/m5K8ap6iJM1k1JpMRCrHF9
ouLgk6RkteqgO7V4XFCijHnXrDuEfZ4OCfdYSq30X2lDKWLBEx3uVjnroL2kJ+J/
uEGlqlUZn35dOsp7262i0+CnJMdY57we9agd0WkKV4uDE6e+97i3VWqogAMQjNDq
xEOx6YXFtOXOHZaM0eAT+ZYOi98XV0uy5F8CROUM+8PIbpfiH7J8vvNFtMOym8I7
2uQA05s+ngzUEori0RNoqNNshdm5gi+phZ8ckET0R+SwOLjnUkE4yz31+3foze+V
fTmOJtkefg+yvXAO1JWTXTVCaU5JZk1MRAIjFJQgT57GV6mBllzC6ZmlO8pTmF9a
aghyfS1MU0s1sCMT7nEUe3p4JYAY2h6qrQzyfDTv9a8uRNN0SJ3fYa+NWnz8tGDn
SgOFLLctcjaP74m53rb2jbnx/scGnDf030V5kIN8UXHRzEfhvuCWPKawpTW9rdxf
1F7dXGLZXw5g9qFwVAGw3/gtfS8FwVjbuE9CnxY1WNgoktStUOF1KUZsKL2z0864
AV0DGvRw0eRakbEal557mfLTVIgQBWC9YP4vMWlk4+unX63ezEwbefC0LuPLCykk
ehMQrlueD2iqR7evjC9f3Tm/LPqlLnFRVpdPjDoFjX8YaE1wnNHwupa6AXVjz3FB
uKe+Dd28vF5V3MxV0xP+zIBV75JlOkMV+MSNGg1ngjgl3vKW6Q1BSOygRb4Dovcb
wR4r/1ReN0wNtMgC7T67vLrn7OcUtKzjaL9+eVJvfyRZcBq40lBy/tYZwJlxX6W2
rZDes0GiWtWw+efVzZXjZBI6LZweYTwzse4UXczS8Nki7rhoP/wro0gA5w5EKaOF
TV2VrMP4PhgaRItyF+qqORdTEkXdbXe2APPTTXTMRQNOqEUygpzOMR/wP8CwVavF
StaJ0tUgTbhSl5iTpko8ATTGMLswh4ht24oniTsjBxA9Bzwc6Y7CrddlxbU+Vx+o
5TT0sY5HiS8zoBYgOLmJkMAXkc+DIHTV+aTt9cE0AzdwhiSfvDP6QpU0h9r544rR
P0gCB3VjT3ujYgU8EVGehgQbI2d/MHjVFxi7FdqQvo2K1RfRFMDUF4o0OPZkrzyY
eU2cCUXYRmlUSi/pWfVhxGAQB03TKRWYkNdKUPyM/T7gQtBTuLnqzVAu2bi7eOby
4/+mRTllxPwgw7I+Nt3latbFsa8NgATT9BFVYguVbAE0xPYs6B/sbNxBVYxMd+zK
AJi4QEEvDQB6ZGeY1SbT8hWP6UGHvAgsF7fmRai2255SX2Oe49QLteupnv2bBvwZ
JGZf0ARCnkmiYkwvtGKEXpWT9+LHoeoPyAr92lCsTpdkJRl/XSOt5q3dpL8158tJ
a12dxu+BWGQ55t6mEQBYSsYQUuNlHnVoJbLtB9Oj+mE5e7DG/M+P+4eMJNRsWIic
xE99EVQWZC4S4Kvs/SxjxnA6bVZ/liyC1zayrNBA0OQJd2afFzGJZ7dkY276Pohz
NsYQjAbTaIn3JnQ1cetCHJWggATVgPQsTyK/PX/oz/dFZsMcr5YFf7kBQq14uSWL
AdjHxLfrHAmkgpXFtWYCjhnLuKOb5E7rmIVPgw2VoL8fku0KXmE60+lD2ueVsY8N
o8T1ynllq9uuXbtDtcTyl7khsqjwOUQV779rkcxyHXrF4wNladIhSJuxo96vH4k9
meEkRjKDd9p1nLjYmBFX46IXH6NbHB2/xRFcbRw07ihyUicw1CZhTD/LMrFdZIVK
1UXiHd9OtfSQvGWfYcFSd/+VStBNWQMtaTFaH5vs3qGyPQvRNPbqGvbB11eTt+ni
kPSa4wErcFVC2yc2+UWu3WQywOXjO06ck/9CkQqJ/fmx5d3tQd2wEASCkiuze7UO
mxlGOWkxmJjCID8NEGVWqLryzqWp3REPZUAQSTK3LX2OQkBUO39Xl2qjeVlkgaD2
zIU4Q27iKv/yXDhw8lSIBDhT2u9z+6xpC1Jp+DgunUnAkRry0i93v1oN4a5FJmNn
XazZ04qkyYbLJDF3N6f1dYYULf84UK2iY3Rn71Py1V0BeivGXE934e8/mLiFPITo
dEQ1HGY03BLnEPkKe9ns0vDIPK2oC9lzVMLWYO78QEyb/W3lFnmmERDxgU29VEkm
3pK29aK4eeRxrvaHmpdjyuLnLCObn8Bvam4Ew5l9g2stDmAolSds7LLHaDxBNSu1
sPfqeJovgus5K+GhE5bk2To82Co8iHhCrY9mqRgFubuFrviW53RgHvkeIm8jLnIT
3mv6vA/byjvomD8YdLpedUjIzZzp2w9bOUzbIwwDOxI48kyXpsdtnsX+p/6f5nPa
3I3xlx04rLb+IrH8niz8KSd5Do8PIDHEYIC/hbNg/sGG2vP1H4pb7a7/6I5+8Nhw
7B+XcoMg4uelmCeI+lvID8IfwDsU+7akvelb0KTlr4bFIAmThE1cyhkm354YG+X7
el9s6gFXfNix/6mjZKSvK0sewyqODybP6p9dhz2U4QIEeoy07ppbETlEjXZXQ1vV
EFgGVkqI5dPWCfmYQGJPAt0UNvX1/yLqso7vnbVqQBn7SfYJSiUcLy/pcxDfVxsd
RbfmtM2kjNn+8lxoufbBRW88MvOMB0OmqlvUapW5Ckh6YYmLe3vds6vrxKyF4D1P
k+jaOtCy5PLak+UjgkU6/wCM+cBsNBn5QI+YtV1T5ty6rxtlXSNUZUPin8LDLKV7
oMW9FZtmWwQXP+MANcEfPfcISysCFaFIo/M+t2s0pYOTPH0aR7N8HZ8dVsLlUDiZ
O6qE7FtA75yM0IhnzpQfLpXGumvF3D7bJO8q1iMHchswcQPPwYXki2yb7ujG4hXH
CYbdSLNkF66yw7SNS6HNrfsxqez0GAircs+WTtqLZnOyZcXKhLlgnCF3WWi/uyZy
ng9Vu1dKXEpGDJwqZjyWRHtN5wl/02GNBC0HSiOxMCea87qItCZVDjjni0FJGXir
MtVgSXSG3tXcJ51mxyxKIAP7Ov/yrWk6ilTh4irYGaL0nxzwpcGX6ekzgbl/GWDO
rx40KvfFZ4jWJ58A7/aTHSrp1ZGJVQt5o21ZK73YtKZYs2ij+a2tz3nQORhCznVR
g7OIkYoFdrYEe+lKUDIsO/2Ioiq/+/9io6p5WwTRqCdDTYAWLliP6RUFFMOTrP7P
QLtEZrufWLxn10SRtfZ193kWq60adlxeZRzYxUnhBRWGdmeeKyEBZYmxgRpajhRQ
2sNvZBv1ejZmDj1SbqZM4CsjsUi3V0qTpvW3lFsaT+KVEohOWJMdgfJSF2C0RRDg
cSgOx6BPaN400OcRDnAaEpK83t1w16zoBq64PGtgowHVky5YZZcecXJsEi612dRh
7MbY6T1UgGqV02COSrgXVTB7ChHvNxpLYNED/b/6R7ZAbu4AGKsvyCzqAKv2zMNO
G7vbPR+p63QQw91kR5NENT2+Vuw4qKlC3VNj3/a7vOwnUZi3Q8lFcOLpqf605TNd
kZ0zFG+m7+Id0puVfTVP1r2DlGbck1I6Vzpnp9f5cEaM/gvp2y1r7I7wrDLN61QA
oJQONb9VmUA9p9El6tT+USle91XTyqz3YTNLtVjKNajEwKw6v7caa7GSh6p4IymU
pkdWk1mLeCEgU8+KRvCwbncuoElyRqh2TraEuC7grHwnrtZFzKx8zPYa3abI8kCD
X52lN6ydeGO/cejcJdxMRaKT/3Dti8evHlOSBiNbd8mkXqraYSn0SAb+ZRiEuEwP
Xxmtm8d2HdO5uX+SDP1NqHdDxBebmuMHbhUFxAvQRQZSPdotVnz4pHV8ftwq1HoW
mnpDBYVZjyTdl2Er+4i78/8dDHwl1SSgKGNHyDy1EVKNZbY84CtsrFn9T5y1sm1b
RKUU1X3qQ65k1vfkLbrR6hkzUF7uQz9PdNgo9PTVD4l3EN9eJKUAwZHQnc1VUE9y
o5mol6QfbtpPey89JZo/NmOzQHliMKFYc+SLHX9txLeowXI7SVyqV8cWgvt/O18D
rRP/8eI/QdIc9Ig7lQ1NYQigOW42zK7RdfOMI6QUI/If9uZtGODSIptK20FxkyDp
6pP3s6KKMrR3FQfXCknrIPlj1YX7Ilusxsr+L4KH7hAzRgaXr0GPMK4iX03JK1eZ
makcjMZEvQ6jrMr4fkitko6isbTkWWQA8xnl2mEIAaZtSpcMYMP0mjf9UXYhduPh
ihbN7LIkfOZ3/gbP1rPsQvzRepfxV4d0muxuU95pmPKbbHJB1tyg0rzBBCL8cJFa
gke+uhYDrtKP6N6r/huu96BMdLwW65lA3yoJoYaHTJWquZMwPwR47uX3iLLs6Otf
4eBazBHCGL35+LfdQjrGe3abz/ZpDt5apQL2YQgzhmCuDrNIcU6lMxpMGFcq0yi8
fl5kOZzBPtnz2jpXFM4kYCMI94L5SAcrF4jAltscuxsJtUGsw4aftq+bO/SaiE5n
m2/gYE9cpwE2nZrZDdBYsTz+Zi9BfT0JUN9rd5C1wxVAB7KXq0XdQK+KWvZ3+J9d
FKyDdL1oSx2GwDkPxYO0BQWBMthDjJ8JyJvGIWs3Qo6ubt4GlLy/nC31XF/PghFj
N5fH/JsIowkpHJnKTCDROBjQHub9LZxVp6MGROMXelOxhA9Ze08XxrjuOMrTA7XO
aVt4E9+MUEJz7fPZy6TQQ8WxBgW2pTRC9gPUXYo28q8VbkCWsnQwCRhwZC1HTUVU
qb0gG9pAHgTR1ibk8r0cMDxnK79Ro8fTnHDP8A/KcghElowl1t6drN/9Sev59Yh7
MVSB6n/yyCeF6hJaX2feS+BSvh8bPSeXNfFFBPkY/EHs94q8YchC9fZwNmTq9sEP
H8mYn2TEImMx2xw8Gb5a37caLp+GEg5CF0wrO+BYbIlrCNyFzZ3J+ozXbCBvaUiY
pLe41sBVM8yuFgHgX+OBhBwoWd03embBmaPkZN4idLmnZaG/9OAf2LrZm0KPxVOx
cOxnBT3Gw4PgkEbRfNzqNg8ERqp9ny0amRhKupEkChBPdsw6s8WtjYwVDhyWpEoR
rLAIi+eEIQlYAx81xSlN0imkBvK6Eqdq9ZD555Mx8iK07ge+CQCxkCE2saWYecJo
PTijx3siODlYqPon4Dsk1FnoXOsUODoNYgGd5uW73z64xnnsfATQjSs9/nyj6orc
4TdNUAX54Dec4nP4ogYSOk65kFmZyxtMJOnAihltZPmyCvooy4o3u0Zbycg1NxXl
aSgKryhGLn9MmejaoxL0E8RvKo2WksnyprgLIQGlhgTjM870tpBg7w7kJmcJOijk
yjwkKCEn0RWnUbvVOnS51hqZOjPv1+sR06foICH2oqCpF5j/ZWiUSCFbucOzMuyF
6Oz6QH3Gb6sDrM3oRKm5LQZ407EJs/HcPw6ybWyVaHyVwddTciU3Ap4MDW8M6Tm2
v8H+oIFVu42ScCFHhBfavz+s1vUZ3q/fi3hHqQRSubPGwn+RPtveCzsTtDd0++S9
l3Udo9p3327usBQRi2eqEXTpJJ4vrD0KLWhCNwSuSOZEPqsh2vWX9vdL+bPYHfF0
gr1+Jf+yiF+I9Cs4NJ9FbDoEkX+TKslHVq9OaYfGtZToTbUULILJyHbjVi+v1YZX
2FGExaZ2wKISn5kq4cEJ+X/6LYwhDhsZpfBKUpGpy6Eizpb9zynVZUgij0AcdnmH
q3j72aYfde+0BPi/t50nOXNU83VIbCqxkKwrNqVn/lksOQ+2YA9jgefTKPjjhUY0
T1dnKxcz55418fFGt1J6HnxnwD9GE51D5d9HvhUT/+RDUhaYAZ6ApUDsjXvwSChy
KVRqWgX99TeHYHWAb+wVeTItjRA6c4chEQT9SK5NHlIPHpq+cPSTNSlxmzj9UjWZ
QWKTL0mKyBUo9qKUWhaxrM5rIPYzUG2i2EYjOOUUTmOHaZIyPicVagWWEM2AJlvL
17gbN32b01dFl4cMitDdVL7iVDuisd45y+dQVFIWjXdgGibQeg3q1oVorF7zGYEL
hg1/PROmnV7gozryMqme1CinzZDPzVH4nA6sPNAZ1rvAgYMjXI7TQQWzzIA6yBTF
2Y5Ga54iDR7PV0pUSpN9ryiHvIONhvNs5SS1Z3rsOzJBUHGmzWtxRxQCvOvAApmK
g7Ruhs56uyuwDdS1noeT5aKXJrRir5aTeP4nRnTmUHRWQVbFaBZjZYZNygdiOs9K
1feODh7ugRbx+aT8NCuQyJSDZF+Ltlltoceyx/tr2cfhUWFbW7ETvr/u4uFWrYRu
9k1V4a3il6gL6+yvo59isOEeU0cHbVnKUUnhkQF7UUHFmDq+GVmDa5A70KDEysbi
J+xDZDZsOhppEhcjpGeUybaR1uEZI/yy0VbeVEoTiH+YL1CTw+4fSHfRJaMCtYTz
5ovrxYIPMZ7HnrYnivdibucpIqQLAGqUhn9RZtEZj+/COH4M6H/pJqjTODZBrQT6
LwTH//dq4RLqU8ZhLmgxteex1pDHDOqmc9lMfFhtfxgD4K4jHsxNy4LZGCH4ssci
yZh/wcIe588WuA8x6UaR9e/E0R3U++7tAZ18qX0U6Bx5FhmPHjyPwcfYnUdvmdHV
uxKxif7PRMDOI2lxDdKPQWHvUyKxyhNQN48MUMeDsCI/saTGraJHJ3so2bTPG9A3
CcIMfhWUEWaAqBUdZpSl7RaQStiCVPyEKvaCEiNyjfxNUHrWoKsRhvkvX8SeDcbV
P6/7YBxsIPZIf2VEoJEH0AOYJkt7cugE5k9N4/jBoCbA5v2/DRvOg0ttos0Ed/v1
mqcXfDSruiZAsKzStod1D2vjGUQHPSf9gL0EEE1ONNQIPdJOHSqqDYljl8PjNDX7
ECNW+Zt66BpOnLtQUxwztABCQacLBPJlV+CDnY98hCCR3SIjt4QmEoReB4o95a4w
Iq804H9InpEHlpxhx4gKYeBoPbpQ6qKherr2MpjYmMRta8g7IcntqWhsPMxwyvTA
qHUEPeIbe0YLFgaSGnGQ/un+/V1fBNOu3cu52Y6t22azfDdNQInNqMS1BRJ0z9Lu
j13ZQ7YJlvEBzU6buSDmb70f2nc/tIeGqP9Z9msU4ojF13DQREQhiWL+Ffax5zNn
tVroP2gN8VsjxerwvREFdh9ec8QOuRklRd5NtNiWRi+pmi515VOD5iM/uERi9YnE
LUqXjxuRYUGWGZbHE4zoHsCs+QjgKspFVKnigwo6j7x2P4K5lWhbxwKSLBEDZZDf
1LsZ5W8ICbz+a8X9G1DeAxPZ2mkXmdXLXn+oEXeODzoDhH3DGFQ8j1YLORogQv64
quSuv8XiRyUweHXTVT+nACIk0tJFKeuDUA7GDcDh9RV9FUbQ2KNQEkBquehjIeUv
1d63LR64joYk+FNKhdJGz6w1+ghGKxXndGPFfJT8FhpUMx6Af28rUAVxHQaZ0Dlh
JqIzoYlcWiV1ZB8YSf6wdoiIzyDoPsBY3s9ydNUVV9+syXgg9sfUYI7Im7qM6hIm
nZ510xjLmYtm44wF4aGENOD/eHTEevHFHGIxwsgIl4A1kj1OoN0siaQTSD2+uuuq
XVkbZah19Yur/lvwXfU+WCQvN1vCkh7BgJv0KO2zWkmcmT75YylT3pI++iWdYcBm
1QM2XERL9uc/ttD/fBSaJXUPq2vW9PgbqhU/Oysu297Q9OP11XaGLPFl6ptIqSmm
Bu836kqPrcehlfeJ+O+InwWQJg6RaqIt7md+eZ0lQJab7m/yrSiWvPGT6535LxoB
i6nVfY1qRiM02WTLHuWWvG2swhLEBqw2d8f0TpiMeKK4zv5ZT1FDHXoO0bERKG6j
rcnXft195V015MZwu/zlAnaA01CUdP7U5+smqxvSthZ0IfOXtU2vpJFOMKoSqHCa
UX6yuFgZf4kiEDAQLpsTg3uh6LcqX8EixBXwn403LlWVRBwJDjXNIierRyBoYzbs
hvyak2m2+AlZURaNZv2SIh8bKrycq4Bw/jfksmqWmHb7MMk5wbj5fsMVBsn+HOxI
0coi/LGmA2kbFjSbaup7/5fW4UaCAHopbokpWEMrXktpzRS/9iqM8LBq3TNFvYAO
LAekop66+qaZ1vK28FdP0H07mnmSgyyO4mOQw3RCGGVvRMGqR3Y3tOr1C6bGE7CW
pAmJbUn/J+NBDSVrqoTOT93Fxgl/GczgLBY6CjeF63cQoTfp9Ea23UG2nRJ+V5IT
yzA/96CaxmrvHZskoWTYUzE7Sy+Vt0KEu79AL2vw1JLI8/kK9shBjqJf2zGYPGIt
9RhTDwtznKWJmPn6YFlRWenw58u6yABvOJlhHB1awAydHK/faFBemdhFEqYbG48R
FXiC/D74xzsJ/iB97Y+cq4VvkbwgHM6OBFPl2rOh7jvmdeE2gHetNjomf192zNol
BJdCafYeP09n65l4YxTqdLz57SwwotyJlX+WFd/PL+pxe0OnTk5csiL1kTtJO3VO
o7U5HvPIKOxB3fyltq1tNzAaqZ6SUXpRW7hMVnK8SQpTbxqQYW3rXI6QL4kAL6aC
EbXIhcD82fF1mpONy9yQRLYsQSoyw59aRhtp2o26kjvLvKvXc/XHxr1yIUFagaFv
m9NIGnS3yWT4D+H/14nmrSeUAXtKVqESTuGefDXPTy4EFFEgZpfAHQHapLbupHIQ
6a3iZ84QIMFTgUhw7TiRyfZ1eGCm4h4nOXhN59xq10cGj/sqgWUfgWltQVajepPN
d6vCJLzN/mifojZiNtzZYJHfe1tA2QVomw7WJWVJ9Anlp6ed9Jkw0jLmOv2wV0Kb
nVQVPHWC9M7hAmCXQz/1QeWTYLdOBSTSCtPGnC1J/dCk58V597cxQ8y6TvXaG5HD
PXMq/i9GogivK04MUX/c8c+2OupXF65mDM5dj4/4WClQBFblje4eWRYahl4XUo/9
+NEOxBVh1a/y279m7gIoNtCPxj1vGaTydA1/oMtQ37FBeLHvrmFZukb8wBS3BBi7
TrLzIacAVQh0EP90FY8SqpVl0MZvyXGnMqQkAShX1BG9VEdgH0fN4T6OrRNjfdYh
6nIUlTDdsGFNwYTqntVDLNlUjjD8tT722IxI5MsISxWhuQkVMKbeMysH7eCJjBgr
PwecV6wMnZM89cH2uVj2+ZZOoRO7C19uqkIgEWsPPPJP6i4mPZ4h06m46f4idy5h
1VgghEB45BlrRzvuI942M3mNeKG6xQqURnwn2/wwmO0WFfqS2YAuUmemgc236b6q
R+C/Q2G8k9q7aw/jWd+z435weWbi6p2skN4c6pUS2vjSPTalbQ5aTOUXBZLnl86J
HStDKIAUhR/skgBgodh3WOcGoytf0Kw+f3ppFkMMS8S6RtW/p0N3wsICKoLUGuMo
Aq2kVz0IUTlFL8styUoQA2tdipQHJjcyBzsVq4VF3iK1rHe2zgseV4u29gH/0kC4
dwDlXJgMS5Jm5H8Cy+pRqRgderDPOcA/H6kYSp+PIexbFYcBHN/MqhNLa23bmQHf
j812FjQlWbL2e0ewYzj3QqTPJfZKlNlDb7c7jkXWXFylzNbc1NgmFiK7cRoSBXSt
jCb2EZxOH11aYSYMI7jEagqYbGBVAA2DSFumZH6onZIUlS0j0/GFC/UQP/9NtFb7
fFWsyspWChzF719FMDUTq4JASFowpPWuyK/wGh0TSq/WtkPu0UNVQP6RAzzG4yCD
GNiS5sx32My/rh0mPRiAzEijumowr+QCsUEhguadF5cAy8bKWhQwtYgoMIiOPtVo
poRsekm285nwJRcUMINWAO5HZPLuCTxNgSlZdycy6WKG0ecWNbL32BVds6BU35I2
fw2/ahTD7Nm+PeMw5+q7digmUutQFShlq0+6njt4dIGgFDcHIAQvoNUmVr6w3Amu
NrTczXtt2/o+ctMlXtwSne5tTGGrHjtJkcllU9uoMT4fEyZrtZXlQewgils/hmdi
DNl3KzqJNuh1M3Wbm0dnruX9XrE1cSHhjbM9ou0DvBuLvD0BpFkJ9A/R38rhM9ih
zyUH/5Girg/Mu8IXFHITuBnKzMcg9CPzN8NmcNlMQ4/8xwp9dQEk4bMIbFrHYTfB
vuW+RGWwBHAq8CUtRr+OdSGH1+pC1YMNNOejvJSBQt3c9BzIVcJeMjCB/y3KHEsD
Pm2Eabu7S6h2xvtf0GbrVt+kdQCiLInCSB6xa6H8e5I6upyKDxB8Ba04sjqg8MBz
CmfvFbaRUFHgPHYAqazkfnSS998SiO7SPZYdIrTWa3ykwnz9rvjEZqh6NS0fkPoT
CLvciiylYW29CASoWDss7TJZf12koINt6FSSywOicrJ1yFYZrY5rr1bgU9LNVGGq
FFd78gNPEMx0H1igOw6IvrSX9uyM+/SSunLn9HAeO8Tj0msnXx/+ONThd2m3xsZe
hWWd1ZEBojJ5UNbbAJuP4zFXYiFGJ903hjQbjKOzNrNZGfJRtRozYZzyMF5SrmKf
aoVN9mH3NPu65uuQpwIWGtJgoPsv+52aKQdKQj4P0oXnQ/A8Pqv60K3nq0FwTB1e
nhjn0ojhVq6+zF0PAXPFTkt/1ytDjB38NIpXJ/InaEY0V6HC4KOwFM/UAMAYj/O/
L/Pj7z5cSu9qSkwHNP53TYTHUG1Z2nJ+USiWYM2CRtXhg/3MWWZtPqEhAuxrGmkc
N+qY/imni+HQ+q7ont5uBZwMXdMCS7e1VGcS5VJH7OiPeLP25YjOP6Xw+m7mXlsK
h1MxA9KWQ8jWCASEcdPPKJm0BxFsGWoSMZu1bEvWAwE3M0MuV3kI+EQglRj9JTly
klCJRGFwUfrthW9mQ7KRXM5x86GuzcDQsCQuOi/Sp6dlpA8bI/AMcklfRsIXBw3c
3mYkLS94Wg3xCU8V8Z5WP5mp1wf+NVPmF+KLgOrrUi0hZSwiJTfccQF3lGzzNNlZ
tefhq3ehU/1ZNangHE/fIrG0tFMWuB4pqFaKtQ1mM3I4E/B8ToN4PKeuFZnts3cJ
KqmpUtIw2ZKk3mRXG8b2FhKjPNxs19mzKcleeBKLMY423zLpy7Upk3TUnFyM8nAQ
GSjCUOH7DW/diYBPeruo9t1lirdnJRjTQHqXeMv4ruRoIe8AHeJV9SZEgDCAmo1k
JYu0hMOIGpRZIV1z7tzNMvB91v0JxjvSkxcIEe2VsVOpRHsLHHGAE1xdFQNt8kTM
xxB7bRfghHRX4o936L8jQv8IbfZJARwggOXJBN23p1053qaNf1PN5rj51KvygXRC
ie0DRpSHvLfh4JTJpm/uNvfyvLc/m8AM+OJbhH2hUhHX0DdP9TZ+0s2VEr5E330l
kB3oJAB7uR96MRov/syp9pp0QsZ3zzPSGa6OjpomIQiAvxqxRvFnZ4NlQXEeiAT0
mKXd9uUGtFTa6bodSFajIJNGSo3DoM7Cty9ao9j8IuyBj8emngouITmvodlD2IHn
myfociOc3zdm1m7dwXCp+yU9URrqdX5cFvsjRQy1e9TfTIWEi68xzRRFcPzeregD
sZpucvE+RIN5GHeqDH4wHEdYsCm9bNlSmqC2Pd5FVZLTkPW8NqyuWZ9aIKOeFSRN
UcnOnwJcGM/gOXOxI4ysHTCYNP7Xgztp0NcGR4fekpwk+X9TK9ZZn4r7d5HpB4Fy
RGujGYMgIWLoowossIX36RTgYPgmTvTFS0JQwlCrWP2YkfzIeupx3sdv+cIBoUqI
8ZjRGScSTlCt8O0rHVnSAqAfZ8RVBWl2DJ9KXCAzMu4xNf77qXYgYLY6G1vRBwwa
HP06zi8XiT0LG+aYf8KjhLSJnfhVvtw/rpVw35hkVxhXlohCsSXJRJQAf0DsccjD
xYM76s3FqFCkA2bd/0SZco3VIsSFq6n903WtBuDu5JXci+1aGNplHkN1brPS1FDh
L8vV3jYhKMlCVhqRh3ZG3RQLkSD7IljD/B3F9eItuUsGK0mQJoizDgN31BRwJPeq
0j6ovqF1WwzxEu4l19zBxGMyJWUyKBF7P43FHoHsbQPhhhBNEU7oz1bG5NWBT626
LE6zgvQMtgXnmYoQcxvN2gGW+Ysm4ljfzaMNt8rPNcrFdwUTXCCsnyduY/E8DGTn
4XC2hYGOSgGQJ2LfrDIEoMfarNhTYI7fc3C1XZR1tBMqUBszpm6htcP4v5RS2fwE
cP0PJDXXiwyehWoTNTQI49NpgZWSjAknxXSOaA6JDIAwKYNWJr+CawtuX/l1/eHs
KVgQVMrbl39Bk08YPNJuIuO1KdnkgWlW+aW7eWnrdfIm5iAIm6aaCJ6q0yt+Hdgu
pkfEkekRd4FNFlHrMLIlSMSWkjveA7Au7SSvfLuKPBmKFmDEQaWzanduxzfs8y+N
hvXpZ4BamMqF7/uX4AyXWmI9XnVSTS5cXl3CWlyYHQ649OY0qq/1qOXuxUTNOW4l
88YLYhcDh0QOFFL7CMq0Olpu5dz4n/liBrlgjo8xAl2XERts0cHK7pJn0SpHyKFk
mqe6ALUE0VgkZh9yPRFNtpeitPeviWAZUr/ApihPEcrj62VqIVkbWCMzm3nOSYRR
WWUTvjAxDkt6sC+ENqCK00pXDiPcrod9XnRvj2jlZ975J+yaA4jOXqT9FUPEiQsX
rXJnNbZzQlv14DIWuQeKlkTyLkTPkw2G+9LNSnDAnPx7A0yH0XIf2xgFrzrLMXkn
p8NZG5/z3gSm7zK1P0JD2/m0pNesJpBCSQi5AKqO+w3J3o0Oml4HokmavKtxHpHC
gYhmv+0IsoI9hCny2hf9PT5cGDWGSQ5rtbYjt9Pjefa0m8TNCwPBjGrdWxyXGMJr
WONLv4lqzlwFEzOHoGnSwNrnVQCf8Kt/7C2zn0sXDC1UJh1DvZLjsmkLNwcNnF42
vY9mnONpbvjgkc/0aW54CPZSuxBLpK2wVr2/BtrbBFU3rpNomEiTu5PK5qElA6pS
R5Oskkaumzwcvs40YTzPT4eLI3P38MCZtgOjeZZPNJGQHwWEl9SPnszz08AeRMrH
Ru3dI+xCuTRJ2FQYLuN2Q1Bv+7N3s79kqDWMj5YVFPZ2O+7/cxVP1SbzKDlHorrb
Rf06byYlFvL6PAAvM6X9IGgYlh4feHG7smJ+hTSbWXGvXqZQv4nWmNEGRfNJ3R+c
nvAkhHhQK7/pV2dMmm1Vy+iKlmiZOeeRaxVyh5xGDw/rn7qdgQUrUTWY7hj4EfYK
C12UHZ96TEspdb4jrzETGPnfNz7jlaAOYKhdhJVZvnVGNCzNNugD/kXvYsrMxKUa
MSrBJIrXvJsnYM/ruzHXzWyEhlqPCM7HRDN0UQSVW3NB0nJKUIG8dI7gDe98Boyr
HQQjz6for13V1KeBJLchpyG5JheiODMnPl673JhhQVUtzHsnyeqiDlu2+CzowdX6
CwD0N0IyV8+ByUSMQ9V0IS7W6BCnH/AADrSAvPs+bvHh5cGmot3uOZz7lsNda2ct
e6MK1atBIFFdLYH93dfwL0Er8BlKFVzKJyDBXj+oHTvGpqcIJ2yjqpu+MYn86F3A
zp9PzcLhYSlJW9Sa7rf5d+dYZE7YBXlcrg/o3N4apwwsfRMBfBpUNm+N99cF3ROW
VKxNt+gd5x2AcUDsQplsuMkriqNXvDWswd8drXrrpnSF4rlCkbDiFP8On/QTpTC0
O/1X/i+DoIZbiKQ9hIa1XGwUUfWRmL8z5PBEVB4UFvWd4VAaF+M27/9aREuXpZiy
b2M3HFCRUnI/MYvzirLmVV0978pTZsgh30N6pxJyonOOzQuObGYz3mJ20lOc1pla
7qgwaKo/VUna7d9aSoieYjhfg9zji8Mvq8kEtalez3Sa0AgqKtvCOK6tdPvsDd3S
LqDtod04TV5ZbuQOgbsv/zZuXwSwNHJYG+ApU7eRvFvm2zdpWB5uDNk+5vqnsxVF
6OsxnRSP8xUdd0i9cpvER4YViR4DwpsNYSpXtyJ/7JOG5q9ppTq0smx5a3ian9n4
JkMqqT9Yz0mvwXJIVNvAEuXmye+Mc+bsIFYMtz02vuq/sfV/QMbN4X5klXHW8X3E
AS/8QR8WZTjYwnOgD4k2i7IZiNSu4jyK/yHDjcvzKjw+MF1ODjPe7NfQb0x/DjNV
1Qqt0yeOFkQfZOcwwmePgtzBB8sJWi5FKTq4eFpO84BJkqxcAq4eA+dW97bFlrvz
XD0yYYQVxQgb5C7Uxlx3ae1kwFZGJoHhf8gu/FsaMH1zUQ1sRu6lQnTN1mXsjfcG
Mfl566uRDBq7SNUMgATPEN2D/3pYx1T3X+Rqwa/JC54KIu3JNZFjdxbcCX/NoHkD
uYWsadub+qoYcKn6urXJjbq3U9ISyPu8ZMLoismHvQcWqu1o0rw+S4mXlQoercG4
KY7gPlo0BkRY3QCS+07ggjQAnEtcdBa1MLuAIR00JDOkr8iq07PjLZl47fd7dFRO
64kzZvmojjfF/8cFI0e+1JT/LkJjGXGpqnpMfwMJFCuilwOaKR3lbJaZTVnP5TLw
oGEkTJLQgiY0Xz11CimoC4iUxDoOt/ioXWGdtabF5CddVvLGMmiQ6ohCT38OH4dm
6sR9h8RSK9gLIxxJ1O5HPHEntMSSsbN9IGYRBKTZKXN7ZIx8i5DGnGbngmzd3aNn
5qxExwtFMD7aSmVbzOmFd8k2rGvcucGMBBFNCKWp2Q/9jAysj+bGQLOQG+jhPwqK
p0GV+w6sj5fVGeRrhirGhTvu7UrWO3clQvJ/1hDqRJAmLN79nFb5IQvVBvdRj+5+
9OT7UqQsGJzPGIUGd29CwDQvF+466YorVMoCdZBPxIpR3W9moskxPjDa6DtzD+on
tCYZFKq2vCoJ5n3lkW7JmbeseJbezcSt2z9N7ALEzYyoliezkSvcu7naVxl0b9TB
ARWgDwcG042djG2qLIx/wXXAzqpCMwuBZGnOVHwDuiNtzXO915V09kqN3UhQFujQ
Nd5lbGuozRPVqVwZFJcBTSaP208fH4J3jUGfZ5Bn9zcwili4vEpAtyq8pLXXN/4c
QjCopoRB2mVq6erARkrlBf7++a15QMYQhMP5z2ktuHVkjPDusL8cuwfWD6uvTxLL
UrG38W1SO5PQEJ+82Pu3l48YfmkTjzha8ckvHfI3Ae8vlNrWHOLtLbQJLUqBG3zk
sBfmzdL4d0qfyQ5yeega+qqLW6vsYpb9BqtJS1rsv621+a3zc9zMGc78P1c96N3b
1Rb7rqxarYvxFJoOI8tRn3DswHglUQXtH/4LG9tjNdLRT9E/GnMc5fwy62OA0gTp
qgZg85lkgDCf2vfF6x6+77hlHd3x/NOvrLOFcd16TCiRz5sM7sdhEylCXSO9BtJW
CNz9F9GXYGYXDOdxdt5MNXnXwjKGCe9QF1Cs7+5OGknykGkKxHvdBn2MJ5Z+o5eK
6KoHveoiQ0Zusa7SmDd04CDIsQiVvOgHH2jMTLngHzD5pI4lhzHNXKfWANSC01CW
6LQAHBUSU8acEvh51pFCl/YDSjAlzHkyI6dce+yunaxn6GF3Vo5+Vm0YjF/DJRhh
wKtz7hk4zZde85HfkAsdQv5Nwn/lV7U6H3k+gVvR3UvzmgfJD/ZW264TNCqMlhhL
/Pbi/uONbqoXIFk8jqis2EERlXudtvBwx8Mg7EQez3zQ1l21GaiZkIJtZ6L6C0Bi
iyx29qChUMgyw8WRV4xcjVPTXMFfBMNibL9nJkg96jraY9hybrjfGNwS6p6WJVs4
E3TpB7r8vArqJ/lqaX7IRNM73Um99P1IDVP4vlRK9cb0t9FlgzjDTUh6OtzHT4/0
36mgY1gVJ5SAjgLMaEulbWzjApgUJKTdy8PZvbqUw6d2lItdWEyiJf/5ZyLS75ct
8TEOPYgSsg1J0R/KLvVIof6GOdZvUOqVAdPQPW07u9HTc5qe7w6kb7DiYxqJ1DBs
XFNLio01nEeQ4V53HCMA+jgg1z+S38SAbzzlak2XLoNNpS3VtoGBQ8LABakoi7Or
cPez5D0eLvPsm3+BmrkKziYn4T0Sa7NQ7VUN1a+mA0QtcGPH8wzjID1qz2Q4vyVr
zigFd4rOgbUqTli32IcWlXiKIGnv69ZwH+s1umThtabjEyjpihc4OKuJqSA3gNCx
EDAF1IiN2xaps1SH07tpi4jCud+HzKm8KF64YfRpUUMND945DEQINohGLgT6TJ7d
D1DIEyYWtZVrcf/vysvkrf5fT0Ym0J2ocY7z37FnlMNznRxdbsLld6KfOhXWRlgQ
/39YVXPtw7sRWhluiumUmVxqjWRebxHzdRKP9PV4f1pH4rNunVKrEus2tPnHf3Or
JKpgIGUzlD0SvKMcuorsy3/faP+py53r2x47feB+A6aM4iYD0Y+h9IePFCqe+NmU
UuZC+JlPpILjkTommzbf4ZitQ/zets15RyY/gg+XINpZJUEdz5wBUkyYy0qdsrkw
Xnf2d1VfqQHlpNQxAhSSUHLpNtMIuUK0XoXBqozg1v5iAxxvaOEuDDEKRtm9BsR8
MJkUxxDjRock8E+aKlqMZgFb/2FrBkdiZR8b5mY/CLV+vwhG3GzERJIpbcwMF4V+
BEmTSlFcFOZ/RugLLQ0odkPezI3ft/3u9YE+tkdjgWhZt8e+qA19FdpECThzt1B1
SuCpyGm/U7w48tWo5FwwekJybUrgRfHkFpEwZQjwP984GhqsZR/eXK8mX5H7wAjn
3S7MLwrrTGmnyQkfWPfLZbeSzpW3+OVK5mSqV5cExVDVmGk3koZ2r/7PGGLGFnwD
F7/4uvPf+FTv69D3urlHGYP8B0bvylfjF3wPWrMhuFcPB1MhoDUmY3hSwezEYn7S
OCPXXOXg+kGgp0l2C6vFp0fUmemszpG55Ym5Q6POmENravLwvrPBC7HlH6s5/WM9
TJn4q5wKaC7KEfzNaiL3RnJg/3afMtmqxWlOHobJZGkVEs+UHSj/RV7Qwwsb+HPg
SxvDP6JqUTfOOXw8U2wfVPemDf1vKR+SgZOAhO1BE3kCj/e3rzBQT+YuvMhDyXmj
NUT1Ce+63VgfY/PiFgGcSN/g2uVj413bYoVgf0S2LKEqlmc2YiVyul/k4GpdCHcX
DtAMLOgdYCnVeT5YRxJRKRTwktzk2nHTHo+wh3edNiQNE+K4VBpFR/TBGRnf8K01
TwCbtAQad0Vcq0bSvDHiVH/8uqmuM1bJ6LCrYcgWl/nFCjyLRs/W1yQ6BPZAWAaa
+hXpHklPxFpGHuv5YZRI6Xknj02eMmf7m7BYjic6zMMoIfg9+bt3Ci4V6QFyH3SF
S7n0E6ZlkfLVunX2K75w+bDq2Cf6MkpT4h8/NZj0sYhw4O1Kr02Of06pqek/jWYu
N2JZzlZuG/P0qNPi+NCP1RzUAxj8u4MUQVqXb/9gy/6BqmRy78H0XwGaKNekbMCX
j605iL2dPOids+7ko6QGPf5eEHtuKfa889gep1oXTYuOdvJEXV6p7UjmSNe0/qcm
CkuFHxa2uIQijb+6p2mXJhKISBoXH51W/re9087Lu3ndQya/uqKMT16kY9yO1/24
d/w+iMoUudjn9zC230hNf5nRGJLTTju9zYv1dRfql+1C1tszrzWl/MBGQF02lMJ5
JM6jiB838kqrdh60v5/aaFXDELfUUj3UjWMgDlYHJAw6cje2pv+HqE6s+d9tERWZ
4RmVgi41zCnu/a/ChkHFBlmK42WVqw9zaQe53FJwlfN59BavgvW+H9udoRmd9zo9
kpSF3zEX69SxoXEH4d3Er3oM0ZiLVcXRmJTIE22sVTP2U3Ttk5KbN88kre2Mr0G9
PuroG8s/dvf4svW6njGNK+VhKnhubt+8WuA4a8mHXQ8sVGufkbzdcJU33w4UfzOJ
2zEag+VdoEJoBrQbB+YTwuIwOBEvIlPiEQTwxYVrjZbIMcqTKvvIOUOj84rQWBa1
OiJJ3LxdbkaEWbtfaBtnqF1IsGqlOfugKpUjb4gZVyhF0FhjmFrBjqB9XbxPDlev
W7Gb5SKmeeG8FCq6CKb+033tkQwxaRyXoD+qcfhg3Hlif224BRt8sBuZDwnSBfa2
WSYBC/PqfMAH+PNb4Q+U2MICYBCSGnDvVFkGiEYIGxHXmgGzEY1ilO4MAQgdyU/C
XQr/YGaFU+pVcs+dcAED9rzUHFivnj9ixZhj4o7nSvTq4RV+fhEH3z5b8rqCMqht
qs82sz8w1/IXaaE+uh/LLntIugNUcdemMeIRj+NuelBA2Fa5pcqoUknQHZIxH7bm
Vz9eFmahBdPkoZsjIC2dZjNz4RFuKt8+xg3AwGxkT2i59IrfQCUxNuXzLfpWzkib
3HppEwPLE89khyKwbq5Mdn87L6bC3Pyv1EBDWMheQPzOBOfOG96MoUF7leQueB6+
Y1qWfv8wirnec5MZfOYew7jc+/zoZ4FdH8/GuEQATL85JtITeebZKc0Aprvx26dq
F/h5ViRrcAPiIkFKY8Q4bMXV1k5nShcb3LNLU6YZzw60L9rX77hEOnuYMhRuvoFt
aDiuxx/pSrPD23ePR01l14XLoB/8W3c/yTrx2QjaIwrrCeUwwEVCmmnUPuxVpyE2
e8Q75CO2hJ9sJCZxgcFUWrOrvfpqpOooNyAKm5L2f214wwIF3Yijh4FEA7gMePwI
CN4aBQuvgGPLdd8a92dN0B8hZrDjdswADkvVERZSX0gEJMkBJOSIVhgh6bUYCR/t
qgoHyEO+DPH1VYF5QoTlePvKbXRowMMCbqeDfhyQ/SbvMx1QWSq1vIquFqUS8nao
sdXdblMxPsGNIHaPOO8XmxJZVAfRqvX6hsbAPrJP7FZ+nwiVQu2jhlXWSrXoPZ/R
/DlsizKDAtF4TU0SDGk3vmMPHi5oZvBu+MQYCrhfQPHO7U+rUUr23XLF9+QcNqIf
dOpH2XCZrgrWsVSvuUkSQGWnN/tPSvxBdyhZH4LzOzT3fQK83U4QjtK0Df0ZY/Lb
7Bo+PM6Fb99QXMrXHHMp0i9TBQasarwzHvnwZFE3zxuMY+v72YE6HYvCrSzHBDBp
J544Ua/PtahSqabCG7edjbnIzbC2MiTK3BBZ6nsDAHMXKAIChc2KXV8KBiLQcSCT
YxZkSa8v2PirW8dfP9hCpqJ9dWLZ7K9tD7I8N3XPrQu0mbYKB2j2QxBHEPKwZZCC
xWO9RHgKGXSwke7ucwUPDhcIAdlzfiLD1owUzxMPKuduQyBaqEN1niszgRo1I+4g
CbsqXNk29ZfC4iZqNwEa6b5DiPhR4f8oWPWuCAtfdCe1E+9y7qYV7KFpyccaAb+P
pGqluBgIEOuEa9kH+yWLnJon/30x5c72f+Tf3pS3VsvT3jAPJbyQ+rFWKX5K+Tic
kGa8yhgDcNKMGfRoywPr/Q2aCXT6LCqnt31Dv3QkZqdtEBGgEkGzdPtgbHoG3Rio
GKhMqj9GYub28ZjH4Sx3t8ptf5mbEvBnjw3CDaixjExLCEs5MCoKRZ+WASTpGz8k
0igCN6rDv09VuLd9nbX7WPVzZt3erqSJThNjJzV0HL8cMmxwbWqnM1mR+BAIe81m
M6R75J8sLGHnHBBCp0YvqH2xGm9QTtak80WwWzaGCcrhxYoByaIyDGqenhG44/z/
42zt7aMZY8CtkAexADukuyVVZiJbwBPZ4TRfWbArMFUBFqBOkFdmPftNZe5tFqOV
V+ALh2F+cjb3FDGJ9o29cfW61AGHipEuVS/J+QbaHi3I7Pp0z7sRwSlLecChWLYz
Q+eG4nQNRgqFrMZuhWwsTQQSaFwfvxp/W/03XUxAa/IXRmatDgpwUDdIhyo8vv4o
ifKKjoqUGdo9QAI/j5bSqlqIbI+79vHwASNsxifW/uSNIDK9MuX+KjTvCprDl4fl
vGYu+43Fq7PPxYOVzL3s0aAou2rxt17Y7zhpzVcOvju0rCxUyI30b/d/k81WhSWJ
uvFt8HOnl4nMIRKmCmddw+cpoKXkZ1zkIE4XbBb86ocNznOTZE4CHqid09QFfq1W
qkwYaKx3JcPS6Xr268rrmajix4wWYs4iJkkJdATasbGylSUhPL7umpkrFm6LcUxO
Bp6SSo/MamtsZk//noaoKt12o8ZKcNNRHt4yikMTF7uj/Q7nUAecV3BU3uS9OWsV
bxEApJK2SRWh5YpsYSzkhRyBvhBrZWDOuRm5qelq52eptP/JtFnPkVXOpQm1Z+5J
VIUso3iXr4kAlOfdRg6ohoGGSRUdgOHPsdEmJWhPFbQOnnDFn5PN05qns4yhuzXZ
w+PuDmkofYNqYIluN3YxhWpyMdyJIehM7Al8i+klX+7VPLSC8kixraby+ICY/b6o
mHRA5Ak6NSqGw2JvJGq0tmYul/3dFNlZioKb73RmN1bKzrmcbbfLIAdvArTll9zU
w8C7teVVQkZ7zgP6SVS9WP1KM5K+PfgahiJZYQA8v2rGG/ovPvn7kPsSv7qMUghJ
v7LJnzMhPvnmV1I3w3N2iZEs8lVUVMI7gulutaqboig6qnxcjJQRqtl5x9eC83om
cOjQj/okvuJsuN8chg7K7tGXucukBPXYwm+9+xifhmwCecer6lW+geqJk2YxAcau
Ki8qCR/u05PYXr2RD+nsEFxM34GwBbjrdaq1YEFUXh90yyca2X92B2wvK3z0KcNF
iTjozEnaGB1DdYR0ZY3n8lhnC68vMFUCjFiJn6rmPOPZyxtotG2Q6R01JPnTmgEm
FXoleM6xDZ4JwR54u/hGJbaPqaUsgVYiBAN23889neAs+JUodEXEFSHpkHDcYPL3
YXNdV3bYy5x15raBWGERduYIOR1amKbERgluGPtW6jTxAXow8I/c3gg4TLd7FJ/B
mAxLAZPOGbVwNtr4dYxjzELetavIell4EUl9W2wF97EAaDhP5gJBSMqTgHjakf5s
EQcYa2/Jyc2XY5Qvx4T43HuLcwTUgNvH+1WddIw2cHdMaoxrUQbHyPDTUp7pYpN5
foD2l1l4LkJWS9iky/aOh4/EvXLfaAC3w4zwIPe92b4wUN/Al8fzucqChGzlktSH
5iEyOr3W/FAiEy3uXre/zMEolzenkt6na8hRdgYd7DwlBHJNUQ6qRAZbhkaRgLtT
qbhQ+YP8dptNTyU/2TWRuSz2zq1lhAszu+urzweEAfZZBeirUayYNrwk0/Mx61CQ
MSHPd7j6eyG8BDFpCN8PiayxURGiJjlYSOyJkcjs608/RCs5kp7MWPmCmtTG76K4
J/jisqLHqhV/mc4+53tYwz431HMDXxkA4fsZsDa1iXTxx97mgsQFJG4otyQEiDtA
GW/qX3WeNWpk7diD/rsnOqY/8YeJ/amW4NnY89c3Vbgs5PmjYFmdA0uRO77yaYwT
13sn22tIIL0InHIX00jv137UPPh46OIScuqzJdCbN+y2yd2WDv0K8QJCVNiwoVfO
eTwQ+MUD3WSjF2V+P1cSxTrlG3oPOxiRUVaWN4gjhwnhg/SQG02stKMWcFF/01VJ
M3kG8S/huElDKmJF5pmWGX3zpHI2tDlzk1tcIjQXV80aPAhpVtjpjH9vNMTw+eHd
SsBAXi1FhvFw/BP/bSoPmYc2rFoTMaAbludC2OMiw3NuLGVUJdXwvCltkURtPq3k
oF/kL0wTyRfaAzpTyDjgdL8BofZ7B30InV8Eh0tIqMh+tumogDzxl98yzDeVZAoH
s9L+F0RslZy3jUiKSwV8Wa/dZEcZT9ynmc2BAjDgExZMgJio0OkV4J0s0nQF2y4E
chRE9CXMeZt8upHsafWLpMP8299duSaOra0239wy9Sns741XXGC+JUxht07CCShw
tFvAAeCRR/Z91JQQshcqW5E/bXvudqg+sxFTbfFSF1ARhwBtFl93W3TpBh+A5Wgs
eP2P7TV7yovS63nep+FuHNJ/fPprPFA9iJMbpPiTKdbY4ux/aZ51hm5y74IVFoa5
s6ZSSUNF0L9h2NMjZitgPzk5I5ih9M2rkA37XlwrOVefWPxx/oukwKJpMTkKb0fy
1GBJkxjQG5wP9SNJArmozixPXs78HSDGt7mrsp0TKS9chn/D/iMa9SSRMqGbi23Z
SH9S8YT8P0N9IrR5H+l/r7go1z/CQZE3RvkKNyTy9Rf6x7RwucWVtnKrLGQMTu4Q
g3zr6SjrdUwMS3Lf2Hf9tBeeZmZ6ohVQTt+RTBzGcxdRxNmPh4qcgG9YVL43T9J9
kI4REAS0BXHxpVQ3orHmQOzg1pqoT9UHClg3ohBmEQH98aYfhsl2Wz3yATKjXFpU
tyfdNzw5uIyVIlRxA4kRB/gdZHUuOkpsWyL9keGZzdZ+6NYVkSvCtAFZxAKhM9AP
+UmrFxZSIUys+mM5qw23rsbVj3afh+XrNc08GNIiEipi83i/9uSg/2xUWrlajtrV
ZkQI+GC7WE9f7TJ3kxs6dHygA2MO1O/jj4Qpiaq4Bzu3EJrnP+Ay64PHWauyvMhR
r8tkV596/hsoTz50kRYzLhXzQwrO64LLUpbk7wNemB5xbpNd/hslOYH489ZogcQj
yZFHzksknprsXYxwdCKoBA7uzCJ3F8P2+ytqTAgcNzrKmWyUrWYlw4p9Bh9E3jQL
c968d5+bZ97/kc0JFS9f+SMAhj8l4IEQPu5hA+x6PESynBSwn+IC1g6+Te0ZHQJt
d6CdDqQUjZTZqKcvswIgyTra3HSl5ufwQ0aRhFXgPzKXRpjoudCWYqvJR20v8Anr
4aezXk9BYaun6ijKEp53SnkmcYCvBGDyRyF55zvSEBw7fsfp1uD3czYWVOs26sfP
VlhKnQOKXFEVZffZqBSgQ365aSuKw+kRIcM40wcGcyr9fcklLcV9azFij81XAfLu
Xuxk01w9XuzXJp6rv9qbJA6xm1/0mAKGKm2/4MxwRVRRTY+R6XDT6inHJm0FNMEx
EIqtTBki8hZDipfxL/IMK9azOJ+aaE78KdNYl1M5Tot+iDoZ/AzlqcfCFKioPXU3
ckpjTgmJQbyxiMrxOIkdLwIiDDrzZ0K6EUot+PaunNbtYIsVvFXDbPFMgb8rdBc2
M3nIlBvVjsJsuT4o7Kqz9D9sCdkV0LrxhKyODMDBijIocX/W+ka4482iJKz69vXq
2vIecuaX/8XxZz9E2IO6qsl0YofpUm4s36+XndhiOe66j+K/HsOS/lYfgixBTwaN
4jHOaXpRL6LcEcm8lySUnKw4HwGXloFiD4Re76XGMJCcRLPQ1A0GzOKytCL9KTPT
/A79iwIU/nQ1bYbXyomkv+WH83zhKgFEAmz9FOzonZh9iQYsnYC37d4wf0eUMjIg
YoB8G01oC6hj3cbrXO6TNjiKVhtfVLGn1B80+RIKmTvoEyEXhB7lLfYAsAv7cJM1
AUdryL7xX/WKNcQcMuQ7fZTsCLIFurIj4mtXiDDCkKE5fd++jilKxshK8aQa00x6
RBUVp9GSwVoapB2SYlQfgrx/eZRNswmIMuMvjoTeL6YFJDhGX6HUzV7EYrbCrJEB
ou9/Di/S1fwTkA09yxDTYYedXKQfKhecTKGRKelWDOv5H5D7zlGJv9ouB+OwoZmo
6Ppg/JU/rZA5j173OQ/5dq/LBGRt5TyAt67V/TY5ntQiMMMGRbSUk2iuLv8ZTIpr
r3EjwBNE7ZVda6uppS0FP1yUWjM5EeEuL4m/uu9JyH8NH56Sv7DA8qQfVVrnkdSe
AC4LmmyEw5urIykrTXyYvc2zhCLxZBhK/Rr6LFju5PZgxdKriXf8E9CdA5x/Dfrk
bvA99HR/7J/7QuSBH2sQJWnsrGhxQf8tcks3fI3Vz+OFPkrMYIIl/O1JsrfkQufv
uPTAQBFNNyRnD9yNyiXrg8FOKeNdk+KwafpouxDnYl6OnwKJBRhWKml/jMq10OwV
Z/ut84lT4wBhtU9WCWHZhi8dOikg0byZ+H0UJvEmKpOf/JCOoBFuzW3m+YMeO6BY
s8LWk4X5zc3B02Vnv1aGQXuutD3ggRhvlGhJ1kJW6E4FTVJYnWm5emR//mWrr/sY
vkKF8bzFFjwmIz2xCBneMab65bkBU6Af6EbhpzMycl8VSrKcHCSssrff3MXTfru9
r1QRGhft/tTh7m2/628H0b83DWzfZl4isczyKAWbmoUiyunhJA/3/DUYADcoLBwh
qmPAh9Q8KPkYAvEMuxq5Est+Q7LZ0Cy2oVI+N473gUlexrE9BJysHqW07RYjXP/w
Q+C4bJXX4s2vV4nKwaJTOESquJDcm8dIT6bsfJJ+pl0XH0bawBPjKY/5deCPrudx
UEYs8LiRMoy4LgPxVmgtJQgO8ytY3MRUfdMiGjjWOC1Pm29bvRP2vXfsH6pdT5Tm
Pz4Sn5h5M+k9QvDwPgVfokVV9JwZ7/YXel9L/dJmTn02pinvq0568oO/l7iqRzs0
stwl72R66Idq2D4LCY+4kqJjBYExxxv3UueU3F9A+UvVUlEPCTDiyYDeSwMiy4mk
/aqnK8Znwk/gnpAZLdvaKbHInQSa9vWiFvs1YbCHDV4JXtAOZWc3RfIJ9/7lhCGX
81QWJAINHqSqT+/afgtT80njoWlixvWU15uhRI15Ssetv6Pz6Mk4erl7wpSVcUvJ
RzAxucVJZi1hcC0ufAQJjaCLNleOYAz9C+ycFazmwI7zvCV3r0q+OY5+TOhaMSmn
UF6/A956C9RqB3j3QORTn7vVWvgnb50/Qo7VxSfwXoZbzcOCuDShlgf/BX2v4jvH
ZSdXbZlrS3BaweXEUMy3s9isa0X8/xNH9/BynE/dRpnm7kb9BnN6LzFBNA5Xv3ok
CwO6cE7jw+fGv0NQgXeTyCPvJ6jTJKC5Hxj5U1qOawb/hhKwVAkCSIz4CLD0e+jC
PbWT+76gNWaF4e19N1DH4f+ZaJgsAeZJafedfONw7DUeSvLUotOKb0tScGMFGkec
Ja90o0RlvU2tn4S2F7/+TrqBi3ksDIxwd7qTsGI1x04dMkFjnhl57dZs7sT9GONY
ny2au8Pr1chDDn2O4/HaNRTnO5iS8qiy0P4vgWLI8khaRrkYn+YPekdn+AydYYf4
yygNKwbkOK26VKG1ao7vZhdO8mzZNDRMW3lECAb6wIB1IJJ0KXoDCisXwV77Fjdi
lyLSa3xfqadtIGUUwZ/bIcvmk3MM1oQWzupvOZa6HnrhIexvrnHwyY3mjRVxUxeH
Y6LVRONrnJ64SWqgMpp1vKvql0qkBma14uU90JfWlKbakef/cHbdqfVSvVecpXJw
Qxyks4WieoVdfmQ6mk4W1NjJcG2f/77r2TZQUcZDIHI2C3nnsxB2Wf+tlQT4j+o5
3BHWTA3O/DXlVK7XEj7O4n7Jldy9roWwwf1u3RD91biT3EctCxOOLoZwHqr6Czqu
dYCgomtqsUVrwvHq3WzWEE1vWZ0r/MO5eC6KlGGQHz4J4T4HpoTKZUduRlbI9pnI
5GvGlgQgw/dKj2uG/+N+i3jamr78bcoBE47wHVsAnbwWT05pPlgc76L+rhPlNFxY
tBLxwiucf7z47FaB0UHQOyNLHXzb+absAGvJMiyJz0utK17Y3TjXs6OpL6lUwaxy
W9q71MJT6iCzTlWWLMWA+JG8vUjdtYxGJojySxTjOJxn1eX6lRQ0gwawzFpdH2TB
2klBkMoNvceqZaohNQ+LVYQSzBeXbT+5ftqTyGrk9q80uAOrSkGfXl9yKEko88qT
/HAF68bu+4FpSsJZg6sQNJvuqWHj04rgVVvT8v9Z8BSGeeSOPBv8OCDJ2cA6AtTt
N+7JdI42Gf9Ifk8gaJH6Q9v2tc6KJG+osjJym15GfBnrCTjseCQir3uZUFYDr/V5
X2aiJ3vF2CR/YOC13EF4H5fjXWW/A7pFb7lldmPSzXmn4klyRDWO44s97fap71lV
FBp825dVgT8QEMKLAOQHiUe2o3349WfUqc5HU8OoJGsBEzvo3wkBy/Pw1A69bIXP
kBXjKHVlyWONhbD0deVOeZqubHM9yG7YuGQEknQgKoa2s4eAqMdq3xUB6GFzh61B
PKIzD7E0/LEnhMhEaEpDnE2+aEz8bsbTfTFe07nBR7kTqJomNkgklRbqwf4w+RsT
13O5AgV2B144GEUenEWZ3l+D6q1KwHToJn0FDe/rKbYAousd6FKuEInXdk6PxT9p
2+US2eS9hrXRNMG30RAk9Sn02qSZqGVjiy9RI/VsTAgdUawn9KhlRPET+/OMwiQ1
QMrKIvqUIWGLVjtrhninRpGe6lCHTcsWXjQdLsQQ/fa1DP02NLLexDomvGLYDZqR
rf7xhiSKN7b/8RWkFjp0k4XmqJPCtrgykjZpdyUbTwe+DwGjBDkjszwnKX0Z2Zbo
LBh/evVcuMWvxzrXYTOSKS1tX/PRlaFQ1KryIas3R6zi0uhMZgzhD+/dnQKc7v8J
28JsuyRjxU2JNpTGL2fBDtSVY164X5no/XTHod9X5ByvPB8YD/kra1FhssEShbda
PN4aVmKPvZL95OSs9otDqPzg2pmb3jR0BbBNEvf09mgD0UoO2U4jzVMWdZXJxNEh
e+kDhDLn7ObRXuc8EW2JWN/P6hxc1vtxF1Qz9igSOj4kkqFKnFernIIY4dzrTYiZ
ffpbP01ryBYD2FF7qeJoIcfhRN8fT6xZdqc+NHDJA006Axtkom9IGGJgfxGMZg//
HwQt+p+iyhHilxp74PToo0CuJaCJLbgo8ZeuGDC+4m4jinBD+H/1z45N2THhhCle
D8rFiQ3lzVaJZvtyXPIq67fVgu+OgGB39xdCym/WXNyvf6ntZKbBlMOqaZ6rIY4W
xPnRu5lipIimQUpf4kvpCCe7Sk4utwos52t7ekS7l1y0wMYEXQFbXM8QQ3X7FVk6
rpVnDzmnhOBDt6m4qLUBKnY7VzXbMlC7LmoYxDeY5TaPxJa6KCP+CFZZ2r+4dGM8
Mm5uAA/gGxVXksTkvMdjlczL5qk+aBl4XnY3WUyBPhyMbF4XL8IGuU52uuLAzfhD
mPKMemb+E5SBpCNE0I+9phDFC9CQwCiqHxOjZhNzeRGx8aOwqmL1qYgtCrsWMOiX
wEObBb3c/vN+5qRItToalf+czlNICgcKNkkFBD1qkmja6n5Uk3AJ14MPRyvxhhPn
RRd/lY9CfdvtY8/Ho5GWnS9kwG/kYqNSrVLpRtn4RCPBrjrttFFDYZBUC9YXis/z
jCIf2YuE89oXHGF5LFn1UhHbFm591AkBCwFINZhHVreptP1lm8L+WY7T9MM73b/7
4d3VnRC/LojJqdZunkcpJ8y/kTBLeMu+46hoU6oXbH0NiKUbG9l6AlD58UhUVfrQ
+12dAFwBWK4rIh7ZZZSUkLHbU8hkXS9x7RXz2rb6oTradWuScmStGN/IRJkuUGr1
gPXLwjz3uRHE/L3uXaJWvJJcde2OMvCYCDGcQSpkefm9vVXEYVZkNIx3U/mbDvif
JuI7e51wBfLmfVYBnHwHfTdSqWA/v2n/OeqUd6LUXY4IDv3aAXcex54IIqgcNABQ
Q92MQ8ohpRkH+5H36EBRkiI0HKj1cxnV7rBE6D9HwRMv87khFJHjvtbg9U0Su50P
H9vN0HZkQItodak3lJ0gk3JVVTzK2xNt+tF79pf5NT6udMdaB9gZ5GITjvYtr4m+
PQwiDkBWqwf6MiRNwsMeMcg7BBI1qGQXIyKxxMK0A6aFcLTSJa3h5d+seu9H6+r2
vbkTQ3eSEPyg/uQISiuoM7N4luSSgyRb3cfFfw2Yb/7BoMG34T3O1tdXg2YYlGVV
iU8KSvjbD/TLaURAOXNtMjtoEom8bg/ZSYKLBerlUfZUcHqbGHw3KncCchI4LwMn
N+Bt/7EbL4C4T2ARTNIEFgjM6k4AIpBn2w7xxU6INJOlOd76k4nD6brqwhczPS/x
Rw4rcvlW4Bsef+LIm72YTrz/5asQebbwy0AmYjhqYRQEIbcoJenjF91cMK3TzsCf
ZtZ6GXRYMfXx5h1/YEHERPNaLvqiViKayuAjVjS4spt+oMbDAcnypLyRloNSCufE
Twi62votn8e6JAdNN1I/N5vxTzqSLiZrsrdu9UpsaF/sQ4SyNwwyXzpVtM2nIARS
3TymEV32CciupWz+PKC0Hbp80uR6sjXigC/+doyU4lfJlveRKwAKGidYkAOxF3ZE
olNmTxLVyZEy5EwtHc05w7ITRtwHHCvz1TVEF6WMBtuOf7TJuxIYNNhnKRUIqT9L
yDPFIE/b/3a8IWk5Vlm4d/w7SBR9Qc3ScBPjsS2lQMEE4MlMYbwB6otVJA3Sghsc
1+EQNqqkK7AVaGqb3t91fYFvrXhL1c/g2UZsyWI5n/VdumpDKU04P8MAglARGEO0
nyQJccAokfc5FP+bLMAFhPcPhQXEXgLDuCbvi1GYs3bHhqBqU6PP5ewGq8qnJA6C
7nT/Kg/ykHZNaFt2X6rkKLJONAOyiwc+TNIOqZRK94quJzTxS4KmsbG0O2j/qrhR
RVOL0n7MQGIjkiUmZG/so9Fp40he3s1SE1HFEWE72zbHiJMlZOsxppzWXU8vBnJf
CbwP7OX+QMRjERidlO1RB5OZXnLjCti9HrYPtUFcu1CWqZ5GR9NvI8yi4ovc6r+e
PX3F3+2UpARt6dwkkL0FDX3XbT23C/iI2civQxGnWeHLxauZ1skOb1d3EVR4WqSf
QhB7nOu40N+pCwSw35vxOYe80zcCLMc8u8Gzymw8ZZy8yGdOXIR2g43DSh4gW/4M
bh7rG4A6PJAk/MXNZE+xz8lDb8P7Wz3OCtUe20MznI9pcOU0xofnssxR8Y01mJzf
sfYWDy3ZuH6TOG+LQzeIah5g2k2aOzAm6JYh2Y+brmjmhbG/2/NmcYRSNGuThKVh
ynoCpJHEJjcfAaxuHQi/ZgDFEUoeL6+SCQ+LE7b6t9n9tN1u0k14ERnbR935K+xL
zdJ4m+kpIykh8WpcYyNyYrPJwvtYKoTRu+6V6aBBtoU00Wts3mfcR8pzdpmvXICz
GY21ygvsqlYCMExsgVTG6v4Uk6ynq3XbjWHaWzBVl7qkOL4GmZs69i9q7PYBJ9TC
XNhqyHKI4brEEoecTfu7FP5X58/2Q0ArYfxJMZrpWtuDsp861y+0H6QLS5MExBJJ
HoLbHPOEe+k2vZQOgZ5mkhI8D+gRCKtoFz86cMCX+fUs3bcYbDXi8WtlL++Bx230
qED8q8uIcsir3VfVbltH1yqwf2nF6zqN9275qOs7pNyi6Uppmh7mz7QpxcBAEEnu
hC11RhHKiGSWczQMp77bNkJ/5C5Tzy516qD3ebgu728GflsgyfvIV7R7BJ9ItNuo
YBCLTyynEXjWR+o9CW6LxmKpP0U6UUvu//DfPG5CSBu9owhFycQ8oAlK9xha3sZ5
8j6aHt4IxQK7aBIZAkm84TD+8z+aKbOxwEAKFKiZTsejitt6urz0l4al50c7itzn
KskWRV+pR5B3VIKmPoO7b4OFlRvFk5pFtvNNu3C70kysOijFmL+s6g6I5hpSrkBg
F0nJ9YbZp4IiADcWokaQjmUVQYMelOaU6a/FBuIGCA+cuAh1yliMYgNT9KPL8BCc
i9j4/yoX4+6x4/RK+X9Q6hSJHObWXrjWuNx09GQi0t6VKac1nLQndPoHBnkoBuW7
yvCYayuOFEXwxvnaiYjKvC8yYjtLEJ7zSSXXkf5A8pySgTJz2LWfso8ZZJM4I7yQ
8HaPDNSTAWBilpwXEfSjopQnIRQRnrEqNDFXrM5aXYMzkcq5H3KbNDJ+9UY9MIiI
qkDXVx0A0gjirI5jdDZEjqJbKRCRS35ZAiT993b9CRlQ8KVeH5ExQwyX5Rr9xlWY
4GwSFgcGq9TtBpc9ZawJnnmQSTNH0iXA7F+FHmMNTzfRT3qqOwfNwdqa4Jx/J0Pp
gsTN0BPTNMioFR0jmKsBWeOC2W7pSf7T3IN4HLlaXu2KsbndxqtNGkB2cnTY/WKV
wDkCOf1RpHcBaaNxUSvEPPFFRgCl1VItEKLw8tMvnhmuAqhAIQ3tPHMxHCH9kLeX
5CGuPSXiMPxWPYf2vn99+x2Arw7nw9pq9MJ/mKVcwxbGF95Y/M87eAEEgdl6ebAo
Hu7Wg8ku8qG16TGWb7AHJIle5oGNdHH60+VEAvjIz4O0pwkVLLixfk9qMYGUMWN0
kd8MxJYpGRO1vQDTNDD4BRYFrUFRgfKl9UXEPqgpUZt9Tx0uPm/pZYHYxj2lNoUz
SJa8ePPnpn6h7IG4HGtbgOnikPIYdOp+mhfBLZIlRvSI+9/zB3TVGF7HLKWxDw22
KRdm3xnKnF3YksYBDfFjbOw7x5xXbLi/mJENJEaPzsVY899UffduCZBTeeFJqLNr
pjGNWbohfWprwF82ihSHSDJ5uIXRLEwo6NLM04O+7/BO4TgeXmXcUUHUu6CbTF4U
ZAoNXEzKn6Uw6FM1V2BCbrTx5H58gWOJE6b2UsqZ6NekqwGfIdjEA56mtlGHfqAF
BxOyInBcS1lfzIGPvbC7f5SbwussxjmwquVTw3Ax+McN6t+JaDo0rRAX9lbjZJAR
z0r+AvQn9PvO7jPG/J3OGl3orxJDNZwmbP5kXALlUL0Pb6EcSkWcz68F98G/NzAt
CA5mSLMmei0rKthjclGJr8ZpTuabcHvS+FckJtP51RdMK4e3uLhbTcsjh7201BPd
7fz7h2i22BQ4QOyDp3mjdbmwgzHkUkHan2MnwGAWQF/LgIbHK/gfqKGCvCvyvYDM
yB3IFRamloyYCGgWdgGukUpmPnWJIipq2w/DAE3qXHWModW1Z/H090cfh6friXSr
S+csSBBFt1UoZC1qFSLdVeVSztsi8p/haKm+Iq6wHUEuGtIlpgtnlFvTG3X2KShC
4g+y0I4dVJjAwQ7R0IIQAluGQj8qyU4CElmgzA5m1yXif6uD9x1O3W+X6ROBGGK1
HEbwyshqtJHm6qHAWhwD9bkFl8kgdNQcEYyeAKgPPo50iBCXwgu2zb/cSukPUnPL
4DAl7uKLJpSP5wIkMMlHQ4E/YJz9+O2Pz+DYx3EEPip6u9tt7rqHOubwe3niNnkL
bJ2V1mIEeZZc0yIj3QNnhRcxRnxNFfvdN4qmH9Ifn1R13PrUAtXiv4FHOQjyws4s
b4Fff1EzqPKFD6BePENiDB5lqVPHni8EViELKFYuCs7SLs1GrFz3PgzYzNtwQz3i
l/IZaENP9pg2MU8MXNrYM5ag9IXVmIomeWTJXR0QWqABs9R69u77Qeu9kuJ40NGY
lAlTUCQB7ltUH7uCVASpfHyNFH3XEWbz8Bi4slOUiTmv6++cGRhAJZ6uZjAdum+q
uu5iL3CaWfLUVk+wp8jKfupJHQ8wqkHOXygHy0IN09JxZbyMTOT+PEUKUUzJTMMR
cfiDWUta4dmzhipx9wL7WufbSNLqbx/oP6e1qdoQEXjG/OC3Uk5E78gkTeNwgEyh
YUfXNmxKEy9nHnRgq2lgUzSRHupgYDQzB5Zt7jt3aG/IC3jSjoU4tBAMUsTd7Sv5
Gm8i+32wA5UHj6zfZ92lRfWzDoUHRrQfNhONNAoAbMaqLtkjFXjahVa6Sa3gpLhC
8pfbYZnVAVKxh11KwS8qMGcRunQvENjsXjdwZ98ZJLyqO93nK5a51KVpHhFhYbLK
9UstznJujlZmk/yDKx754wgVnUSQhCqkanyo8k+fvi7pFIRMbP0ePEHci2yMPKbH
vzWVFoLF/ziEb+E9ksW8Zp0h9apPPo4zth1+bufaCb0wsDgMmG35ze4uMNQC9f1J
tvsJGq0Q/25aQHJt9cSEtCqWDFNTbRddwuH3nMdEfQigNdMqqNsB48UeWfc+g1mI
CjvmuXV9X1M/ZXQirdFD2eJ8vBPsitzFky+P4WLbDEGgB8zHPxplL/xqcdNxptcb
aTgrvEvaOJHL4ERCuJxJLkjPs/cwNB6Bd6xmo/gm+Xry4LTC/EfK63OIP6fJ4jgu
7fJeztQHBJccmSsT8E08Im6hdkal0o68t8b0ePKBJcGF3UOSJdlje5T43cfqlqch
H4ZGf768wOwIkyJbff0H1U75uTv4GyJaRcEetw2jbuq08kEGmg5e03bnGAdbYd7C
kzpiI4/D9aha/t/MjfIE+WkjPnmDMTdjKP9xTYVTxsly91Kw3AZ89WI7vkEqtNnh
JJ5/w4BBNiJOJcELzkVDXvLeawleS39ntP265spMMTg7UUdTGrlLkY2Pl8Gplyw5
XsSLH0a/k83fH7C/bTStMsDbuPqkwzE4QPIqZ/fljaU4E8R1BW7JimlE+rhr/mYx
QWsOUxqgJB7uovUSE/Hhm1Ar9CZzdKG1fEY9bAGbE92T/0+nVry+XrRda7w/8KNF
5xiIWIpYCyHi9ZUJaSbljWHtc9pKjNsY/eq4aDM0bBHw2UZELyzUPm3rWwYF4zUp
WFgpZTPFQSGcEM+cm4FgN1ycS4z32QbBxbQThnXDBdt+lkR4sv9S++OcWQxqNmzu
6Ze7f4KhJJ0K13LyIHUDoLVCW7RCfzSYZIDG8jA1K09Sk5/sANr7mG1BBOxNXJOe
uZKc/psecrGWIgKn2cl8Uf8G+s0cIr4l3kzxzU9gE0b3/vHQWkgW73FN//pKrKGY
DB3pbKDY/RYgueF+EBjpSAGNJ8lAtMII6DjXmm6Gk4rKl9wdpJCfumuxe5AuUyzP
fqRr5N4FPMvWpvcPXRzPyvf+tDBJm2IMACceM4B5crkq6/tdqPjsWqco0R7nnfNS
g/cutIaUF7AqNWTCxSHuyf9WgNrnXZlcrLzCLtlHn6PO4LCmMplvjGC8lOJTQSqk
ArDnIeMuRKyYXWtwi8SN3q6m3WvIzySFY9fLsYBpyweu/pUL66Kyw5tlkJGEPyTu
znpQlE3GJJxJaDqJ/zO53Fj92Ayv4OsjupBByMqWs43KRfweToUjkyyfphxzAzxr
Owc7/j008Aq9z0LdJFLOPWAMyi58e06CAxFh/fyL+JApEJzZVdOA9aTnchevlRbn
9g+jNJtC1F+1SizPUNHJGn4ygAHOJmegClnh01C/VNmmVxbLRCJuqcAe+d5SgFS/
GH0vFzKGfUuHKP/ACqt9o12RngQQHdenM21nQ7rr37w/yWCIbjGyY2tr2G+tgC2J
cDLtAif1q8Ixyp85LnohwYdLzx26oM8WWSXW89MaWMphFNzqNXYwweQ6bmcGMrnX
CK8p1oiWi2VLm3U462QWZ8JP2toxKHnDijq6k4VBH7pihj6xP905pQ8t3Rao+SID
tDGqyeOrUk/4U8QALp1s6ONzczeQ8QRUFz/05PFEBKCIO4RYK+XgWz+pks4Mz4RA
llVj1Gvxq73qUPPDGWymtFcxku/adFXVx+vRQRLwgQzl1cfgbvQmwgAYRMenWVL2
8jyNPT5joz6KwTRd5oG6siN64P/FaiuWqJXKn2oDW/UE4WE6vwq36XdC+OYCNTNY
131HlcvJCubjcGw6lyBUvra3DRg6zqnxUEoKc84z9I2hsxkwfkaqTpqOVGudmmvg
XeT7yWcTic3plFzPlK0cyIlErStnxiDxhIPt41dEMwMGTpUNaPcSWdp2Flcob10A
9RYyueGfVdROd4BA1QjLpYhbNCeAPITywFx6QrIb0gHX3PFBl88Gi1Pf26fbRnRW
rlAYQy4s+qmwBRdCHD5WSq95JDUakvEJSOtcKAo4P+bzsGu49SgHfveF54h9kya4
HUIV766GpwChcc/jdZ+hheN7GrpGeLvH/K6Nni4MWsuUzrFQtYY5mHqudPu5GkKq
ngS9iNihvzNqv4zhBjynpCbbTM1XAQ01AgwtkfEiP3ZHwmFcf1PSV9umJ7iFpV+I
vD+oJcx+b0WMIqi2NXPIA3IP5a0ckutd+cDS8x5pSfirWet358M7HUbllVZcxecO
QCxM1lsziMUIUX4N/xxJLHVFgYWnNDZtHkd/Bcd6AfucowdhcooboQvOZ0YxWnvh
LYCPSODKya8W3JMlbbfstya1qRj/QHxi8ZT7NOwTza0txoYL0nJpZ1Yik99QovtW
t7cfSaVbqCIHtEFGlScLo7JfCG+e4+iIHkS2mX22aIHVezzzQDP8nxngqxN01uI0
AmvsOJaEVgbU1mz/dynX+oFO8kypFaOUCoytf9zFU+D0vO2kOfO8UTNa/iUMn8X2
z6qm/VPlqLSi4vJhkGNTOxh8LRKH4vHwbFI28BxDPaiZHDLYb6aZX80HBE/T2eGG
0y8dBKfxNwknkIvT4oBVLY06BDaZ6Ltk/ursR939EGogCwcHkelHe9PCFG5347Ap
PaqNu0DXUzGuc9ZJa6EfRkpNBsswQmRkiI+CjgOVOKbKSp0zczUVfRsHqRYU3wt6
kS7mIcHvWF1RBgQQK+6NP5ushVs09CPgFCn2POb2yV0uX5WEb8DRYqGIROmWfj98
QS37ao9ct2oEkgaQsaYSvyZjoUjh98sRKnmFH8BTTfXiPHfy4UuO8nWEuR024nZR
recinpRZAHEZGfNIrtdz3R2BHsdt66bwKIdbTqg3TjyubzoDgspX9k1ydKVASrsO
D5bxhF3vSRqe8WINpUAnhho515dY5NUEdSxfbKzmwz/qc3jjPa0iLaOB3pY50m+v
+fxjojtligCSm25vGIAWOmWVDohYVnLhmuEP3rs8PK62MPvvnNJ41z8BW6U/gTgP
koWE0j9HRq/UY3XANSg8Mc6Bsc6AhKPVzhY16Z2r7EPXbkY/Nei/tDGBbGfj3UCK
byv9dksMRBy0Rn30EYKTuW80jtd8OTYp7L/X3J2SsyjsjFqPqlqSUG7hDbwuno/c
SLFabgCOTnxjussnDDgH5Z49LkMjTMNfKmkuOqC3vnqfJEKsFUU8mZev0NOH/SoY
y66b8b4idMTgpPDZ7d85jOl/TDWJyq2Q9TqOm9ZmdjieJnntgla2/16kgwxEbsws
ALsFJnfYcvokZhyVbrXzFWpi5eZdTBj/pBA8DZlkd9D0u8YVENQbudVS09AKftaz
xeEMCoBOGL2IprttCcjBu0T0K6ghcixyhxJwfc53FCjFC51GGtVrofz1oo83ELv3
G+RYBGd5ewKGxcAb4CdkDFo6KtwlKsbSPzR5Y0UpbfqpL1SNHPRnzaQcbhsiybG7
s0G57/Sq3Z2UeRdCPS7Vgkl+OKMQhhvA5zsWuwOSu6dTEfYLee8BFqTJUilMeTxD
JQPD+inEPyTl+3YJw8YnQi/TJ970NqpJDR0o9waEVqPvQTHU96ev9lBY4y8jj2CJ
inpj4aBHQHBMqFziI4O0xwsFUNfThh8M+eDuRLEj/+ib4OsfU2pY0gH1A5XY9m1b
++WHZNh/jFaXSseEvL9Eci1PhDGlH8D2ch5RKQaS+e8UoOmpJTOa7HavUWD4BoSU
OPfBWyFU9cJfbbaCFEEl4eV2FuNMAmQ9TWVd0pYPWtmTtYiIu6mlxdnpohjV3uTW
UqSo7n68x0D516wNfFmfmYqmFPMjmyG5NTaE/v2iYT97q6NG6hGBqVSl2Iyv95/T
Af7ZUBPi3oCXemY9ktlBWhoeLDx/w0m7RXa15G01c7UP62dzZyWBh7KV/QDc3PP8
Ji3Fmd+aPB4uYT1h++WL6JrK987uTGkfgatOhempxUGFl96adOdM4vyCEaz67F03
yITXdkR2uF8y0vJVdvCw6hGVwhldW4sw0vZLYXgMnta76+vFbzrCucIK4Eoortl4
PGgAto+THVS09TTYFfK64hh0m5mtCFiUbqDOjKE4/IPyigEY/zBAKe6wuZUVp14+
IPei+l5mdOVokTtMjKyBb86CbOq3V52AcvtWdQ8rboWXjz+tnw5hFEu29iQWrWt+
qoUUkm+aZr4rivsgndcIDyL77HMmd2bCSdiXZRh5+WRSrpKu37jLUUiT0lds/j+e
jKblBqnJaRN+c4rbo6o9d1vdhupl+wgLCdhwa94V5Ofe1BmW1YWXj6DAB+9Lpf+f
GFma3sbToOFs33jHZdiP1uAakCUlK6CRp5xjzHal58d9Uhio/hnu7/sriS0m+f77
9M0b2uNKU8RoSE7r+GjLdPnqTOQ/30oLHMQXLRCJ2CCYkEgjLVuUuoiZCcje4NNm
3n0iYBO24tTB9+kKr+F/i8AUxRNNz3a+JoJ9QQGxrctufunEZ+j5aVawLI1GFY+V
hkHjl2d9LP74ojDEo3ZQPowyAwsF57NGDZhPRP+OHw1KSzzJLr2vNbeLaLTGHtk2
dmkIvtBCiPjkjQlHk2ixPtghWdhfNQnZxoTIBNEXggOWK4bL82KVSoI5me+30oFf
8d5R5Cc6k7/7xAbsI3X+4L1+9AHGpQY6MtVItLVRSrX2zPuSJtqBEDdi0tG9NXlh
V2bycsfAKf3r8QOtZDlrz1MVnxpifkeqykFetyXIP3809i3dI6OsRz+KSpMbvViG
bhsuJuwpQfLVL4F9oGRdYeOOMPNPBDsWh4IanmnT+wPrO7+2Aix4BOeQOJKfzTi1
pzpXO5HC+1nsVMG1euuMI6t9XE+xR29G1WyfHiko0cw/f8e1aHrFLa4Nwab4QDrW
zE9hG/WSQiV2j9kWcTTbXrJY9lJgUjO6wY8noOKAmj0l7IY25aD61IhUbMlbnGiV
0rXwfI7PGVUiPIFCkc6PB+uVON6lSm4HT4YE10/EkAsUbnI1nptSdWL6e+2dowJ1
5KKEUR/QaksIir7Th4PLLlgvbZ1C7b1vmaAw56tONABb6/N51qOfLrjHMsg/01kc
42hobCin1/Z/wVLSVoPfYRrbd/MU+PdgwkFO/+VuvTVUE+HRRn8Y7stTne6MgZwD
azZoiF1fSO54k9adnasC+tShe06idlJrQOflcCTj18Cd/U1ClY/sE8sUfXs0PL1j
jmjbLp5h+dltjUN0vfNJTA/CcEh8z0USvjEUt3j8YpHS3l5qxeuuQxHdoCNiS22u
g5idjKd4n0CmurmmFfGp9zrcFP0jxUcfPPYY1/WGmYurQmq/uUmg0dgp2wFf8FKG
Hd5c3z+SbNI5v69Zlu0voPAAjpbHpJfcvXgetVA+VovR3uHpoCdGA/g+zzaGn7sF
YIuiTfcCKTn4zLDH8fJfbZFdtn9txwCTBfbb2UEjjpkPnO/kdxXSckI9AWtSfLPt
L9pO27KBVTo8xmFS7uoAMdDbsswAyEETE4i+lhMAa0U5bWTaS/fRU7tYdTDLN60h
/3uDvFgPATUQnqbtwUWeCVKxKla8MjhCDCbdcv3JYzeh6GoqpPblvwJwwoOX/6Bh
j9vbweP7yHCUL8zmL21agwG1otmSvGuIpeg5aQw2SM//TsAkAVVOYQWGR4axmVO7
e/p6+xvwJtubVSgGuunQQ6bE4AfAA4oxfqSJHnjuncjBowVTRfMx2dlbph2WuWDG
CCdToJYhNQFn/FvLUyIhf7kwyE3rFCGHFQV7i1lN8s1QhmAUxonXN/d85RXU0x38
9HS36V5gQ1L7+g6dQZSe8uE8+aNasrqJhuE9iPAPo6bDYUA3+NQPC3pJKpgsjZqB
qG+pBH4SkgtHkET2YscbAfIj67E+ujBKROE8Bl5Td3LReoRCP/bHyjBGhvywUzoM
ulyQABRet/pWb9rQNyVyWZhElmPoMRQEdrMgfj8Aq9IVDZuOzfma4Mlk60o8oCGQ
b3Fq3Kz2jcNapVRa+B1UWLBQBju9so+uHjkUidzAgy0mMB2Mhhm3cRXC9Oaw2gAp
w78GZTquoA7hYrgKh6Yw+7scyhj2nd+WTRc7dAMNMxm1uI+f9gm7Ea7PYvdgHAYj
biow0S44mGdN8swohgwzfNRR/TCVyMqiDAL39lvtYeTTBbwlA1R6mSJlJT2jGCGT
rhhkcDHBGMZfPnm8sq0Tjw5yHFw6hUdd6CT98SICjN4gAyr/SXv7KbLEOoLtDasy
EfrEothxSNpXRsDaA1ykEqcA8h4/dL6PgLYfQeZsdvdzx2jq7Y8oNFLxwyNkw6ge
WrsunoWTx4YoxISyUg2PFu6JlgSx0e+skMR8o+nkh2+bq7+4Y++Gkk1WSSvj9IFD
fgeHwEl7y/L+H907k7kH5oVgQnqF9vWKEIoniWGQJWKA837i8pfhEVow18xZA813
tuKa3dneUDMBZnyPXOq3+np8oLtvAJFu63519UjWsCSl7cjLnxi2lPVDVHenUwdJ
LKyO1hqUY/aLQ6JHjTwr0q4kw841tDYGD0HJBPVrECO+uwt89RRjqPhJ049ubf7z
lJsy5HNuOuxKKCv/2oDUZLxm79KvnR7T6UyZIxYWNiqXrGFU23sBxBEJDGGp+FJU
Zj0FdFxMVudxHIg2G9V8T17S26vypRWugt1Fd2ZjgSP1b89JGJ2Ju4dWOmD/+PRp
s6V6tsp+d/m+U2Gm/73BAr/Sgk3uzD+bDp8af3Y7KjtQCax/0NEXk8urXWZ1nzJ6
UQwRuKNgibcrcRpeVRTv3aAzcBL2GQd3gDq7E3ZdV5LSIXBc24o/xFKeDyE0U7fG
Mc5kMevG5e0382ncKcnv/a7lXcc46rE/eO4DOg+zf7ddj/nsodtIPpdz8wRUC8MZ
a6sXCcmZ8/R42lM2TVLAe7acQnBWsrdMWENGPmTM6MNjfkvjOOzNrHKlhwiQYLF0
27gFgrUWsyFP8EcsHiijF8eBTeNLUwMGRnJT93rpNsRXN8hi0lRAY0t20bhRHhoU
jFaE+4rewy0TdcD8ydSMxJuKQxL7JhB9UqzvU1FwvbEkxJAVyr5r+5L4P/eztCyT
q+M3j+XWmE/lQtDWZOwakFHnGXkxs8+n0usctMTstFoRFJJ71Iw+Ukh74YhcWWze
CSH4aD9LUIB3uV37M7GPdhqVQjsL1S8ydPDmy9RauP0a5OpcQ3pMG9RtQxW3fgD5
T/aISqndIKrkTKMTLmEhPDLXLG2g+MeXJ8kYeqYM6kEFqC4ZP9TEBBgyNB4YeFUU
Ii7WEykN8f88adRATcTHRsZuyrGfsYfVXCDd68HEX782FinaO5/Xqxez9lPYmXzm
WPnLJRZbW7FdZTYqCchAzmrI4HxnsIYR27s3lL+VXh9sYOP/ZHkKxUN2YDPyz/OV
y8nwhq+nFYuWNxKMS95lABb3isMsE+S8BSCvrJYHe1HrKEVWUeYUKCncWGlZRtqt
iN5V3vmc4kD2nHIERghZxgnE47IPJjSu/PF+4Mw9YrYvK4RZ6HxsONj+MjejNZqg
/tOLrgRevPE3gd76eD45NjzPMs7O+zl+9zYMBI2ljPmU0LNGrV3eKRPocQ3v8q0j
TRp5aeCnBu8L2j3dyZ7tVtYDvXr4q9yeFIcDgQFygQIAFvQlwv3wgjPc5lttoWol
+Zft7TEULMzw7gCcPeLA93MJKkO0NDnKx2K37thc/VnfCG8W/A0NtPeROeFhM8kM
uzRzuZUstuMYrfES2EFJVZjJtiz8zb5034ucC81qbLq6yziYWpYFKTyQECtLkFW+
trfx5yHlwzg52JCJhQxxlOeOFdxV2CGKud3c9aZa5x3SZjfvqMGaabtFiL5raHCq
z3/wUPiLMQCYRZlU6D4Qkb0NbO3lymRJgnEnFNbytCG+8++hahrsXISFqrpxnV/T
/vb4VIrYea2VcqHrADjzT4pWT+8DcD2WKM3nsCwMSw6GXYTgiKRVCaJNX8TErmOR
0hWSPr0o0xrNLl8i2D92wwQgMS+sK6fhYc3/yVO4gTNfYDkaXUSCsEpjmjYVkSCZ
jy4GBYDhbXhu3QEVGcJS9SgmkjpIoE7mEEuGPENWDiYrimjFoOSx5HTRtU3BxHf0
v0J2nYBKgTJRPvOSWcg2Q22VBLpM8y2ijbv0nfP55bLGi2Xwi251WrbSybBROmsk
7q7pWxmrOfYy2LYijVah0Uv2IuTqSEkwrSoQyyh7iiqXKAKVIDMyevrfnV2B3BmI
A005jJwzQwqvbnTBbH4gji78CXcJhX3yD2Y+851B3I+7WR36NgOcBXzvd8aTQqHE
K/kU7qi/lgxgun733HxR8MUauNWqCKCJLkARYi8Vrf1wLqCWOUGHPR+9d+sK6zX4
Nhiq2sA0xPGCE0B+9qW5yITVC1I+RmDf6g8ru/03GTZOrdO8d7xa/la5DgraztQu
exLOsB/l7qpgBfH/uDKHCduFJwErMyZHd4lr5Wg1Hjak7U+xewK0nuC7JTSF/zMb
z2cf/tfqHh+gvaMLRm0kxzLaiIEs43Na/LcYwyJO3VVBrnFSRagjOgxMIyWv4PNL
pJNNmESQCZqmH39bqwEY7XYP6V3eK9LvFVoKbQ5N7uzP+C9aDdUWdJdyjB2lX5wY
kBjm4aea0P682R/Oy2ncWJPXxaHz6T+RXttGg1HKUiDkrHjs/9xK60RJFWioeRnB
jRZmgxHlVHWcMejRopD1d4DGoER3a6nTWHFq0Z4z+dPMmG4kJeVEpOeD7fxJ9TFK
k66R2gWVh7+JN9LKBhxuJynmfZr/wajfrI2xbrII9JUZtuPjBTX68UP/voR8TLEP
UVH+kUuwpDHhg578l5lKlpldf6KrKga96jVGCJEAmew9U8SKIzLYO6IL7gcqK1AE
FjgwUorM/ch3l2fjKB+pIBTeC0fn2OEfPrpANwULQhRaUO0wlWX0IdNq1EaScAQL
5fy1Aq5npjgEH7WmLFyqSSLu7fVB/RfndvSanv2yVbFVqWvByqbRDxxakSwIYfVA
8+ZmJfiuqOGwGjDg3Jeym+T55/DsuPZTkyKJP1tGEgJHsTeVb6Zdj1HtAhD/36n8
B/ssAIZ4MOI0C6p8x8w+RHxComRIFyUN0BVEYnXnt7ug+2b+yXdVePsq9mDPzxMI
+wF2ZfxzyXmfGPYkK2M+Jc2/gg+Z2u1vM1xhKsl6k8kNZPTQjo8C6CzGA3EGzwA8
lukMFLIrv9WrAZ7HnpgDyQvx9mFeGVejJXPeXVxf5HQhaDUyz2wn0as6JB3KubO0
UHCBg8FQN6FYYZtrY1hO3MfSWZfLwLVGbUKbUsGyig7/2193kQuEFtmsiOr5lVln
MXVuO2n0Y6VO/GVuJktzZN/x8Gpn2W/V7SXbWXiSpXbHgvWJr/BbWr6skPaUJun9
t1RRToo45j/R2weshVNmdJw20TmTMCw/tCA9MVuu7J3gTYU14BtVRP6daShYg33S
sZ2AoXdOu9d8uZ85sD8luvQSicXSSpiF+CSbDcZSn9VMBbq4I/4rTS3FKUxXPWw3
Q0u4XcXmwPJPhDltC6bPlKBxt2pikZfo9IjuLo8siM2kHI4kjZH0/SUiP0AlU3/s
/xdv4LJQEA6GzoQ2LWT5B/cSB2f+9zHBhNCPgCRhkM+f8LwqFNz3dnZ9d8bVhMLx
oh4KiLWBjKIaXpY97Y1AOiilsAyEDg49qguFZfAplF2vXmvpgFxrQUj1w/h2WsdD
5KdvCAcmTyMCNuy0k1sM/NmPm14Syv8GjrSUkrE5KS33nRSBzOgCKhR/JW9vD5Is
d2RoiOebQu4PBprO9UGmyPZUzqsmWc4aSr+jx4hpcxXyFdHGfRtOpAD53QtX1rCF
Xfd9qJVELxvZ1EJ9b5hqk6Ruk1seCW79/uKcpGvVqKNXCI4Pmg0VriH+29mTGQ/y
KrmQnYNVcZQ6vldyJEwNgo7c3vZtDhlN+PHHCkm2qwUAg5DNE4A9jT/wyXDjaeTL
5FjyNKdMiAddngGM6tewn4DGXV4DEbiLC8Dl1cLGQq4N7ebWa7+BD1CKp3Ig/Sg3
jvN1+NJpS0aeIHqjlKc7P+wan47x6Twnqy5KQBkSnEUqvh6jkORpnfAy0HAxLZj3
uH1GWXZa87NNi3E819nkvR41hlTNt+sU3mhh85ZUGw6YLZeF7PDaCOtrzfqwq1EH
iihnALbaNydJM6SW4YBqbYxgeOsutkIxDclLvu8zWD3QnCwDFDWYp7a35w1Pk955
YjqbJEBxeMnNux01roWtd6dTr+uWtE3EtNXVyi5CZTFe9cCMYzSRXyFAVIBeTjqc
JyQJiuLtxyqVoYCnOOeJDIewnGb4OAC0cROFdMbNEPL4T7UErykE5ZXwZ267/hNi
n1GDanDdady/9pE+sVH9ZCeVZSfmK2XVzjtP5VvXxkbw6UTERj5q/oMbj2e2srGr
iNbS7M23ps3Vik0jIFL18C2YGgKiFT1COmYh8ItkgfjGLSYhjW72djJzHESoFc/m
g2i3XV7l7+Ig/wT9NBDn6RnyGJN0jhBSRX66rBjVC40isoVejPVqsnEL9wqKN148
aF9lu92G+sCUxcvQaJZFrTZ5E2L7UGqREOvHd2DNEn/xeOa/eTNqUJ3xzSoH8n0d
8n7KYBea6OG4AjezhChiMif0xs3mI8gfiaddwrZCOEnrAbsQmdNWJy2ZLey+he/j
9eEcIAQb5MU39UEI21iHsqz3x8QSUVOLJSYBWxSHaibJK3j24aQSyt1nVnNb6Vrp
cV/2zafTljbHvQXqBEtxsbhNzinL1KiTC2pbppg6L4eDAccAqhBh7pA/KzjrH/sp
VUBnJ5EFCZTwVYDE2l/thFay5IExikQSe2N9aVqf2TzbqrKP9UocHdbbLgHLyRg+
JVg+oTnaQOYi6Ld6l3kC8dnMLpBHQiHmJ4C4//lHH9fYVtzWcJyjF2TmlS6qxisD
WClXWTwE74RnnXzCX6XmEKGLEzoK+G8nM2c3fkXvkFdNEP6jOxWryuUI3qCH6357
0pR8XjqCMHnMitFWgeTjuqv0/jtPqlchIUM/e3Oma1tgkeo9Bcdd+QBvZGCdjhsi
CGkBnYje09shT6lPidUmRWrTWJ3bYvjJ2MM/pchjkxIycc/kxp9N/YzhCDcpiwEP
6b0DVUvWX9JGIypo6d5L3R6+tpZTo4g/zOhUS7zOmvMV11dVy/hxlnkdEyrPS/+d
R0v9dAwM4ATyd9VFs1xgnQgLFOMZu5umCUt3KL4xOIVGDwp9gDAs/+6BP/26brP7
E1m4JQce9d5x6y68KAl6XotXa13hPAjR+xTxE+Y5KyaaKrxB0hniNe0L4cGnA09c
oGlA6CsoVuChVRcY9e7gwj8Bm+uASYFKqguBTSwZZANDeVoSTaZe0mFKRLm/trSm
Lv3jMJZQKXAI3Mh5QiwCgVLg6sPHWEJtNFfO1aqTktMOeFUVKfRn3hXDI86uzm9R
OUFAflbpfN+dBVG7FtH3bdYA56dPUvxSMWBi9J8F2E3Otush8XXm0TWn9VmclNdc
TXQ9lTRYthpTeV+3LAw2vJJ0oeXPFWVbcK5dzDUchxv2hTHiTWg6tHh1ELUJgLEz
S1Wi/UX6qSt6QrzIT0ruzaYw2x/NFzpRd5oO1BHGlCs2vIjpzjf9FY+vYQa9B4/P
GxZAQT/D6dLWJ0/KWiD1i2PjRYA+0QaxODF3TZlV9QXgan3yccTaWdX/r5EGZeRy
hn2qgSVTrvb1TFElF/tdmt8byMDAZjla3yLSEEAAtHouDT2fhsOcNxSrFfJCMVz6
FMD+j/JTIm9Qn/yNsEBUmKnQHdnoN5wPr5lBQ8/OYwalJ/h+npuVqAUrNaSq8j4u
KoNfMgzuq9Am2cX9BPUKtsPu/bdFem83dTS/QOAl2BIVgV0iIAzdHs0+tSvvGn43
WO5gEfLVdOGQ7miOvnVzUDCuNdSYGpXmyj3PyTWcTDQCKUU7cPVzpgao292G9HVJ
+Q90OlF2jLFVwdTBUws4Wu/mBDGJAgk3I08bCkZUyhywxgcG8jUlqv/jVCuiJIMy
0Bd5X5TBKQDDBVU4mp/WALymJ6wIqzAkL+YAg11id4FdKPu3mk3rZWkL/noo29ir
QmAzM9gabWYWnWjhqhEHmB6UeWzpAY7XYMhMdr3+p11EyDuFejxbhz7xJov4+Upt
ew4MI9dO+2bAUq884bnspHGGyNPK9AA/jjf9RXrgKZjID7CHE7bIukND5XSCGY4+
oMLvy9ki16yyROPvdedoyCCu3dtBB8FDinnuziruiEDmvp5fallolWjBPFRhSVfE
rsXBrIhTum4BJdp1mSOBVFd+gzi1o47hzy8pD3XYlPTZHUzLevciFznzgmlwO+wR
EA0jN8QxVl40I8JJOMvefYROmApDEBzxp5lbgzGxwI8pwYgp81WFIJIfH1nOqznE
jCDGfbUMD4ufEqHK+rJvWz2Tin42ERB0a4794uQACBTBFPd8OhzAWA0JSKCozOyn
kwDfuTNt4610zc6BP9uyfLGGHSve81OhKLyJX2XPU7oRqF/aaZMndpxCPfz3Xeuv
EzKWKPViTGA6Bpz4ow2KTodr+tHrBvQiPjXb7eaSEtCM8KL0yyWb+R/Gopb1KMy7
4FDcOae2z88634HLuLdgGPVMZB+QtyXmVRang+Wyc9+QnjdP8n5kbihYZCOY5Kwj
rM4fUcseMhVBiJOvSNvmsf4tpa6GxmgGdJUN7LzpTBiaTd+MBAsKcpVxtmvn8ORt
WbcxzpBDYFcyCfxWktKH9kGHC0QdljnVeAgBYXFZ01aZwPi9kU2q3spbARkoE8E3
gRamb3Ot0/x27IOg3dVGhm230plyTloWtIivuLVVZmfbYYmqLc0ndigpR/nfFvUt
NEdBI4/GShbT4qsH35U4K5mPVk3mSl+IyuQWI2LOnl6S9BDCyMg+p/Ctx9rknRe9
3P+LhbgMEZFuUkfmoL/BDYr1rlXstExrzSk87+vpzWSl+mBRnrNlJaT4jlaki+q2
n3b1cyKcFiOinSTxLv3zujqBXarrG53YXruTWIGc68bZTQSoElPiHD6h/OEibZoS
b+hibPDL19Sb8wMUqadW3a5kUQHxb3Ja1pJSBLhXgul8TCT0a6Vc/USQA9/8IsOW
922oTh1YNQbfzS1MoUu6KYrImbobqWmx8Zq06FH1SNCH4sU/DErg5tihroElqVOt
1P9wzCIUps5feBWt/Tv/esGIIFWS8jr9TMdQqRHnSdor4Tg/20NhQ2v58P3s8tAv
zDtfQaZ8UJFZPI8wq6mbjoixiV+0OIsvUt9qqkthJVrms8oY7oPeb3wDqYCqHbBw
D5EQj1DuOSDvA3h85CfgSLYoXBxlPbgQeLsj92P406q47afotOvKtIFqfF8S67ee
0wkzkJ/dHUHkWqu1S2pVaosTSJnDr0jtxrT70xWfoFmiv4TyPC8wRntAQzUp//02
Z8ULeplQ5gJfG/QjhLRcI/OknclbWc8ezB9dddLo4sxpsRD1dJ7KhTIYMOjZItRS
YWjderbSNwbpYAXRnLndlf9FpsvRH6oDVFqIXXf2V5XkUtRC7oKsZWypkGfiO+t9
MmTHQu8UNPK0NvXI9/jVn7oXUUxBrX4p/YVX5gu3lm9Bp54rZ9CvXmcSVf7UsvVX
ZLxgTu0uBR5SWcYDOQQLKnDnonfE7qM0Pv/FhTXxFW2cG3aHcWss97r9y+OXdbkG
sz9/SokbibQPNjp59kG2d5OakS+9s7Ho3UrLySq0Ml2XxiZgKlYDnZZH9b2zIPi8
QJ1ImH/DgUwVruqcl8gLfWFmZXDBW+Y9I9iJ0DNG80Rz9edTqQoWQfKvBAgK28OQ
jOH4D1V8wt1R/z5N35BkbWyDfw5ATr6Fg/ei4hNrARlfndGtF04NcsqKseODCtWu
xy6Mjs+w0izZc1Yzefc1CCbRXTiZ0dXvfZ8+ZMb68w34xOq06mYkXmHVzCbg1ki4
LQnA6yyvVSOnGHDLeTWtey0UFsb4aXkI6E5kyNdtzxNT8BXXCCypaiLyjDsTyEGX
592vbdiB/nz2omTuRtxTd0QDSEKrF6Fyh+ZGnr3yKkvSFfXIS09SEP0d2+rfYYfq
ndXMdva0DKte4yqbnPBozBLDU4UkwHm6NA8bLzp2ZsfaaYjugibvk4wW5hpSyH4b
9pQ22NrGc0R54yroAauULjdwop92hP63AA8dr4t28yp1dDeEmKR4t2pjzCwfL00k
4GFLHJNWb+yb/9VEV0OVC4fe7IB+LLjdLr0WfcW3/zzv4TJoeDYKQIyg8HtmPIHz
IW+Ydxxuz7YABrolJnofCsmP3HlOsGu1/Xgtbcu3bID5ndANfzL/IX8QrQm2O6j4
xCyUNKT4kSXIUuiqZi5sszuXzttEtwQkCm4nkW94bh277n+e29Odv9/vshfApU5h
P4YHnpHCg95jvLmqq5snW/NUAtrFHGxeUXyCzptSdC5fRO42k2M52Ean3YjDiPWr
QNZUj1WyAHt5HiJH8l0YPLLbQOu0osmHPDQMqG1UdVTemnG7Davoq3VU402xTRUs
mZQrv+EwOxAtb+mGJG2gEhuNThrNnyzXjJeJcRlGYUtDA+TjDZsQephuWpHwFMIy
sfD3nWrGiVn8SUvGSllrb9OgE+Qh2dP+0DKtuaTTTdPMXbgnDTwBpo8XUk6VOMv5
cw5rNpsmzbfOaRVCtTOWBahEyIDqbjR3/j+/qtvVBK2arOirC3D0QLqRYfRubTRS
NrY9ulGNWghzgmabZ2ojMgiEhOJp2UVeGVKPYxvnC4O4ghNSUx3st5+4Fb8A6WIs
5mbN8Jos1an0f5EdZ3/C84Q1rWxyRHxGuF6Tpquz49G2hISCO06vvl0MRfa+Jacb
01Zv58dJSec9JB6FqYlKiPR3VoHoWXVJosq7cVMeN10YW5+r4QBa1UN9z21nwoI+
9DZQyGOYTYDynF/UAc8pp5/7pcL+iLMiXdUd/PuP9lchtkluhK3mrW3nwyd+w4QO
4uT4qOE0OS1WbpTlLdqc9VmKeuWWW5at+nPS+WC1deRD/6vdu+0vTOfEjJx2n5/O
xm30sqpq1trwKe9t2lXt+TY5R/3YWVMI32f/Dq4mPt+lkA3ql6ivAHeRrlM0CKMa
3nCmFrzDhxpjGrqRD01y5QNGLzEwssk1JE5x8GWTGiMKwWIwkH7VTt6YAaA8hKW7
VG2Mrm/lA9HXt9czX0KSe3vwV3X/PAeYmQtsuQUbLko7WTQk00eDuMCWQwQdhit2
cpHF31Kcc2kYLkx3MBJOu/VYihLqevKtYd++n54uAymOXbXxY7bhZlEPQyBpWUgj
NUcRwv1us86mtBDwvkBl3Yn/AC0erLGMqwWijZoB70LnQp/MDMsltmXS1F1OIHfI
+rczr2Bw66igRukA5yqZxDG5BAa2htyu5RNXWLEaXjmqPM+hw1ZtQ7kjiQBuhO6q
pj94lWPNy7gzXjk6XrkhtybzFpTJaBipfJw77OEUgVbgPHUqyvYLhtEmbruY9Rij
NWx/BAtU5ZMn65p1JGI/7lyaUAUNYmKi5wuwy8PR5Z3j867vcU3z4tT2belfkT4B
XC/8sxdhnGwgISTy61Sq8JjKYW6UwVJlxHD3spCDzICLUxGbB1EjO6Vr+ra50xZN
lfMzcUwiKEBEN+0W3TWYqfQmEbT6CW77Yr9U8bzZ4CTB6QCSfxfJfQppO4S/bnkg
fXY1KRi+pfSq2G2R/3fJVw5b6Xeze+2tuarSOAA67YZAXy5smWwvJKii607EfrB9
fRBAi9q5s08/fPRXE41inAtrG1gEW0QKi9JUkTr3SobgjRvH5WOb8EP6FBaIlHOZ
Blnt4IT2FT0sYMCP7RoPLzEusoLAwsP1uXcz3p/DUUhMzMCLQpkFhs7UFRe/kOgN
eyIKpF0L27fm+w7Pax6tA+hGbiMOxVMfXAa/l8TQlPL2E/o/WyS0kZEaOa+psjvy
ZkFRylxJMy/CrKE0UD22hbL4aZnlVxggpvKCMLSPzIQkeatQC58/KOav4dUMVQc6
YQsckCbLIMRGuvfTmLzRVswWRL7V7d0copfb3cG210mPpSX1d/H/81OcJIAaq/JA
cgE0BLB2o9hTh7D6E6TIs0DLWHXcRyHurOuJgYX7s5JJDazCDtSv8hEaFUMkXXd7
POZ05GcQ3ynEs2CCXHKjexGxcVGIWaitVwc62vqMHinCtouB0SqO52N3mFENw57r
MPa60Kd4vPDa6pEk7enECAZWOZnOxvfKgy7PP+YVlZioSdZtiaNg03OMcI5IfDld
hA+LwXLmXObnD+iR3cZgvJXAaSwCA3uZQLtOifLW4CSbbnIicIUA5xSthbOkUKMa
dO/xxGTpPsnW9AqLqbF3F0OizN8LPENtu49onnDl2sUX4UCEVBzc9Wt5P3jFGWvr
+1qDWtzjdfb01rQrkuWDtU304NLMH6HMRrEtEUcho+SsXD+w1D/AVy+2K92cv3Zc
0UzuzozUVECsDsPRSbvqzfMfY0vZR7M4Q1pxdCfq1NRiPCprb3X47OfkqYkuQnIM
O+QdeuIIbhTrkXko2ZVJVZF92pOAQv12dnjuX7KPT4sPC+ndOVanA/BejWHlhMDO
RwW+MUqO3UCvvhdnjjjh/T0Bww2zhfp6ogiAXJ2fiFWeCR+f/PYw+QifyqaUJDGu
usCUTZfeaXmf9EwZBE1pbDDSYfFEdbhUuG/xL+3iiyxUYfzcoAKQlzE1J4L2Tt1v
LzHZnqrAzWTxab6K8QLcbTO2k+suvQ0a7RmnUuZDzYyPyXo8a19WnLYCr0nUjMqM
sOmoPmPnrgtvSB4BwoT9yfSiPtTyQaCrEJ0mItaWPVUzuzyzmxKfrkdlzvRqkqBP
ZHvuLljVrnQVIdCh4ihrjcrotv3jz5CKVq3kHKJ4ECdbzZDkTivBgkXjFxqaxSyO
uA8lLRkiYjrqJQ+eJAhnr1d0adUQa7RXD0Xk2Mup2VVqyFL8XtH+fW7uG97gIOtJ
TkdQ5bPbgQ1WE0RbIrEh22Lr1wH+/czEAvSnwyECRYCFMJjPANP2WPP7q7M0RgTa
36zSSHITcev9dwMlqbwtAUI8rYmz4/Rgk7ClNuLSlbiPG/95y1K+z5sybLhMUZT0
5qzUfMKdpv35np76N6DWw4X3dXrf2/kO6k8zd4+1JCgvtzl6meqsd5+ifmOB4D+X
OFn0BklIIXoYCp7BQ7TAxyqz1pacBCa0wQRq7tzDK7YT7atKnXT8ZjlEQz+sY/QP
bQLLYIpuYEJXq4VK30O0bfbJdgPXIuJGdPNCw2Nwxjljz5EklTswzj04H+CUmR2/
POgauvQdFOMaG4IVZhGWhXmJIX7x3C7j6eydT25b2FqUb0LvVtsX5He6IGxx/sFW
D0D4LLSM7fS+lDJptPS0KaJ84LZUnVp3qxoRpImVcm4XCg7GypmHbOzW857fRLaA
MrEysyhzaKcF2dz70yZaANCtISOZp+kscc6tetBdpnx61w0jgSUkb/Y055SJ3CMM
/f+mGVn1njESkVaJFTrlPSnbPumnLc+buTQEufQ4hO+BtWPVbuLwZNzc0ar9nHDh
ECF/ZATOd5oObAE/EeGJy9O+gf++RI5eP4qA+ORVsli7o152RpGOolTVT0+LRBG6
6v9CK8F3XksWAtZPIrCXsyae9MVd4z3d1ujN4d0V02fAUxBp6jib9Nkkak5H55JZ
gZhq/wtiIb+hUvkv5hZ5AtuO5bg/OdPNr/XCbni5w7KBWvAsGa5veOIrBXWqedXr
hX7+cJRxiufRj3fw6kXuZdZVoit1mFYCGB9MBUmYlkJ1uFb6rguK4HihnFY8uUQL
epA1D6G0mQL3f79hh84ApxZ69LqiFAd7EnbkvBliUiBHcnQ2ZrfUulD5eTBuDMTi
/CwtuYqhRBWPDrHUW1eJINBZvXiHi/C4qifh7T7vdt919+OYCJFPsKMDr3t7b0bo
u5gK1sseLEIBryZ/09Dzk+dbppQExFDwoXkqaCamL3U0Rk4ODacDs0tn725Bii5Y
PQN8V53kjL/+9Z3DKN1+ScXtxwPUOiOckr+GvC43rAxW4mP4bnPDZPW6SBmjuPrN
nrPk8Hao3htYkMdLCG/ZoYqw11yjCk9M+dLxBfZJ6T4yxSbrtI6eoEUz77F/Z4t1
LtwqUfzqKV89mMIjN7WZVhfQNAhS6BTcsFFh65Uk1N3HZ9ERtnnFTLpzOPH4nk7F
jFJiOzNGCKerva2x/Jn4b/NYQGwzQ1pf2c6TQ/OBMhIW/IKcrBP0EGGmHNuLhysQ
lO0rA+U8qGgB6P5nxAEFxLXiIIAX4xVgQ0qTGVkZTYdVKHwkjDlzjT+d91xPybRU
neA2G6VhbWc3Ey9nSAvNcO5QCCDu0/Jka0ug2a7cj71lVyGCXFyXBQmBgi8senOY
HK17eP+2xDbouaWckai6yhVsuLlU6WPBwexmX7YnlD1yaCwnZ+755wxRvhA88xlR
77Ny3O88Q41oeda47IfRY6fxYSsiMYY6uOqBBgUy+W4x/sKncvWKt+vijnHvaUur
hYRzinBurKcWjF1yYakWAgEsqld0LikwMgX8sgxv9rAe6KAGXD79xlk2DpK34ayv
R4HwEgcMKJcELCAH8D8lq3VxpYf6q5yS7yjUxBeaW/aSxGriRkJIrGn7dQJZM/zW
8fRP2TU3yKHG8W0wh91fRtoUbQTcH+DYUauNLDaVgti3F5lng2pO697ycNv9edXT
9a4BxqlsqS5DuxjccvtjM4M6umfkab0nmDLxES70rrU+K4bTD8tCBcP9IPQqMjoI
KXmZfxB1Lcca7SK+4cI5sqc5OJRLBmZh6VV/NcC1BlcoW2X3SoBkJ+CZ48GwvuNw
17s/nzAydt1uNOtp9XJCh236qrVTuMnj0UtuHH1BYoLOr0AEqX8SQJ0LKqKNSKgj
IJHPPif7xk0eWKpNvBnkwvgdiWzw+qByuWzGBrEdl+D4KVOKY4MQTchuifQW1vjc
yaGXRdqBWQ8hmeIgSGjKeNzCIo36RFz8e3uy/Xq1su2LJc+30Uvsx6dOD3y4F7ay
S1ZyF2lQDuOVH4Gt3QTg67ewdD/oYXMswvmvl2FbTkwKc0j8l4U0tjz/r+4lqTtN
6Meu2l1OBRr9eq16QCUiGUzhPztwfH8KO9eJQwgnrMYpIRF9Shct4xpmojyWQmEO
12LGJWPdT2k0HjgUIk4m+PgNITL0pl0thupO+lFEQPcSqJykyF3SA3WNNhinKlo6
DJOTLI1+RpayPiIkEagMMOltaoe6+CCVinkBg+JSOI3pHGZA9qSYaixsV0+5H4u0
50qEn2PwPBf0uQsluXNXi2QP33hWprNsiLwCpiIV3Shm8sLStUiFS4Q/vl23FTJV
j5GoY+sJTBkxT50swneohSfT0Qyny/Qj6jtYNkzs4NX0RtAfo/9LcyeFD1l7uC5x
lrH3ZRr7tIhDHP/PjQ5A9dp2OMHn7JX92xEfCSrJB4TLW9VxXiuYYq6wPSHn1muF
s0xol3B6/L8wVKUm9Szf50n+R0RV6JwMbiJlQ3Tpnfc05jbu3sVVVpD5ramHgWi0
pzVm15FYOLFTVJHGOsI0mDPXc/dKy6PP6wms+0G+zA/aVjWst0cdV3ge3imTX+Ct
C4wHHH1tQb1SfeEYgG0LTT1ggyCTqpJzwigU6AOKEyV3ieM/HkOuNDuk1xpDAeHj
/6zY4FSzQqu8jQfW3IH7o1upxioC1hAYrAj60o5Y2ZoHDAJAyPoAI78T76uVGJ69
SV3W57BMNpr94DsfUlhbV4guzK3r9oGwixqQqnZhdRTaYktLrjHPQTekkWFTg+RS
0VGgXVwyatcFQ0ar1Ty2KDSBQZnBriIrzQsh0erWY1crY6BxB0IotxO00wcTExAb
ztMnSufElU7/C8IEsKzCslsvk9xINZ0X3Kb7A/DjZeA5agkvT11xjHF5dFVcgbuT
AF/1vzo9FzpfH0dOgShBDUnyC9jd8s0qPWMj5TcgNF7+uAMMpgfEnWSu8Ji3nGVv
YBuMVcIhNQspL3pJIKgFwYTiSflEbCYHzNW8avGm42Hm0FofM0wxbh4CRrZpkT2D
e1r4I8W/HKgO9xzEsT+2TMGVz2BnZZ1/qgLwRHRxFzIVFxjwNzwKFbnLkSOxNEsX
e5oQuaQxfBJ1nRtkTAFFHXN/E2XVR6rOzhOFdschkKLQEoswpeW39byhz0u1GEVT
azb94WQwQ2gC7JwyEWHr7KY5i1wuwHkEDZHplO7sm6AOFkcAJREuzWvBnDsKSv2s
MbSLPLZN0ha/uusjqLMXHGEwdYlaBGswU9q+rY0IajZOGKhYD2W3qxrpZsbWZq0w
2gLvQpYEdHGJaYVmjxufXaiGn+JlP8PfusDhHa4+tYiUDFgsqJX1vlffDuFw6IwY
l4K2UccIbmrHWQZiXsMScqQQ3p0IkVXBRuYJo5XkonOMX/lMFFNLsZSLEuzBepfy
YIPLJRoBKW1MZhfU6zYWMVTjeWCfla+IomkJAGkx+DPfm4e8cU0Ulv0AFSm2w7rM
i65pRwk83l7wENWrI8ONLUvhtKEr29Lmj86x+NjcjwLnXmxyQKJ18/Fzl/qYkV9X
gKJO9P0QvzPg+ZqYy9aB5smyOqqyQ0X8KNo+XpjZPTuTezO87eoOrLVaOYIsNefJ
0mptsQiK2slElLUnnTKyNIqSOtsS41CYtzYl6wK71wr5VztDFd1alRXbTIHELcLx
jMf6PsVDzqb0JjPol7TPu45n4CUwyCT4oSdpyQY1HI0hTGf0ewyYUareQADB0X5V
lSoeelk7O65wb9SQc8JtJO3+F1p7M+5uLAHg95qmUnV88T7nuOrFyg2f8agbGJNP
e0AXiK91hodAXiXAry1y2GJMJ9X+SutSOu0nlSofAr8WiYx8OCpgT1TiqvDt8kVT
uvyHN3aOoOs8MxB1hWQrzlV+1MkZ6MWpFqHZNavUX07kQVdFNe/QxtT2oR41/6FW
uqyj776kDkVwx5+f4cX74h7FC26HYM/Lft3+qsgPTjJabA8hk7iBhPwXQ48YWo/O
1Z8Z2P6I3oB0Y6yxSLaOQc842bVJ7IJWLHFahDz0XlHmUzEoqVFAJhaVdcvDze8m
7oLCfibHlDTpnWSQXUsUFIxxN5FVeyf/jn4Tyk1NFFaiWo1JD1O99gJpA6CIX0/h
JOSd1qwJRRhel7Ouxp5/avTbSRhBcNcG6bl2ODqP7MD3TmZZ8bH49knewyYylwjb
QOyGlI+0xdc3zpBk9cavzM5DxqQkd8IaDevKwwMRU3/oWwzf2XSfu+IWzQ7yC10w
81gmF2Cid0ALXrKge3eSXH2R5ZXEiue+3y5MMGDeCMfwOuqdmzbouvE9OfbNhSgX
aIFSpVkDrxEpUaGjd7GHtQdAD7fRDoSjZSpx9wycPjEx589DBIA2CjO/Wbm1RKCp
gaRNuoTa/fBq0wM5W8+8aAT9VRGE6zdUreJ5uOHrkGbXYMohDWFm/ufEj78lzCfX
5eL8FwXbxU3dDveP2v97B/65ys+WXMbnprBbmWIgNrs5Cf1EuES5OLCDq7Cfx8un
Zx1sLow9n0cfjOzJfU9psU4Fn+ZUEUl+jKsFe9OCgqanGpNvdR4TkysJGeaAJ6I7
VmqT9yqr09c20+MtE9m93x/JlTmTAd8x302fzM+3RH+/D6nrJpES/cWbuALdc4/r
uXoZjVtAfPWT10Sm0KU9ZcvTQPKFtXUNLcke7m7R9Xm/UyUIW4i7/2i6wjOA147F
jrXs6+tEduJt/JIlRmkGzlRs2dngXTEEsNd+SJ1qNEP8J86WTWY1aYfqfWnxOX2Z
/prxboe+XdN4wIiFl7JZ3A++Tgo0ypSp/KwA2bXBWqT122KJCsj4gKD+vYKnlTjw
KsHbsejstqpXhrlwudEKaQdo/IhdGFpClbVQW/VR1rzh6WtHWReycAkbCvGCx9rE
K2s+3SP3KuuZtLyIlGAZzPz8D57jbB4cDk17qSABfzmklgC7pqJRWEPmnC9paKuC
jYzlHs+b1/5/u7tN1/CXkC9CJstdfA+y8VG6x+jhvMwLVPetOtb0traSVoX/zWqY
S1i9u6LqMgS0/Y4sKtgmnt5l+8tQCxjpOKK40+FnyBMoQnFBrGkvMDIegXyVABpF
cwfCCejPo5ORi2qH1xxm1e/3TcUfXdeGJYfqzPLIAHow4OiMfhz1Sb0jsjvu/Dyk
9pRh3a4h+B+n+Dj3lr4x717PSzoYSXS0zKaBYLCeswBnhM1KHr6EvTSyp12BJY9z
SHPrvRfutjGwWNZlZLjVvarOc2xxZ1kYztUQp18NAjxTZdGz0saCLRwTRE+xNrc9
f8n+0Fx0xA9dsHeUM6XWsymjCMnAZQzKhEvkbB80TYez2Ln1tKnw95pJneDHroH/
X9ojJy5vmlAtmwJr+a+t3jQkAN7S+hAqZ9fyDIBKBAXkeT7wfdUshE3bCWmme6Pu
sw4UdMNCwnTStLOWtPzonpL2KQ7Q5NcmMmLfMAokY01B4X+Gc7ZkDoRGGxBU2d+5
lfCOab0o3/H+gPkf/KNQoLevwoYzT2vClYdzol1nBHNA1Rs8gteKw+BqsPhno7o4
vvkSPXgzZ9CXWaXADC7+nBDNY8UacG6wVxSlJ2wS0XjhDb3MJtQpRmO/FaPVawU5
f0aD+B9nnWGSzwL0IsnIEQ5d/gIy4UyH3xLrFucZT8egy4oh3SQfQvMNalRc0A2t
KQcfL9X/f/yAjLUE3CBdtFu4eDGJSY0c4RQ8z8AWyvG8HW4c1MeUvAx88Y7HHSvC
x6iZIYjMteSVz+KA3kqSY+d65jTC0uTpIVSlEeXDhDviCMofRC/02D2nA1XjRLZH
oNT72ehCF8l7EVyFKYtkEcXfhAZaOW0BfzGphM12nsnQIbvpyosIIyX6inpeOFPO
wc2cUKL5W4M6Mv/Z5fqt6QJ66YIM9VGU7ujQ6xced3yvvuFPPlWajDny2GxGIrYU
xEfm6bEhwpCgwsZi9gY1xg6fJAJkR+Env4h/g3DOnGZnwvetiXWIJd2G/t45OOzQ
0rp0Z07B3Rq3g3hhZD2RD1c8s5C94Kop/u5HJ899wArqI5wFXOkiLngo0+Mg6Sql
kFa2k6AcvlkPi/SXdFNsypTCcgZtyPo8SV60Cnf7s+qda8E5Iv5HPg9wi3QO35RK
Eg6/eoHmu8CNTiaefUSwlOt0+Wo+ZFF5y8GeA83nrrFC/eIo9UdJTZu85pdkIjYA
40tSPOA5S9AUi8C2rQsabdaorfOsHv48qzVdBrI5wqKTEATuVICqoHGNY/NFyEeU
AecEmipVfplIJw97T6An4OCl2d+yX3LYAMpmiVPL6GWLcsKdUg2Yo9Gbw+fzwITQ
xtClNdNND1CYMJg5pBx1xEBVraxr6NpMiFz7oBIn3no6ZJ/pETAU/xyHQTH7Ts1B
4UuPcj620a2U0teVLoxt1UC381RHb4QARDqvfW5EYE/AAylQjRmH0pbk14J4VgOc
COiOzZsaFvgP+G/mQhwx0/ZXnb+xmYGOQjjHhMQnNgAWC1fu4xdEyPKMRJmBwWti
mBohtLsXojzw9Edhu14NhkVRWXJbjlf1JGU7pSFz/alyqnEzengSQ5BnKfcbVJa2
MGPayfk5vt7EvRjcVrs4Fzo2CwMlmtgKAludj/HdBcE05MZb87nenGXQlrR9osNb
xSCIvaRGU37VcIX6imhSAFN3R969dHjoffJ5Ht1Ll6dNqEQB4h3lqrGySBmwJWqL
VM9M+lfpcAsAHVHgnn7zLdrDHVAgpAde15Z9hiPz+p/2ML9SJ7UukMGcsiB5PMaU
Qamp/kjaMZf1e7onaTgpgTe1fjN/09EJKT8uACLad2mKd6iLRpUSjMS/XJotoOy2
zu0JoN6V/sHc2khvjIojPd2TJARfLnYWwVbZP1YItH3QxPHze4tTc9m8dg5yJ2G5
wTnreBwrc9oABjk3fbsachsINGw2pG/8oo2bwOJyArRJa09cd8Oa2xHUEKjYMH6z
4MOwuigdVh8SICY49XTcCjwswl9jhwa6og6EtpoI0hB3f8mnSUviJ3fDFqVOHExo
zsGESSTedekf8fh94/eUiCLjU5trg4u9lxcMjqI1icWx0DtNyP6fjmGX5F8cQzs+
yI/UGdoOLdVYMyTXw5N7M6eNtDly5woQF9fOLcWjgfXBYC0blOSIEcU3+B8PbeSF
VVFEkvvpFoQMm1jdRIZcIY48pA1DBPMPApK+VFf58pQToyWwUS/6mdLaBXwHb20F
MwAmVlupxpYqVW1KIH8y8bF7nNrNTD+fbQ33EVXUiuNzAoJpoNrlMAMj5agDLV/q
6LxGCXy4D4QJ4XiuvzBkecU5aGyrX0jnmHgJan3wiD1kJcpB2qA4N916+F46QBld
xeIzF+EUvFkztUVCSKDZE/c9uTq6/2VSmO88u6fDrtlsR1Q8bbJiZ0hGCdp/xAc0
XxUo/Jq0h4pG6aPweXvTRyut84sk0YSr6+T0ibBkNNftLtjA1ApcxPmwpBV0Ha4Q
xUrku3frO7b3xGHtHBugdmUxnHXfDeiQtZx0voZneqzBqe4SrurJhgkImEAhuVYB
twsPgkIl9tCCM14YviF7J7kMWKD0PyILhcOOgTMt5SJEhwQE85kj1H+WtBfHCyXk
H+3rjNEeEcBiavR7eXjPrdF0osTzrkV0iRrZTM+ihCKJA446Mg0ERLrwsD4NsrDL
Vs/3YDv9SNs9gH4mvzLLxjj7WbopE3NUgpj/f5PZQde4XJTHFoi4v7Umw0RqHXoo
+eSwQYEP1wmcKZtI6vU5rcg7pTol2KtTyr0IvOSbd91CK8/uTWZwIwCb/qGz3R6L
+91yUuxCenE0C5IHwwyIO0ZTD34e8avv2zW6g9Yqcc3WeV0D3pSAjd2PMTo2+eY4
mfl5c0wnCYHtHUrHIPu3cvrLxFjzsYlo0iuEI01Y8gREpwW738qLsBzH0eQyPLL1
XbLD2lCcOcW3LGL74XpfHV3Xnr2zxfqNoitJIrlAHSM5xoYDPSPz1waA2l7Hns6d
CyvXY/rWBqwi7hAwuk0rDRBSZMx3Q8Ilz/zVPUCLhuP/T5+bNyJQzhO92w/Lq7VM
5udqdTGHoUL454sx3tXBGz58QFaKiLWijn0gO6hociOo7yVGpLREZg+t/bDZIY0l
VSpaWDJTiB/xPteNyjVAOmvXUmNeTz5D7bHbpUTkpLNnwRRzHAkVxIwD6/+UiX1Z
BzGfIHFsji5mDcLNQETYLHn4zMTUV6YbdfziQe/EhpJ0LyZtaL2UfEi6uzVkPvLE
8DZyBE8F3OTnx23oXYxWXoOHGe9k/C8ykD6qkJxJQPuIL4RCE6pK0nEr+86imLHs
tslBhHY5m27/WtO3x38+shN9zTc7sVeMeYZaR5SeMguzO/XTCvKBQk5xCdHBo3uD
T9vPR0A4JE6O4WhgYDbrYVWePLuNtYQB3mnVOb0aucnbcQ1QvhwPhRHFZqu1IQ85
xiIl0DHYpOdCDzQBrLk1QnCGo8vywvimK/MfmR1Db3zeeikiTAVcHHBF6vb7T0E1
ME6UOvvJXz5iAU4NE8ppM87nagS01GSalqWlU2dRxh4eN2yekl/tcURArDVakWzk
RtBBq26oV1pbfv0n6wO3Bemwf8DlRBc026G3h6ehWRsceNfKgjLTqLKWHZJ0xWMe
RZZZZIo8iEzhICcYgLmGYmuj9bTOZFDu8iBYrnPfhj5g4a5TivtMf2f+Wq085oxi
LFenyEy6IE9pNBB7pPZsPq27g3VUL0yw3N7qd19BOxByNWgaciIZLdJdvYbdXknb
FC7u9xxSei1nNXkrTAh1Kxp787v53FBCgeTmrjbfczUZpZHRlhlPMIRuLCz7qIxv
KuAGh6x5VGy1zYDLTI2i07Er3jnq+1IPVwKvgB9zAbWQbWOrDh+uul3Vqlxe0Piw
1NWNuzpE4C8JlANviTe1vfeEM+243N3GPxpzPXYbXLFmmcbr3YEHU/uAkJ4ud1vq
JzZywH6PKgGSW6+WoaMOFSbRuU+aKj6YztJPXa6h5TcHYF0z64gqReuuT1zuRp56
iUslTumv2T47qVnKelzOR0xIYQ1A6vQeZhUsRg9NypsQmbc6lqAW+W7MYk/+Q57N
b8XQSjgJ6lnpPpQpdre9a+IsGwxYnidRhJu8simnkaKigkx0K7CHuY0C7LcVA5r1
5pu/BtP0Ep4e8TZFbKkNY1xz6VArhR32ON3DcVz2Q0lOvKg8a/SyVBTXRNBM6Ie2
DNT78MH4SYgJS2dAxI0Z/kgoFGXRCGSupHAmQQMCASukS3tKC95T//FJ8KYgbVR2
QuKWIBcD8f2fk0N5y0kPZuf/DM/EnA//5KV7/eJYywo1OPYzqvyo5TACFysakK4Q
CIsxIYnt/NfmxGeIRByOijBBSaY2ZexNV1CU6Cqq66pOq/l35y9K6vVts2aOOICm
KsMbwI9+e5Rc1L3oC36XHbvqGG2YJgwS58uK7AJWmICafl+s3u3To8xa64xc3D2Q
hPcV8ewVWz0rdUr5GRS4+lVAhMGCigKOz7lVqbzS3kXbpxqAGSlnEBBtgVpkhpSS
72gHcG4TTrz+7X93alc9Fbty6zvhVkKAp6qT7BFL9fDC98zyUfyYDx2Un1SFWh5C
G/43tlWV/ZIggKct1ajYskEbWE3ka0ReGG0HBu5VOqXEu0rmBSlx6kaS1UOuPrvA
b1f6pDsOpuunf57aBVbzBBLQJII1egVUWMCiIMx7bWQjTqDlne0bFD07XetyYRyT
Rz6pFT/J1IOUT90jfxJVIozY7kA6Ca4JvhBavNOX/CCkEUYPX6scpoKoTlQnV7JX
66iSBycnZkq9vBS3y3t5ZOce3+uqYz65dXDeBsI0rGBG5RVLdMkCB8FskVTzGA0n
RZRQqHBc4umE+lhc0HwWa3Yiq1PRZQOmWg3ZKhl79k8I1wVHJcA+4s1d9j95vWJG
s3LhxtslmuijZHci/uFHvEOVq6ZAsC9yejdfvgQhGonXAqgNRz6IvNj6bMECis0X
bmzooweeOmS/xy3phc0T92N99tRewpwR5gt+lhFdIndYSkkqKzBjlUusMWaySY6R
ugnUBgkmzS8eWd2nu0F46iZEZ3XK2/OYPaHNpf/2KI8VHmEz4FJo1Ygcq4fNs2c6
AfQ75WkD3VjYNOV+U0SdI8qIcR2ixBEetj4dxISmcXVfhCquO2MMXZBM44sgbmAZ
KCfK4TG2zqMXv7AoZMiPeK98PSbb/CkypuPGf3StBH64rZY6Hj7f481NHehDH85n
JQXB6MTcM+YRUMN99+4R8EJ8bfusDxm+6gcYPgfjZCebYYhnrJEpiImgOPVpDOWf
/hRH5YN/225APBZ8hXqVYkVKKyTHJamOsa1owADW02lV23QJ2/z58GtIxKK5ccI5
3L1uCDGKkUeSUI7LW9FArT4BaBlduG6yiAXRkkt/r1IV+w5XX15qCHJw6EthLYXH
G6gfG0ZPAF1BaekBZxxAnBApQiW057oFIqnw4BSZjtw3HEuPlFu6U9TM71v9xF2n
VRXFU692mCrSm9xbcuurOJ8kVzB1Tc/+IQ9ZLVhnrTxr3dYL8M/+2ogyhuiNCPLk
tJHBDE3bu6mQuKWk1HW0I1EtE8G0/ymjf6afzAYtSnygqBl8qYzWILMf61amMK7z
EGnz/poWBlY7otJAulDJfIaD2Ry1BfR37PSMQSCoetUcaKGkDX6B6smxFX/EndIH
0h8u7N66EMMTtkerfLvyeSVuw3gpNTYWp4XnMcRQSlocLuDH1inVKi+EpHUrCusd
wr7gwAqca5qwk2B2Ax+NSCKs/r2T+amnhwPTNsBwaykTt3IDTg/QCbmoCwB807u8
o0F+P+xnmnkQoyaUdq/g3978Mi2PHK7x94Dqmsw+JfbA6OPrWy7Oe+gbjteWSOJv
Zo7j28Qkaixi6wgXQDvgzICwR1sfktwTewEqlrcJnNOqpv+hOpgEmQCCEoA6uaue
plpRV2Pr5VzvfpECWy+39ywu6YBxQno9MAaXEUcOQ3GIpuPw/H6okQHS6P3uIGS6
4xnqy2BNg5DyDKVX5UDUIT9nUaxiKG85w4b2vHBkjnuIeenUH/D+JKx7jfyL9B7g
hUYFlAVWDj2Nz6xKnjuL5L4DNtut/sJH6NCqXa4PC5dT3PK6oJOaz1k33OGkPms1
7WEv6U7r6X5cn37P/dG6Wqv058Fneg9MfIhT7uVtEicfoRrIhP7oFgFCTq4Ml8wn
Tt6+smZBDk4epBNEQGw2fOe5E1eeazGmCzpWeBqtN0jPVEVsGoHn5tnD3WjioADZ
6AZH3hG1N066qpj2FqkFCTr7eXc9cXhuuCZlnKvySOAWbnV0cUoBPPBV/DFtxqpo
B3cjY6YJ9g75K3X715N0IWj7b4/FR1i5uGA4EJ78evYS/iqZEdCoJ75AgN+MAOPq
RdMmGKGynbbJUk3a9mCfmxS6eAD466DC/2gzMibKDxUA5sMiq5wT4BvmnbPGq32s
7wxy6pvEK9i2ATo0/L/CMQ630/Sc2JjyabhDBF2/3oNnJBV/KtqxHYYnlPz9jg5n
99FspohIkkCUYwQqHexRVLQYxj0MVAoJM7u1B8Kc3+5GsSfaYc0iQPh+5BTRTD2g
KoCIrUeH8b2bd0GessUz2itwJtpJewRqmyGIX4s02KTOGbK08moUse231SYubbQ9
O+RH41i87jmVRZWmq3uagYzAHR22XlW6NZLVNKnUDl1Q79n61X+21nCmYo/4ML1d
KCZqxDBeJKsv/tYIjX47WVkfMscXWuI6gZIVOxz9eq2DKXPOa4OjRgGTXSEbo9Mn
9L39VOcQszvtCAE15uVEaW/NjJ8Jpi97kokLP8RVDoWFA+Yi/pk9ovghrsgB37QZ
+mjGDPx3URs/ZhjuUtKDVmYHdg5zpzbHVXkA7LvCrnDhnukVaaKFHZWLcIsqZoxA
YADpnBp1ztcfe9KKqA/nxt+ubQhb0twpQP9eXJG6/1CWwDn8B3LrnDiVerUjdiEf
+v7IgFmNTDExTCeJTSIY5KJVkodNZkElUNALzDgoB/nPINngZGHYnU2scswP89SQ
Ul1xa71H+xoD7w+WDcQggqDSupR0jexzY1Lzw3jVBABcnBJu+ud66JaTgiapNaZ2
4VSBuCrbDxHM6BxEo/HQQaChTA3k2LJqT0tBSycBqSVv6E2OKXyOzmnNZJyn8y7E
59MpK3Un3zVuUG4OPrvBhdBtG1YBfkaUjvQm3XKZm5IACOehE/EACuSwp+T2vnsC
ZB3pjyP+0si+EOjvlSUjb1UoWbiwIqRa4/p40OQdQf4XFyIET54e5+b4qnyJEGj+
iNrH+cU3u6UItls4oxyhkuyqIF9GPJyBBPsBB5NhNfuIxlcbWLWC8uHo2HRftISn
C6kTazJDNo9wNEe8Y3Fp+DGJeXPnu1KLVazOgZyvWHdz80V0+IJS0ZaxnWNFcDwj
KFkU+dvJ7z6eY68PcGKHLeC8eE90Gg4R40pk2TvjqE2B50wZW63HaScyrgMW238F
9Z8Oa0/4itj59qVd798xG5c6GY0GtMeNmS2yJ0Mv61rggMt9VkDi6h7iPmg0YfwA
fEjULDqdG4fJo9jyzUuJ5k2AOdaTiCyeN3+lWib/K1rUbhvBbVRFd7lhIXbGAO9v
O0f6T92R7QDBeIcpWgmUCZCkk2on8YRMaOFbEJM/Rr/tpu/h2qebz2632s7w35/W
Rxd3gJtknek/Rz5RP3i+gwObqX9zrD/USh/910eIK3/DC1aCseCFuz5ZiEenYgx9
RywYoiapUIRIANxRtxwYeVtP5iC1H9AxOGoTgjep3NCAXF/W/cumKR2Msm7I4EmV
fnnMR9KTRZrRGsx3UD/IOffrHstIZJchpY3I5sIG5aR9iuUySiuk3E7IZp5wrAdM
n3Ubf2r0L+DxSUgIcQ6tmYiwnRcLnf+BcTORqX0qj96lVHJLnidPHbt+ni3LUQ42
GbrpPw/qotGcdMLmMUMSCzIDp/fS9g+jwo3MK8wOqlYF7ziCJ3Mme0dUPmF0lrQu
CDx2CPS2GxvDdW4wJVJFUzdzP3T9gkXhwAcDIkQof1OGhlDkpcDw+ukZKzTFzYxm
Ulnyb9/Cbo+kcVmPRrq0sVRnZMf6TAMJBcmYvRQ8aXk0QZ0L9R0ZChVzE+gKDO4A
M8S92lencKNodlFgwilq4RymywZ6elaMB7jBnze5VpWtvSLvBCqvqDA7gHM+XQFW
BmKMTDSjoLBv62L1+gg3+XhZGSXUS6PaVDE1WnUykCDHQ1kPh6XnV12AgMCN75/8
wHFpvhPtl4G+zK89oA0A+Ag5iOkSjJLH0ROvl3w5AW/QdQJbSaJTIJ81mKqrkNML
1w54+uAi1FSXV+iQPZymA38xkWRMlUz31QYG3dX+x32tmzhunEMdJnEmvlWbWO0W
ar2teZrmy0aB5Tei8b9H7QaocthtgKGz4ZwF9X+OF4gt3d1/H1hW+drVb18S6hiy
XlRImqU4O23eFBGKT4xL2wyTO/v0rCC8H3C3GwcAD+i36nx+YYBAMwgLOkVFMc+J
oPAHtcUKeGatWqOSLuInUalQPeFgH2lMlSyZRmQyXCdxA3yqOCdpUkLO+YcPsMiQ
TXdpIvjGNP2nw165ej8rdNLH3NI+Ki7FxR4t1g1utpKqArgKk9vPLjzZaIKo51fU
kBEMGDB/h+uAJDSfF/+LBd986vW4ylrGyU1LNhitVSBXyWcRgLH4w4198c8HiHoM
+8OhDP4icP94gIWu3212XuHlNi9VkY0sKpjRT0QbZbyIxKX3fn4Oc57yUimJnlCu
PlPQ+AoM8LcUbd9QteX+8YT59bnYLAW8Q6YGR3Dc44JlKr8b0vdhQ0TAok9hLyBb
hsEcNglhs9CrBxqs6i7nF7UVd5Na2ckKd6PHE4G9eMrmcrWcb6k2HGW/xtiFOg6W
jxzDkb16aBmdehNsaIIF+o78quDuJvWupLsVb0DXQO1wPSRnCAIkeYhacw5455uL
ae18o5DDXw3uPRcB6gagfVRAM2LIhjaeYb1QA911eXZV0StEgyB5A+S8yt/WbpuS
1f6xaINouVTdSmqg/ETUAnVSmMzIsvngVV5JHIzSQOmbKdwDrRubDzxdjHscFm/G
p3mpGoP3S926B1I3X+6+1DBbuZaLZqu1d1WN6hXqZG9YSzhLm92ufQyps+F9Ifbq
NQiOaqH3Qbl7NBDhwgFL/kDogDWtZjWizMHzSxx9iZ4vNlQyRSrOu5YMoCsu5F+e
cbotLjX80PPDglizBv88mlrvP83rOqvPYHf0AJTTrGdScsDs9IXEAomwxS9P8+XA
4Y6z81GlqxGJBn/WJm17kwPSjloABriR9SuoPTXs7+4m3/XECaF4+rF9lqxK0Wus
lUZfT0dCByyR3jMJEnTPohdh/7sUYtS1KGU3trh4ie+xCNf3KicI2XANzfipkT4u
P4Z/C8b4CmWIe98jwXET4nr4n4wOzOt+NALWfobfxeA7BGcctMJsiv1ZH6Cu9kvC
SvHgqqYeI11baeapShDezUhgqmzkOU0jzZCBxaBYGQtvao584Mlv8ZI9M0oQgP1v
vxAsBdVR3LFXDgrxeUGtT+Y0QrCHm2JZHp0SyKnaGBatrq78am8NUH8j7pcbq5rQ
+gR5AqL3oe5qxQjVsl8CMub1jiJjHQNDP9Flx4L2wE1U/tbTpmoRFtDYt6zjPNXy
2l7h7uJNCFqN8/2Co7W7Qz8GWShFF8QA0pMJIHgTDdAunG/MItCdLdM950cuxffX
ZqF82BwgiHzhevYcTr5N10CrKQHpd5R3Yz4ZoPwsZVPBlvvgFIaSfJNvPbk8wcLO
/Nfp/KmI2x9J6J3AIFJT0N+Dbqv6EIRNKwn37U+goBS+zlwWL0c3ZPtWj7aOQ1kD
e96Ml30ou/FEN/e9aj+Kfd+xXWOkGbG38XKDMAUFwDSsBcVl76jwXVrMgNWtGmA4
GRae2NBWgHNPoM/oyhj685rPchd9sud8ArS685rH9FLbys2MUtzKqVVUMn59R3Hp
JvWGG1xjFwFUBKj05+JOOSPUJLBkJgiKIeUa+owUrWuVsAH+aUkjeITodkn5PAFk
wj6gbC3hs6q+gN/eEIidlGfO4H5lRvF7YOJmaIS/KzTQzqgvgA5RConYsO+f21s2
F2+awuSpz7goOgV9/I8pul72MvYHFRx/fcRAQqCX8yhjfPvays10Ybl6GLlSNgm0
PyKXhBB72e2bm1HsEMJY3gXdsofZ22af1tAC72jQnxiuJAe6wZL3D06KrNjYVVmR
hjScu1yKU6MbCxRN8oGDRwLHYFZlJ+H0btuau6kcnOeA/zdHwDyK935ZyjMlc/S6
C2dIUZfM8KVAK06DQ5xISAfGYp4EQ23K1NbntVExNtekf4/DR2tltcEeMP8/6juZ
jQGWdF9DymqpLv1Uwtx8uWbwOhmLHZqc+o+L0XjSSVudvqIAoBlhbwB+HTwlVx+t
12UGNAesqndiSvulcn5F9xVImB3fTFbP0+amqpG+j29DH/fnUXGorStrrYaBVID4
0H1V7fXs6+74wo7K3oZiORICHflDhBQttQipVXlhqHyqfZUQ0Zhx+ssbLoEFmMQI
K7U4KUrCzGv5YEqzxiUIpQEoJB/x4eeJvBNlOKUKwScrQm8qszmBW1subMiPw63X
ILe6kTolKRdIjP8VjtYe9JejEdDXpXk4U/O1kQJjjEFQw9+AT/HC4MGFyzrxjXMs
qZC5OIaeq3PNloVhn5VTImgaavPcUeK1SQ6Ockh+YzJfP0WlLw1Zn5nZrnhgPNZE
4ldCXyxGc+VZ8G+zZYajcHnJ7/PbF+ZHGSRKOkyuy7WBofr9pBOj2/UR2MZbppvw
21FpUpQmRHf7Zhd5hBhzwtPRzuw32ZqMHoJxtx7gBCrDuVzx88mobg+L4Ba+fC/R
yqI7ah7ISKd9fVr8sprx6GNp/PaqX3rSWfTrDVy1gnLfzfZMcjaOMdhAxeeCaG3e
Tz+0EMH11hDOnXLn8WJVm2xb3peKxr9Hn3N0RqZSUHilRITEYxFlAdYNBeInxHAx
RXH2Hd33ujBwOj6b7igIQfd3xMlOKkxMtiGLz3Km7+OZnxnIP62mMQqkBwz2W0ur
HWCxeSUjeUAPTCawMeAJm2MZhKSdLkSaGwc72h0ESuOjNlAl69xXASff8pTtpWF1
CVOKgP4AkoeLzeRdjE1i7utPewvJDGetxU8zRaZuqRhGrjpUzRqsNkQx2bMoQ6DB
XKNFrENJj+ra/leOUtSjgWa/IIDDuLDaP81XNkBbI1mLpgmPTD1l4S1dilZ/VJeU
uLttSvTjbXW8Yz8lfM9yQkIJ0G3G9zqVUJkvpJwA5yk4qqmoDf497LHI2fsLmWg3
QSdLEGye/M7ycfrPxmqRakPdmbCy/0j+FvYJNjwCvBdhpaUj/+ApqwzgUmisxv9b
cRl10qZgbiJTeKNzTGPjNVm1PApc4tqPHhgZJ1XkWpupr0Wk09zQzWgO638afnUH
jwC+l2zzZ9m2QW3UOEJYm4G01gqj0gIa1JvSUQOs/L4U2OKrjtr2TNDtFOpgmfaw
H3Cj9ndA+D4G+kRk1Lj3YS76SG/d8waZymTQppHtReMK4bSg6ovPkZleW8QKZqWb
alNCvu7IER7xZ5kqL4PSNQ97mXtGYx/+vBKzgT34UIoWkfWwf8s7u3b96YcCTx01
POMPnsnDCgagiMvMPXHZDBIoemRF3qvahrOCO1PUQMo8WrFyDrZW41wf0nBbqJXX
8R4xvLDP4az7w7yQ7I5ozrpwWLHC5GMf57icSdN6qynTwa9zI3A9rSZJu5WFGCFt
owCEpWKl8yw8ativOdWYccdOx1WQSVAtEo3yx6fiozrM0aH+jwjVYne3Rr4Fkynf
a4EBUgF/7L9S5C9dtVJJKiVcDY2lJ1OCzsX7hB2bOS9PZ6r8YuKRWC/fOQUeBsDY
2HKeEx64uUkwXBJdVLUh5prQNfiSVPzgumKnkovKIwInBXNLFq5xgSseDZiH8eao
51cKTRf7tTkD/FMc8B3UubndVHWO1frTRssWY8hpH1s/xlquc8jfe6SqbJ+OeZIR
m1kUXPcA8EqaakMhyg77aTSbGM0Z0NE1yC8ER04kSzX1ZBs5LBbsF6bC2a9h/61s
oEvHW6rfnFDME8M78fuwIzpxwR1WAy0VYbXBpMyZKwjb6FuS4Wo0BcG/OHT231rR
dmAigNr++WfRJccX00vffvO/1uWeVMRSsO6sZu0AGHrExeXUdmwOL+gD3/o+cpEq
c4wGhcyuWTajJk1G4KGKyPpEal5/30ztQVTnQAZMLE7YSmy913BoIe3z+IgmyDDi
uAfjiluZTCrIpV+0Czqif5MHr5GJ2tzbRLQ9vVkUc2Sa6mq+/inhFIYGFSi/8LIA
i2BaUT74X/8SM6hGoQFoqwZZy95NdbdVA5vaZefx+ae2T/V8OVG/APXWY3OzkjL5
yqrCkImcuSXNEbeHe7I2Wyi/TZNAaEhETQvQa/bCCtqkcynh6wE3i/WduJIVHyhI
nzyVoEADd6r+K5Op+xS5MtFFC0hUPPSmI10DI5G7Ihnlah72XyQi9IsImAgh029g
F0gdDG+IQ520YBbnbkjJjMVKiS1mfq33bIDyc53WvLfwi6vBNbNz7MLhnWhjV/EQ
mvGNmnTNpvppmoqey2XIlJHMGm5mixN505FtlRfrnQngOb+mmV0K3WFNqx2NM8HO
V1zeQvtLNZeumXuZ/k3kh9s1zhiwl+8NuKwtbQdQ8YTo7sG+1pAafVvgoNFK1x7h
iqlnTw+CL8GTHBmo0ZrTzZsqJ7XOQXvUv7DxJAaPN7ucHLbeUrLtJ013nxN1OOAJ
ic1iQQK/RxOoxj3BILxT12SG1AntyYr8llAQtD/exqrJ3qDs3lSH6G6s2VMNOGxk
9/W6OJcaDI/tDWwZ5Tp2+rHRnsAbypSfFfIoYgbW3TLMIp+rQ2l6pAxNziU4987d
C13a9M1DpKTnsqEPeL6m0HmXxAYyksocXbQ1Uw3w467EFP4rXYW2NZhRuV3XliWR
WuykxtZTp8HIguwJSN5AQxCPAV15KBez6f082X+V7YFKcoIp8sBGaXAduE67vFew
V5SQclNz/Wa9Agx5WmChJjfR/kE4Z79fhH3dz5PLipHQGEGTtG9ET/RwOTaLzMhq
gEeNkOppah1YyZx1WXv2GsXiK2GU4ml9JTv+nH6aRQjUHG/Aa5mbkoWXBngxqdrF
OhoTIhjRgIcQ/nG3xP3qtVpLJnTzWHTN24HRi75z1uaEnKwu5Omp6ylhlCppZJyu
QFIDC/JYu4Mrn/YCK2gtYNVoLyFiHab7fw1UuyWowLi1mTvvD/FyUaxRmDH4cjzr
bnyYHcIpoYaQFeekJN/93AM+Go82eaFs1k5Q9JwJOHyk9psvtp4bGuIb60pyCRM1
VPZr/2Sz0lxMLrtOFYYU6140cXk4uR3cDNnJAfhMSB8hzz/dd/ji8S3NGIApIKHg
QipVvEj1g/SeC19IjscZBOwt1WiaR3qL3/Y/tuty8bB0K9RFrYPKzYJQPuBVX99Y
woqJx/W/4TDPRBfc0XGXTOzt2Fvm3fb6lZRzN66bTT1MtZLFAuTeC+R/0lyyKjKt
rGGWV29JmvfdPMuABFxEwTxqhGa3sbBe3e28K2Qsgtko/yYTlgPfEhEYN2/+tjiG
GKMSCdI8goP+eEdDQM47Ywvx8ZPf+LCkZjIYKjp+pvRu4Jcm4QsrtSd8JTilvXc1
WslE7j4QDpKa34a7U06GUa8H5XOhjmuEKgMMPHCCFmOEla4fidbCtjn+P78UMGmO
E7HvXEhlvQn/0hlPejlfTlp7D7pvm9OIWqlySAYo12Tz6erNOfYuMY6xmO1gbs/k
0ZMvjjQUgsT5UwDeV9DyUPX8kPMaSaoVXqUWAlamnkJSCSzbyMHacEuT67YnXQBN
ts8AvNN6jZh39/niZUN6WrapLPRkL7/m8w5Zv0tdGgv4ZgV6/mI6mugupdpj5AhP
pKfR2079mIwIDZ9w8IE/E2G+7guTfw0S/zznD+loOVvHA+iJJkC3pgLAl3vxTmVl
Di8hWczZ0jSgsr4/+1rhMY+aerJcDhyVMZmjirauq7JVWww5yGVYEJsX7pLBZxXE
kbjp/pGrm92S0soUm5YJWpyv0MnO/AlD1OAPkYd44y27ZftCPQzagv6Ou5If9fyB
Yy5Eg8RWtrd+wJdxxzWoke4AcoKarHZuC/OKSEo3iu+tEcTIhS/lYJBpWvdnu3Mf
30uwdLr5rhewjIwmvcyMBwxIud8NmeZ2TEnj+4Fbh3vMMAIi1dugXyuqxbwqIt8m
XlAZssIGmpVC7e1o0ro2hPAzSUyR9qjfrZvLJm7lT7Ob9ldnMS39gC3lrePT4ht7
mee/krmx/qkzllNySJhPtjwsZByytXMJXBzlIKvOUpHU34PrH6DoaOh2fxkFh/06
rofzL3z5RL1iGG8Yf4PaTTmIhoitR4NF43M3UyO23QuIFl9P8MibWTuKwj4yrvXK
JOpfkhRHLuAl3Z3wNM0VF1MGLFTtd8ZEMWtBogxXlM9QkyYKm3LT7jwj2a6VVt1p
THIY4iiq0i1hPDVUpGwRLDE/6BP0BRG2va9lk+3dZaDh209et+/2pB2hvsJzfeiu
BO2QXGZHEoFREULhf9cprtkG9rq0r909IxWepmx2pSG6KyyF2040NmsyF9aTotdU
y9qf20tP0rLKBk+5nmMldMwj+pw16endnfDXwTwRdEPheeuQ1G0iYgJkROuaMIt3
74tli7zB0+Yat0D9MTP8gFHdwN1Nlwuw22+jcD9rZArtsffIiT5fA9woR6ytXui5
PWSuDSxqUeB60scE3krUP0XSomDJAezSGmIATI9+mBAp/Ywx+MejqqNRD9thVcjB
BVmqK7GU90irvlGOqNDKu1buXT+8AEuarWud0O341f70qUFUeKXzHtaE3HHr3iVT
OELHaiU36DDvswS49gww2tB6bAzsZr/qC0mzn12Z6TOHu+LdHo/uwisuxSh/QBRl
igoicYdZd6D/uKhALrFtYrxB+zKJe6IN4Eyj0zMeqF5xsG1+er3yZUhbdBmWeTeq
v5l1TfMtKgWELinLhN00Fi0V+MqDZFaBfJGxf/l/D5FE86GcAIjt0xkpZjsniPRL
PORTwsS6mnFbu+veP+JcWdvMd33Z6NvFUccanKp37KFM/0Ogd2U8dNpWf+o/wXo+
fGNtl6JBiQoMtQ9fJijsGG7h4GdiKpzqwXpVkvHffcL7QlxrKP9aBL0LN5tnOe/Q
Ci1tujvi+/06Cp4Gsmx7Lce7k1VdN1ZyTbsQDE9M5g510Xb4KYoZHlnXpsYbJeE2
t57V5vLoJpvOqjmoa4GKKZFuMGI5UL266f1I9TaRXfWfQXjvJmQgBeCuh56JoJ6B
e9qBtkE0mrvAQk4prWFcqmNm0nI8hK9o9v4XeAR449Sk2JrEnQvDO3JVkvuImKNq
0CAc0U4ndOb+e2BIF35YVn20EHd7yIZ0rs5MOcfkkmQfwZocLJOdpjaqza20EvJy
+eKc932c2HB+dE9mTbuSeCwDJzCwkpqDuWkMnFVhEcevd+OmgKxZxNvvk7mFIkgT
lGIW6UftgXHKM5sTIzl3xgL+kmi9QupY2nXDl/5F27jAOZ2JJAF7LO8KccW4s9iv
ZfQidCgOoUMVqV3QVjOdDHBFJyIo9+wne9xH6hs59Z4M7qFy1WQPGVtl2fkPBG70
GC1u50lnD28UMNOUmkauM6WqUAxY20rzvAZyNrBEWMmklmlDiSwQiWnpxTPvl9LQ
OIbZqbZweeKqXsyx86HZ11efU5v0MfUZRs5e80PZc8WDq+xuFpg7XFixmLvJMf1+
b2GVjyBtTm9pck+K3shKRFx93okSYU+oEGodCWdT4dNTNCDFk3u3zFb+2O+l/Ab+
VIZtzrbe9gVp9Komztq8lfVICCr+6DuWb6Yff/P4Hp+yqfZMzzhMwA1NvWpETwXz
EBeEi9lnOEJCwHG2K9bL7zKNKVMYL8XH3r0mDCjGkyudaVnr+kJ9IDu6PYebf8D+
dJSmziStI5vontL87zjI//lzC46djmP4L5Z2o58v2MlG6UxmVcKxUywS1UYDbbxn
beH4ZgfzTmEJ4JT//bP5PiswWLXQCVDfUqGchXkbqYwHQEdAufoLUQPQrYzXCH+M
GY2KSRX3+Ss4K38QtjpoA7gLKkdZlkgTaLNIj5upRtNBC3CZy+OZrhZoUb0leEZO
J7z/6T4JYgyjrurRvrB700WZjWY90kXQbjMBHnnxL40qqSHZv0QXeW3pkTriQYFq
6FOz3aN4jwsnh2OJifSiRnZSMEfy3jY0+1hpQgvquRqMD9QVmmEgMGs2CflSqr72
/bvoHdEGZ4v8fMndIvLm6VR4pFQ7/kJBAxFi1M9EkIgKxTKhSVXVrlPeU25P3rSm
h1T2tZvNf0xra9Ap7+Z90V1J4I8mNF8EhzhYfU281BxKY4GHTGrAbRFNNYVNfMat
WyhnPDxJ6TSZ2MNJIuQ3QsngYcqbZyZzjMJb3/7xgfBMDgqQ4x+80uzeQxM079VJ
ApB5mLNyOpT36GNp5Z6U1bc2aQjZIoKSqQEYpTYN+tg2HLp1O2h3eoFplTU+tVel
t2OHUYTQOCEHXcRBc5BuO1fJAAjbxiXhY9DPl+Hbm7QjZZmOUGxu3iu/2/XzFLeW
JfrHOz+PIFTIc25WDH+17je8hJCBcM0eB2dMPX2xmJENw/QnQYivs6gcWU4G2hih
NeWLCHLxen7JKKbGXWGnt9ygtY0THpSQzKf/Jh8++JTVWo/amn134NKyOD6Ty4G6
GRmxKw3pzGwbRDN8JVbIfybae2rnE4aP+GrNg0VfKWwqMsWPU5j90YffQZ5Ont2E
UoOPoDCAJ/RiIKrsSt0En2k5ssLapFjVQfKGof83N5ENUA/E9XuBi2QKtCYXC1ac
V3rA68KwG+mTJVPvzcORYcZqaGnstGJ6vCIs17e2AzhntwijN4n3WBnP6XXdtX7y
TcRmc95NcPK/ERrXRwids2Zjfnuh05bi+QfbwXjI/RvcTxynsampgH0H4EZNZ7FL
n4D9aJivgNuw2v/UkFVD9LFjwVPWSgb8dNLzS7l+9gueWKFv6bekah6ajV/OBWfY
6xaUfrZXbZ9UR/uHEr5/EpsrF9ne8pM0BjNOJAsRaBH6uorWNeQWqtJogYCQ5/uT
KztjvT+DTuHf5ruS5sDsvsuOKpMOCE+Zll03IhOPKR5xc+eFZ/H+hWHcueunNmpV
68L3DqvrrzK20zHSb3yMMlqt1jvjWHUQRnLNFLxDp42s7mZ1rtph1E3FASGEIw58
FO7ptqun0kwGOO0whLDsck1y5D2iE6Lrvf8BE7AWiLEHB5VXRUD1oSL/cKXOBuMm
1iknVFrpyG0uH0LHpxie/c2YXFxjQ4Fj16yzfBSQHWDrJxmQuabKreddH/AR0iiR
bYY0rioyKwhufag4hiBSeKl/LVoZZto3OvvegxUwaDmTifiWLT4hFsJg6Y6aO4lC
zWC6Z4EhmnWLXLgV2xGHb/S6i0xEX+odtbGQJXhlmPusMN1LL4TFu+wl4Waluabe
aCITDhRg8LT3WcKedTdekCnhTjjxiVjEFKCWMvnGiESKhDjRlPmCAFD56kdvPxCY
oGaXzkjDk4oWAcLvyBy8OSvBHtDCteddYsaXmy+5bs2CEhF66B2KtsKadrl1U7dM
b6qItWsIkFJNp9/iIQZcexnR+Zde3mN6FrmA0TWplpMFOPjPb0OoioPrqwTp9NtB
JrEcXHMLe5pUzvZVvroSWybxyw2qyDwZ1Gz3W/pCfYoAu4u4Hr0m6Xjh2EKGimnL
Ae6ItmwsmMcrjT0UdmdIW+ml7L9sYc8n8q3B30kHHWrQKND7KCEvJ6Tsocw4CqD/
86mg8tUkMWy7yu1IyplSULl+IAc56VIxuO2nGnJdoeHfn0fjB1GGJTV2H2DdiiXq
LoWKq1032LcCqoGWPUzfz17av5pnECyYYz4aB+kONLFjcyg6LiXt3iBx6C3vnVFC
RAyndxcZqdZ3SzyZLBSQ91wMxDJrWcA7BBZh1QfGTzm+hdTI3NiZwzLWuhO9ef4C
GlrI9K1rMQXSPVdntpGBu+Ys3GU5cgq6z2LEJvcrPuyQdyfmgUmGL4+Vi8IwCnwV
5WvP5fHL3Sqk+B56MkCnzHWrf3VN4DGAOVFGJ9yoSnVF5r7iX7pA0fJ4FFgVeS0S
cobRSQcbA3EVsc8pvHQKRXN69gg88cGUDdVvT2vXSY3SFGJudqWRCpCsvsGlQzPH
kFX62QPsuHqzE0W4r8ZkLSODLrteE3qNlkTonQnDDo7rXhQisj/fwPhChm8DRUTz
e041YibrQi4VBY9Jk67beFUCTVx2JtUD/DGe3kKjNr40Bi+cLTBYIZstpEFbfv3A
kPCbBQAmzq9xoPQ+/C7vKd2h/ymCEAzRjSj8AwhD0Xrh867ZZE5lsmHpzdOggQpR
IzOHb8/lBMQa+ThmnMtO0Gr+urwR/3hZ51ukuP3dLnTh93vJcsE37zH5CTYp2cCf
HEjUWr7YSg56ocNFT7j1TWA5DMOtcE6/6sn7e3UgagVU43l/xsoNoYxtxDWkKC5q
nG6OJyfW7v/KCwbxXGFkh4UcdsvJ5SE71jRTEThk02V4Z36QBdIrJ62BCsEviMm1
kWM9cQi06g3UkLUYFeNe5QbDi6Vm1szWgMWmuAciAgac4GXIOugbMc7r1pkmIDg7
RzzmjsEG/sgo3spKnu+e719khmqmlGo0v0eIQ8YmZn5ofQcTFzFG+sjaEBeh1GAB
2cFHv4DYtVYxVrjJyqKvVZrS9O6U95BA5sBgtbS4rOEZKcYEG8dl9/lqU7dHvZKN
whh0ikqxSk8Lc/a8pghtiLCVZA5JC4mI619A1rNqIz/RwqDTVIAzgDsEQaGXzhCq
xWb7xsjy63DCGKar+yZDB5dDt8/Bs7cLxpGFwcSu6nn9QabZnkfK9xzZ5L0YDV0V
e0A0O7SlkTeaXBq1YmdWtjat1HhA49IpzSzs1FzTitY0SmPHrddpSQQGYFuhtp4a
rBGGj4DZDftqgUkmkcuuopU/ZoQQfbNZMLGbZl1FazZqVzZ4MALfhD0YFpHzt1Ym
m2CaDuR3yA0cD9hb4V7521efVtz6uky/Tf/4/sdBvciIHzSxrvdRGaFVLp/zmiYP
RPWLCAn8ACjkNH0nRjhT2oxo1pFoKzCGGnIzqqdqcgVpBoMRXjgR6qMsgXVtweKR
xUeDOh/mK/czlRwE28ufr9dONmZWFNhfHX0vmOdU3it0y2LckHf9OlEY4u/41CAW
Xxvd/5Kiq9xefe8X4Rm9UfZycRB4x7nhP9XiY617D3br5ydNYlN8D3GDJsfGnN2K
bKKqQB49dX9RBWdNRx9qyjIidWNf/OaRpUpfJ+H38dM43/GBuNo3xRBl78Yev/Qp
OxUUfwfnhQDO8cwRfHgbgpzZh/XpyDCbm5t8n2L/Eie1+zWsCKJnAndMkfLMPNVs
L1oLW8Bd9V9oWeGQ1btUlxnGubwFUDeQmtOIRidrXfM7+EQnXzIeLE+N0nsgf22C
D5TrEY0+C0y1Q2dPk4GZX++GlDuE70ftfQTcIYfOw70Af/qJ2xY80cQZNZZxRvhh
2iU99fDXQ6lOdVQGfyANXOc5u1aD6UFb1JF6mbklDc0/tKK4fsYsbYKZYzAaihD+
BfELi1p8fraTlN2lzoBUMN5DLXsnbRtJUI0pbSHjuWFma+nF8IETTFlstboS9q+T
PVww3IfGg98xK6OpoXCcc2nD5jcotwb0ErebllSjAgn+p382oYiu7/jyaOR5SxiT
apqhaJivUOxwQYpFNzxjeX6hFTxq1oYepmGcZ0J7bvhWmeffI8BFRWSqvLwtG+/I
psVwjKl6CERBsAyiu+8vnrDmd2SUdItk1cnWe3daoLqzKlz4qVaT8vJ4W0xUpGFU
7UbrqfY8sFZiNkvqtJ6AazWVEP5v2SFuZy5dTc7QAPssRNWm+OsHE/rz2c/sUXl2
K70ESymujKX3JQ5B4tFLNqOENJqqZys3y++DFOFq7nRWqCS3kmavmKQT+ekVNO/s
Xp8d9P0YTV5EBlfOqbXaRBrtNSHYPtpX2j8cgkwpF8OMZ84FcNzFIl8qOyd67N+I
IEm6GIcOHI97TTBNucFbOwi0pMYy5RJvX3navnmKPHfoc/0QECzHy2qh2W6dZQkj
+6SI+b5Tc4h5lVkRyILEVuAYH5EOA3AQBobcaFtcB1dCkAeHnQta5aeYiP00pnCc
m97gReu00f9eDIOzL5OfJ8WacNJO922NUD8gD/eItzV4Lqk+xOLSrESnvr6OYHJX
9IyhSeLbvq7ByCunD6ROTQFA64LuSq9SsfXMq591LCesu0xJyUG2DN7cXk/WE8MC
pQuN294rnbdlTYJoeItOPcrDh6+E5XFdvR/p/o2A/ISAlW+/x6sfmE4EsqmUOp26
RriLeMpFQtgQ3yXDpyuatyH06WO4epqeZCejczMH/U2CNx0cUqsyZlBoZuqPg6HK
MsafOesQhgUtesrqTv0EtKnelUhqlw/xBD6PdWE7+gO301eo8KiLEwkgwIZ6pW62
F8Me74UhhH8wKj80PFqdx1ntZDriVPeRXL7kc3UkSJeS/gdxfXI1D6xMD5f2c0H1
p82WbCzlOBvbJFW0okLBxLF2TzB4jcF4od0n4/vSkbhuDm1ABksoy0vUzB7kh3h3
WJiuf2Zfh/2t1QLobtx02bafq2hgTftj3cVx/4U7qDUdh0gbB66vmJfzfoX10YnQ
+zm/NVU97i3JBCS8ISYIvU+8FgXSAkqptCB1wM+1ZO1CN7zo0S8S0AKePnYhW6sd
Y8QN3DQL52k5h6x0eMi93MvtjcHBq4BAKGFnnJwbbZ20UJKX4zbjQdt5/2zNMyaS
nu7P2tHs3xPrKidOpV9dWaYb9GxljKzgwek2VlD5gAfjC++2uowI8rFfMiPkEy0T
CWLllgAFPUB4GEKxcAo6/ip8ReKdUa3QG4otRGVDlvYCcnhdEBpUuvsvCiuJcP27
TauC+V6o/3sciqib/mocnAwyJnaSKuA3xFfjZAnrAk091OvZxfFVgFPbe9YYQdLt
5/pFIGuMzZc6PZTE0huUzMT4apSoACxneagK22CGc4Daxom4X213Kx582iezqswy
Wid7IJ0fhZU1pOH9/Uhz5ER/dGMs6ec0YpvtGyKkEG/QRbWUIE0FyazDAHb8Z+oY
393Wh3EwDksCa7qL025D96d/yNel10FCo1q8401AUbNlYTLC+j7nW1OeXRS8f3YZ
Vc5Qp41lBfXVlqLYUs+uo0xhe2hL8PnQdseQym15pGQKxpFs3z0PDXwRZhI2+VKd
PwVys7TMneh4Vnb7pv5k1n4DCZnn/NrZ+WfL405lu/AGZa0L90eYsNaHVBkwVuc8
wIhoWanVyDC7AZZpv+AtAZHydpaffZ5RLq53kgoeqdMq0g+e/DV26n15F679v9KI
5S9ojJHIsFHNXELQTlrLefzoKktHauDvAmg307siT260l83+MKk733yDCEEzfAaS
LuR2+0JT4FDQzyfSueFWOZq3rgNPdFChXxjR6QtLNl11y5TJzNrjMilvZ+5NSRZr
4N8ppUC6Mcg8mr3/3bdp1qyF5q3gADRWCc4B2be0oGyCJMh1vxgZaI9phRbKwOS3
hju6FXK/MwL/5UMXTDX0Yc3HQBjdYgpOI4+lw0f2ab+DpB1q4dRu3vL2JLGt/k4W
xFnTAr93GOVed/TnwwbouqHEpH/0/lO5pMmN2GCUWdQE9HabhS58mlo9xYC8Paln
i8v6qpBEyjw1nmj6ULJAUhZ2+9Rr50NN5com7g3b1ww3fLJBBjE4PXOtBB/vzZNO
9NbQgF9msfCZnaavDSF8G8cP1gFCJwqliaxZ2XXV7VwrIBYPsfI55HP/91pgN+ci
T0oBUdik7J7MnKYoXPHtS4SquPWwjK6PVc1uCAHETYiyl4TLfDKTfhFRdm0qq1By
S47hf4ltb9yGwfP9wGLiBg1OPrZ0+ym9wMm5KJdvQg512Ho9Jy/ePyynhFLrcJeN
O5v2x74kOv2XCN7KLpcu1dm/RC/K4vZPsY3SCPNsI3NwR5wQO1fJK+aeUERwei0w
yXxjqXm6KDgUikDkEMzT/jpU353J2p6IDleAbpFOsgxi7loc14/dm8C5RjPcq9OL
QrE5U/xNdX2SrrQwZDu9XbABWCLjkDm+Uxx3Qw0MXXAN6yu/6UoTQ5IU0w1rf06z
QpbgD88lA4yVn/GB+DbOLRa1nlNobCImrSXObxzUFoXrRM/RqW8UecrZsllR6ltA
AWWFPhCr4YN0NIzP7MuWfg63T7SHCSfWv2wa2T5NreshKVMynf+HHNMJaYqO48pN
RJ3UpyZz32vCJQMNjVIBHOzbO2tLzdLDPZ1fcGugnbneZDCD6tLD8PS9gosOyY7W
U4K/nsC+yN+WKPz6ecJQkCKkeiSWj/w5tNi4INLN40BlBwc8zakVB84dxY6Sj7/e
QWOdeZoc+YGZGhcabMol09Zoe7oYiBDc1aSL2iyi+9Yn6Mh0zVIA6meLasv2C7bz
NVJD78OAtv9RaxP+WiDKDGdgeDzmENzd0pekZxVH5RBYA/SrUMvvQSVFu1ARSbID
gEiCjvjbM3+fiwKMkveU1YnCSt3eVnhkMMK3sOY6rwo3vmaH356FV3mCZ4MVPFHG
HjHbT9GWxpOA5LRMyhT+r9gehrKn9spZWYa0HeQS2JM4pAg6GtJZe0h3h1ZW7HF3
nnLZMjpDRWX4c9bgr3i9awctF7Gq9xPD+48KHU7Meji7thT38Efk01datbsyXV+2
/vWGPPSItbZZrixQzuvAfvMqks5KWSLSE1OTmi0G3Yi57WtG79M3Uy9iQkStvBTe
gvdsKXvllcX0Y9E3f/L0h6pjRaz6gKnewaY6MUjaIv1SHf7ZhC1sYstq7npCK9kL
PyQio8qwDWNOlpZgOd+O/BMeXxrLb62ePAMkjFzPg3tJyOV5m/ypi5/ThBK1SMW0
Y28/VsQ2cFXL31jqAq+YfAorO++Cy97SOEzfTCCW0e+Er8iysbXhkXCCe8bkVYuv
gGMdf6XsXqdRmbj+P2r8mzKOr47aNtHCXrJqCv33zVrC1w9SQUGfFbAk7NuARtQU
wF6K7fbgjQ+2CEUnr9gdffR/aPBW+udpNJKqKu3aMaPlMsWQTU2FC0DHiWvrNPks
/SpuhnqHIJNDxechclbcFqVwBC9w3k8krZ59Rdbd3bfpsoTW8uZs23M6EX7SHaOi
W2qvEiGGnXMlCvY65QaVEz8vCDDtTxAQ0cXWsInLNWId16DQnENSpLTPtiq2I/AJ
zpup1AMFl+NWSbr4olmu0MD11deiB7GFqwR2LoM0KXZ72ZDVXg3f0N/Z5rPrEfSi
GsldH/mUZA8WOvHQ3oCslNIcCOV4cYg/zl3j4nTisVJY6vy4atS4ZSSbwAxEiqpX
p2BbkrEsy46kBrLKxqLQ3h9qejxLyEHNeMtcgrcj44JYYukG/uFlHGcFYP54FKO0
C4kjBo0bZDZDdmlRC56OIV//WdzpZ1hiWEjE8akpc8oNi2Pc5F7PvZoik/93xpPk
BN3U9lSveZObUPsfJ0c6ztmQXgW8Lq/kWrUuKOwQ3zlYu+WIWq2XCwGehM+YO414
IhAF2Rt7B2J+I0LoDOKqPg9yLyBluUKNaxoIAVko+cv2FZZN21+cDJ+yCKDyWcmT
ZY2/Ip4NRHIeDurK1ghYAZ0Pjju3uQzDSPEsjGypcUrUc9Y3kHphp3e3Wl5cGARJ
SQCoJRPRE9d0YWCJemrO2lLREmQqDFwC7A/x9PjDCDW6if4BJySzgp6PS6zINKPA
VMIJJvzx8h3/IHjZJ3gf511WFGLIPAwW3HfWR6R/PzLcVrsVXP/uiPx0MSTI2ZLW
kaSLNg4K3eMqd5daBsryGTjZNAtVOF48VT6NRmVSuHfWxHIjIZDMppAuD8AslzTp
qvjy8Ct7I7AgmKbFnyeksLRdFeg3N0Mu5QK0L4i8PtOxnJKQfZWb58bOWeeZRgB9
fRGQHKHBdrORhH35VVDQ/IekafjV7uqPdKNM5R1q/jiiBmiq12x0m6LD8bsZowSm
B1i17fBAm0CmPV6R1BxSLNtjEhYvzkLWxKQBh3DAZGbmHjlgd6Xgy+yweuOQDCV2
bIEYvOw6Yngt23ceVeZ+dXyQl44isfNxoId7iRxROO55kB/Uq8RdAObRZi08Xxct
4OWrzvJZDyp8aMWDyNXT3dsjr9YNwGtND/718ltwVbP+j9y6N1kopUoTk7wJu3nh
8uvt3dB6WKHj7BQNOS8LhbSUzrssKvndlFhrS2dpmlOD5tESB62YJ0c4nggs11sh
1Flm4yE0oHN0k5OtynBeetQUo7ta33yw3PIkPIDjLpJmoMcyxxL+2QYo3aZJNoGg
J6AxotfyFsYhKX6M0W72fmOJr8BGZMFxTyZF2h3a9ix0J0vZmqt7rWW1httO2uRA
BpdO1Y/KS+OCDXvFPXXEgDCeEVkJEOHq6PqXmyVoc5azfhmw5lZR8m8Fg03QAAhB
9DqMdKm+wOUE9Pa21mormk8ZBkfVKmMN+HAblH5w++w92p0Vj+a+JAWuo7n5WZPs
9Cq+a2qmLe0YBEBxCG/laF8LeOVGa7A8Ucs5Q277sdzy61cPevzBGocGVe6KPyHc
BDqrL7xhqss6q9GB0++ZKQ3J+Cb7+erzlGOrx3bBjhQ7tUogdji4E3IXpGGen1gn
wmcQLkX8X7EGEq/VSmybJ6QPx8uHPbPi5/XCTIf3qkw32uaeqTNlPs/4BbZuVxSA
W1sTXz/16eqp9sdeCKIkaBdgnrLsDug+ADltLg0OnCB21HdjXJoshbj1cJHlgOda
VgcOEQbVTaj5U+5VFRDLFZJ8gOtBOUulQFILQA/i6VWT4QzewttFG191bOPlv0RQ
DZptTyCxGIwTqptSt5TP8e2bktfrs24EseeJsZqIEp6BjXXFshuBLJc6J4knbRv7
lcx7FS2viRTWvlE+IeN8iiz+/bD1Mp5c/QtW4IH6XfCykmztE1QX19heq0ygsgi/
0JFxwr53XHvcTKy4yfBB+Dk2Y69WB6QDA5v8tUI7cNfSYe3byScXO4jFOoKpmen6
Zo3ny11WccL8F+Fh9lUcMOesG/Awm7K/lJhbvIXbm+UEtVkOB7t6L2VSERS7WzOT
50wpCnes49rog9iS6tQGrMkvNmZRKMMjzAFPUz9eDE9WhOcq8kLylfTfD56PL75B
gfaxQU/MjQvZtLljrtoG0jxFrrBQkGtM1SRT6NEAvTByC4CtUkAtJ3YNBfBXzo66
GfzpcxWRQsqaRjicxrWflecDjfbkFSDub0vU4dE0UHite7GI1mKpmO6/HzRWH+mx
38DRPObqjkULN45M5AjCKz0b9HhdjMBmdNoGs8ZkHF+hhcm3opi7AAEWR8EZthKs
2grtYgd+GkBk+BAUi1bB2nFyp6MhH1ZX9oLym8Iv7fT+RgPBy18A2hDdwtR1D8I3
pw3Ir0INi+I4vYwIoCSNjJJFPaXfwH3Z3w9LnzvvuccLKtentBsY8dKIfPYJnxGt
NOh621affh35hOK8PtKgw+dvgX6EMHy3H+DWfc/dCc8pBeFeO+QKlhHBBxLX2kBW
3I52x96HjY7u+Qn79KBP7Ke0O3I6RitrL9eaJN2Ho21KUIfOYz6kDJWSNOLXp3FG
67F9wDKakB9NicKGiU7HJHqzk70b28f/2WHhVc4VIJqhyB6B6TawLOSjAuFLmZmw
sI7IR3B3h+BeWhjPbYlJRas3zzt0c5j6FueSnjc1iuycPdhHsnw9HLxu2p2gQA5m
pGhQVMG5a3wP21pQuxFphMh9q0fNNiCaL9v3Zyj0TaZmD21S0XRrCFx6TCM69Ih+
CEXSotQpckEZV47KLlZtpfqM9dQWh20NZHPPQveCjAO4A6XAWVjp7EH+ILl9WQKR
ouDjd67RRz7pYYFPreINzpZe7kqdz8jRqlSNJ/tvurDOm3zMfMn0sr6hRntTQZG7
oOwAhnp3S+7mEtiGCty0OA8ENinn7Wif2YtE/PMNdhGrZZlrfK+pq7MRjSr3zI/B
YRUyKG2dEEojbITMC/JymFSRVra6hz+al0+/1JdtgO3E9hUOXuG8me7/NCKRX8pE
kwXvOTHNcBk1EmhWj/7yf1R20Z7ANe/H/oOT7PjxZi6zGdTmap4vWnDq7N7K6Yjx
dQRUj74TSbewZLlJwpRbXUyjj6rDEVEgj9JX14CPqIQUnmb1y1CUeJ7l8kbkc3A9
ZS11qkXGsXCS8rOrzuckv0Z2u8JUddqyHiIuC2229JdUu/ZXNnmCqNrpWSw9NCNs
jevUT1LpdxlCq+G4gvrBdd5QtYSjFFTc0jPRY1CrPElNHoFITYBijlaZYUh14Cmk
xbONjx4A/YMhzMVHuYzZ+5xc17Zqz70Pd5Xspey6KYpwse2UwbZ8w5bwDfw6RVIK
zGmL+fbFiwNOCkyMbTrGCTW8BT/E4F03PxCSPqhh5FaIriyAOv0Hf9oVAy+b8rul
ZBCM0FZ/8YOC73TFTO3MInwxqWq5QSpRL8qjJk3ykWUkdPl2AJBC9BWL+Nlyh4rW
ihErLUlK0+K1K4d79DSb1qLf2gY8SiQMsx1dXfyUhkFFcAA6XW1q99OJ98m9SYnl
8GEUIhWkHhRBingvdGa6h7ub6NGEfVB8HP9m0gfwLmvDYQPb90NrZl6KVBHfiw5r
RnjdVjMounGk/tjXyqTTxKXqhqEEDr6it0pu4MI10JWPMysuTSEhaMmhlinCgYGf
PuKcP2z1DGQYsZxQrvRr4unW3CTxyymUazgYAOFn/Ykur1v1GVIhcRc9X3q/LdJT
Vh3xZgv0uAIHfBQ1YN5zrK9g/Gcp5LLtGn37RqW5vNyIAu8CbwgyLEXNeksiv0Wk
IYHq5SnTq0srIX2/JWEpuZe3A54CVYPvRnfDriVdBeSkblC+/dbPfd990LeqZ4j0
Qdo8nCtQBNorf1YksZuk4duR9lz4ukcFmUy/VemQ79ZIVxiqBF60aJIi1868uJPQ
WZwtu1bAhd97xwvqK6gXrho4OuflY2CEGJUbCMi8wQMd6QyvFc3du2Bk2dk/jG9z
fV18YbaeS7F0udYrQjzKOgSV3OSVzERL3jF7eMPTYayChPUwAJHC7dgmgtuTJcuu
Bk/PFggOK+z8fiIhDSn32TtJezq2XEemAvd1yEQIAI9AAVjjLCm2VnjQnTa0DrkV
1mkYT0FGvPiph5rHkXrH5haorzgkM82DP8THofpAHWWJ79DK3RZKSuN2w3jn0P5i
RXHOJ/0KYJeNhxkvFIBAT1Al2Reew7Y6qSSHbpz426AI0vTqw+8iDz1KYIdFNBIn
HrNJeMEFnbYG12OU+VEwf74xD7O6vFV7KzT+ygrIDk5sC2jzCVWRyGrqnYvR9yre
am7z5fqZEB26tdKN3D82xOIVJbd4wazPuroujdE0ITwkN2Dm7Fu6IIe0p+M6l16R
lzJ2fV5K8OdN5UqNbuiNemKNgbcAiyE7KA5pKGzPmAgke+qsQEe4wNE6xwHwqmzV
zYtPYbz1mCGbqWOPFOi79wfISDm2MEKbPCwnwXIJge9qyGxu0IqJ2Y9v8S60ttrg
tr0p+uo4jaaGjrKyOqyRDM3FHK8T6Nx6koAMXcc05Q0CzD77HIkZ64KXSM+tGe5A
R+Amx6uBz1xLt2t/qrej80jylCPt+2wvdudpAkXGoEC0A+DnF6S1zD1MRN20SGaQ
qDdtCIa/p1B7eeYpDSD1jAXieW8z+CPHY6rvXNWgkTgZqh9xiA03WQI4hDKh0Nq1
UMjPOO3BzF0CzkJ65MXPaBVrlVc1QY2f/2qYFfeUJv38BHt6/kUo2DV9v+rPAxji
0MHAwY5cZXhK/E3T8lQC1xVXZTD4zqVIb1R1Odg0nPxtGQmfFAZbTm41WnNYDhl8
YZsLoX52yHxkqnayNphqJPOSL+bxB0KD01Aj8abpkDzPc3MMf7GrCuLME0gspW1L
DXsnsO047wjV2HPmib7454E9+pJb1ULuFU64PB3RNg1exM9jNZ9IklyPE8IT/Zpo
xzBJLZaTx9ZIlEoCWAxbkDmUZq0cY/sOEJCa3DfkwpUHOVJVXMNFMhBP9+y1n84O
WkzYj7Pn5UMwFhgbqchIy5x6/ooCxOz+MuJ8OJaG++IkqjpuUFoItTM9pq8Gizss
fkipuV2vkXuJllK5B7bVBeQ+aXVlx8kvBomV3dTYqxA0oQlFBfukDltsdsNWlHj2
I16dPR8MUIco4ifqEnwoSrcb+CD/4vBIYN9ZWdCJKFn8cnxSm9zgDGtk7EUFUWhJ
RkCzoxg8fzUFSn1ZEzIDV0pVjfxXz/c+dDwLM+ESi1kL86GyZVOWQWDjMCQ6N6ft
sr/xNFPJ9FCdei28dDgxGGufnWGYUVlRKrl/+sdJDOwHI9vPPKLbyiTQZ/82bNb9
/ZWSbZqrBtXOey5CMjbRyjkz6aUZE2Ej/iYb0TE6+kjL/CfuCer76X5dudbPMQaN
x4LYTyAiN9DCpW4khoY0C2TMRcdHWv9a/OL2+LU/48db7OjALud35HHbbzgwI3y8
bxdmEFIptWVX1ceA/OhJhOHHqlT6eUguz8SW18sk1EqLJr4KD63RoPcELeW7ComY
3SQm4YhrWMk4i1T/54beSMIrxK+m6GYkxzLv/IJyFlEcpXTI5pFqB2caUIboJLnz
kesd+4afK8Hi1vuQWaMI+q72u7Yskgz6wJROjeeVcjO8s8fk26MvK6EqptnpWZnS
1s6evFpkxpV4ahLBWRG7z6uXLnOwkx2rImLtqWF+G4kFxEl1rdw4dSbZO/E22ryM
OPPSGdPG5gk/rKVYvcUSwbdEcL6WGm+++RqLy/i/mKtsnBPWriFdu433TV4ialLC
haXpvnAvmHsV5s/T7fd2FHkOitjLpnkYG1ZQ1ou7tKozD3EWnccUqCAuVSFmZ4YC
va/Z0i1UkU3v+x8y/HUnApwpUkk6+GSzism6gYGFXFwZBTY2atb45+xC40Qosv2T
i3HFVMwbMdcmOppFDKBCfrY3kKFgOK0Rky6vY33sTjunYofjAMuNu6VAWRxP8e0O
CpvlO8dCJN1Ejf2UtqlJRcJIwYEi3GY6YO1ZqT2BPoOp6is6O78RBpwfqp/pf5ai
oZf++igp0dKCuwvmAf7LJxhcXijS1xP0yhIh8Oyoe1y3m7X39egfG0mKr42ammJ4
IRU1vfqJ0tEEZIjPM84BwAwO8XhH8DONv8V1wU/kA3Y5XQ2FmGOOJRQaX+21h3Ct
ENVStwLll99y3L5T6lPt53SGu7QGrsKGSd/B1pmVj5r6kALpczO8VvBS9l/0yWIA
pCZKMvvj4sRLSxYQhIm1Nqp/t98V+/PX2A8BULGwPPLbFqYlxIz1NVmIVnMn1xa8
lqMjv+iZ6YNbRMVuUHCfFDbkCjSPppNa4dgx3KDLIUHoE79cmq1OreTp97i3eyFS
aP4e45e/To4uX50svxDhidhVv/3Sz+4faOcAF5VFTR2tLEjj24ftZ/yIe3WCHawK
4nTNdTb9D/jZODr9fNP/8tAUhwbRBekYo1Igo5FUe6xshKvWYEWz+sMqIvB9VrLy
NwUFqUZK4axc2z1MAVH2eOJwmdVjcXWoEJLy8ek0Dgr7xngkMamhoXFHNOQTlsP9
AdS7N7hFh1fWLJdqku4BX5SurQvchr0F4QHFv+cZeY9tnb8S2XZA/g+EMDpxWYVV
CIQqJ37cGIH79GQxYNJAw7eDN9PAtjF1e0qufoA5ATPMVhjZhpvqzEZybcQgrGte
S6/yIUM5c2GGHVogDKeILrtYJ3h/1Un0a5VdoqUq79XSmEOUJsxvxYGAqBoK39f0
/xPAS4V1pMEJsfyqVv4BViFEPJA61UcDTG3NO0rfR7jnbDBxn8Zbr9sQj41rZ5Xd
sPSwJz/uFaLUhw9EW3GNsI5Hvoy1wpX8YUbVwOd8atXxNyb04gygFSFe/3oCbDg/
WPKN9eMa1yEHzK9Q3CQbhnandO77RuRhvAHl8fvtRP7v2L6khQ3FVb/4cHfQdQwp
6ZKHxE1vFQ3TQHa1Q/AdjDKg3vd2AzouzEfS2ugNxfU6li+bTf/GBXnC/hd75uaj
tQG7Y2twZfNPpQkQ1R+fvsjHEqVsQppS6rr87BXkunynmEhfPbT9DS3Ft4aqKQnI
053Am4RJsEqjnmK1zEJKqF/ugxDaXROif1Q4+3wSyXWRm4qEEuukijXQzKyLVAR2
a3oTA6DyuQK7o8GrH8bK/bgBqaNNlDz+uXQX+xvbAD+CibimvZtgR+oF+7v1rjmR
pqd5+Scm1FXfzqXX9N8EGlPmUtXyWAo3CPwajb0qeAjms+C7eIgXuJDC84OenTXR
QXy4b4J0MmIs77sDV/LnjbEKued0b/SmokDXRYr3P3j0/vUAn1uqBX5oq0vlDGzm
0XrvBW+/6qEvpokHwvRTyBz5sFdqVnuyfOWt+rji+1cKy+S25NKV6aLdWL1CPdWm
17CPK6/7MJffAaRq+ijc+IhPXjQUcLz09Lu6K7x65MlVF3Ozy44s2WfJYb2iX+z2
aRkipvC1Nzkfy9n27G6GDWhxszpWx5EW5fC9C9We82MzYDrXC+t0fykXuv+oPQni
zbss5B3H1mLCWqHi74fsnMi1TE6clJnk+zDv9mxjLchg3NIEmXuToUsA1oO6a/IO
gmYqjAHhxDwnneV7hHSt4SKnVs5LXzw9T125ZuJykwNv46kVGpps8OM3cS57ciZy
7qEp26I9Pvy822DaXGTzW5s8Ylm5an9MLPcOtsIXAbOqunQRTIGVq3cgtMZtrb/4
AXg49gMPtVlPkSkBYbL0JbmRXInRxtGZdTmnMEpExyacIRF/EvhVdwhwDxKniM4D
qEk58xnFcTVnXgUz3mpjW/ogDktBaQ4SZKtKJxTN3fDqgyTf2FPHvCP+GTJeW+fI
UIaFVct1WkZI0jQqhubeiUhNgjAm7hOAVRdFHK4vOJbICIAJWpvKn1BMLWzsE6u0
D64VFE7l/VjZ5RwXEfdDuoo4u+331S34Z15n0EXV4TlQKUpJRjC5jxGL7Rs1RXRf
pSKMfM+L6P6C07ZnDrUwGQCGaBD6JMdBzvhhJuUID/TaGTjpl7c+tGf5dNgdgrs1
tbPZ19UwHC6rCCsBeoornDnqNAuVXNVJfZMWifEhSvc4wqAMZ5Rgy1q2qvbO+j4o
mK52gsNxGWVwrTQX5A6A5GoiF1r/6n7n04Knn82ZRtVrw5D78/7QJlV7btZOdwWb
5XiK5EJch9gPhk7yVmsT0gdlX1Qq1PDGfktMTmh8VhgAW/BERTnAUvU5KZIOEayy
kiKN+DLLnHrKlAsEBPy7FCEJQ1q5QBM/2OP3UbyjS15O1/zU0qZ/kz7h6zSPp6Wd
upnG/ez4b9DeG3R2kKNpDjlt8V7+Oo/ewRvyhfJNMiA4utP7kP1YoWPm5Sw+tavK
jXa1hMi7Lih8Tii3zXUBgfZNSvPghLgaeHV94LscWp1MrNcjd0RI3qSmtYzRlC4w
NT6MnJYLpmGHQ8B38S0+Mnge4C0sdE6OwD+xNENU0Cv7DcYZuqudRk7aBzChyJS4
rQABnoNdVrpPBY2ntDoqVAeSI3ZPmKLSKRWPJnY5+vwDNUX0OZRst7733bsIpXF6
QxQIDa2M5F7eSf/ApjUFFlKHzPJbriWkBE7aodRPaymjFk3QjFaU/9VDaaE5CPtw
uvvSVnLBTA5/z7aflp4mgAv262CDZG63mcXGqDdH+o+JJyzPESbVwSnj4Eje6k2D
OeQX7v+Yftx8y5jyac4gsZwrBb/huAqur6xTeo+GgGbXBHy49fAb4CRfVKkuSngY
UJKs0GkhBtyDMr9VEAAzj15FMP45ue+lif++PAs7Tr0H/h+SaEev9mDeGVCA89jR
9MGKVBWBpTOEhZF+FGckeqDxi3Il3vsM7infPZ2t2BcNgr5tE3QnmW8cdgSgfiVT
SgkCDNm3qfSbI8VXPAglFmbnBXUdOj7Zhak+5cdA+YgeoOWdDKOM/o67N9v6ko4S
OYmgCyDHK4vwNtW3mdfrbu/lR0DrklRy1+kAtGf4czBobxxKqZ6MFZKu8434DKZa
P65Hm5KDaGm363/21XjoLsJU6LKQdXKXPjp2KOHcBbs3ksqTw3Xa8w9XQlo5KSE3
CwRr+PccYcP8YmUCb4lAb0gX3L6Kc2gOYx8cnx0BLDoA7Yf5XmfpcBn/+JEhrs7+
H1HdxHw89H9UfJC3hPIM1xMhql5a8sRmElCFzy/MSVIkF0I9Ws0m6NKDoMqt52rI
xcpSDbcfHIv6fqPSCAjzNLOHq3Dc1xXc3kqQniO8tFbPnAGk/XtBo6C66KvEdAea
aFhFVKTC8w+RmJyvWBYBxqomdk/KGaMkXMy8E3AjehjYHvShnriofPuUGHNGPRIu
3mJEdM+dapDEVsnsklHvVSXleo9urISnO3zVpO/3iSIH9I+okWTtVVyZI036JEvB
ayP47vXTPTBTHdOrghvhuOsrta0wM7xavoBW6tGAkkl6LTOnLxWx9HqviKnGbaHS
xvgaw2hKoZgUjzQMdcv/ex3FDZmjY89HBh+9+y8ps0QuAka8V4gGo2CK/MynD2yF
lkS5ZWOGkDmrGYBF4l4OpH37hOawq/2QamisQLS7Y2vUI7CynNT4Sc2X5SI0rFiq
f9aLra5Lr1HzZqV20eeRiDWgV/vMDERba6B8s0KovB59tZ8cZ5mn1RlWa7s6/NLj
fIcHWpWqmDL8GVMRVvUnvxYsTa4nOIfElyYSjt5iGvG717gCX36N0WPruSL33wFi
LLv8xrboaFK5110kjQNQN3+i9KnJ5eGrHDmofAF4Xm+KyLiAZ+4XnVxSRoRH9D4h
SW1tkMW7G+4IHHPLMyMIL0DUYyCye3JxbAge6OJV96bF3ieEqEEXsZ6BKfSyfrDS
HyLgJiPfnVKH1qjjsevQKaE79qwU0THp+Ukiy/Kti4v3N8OEQtgn5Ja0BxarlKrp
TZT5HzqTegDgHSCpvqcpjLgevU19mt1P2YGAi+FZkYXRQonzpe5AGwYCkhuOPnC+
VoBMZucGNSL5vqlyZcf49Vgt86hXBBXUQLiE1rSXIxiBwEJlcJpEMPez+pmjIM0F
ih1Ka/HK4mF1b9Fdf5EyLAiA8PIbM01nmRfjEeTuU5dkoSPEzs11dpG9NR3rNhib
hdPQhvqo/hyeb2LSm2egtmWJfvvBYA23hRauZmci3xpyNdvopzvtZzIcScpqmeGt
9wRZsVEREevLmzKM/YFrHDtWBRtaYGbJrig3/ZbAcxAUwI/lBESxFSqkpCDFGpU/
Mz/7KrS2Rqy2SkaCCVowHg84CIfNoqgameh6n7LDofsDvauLeDgZDxEVaPR1pdEd
AssOvoCQHKLEhhyQTm/jhkALFYq+IvxeeSw7h+8VkQ54dmEp3wdPb/OuKzN6oO8Q
zDccx4Vh4dGhnbGipqdJZvABs7E3z1gOM/5XYsGbQ8nXAOmYSDQ/mYK9xAx35Gg1
RPXfTAgS0NSZZxnajdMyUj6EBKLIeoeFCmBNsKjq9MxalMmzoNbWBxyCLiVj/e5h
/6qxNI3J5IIYyV898zaoC4ay2XpSFI7PeQZBgpvgBrXI/PSS2uYpUTK3oeOvnCIr
Gct7sX9ToCoKo2aTqz+6TCOOiLinehr6vMnQoxc/15Oty2urwSXPo/mtwZrLXGzc
7uUXyrlSAdir9IEhkMWq9swRGLU5SgnKz7S+SaFA6Kf5Q6xdkLKpi4+Rs/1Yb3E+
Y5v/Q15p10ODmCOvJxGSypUiGNB2cOOgWNtYY4KbP5fu+Za6r0P8vx+aWpvzj/Qc
5fLrTGxAcKNA3oZsfqWNt8WcCkMuJSNLKJFdDtk9LAYLgLy86lhDYmyj4fFKo0s6
wHhGb/dy+zvhuntNfPMgkoE5rc30gdzwwIrmcOhZDNy7nWTSa8uyjZ4rjhC2BSFI
PSkYCTBM5X0AfKPgC+84jMOzvNIQew4Lmy117Q1Xp0BIauXfB82ZrhpRYA7fZBtL
/xrulj4teFu+4BiHdbZKSmnr1EpeaYYHzEFKgl+1k58LX8mgW/JHsukiQXsN0QTR
whoJkV1/sqJGv/Bjzet4SjUjULdBxWkwrCG00iLjpJ/3I5Gl+E4bvEjNckzvEao4
bruyGBoQlb0o+oT+ylRm655qooAcxAPUDQx9NpY0gTZZ46moxDW6KKOUt440MRKz
k/j9M2R/D+Po4qAmjoc7cqHPL5DurQdI6+KhL33wu7bniGoB1Cv7KpNbqQ6GuA2t
rdY1ysBPcwKMR1w+1kNXpJa+PUioIrVD2DKJlaPYDPU77aWaR51FhxUtY3anPM8M
8A+dRMCejmmwXvScF1TluAB5RW4XoNHqytp0Bb+e7qpyQbnsNxQOjQBlTDSt7nAm
iKBeSg+kY1bZUZRqPq7WLwHUt9qLCvo5B2Z2GWlw9BRjpDLiyjFM45PPP9ydKO7f
8vCApXdZxMlA/6ShDLpnxL+uScPvLmTnCOkc8g52lkDlO6UDK7lBjig0QzXbyOWF
CcFE9fqoO6+LN2bnr8ATaC7kWXLBnhPXcRrXVMgsNorCgQBwaq3DjRjpRKbgzEfW
FN6d1Q4rIJb+QKD+tzcgF5ceJKuHvmA566VtOtxWHafgiLwYcZqXa2jKX+K46HSu
FFOv2FvnryolMqpNdnrzQFmFbL6kYsylKzDncyjdB00LFRrXMeevMqbo6J0iUcUh
ba+WUEFqa/dR87n976cNAV2oVKz31eFwMwI9bPiT7NDWqcoePbhR9FHfRzHXx0yA
A1F7+c5si1Fw1LXi27c0MaSPZk423Ffcj/Bwp2Uploeh0AojBWVhYZ6s98bohBiD
o9jGdtG0Gg0QBkLEweyAxycSowAOOprGwjtOV3tWTPIl2NUL1e4uYku28MnjatE+
MyqyeKJhBwRcEUg+zELUPQE1K1Knd6nXOrY7df4vRrhsrW8prPt+pZz8MnCMgbNj
VC2YjavbZYUwoO6sQdFmwR31qNtUyuN1DJRktuedRq0jPwUt5yaoK5ecnV784Kay
fOAyUuTCIKx65cg93cZp63dSS1+70X2uTib121AZ2pj0icoAtSHWzKVUURoe48LS
/mqJD5l7siuutlbu5ytxEhnKNkD669jwTUb14iF1dLUQOUMdTQ0QVdxEIPcjkUBm
4dY/SnX6SZoHZtAw7Wv2b3AbiwfWt4s47dKHNGWuvJKpKhRBbdP36Naf/mKFzp3m
GOsVcbPj2tKzFQlVfAM4IXhAPasNis2fIJiVsKViW2Ntezw8agd2urhVGm4Vg4Bq
zaBT4jHtQ9RPi8o59B8QE1sBevV48+IFRuoxWGJk6NMGIIK5LnpVMii2dp22iXqJ
5Pb8xmuZhvXGe5HBcyfdDgkYmbeF03jfHYw+fo82NRQGqlAgOhnnJ9cdWUodx4g8
fcUeBKUV/0+M9id0JLGHqEcYHM4C9QvSiIr0I73QwbEts0L5Rqb7WsJU/5WA7P5R
vb7+MiXkBHtFFvJTzQ+SPT79haMenUK6elfo4sOa7YbyeGlpHBx+usp4EuwNuzIT
a3whekUolzhOWhLVoxYfuUPy1h1SEQFA+Ozjpb6NAdJnf8yffDFlvDgcRgBTJueF
Glz+tSuPdZILCIoNP4cJFiM25ToRJsCnh1Wmm6NhevkuPDwrUYZmoteGBKzKnC/G
w8SDkWDMFrR/9fPDLu0j09tqGAaKUHm3dcBsrZSGXN20GO9t+ujNy9A71Ea6TbCT
JsJjbh9gBFZJ2FoIPiEOuSi24sX0F7+nFukhDnP+pM/tiL7sa7nE11hLkOGX5KXC
RkJqHUHvf8P+1BGEnXBs7vAjGUYU0Hcsq54BC2xfRF6ZPeQi0uyiyC5X3Aeia1x+
RGtwVrNnOAi86z9kZFSg8dpHkkYW42jwkClOw7vuGKH2c65oalxcUW4O2eqjAcKO
xL9bdmPb1vJqebhJjVAsJCscbTNFM1cnYa16SN7ehAH6OB7lDmYV1TtCtp3RIuj9
rSkHKOo7UNOsTd51sGuB2F8JHE7zwq/flaCfpfu3VQBLbC48vDP4D8CvZfdD1duP
RRExbLGZ2te00CpROr2v8Kq4+71DMcqzkPVaeidARyR3can3KYFrP2sN3HYk1PZU
u7bk3PVKZHsJBbYYuLp3IPZzRQ/RdOCA2M53Mzte/URv4YxURuciuyjADTlZd93P
l8oR45LZsKsMTKjDyf2OFqWoO3qOXm8yc+2FkzbweTYAiEAaLaIgCnbYiT7SEfWW
6liYLzDnugnj0L6IbFu/prawrEB86HUYR3i+hI3hwp88fHQtwy9C2Fi5XHogMAyX
UU9nbcRutvYmyn17zdeceGjVdApenyoSKN9hTwPapoYCUvRwV6/mEFw4bGAWqsnM
Ht15crdWBanrb60c01UoAd3VAe/v+sRVHZSXCC/XX/nt5pa89j4dVHcbiRdVFbka
HEBqjYbS/vjBOyuN9dHnMAzFj7IKrnuqynmQOJFdkc16cIjlpuPYk1wst4F/+4iY
ZxRltcp2TucrrH8xoHTpeE7O3TBggb+wymijbG3STxifk1Wt485vyXQjEzViOkql
1Ztb07Ot8VzyqksPwd0UsM0iD4SBwzhnuB5nmlS/vz75XVlVxHkLmdfiZ3bQMaU5
B2NP8QadNb8FykGYYtaw2lV0lSwxOZYnrCBEOzz90SqXV6NbWfTgUakInqBZYrp9
TiX6Ndt6bH6KuXlOxwP1qnN5fcRpOTLiQi43wtJbIJvqpqjZ1fZAQpJWeXtVdUnS
yWAlo2f30K1hMRtsKbQ9JImkk3pjXVjmaDwJ4ej6aHrbHDtKiLsMm9O9b0x8Rtg3
s4paXnaVAA7GuxzdHdUuqUHSqbj8CsObMn1j3EKqimBCAe6SK00kqDOhuDspt0ja
jLoPllAeIgQehd3Y5e4AA+uLzPAeDa/OudAkidqaiU58VRqECutJpHaQmojOc+ro
nzbKz1katVEdUllO07RDbmwLZQRmiwfANreveTRPNji0PgnqKqgsaIBqNM0zTVao
YkAXwnwENmAydjIPNfLAm0DQb8wzHSUCBfBQwRt/p6rYVM/1oLWi502vwjCP8eg2
w7VIqfenUXOoM0NluY2JpIufcAdNvXfq18fak1bLX+uT3yC8LhJ1gF90xhq326Bi
pNgzyb743YmfycjbU2bRo6ROB1YLHOCy/dAaGlZu4D35y6gwtoS1q26oVpcWKxlp
tAFLgqEoP052wYmp8GLYuC87yg3nLrjGV45ZdlCf1rUH4ZS/JN6DlDhw03L+32cO
9+gYIb3OCRzqBHma2COFHH4FrV12RGMfftvkth9DkbKjAn78hoGKuxwJswA79leC
Me0WajQ4vtuB/sgIx3NyzqlgMgqxp1x3tabU6DqCkpNAyUBI1zqMhu4Nru4+KsTJ
ekzVgBS4/5UBUW/OGo3HKUG1R++nSxO4+IumWgkNRo0ALUvgnZig5RWu+REClt7m
1iWW7pHGrwFrxFrxDDqUbUAZAUxuLsD92i+zGxH/rSuE0Dh7cA4cSCc2sf4kHHe9
abxXURLhoGlsW1UiO382ou6++J0jYmStzP0u0QI5pF9iBPTdYqxXpynwB2Tp2K6w
f7+wSBmeZ+U0+F2tvaOkUh+780sPRggpJ0u5bP894RUW3jfPcb826nU02nbjujl9
ixPg5Mxhp+tbr3PO4Bf6X1mmZG7zfiUifmlnA0hoBBIF3YidCeLbKWJAoTX8QmSD
MkCEte9rJi1SVkFGkX6JiLu0YKAbMEQDsQ4+tMHN3KCf6Fw4tjsY6xNa+tHonwKc
NyHy9yCcc+ic9tEUaIzPO11/BKOXpobSV9k9/tIdB+xmSy9Zr2cfzTEfK/ubWlwm
wmuWusSBGXdwxi1quFw7V1/DYxDzHDjWvUWFhxjJ9t7JgFO83xQUUbVflAjE3f5x
TgaCMUpKtz15CzKnvtVgs7k2bKrLe0EJPJE1BkMlqk6gmpdwD/KteqKn5n1wBGcg
vv0X7atcJoCPOeazF2zzYdlHMDksDdoNiyBGsEUd0FSZ1pXAf7kzLkxeVB+4RlbS
LGQhdtEpNloAk7jatZCQaJA71sFbXqNeLcpI8Sx9xzxm+OZLUCeqR/sZU9ADuc/b
fc3OzVnvrc7Pzu8GuCwXdHEijMHwHLXEU/EeWnRKpBpB16SveUIQALowQlJwKQFV
j33fsrCsfCYk5m6j9TlztmnrJ6m35V8lyEj19ULoAEvO3gI3jVd28biNmBXiNZfi
BbaVpd98jr+f1h6plRZ6g9r/e5cwXxujHS6pO356n4zXYCHyZ8aA6qCqpTLzKXbG
0ZQWeQS+c9sddzWMcdo+/FOX+YTLst5Gh0iQxF07WGk6/6Xzc6RPlX3UqR8Na/F+
QvMEU3k3aZR277Y43oTieqNhV1UjusCwoB2gpiKoGbBMTZqOkPWA1GN9MN/pe0g/
1xIEvLpCrnqQgpsxbVlV0++gXVoeg0cQsM/2sC+jj/7eMR7OC3D7tGNfNASvGhwW
j3fM8xUW87KP8bPdI6WfzlyQZ/NE6KGaHPTSYQCcDyBXVGhqCY3mA8yzs6pOHQo2
FV5zWnqYQZ1Tnc1TyPpnclRTvCX8T40Y1GTj6UpzuxXKZxqx5OxBsN93GyaVVGli
oOQ/O57vJMYGEnzNOGGG7oXgvb2UCA36BTJt5+BIsnG8hpgoGIDPUG/2UbfE0hgy
xPx36fw88gbccN589HNYP7WSLeJFF9OyBmyT4T2ScN0EKky3fouN06pxZ77ZrR7f
XXaY4/RgWdGGtCxNZ/w3r+Mxa/jUWidK5ms6W/6JxVrwwpGisx316m2fd0In4ZXN
z9X9ogofbChqmrwKCrzPbgmeYsWgUx2VI57y40xzQEKWeRkMPQm6bc7GLiMuQvMb
IrLAj3r9n/uVWHTz8vk8Bg3ikcYe1VTBMl5ZJwuEvAYhkvfxzdI+cL+Y4gTLC/Lt
1f4LEJl5BhG4B9pWPJalRDBxI/kmC32k3y4x9hEIxUTOOAX9/dxIN7peSTpMHzIn
spVS46Qjb7MQCfsSdqyecYibCH8UxOKfdOY1KoIqW+fAFlTtNrC7AspED5JoXL2+
lGC9TY7nOg07fLDPPr9O02zn1BUMPhtumENBrjvtx0JGKmdW1Pnn9aMp9pl4puGA
tpYefqtNuOIhZcbAoPch7jGf00nt0xV16K5nRhK5+Dt3BsFOoP0IdZFIXxKws5WL
cD4yUxHZzSx0m+x1XxOBgPD66nARmKuRu0V74Jc6/KjUrAJqVZwYucXiMJc26g6K
YMlOqnmZX8YmAh3VqvyqYogb0272/DEqy5qlPthHgo8yxtrwNrDkqSrrClVqbSMe
p/k2kgPpRTaLBRl1RD99KiBRjMs3Ea3Zl/ezKyctUnhqk22rn79VfzUyhoiLr8fB
d8YOdv3J9HJrLtAotEvexnXNL1R8BdG4zdSq5+pZ7Ymqb/NN6y6InyEOIvpfjFvd
vBjWgYVsAQGzuMfefNZXcKQgp09HBJdVYE3fxzxyjgDV1xqt24RhUj2O5VpHYUFJ
wla8YInrkKT8GHCj1XfKFbZGDUR7eJ7wr5JfYu1XICBRhK5Sa62IgvLi5ryUGKN6
5p5L3XJbd4CCwViCoxItZ41ejPu5njJHKKVgwzeAv/tK55HKtoldzkpBChKLW/ay
o4dW9pnDkJr11r3LFNhpNq5TacmLnWrm0sD9LfcyBMXwOMERX0Xntr4C1CizNNil
7EXkH/DD3t//L+YPStDkW/3L80FuhrWTeJ/xVl6uNaDHU/XH+JAODO5PALGI4eIX
1slenB/TTz3EqAeYUvC5aPo/epF62mjGK4kck3qQ/HpeW3BgyKcQ66mEnUn9bKNh
EwenGYjKq0BQHZ8IKobBWb/cDG4ZXo/WYxV0Ia6aFvzHBlHZPcWUcjxr1K43zvBN
Di7QgIEiXG+P1jEPBOSY7jXQLg+CLKSoTWg6Vbbjw9XnkFdtGawie6WPtAVSKdLo
MB1ujMES905EtKrmHbNEJT8q/KJmkgDaPy+i/Y5fUB2nES6pvrDvlfndIACHtVNc
fE2E10D5h0OGjDKLfMal+PM5+KQ91V0jBRtHltoOJoezo2/BQMqUTb/Wza+obf0C
CjTjGJdO43s69qjc7FTceBsBmd9qIdPWVCzN2Uk45pa7O16rq0PjkWcm6as12prN
e1IXEZ4ZgHeZwoVqlrd0qQwRxQiPLoewH6ifO9DWkpD1DqFPH4+H8FCKGGd3z8uO
stu/VGK6pd5zEPp+pLp9EH4YD9AS1E1SUPIqQxmeEhHKii/OFo0naIbALhSIKY86
GbE9OgWj+Hk4XFiyjYbRLQJsWFQFY9X1EYsm2HE2W1TKi88RNYGLKNT9B6es0YSE
kyXP/TcsRF3bWslKqnTQQUvRJfXFQCKQkg5HnbcongAkFJuYLeitCzp24eHG+NEk
HdYtEb5B7kWUGu1VH0NVotKzunuXmkOxUtyxJTRSM0PJ32W+9iKvylOvg+AR/gJ+
39c/PmJKk9A1RWrHiqXKlXda2ZjLONf+iuf6IDxwlPupireMyXeU/41+sCLQslVE
Rt4DbipfmAzpVCIMib7B1VAWaDUVHSeEpP2yhgPnIcW4kduVzjw4ae/qCDj0054Q
BGOuzDpP/HyYS3gviizLJbbDJVc1oUrUaU24zGl7FKBBudE+6RZZ3OAu+p/YagWw
D7lewfWjgmq6eETfm6rCBxNQQlEQs+eQvJZBafq7I4wrTfwxzwt2aWcDAbB5r53N
DpsSS4ihZ/bmOf5qhQt/6e9r4XJ6vMhDS40l4kSWBUW1EJnxp4Fo6nx523nqXcbT
j1Q/3HLMnQvT/b6wrYSiJBiTFHQrVUvxGUJII20FY7P1jtBnheRZVxwHtslIwx1+
TATGKG677oOt2UNQs3/RM6PHXccSrZ3DlIYj4rlVzd1OrHcOeEFCWjRJqVi6sm0W
Q7+DaRlhr9cywIIdJD1+OufbQF2VtnyeIEF8S5Wza6tIX8Y+i17Myv/nnKE+nLKN
5tJ9Ah6gHgnvFEFdNycmVxaJIZo7F4liCygVKr0hNeHReES1bGOYcH7OrCPaffCM
uq/wuuK6ZtCLgMkKouR3Ep5ZDvlIqTykDpms5moD0AewWSvqfkoR77tBpno+2Z7p
ISeiGNVPOSeuQXlP4oLlgbAr4eQ1C268yGQAyefI9nA48374qbe5+J7CSHeWTWg5
T9zvXUcrhCLc3lssO19A88ZOdAaaxwkWqRynjXTBb3drscoy/9XEqROVR5MtXhjp
13KA3F/bNYHYP3vm1gVK6XDckMb3X7XzD1OOregK5jQWpd3VciBgmI5QwYtzuhaB
Kncs+9RLh9pfqOkSDfSUwVjpAqTe12+CE4BJ5c0VA1LzV5IH+vaYFH83Fko5q4IH
EEwjee4SR7jrKXAs/l5v1xZQ6wuoH56pfGy1XjAIcuR/dbps77ZEIOqwGe6Jd8cn
IXYoEB80aEFOQKDHLYiWwBZsT1ntRkGL2R43Gtav3ksv4OX3+OzpHLjE+uX6R952
2IZUWY5VcaJ+0CJP36zAxXgxT76dC+iT5LYeC6gtYKIuEPlzrmUiHxYGNacsg9U1
AbJ2wAhozN+P8+vojDNTqrFsnutboMsWR/iMq31OJ+Mh0S8uquI6NkrxVNE2mm1f
dprV8/f/73/Eh7hNrjWYkT63bAhsvk3wtRnogciLdqFaubaa7MwUA08XS1viQmR0
O/REO3mrbQoX7Ldlj6w0zDCZDTZnRAFlhY7RxG3OQLIcBfo8Ige7I2po7T75SXqU
apBO/rTEV9ocFjwGMUcKT9Lh2hal4WiMFGRF0+iC3cPNLb3qbzNstbPVgXdwARXw
AJJ5ERcFJ+rCkpiwyyN5soMPMNBIpD/y/R2E9LcsVo9+1GFZ3zqfnzll8UZ59+mD
reiJvV0rLoeG30pIDwvby9DZfq63KnahVWQI1VC4WS6Atj3GPp4v97SpjVGKdwKM
rRYX1inN06tiuHNFhcP69+aOArXt+M/t8TbIr5kBER5DILwiOTEVqNl+wozjvCNU
7q2zrPlpVPADKRJiEbq7zErVBk89W2CkzSaQME2TrP8YgBpSF2GeyrwXkSFcoNTv
sPu8DIGkMCVZN7I3Gi1v/M8nrpPNyYvCR1yZCJGN/ZIcD94/ASbM2Z0KXZ+XQido
ZaBCazcb3V7Z7RzoQVsDY6eWUtD4isajEILhchcewts2g13k2AgKg7pawgXVGdwZ
5zHAYCBUVoJ/lM8CE7GHKV9I7WaoytZ7NIJSooCE4THAX9huV2WOMlOg5DG6Bksh
nkzlx9C5R7IuUL+YYDVSlc9PDv7EcuMN/T3vR37K40bCRarCSbanDLY2YP1jb8SF
xzo4il6aT3IYSR3gjm7GTj7uB5LPBVNgaGKMjHh/dqJ884aC/VEMVQ49RaogCj5u
Yi0lZZ3dsk1suTyKaE1HOPdkKJEBr7IgtCxfFF4pr9kLKR24T4u7BcJaytVjHMAo
MUfl2GcvMXUmGMZY64pqA4f1bGtJX79wQbLBU4HDi7ilcmgFs9eV0hcPk5b/ogHO
yU6JwqtZNtOBcZeMeYLkqLtsz1wQcIVC7GFglli3GFD3EjsZwO66Ii8dttYqNpb0
CbP9lqHw3hLvgNPeyzrvFeE90qeJKGqfHiM3EqwwKCqxWc6XEOKzH5Hnj1RAtZf1
RzmuBLZF/CRBEJA1iBW2/zjMW2TkBIYC4b1XHmw/LK2XNgIoh7Ki9Rrg0sBZ5LsV
MjbJ849mMzrMa+eYYmnM6hwNjwxnBu1syvkrGbLufonteZH6A+RcWM2KdPV3c2nH
pVgleKFxLXbVNKE5vZxTK+f0W/ZrZjO3yox0l1EK1tIOm9X9vsvN1YUOHOyK1Ke0
PsDujfAdJtZYfmdxym3l5SD0l1JeSIoo1PI7k6kVkchM7Po9owWL4rYvlQRYZETW
N7wWpASCLzMZOpUI7M2ck9KXAv0newyg8Oh/mmp9AV7lEsKzDFdnuICH+bl3Y0S2
gJdO6xVWKbe5IOe+/NJowpS7IaWsTpo4wLwGTUtImPMwSxvJnZBFC2d71mOjyVCY
D8/StL6pu0SVYPZ4NugqgwK7UjV1Xx8SJ/8Akcbz9AOG75c8AuAEQHGoAKHRLMw8
Rsg4+h8PhZVIh/n70u2IKC+cIQ8K7s2B1LhbSNz0Ixab7OTw/Lf55eVyGDEBYG6X
OloORsccQPoK8e/4LO28SdZrHYf7jIVk6m1ztmYfdxyRuv1F8726jAAhJ3aZ50D9
53IZsqp0zog/zSJYi7PR+Y0v77002PREujrAQUigaGoRLU752w3sO6JyRs1PAlyE
P6Ohsst4V3ydkTywzldKukH3lUi8IRXl4bCg90t06ynnuCRrvcpfD6zaGN/AMSfy
Qmy8rn+C3mPuaxsAGr9v9xSLKSIinXLDityWyaDqThp7gT04ojMFpTE2UhO+JNjv
HvI07skpjfGQvbmYhDr+8VsaFjL+E7LD9bqCooUin0Bso+fK9boREauzQakXl3az
+rmWyp7D+otKowUd3hGY6uQXEhY+G2+Y6lDr4MZkXqdGn7ZM8NceN9RxqcztQxwE
k8se7Rgbh9yXafWWa5EnBSDDY5Y5BBFucxkof+K3HAmaVpZGrElQ35BgyiRkObfc
Ic3l3/8e4OvYh9zORFfThrwbz5nHUe2TjmOFa9yZ2q7hC0kKn++eR0jM3ExMeGtJ
aHb64p2F4cqAl4yhVUvAejUneRDCbq3EccIvEwvPIduua0yqbowrePKzDwNESIWY
EpEL/FkRwvoWlQSpdeoiW0aQIig7GFCskzx3cLp3rz+zOo7UD/VHGgBAK+bRWwyZ
mCUGcX4QxUZjSiR2a736yHKxxrPVpC9MxzDV01a8NS5n6As99VMJRrLDS7Lhl4kq
LyK3LrcAUzsserseGmHEQ7fJ+q6VXENH+stoI9OoemDUqxTvWucH6wxRQF7VxMuK
+FJuohrMtpnRCD37bqVbEARxN1esg78NBPahtydad33J230u5H4mZOOeZkrSgVpl
E32Zsn4bNoxrxvHxG7BTMwNYABdEiMdSSajuqhB4og9i8X/D0BwMkIp5ANcFCq6G
xaDUFlvtLpq7lCLUNYXhGl4vzZGxK13C9dKycMkPVIyMONW4l0ddJHv29Nb7ksXI
dc/kN9oBL33YvWn4CeNmxxiQpK1hwdASW7fuLyrKVC9jNwecF9AgVW6u057q5ywR
VWaDUCzoW+y6EKA6EpNrz0Ws00vKIqSOyXIpVOKWFfObW9YXIzR6cTeTzAfHfM81
BDWdhNmUGpIPjEhvMltxL5gpNaJ2OhNAtiN0xKFV8OexSPThCqDAZe2mEU3OFvuw
3FGWt9y76UORmz1R05t5HrlDshWlD2RgcK+jV17ngfmzKVQz/4cvlGAiBto30a7I
6gHO0wzgYMg/Tqul4uSP99iDBZk9AZOrMVl+wIJ0y9NqcOQHtjVLVDbVANa1aM6S
94LVK2mc8KAAbxdcdGukf5UnWiZBJMZ+pS8IGu20LvBAVEHGsRZxsh79LglIaV3Z
TNI7lkBaT8028ekWltT6DENPzgchyLeg64helntHjYZVNWgHpTKb7RdWVrZK41nG
5g4gkJTJ5KHzUYgCeBD/I5eQIv3iJ+/CFX84/HoYv112sV5CS9UlbHScxdXzhzzE
Z4uv28oriDT3i4Lt/UwY/yuqnkA5PtLq2zbDg4ppxK6JQ4KnnplWkVxLhmXYqAsF
JskKfDrSMaZFswqWucJkXKj2mqKiTCargt8WJMMlhwoZnYbDT13GBJ23ZmVJ18TO
VfG3Rt/j60QLRa8qptBbcxvBLrTnO9OArGt/w77ieiZuC09mfLh7WrnGnaGs2YzF
NBlYWxpS+p+i/dwsVnYWEkV7rd8q3F9r/+ZS3Z7aY7DspbpNrbXQ9iL9539Y9zct
+V6M0NyUka+fcrQmYPf0OaYYjVuISdDMT6tHRRl0o8xMgy722EU/Xq1wBDZDqRlV
VQ2MskhCZBYfxjkby8zVd1FrK08RQAWjiSdZvTOiHV+xmFmecjhyyh5ECYxKzKnk
ywk4JM49HmmZF/oWHP1/irH9mMaUg1PxhRl/QA//FlcJI6Mz72KsGQHGRYhPjAMw
UAHl3l5uAYBsUq8U21HfMflTw4INQuhJ1oW674OkAKUhTUtJ7nOMxe4DUHznY5dK
9ybk9DllvQPx8Qrej1rdxywtwbyjS2ZjDIR0dHOcV4mBefDV7aPOePSS9sVNUO7b
Bs0KXN6sJ0uLqkjiqn9ft7yY9T4oP9IVVzpvrI7jtsIo7/2Z/rDP/TgK417YgnG/
UdIIcA5mMg4QFRybuIhD9p6SStgm+96rlQrPpg8jsEcJ0+EJw1ZLvGgUT0a5Mf+1
r9YZZjHacwQExNE2OYDfGLNA7IHnGmQ4uhJNjMetqXWkiaBGwkvhy9lXvu/CYo27
ki/lQeKLH5xElxDcWSwF9jIa8IkH+lgxg75QUP2V1aJ6r9miZECNenkO1rqaOb+v
9ZthMX5PFGfuBTbqwFz/eKZfVp8f4JJ73Z5exmXX2FZkKmqweEeIIEQnKh8w+nPP
fu0UA+7EvaKPaDTe5pk1tR61/o4hi9A02XrvJJymqfMR579kWa202BGU+oWZmODL
/3ydx52nUyqdGZ1rgdjgn3ZvOHwetShDdQ8ExdsFz+D0Jq9Jntx0QVHWtNAnsVPl
++ZzXZPjo0xNbK+cDcko0Gvg2UMTixvfgMINZtbqNZBZdgRcm2dl/2BRMLXwz/TM
1k5gYWBKmpH4SCTZ1Xj/Atz6znaW/VSpiRO3RjYgOG2OSjOlaniSvBXlOSPGn6HE
BXqfNBto66tuSz/uxfQ9TkfufKASiXfmXwyfqsrZSpfl3aPuV6R0uWPNw1ij+rY2
ank6DJHwE3hrSCoXuHxSgwPc8MT1XwXK/lFRXJ89/aVApKqyjfCz7zZbaQnuBO7K
yr4MhDC03CSyYKeGmp2INflyUQX7lsQCnZO9YoGr7/JkXsxPTnwg/huou0XdpoA5
mkiJ7SSDSdTPPRu8ZQ7dqODZF2z5sI76vy6D27QBTATxrh9zXJUQyzalnfog+ses
adTDg5AWj3J7mXHWI7zoSvTRg+OmkN2rPlY+x6sNRaNhXgnTwApiZC2zC+9DmTB8
AdU0MP2vEM/LYfiHBamAZjrVA4llMJjW4KXGc/qBbaghcP5oXNykbmvurzRvILL1
7StPxMO3z2mbssfxsgiqM3cg4Q9Hy6rdgmOe25Z1VxQnM/JHpKSM1/lmAxMga4oj
/WAkoa8JoZt1kiS46fO9Khy9wmnbrd9QOm3OWx84edqN07ZUhMeaKsJ7Jc+zuHAs
voqi0koUgF6dnh2YhRRzN77pLloez4oIQv4tXmQ2RlPfOChXF6xNq2LMbtXLXJcE
3rnyNmDn4y7mWtDkz2EF2iXtxCEXSeY+7gat7Dg/ok6vWPTwDaKTAaqy6KHzJ/m5
/pzFlbzCWWAnvYsaL9OPUZ/NnP0En9yzpaa2kLgkPny6WqmJV1db64bMrARQERlN
CjblL0U4ZPnlIHZSo9L/5YtwNc2VZWKXc0DBFW0bso/X8NzdpmWOPSkVAa5+HhL2
Nf+QugRugApN337czfqQlgqScKTQYVT+qWualDci/kg1Yq7mjqhOj2cIpuOpkeG1
32FC0szHxjID8Ftf0hJffqvAXTdRXhpPAgkyg6m5QCBnaLM1fZX/baeW3Vvxmpu9
f210Gw0gB0p1sPmUHPeXqN2ztk+pI9lFNPLLf/6XPd6xo+eHzHa4ePnyDbKRqEua
DCqkPgphZ9oGcAt7ZgSE8mdjypK2W32GYlnHPT4bJZKNPzO86oHVgHZOONu3UO7R
spHkqanZUhrEsZkYcWotYoOnnAWYzvGdvCPOy1PkImZ01eTa3vHuhpkh2koJQpmA
LRd9r0085aS4AW/lcpL9J2kS/RWZDQo7pI/I8CgAaeyeRQfqCtKG6hcsCr9TWlc5
0eRN7KNanQfg8vfmyu6WZSLtF5oOOX3nC/cImYcHisFe8poEcI1EpTubjLo8HtKF
xk7FcFCl/BubnpmvVQcU0gZaAJzAs0+cgJK0yuOL9b5pM00KJn/u3p4SIOqKevmY
Uh6W8zT19Zcun8QvvWsz1c1rWlXBgpfQAPK69YY0Dld8mJNCVqSfyyf6FfphTY3F
WG8HPVOHneZz89+rYskocU1XtKJMG6YFNbK6jrSGOSM1Xmp3QwymVHmTyU3ktB6F
kO5gyWGUAaBNaEnv0OufBD+amIQc85UzJp0pi2gyV8artPerIlvm++CtcBtVZh+G
Sbk0b4Bi5W6NH+Uwn+IL8rj+rg3378mpbt+jEplaxeuxT3HLPjUP2Gtk7GPDZcbF
8xpE+cuK5TJBL497RlWzDMA41zJlu24hryfHcPceTz0zeqzGvOyEAcAnqxNDB0KA
caOsRjytFRue64XPzXH0cgl9loWQ/Bzexov8hiF2fTrv2uvHxxBs4DnskRqvXTnS
FAoS6lo4Ctvu844tjbn6VhZjbg+HLnChNtVzFIuRFWr7L8bcA1C5kyFSXSHqzi2g
Kikj+NlqiGy7m/JXqBDJXAtplBN5BBgn5MEMaYkluCmNlzUJqe395uMKdU3SYB/2
h7L010b3cdGRwySdJr25b499jcrFn83wCK4YGpsadRIAIAEUiYktW/lcp2ImnyMO
OQjDIzXBb3ppqv9lAwQz4ZLHeU1oYot4q6XcRoCJ2Tjx5gUSsmMzevPn04V3iUbS
QOQvws0kM9/OnG1uIrrj+NzAT238d3Ly+QU8S23nUFh3sAXf0XlAmlwmk6XDivHP
YEYs9jxu6U2JCuM8VDABgeCFchh1rUdIR8NjkIaYyutzan7XibEeBs7qwu6p2CmJ
RV7LX/nXjlO1z6hnvm5hBjgW151IxjSZoeT/B9SVRxqvEPx71C3zvj9A7Spvgebr
GomUr8Ot1E8a55ELwSug1tdWaeD0emeR+GAiA2PrInjtvNMLJmJ3TW56RjmxkPF0
oH8vcsdrrepQ/XiqNgnDJ/yUuwio5jplarHefqYFurlEhssZ2OC7iM8A0yZbmXtQ
P/M2VbI1i5UkljEC3Kxn87FTyP/8KhSKIdCaDbHWJww2aEvdXhinexDm0wUmEX0I
ob6f9eR4bWZJVSOR6i+PrHPUnU+4Wt5Fx1+i14X8vtYesi8/tegrZo5R/uk8QALt
uziMqW8BvLz2IgzHZbZ/Ya37hQ12IdJi4XUKDTodfyvUpKNr+qj8srOHn++L3Get
sinuobt9Xb0OnVzIIkHAnjLIPXJJEOQHQPAIkRun1Xpb4Hm7nC+qhRG1AMWv6ZcD
ukQVjMQ6eGxvKga6Ye/IqTEENlD5CRWWFtMbLhYLvFk37Hdb1OV5lQDEt7xCa5K/
8m/Sl89/J7+HIDjxKvxBaVT8lHxnwTH/ormXqh2cFQ1jgKcZMqlnsF0HjxSTZy4T
qaapCtWyoMofWQPN8GVAg1vV3llvTvPdX+HOE8fIvV+SMtawgFpHD31jAaevAX22
Ho9BcSM80rUwGhTJJ/hm0to6qxcypT34WJ5CsUZIgSY3Qw33xlLb+Lc6+Z8p8olk
HM4t11nN2W0/oavTKQxPXMDm0S8kQ6a4v8DeiMrBzhNUMjBLulyav4b5GXcTVHJx
aKPQfxYhQP01E0Mc1ZNHSCxfPLEW3C3pORJQBhazM2px7NEbZByIsR9DX2Qc8+O6
1ud5DkuOH43vEjKhn6q23RjE9yfuCudxixyXpi1Xi0HhuBWAQA8pi2ct8vPyYD/d
tPnpGEcfXF6if1LzOSjbefygoa1h25aWAN8fdbrN/qLtPlL9lAHSnNdh9zzHkFaZ
/c4JZ/frQQRcAdS7RvRY7dZNDzsIp6zJgDZNdfeXKi+ly2JB4+EJG4nOW+5rhjmi
XXG7Kaump+tugjF8XCknPxXsJGnbvdWkPbiXiy7VocFf1OUYBLRwZekhix6MIX6v
BPSotaBV0N6xAsFjB/bxZtXqIGxMcxyi4lVvZSyKraGnHHZH6FVWlGXl5b/SvmOW
QYvZDT0JH/YZPBfvB7ZzNIjAcGGcZh+WDHzrlofCWedmk5KAZcxPDcA1At/A4eoh
VCOo/USX0cDWopgcCjurXcM4IY529RzApe3wLAmZlGM16NLt3GDqRYgXCymIqLNI
5rua/cUoaw3ABog1OSCsvAFNiEUJ+77VUI0NxC7kIjRBPrA5pUVEUffYMrkQtrjD
WFF7jlsQgT2WGaak+hQSYnt2jFT9DfG6otwq5KGDVpS0jbO5xHM8AORrWz64Uszl
W/g9rr7rEWBVC8pLZjm+Y/q3DZH9JHWlybjqXRHk4BIvyKU/Ucq4XIxBzxCEnQZ3
hd58p/2VtdearIJOmKM5QJE7mltMRMyEowIcgLtHv50zGrEQf1CWQSerhcNdbOvw
zQxnWrgrGujR5Xeak+98Lp3o5x506/U6s4pypVwjQFi8Hjm3Kvl4edfwNF4IdwLI
e+ES7wG5hkewAhhtWwMZg0X4pbbuRBk0FY7Y9ZOKWpqTPK68BtfcOS/MsYdXGotM
j2esW6WihR4QeGYyQlbMwps3oqjLZY9FYyyceBsx1e+SlDvFLrHvgBX6WKuPUSaS
+U8GYBcTTN6PFUCp3ai4XeLyER77Mdzj2VSluc+HqRWKmkzn1aJ/Z6uTmUT91Nh6
m4utV1wqDBxFl1J2WpEYx4EJqlYFn6l+FaYMukiv5zJL02WsscYJFxdAF7wYjBV2
3FIO5DEhtqq7jIklJXQREcfu00BMcR7nSqGDTSXWDZcYX6iH2OnzZ6igWfUovOFf
NU0O4k/grJxNI6ZCscc25isgwkMEQ8pQax5XXxjhzp5DAikOK2/BOcA8Uiy/C5CW
yEyDObFd2tLgByTJrH2+LpY2EFMfECdreveNAnRHh+XB6q0rdv0ejiiS6SxmpUb8
q0NJq8hQFdjjAb+d9VAxH52vwrvwNqfHwIRg3+rMas9xkRB063tc0sLg2rME+kii
OlDfssG5ePCSmXBMlYooqbXyoi0djVF9Mmp+aljPtlFEjE9ozyiNaUDHOsD7DoO+
qJWNZmBKodX74HROyadPYC3tHt0vNKMM0SWKIUjjsIZkMs7pZhRZBiYzgIux/f6c
HMNRPJWoCeyzKs8XdJJr5zLJtvoM/3cz0PzIBl6wQpU/yXmEB59yCnVPIflJ1OHM
o6hQ56/ZtKAbO/XoeXBHlB4D2zPcB2L1sVhabo8fnZ6zYXqjtv2j09f71Ac6eqLF
BvPV1hT6gGnrdYDr/m3OGS8DVPKkm6/4DnFbZxzjXIflXhwbBq9xh97rmU8FC1Fj
AwX/5W1A4FdOBaCMJMZ1FOlJ3qEw/AZcIfLotU5+y5CLXKee5orxQVqPvu2myZbB
Hrf1/FgNekKOypMduZ7FfgfLCgoHMI1WFhuqPFIjHV3CgAINaLhacm4pAJAFM6Ie
9f4NfVEdGgPUyTT4BMB8X3v06MVTku1zxiT6Y5m8b0gbLgqapw7ykOHW7ccQby4E
eVP871IGuSJsebqtDiK5gDHoUDbZSS+Iie/0Mb6l/D4FO+2AjsigGpwJYRdkmta9
XSpazcmNPtsRKRWrAHvFcfVJcNdEOt5W7Ug4S8gnidPf6On07g8YUG+ygkW9xEnT
PP2Be/dbHBN3kJa30fhxnUfNhw3EZJH5dkGZBVTu1NemzODKbph7whGQ+6PZk4rc
VNE2tEP/4Kqzkkxs1tP+9MaZVDW4S2kFlvgkDB8fk8WEUwqZCxOjh6ze/hYaH+Zh
ccTytVBtPo3Yqd+peOg9Tx6qq/EWFf5idVTNfuQxUvbSHLiMAL8xiZj93G7UTg10
OnDRzaggMJ3cw2u0oSd6pkn961nkpoKKP86gyHCf0eJkuBYoXGUgU57xG/HrH9mJ
dxsNi3tr6Fu2qpQ/zD7KEeg+iN++yTW3Oml4O0UK2abp8/6E5RniJ3o+Ki5s9xbu
VNvdVMLnmNS4C7f+E02cw1/wxgHXLR51UEzTrkAU55U5nSByUm+xjeuxKecoS/3m
9moj4m449KuaSu2yZf2wStB5BVYlcw9ldePLAceop5Uer2G5a/FhCHHO/OOKIILr
4KDKInVUe6QQLVjb0p42Mrr4jyGjKmseE5j0xAxC/krqUXFtjhLmPC6Fo9R12zNp
hZ4tz8a283Nqm+73h2Cn1akdMQuLsyYVLSN46qr9xkMd4pf8feAQtzhvj6AwfQCA
Q1/KfBJ412R7PdnY5D59oGpddOrp/qIqAhLINFDQ0wYLfqLczfO/v5D7Jvl6QEn2
IrsGiNCvU4lMABKXCTJAXwjfvZ92eHjCksGYQHg2sVx5BxoTV/XXV+j0ydlC/Z93
eq4ILqrZ39na27aPLfO1e6EZhJb70RNa/gndWCEXtUYrpReNS2hYzstwo5VzB/p3
ukMO76SoXIYwb7EsK6CnJo7eOAQeWlmHk7mIIDBQvDJid0LAJL19fA8EJPmSjETh
P7H2kLt7OgrmpITFbX46glmN50p/G28BSFKJEVXsXLagrWoR12h0nvYXe40uDLRX
LEEjjh3lxGSdst4wnUABXCCsLGDjsC9GJUYuQIMWi2PD+0SfyMq43b6yGD2/xmyz
lOcY3o0ALIs8V/x/fjYOJjuIfefrlSManeou8mo/dQucAr5TpdDC2m8Ly1ntZC/t
1TkS0KueJXN88dHM7ee0JKjrtGxqlC9uPwT2WavVVSCkA9ZhBjusqY7g+oVIDlBv
r5PjkvjckPScUWdFcmaQt9GdkoBVaPRCAT3MVbEox5yIncepz9HxHkSrr4geXlZB
BX7jZdpq52YFu9LmzM6BqCOQzr+yjKZFwrhzhZJhVT85RCpHSdEpOeXeT2QHpIQX
XSeQ9U6tFGdE0tWVov7lQscZ5+outiswIPaT4d+rJD3ND0zhX960zalmh/0QjsOp
gA8yemawJ32QtIY6i3pFP2+QPT8Zft9qJpBmsK3albVfKlHun1ANrjOfsbegcTG3
HeyK1FGaOUGnueivgpNlg+iWCmW5b9O7hZcXdx2IIe0Le0qUL/4mt8T2ozFWrTPl
8xQFHDnxfhEVZMD0gI/ke+jo2tqEFNWTH1O9qTO5v6HWTiKLUXqHSoSQN1vjyO8T
3xVphRX2g288GQCr/LFjVPF6PFxmQWPBIVLUW33Z7IOJoigkVwV8aHMw/s2EZhqw
6r9G6aZh4OYNgb0c2/nXSbfYfpEkWxFymyQmHtyExaEkxoG+nsHFrUFV8YIw3+rm
j+O0c+i+fK6YTKckJt/+TNmO0gJg3dFfarB2vtyhmQe4egZSlnX3ETmA3m1BzHEC
r1xeAz2RSps72HP9GglQw2sDfMzeF6TKoMjjbxFq0ZCMobGLxVR8XOBB6yVxNyaw
4O6HeG6rMJPu1LIX1+WeaVG+SCBHQo0lfhmUBnbQTGrRuKcMeBkjTwLkQqK2+6Oz
4L0W3cPTxYX0g8fxUuj7AdHr1bIfHTn0be1e+JLWAFyYQ5N4hqcd7g3QHZozvsIO
xqrr3Ug6HeSzfahiD2QKbSxpkw4aotaHybdy4F1eur651PHB+xDBR5Gh/aNEWTty
7D/Vkvc9xuqTC36pv/SGLm/JzPTtuIUYyNdqriNOWX2f+WhOpZmRyplj+Htjnu4f
V+xO8baIcv2vrJUqcbSEGFfuXyBCqPmaVs2Y2sh6PFxhm8qSOGqpTSW247Mp+Aty
Onh3+xKh9YdKarkS3U8Elhz/eZtbpl3/9lQSFCx8NSn3sSPyVrUQL6DEIx19meqe
NVSfFBUHqRaOfrF1d3nBvH4QppbZKXHZF2vw26vN56Td8iypbGLnWGD8v4/hdFJx
TIqcQLWSAssPj6njXo3IzksatYIwg+095Gn9reYiQQMgcLny2y0rjutc/lOcri5p
4oOB97mFLTl3rv/MG4YwJz0aJ4nRUjqgq0bBpJu8BvZog4HewjK7aQHzThZFYQZt
G/9l0gh0L4LX9rH+g/xuyKfD4GThYZXy3A4Yfs0GhvFPpfocH6vOetuNTAD7ZMyh
Wp5kewyO9kDnvCkiwTU82VhRVuhxBzkW9Asyqv621ilLBaGgp6/lnBJsLw9TsTMU
RFr9LTpu5jeHju1jYMzvAugzqjWqMkC4Ws5H84PQtNM2UBwSNbLmZCmTMfApPIA7
Kz5/wfk/WQYOJ/kGrwdfX+sD3d+9StyDwUAQWXpsW5zjoXkaapzUgpdOCn4DB1p1
eNdG/LrfQiAEAjm0zDhy16IaBWXkHjSu2109QFh86tYMmVPKrA278BtojS/X2KZC
WwD4hA19jV92mm+L1Td49nlGd7lbdKtD/20/Z4SxZgB72Qhnz3rbUN9TMexhRUMN
6oczBdVKeN0YWrwyG2oqJZeKaL1wwgs/5wQEIBrRbCbZjCfTes+INdYfvv4pitKq
+94QZvpF+eRY6nbabPOiC8+8JtNOEvrtZsyRsURtp5qMQM/ZCRV3lwmjztNKTxkB
PYYMMGbMpWQb+ZgouovD9zfqt6B2JuSc49bN5/QwOUdmy53i1kZpU2x5zeY7/Wsk
9r3tvfioymwScqPlBqEVprwQgsh4pfEPf0XbzYv3rYv27RF/9/ugAGvU8Srdj0N3
NWixmkhrRpnwzwP977bzvCL3PB66E/nX62zrm8E3GjL9pkhCiOEn3xiVE8n2HgBl
TEe4uqzDhzYbGFe6fCiqKhOvuXIZrTBySLnwjBvQURgIu068rp/ZHp/BoIOqUlUo
sYcGfoS4jOeAcX7DFPtXvlYSlu8m+c3D4S1Kjo31277bnNefSC9r5pjiZVTCtTTZ
0Pu3MH6GjP9ajbeQ0GIsYxhiHWjrfV81ufWAQsj24lKwYQ8KKFrakaaIxsoOk1NT
xg4PFYwd68VfygKSrFAiyWPvehzoleBLaPeM4MehajtzSywx3UHyRF7nw5BHpYUj
SRK1WIAhz0Fdu1wxQ/eI3N1Se1qTlAOW/rKtuETETul4Q45hu8tI8naQhWWlq/QP
i+KblmxRjCBawGBQoplAULvGadfKFmXtyVewShkaLKwfLws6xHmo62IfnXZk5e7t
amCfcnEUEnEU6gYRab4p3/lccGg+B+DpdVuLDvvdOgD89InoHPSf7WgkA+/ZVV3X
DOBA2+C75lBPg3zSoYHjVtqWEOwU0BSxxWcwR7UK5/1sCvsTvPA3ZLNy7nej/oDs
LjbAgoXt8F7JJEGWV3La8VH34HHR8DS+/g2yvFxpumUlRPOFXoTyDqzwEMMyIoS+
1b30w9DiIPz3SHeDa22qlfX6Ajj7wx+4XmnLTnx+2FOTRgzgdk7Or9dgQzsU16nT
xqgDiLC/NPcpUMYQiEhBlnF7qKJ0fu1se/W+3ITYFX8TPmms0gCA8LREe/ESNPzA
GLl1CP4X2ulz9+bco46sDhmkwd0pZIuOZrFmWn/0SZEdLnJB3oF3CSuZT+xjIRj5
qZv8WN5HM+cuPiEIxAmelKQOASHTeX7w/LZm45dbzICaLwSTQslehWYy0OBfkGYN
hquivqCLTc4ZTD/yWqVhEjLSIhnzSwBrys7gnDuUBs0THMar0cpZTWg5wGP7O0Br
jhZhnYLRu1h+bk+vBMUPNkgmBCMRbYlr+ffsyguIrdonAGWACMmo2dEvWQZmpX0J
5eQ1ABA53QA9j5+hQ9sojlILnVtgqzrJtpKeKck6lych86b6bgES4QsZvaWXuPuK
yMWq/TyNKiG+r0d6zwZrh+gHJVpAVUkvSelNBtUG9Gsn2AMf0eodopo4SpvsJAmz
T9v5mgNXJRJ5I/6ES57o3k2ZdMal2QAlLd8t1zNazddJa4pL9vLlT4m6/+j4+adK
k6WQw+htdFMsvMAzYGs8VU3LvCjF1xwLsY3eAy00538Ub4neSHUqMdHsBqYaJQn0
y+AOEBhovGy9s2F9RrHpQ4/QncVIeQUFDt9z7Sgkzwy8kSz9cuIFRm7brOQJGNzn
+pgo4x6DtG6ABJGx5ZexN10UGW1Oh5fPuZYgwsf6ruJCKyH1eGN4yeoyn2X2YCZP
tCd939UCMbK1sum+hDo3JEeEvemLgw1kEKILgjDcUkcC5sF5oSavNTEbS1wlEScQ
Ou8NjWfQIjYJVzQlYbc4N/M7aj/ZH+erdGH0R87c4cUpi8Lc6UocakmcYXOAEu8j
IXFjZnzWj4llmwBI1WtX/hyyqzAuWb2GhmDejH/3jXswU7fEO9KkZpU9BK/yAocl
m+vAAp6p+0WCHyWKgZDGO9wCWZBEQra5cH5k0z8oJSsnNQkz5hcOo5YD9JjswgN1
igtjpu399tYHbfNnu5ljynm3sDVqSCjZfczZG7OQ7u4+3lHyJgPIeYq2J6mI4QkN
xo2FROBPPI7NBZqC8DJAgklTzvbaV7NletyyqcUtQn7YRUcYrJYVrpt3Cp7KySOt
U4l7YmriWBH41ok2Ls4cIK86PWNCjxw4KcPbHOMIWCzaNgopI3Dx/P3/l8zwqrqs
6DOy6Y4EZHYmgEPSjMzSGQ79ozFZUSG5oIN1xW1apHoSiBuH2Fy/jVBrsoOOLX2R
A+c9ji16S6OEQpbXyJrmj2rbeZSvl8kWfKggZknYzJk1LyYTQqUkl91EayDXRz5B
Jv5+v9bqo4RuPZ4HdqRupmIkw9OD5RZ0UvCqcyCZN5TuDVmoqRAgjre2Nb15hLUI
/ReLQGhh53OCd9yy93/ITkJbIvqiiA7Q/T7rKkYcmrNBy11gsz9reuYPp0KXoxyG
TOVrpK3otb1Y8tigbXHU1E09eu+tzcTUVJT0BNqApdcIXRzc5WoqA0uQx/sviBFx
b0wgaRh6RxSUaQ+aNjN+vygm6vKkaIud+/yZKs9FCsfnyAkM1oaMTlwE44FN1EJC
2sk9zayikDcBBnD9vWDzh2YlBc2e4zN6JpCpylAzLisLBK/4encR5HL1VQjKtc4c
SRum52xtAUyRHOQgwnZ9xcMl7DavDVIRTorOc+lYOVwJEQDbcFoq7pkCNEYYDmOH
1+4cSnSGVErzlOfCXcqEtC2qqeE3KIEfU4Pr2KybPJ37we0xwgqWqtrl1+XPVjLm
jtuJggwpHkaS4xMsWma5TRxRp0PRthNmSxwi2FLarLY67kjlpr+jJnoebjW/2pwH
hbQ4+wp6CSYfvK482X26IrI1H8HmyigXsYBgVt9s1NCmQysewq7aRbSPNvk8z0PK
bv13/HU2PUC3ezY2+nFuo7nt42QgDPenl0ur9jvqCh1Weh1b6VtcrNfvhHXGa3Vj
/HF+GXQVYXc/Dbh1qQ9K3bFLre+jZFH8wCKw/lsgjK9vtBrGgT+XU840cqMi5qbZ
xfv9F0xnA0dIhg1qJhiqVCXAXIyqpnu7Sfuf349dVkQNX3NzttSX9Ap36hVci/jY
1LqKyo+8bUcFPYtW7pn91rG21MOQJ9iZK0ZtK+gjUcOiFbQMr9wsUAn3SjnL9vWV
CatIVB19H5b5kGmtytVbnzBlJ9VbPR/pBm9TuUAbDxIMvk6voGmn9bu2wFM1IQhn
GnjMYNAmJmVkdH5X8H8PdXGMKi1NnWv2XNNiZXHsbKYR3EEKJDp6oR+fcgaUraOa
1knHqnYn0az9GM6YfEhUBUXibeSiVRazZfjUghQx+jLXsr/9tjm92Hy5RANilYoA
HkS4Zojgghh7V8Sp8RgcIrUTx5lixxGhJtMXiFQBKXO4NZJY4TbER1Nl/3Dpd5ad
H//WtkoZmdSQ5UrffDy1/9FOTQ6F0XnJfCfjCb5jjoiuI3Swo8sfzgvFrfNhbPBy
7qS5XTFOBwwjI/EbPFn7kPry1O7sGMBZ217DgrbxUFyY9k0V5j0tRi1C3i2Ieult
j8VFN2NsYJUYcOj68VwUwHMiytfPkj+NdGwfcbxZpkqnb6ODFNxKtv2rFWSrL+mn
r9J/lZ+NS7pI3qTZGiFs8wV41TjgL5DG3m91EjAMxnlqQFJpTqtGuPd2bXUwBH0a
aOc6m/kSDOT8vyceN4z4ahe70gVUrLhtgrAmtN+Ir1EayEv7wCPHwaLGvzT8Vl5c
O7qx2PZylSJLuRaFc3oBO8spa0Ph2ywjd1woqzz7CReANtUEh4D/9FmD39KZwCiZ
xD2ev9RbOFL9n5F2GBY/P7QJwHRd4/owXJWMzK5m0t0WqSBHDhgdiIJ+5QJj6Mfm
/6CnR+ksPnOdM7a6AUWC/zkPkNh7XNuM4a5zZRT8lJldIYO/dswsh5knyNmzAcH8
7gR0GzoeNoO3sHhMTUvxE91+SwLLg6ox9r4qLGmdd/I6jyGGd70VoD413jLnopNc
Fq7w3mxrw2ltNOGY+sakqi06dW9dEbKx4BnGCkCIWtNOtegjzjK1bp0utInCP65c
AHJmBRCN0xw8glw+DhffS/+nh1SfuD0Cwt2dz13p/XXBRpA50la+P3aoJ/v1Pv2l
vQA/am2cba5HXJTWcmYgx0tHUDzePHBnVJDCZOoG27Em4z+nl9h8UL8Mbk4saVA1
gkaW1R88sNh1oW5bnFKCsSwJNDJ5j3XDBRsY40Mp5GKYXFUB5J6KmaTnQxWV3Hc2
K34KsbAjpMFhpBjYfchRwhTYCU3v+zR/HmAso8GapawVZagyMX/3avTUm2l1vyb6
GK2qVgWj+bhBRa0iWYT/ZKAhSzdk4a0uHFh6J1ezWDaWELMikUedQ/R1mCpN213x
9Fg2RhPF3r9UrBiVyrelTWaNJGP15zLIif/im4r1Fypxv/OWfme+xUgEI7oXu3dS
US5vu01TIlvEqXClKQ3IYZtUoG4gvnbsCFr55S1LH45+PlFaMSiPGg2fw67zQj5g
2KG8JnEDGAqwbrGLmFrgAKbb6FinxCN8Xm1Dn5b0NziPNwWBPRjY4Vt1fkKtyK4R
C553f6y6hlbkK0eg2b7a5T3fLTTG68BNoCT8BMuEH3zB7XSMmGKQZ24pHbQzsnE3
pY47xSBljAG8fjrkfG39dpEgDu2AxxksHnGQUH40nfuIXnXXmZufOfBslancix2I
fMdFAQS8lSMDc2fG8w1fsC573K+X1nJFqIPjvAtGbSWaMOncMxU0uzwZDi4SUZ1R
nM3r+HyJvxnJmpx72vZe1gS2ysf9iwv4d1tXiM8l3LqBj1JYPQ6+mWJXgISvcFn1
A+9UbUdl3XdlLvRwcrhNMIfgqpiOVCB3ciojglgnwRDzer+wcm87PagQX+8eCcXy
Byw1tXitxEfGFylUNen0ydsnurm2CMsKmO+w0F8qjEusuO/zn5YPPw6eEbWqPq2K
BLQWsmaKLQGnTf062lSmzAJtmadIOk554tmphm+JiCsKoe4/U5LPauuGTtZprY6d
C4cWIRP4LzRaA4LmEkqfQMTr8NmJI2/64xZAzNmGIBF6OF9tA9UPPXIcJbRaAIjm
rIn/yQUc3XtvGae9HjrMpoHY+8gVglGmlmGwPZFi1IeofsszWU54Bb7w2rqHDpCe
jdPM1jBceoKfkNvuMLFT2ZMcoVHP7j1qAQliglNp5KJtI0rADdMP3AkREHSgq2+6
j0UxFOGoyE7RQ9bnFH7tfHrrDz3r6ABOZtFyvjW0AdIStvLgzstPYvOcwBDJn2pc
AQ5vvNxEOq+kNPCiFjm3Rfu8j4pIqL8IZRIe8PiBD6rLE5dlI70ye1W5yRKhV6nM
V+iyLMNGf1ityP7nDiCYnsJPXHcrZC/qgmIL8B68NFL6A6DuVGKyT0bk04pnRa1x
u7GR5420q6hGctKbBGrBozQlD4h93r0MMALAVMt6InU1d8gkGyHuP9AG8EZJI3yx
ZE6uioh1XqT0+FkBPHGaY77qdiDjKlZPOZsfJPKeCjjVoOgMIf7YN7XbQ+EwDY4C
6S6J4LHxASr3MknXq3E2z5aTHQGMSkYMnJ33R2aIaqQ0e1uZZPrD+GfuqqgVFicW
lHjvY2IuwOU04uBzRtZ6hRt+k88SvFJPpA0C7JzRMZexE/Wih/yatGpLqyGDl+f6
Em8yZOIdhlHslgJnUe8yNOOAGkVP2vwEhAzen4ztcNmWD0YGivHCm3HsKloc8Tdh
wjUaN3vgb5DfWsYmD6bqMrotqbeON8EFs4GInVDFD/YL7G7qCoMsfCfGC3cQzPta
eIbBeB6CnVmLPlvFOw4me2qZr47mll+jezLPI3nWA5y6504NSnwYyzb9BcMNk52y
EpeaEYOhIH/Gx5MsCWwP1Wwydn1oXZRgYgUSoFf1jRL2w2WwLzfIFDmy9l0lVR53
RbqJ5IE0RzNvh/+KJ5Fr0OCOjQU9NGt3/qkd+PtJBCTW3GoJ3FHytxj1aW3Kgldh
FGxNlzdFwMy5vY2I2EcR5Nk4esXUN0SeB9pPfpVH498FDUr8/B4n7Mw8LjwxK2o0
aXDcGbAeSeONZauDEtMsNjUviO8fUdoP6ED6Ptcsr5TO6/2xX8Sn5RJQ57xqgVMJ
SkP+P8ux2tG1Lg3bh7buNeLMbk2Et2wAVmLLgGSTZu8mxPtrhtUp2WWV3p094HPu
6Hndwy9R7ep4kg1RKWSN7jrmgSfvebeK6zhPbiwo/EF+7+iyFUJWRxrbLCsFhT/9
XHF8gHbjfK/ePlGxHypo5PtKP3XsTtF8gYM34wMZuepo0pQ9H3JNkyMPX12Gj7N1
yZOk/q3FbG2cmB48zMkNf0H0yrCKw2thHBHCOdYrOHDy0cAlPqGZ7Skbdu/Av+ou
FZlSNwBAzPo4M5d79iaVoxcozyr/a29ieCfd+JNvYT689TdnBH+/x0c4u6Cul7IB
71BgEEUo0UHe6s2pn2BkjqTVZlIGzskM7syuSq/l1OwGwQ34JHPUvoF/mE7YymwA
2e68OrT9MwUHxEh+EwPzX76Mu/Ywn44R20SpMIAUL2wf+AGF7w7fMO6p9S9Qfd7v
jTXbzfEe9t05FTzRm8yopeNOwcEIATziBv1NmxkFvJ2K+RemyMfPvoGsA8NDq+5A
00lMM79tUDyLK76LlzZNOUs7dYu6KE4FyDax8NnyJ4fAtye9Ye6GglHnzMQ+uEet
QzqVXEWjLMsXXvzkyVl8o3/U2IunkSSvd5/xVqGZNMrY38weRLlboIFKymX+Zy7P
UnCwT8qwKANKjApAJdlaG2xOFR2TkwbJdLNBHgtw3ZzimZJwaT/tWMUY0OQ2ML44
gDYgZR9rLj52rkLlBR0a4eBajDhdbXBtK/OGWOCsgwIm8C+v1XJSB6lmngD3gWMd
lxh40np4ZV5Wda99tE24J0gKnEwvFcCyZV+CzbI9B7ZuO0lBgmusBMx88HaO0XV4
bDdW9JFxjstNlXtvEUCSO/IUDuYyeYeW6BiSZuadbic9LMNB6gBsmIAtBtw9p2Ue
0NG1foT7YI3CeyRnYYBfYLKm8IbxVnkSid4GX1YpPlwd6qQAe6dV0bhOFLdsVNvn
P/5sfu+09sKHETrJaunxlPSvqkCMvyNChPJPnWsrz/cj99EpQlQqWdJUrqdt7IjO
GRkAQSNBVRNwlJkAQYTgPm/Cbaw3F5cHaS47vmtv0C6SDlUcZxNcB+thGT+mkNxt
JQZP6vuxN4RqYsmd5u/hPhXE6LwE4bSjplBK01fMK6SBsscp4Ma4FuXuXUmFh1jm
JHeff9t+3x9bhVsJJEmLhpIIN0o8xLQ7yCM/UuNWVtbJcfv/i64pocrXPw2S8Wd6
YvhrNSaDtpnhazAu0hZzlM9nKJVDXwYhi1Uxjl0Spxtp+v+eu642l+Lma1E8JBhy
lhqW8J+BagAQMIjJhQDL2y/UZzny/0uB9J/wt6haX7TF87ubfJSSx/KfkiYyxcku
oi0mq6xJSJNrCPZItcTd6ttOKr2IMjkiHkFFBs5GfssipmWWjccFErofLtNEDkIx
9oVXZoWZH56PhFRx2gjKJ+VUvqcmukaRV4RHloZm+w7Tmyby7iuvzqSpCzZXpJkt
w89GN0E9Avr8w6UXD8sV8eoTNoYop1SKhn3Kp8LrRzv9n9e7tBPYO8YkUZq/7UkU
1xh/HnnmfS2W9FMo70XM32U8tnTmgqbbDNTC/mIqVl6UXB8TQz0H3htif3MC/f1u
dcjp9Ar6g3Xdbycxea8M4fn1C05t/TmRZorsGcMCWrOoknoFDl7CtGiPXAZbLqVf
dCPTVBJfOrfVSDwTCGR/rMHrCB/Iv4CsfKBAPnpk1PhSoLaaGFNvopP30q3gJXG8
EyERUNIYotnD08N1vlXQ9MZYct2k0vvdAOHrRzo7Pf3KTyHvLTnphFXlYcfJs5/0
UyKNQ5bVY0vS2rmf4FVdQ6UQAmb9Krv3hKziKr60pOjXLTrYXb/fJsGkw1mljjyv
q0tFSWIeiQsjd99vdlo/b/Rr9ORsJ8/JC7nLwVGJ6RhPOmjGkhZlUuPY9+k7gCRN
g+5jCdCa6/CyeAgritngqgczGxJYP1bdhLIc6oNYsc8G3VxRv+PpdBvUeM5rCBYO
DijyqBb8mzRoddzC9BeSElaL1hosJsCkAdEBwrwHPbDtnlYLulDay2BuZfCNAE8B
yOsr0s1miXr2/iZKWsHQe5avyMTHr+TURkCV2RnA3UiPfKFN5tfBltfLAviyA1+R
rJDAOhvbYeRww/r9rmMSilszLQJh5GO15wVDUa1hzNE0EjFiCEIcbqy00aTOD6SV
fwcmfjnDcdg1ZkuTdvnD5T32gybCMEWLsB2fGtgrnELnZ5YLkYcsYTkJAWrdUBT0
zvQW1bwbIBvJWKVnH2br7tBRhwpqKAWhkCrIlwfVw2hex0YKM2kTJVyTzZ39TInU
QRWnAk0QNWkiuU5FiWwkop/7gYLkMMmLDHX3RXJ4dIr/uxPMWh9Euedh2UAL/4PD
XYBqZBskIBlMjxiT0iDMbR5IIAcJ8ekKOGFzo6Pd6h/wTKmroblXuCg5BFmROawi
FNs98TVjnOaRi7Wf2SUF7mG5FPiyVSK/qF5WP8qa1yNABGiiRJ5mKUqKRJ2OR2uB
h8B5bCmQoyjjpJpgakTbdKizPKzat/jotG12mdcLGyaq73UBBLu/rmQTWa3mslKH
76g9TWhkucQz/kCivSggfZX7+E81FuK3vq4s+NY2RInIyI0ud0bpFivBlKzLFgvV
SzfUE2VHKTlXoAywBa1Rdw63cN+qksHuGLf+uUcRCldwi9rCOtLbrhbsdtQwxujS
r8kjuazJQ+tjOUhwCVFWYUesIT7VpPU0RsD0JC+XQPUrGRCwbFL/JLZfRknuD1Hq
TA0Lvk9ZpUoj2/GTWJJYnVnzkK0EUihPtC0YmVn5hkT3XegnOcWim2PA/7UWLdiO
qGtQD8HjWx5ebucdQ5gp/ji7mKJiQTNlu+2ra4+G+qW7l0l+x9ke4/D/0ij/4I5j
Otk/GNvVxpdvFujuu2pon5EQ8eXqo8oJvZ5ZcNfdBof4vjcqb5vzb0d7D8rpxPMc
4GBBC0CooRM4mMYxPacBWp+zMmbtscL4T6tOdCJNnnaV2cLqu+VXZAbMHdZMQe35
Fi5twqRGD9SNoiJPFvSX8pxY3CSKya6GZBFNGCtMspKVO7YptypG3Gv4wWqn3MKZ
s61p8dQ2TOIjXQjsDiDFeFDQB6eMHW9osvm/RqVwv1JfKbUcw6+QFgkAPOV3G3LB
S6v3EC/wa9WkgWX0KCfsARucaGGl1yiJ6huyjibrOzG3Cpzg5JS17DfBvYpWK7ty
yeSV8YkA62QjwQebUGhOGrwdrMAtPVlO6msFCEloKpWCCsm3L+jgDlX/hoJJT0OK
CLeaFFG38akTcVU21QefHcdJDHQc6ThnyV1dQsXDXEvzV2J54R+B3FqP4rKN+XWV
qE9dO9x+dCsmFXyLikVB8GtsVyoA6ciT3QtWfhmwoa5ZGEAE6CGcByU3eVGefa65
Dd+osw8/6hnZi1CvZZOU2I4LFtImJtundshcvZWOw+wCwqqf8iZigY7Cs4YWiNXV
vrQs8Gax76ZAwzrLwEoRo2Y1T5T1aLFkKCpylS4GNb6JxXmDpnBVcrFXGCqpQtDH
sx+FVlX+jmCqgoItUrKFSxMIJUBTxCr8uE9y80YRzjVBeGfKZyJFFxzuuS9RBn25
DoLJFw6zWbapq+xPmZHHHbMKGkHXWC8mBS2XAX1wkx/H9Zvs2xOSmofCKNe4QUXp
a3feIFGVkjx1PE5q2YDvP2rBNODcm0PiQaX66RLHOHWzDiKlErJHR5D2pfMet2QV
3P+138AlNVo787EvdKXAngoVNV+N/kdzJvghTN7nhcYbJncthnNI4u/R3SBF/svK
qHB0iv71uOW7UdhmORNdQgeNxwn+DqLs/1TP/yHdQCH0AVGNIsk9xoyz5RUYxOhf
O33HW60VkSBeViMXB509RX8xL1hIlPnmAY+45HHjULqoLNj9p0SQLGM0KSe5JCqA
FFfkciVWxcZMVHx8/dOuADjTgsKS1vNZI3y64xxgU47/1uK3rATHtoJJJqhA9gjj
RmJb9BBBMoDXQ0erhARxPrBgoh9ZCkR7nDLU/Ll5EdZwj+Tngh5kgpVlivy91obI
fJomNTJfJkhSBiqgWawPh0Gq7AHt5YIs4WBZtRp0gkt1ScwuVYadBSJ5VAtY9A00
1x9WK/7xfmMfuMO0SAtsJA5kRpt1Pog5w3MMezmNy6i3GeN22uKLKVzl5U+mPYoy
wjjJnGoue6U4pWEdQHomKyfa9aCbFF9JNv5/7LqOQIrfDY9WW5tqTxe4X487hXy0
onQa3uEF/hfODFC1munHAKSxgKd8LJ9cZlZe4RKABTTwgOw0pggk/cd5OTP/m1gZ
ZET+q8tpULKwXYH33z1nQJmPl7KcWaBw/Z8Zl6MTNYqqu/yUD9i8UjzdO+uC051F
0SLc6aED8DvBD0NkK12ur2SguQlVL6i2PObgQMK/FJvWaygNie084zrZua1cwIWK
J0AV34JF3T1dO63RWbUEP8vapS4ahLwzt6nFKd+Z693Xe8ngRi/AlXjZzrysvZIl
c6mcyxctWJ27bebHpvWaxMWa22gxh5VNz/Z0ZNBJtMgAHk53uDf5VY0HmgXSdFsm
0Ff5K/Ezx3MaTth6qdjD/Pe+rqUfxtSKZQnCt1kIxRnzbfjrCSoH2z/erVWRekq5
JDvLnMLdBwWyXLZKMu24oObYJ8RkRZuHKtqISqUQvvDOFdApyv/3MHmIORfOaZLB
YHFJogPvqV6TMyG0iUDCqe9H388HZ+B3ZofhGYr2U5eF5Hk1PqPzMrsY3sfJW05v
jUmBkmvjsNO/JrUpu4V7duIaLGL6OnjUHbmeCcwUEx5HuwTkUyNKzXL4le2B87RM
gmqdtvftLq61gJ/w7rMEQzg0IoRwgbzEuZC/Y0Fzz0QsY8vix3ANGWp7TvfgDAgr
TzTsSCJoixCummi4+GH02sosoBSJxYD+yahtdWNqal6ziEv3NbqST22OSJkQLvy3
so7U+gKDbSulp7Dfv8YnzfJCdS+ph8gevCStK45kggyENK9DnXyoZM2WkHwPDlDH
OSj2AJKnxpnPi2RrknhCy7pYO9U2evtXbH8T5kL6EcxZHi2VA8Gt5TQvqiu++MlF
oR+oBV1bdK8DZhYFle7SaXttZilr3XeNUhCjcASyyaa6kRzkOQzB7XjpqtunYBiN
h4BPIAWJWKc39ZhzE4J6Jyf/Eb4ppisYtWGSI2mtCUqtqyOweJ3dwdv8zHW1cs2K
KAhmg3eo2y+8T2/8/omQW3aKAZzV4MCIFEGxa0xXYcYqK1S3y8LVw5ztVuBo4nTC
qbc8+n8mJvemjpZv2Ca3PZl8lSltOFdb1Gu3/HPJdo0f39BvZDShgQ0R/HnHt3JA
HHgMSUEeKsMWt6ERMlHdhICFnDOpGrT9CPWh/NbZFsmxkSt+YfTUMJGS7zwYp6pY
eX5wNu4309cURZpnRIfTT8hskNmaN58ID/6fZL09OWBygictWdIMjkyyvvPH2kGq
opGvbMoZfbwQI38mLX6LQhp06NulQjaKYXB1AmQpQYJVJVoxTc7OJ7ucGrQ+r2MB
vFMR3wDPsQbmqhhFGwRjpc6LuPJ21okQ8238fsiZZ7AHGzvcemY10K85M+EfcqbQ
76scCfCHpibrrC5bpJ4LUDGOa9y9/tyBl6MbxDOjER52DGuKLNGAoq+ZxD7TZAxo
O9SeBEvd/pvLm4FlhIRt+8Hwc3RNHYKph/ubJEYknTlQMol+c5UGbtiqxmpgXkCY
eZ950951gmrqKkHWumqBwwbVqQQb0MfmLJLRYBieO5EPQak04mcLgNwBz+Ytn0kE
f2S+VT7I4j7KlAEdSgdaFBdV2+UVGgB0YTl1jdfGmJ6KeNrNBpHzxjxkU3YW0rQ9
KVLEGOu4LPQxYWyoXfO1B7aZZtk3yKc8ZhA+qB17CPVxDsIPRBjQggShEnsbXOOJ
M8XAKGTG+ZiRk/NACdnQZemM/Zg0dh9YndJA+/a8udFpALxKPIYiMkcy3Uq4IQKF
+CrUoiwSSKY2a8+XcmM4FT3QGbqlmC+fa1yjEyUOeYAbd+8bdyLoXP2YAPmYwHNI
yhAfiogfNEK17OOD6dhWEvyZcIsiLjzxT0srPr21Me14slYe5MZP/mrSMymG2iPC
bZvmq4BJqmkoQp/Wmi8OBZZn7fbtazsb6+jCy+T7u+6H4XcpxsGWulWnzTjsj4Td
kS810SlSOBRJytow44ZdFwRVxzbhWBYIncIj2l8VI7KDpT6u6RtOWdlX8dcVqbDq
HvVH2iLM9hr3i7eacxgGcHNmnW0FyKe6trB5hsCdrGQKgeQmGKps2zzg1OpC06rw
EZACOxtoYB8nyMQiQU+nYM3HCG/w6NOcoNrUbeMR/Ycv/irv+7idTn1iK/LErsPE
KHZYjrCdFUOnDB2GcvNGnQknXaNLSorD/WvpCIG4x39UUhUHp+/Tjmt6BElkB6vi
CnZJyU6MDF/ZnlnKHnmehpAdvxtCNeFuOy/yFLjS9cTgZ6lYYt/wIOl0aUjMf5MW
IgpyaATRBGOhyy4mcfINeq8hl7eTubRQu/95BA/n5jmbw/2Y5Ql2ueQ8DFvRug6s
AwsoJfeuQE2dtQDFknOVqWuDQAB/3GqXiTh0Vun7Y+WuhE81ozTsuuxTzNfhre+v
YL5Ap3LfP7HOu5mY1Kg04eHT288iDjFBb+28ofdL9UYVVTDayHN5ckZoMG0JubfT
A41e56AWjzVSBW1ICiWX3U7UNYRD9OLoNPLwmRha/gDXNk7G4+u+/447b5ObUlY0
kjpzCf7f/8axd/HoObzhFtWP8oKf9zPZBQtMsu6lP1l9fwTKbAHbpfROt3mVWTdy
MbqdWIZgm9zv4OchhWHa+rMDEjX1bqpDzbadogO1aAW8xc95p6ggHK1Rs1AADhPl
NcWPe8S62RfHXHcHWQDQBbAeQWe1p/otgT6o619FWQnmwBASO2DC6DhYwGKTHW8o
2COdsE0qmjPflnEMF50m/s7gKULJTtzb8cHEI3/1G6nBKIbCe+bcuKzWKH0s3ecl
5uwK19I2umgPGMlBDeChNFkZnNOlilQOn1Vrf1VqEzWpqCuWw5IUMDeKnkMhA+/V
BgEVMHkdqLtfoW2UPsVfrob9weGCefnDZt+irg8+S1kKkeoYjnpE58lfKSXC50gX
qAwasRcqOph78038oAfaGIzt3LAYLCSX7J09+2qFj6mnPOBxYNy0Jl8bg3YFYzGd
4UaBrp9wv7ySI6sNLZqJErzzAg009/tNtIrtodEP0a6bkptVFNoJV1wduI+pEGrL
DczE6EEOtohlFPbA8oNgfrRc0EhPS90wvni4nm905ujy3S+xxxXo/95bAcnxPuiq
4f3E+dj0dMN9ddtqntvVFXhJ5MJY6OIZGruYpy6/898Z0kr4fgp1g15csEX7wxF8
07KBT5RzNawYdUhmIme1vu82mifQNG890n891Ji955tz1CNerz0h71mvN5SP52Gx
lLWRvEJGoC3InRttCDDuFLOQauSpvgBUzwcEjXQx1o4AsejxXPAEk00a59CqbF7x
wL7wE1I3D3fdwTvyEalB/MgBx2t8h1Aww8Yo3OjQbe9XStCgPlv/mgZqrOtMtfXf
vLo3xUpSCYdnBpjNYRZk8Ci9W6eTNiShIQgTTnCoidJGHDi02cRY0Pl/co8JU3fj
+J5C31Mw5FgivNsovSFIh6B3yh4uA3oBMttxDs+tIMGjdvgl75XBhsq6X1aTPsgt
ynBQ//C5JaRe3/nFkT4XIt3IreCtFROkzFsxBGdJ96D6B8htrEA0UvI66h0r2+EE
Qka5eenFissjuGajEjMJPJNF/1CHCca54QVyDd6R0rQlhMvD30Xd6eS8K/R+gM1/
BX8RXrn+e1NInaUPw9eSbiiLtowsWN+CoW2yEkwheLyaTIiAB6+UQQG38FvY6qO2
BVgLM4teLkhD5DjDEmoNaf+L7VlisXp+17eIVNSOlbXvk0pn0gQT8pfn4cOxKX30
LdDxFKckyudVvqD6wAPr47llJRIe6jC+YBGEPDfM1fworEBS+T2s18oLJ1J7u07H
jJFPo85Wir5+kSSilr5FV3OlH3iF03y2Cf/pvHxD/BBk7pDfbQN+SoMPBA5EbnZA
BKhDPjs6ZVh55IfrMFgvvMP8OA4B0x755iRpQ3qRGsgzyWymFsgmH6NdlP22lf2I
S7MJOBFAuA5EqHiMx6nUkhEesg2ZX1wvIDyqXjVGY6ROiZvasVnaVHi7enGjfQyl
UiG99HbdqBuEx4n6beQAmxPGRFlhp39X55dEwmrSSjlK0EdgasRfqHUvzs8PyQE/
+chXsIKHxTzcToGMtWBKHWrcRqGkz4f/w7Q+Q6PspoP3Ahy/aKCj9HcxmcsL/Atv
MhZYDi95KOUk8FoyFGSLzK5XTXnY3nb5y5cdtDz0FhojQhDKet2HTgioHxf1wi/1
Qw79I0dFgRm+HJcH7SOxSQ4KYGOz3K1pRcWr2LlTHaoMvQfmxB+iyDSjwaRdTxQh
TR+4ZmgaLkz/d8iH6JXQMjkGqTXOAxcqI1VVvA9xG9rNm5P+A8uXd7ZOruDQg9++
Kb7wjFIBMAFuGx4ADOQwk5MURx7vPcjMzeEggZWemcga7hMLbWc9oNHtAkuKRJ2t
+IsRfByjqt5EvX6n2ui0VtHzdTW0oe584EEewggnKHZO2h8RUN/yCcla6JwJQuL7
WubwjpmUTdEUJqt0YdBWDFPfd89cRpIbBE7wHTql7cI0OxjfNLDgKAaPLNaJXN89
LvFd6RrunYZB1XDyGTFl5yBtLKjxDzzkJkGD7C1tAUT/K0+7uxf50wrZ/FI2CalZ
bYo1a4sOn5a5c3ZlDYx47F4jO7Xm7fFWJh4MCrnJTEpnLy5yeM/AP/uCxalajdBo
t4O5LzoM/nO8SE0rQkmsakuCDaB2poOzgGJhrpKUeV+abEB3sq7kknFqzqdV0xYx
Xw5pmBDlOn/K+een1EQCUqdgyyM4hHf/SxLQveC9L6Y/fEFQeO3X6ipLSJGZwqId
irqn4bvYcbz/QpkzmygyjX2Q5L3lA2LV2BvVBQOSw9UCV0f9o0fqXgQSxtH8b0vL
cIt9Clx9tz1m/tKmHSiGnsi0CRtrvjwJm9vli2CWp10E34WlolGPg4GqPXiW759H
FRGp9b8SBV8xFlS94YtBefhmQkupOwP1B5fLZQZhv+ect8pBYTh4sZ9exqPsaM8a
bQWT0LqzRxyR6VghcSIZzbsVovnYes7UshB4UcmfmGDksbQorijm9Sw0jZ/RYYOw
CN3hEgZgCB8FnCPAuVj71qDzezs/4dX90Oogej/i3OueLNZCF/0FWTjLi+y/hogc
vKLVq9mE6YFVIZWuP6aoEHQZHdsE1hKoUkg37gxbkCCb7obAa2Zmur5ki7nWAcHq
zANCi8hw+Xb7tAiGbottQB6G3GBf5qkpBOoY38SvkWHpnXX+r7M/F1THChHKfkiv
5VOhsn3TAXR6RdJ4HQkTPUOxiK6xNPSAqleptGGqA4YVDG2SRpwu8syuKnKV+jmY
erZBxNwxDbdXJZox7mPnOdV5C32zTTVIHBfkEmOKQvsJoxP6GwjQ1z2a8gg6GFvD
s6aV1OHOm286bcVfYnEbtlww4z+wzbRY9um8qGr00JgBKphVbaDbHmqlG8iAzk44
PsTrsFwQKS9G2qcbZgOUdrP6TEFTuEo0imGjaW9OINKdzb0uhb9hxj45nlQ++FiF
5XJEcizMoidAfoSByRRp2RWNfBt03eDGZGNJrZDj+XXnzds2nlyKsSs8XCfadwuJ
FPndU28o5nqHoaSyNcDmkpgFvlalVu2mPJ+JKo1NmxeIvB0HsQabs86YWcaT47hO
VmGsuBX1dmUoZ7JOURmF1ZINkJYUkbeC0xNEwweqs1r3sSl3j62tlvnRHkAB8Q6D
EG4vOEAo30Ug9NZnOVbQ8tvan/Jn77AvdpnViGSHd6mZraujLcj0OgYcOXb6XLCY
j3O53o75aZPdh3g5Gst3nXIwU3JICGHHs3wAkO3Pqal5hmoV3u9FC7qZO5q6r3eY
0WyDpnqHRSJracma+6oGlnzNDlAlUhqkw7eppdoWMRp81c1gjD0BLM2/r2jNfJdg
Jci6cJIrb+nZlvinAwsWn1hxnYO3v4e6qWH01UEna84n8FMZE5yON+1mkRRZRUwV
yKk0h6/eB+0IDC4IMIkIziCu9V+WU4t5LX5YM8WmR2qAZduC1GbSlCRBW7utwbAS
0JzHWXukE9ILSuu6veZboqWM3PzWeb3Mqzh5bcZl9bCIrj6Hw4VQuU080EKhxCIt
zBUdqn5V0jD+lNsEGraq77FqYI5uk04RfV34ToC8cZ1R1weyZ/akbrnAFCWckH4z
/Bbr9FYgAFRomUiswKpo9bD9RZ8Kr5UE6z0gXf9bgkqkp9LUQq/XpavJuoXWfdle
Uz8mxIMSPyF5zmKMNtVdhfAgJTXPqW/w1NzR6qJNDghcYpfeBg/2rCjuHNwWBJ8L
5TsTv/WGKktktlPBqpTLbySVnQ0TT+rbjsZULOyogab2kv2tDVoqY3Es3HIO724s
tQcU38BXhMb+/CG8xWD/eEAxPmWYmbjfGE+AbokCpgRSqkjxC+nqh+cWvMUeJMBe
OXPAi1iBRtj+kQZJaJ6FoeXj9VsIqlfnhj0+7UbHf2NehsKr/Rk2VPe98nJRs2j9
4Io7JOvJ+B1GGrWWr13y+/zG0QNk/nwIt9TZXXQCdn+vf7OhD3OKT47cb14miDIP
nqA+yyhOzEojigTeg9L4aUXkMbQBxffly0X5rdTOySlLd5qcd25B5DC0bbvFq1eY
tf9EWPjdMxzAk/i4NNIpL0X9bKapaJOReKifHy3riXI+PKPy1NZCAelNj6nuCODs
OIUzE9OioasGlA4TsWsCrv4tEjy7t+xQLZ+svBstRUziYxoPLDkfEce7noYQaCOU
EDvgJMRbUg3/e0KX2c3TQA1bD1Scmt8uWAj3eJWDrNaBJlsV/ZR7yQCTd8lVKh9S
B2Me8vA10SSKQeYQ/UXx5A7/En/E5xA6GyGmFDLUGCqlDWu7LDuxKdbr+fhqC5ne
SnqK5XKRET735aaBEPaf+U5Z50WFq9YlWZvjKOnHlYUlrUz1oGAauO3HVYxgMT5Y
Ag4npyuzUm3HV+02s9l2deYeA/ySFTUMBZ0WKh0MYbdp8pnrNSO6SequMkvk6O7A
N5Rq382MGwckJ0Rw0QkZOvFay0Q+Bu4g4NqNK8pP0kuiReBsprTKQBl7IrnHRTsc
LfI7SXCsCgLydFDknMWyjc59RhwG8xRvEXXcwzfnQns2gL0xtHOkHjgZ7lQDWuyP
05rJdZWpX9fIr4VDoaOwSl/qcgpLv4aQJuxhAC0qyRnSrmfXD40V+af+LTDVK3Ar
L+6Xgk7cYN0GcfJe1leX2VoLVX7hvlVDRcx6PHebKxlZYHfmOfRc8/Mv/wLsBiDh
bSC/UhUR8OlO51BgTSr5kKl1aCZ+CM635v2ZKjuhAh3xNgBAqG+TiEzY6CvHAlko
8qhixRXWEVjKEBfwbEvK0zlyvnV3BY18Xi11y/RBjXUszQwgA4RMXXZU1mwVE0hh
NIzHN5ajtKgSV34IPehlff4iJJd4CrB5Fj9FiCju2niGPxkd13CAvfNzgJzuu+7G
JMxw5Rou7Knal30Ly6wg/agCqa0OEysOBVagu5W6xiFRIH1yxkl9mfRWRjnqNqXI
99GP0HmoplLJaHhqPRiAj+9J6ea492hnWnLjgfprEeJQ0kzJJ1EABpcEkn/ugb3g
Xa4Rqu1nSwQTnRIUh3qaktVsVulo5Nhhkyw/o/qBRgEadotFy5cmn2wUF0WbPi2y
Cvx9WXbM3g1KqS6qam2cyXschDXR5f47spWro1Ys9alFl5Yl8c8ZFcTjccoalfje
GiKB7msIaLqrJIv8XznYD6QGxDIEtw0tXDZ58Vt6T8aH3DdIMyJs+WQBUTYzDsjA
Rrthdn+GDmHyvIWwf+daokikEjboVXxCcOl1+ndnJ9qhH9rnDc1EpHilB3KLyxm+
oD5aML/Qz3Si/o4iwyaYVANR0F/XT4T6ud3rzDNlA64sOAjwOEOiElpEYcOVAxtc
YWOSP7HY0nlkyjvWf53X3E3jmqjoDXhQJe7M3nWmB3xJGxcL+Qzqqv79pDK4zBak
d3XmWHyhF77Bfow9VcOzV/hIkPW5GDZ3u8jTzjHxQJE9dsDPMKyb/c3g+uAuUYKi
sLlA2I5XqfwouqFDefx5+x+Hd2W75g3TKGj3J0GfkIw8IePLNbatKvakeXYlJAGD
cNwRRZbxMpC7XsqKggmB1gdAvHp/VYVnbtjE1XZaQ5whyj8iwnbdoJw5kwZ3WB6d
FnvgVN0m9TFsl9nYdssvJtmNOWW245Gc3DgzCJN61o2brQX+WzAChvPpKhrqgVyZ
FBgX/aX+piJyMmTVbplc1itFFRxQEY8W5tEu/Jcfjwk2vTb82d3MZU8JlaFjORbv
+aQUI2+PKGuF3ZRgiXeOhluX3yvtrWYFAIlZ6XgKwPYMoQSTTSaVxbOSR7WTfn6h
r12zBVYcBkNLLnIfYCUcIpFV0g89tPoNPRY97sRTA7RklOWFpFOnJz1zD90ZOgJz
OUcrMBBL34y/ki2B8x3cbzOfK4cIruX0ec3RvDlcJ9y7jfe/0JPIAjD86c5tg7e1
ArkPv4T32D8yuUTNNCV+fwN5FsN9MT0Efp/pKBCf+MUD3jNg2kjlEMp5rb4ww+gg
Ew+nT1rA7bF4cBkNPMwDk+CL0TV0GJTuib6gywWQLK11tySFfLle7D3+JFlBLeIM
mnTtWSMwwy5h9njGUU+XkhJwepa2EKzDGlX1MdBMngiK1CfDX6r/sHImaEyHZO3f
+TUf2WNZ17GGPN22392JfgE7KZvOgqsJ+1z3wK2GfPQVSTFlRFHtEa9C1x6azPlK
ge4jAHWVy0EWuaPsdThKhqy/CDxrQhjtQyREnpO6Vsqp9/+kRbmYb3skVwXSbrO0
+joA2TG9U07CfXTmm6KpbVRUR6kEdBTH0oOZ7OewOP7dC8PnQ/4IWeGg9/y2xcWe
VeiqnvwBFVvzD/odx6CmTmEAqKzeRPrLJEQYxKXU2wWHp2k96eKfLmn7eNLJSC1K
wHzZORltJ014oN9I1OF3fj0yE3Q5GEKqlPYIZDEsSYBvU1YokhOl2EcV1NcMldN1
PWS3Qyqi6dS9vINEDLlz7dkfMukSe7GSAowMzFAmiamHJlp12gNLeFo9gxqrrywQ
V4yGrlwFKBimDV8flOwoMPGBozt1JBFh09jtprefnAnHIn5wQVLbnZzuq4u586rr
KIfa7ptpCoVLGKoWhPFrRCR2ZxDkXY6O6bQKUkGrlxuo2ksGiW7MXz6F5Jmx4ftp
+BAJZR5xzIruKyLMlPS+5ZAmff4xpXhuN2fyJ8CedCpQ8Xa10jnNCjLhbq/9B8/O
NK0kjQ6xP+CCr+5MTaGWOyDMVRapAred9zzRVYYAd2o7Lh+N3w/LZhEDr1JiRaGn
gEBfQmk6MBI37Xd/muU/JTezyMPDuic6NQMVdpmO8nCrIMOgqlQIFg1KxAoklP6c
YIO/rN1oLFYCG27B9oWL2pYVsBL3B6fD8Z61RlYV5HFhAMpT8IXgYmaCRyvdzGnh
AbulYJsEO5mMYI9m1ej45sVrqQVAngvb2bRSzWZTB7hTnPgk6/WIvarbX/zi6Lyg
R+Z9DhXg7Q1kWOYNzSV7PMA3/2N81rWMNWQDfgabMAp+mzBzWwqXTE9OChpT/02e
s74PNIW0oAJgoUN5OYJQbHxX9QuOEFZ0t92n7ga24xIxufiRQqIgIsCNqvJpNdP4
8RCG18Esae0raa6suswnqSLSLuRsErRfuxajD6iiNbKoc7mKfq/I23EngJ3jV5Eo
cCANteEUkI/HrqwQaV9pNb3ODlbHoyLzZ/2jAXrEr75jbHtQ/hwhc8yL2xuhU7dE
8+Uoa6rYddXALhLaz+g6FuzfyRh1VKXwEk4OSjXoMT9VGKIRzFDt5M8T66Gfroin
ieXpEKp8xNb69LEa9+6RC806cSSvgrlr2Oi1msIrGpdEcOwNXJVH4UfBdZ8K4Fs5
T1XgPWID9D+bZK7ZB1GbWe212cWi8P6Wp2vDH2fypI70nZUiEEpri1WFMt87hckm
RKDNUT7FagKMGtycQZEE18FF5vNtNI6pGFta0Cp51pXPw1hDPLP2//vzIKTrCSUr
sUr/uJ23uBEnIPd73ZhFcI1HR7jfMFf14ucBTB6cq7C/Hkp6fz1O0hAadaiGiMzE
81oiAVXGlL+kCqu0JWlU8V5IFN7Rgv9Cc8v7cJ5mWfeSXsgaON3mJtUnIjlgT+ea
EMiKdlxMaQbqH0zN6IV3BfPHIw1Mp1fKaEMkz4VkxYrv2vO9NHr0VmXWw6+AfOaS
5cU2va6lpKRHDvCW8EqUBhmB1+8NEY1ljf9QDg+v71XHhaeJ7cMZfOY9kKWGhu9y
5EU+sIFJnewgS4phkCyMN7KyrSWcXtRclZ9V7myvNzju2JpJ4C0gaomp4XNPVK6W
OmVsD/3ggRs7rLy/G7fIrGlqHJw9WUhHyqf7b4dvIHkflw5njdZXNM1CVJKGdP3e
60PuMxXcbpax55ldM9qEzuyiEKiMqDFsnbV/C53mG7bfBXo00QxJua8+ilBfmTdu
eZKKUzd6vwyiNkr3JX9qrgJnbIttaXl/ZsXlTrMDTvL0PzyKusCd7gwIUdZyAcgC
REXW1aAZHKDEd2mJGnvkcSCrcwPeKoUhv8syOtxecy6cPWCrVbegINp2YB/zOv2B
XoeZsjtziqaUROHJMiX/AUZxeZEUHfGqgiwLY7Y+9xO1FwQLL2pC5pqxgM9pmrV0
Wled+grLCD9MctNEEXNq65TVGyNT5ZfTMriiwK6ENwNWl03Yklg8pYJ5KFXmB8DW
WiPNl2AfBKwqYO4Z+hxpaqKnquPPO5Ohd2LL7f9CWFWpGQU38ZiZ6nPab49kYjhy
5UZe+JlwwNoSdmk7mdIwzHl2OtxBLM7bU4n7Cv6b7HymqYzzL7EOffUvi39f94lL
JKi7NEpGN3EaGiYxzsS3JvYPHwsbRcCiSPG8x/iwgwn+qs7tF0xfOSjZHZbdPhEc
Kn8qV4XkiWTrE0hzOIPT+38yTpR44nvOeTHHoi90JzeCsvGzvQ/ED75e59TbGGSX
fOdm2Sb2UaGF/Vwv590wlIfGecBHh9Q6q28icPWvXo5aUt5vqETPjkebluRfCuLN
gX12DY1X+pIiTaDHXK43JfQxFuSmz3efz8vOgfT01U4BRk47lAYeWU7avji4jgXb
pbkFZ6Vd78NKElrxnL6JHWsqfE3ZvyqyPBXWwC+TjggTTGk1uZ7r+xxyAU0rgpWk
C2459F3MSpLx61jBEF/w1n/risF5WTI3rfV8tcRYqwN8i0oeFGs2S+F6VkycckEK
RJkvyK1Qp86Tj4QWVs+1OLTClMUv1EtB2x3WS29R+PM3LKKyK5jRY0j4gUw1mo1Q
N9InMUv5teRZ5oda3VzNd+GLzzfoqURI3g8eZxIiV84ChCAffpXVT2Dil/VGeQi+
hfKKtYghJlmbIgIYFpTdJN+KW4cZkEnIWLLZ8heb3JoY7lKakGmJXusn/hBKPmVJ
HZqWEQk65ZqSavuWmyi9tYPPVwEciuZp1KNGoGaMLTdWQOQoertX4wVdpEY9Yg04
c8MX+GnPtqYVsfwcbuluKYd8hyrm5BV0krSSBBk9qJcrWRu1nCt3JZ3RgqRn1vRZ
rp43BWO9W/LgALG8k8F9VuZ+dTISckuEXjpSKFSZoCt9lUynC4Qf09NuMnw2HFrt
DhJMuiIb7WUiiNU6l8YVzAckSKPk25CJ5W4cXmEuVU3ZTgdxw2oE4/RdR8qzCWIi
yXTdLPX7GMdHEo2UJbhkS/D+HFEBtP8eZ7V1XTwMwWrKkdOcpdc0PGGrrxlz+oQt
jLuTTinKD6fC0mhtPLEf4vSFXBMQCZnzgJyerQMO8teWOyYT/r98SmA5OiehIgce
GZLpB7BX6YiogoqJOxnkDqgt8bk+gNt+i6jy4YBczeJFHS3htYnelBwLEFlFiWHt
DZYuUEEjwnKiTFjwK45tMmyehXGPlbQ+MfpT/MPRhI8fF7Phz0394q7/cxOiDP1+
xAcso1mXY+qBxUkmvNgx5fUVWd7y3g7wVB9KAA9QA+UZdplCQeZlY6GdHdH6fyrk
gk2LZzU7I20N8NGChz3wkPvE2lF9+YfDe1UAVIoEhya5AieP50kxTAxegbW9ioLx
p/KGwM0SuyNSswtdlPvEYGFMRJ/ouHe4fMD3It/aTdVnXjXovbTKNoN8NH6N9lOM
8gsxzawieQFgq/waZ8fKdHDztX1n276trXIsyHYBwUvPdI2SMXvXI/G/V0d8l98K
P8ExazASFKZS32O2cEU9R9ZVBcqO/wElNKNX/2MjeP5r9mOHN4fXriN6AAlMiptM
u5mmQS04exI1l8ig17KyMD/JzjMk3jO4/osFfKFJDgjpzBTxUvKTE9LP4GLOwJvs
YKikpw3IIF8aOm4+JocekaIPerQzrmHFn3omjQe/qkwmr5x8Epr1vBvIua6Rp1ww
U7lVcxKc6DYcVPoC+xttomnJgS3uMZVg6gumHIKHrmX4BPyeUCHBUAZaCe5bUmWG
tWWxD+Vqjj+6YRJOyiqVweC1tIBjiQkDRNPjOjTQBV8S6JOPZbhuamS/+iX5x1rU
DvoVfS/yrz1q7KL9ZrywqT1BnQ8bpO88+p8w4+M8uGF8LgPJDvNBqL/FR0dVHqRn
NO1gyrizMyJkvIEU/ai5mPVIGAs/mj7KenSI5a9xWcbNvEPvgack5RbBes0hUP3T
6x0CqSTjGTMD6mK3R8b/In0kgLgF9McGYyRRhm581JiF/5OgT+A10M4VScJCajMX
o9Q/pwokPqCczGbISpN4QCiYXsVLwpjn+IqTzbKZCXyqM7JK8m4bsPaTYns25Rte
P/XgImLPMd6kZnmaISvyEnOtQ5wZwx5xoS8bLFwcT1zqnqWUKnYYPXmJKqGuwFWh
c8QTCa/U0bbA+x1C1VSsXUa4xQ7IzRVnCb1KakJdojgk8fcoZsQni7SebX+CCpNX
pmSpfHGZIz/EJmKW/ET0V1MkgCKfkbYh3hBAL+flMaljvXjnCM3r36AgswKMrJRO
od6n+ztX1EemEZ+PFB7GqswZEHanfGKJbBiNW5bU96nqNmw1DPUfJLYa9L99XDvT
AUVTDBg2mnfvlnAhMtBqLY3X90SdDTVtwHGiAhsXZxshj6yh6n5jOyNMeR3YWUT3
nwHHw1nrdpllyJguS7ZZ2y5dPPJVZWkO/L7pFDcyfdBzMN7NMB6Xw1Bj3i1mggCc
ZtTUzrZ/mkJA2ZhqlaNH6Lo7dtrDAu+NC+ysLZwesUKmhg1JIfyql2vJlBU+eE3f
HgwKQFRYgKLtt0LTTC94TWvdVSEBjzAH6GgyjJfvfHGI7xH/lyEm8tCiQ83mk0LX
IIgvnmQbncKIonWLT3Eo9C1zJgMiQXru2L6wKEoAFgfYGLmDhUQrheC+7DjSCvyh
QmtYdkOpzICyY2RDy+2VLPs0o1qs9ncSJQfYudnOP688BvrI01tg3LzPZMb/sj8+
klBUC18l3meXJcaAx6DmN8N1UbTOJLGnfLw7F8yCCNvYocGqG7OSGts3OH2CW6nq
vFcEzMdt8xtY8+f6jHJ/jC/Cvd+wR8kxf9dftqhkJQ8fUcXU09XHSdqOHVjuDYMZ
VGyZ4+T59d+IvLgRIYZEJLn1GLEa9qHbbF/CnhT/qx3Ra1csM1/JYYtW14nf8paq
YLKtaRBCy+W+DRClNLlcDEZDBZEB8IZuDadQLn8YAjo/ceHYoZiT/STQuDI6JTGs
o9kdyl0rYKxgep41yie8izpJBEj5R+vhurHTps0qCSF6HCOvReMSJElAf8vEUD0C
W6d6ZleofGECvwCAzrhDtdI4Lq/5RSZMSaZDHZaStlw0QOcVNIqYfV0nF3g3HO8d
KrX6J0+ZCqcAlv0i27ZFXNc1xp7qNzjwyvZLPYW5WA4Rhw2wK/Ejoiic50dWNaTB
8MCLWtk/MGxKTKzOvRmE79Uz1kkIRaJ1rAAtGF10p36Sgdy8G4IauRJappJvnV8Q
xYKERnwCQLy7DxctMx3wY6RrzCj/0YV9EeYPp5l2lL5de8ERsQl2FpF7xJqf2Ny9
zsmfzyNkxsS+rDUc7MPC9Cs6WzWPJIxXkH8zu8u4laSE5EBku3VuiNk+kkpbTtID
qM9v7xW9+xdW6JTBHYfotE1L2TSVpenhren+RJcy8li1YgE7yTeyK6uXcQtbBvNI
IjACjpDy6AmkuQPoZ5pI6cWEdoOgpE3dVptLtEzXBRXPwO22B3iqpJbaTAhW4Rh3
A2TsfpXgGIor/+h13J1RfPeOp2tBEqD2iad+zXcXsjSkmCJs+gh+VsoFVMSNV+NA
OjSn878VX7KqgUyBZvvM8CwmC6DoS6Viu1en81ZxeAm5olADJynE5OlBORfmA0S3
huFeO1hfdTw6Zt041CLlrmTFKfBpRvatycOmBekQGveCb/s2+VVBvhqIQX7DGJ7Y
P0tl4Z9p5C/rGhNa5O+l+mLo8dIYoeq0UIRBz9CQ/LthM6VTXioggbXi0+Uh7nre
uUyLXFRHS5Ck/Ds+dF8TXFK4vnF6Zh1pwxx4+tvT8oSSPwARpeicjVTiyfp39evi
wCGk4SGEwH7Di42Ogeo30qoFBHPlmLvLs1hE7JdgvcF8SG0xua9SnjqDnDqgulyZ
SkhLDZvsXUTnLcSE2l5ixiQl+yd0tlI3U3hsZYHZ9nxZqikirhAHijKr389Fy9q/
7XcD+ZhrChCZaHhMT3nmS9b/ZkGoBh4eU0l/4xTv9O1VPNO5pnm6j51DFcd8NWJD
7YgnwVI6s5jPyckn7cVo0ne2/o1mIN915vySrI1cCfx+sFOSQEt/sJTjZo969Njs
PXQV60vgzt4ga8QVqvanFPyBG8cKyKB1uV8r2YkdqFMgltwSEA9fUUO97Nwx2MJT
AtANCw481uGpYipO0HzhHZcC1dYZLDB2TBvHxGCLpzofkctUaBdPV1h2CnpPqrFl
N7uy0+OEc6Xqbt+bADNOnHPboa+WgFhTKa7dI5kf1ek6iMhU6QlsdRyL9dq6odUZ
Sckvf9nnigolBd9jKIzePVGLox4b55VpU/QxvFAGoodE8npBr7sHAQL7PBSTV5WQ
KUfzMH1i/E30Ik+cetk8g2OFMJ1YgvWJdKFEssYNhZ31koE81KqrnfURRsnzL4PI
VAI1dPe9m9+3BSw9/1/iXiQ2YInWSH/yE7rca59LbsTizMTo+bs7p+z7VY78ceQZ
PHU9W03bOId0lgFIDJZA5ZGAcKkAdzcItfCwVbMPnNdf3jSFyK6kW55xAyYa1iaJ
H4xTkL/aT+50koKOlFxkGbnfwsAl41JsQT6tAboHFgSPbl4g7qKKAxaCx8bnSFZJ
jl56bAFO47pVdzKqmrslzeJZlERUeOZ/qQQ02fOQbQDafvqFtNZ+ITqQJEXtKsZD
t4O3sxOADmiFzuj8fX2n4IVutj9glRt8LKxtPSBt8/9rvniYpW6jqAvsJ1DFQCvv
FGHlYE8MLhPX+1IokXkh5buzxZPqNfy1tCQ48sI9ufFpLkdnuF5KP81tSPHkAYGM
M+eJ5htbCBqoFCt2OlIhtZaymcpKS3T/zbq6NZh0XUnnroWBT+N2154AbCNr79f4
iNQ12Yf4hx7xTP2mvjH+Jz2SrCnc8SkLb4PJytOX+zmX27uG2RI5/yuU9DTFQ3bD
qLAH+CzEa5lgIBEsPBU78W6IdKiNFyTnHFanPSekdXzSmdIxtM8AIQ802tzSU1wJ
9b7YKclpiYUWq2FPJPorLrqNE+L6heEx4eqr/tbTrRvQ2e+Vo++SI6XyVa1JPY4Z
gUuQSVOtWoxsCKjkn16BQszs/NFKq03qhhqTR5H2OCRQSYxZXv7xOKMj+avT2lZp
b5U+pOJxnjLV2y7rGX/UjC6rHJ6SeR6D4FtZScIxN7zbfWzcdhSY0TwJE5k+nY18
amRFPSwtT/V542QbeieOGve3AqDC1NnQlcfGszWxspLHVOVY5kV5L9/LBa/x0N7N
02SlDdBDGCOziMywuT09vmQgFlhKZYtgKjULqDguxbSPauzPPjPeM6Z+DU6fPBSU
jfNeYnSo4pcE4PVPG1WyHqT0WCIXaDF86k7VVcvDiAXtcJzwIoFOKllxblvdK6ZS
Wnr4+ck/GXSdcl6CmtYu4k7GlTl8AVsg0DtRwZV/zjOoqngqsK8CBN1C+7W6bsjR
nNb1TNt1FOUYYiYmtv9F8LplbjpAKdmEGduUcfajw/ivTk3KFb94ChiFW5nyqxmT
VHGPptboUNLyXrG60o6CWxYxHuF8dGmRPojQJzvDGZLp8hJUTVlLsESXfZ2l5VO/
06D5RuzTOqriVTOfwMdZs2jBswcyKdfNi/I8ypYmDehUL0Hrz0sTDIx6Ys+qqeeg
Qbmk9I0msZY1mSK2I/cX8pVktp5CyclprU8YsiNNyQwguZcBI+5jkTgQ8pFvIabV
aTSwoqpT9erMLezw4KvO45UQ9OP7YL/7q57NCeYMC2EsT1kTefVO9MnkA0oFQ/MW
+ddBQ7x8inFE626SdXsMug2vix2aj8DOXcoJtktfZX5zAE+EllMqHeT+Ouc1sawW
G1b7ecwQC3KHEgH6zs3DUHJQ/idUFlH40qCmctcqoSliyFufyQXikdbQaypagzLw
Dy3WAj6pLR5cqb79D0mckyJHIn6sEOsx9VlEbHgMmLqz99H7VF03QhIDurc3x13t
ssCBENcdsTj2A78kgmh04UKYk3c3i/NRRjkVBoaJKs0nF5NxQIPXkbWmndy0miQ5
XkJ0YADX3MzPXmiFFUDY5zYemPUncQoiDRHDNLGfL9PrnbOmUtg+2sj99lyVlkjO
rS/+nfK9PDJJ6LgGtu+sYtrf1iagOp2UbuWbQWuIll+OeNcsjKMpFjJ6QjZuEEm1
521WN/rg3VevaUOMCOCN5jxY9o04Mr/bth5GHFhPdOLP1oeddKGouIaouTg9Dd+w
lbEaqIVTmpROXep8OZBdAkp33IrFTWLcxBctmYFhyDq/3HXyNbyDJTQQJlLdd+6f
nZE8scq8gP2A26o6rvmeeg+poWPiqLPRHYz64g1B6+QDgHkVZNgXrKgNoZG0hqaT
BWL4mB/0PD9U1tPOopXiZpHiGzklz7yhhAjoFPUr5iTAyeYfYiKa6cTUGFWxKZRr
QjL/pvXo1MQMrfw1HOZI3mji6D9KZ+szXPJGUhjb1QCk7FGPu4t1ztKkyjOMUfKr
V0OB/Vix7CeBue8ppCMKjR2Wiry+3nqA/WsOeAnZquV6MDKn4QiaRG9G7qmVcFT0
Y4VPXM2p7ywpOS5AyDN9NywcAEVrSSwc84NfeBD6HQW7GmA5Hj84TYH6pgUeZe6G
tpR5l/kPVuEWTVTQW3+xS+f5JPo7Xf/h2omlNODGNLM2vX2eGFwkj0s3aXTepW1d
f51BTf2l0EEBNEqX7guzEZOoury17bl1fhZby5rx+e5+bgNFQH1vtNs1qKXEiYjg
aIBYBJ2QTP5qtoNRX+l/zR5ahXKPikDHY8CZjPwSeeadLlZfhAjg6uqtj3fjCzWc
obpDacQHD0lbd/YA6ffdeImLORk1zaQWKIdjHZdwMFCdsmL0TQsFAMiS7dbBrMCC
2gQQMwUIw/MOr3Q7UTxeyj7POxFdWNmBzjx6CBZbWIVqlAyRq3Tl8qpWzigNGyLz
4lvgdnRQ8saG1kn7nXAKk5WdrpUjWcPBC6I2X12euajFlfU+dYCmA9l4kRe27Jo0
spfEl9Julw74hsv+MN0VwtkDCbJAZSazvTBp6Uwo2g4m4Yxc2Etcvpr4GVrcybaI
KRTUY/tLsSJHlYJPCv8B+0hobn4lNjEfrceMB+bpXeOb3e8p8uMJqnAdEUGoGf93
XcpKpIr/JvR0vwCflDc9B+R6dcC3uVAkB2IUlypi4irP1mT/K93gJZlJYQxVbXhI
uKYEnUz5Rcqtqvzd9d4kpA0Bym9u1IeA954unjGOI8nonmB9LXRxhUY9GfsYb65k
3hIfEA3uSLW54f827uX22wLOiNqZDLHRYqOup+Psh+gXY+DqW3vb2wRezNO9f6kN
3Amm9XEhW7QZMVAR7NHHh6xSy6nf6Y/+BVsKPQln+kyhZQ8vvk4XLuKqFWA8CJHx
2mPHUFp654w8Ztve8y1HV75hfNFQW6lJmkXj03eQnZwCwkLMufpdFFyyI4nuAzAf
qXLdqdYmWcvnMePp7J3k/iqCmUX23icrU1ycyLINzopKXYTj2xDrLIjPnL1TjRAo
Jrt62fLOP/KX3FfWcfH8qEsV0Db/NW7PVl9s5Mv0/HY1s7akQ+7CnGYlWfFk5P5X
Vof0wufnwO0J6+70fGGCknv3XlMtCmVgPeWcSVgdGtMDUer0cTQ5vOrkEqL/X0Mp
3AOcILLpFC33eyaPkPG/b1hOiy0UL49xjNa7/VL5qIT0S2rX8QuQc4tF9YPhuDHE
1hQL1ljZqXc0FnimQwgKAzwb0mobCtUb2sjT5e0i6mn4mmvOrUIgy5PH0K55lfTM
hdWSbDPr6xg6eqTr68ypYvclGBV90LQ4uFAuE1aA6QgZowDzVu+KhPsG9JvwTYoV
LoQUigQSx2OHx+BDcA1DEPhvWPAxdVeXCLxaXiZC5iIr9hNg+YQYFuFAoCCYy8sI
kWF9rxaxlplZwd6faPGuwXSAw0QolIevucaCu9UARK13APrtKZqDb6JCbMz7c3F8
AIwOtih9tKL/h311gy5RjPodbTf44xM7Vdt1aPeCdFP0jcUgNPLanz7kqe4V6YJQ
vxI+4Jyt3GGc1pedyBS8I6ylfd75fcLVdEPPKEsqHlc7zclDmCkg+qDElrUcuoX2
Y/K2Y6/BRuInWc3gw1YInfVvdeR7PIku2nnn0Hc2woDH4xiB+52v4PFk/jzE0VdQ
w+sCI3Gqu6v8iIzqCv8XxpOBPZ0RgzMUJl0obAt1BPjpQDOLuUI7Zyr8P3uFTT2S
f6Ab7BbLyK5h7gh0SxpO0XCV0Fmxf6jMdHVFvm7MDzZyHeEGFdD3/GRZfgv8Ivjh
hZCOmlUzA2R8yx0XohkHtxo4Re4Syz0FqzDjjOdd8E5HTfleKtP+FQq8Mds/BFrK
fktsxCjZwv6LKrzueqm7Q+e5472Bv6kOc5wFYhHRCDB6TwOoQBS4EGhmzl4UYud4
qEFqaMQS0tXAUMdxomHStgtkvVFWmiSDNaeknqz/MA4hY0g65AnDo3MKSb8FxtFB
mnPd8kG4/+vE5rGw3ObCnOTgh/6g6uckwTfSaH6LrpuxwHzA+HU43arr4WkIGkzm
O93G+DtEvu/WtjgDIyN7QMcyTEDmRYNNlf4MtmtBWpXuDwzECpq8TELK8HhYc0ke
0gTAjWYEUWQ2AFFNIUDeHoisUzwEvZkXIVNoA02DOoPmv3fd6uVfxiPaskXstXSb
jRMlpiCL+xDrJbtlmtYlBKJ3/8q2V2QoTBnCTWM3P0Lf21wK9Pvq7QIge526fmti
APatR/ueff5FOdLcwCSSzCZTxXbKQFiJHjnANVizUVhH9DEZwGyDoqopAdXXhcBx
El4DcJwVkgJvRx+vZ4dzkCw+L6gJDll6lIAn99ETC9XZm2vIxM7dCW6IHPPDFm5b
Z/rN2BJiq3LnqZAfMz9DparqhbVWikcy5cXt0uucQKzvFK+6iuevZ/Yz25LnFX+E
8q7Mc42mhsQopSrbwOzkSIyZiQ+YQg9cHTlAGzIyyYGrqXDlvrxprXzpTZ/KlpZY
pRi/1o65LhNFQ5ESeiIzTX051qA8v65zr+sYGXT0KRcJ1UPMthOjJXagJp6Lf/8B
oNLg6g9W/65Zne4Ztdnb1eJvCjhQCQEIL+dQL822J6tIeZQ8KDPdGnjM/m1dkgEK
W2Se61bL5vdohKeJwrNJfSsNE3tnwuXwZKso5vKSreEFQrYnUWlr3KZ0dz3/tWsp
QKAOe6/a7nAKu36xuQZwcF3jGQu+G0TRBhLO0tdMYdWCyecvh9gdkvZyP3HRIntW
K2yATDb9NEFFknos1Aq1X8eVnNNNBT0ScjyD3YFrbAPqCDPVe/UVe2p98cCSlSvX
tbV9zD5cmdDuQR28fKSbwBlItNtv3ruSIMnO+EZ7odUxt3enet8Q/T/3WWOlyJL1
KsAPOp3yY0ZQgvfMsISY+NQkcCMp6A7zJWW+qbrHAdfkS8e9Crtk7two+p4/Mtgy
nVeQVQkhOxIHz8C6a5/u0CFylAFPRranlFiTap/m5MOwobzyqdMgQzt3XRMmDhDc
f60M+2qGH9pROAhNMIOpR//uZtDW9BzmQmdaFVd/S2h+q7acYGzZWxizsGUqSc9u
yxninaLTOtaSl1SRltYtmcsTV1rvsdI237/FV60uFJWbCpBbQAA617jEkT169Pwh
AUyL7KmeKpt914pZw1m5D9GmZVQDFty1M1MRJHc2VOrIDT1IIc+caml+1T0wTZky
w1x7dBFd0e5O5QGwTH/ZuaXORiqj3OYEEaT94r476OgR12Tb3+XBEye7afcgDyTO
dn6fMRgqt//YSvfcYg225i8JVKj3Fic7RDPE9gvURlTztDg3/YgOBW52FAVP/qT+
VrwmjqBpNoYbou1AlkSZa6abbYnJo2xGnMmATRQPCjK4glvIfLK1ZL0/QdmXV3wc
gl+Tcz32s9qID+tMLSP8suIR57wc+FipsVsUp69YH5r641Qv5XIYFRqRpfnKLKno
284FG6HQwrVYQCLx7jZEjlmBoR5jWsbEx3L4Mf5JXNKWAsnRjOy7GCWTsj6V6DUE
MII5myDNiNmBrirMXYEr6PfBqVsjIZ+1/8qDJOBTqiRLTJhCylPqcRIdKbmTpoHF
ojffHpTMga+aqoORfalLSu02/1GSgOaQw1cbI73vSGCujNFa27Xw4RoSERSmrX9O
c1nBGfmKXxcIEovbfnMlnduJAig1UF0S8vFJ6XvWHnJXJXBatgsV9KWTeUJelPxk
Qr1JLoMkZkVHyOyP23gQfjfEJKP21SFyfh5H6c7huSV8P6v53n6gLrMhzptvWbHv
QYAG2vBknChbFfXqTvvXnSMSg+uhH1ZfdDAj0ckDKEjKMWt272VKrR5HDHc4npvQ
CE2/H4WQCbfXzNGgkNcuom3h0W1hqHnjUftBXfg1+iv9kiN0dhmhFuwJ6otBxtVl
7beL9w3VoEs2IEQsw1dZOl4uoD74Wc1LS48aJ4r1dujJmjhNACGxLLZCT6jNHaHP
sCxxjWYgkkkC8UslzRGxNG38dHOGM9xj0AT9/TFSqsCH7apcTI0q1FO1yX8BxPwU
diq+0/dPEb0JmK0v3h974PzwTGREDYepPnGl2WMHKd3DgYLznJFwqtucxRfz+C/u
Hth0Lc07j9575n2adryQ2K8eJNKSMiEP1xdSPh9dbe6Ii8U3xFwB7hmOq4fUZKA9
wv2gOKoghaGtJfeZI5dtCgt/B3FjJiQWeVibeHUJhlGjukwvzAR450B68iZnDNph
odREiIn/iKvJz4PZY81U5lLQu8fLmZIsUG/YZDizFU9cJ4/i0uiY5W7xQDMosKC6
UdgQPDh+wwbBx/iLzi7lpQLtAI1z1hyyHN9AEVnc+3CBKJGi/D/JCLZze7PLP2dq
yNQL/c/A+G/3J1R8rd6TP+OO9sG92wULVnPkzIqfzGrqbV+4iwAEcDykdK2kLAEv
bCeXImoJ/5M2Ks88xHqZ8DtESBTsUVlGQqnuRFkN6VzAWFLG+T0aFpmHRwVwScKV
ydL7btSsULLFCeSjgBq6FWtrmakQLz2Ymjge2rSds2JtOig+UfIjjf64KDPHusL6
8SGEQaprfBky2bSjfzCLUJ5q+bubPYvGnSiNIgUcD+2Ub5hwUoT8aXdwUGYhbL4u
s14LIdATaYzUkYoom1dTa+OuHSsfYkk4gcyOQYl16jvb2apzOFntoAbB0PYUgpyD
D9rCJmCxiAgZvxccPZf+rMFtNJ6crngS4VLV7ff/WeDr4dHzowsIoRU5qT2pZ9cf
JwxvuKraqSiHe6PBVLGHClwxSoCbMshpK0W4FQd2WZljVaOqxMD7DYTQCpEZROEJ
gBgiy6sj28rgMSSE++R9bwiy4ya1bFzud7sdQ6b5svbDrvWyqVyxW4QpG6+G40Jo
VkkHz5BlXMsSZxbquMyPNtxjAIwpzvgOfbdt9TsVGclrUat7DYmKTAlfvjboR5zw
vZT1rss3BaJisDtxgSKcxVmE6EQADVLgwQfiuZF2AGe6B+nYdtIkz7QNCYYbxbGE
swV5lo5zRBKT6yLu34+FqAqvAqwoFn90Iafqh0acVv8LRiQXU//WsKsYKFV6Gr88
fGZm5snc6+Q1chtNY1R/13vBA62TH3UnEshTcojo2A8sBZ8XCsVlh3+g4BQxeyys
L0fsSMMlw0wdDhYCZXHucJNoq01qJCAfAWLGs3D15kFTKOwX9VzAmutlnxgdFNVn
KW/eQEKsm1PtFWNwZCx2eRW7sbs8UlS6JxSbuqx7FJf4PjcRKk9EiTfvCu3nxqiu
SiGTrSfFFF3jS0IQ3Bhdz9kes+Z5Jy+EoU6l9NcMS9JcSUlrLzEDI5Fopd7kQ5IN
8pd1isnB3TCdUzSCnWIapTjcGRx/bO3XxfzOwpRwpW2dT1Bp+cjco/aUc53zgCZt
VoPXqdUPbfgQM1bHZ7KsbMNoKnzr3rze/R9uK9hoRV6I/ldhPIe+VKUrFmyFPWfk
dRmJm4FuMiaWf9YKC/qcF5so/6WIwBoRWirwPQAmE+eJCSpPKntwR8zaszVXvhId
/yzhrRVuErFH3SQOfCq2GHdLi6ydt/XOGtDQkA0FmFdsd6hRgNRJR2B7dv62BNrv
9/vkbhNR5pTH9hBA3lxxANnGOkfbQUVWF7U+yyzm9aDFPKPhAPKsbRPmsphng2yN
KC1UTedd8z713B9l3EgFPsz19DBlDx/bdy7zyZizY+6yYYX20jDLL8ofm719jl15
oaGppFRFQwGkWzSPvmtzKf8BBtP7lqp0qMhf74vFC2ReKkv8lfqONj8j5a8evDC/
PHIKKzk5VwLKGtX4JDLNKxAgiGi7teDyLCkYt88+/1pSOlMk5614XPqDO4I4HC+/
fg88LNRYamzVkblnMiQrbK0ah11d9PHK/BKspaMCIrsh0RFPqpsAifWAEucJJO2a
rJCGOC5TLpIaVoTcn5fGfHCZA8dGHhY78bciEeJgNw6RO9tTb7qNdbyPsfogwX3g
q1pv2JByMGpXqZH2c9mgmlzT8BCUL1PgRdMDgBYRb4PFLImfoXJUFep8vZWlTEXo
XXAERnHy4VOvBff84JBiSnEZ7UH6cN37RhcUPgKETaqOaKmkLbgtaXal2Ny72p0p
VQm6Jvnmk0V2jQPwvMiynJBZ2ag+CBHpxkhI5qtB/JwZ1VCriOV1BjfWgpE9srUR
L7hAKwptbsxk1SjX1dsKxXWT8fUnMFLT9G9IA6BMJ8SsJVcZJtEQXH0KVpGV2+Ko
hJAEOXXEQIPtIDAT4hxvpmwi8V7GsPfj9+Gdt555ltq2pXAYr692R5At+x811XlC
VljdDdtHEUFGostbotqJB1P9N/d4GWeKjMUpx/ETtXEADmDP13ds3FGQVjUDu6/6
0GfpMlIl/MSK2ivl5HqZlSB8eWj8mKtm9HjBmTUG3H6phbMrpGgB9CLBu00rr8sS
N/RQLxAWw6E34LZD50wC4RT8ckjprCoWcOcPEXF5aLgLLi+OdemGdyPUeFJ5RICD
zAQvl+C03N3lBpCMxoUsveLdbMEg3InfNoPOPgBSZuXUvvxNBI9WEMuG7mXvUBBn
QPfAkeI4wJwWGIT+fdZZaAuZdqrgBbouCXkbEIx10BnAB9zv41RclrD33bUd4yzm
jpe3+e/RvkiAhBntD9QfAl34gS6eZon59qJOTj5E+zjnQyY8zhUJmKcJ48aj2NB3
hc2WNtwg8yHZMuP4SFFPJvtKBJ4WPdCxjOIYHYjaYHz7Kr6SNATlml8QDs9E3eSw
5NxiDQRbhSxan8Aot4KjdZ9Xs/2RE+S6HVrcivcJ6TWjgePg5g7K0kzyLxONX5ca
pqtPWS3lB6D8camP9RrnmMNUSA0ENvu8f24f/d+k60HGFKvqGjCip/Pnh/HhO3/K
E24mkDfT53OUlwYwKcdeWbitNqtrUZrzGB3x/ga47f96RX6fs/BPMyNrQMsiY156
MwRKJi7BodPeJNhLDHeuBzERfDXUxL6+oTfTsEKvBU0kczxYd+UB60vsLTJmGMCq
6stIVqzaSbPP/7BrhGViLRPmR6Lj1ElTyk7a+DT6UOf2Jm9d2uucKgK4pc1EpeDX
xp/VAkOBKPuN/bqan6nIqfbbY02/RdbXaubNXF0hYar+45hXDq0sphbuf9jMGcqC
mSXcwMeGHRysShE1Zzx7q9kaFhdAcbvUbeAqKiQVivTtbihEXzvxLmBT+8bbdl6O
IcwWeKn3ViWO0VjorinjkcQ7GlgWUkz3Z/FFpi5KEMjQgdH83TcX580r8HNUP23j
YTTlFSl7V+LQUjtqorvknibleFCduskeiuxwIyaPllfY8/ioB8wwJ+WsFWOeBtZQ
Lyj9wwmxVg9Ejz+uC8Fc1M27SPyeYV43Z5v7jfB+MpCnw9axQogxJbec3E9J739q
vlaxfIz6Ewf2tya7/zrwmmaaj7Rry4MJELNs1k9FZ6fPHWl/L2y9UMMxW6h1cKV9
voGbIiREJkXZygKEmwDaNcBUl2aJMk04VGWfUqt4hLRC7n1G6t0NPMJKYlcUNcAu
QyhVggi9302Jt32eqZrJFJk/yTpTZ1YqWp5iRYdq21dh0n0Pyj9VA9ctjxVj9lk7
ogjeN2Ei1kKB6dzMF3zHB2APIRUu1YtKTHF9390IY0/cqE/fYvEWDm8U+RYREZ/k
mGiNX3/8bnzPoPTb5khJ1syz5mNSS4p1uJl6BUL3AeX60l6tV4OGw0F/vpOLPntM
jNmQhPKDx8zG2bbJF52xzKfDAFdvgKdIDkoZEKq+HWP7C4tHoSoZnStWcVYtzYEE
ewFaz0NtcPdPiYLJ/5oXTzsxJmqZ9HrqBQpxrEKFh9LVRu0cUH1PnjzEZrGB/ZGB
8CwWB/ordngU6Nh9dZ1IarXD1XOpxUmZBOQgZ1YhJhQ/M4Ozi/6nlIwu5wS9j9m1
XnKwUkf1BdmBeKES/zgvblpPTC7cciEAE6O0/wn47hsuWiCnTHN+N/yPyZVZRf3+
dB/GD4hFeANK1na7btV7NPvGTK4qGVFUjVpc7rafGyysA3q4MUgGiEIHl1PwiZ15
0mKRAo4e+y2Okn0jnAEVrRJQ64SLuCWzo8jkermCPyE/i+L5/79UGJQzq2wtwfOj
6FBwlMjgpNgwQu76jUTXxXegIvhtn813fkoZMxfxYfLkkt8fDhjGOiOEqtHAnJvS
uifMjaKb17BwYdihOHSpDgmUdpOUElOwRNd4iS151R+VMlMUXapuIXziIGBeqh5w
2o8RtYdg3npBOmkHdhj7KU+5mBxDzD5YrVQhDur3OgtDSwirffjh2uW6haRzjXiv
AGAqJTKHUV9cCjUt/Q2263EqPI7UO27bQyG+dLM8GV47+V5Ak7sGNcC/JI6LXRl1
aEBLS4GUiSvJ6JTQDxS4Ok5ubJtetr5pPzhkxImbP3JbwFJoe1iXGIGoJbtgvJpZ
xn+D0eCqMbKqzm9IAuadcV3aKtwIUZeAzwbNcCtOZgLmxXPSXTUCZ2CCdUCIsfWq
pIN132O3IXIq/WTxERs9WZ2xz483+NJ00hj9GD5ts3CfaHUlrUcq8zYXTHqe7ahN
Axfx9pymn68vz2J63Ceon8dDKazvJCSJGFM/6K5JXJSf4Ncx1Iy30tjyo4tMR8sn
Mx+rnr5gcxnqUjkqnpfz/i1waJlizexItl16G2+POi8ZptKxdKX0/642lmtvj4bI
iud/TCIG9q8voxQyVoV1CXfBp6DHVcwKOapnIhfoXNwbW/ax9pRCjdc3LnKxo4Vd
vGIwo/gWdBC1GUB2mS2TDgvTC7Y/u14s1DjjwlMJ18qMur7nB7U0I7CX7/m2v7o4
YibQcCIthZHWSejEG4gZWal1TaTfBvXN58n6WsN6OGAwTJr6/1H3tatDVt2tuUbP
Q+JkRysCcNhl6tG9v9+fY4/jYHbgcTK1zyrK59HTgbFkYV+DSGmitLiFhKvq+0E3
t2vERzz9YwWt0i8Pnu8ixDS6XaHKYcf04ig/4QJ7bgDWX1Z3o++3j4CsHMW8ZvC5
zUgUfSXKfwiyKK4YUaLTAFq5uL3SJOJjzK5itRXelAQP9fzB1KXFcLUETx57PWKA
uim+8+rRNWuQDJ9CPt9tMnKGeFlAmyYs9OJ6Sj1VCeZdqef1Yvgr1T0gmVCGrtdY
fC+yN41w6K9zsFTxLBFaA4pqb4w+m3ViPjWM5/U+6D6VgOEJb3HZ9L/2zYbdi8DE
ymqhlUhm+ZYWpSBtI4dElT+ViIV/4LiNg4esPFnXDwTREi5R7icreE+GEG8tSDYo
EqATogn4+ZHprT0BqqI32KEvvjTFVT/bK1VIjUfLlBf/523pUFcodWi0rjK9lL0/
NgyKx/WmqDEr0aHa/Rp2fNABDfrOBvWrzGUYzqFqJl1IBwOony1VxyPn8dctK2gE
SmqVnzvVR7OVEiLilVRplnvLwLEiXSW2iqINcV1e4CZnI1oH72obIqruXDJyjRN4
1r14Yq/UpUPP+//pByBDTuH5E8wj51z/MERaNtgvDbLgHbEV8ZJycPdccB0I/ZV0
r8rTd9RzMMdwTJbf8JZ9fBIRclgZw0T0IzOwns/3febCZwWVJPOCDfgwO+fF8cDG
bvqg8uIk2Mj88SF6pPENr6Wov/n6tRuOXYlaiDMMGO5gR2Oo9aZh53kCkZGYsEZv
Xilvkmipupr4etvx2auM8rCCRmOYOMHeluu8C3CPynPklnpcGvcnbr5exeLOaZ10
55zzT9TaQpG9lLHqt6WX9flBqQgW6aNs7G6aENCIUY5XfnFJ0mgeEtRdVH+eMxCv
0u78tZygH4HmG1AR3awwgBWC7CU38eNInFftRb0aYIjrHXNXWdyHoSqIypRdN+NK
8vtZL424p6iH0C3mx12gXreJ/S21qfT1yFRz57EiA3jdNpb9bYqDHhxKdkFTBlIu
khOu5oq6UIBYUTtUaMx8FoC6C4XmvKUcP4OFw2dB0sOlfloAXIuml3ygs4itXAly
/5KVQXIgXav8bc0ZfXqVdhsaubk8gjNE2j3JyukSn7rAA8MYZsUAupF2j+Me0/nR
4nTOVUyaOczAJxUPoepsjTc2/yQt+XvCSafMEkBEL3HHBi4P/J/jk1uXOWKoyvfV
YliYO2fHG6X+qXdkhE733WuBpqoY2UGRMq6qFb/jcCWTTE6o70NCpb4mFEvdjOOZ
z8j19rt53WoGw7SbOCGDpJtEFBvnupIiUg1fu1QA7YcIfqatr++Onm/tnuyGxLlJ
gSir3xynTEf53xFKra2ilaelelj9hOF11In08Mrc6kmkoqfuxzSXhu9pQjyrBGky
3gMswYruHtRLFxM9qzrIzhwX2j7MDH2/82T6D1cqJ0As1ALdu/aC8LIM7D9yhGOr
5l2dcNFZmljzqCN+GyyQ18R/I8Zbs9peqZjgYnv7D22kChFzbTlbxTFy1h8VJ/aH
oKsbO6GzSEvs0N5S0fhgL8ezywah/cnWtKuP7RS1QYcJmmsmWA8w0tedpy8oEKbr
0/EVdTz2a8XKXNVYP5ROXaxQKjXY0+hIZenk91Q1/ToH4V/WhVZfBcMQOOM4oreQ
J1UBokQJeBHm8+XCFtrFxV5yyhxqAZwUVhPE6fplO1yyHxJbygP3ZPQoIb0BlRd3
TjZ6qilikdXrlMp95bo4hE6ln/fumDboTiyYZMy4LXczT/bvK8WBR2qq7NwUcNqV
GRY1ZEADTXs4iygjK3s61XHXan1wBuwy9E4jbH+fIK0vbDpAwP/KJbwxRxoe8HIk
up0hoGEJ7optLFc4axDtwD8h6Rrc39q7VbeZhVVR0MdC4k0s8wKeITq3nzKMoDxk
o2Bx3uZ967toLBbtiyVAWQrK3PN20HkASpjVLa3XkEC/XAw2PiplehQxyt2tqvtk
EoruXaqM1N9NGzRP//e3XVoELu4AX1o3ZEJjW1YRPttiQw+T53MKOsvgWrfHVu0K
pmaXLJOawBKC1586Z67n+byaOID9HebAlCfE1UrCNm8YAEVxFFbVvg+gDeOKg5Ta
TK6BXlGX1gFPd+jETxGCrO8QSh5gzVZfCSwKDexO1Oo2o4ADcyQ/gNtAsmVhrJ+h
6+AfDcxKLrRFTyCR+2QH7VOkzDehKJrwvHGgs2ttBw4cxJbuPCZ1mGzdsDqnjYVb
wM2AurHAkoXEYw6rzT7LY+7WJG5L8yaOzqU0CHLS+NIUXSn9J/yzWLxT4OE/OWmS
aYbyw2BVc9roEEXayBfrHblxRh0LizkUow/F2sMt8gb6W1QysLHjFlkCScg8m8si
Qa3izgie5glpdisvEjGqj/5Jqd66uxbPv+XCOZPRgEIhUCohhftuOiBzKidpkQpx
doSBM1p0Y/Wj+SeNHN8alblzKKXVtOKZIT5E8fK+zneSPA79bDGA9uLHlb5dQkne
fJ8W+gpMFO4nYZZJNClt/zilu40Wx+xGgKKdUW6yN+7oHtqECEAdqOy1sx0DDsHn
k8C6R8hnl99j2xZAqNqBR+aQ+G5fQcy0i47MBJb1ZDBw56D7/WX1488LZav4sQvM
z+yEx2t4R5VhZxdAq4phkly4P6kkgt8UJ7HTkpjRrn7JEsasE5NSlXzOU4nUWNsG
Ndd5yDmICbQYHcPQxRaua3Xq6Qtdg2mA24d1WALdC7yfJEUwJYfPaXyXrv2MTjji
WVa3GO1VLghVugrSMFppFucw9GdQpdj8+vI+qF8OiIzKeQghACVO1pEKYEFyRRDV
U2id4YDMJ8NyRiENACnjoufr/R70T5I+PvFE8ZlRn8+fcf8NUhbZme412Wwl77XI
+HZzVkbpvJEhpPVpRo53NCdECOmWdFVt/NmvzriKg/hck9pMTQ1KKaydub/KqA9q
kwypvbTj25GJxt6lxuYlfbEPSBAp60C8kUreMSa2cWKu6eercgih+YitSD2TzP46
ZvxokNb1UpjeyJMa+1ry+5uaIc5qPylSlKM/3fyaNOzBZCn13/fbkI9i00koXyvS
xxNu5/wi+lY0SEyMtzP5DVrysMyDHVvIYI1yAlCRuvR0IxMedVTgbcBb6MHgLA6t
LivsDzN01UjPoe/OUEZmNuM/0GUpA3hr6obVZ//X2DxjX4UgmEhhYXJA+CVqzv5c
Y8GaSQsKSDvfnLcsgH3p93iGLV1gCUPOsdZxPXqF5yJeuIvGWqFn1xXmFYm8yZ7U
GDYkfeu2j20LQwBQNXPbhHaa6ogaX0jsab3JXQZv/7lQyDl6MiTE/NIQDDfwbJqa
GmrUJCH6Eq4SeblfFIGJ3YRpnExvD16t1pYkhX8TjjR1dBG9pC1MmZQ0DMuLv08/
fLQptfeG0M3UdQhiaFXUBr5aswveYtyElCA2d6jMRTXb6hPjt8GmLUchXB5Y+oxM
I4I2NCyYoPIKKrFzqH/iLHtImEfAOyylAb+zbVRZJMCxpFXymg24GXnzg4AWQCAM
l6YeqNCRiVqPa/2Y+Ri/Dn423ldSC+nqJ1zHJYk1tjdz/KehMt4owt7cbP+jqVru
HWtYF3esFbVT8o5I8bYhKL0IbwpNRnjNXCKG4jub+OUErsD70wFF2bAWXwZsk4RP
x3CBBdy+AF1vbS1CURzJ37sOhg6oU3u6Mz6DIQmuvEZBYir9yzyRLeLRx1tT7Dyt
yLC3JMFq+7JVBEYrTxh1r8q69Zq7/vmsvYjrDJDDSsbzZ/s8t0SeoXdW50s54lBg
Y/e+fn2tc37pk38gs7cVqbbHfUwjQsT77Ad5fcXU44bVqs2x883pav5uGTYB2T8r
ZugY1mbVqPJFzz9fUIPN71yKQ/J1+elhgfJJmRwYbNM6ztzzYqjB8H6J4I6CP3pj
h9JHJcVn8LLllIPzFHOmiKxrD/ll3aYbkTwKigxEM3gZWCF3NU24FxAYTMYWhu6C
Qng7+xaGHe7iDu0Q77v3syDW5yJj6nwDRUQWhsCMx4dO1NK2ZofkD0Fi5HIUvc71
11vZ0Kcd7M+m9QqZ1GCF/6qTQySSq0uWxGgoR8Pmb/Plh9PXT9F8Q8sSe8ETMyTA
HSYMnHaAMsALmBkHIbfpe5fgQVfEcdCTmvneql8D7XRXDtoP/2nXP1JEDwodRlIE
HncOE2fUiHvT8ze10dXL0XH8NeYcOlU1g1vtkyPfVA9pn2WQ97JBZX+jYq3uc+Qi
gJO9knL/dvfnFof+Jd3AkwTmtzy+XHSsh8yKgkXLooeAJef7O+yrksniv4tkwQ3s
ZM5kAvjfymGSc3Fbmr/yDSy3/Irm0O4HyhTmbiv4bO7YvR0itWT642xh/XmOQq/d
zWel73GEbc6NSDhItEtjFaZg50cXFJzUwKJwS9rv/DxIK4x2JlPfkol4GKijHVkY
WJitJgxvkbY04BsS+6T6SLai1YBMCg/PFlb7Pjdzn+L2kwY4M2N15CcTb13YBMKP
COtGo82qWne1dHcapYP+nnpuLDs4l+VQDALTBLV1BFh5V7iPlDvqN+4q5ep3O9fN
tIvCeO2R38v+omzKGL4yXdnz8nHOrZv+TkP4kuBdrvalZlyLqg9m4toJuj1DMILM
nYEAFvNSxB9tIBbJoMjnbDxTBOzNS6ov6040gPh+w/6nAXKpMVCRZ6swBWvqbp3E
HuBuAQ4Vtnyd/6wsiULFcn30sIQ/yKpXSvTHu1WrNXJspmlTLKg/fgI0HgG2jMMb
y4RPZpxOha9bjPrYvIE1QbsMo8Wsh+y9OJsWppG1tze6hpHdd+svgHBpSPB31KhY
4tvDVcAEmflEQnzk82s0MZlFhjJPCqGK15Jp2TlMYc8lizYF9FeJtXZXrUNP7SaO
tOdg6RdTzdkJ0IMkzhV2zqLUjmQlwALgJ1D7CThwIJjVs14rOqZuNYW/4hyFrlU8
QeR5kB5PDGx4fHYHMZhAAR1LlxGUEkmc4yXco15Fw3peUja1qHdzREMU6Nfkex/a
8VRa9s3WC8kGzh8DFzGf7WEz3MALkxMYhcRw5wPy6YmRu26ezbALwTvdBliD53gK
tZ2AUzxv35Bz2k35XwQmWMgqyC9E9sk96e6HJZ71A+7HVZxz9TxZucjvP1IpIU+d
7hOymv/jDirzwGmPW7UMumqT/7Utg7LHEvmQq8e/wBRvGWJ16d8uukNRbvCfveFu
FGDFMA9emZKZZr+/TI6Vv6I/+6HjLdCXNxhkjOgsopsZQMg6L/lYFrmB1laYLzSH
S4Tw1vTeJOpqTRSXElMj0l1b1qi6Uqe+Gy4PW0kdzrOL6nUProQFr6v5yDejX+Yv
xmBjXlnWQbX5Gy7Qg79iui8F/WsWHUOyLoRo0slAmM0Z3hU6hHNaoWF0ae3dtn3N
uJ+hiy9r+a+Dm34cu0tBBNOBDJ1oCkyaKU+QTpPBee1knIYPiMhpqBUUa1L0/ZJT
VaoGss6X+sgkzYOjZQduWGU6NyJeVQF0FFST/cKGnOc/QMupYWruUpLeWWyFSPF0
A7Ie0idTsr6TZFDAYBqg8/4C5E8EnYzlUbMFSgH5Y7Tr6e3C7ESDqJbwYrTerI7S
nXxUfZw8FF6+/GTvyo9D8VBhDBnVOKSRWiDvE2srAk4RhoqRnajR2ch9J7zjK8Mo
875QT5YDRRR5BP+uOL20b68wYdpyTg7uBSAXJR9xoQHv/oc7nRgDtR1ChqdcIi+P
jKVJY3zScVM6sMH2+xzj/gu/nLBkR8ExKD5Ry9NJwlTbXWStwUV5VKh32eiKHhPW
wQcyiDV9WVoBEMfc2UOt5iCIx1u6qkmxxM1QbAUkNxVrDS3vZfNnAB/g1PgToBtK
fATPhQNUmdnxpEaGzIKoCTQepc45R2a0Iv17LAq6Jxs26TXWfUFrUYCAtmS92jMz
+J8yXRbkl0T20ZP+xFhyOJfsg4KWqX36PdZ4WxiPmrSl2mcD60yQqn7hX3gU+HsU
iVl3VoUeJg6V2NUWNc8mwQ5qBqERCtgs4vipbsYXaV2cpl4iNKhOfkuo/mwVrH0P
VuYRWPx0RAzgZNGL6tWi5KFdgUtMiBzo1EBODU24Sa7/c5LyBpNYW1JgtUB1MSGE
EInn4XIV764z/TOjffjPvVznWsKyoZwKY6dQuvxXf6mNRllTWYS0hf+rU1vde8OE
leVcbLE8TfIsCfrT2OSAUe0LAts2PcQrcaEl3cgrcpu4+S+dLKi9pAF2rnK2k0G1
uU3FvrCJBgxOMkIhpyQFkTl+AdY9LcG1pQ2vJCWClHP/2fVni7UlK5+Q2VacFG6B
eovgu46LNaNROA2L1/oJEuBcRn2inxkdrs7bHcsXEint+T6sud2cGOwcMYJYc6TE
CXoDH7UmDjat8wnTgAs1XzJpz4+FVEUV+D8mKOUAljEfXO+G0+TbnYK1oUOlyv/J
B8y4Kh+JpnBB1WkjgHVLhibeZo7uNcQhn3M6wdAkEr/LNcd/t2nsjTb2uOipwbMa
HDSZgE6U0FukJqjtioeURxDNqy35Pc2qE47hMXh5Bkqwb4ncnp2cdjxaLrVEFc3H
MGSxkJuGk1KR53JYMvnN7ECq04wTipFQKTbklr5zS9JVLjthbcIW0H0GjT1ouDkC
X/Gxw3WfUYa5aCuAKQQNJr+cc1MiQVQR7hjxo6ZRtCDcYzJuh1A0syy2XPoXFGaL
VDdu7rN98/sCv8+PkFrB+6+gTkrD70XUcPj7eAukRM1ghz+1Wy6nmv05LJdYB6hR
QkIUzHJzAj/98a1ckJKY83eFKmDS++CFUCV7VV6Pccw7YdB4i0RkPqAhkfhgMy4v
h9qHTJCB/PntNcd5yY/xfSArBrCNxEXUZxr/mE1YOVCoF0F8i3d0acRJSnSZ/NEw
BegEjGp/6OUv4F+5+iEpAoZqxENU6OvSztT77yr2nQyZ+/b5W1dFY4KhP+/Xemdu
mnX/yXEKalcKr+fBhVPuKzzRDtYSPWiBJTRVxXJdQ9SwG18/J4qpLJ8X5u4SnzOG
toRzcp4EX42P6HIweBAC/DR1ZCZLB4bnvNwrTtCACSRcXWxjK/ScB1YYIxv/dC2n
RD0PaXGoS6YRMdn/O5wxkqBTwg51wFGXd6sXMxHs2wVcfS+M4cU6qcnJGZJS04fv
7gffGa41ConoZOcms+ZIxnURtc+oT0v3bjP7sWGdS4eq0whh9hRI9JDyAH7NGUEn
h4QxkifebPwK+adckRZbofE3+mHcwOEjBe1/IISxYR1l25HghKNTYHxvLanohtpm
dMRyhucF3A7m3JBfPbjqTtHK8bZvUQG87PrUPJLi6p9i3gx6465f8bOZKv0EQU5R
O2vjWzZh/Ru99Wkn1qTaHd1uhu+0DrOh4M4aH6Tb2youd8g6sNvihqOA0pAyQCXj
u8vEWhNNNMMnEDm2T422FgRzqF/D4/pgLzQPuAP5klTXXRpUftVZ5kiLgWZyhzfh
2SlfmQHp0chCEk3mZBvai77amjkzoaOGtnfrBCIRhEfrbZFL/C1EVpG2KJ4hl0x0
OdpdBmVNvNvsr4ZmxDPslqPmMlJnWyg+zbcDPNW3HNYSdb2tsYLjxo6vdx1Q0jgN
9OGD/19R1xxahjyP9hOjq6CBA48yy7My3aDSsbk198wKNcJdvY4Q/eAQxvGyyXEJ
yXHZOkjdS+oYxGr1dcbVp4zLnOSDQ4n2DuUZlModgBapyQzkhJmX1dND/ltFw58j
RySF98ub6cCHgvQiFwbO3zucFudlb3eDA76DASeOjeI1EnTpZ9jONxxqnbuuwATH
sdF+7kcWqSp/3DnoSj+ga+A0Duv42vodB+8piF1C0WtV/kA0jBaXW8YPf84xduk8
SVyjaeYIvK+GuYsJIinn19ftDIfXg3qmE5NF+Y437FpZwks/MrMDVbPUZzglXEqL
Ahe/on/DoYsUhPpxE7SA10uXluuFqy/byxi5y8VpuJnFlnnSZcPckUaq52o5X0S1
FPP4tFf6SI7yarnPfP7B+s11b666aL7ziTrUisvRmmC6xhqh4evVkdWPHAJDG6lo
BQO//lKIm6SVyQMmEtQoJCrS7tD/zD4tyVc20oNdiW7yQx45EKVnrtCdXDlhULdD
6ddODGXVO6jSxnMcnUZv7qESFa1q/Y+oOvdSfbBLEhnsdLqrI93ndz+c7MB9OzM4
Ri4toyjy6iwfghD7HiZAcBEwj2KFqbm7vgI+IjJZcmPiRU5WPHS5M1bPWIDlHR0Z
XHzUWjAaQeuKExpaf5C1oz13JqjZdBCxMbLp6KJhdl8dbXrDVGKBeVCvAkNuqIP8
keoHYDL1a341BX8O/W57CNulIB/g0DKEP75CjveR/vtWobt+Xz1z45u33mc/Iegf
+j4Jjr04L5wHxK5fl03SgyB38OL0S4uFFdvlr9IbnohNNOqwOWlOTXti3ROT51U7
7zt2wzSdyjnrXdIRpDvIB6Gngjb0LmoPDCcElXBJx8Huq/2NaToT1SVhiQ26wmnm
tXz9nhyn0rW2rnJf8lpNLwpaBh+CSqQvyxPR1nIGXd0spatUBzyLocyfB8XmOip+
qx7sK3uUSlqs6R8jsGgqIK7J8GKcYeU/PoSJ03G9BSEZIoXdaFuq0Tm4Jub4OW9+
LVVCpov5BcIIxUzIYjY7yM43ZaZEExj4zaJiNYntMtTGdL27pNfRev/XfCgt5S/T
LYQ1YmlJrvRFZ9UfcQ+hKKt008TmObsC64SVc+ko45mXh45a5NBPhg4y/oOKBw89
XXnTY5el0YlhdWxwahh+WzZBlHblw6x5gmsjAL130Y7MhsgqbamAmAUuVQvQqXPX
D76oBCo100+ilib5KB3v3kuJHXhTDdC7H8RqyaJyEgz/Yxtxye3fyjZCzplsJiiI
MyLgE4uQtE8VDigfmj0K4DO7NOJIq4+Ju58b99oirPAf56cyCp+cTayZDfU7oeR1
Gj63P3pZyKvmd9ZAKNPtUS7PoTSVGGKsifGmrv+jOD961zQM+RSFJhGn/Nqvdsia
NwaZ/yXyirOCV6igN/k3skY01JRUv93wvbt7RmJe+OTr134THANvlEJ7buJT/NDR
iefA8eUXeseIAlSf/Vd0dgJXivcq3FcaOQ7yeR0PlR7NzLcLaavP2wgV3UK7vWJO
zbvqucK8KYhZ6q7X5qhWYwsEP9P3hqwycs4jB1B0gdoMjcEtTPzFolrgLG+MC+Ly
zFgT6YooZPGZzdbh6u5XSbAgLRlefAvV/TXtATwqwyS7u0ehWUtwk1YgrerBf/hB
LbhSfjBEkMh81UFPWv0nE+V+tatV8+0KJ8Ve1x3w5bCI/jXY5QlBj1FAR92LY/8C
solgSoEu1XCnXKcqnhZz2MppKJk/5AsQmhqHEetx3sdOi0wmSqc3QbGkbF+836u0
vx0EvfDWroTjK5rRMVohom8a2vLZBJZURSAT6SOencVHZF41BeHEP2LomFS0UWOd
furYrL7lFcapxSjnv0HY6XBXKTHVETZyBeyMVFqrrEbeNsyRgN6o0NBbzuOinZ3o
jkVnqmuzhoS8JqSNiCqOhwJ3rvLj8334Q4MaiOFeYZCBLSBKwglTLA5+D8NdYrxu
5ftUS8Oq6ck2/CqDa4Mv5GPdboZo80FTmvoNJUObcaOHRzY3AGFjdglpauXtxpi7
BOwY6/9E+uwuwCYxjyQ+M7werX2uOxhYV4vNl6LwLBxlKFJVrB3EqqIGlq3HssuW
xBKJJ6EnMr0OREU19/UggRKsnBzWLTsE5cUtz1xVSGWzF3LgmYETtkuIHV4XpYrP
Y7upSCNWaqX7EKFUakgwSTamMAeUYcq9PY1murWZPF7pibEsVT/rDDSqqfWYalJj
gmPOlgHigZWuz14KFGpWzUBmXxYx+cqP2r5jrYB8+EdEt4ONx+C7oqSNMl1o3/Nd
UAC/YfHzCM1Wqk2dd3MiKzyyttoojvYmwgg61GWFzZ1ZxqZ1yGVdCybq1DbDGmnY
wBdFVob+sD7iin9EUBJ6NHAKc3L5eVp0dssS5LpnX1xhU8N/Tz8GicwEBvEbT2xP
xqkhtGtqZmrqTth5OlJEkm61pOfEh5UkBjWp9tUx8e2k0T8Y7V6b9qXU/Yxv1WoV
QKABtUdTLQBWurV2h7yqyn8uShteH0AzyILvipSY5kE/+Zsrvux2HUbfdiM8dkza
pjC4/oD725p1bsgyikf0oA7/A8wsIgCWnCHW9ADrDDeZvV5rLa5oAj8yvUzATJY0
AgQhA748HU28BWQOuxpkXq56KVEc3eih6gLEGRFp9DhOpMkogd0hsFeEC9Om5xOX
njHiAfqj53fPg/mXxWasFEEwMC3q7WJQ9qSNq8Bdnjkhw5eCG6VQmFVAz8VP6PpF
zdcdR+9qW4cAcyy5RMFqSlipTo21aBWEJO3w8vhVlsZ6pfaOzNBMtqwxo1Sl3pBw
CCTdVy/kSzk4DgqoJAV9VOQq5VA+NbsjDI+myHa/InqPxDttwmXZP4JhzQk8SBz2
gVXYv3fQqS1iToPgfWxyL77wAtbrcsDNbfE2xMQ2gpAp3sUOJeyn+uu+ojlXk/JK
0m+TvT5Pp6eMOOBFszt7AJ8+pXhZYQXMmGgiavVqdSK7LJV9LLLTCZNLz/xFXXcs
FC3VOWgoSIesri98I6VKLMFGSO+m0cVk0SFtLNTulsO6Lr05c0TAszs+8pFrPJW3
DbXQEREXdahqTp5zBz/m0DZN/xc8lVV9ScegLddThxFu6zzda4Oj0mlffpV6JyY1
/1hNBieuqGNiieuzq656gCpyTORzE0Bq9Z5cEvoFSw6A0YA6kMRqgTS2BgXqOC2I
U4pGs/vCWotK23BB6wdVroUvzEn6oETLBmCQi02HTt+BflH3jf2PKMyJBGgDzvgX
HFwgkLkNMRbgscioTInmMG2WWyFqtWW9OEKTbs+egpKVNsJlEDqOvGAL76crvCwG
aoGTZqszS303dZjN0TeMlKKOzRq1OJuYa/mFg7hIEPFE7Vdnntk/Txu6OVyFFNeg
N3dHOJ3WObgPBttxEx8q4pU7c06JNjDQJaGXD7NmYF69l0KNXoU2ShhG0j/Nk/b6
GIj+Qf7jiIJryCedII3f82CVNQNaaoH/d85JMrJVSLE+w9w2gCPu4mAHHB7bFxN0
TV2nBCwPZa6Wm54LZRRBNhkL1jhA+ZAkuf3T08MEYhmsx5FwE1AQqYhQf9OqHKbw
mat2tG2I4Ghq0x64i4c3iRDDkyfqEfXjAHkfYXiBYNWtdS9YfxuopIzkDUBXWG84
lqfIfEgWGxjNpJa0wmSVdM/T06R/ru6F76m3oBUYPbDYk5TtwRKQkWcMfiNAvUuo
mk9hAnJPzBGeFePHowO+0bpPGqS0f48V+O7moGrNAVvpBNdAfkcicmSisw924xv1
44yX53xPhj7nJebkijDJL71i924axw8rP1q31NoOioz5Z4KhaPe3JUujFhxnX7t5
L0V6cCZng7h+MU52RVv+FklCWJQi0OXSSWXJ2mwxHimsjyrKZK6E/5lsgcxq1AYM
OypMlZ5TDDRr2JN3iRgs/eQ/K0jRnyT7go1G9YLgTL6hNcCg4d/MxAeE8QeAlrCa
JXHCAfG3mcKnfM7KK5OGCNP0HYycmn7hWwxi/dWhcoRHx4PeEpGBb0qeDMERwBw2
tXfw3Qykz5diZfeeqm935FufatOXHaIP0U0l9XEanwOOZ48Ayf8RU+9tTwSJKubQ
yYS/D72oWBSfyaqzIv+0RBg2hOjdi/hZ2R22D34d3rs4Oon4ZIgqYSS8yNWxsAzW
aZ5hZVd734IcoubvMn/uNPZZX72uhCfh7QZ9CawPfMUV4Rf4t3pAVTgXrz54SIfz
GKVzEzXN8grScQVY/rJ6UlmBHnRz05BoTGdN6jM2WsvGiznF+vG5c5wu1SjX8OId
A/2hVl0wGQQlqQ+PUGVA8/5K1s84OcAKV/0rUmCDk9mvQUnYrQJqaJrEkSVQqcqN
fdD6AkRV8fs2IS8iHo3pmqGZmtNACfU/INqKMDD07hfikEk2ywFCJTrDatdP+rLO
y4jrBwhUt5kdLDDElrnrs26b0PFMAXzQjfJa1utanCxLrb2pV9RHW/L+5UIDLGrm
k9Y6XW+p2LQxUKvZkZVU3W6/eXv4QwvkGW3T1ZXpnHnfdCJG2v57Mtc6RAPgz2/A
GdqAqHNaCZU63FGy125LPBZZ2HpASSVj/XJpO/KKOGwEMFQChtiOxVcKLG/LxRtE
7zQvuLQj7MpjmsYiNE0cRcvM3L+vNQnkcKRcisYsPTuqmcTl5Ish/N7ESEA6hcMs
Nkw8n8rBRUelQHZgxWnm5mod6ydwfH6LEMYZBQ+vAY9q5u1+ncMSj+yMKhFSNk+q
7xJ+qIZSOnsFfr+WYRLkR2g/1jIjthM1W4fieJebqjvkSAklO3pAOWiLH3PbHcPk
Acfpp5WvTyT8mx3e684enK2NTESDmL7omET9Eoqma5KW6hcAp3IMZdkug5Yfzv85
rAUbaGsolBYM/f5FXZXblJ88Jw8nYg6QyoBqWOzxKGrsVPB2GxGlFpo4NlqPksnW
3j/2KIlu6x1C7m/s68LyLNiGT2A4QyZys5Gm1zxLdh8OXBSu+ILYSra8w+odMFif
AFgH2swp8GxmxU6Qg++riNNpJGVZnAItbMDr+2mfMffE80iPQAzgUPWTc7yxfTaU
xoeuw3rtPWx055BRM+BzrrtSxfCwuBdW+d3Y/Mt5VOVXZT78+QS//4iCep5j8lRn
WqZxD/XvaS0Pu5pNEVlFYZDkWZA6MT8i4jyfSvM1vxL/nWyemJlKSGWpGRs/4+37
ZOVAKWZ4oJ2A4wawf6ACUvkZgujh6qBktTL+4QNRpuoHAmotocqpbV7sD2r9AcUV
zGiav7sWtYovjhA4IMSSS/raG+ZPYpN3M4+fJQDYsdyUqF79/ODWj1tCxplSIEsy
dFPX8Nz1KQNX2nfafMKJYG1kcRsb1I+49Koc2L7IkcrKuSbPJwDYS1S+YThaiHV5
dXSmuCdNd+ci/dt/Azla8Zh9KW9wpfSMtEyhUW8io76VCSzOcGTP5ZQZ7tRoF7dM
2mG4wygJSzxOJFrtjF3q4N+aVwB5+4l488QMgNvmJ0DXTQI0OyR2INBpjc8GpL1S
9TJl/79uqGUjfW+UDTb86ivm9eyd/19Hds5hAvxhV1b2VICYz4w3r8ioIOkNqbeD
q7RGLmKcHQAXtseLLSvcfkYov61rbOX5j9spYCFPLEyWUPQE1aWmuJH0FOm+MTuy
kSMSc+SKH9oS8Ztg8CHEEcSitDJDAigJ/BgR57T52ZCN9ZnkFzn4rDHDBNURYINr
uVp7ZOPnDfYGw/ZJ0uFGjmVD63hMDEZ2+sAeKxYf3nempGW40Nc6ORvpm9Na6qqI
ECxwoGsQLaE9TfmDxw8G10kJj50Taso11a89etMKnbCzVaxbK6+N6Q9Wr2vEO/8y
8MGdDRcdes4IdhZnMucKS8ON2KG43hyZAEW+UF/X8RdFaIklujOuo10XpRjM4Pkl
zWTD//vQ6+Ezf4AFxn2xDNaUY67fzAB358HtLvYkCuCExhGroW8N6Z40JgcUbRVj
iXgDGW714Z97I7doQN6zGay8i7j0pr9O7k9KZ4F/F/MdoPKjjQba/SuaTDd6Twwq
7G52LYQd8Dqfkxe+YBLiWpNbyQgr6vsPLZFpWZ8f7vV2DaJkde9uUJf0RGtRrjQ+
86RkcfXoAPniOFWGzk6iQ16fUdij3sU2CD2qvY+969tToZFZ8W3/AOFo75f1pPbg
j8AYM4h3e+pkIczcnvp0XKg6F+uTkStGEhzPGVwQmZ45nE3Gu548qasOER12vCfy
/nvSrm93/RVG5zweyZWQBFXRqoN1b2BqbbHUCmjYooO/huXLymsh3pv6K+0TKfRF
MsHrITmyfn0tgcMQPdkgcmhML3sMHAycADkjGDNGRP2gwPkfp+Ik1PlHz+jsZXkK
QxmdwTjTa9seT57OgmM9ZVejPdNooE5+TUs+SmP25KZRmWp4FrHGDfSXRU60azad
d5gyd3sZ6pjbhlCDQ1hT3uZ3IGk+0Wvs3qB1g3RVDORm5d4JCRBaW/FRyLbs7G6K
Jug4LbeLc/vdZE6niiNiOLItPUnn3JVgO7+Z2yphzU0JREW+cWfStw0ZO/eptyq1
rHKoGaPBf1HXv0qbQ9Ap340iWgLR6H0NP8dF2zn1e+ZRpuMI217tHzDER/okkSwP
L8rGZe2Q2KGzG/J1Z530BxKuGjKlvujN3zaRqksj3dEr+/ftmQpvoZXfZefDS4/K
71ofKJnsX/lCRsWefK3VFyixysXUCR7YR2cq0jY41gXAU3rN7PdhRrTGymijwKNi
uE9Qx4KDyjYhb/x9KNYGtqUa5LbZrswh0R62dmwzDw0rN/LMV2noA2gDoahU8Suh
x3VRN3mzODENHD+MFb2wGgZwaqqxIkIFTJGAoE/6vJl1b92snJlCtceg9CdEB9B3
9RS+mPKLFcCPwJo4I6jYC0bxrjLebFP0RKOLpsgGNNMyw5L1dw+0G5U0tGRgT9lP
SI2rTimQrnQoBMVOxWtx91kTGFYXeFlVMHemS/ngFB/xHGOM0GborVQ5SeMtmZq5
4s9R+L1tRPVy4FVmKOIrvTmH1Vd0wjPxa36L3CEooLtUQCZEWJWucc1W2NeSehn7
cleos4zFEtpTbSIp5dyQXM91N29qWvHTI3kiCHoM6bFPfJRFd0CLrudjEnXwf/Dk
0QYS4OvYbyP7MikthvS6CdjKD7kE4323fwZnLZXfKi0X7lxIJ+GUpO44KVYizQYE
gdU6lTvuEdbwJKAgDSgwpWsu4Olkc9PovYX3PRJBfmzCg829oaoaPiy86rvI5UAP
Ralye+Rm6+0Jel4LvvR4KFMerx6s9DAoHBHlZ1wArjRi0rFdDqhX706R9Ven3jgX
htWlLsg3iDq2u+A9fWZ3/YXyWdkM6G/wHstU8+KtOTSQ+hFvJKjDO2tPnHkhqU35
n+8fI7RMedmYyQgVtqqGslouhfX50uWTAx5syA5KTEfFJaVObgUkJ+qaZmNIaNUg
W5h90dCpGmZBaR9Sv7Y7UtQvDMa6v7AH3898IAdWAmDoTWgeeCYY4ubasjg0N2Cb
88Mod2Qfr/t636NvpryhuELuXN2Flz3RD12Xj1HJutX8RfdyyzBIt2Rnj3FVdxrI
rdNx4OaG6y24aMagAZaVKuioi09DbVBmBB76SnAQ7gs0jx1D792BA8vFu8ZyTHqA
Q75lHOScqNlaNYU7U5FEEs7er7gWlStwIOjqocY4pp+tAoE382WDhLTrsM3mMDgE
m86PjTPI15+gKLPeg1g9+6gD1e4FxjBGzQ2rpPvwdFSoMSOhMnxnx4ixEjXmFS6j
S9sf1mqtL3JSyFR3u7nTh2H7dSWGyVbwHOzh8/ct/QUEJjQjzUpv7Cr3blRQpHvw
jpw/dnKEyW1iVvw44+HOBayJC+kfCTYiIMo03rgJJHIM0o6zc+wkKYqnQEO0Tnk2
g0q9ttVURo2QmTiuO7JlI/G1QwUda7OXLlZga4h/dpGCdIhfcEQSW6vmp4h5y78e
BcLU4jIAVVNLpWyzKwny1hTMaQ9Thv9ZGgUpivX/bP4K8CmyWzaTwOGtWfrMmVyl
R4C0jHqtRuG297WroESyte/Kbsz0VUQ+TJM0vU+Qk11dMNEr/9oPh3ayR3aIVP6c
oAi7DN4It267LU8q56zZM7iqM/q/IBzs0bKyB23rwGRJ2lVeVJ03TzY8QwzwXBZi
18cdTVHTYpgFxc5bdJfQIio6odjFiQQCXVzRBmj7Y6W6CZ6ZgUtneklqSxUhsgYs
2FBIM72xp/Pw96IjTsVvTprlpvV3ccvrQQNLpGknAe56x82LhsilTLgyevMB193E
Up40QUX7SZjNvwTqRauoWcBzH5+vk7u37x1jQ18lzdABf2mr1mycaouuopNMh2io
IcBQA9lkfp89vqbRssRoBXSHbqSrnIHkDvWpXGp839Ub+dRJ0FQtlq4nVBSTgFEF
BGeTlEmnd8ApA1sJ8po8v5z/iJKsiYijmuxxKfTnFDOPTr4N6uI0ot+wUhAMM9HH
IgEorj5eksN//rOBqKIQkjkN5p64CZurNc7b/Md6SQg3Q1Qxz4OkPjG21ezPYmZq
ZL4wvUgLuAiDzmOABqcDs9LOUWkwBM4AZ7LS/eJIq0yswyCqPZk3c8FPWFiV3i8u
UUAFxgLjpIJjuXV3x5CVKSSfca6DKnApXjKcPF0ToipLfWg++Dqhm2hEGeTrtMxq
ozcoXoyRIaPXufTAu6S41EOZ8t6uLPCWkOf8cZJVWIGpoDb2rrXM2yn+YMTs9JEw
xwE6PZQNz0F8lbyWkjoAM11SQdlSDs8ucUFlgE0ljLA1dMmqPf18jv4HJQsO6hJT
vYmzc7iWSnr9gBe+Lh5bCQfniyhdkaTnP5e24X5a/YoaintghG4wW946lrTKTCQN
mphqKlflFMW+cmLBt0wSXgSbeTE9MEQtBpu22zHWce/RUqs2JzXsBzEC0SDHDWbZ
lpnHc5wYviblKIV1T/8mtxEZ/Ku9mNY6o0tgAMtctvD4CowfxtJZ6VOlLX7yBS/K
sp5GKQ7VuNqOr0P1GKTR2Rn6fhP7FgmXPFVEnpZen7azrp0ibIml0zyL501KFjJN
Tozxw0g1XC15SzqYaBtAclSu371YD77NngY3Mvd743UAKaO+em1P0cd99LCnzy/8
G/tY6/HN9UWHbSSnvW2O6ulCTyQJfJAXtUteA3+3dDfGFUNN+kd4NlowN0uRP9JK
4GLytjrLDMTS8J4auMuulINfMiZ8pgDSpy1HS6W0FmKQ0IfQt96uJDU01Bs4Vhgw
NuxYoqHRlVmLGWzH4XMjXUX6Ffxy8cVQDGWwMRSU1AtM+lTU/LZGFVtMy9Sdrl3o
QA1GBDUxyGsZ6IzgWDIJSAjZVK6XC1I3ejq6BsUpBcxfVk7dP269Wav+iLHRKXVv
0v775tluKgVEJcrbO8qDbD91mXkbXNlV+r/CvcavQDmBR03cpK+lfG4IYr2idZLd
SQ1t6s79kUzNbWKj1lZaVd+Tcw2DZ6UgzWs9Ixo2dxKt9RVibxlNaiPOkgiqe1sq
3Q4Nm4a8mQKA1jarDi9YQvLA8t40B56d1xrTrx1JnwDyhewmgnlIH5HEWnCdqvyD
md35s++QJTJuY7DBhcthUIo628XoGWSwPqeEMXJokCyBzRoE3mGfpp8xG7a+kAgv
Eidoro9fkOIeN/QqKLDLz03QT4Po1rPK90NhKMvhqJUYIyMybFsQKiR5ibSruMPT
zZF1JlX+dzxzcctY6Wx2PoRsLieTaWMawqG3qJUaVg7osEKAcmS8+DlXYVtXXjwd
wgTE+li+pPUe/pi9hJ237Nctmnn68tIjEpS7lkjvAYpaKB+Haakm8pWqLyGWbvnv
EYxyxfWfWKcUqJOrSysIEOaHTo2Ah5YRDA62WAMn+/QaPjvNsPdLdsHSMAvjA8Bd
hBr0fQnWfcN6S8zbcIBA8RhVvsQSDO9t1Aphb93FEBMDghlIwOMTLUSJorw6PKfN
YcpxdUGDtcLahu+lLHe959uL/PzUZfj4LOe9oPIlWskimlwyvNwZt9sTV5FXHs22
qJ0hQwtJx5gJFlhVjXyhcFIXnrO4wHhRGHbAykycJNgOlwy5DZyKs/nBd1GLLL7Q
9uYAYT0/aVItxD8jEZeKfmhbyib2fjhrK53ZeX1O6bUDIa2x+T4VqO150kIWL9s9
QbtapwGx95m4plzSV262ZnBfdQPrZwf5lNdlSS4rB5INrNcNrnYAUNLDBhQmlBfx
6VYTliVSh78mMrG/xJbNKSycmipVUboMVnZXoe/VYHTMSs1ua2ea7Q7KbLd9BxFz
RjCy0tb0c1hIXCNnyOK1oE8VQEJjbRIZm5xgI8QhxDF4zLYH2+Q08+AJG1MrfQdP
WIsfR80MwcqoVH9MCDTQfXyRVaQk2BzD/oF0Wj00GLZ17gae97fT1nkCbeQHO0kc
xZ+Crlx5enrf32fq7DdMKLNyFPj30RWjD+ytg5VUZ9NCZxZb80IZkwZ3WvDdcetL
RW540QJ/a/F/90MZBCkzRPBSAlbVrxfo9R4VPlTHL49iQHBwjpBiodM5d9IwCHpe
TgDR12G3vC6o/maGkWhtpe2a3HuqVH0c0FqRqTPAfM8i4IsnJjG7RYBTaqPIvNP/
RgfLSTxDGVmsLHubb2/7g/qJa3oy39jjiWqipXKnSLF1oXTvanCDqBvH6t6CsE0T
cFdOfyTvQebyQBzf83sFvvifFCv1JdYpgie/4DFAFMo1ALY69FsAmzAUjf9R9Shy
ouhtgHfLQP38Kcr2GyC37qB+WdRi5sHSbLZ9miV/Xr7xkOqwhA/4g4BYXELCNR8J
XgmnIJVPo7gSq7D3Oo7dVE8+bqBisvuxiE/CkbTiyfk95JwPR4Hfw5Yg/H8+1imn
vCh57N9RMweRi8nly90pzKajuHn/t5o+bBWJDoblQwx2KPgry7u/dgKLrtegchHr
KAGP3tNb3pRFP+cC76Bgx9d29PvKj2EAjfgeaH2CcB8t4tf6a4jr17JwKyf4kzjx
QLdiZTptTSAMdXfsecEtGHtWNtB7hfGaJ/8pO1/+LE/pxOeOsYxnqk1c8jw1VQ74
xOBgx83lAj7u7msmJG3haGAuBGbcP+YWFjoOBpw3YWFSgNh5xYvYSyN9heWPtKb+
2ROs+ViWd9qluJpvBISuYlv5w3jvq29BLDk+UCHmwvF04V+9tL3vA+6w3ypVUZEw
D/carN+ec/wUEhjXYCwa7cj7knt1YFkl0oFYuH3+FOepeYpjkzJ1uqPvGq3RBuyj
AvYBfixhsGud+0pKmlKUwXgqQi30AoOS92NcwCAMaEUWvLWi0obudsYlOe1FMTpO
HbpWCV5XHGXf0K/y9877b4iIAk9h77D8xUQE3wmfdsbQa2m/SVa1p+MMg4cwHZr9
tD/vkG8Sxf7w/Hqw0mcwF1VSlmwa6KB9Yy3MwwvRyWhvDhhnPztynk1w0kdkYnOB
WjH7C8a+FBP/Z2MlP9n6xsa48GUTZmzEPvpFn/F12TsQwYvPRN51HvvgFeS3FQKM
MIMbGcUXWxOMfxyNfO+6q33Ihk8U85Vl6x80CQZmssWcjbz4hj4taysDhn/hI0zf
NqO6xnqbAxPiTC66v71Kxo+6XVSwxp2+cKQ+0T2f3wmneXGs0nlgss3WYf1kyAVj
y2VSUjb70gYF8mkV/PVPhBVJcKStN4lUhzkpFCEV4y/ohwiQTPQTVXsR9SJvNIsq
LjpH/jzIzQD4UFJPSaO4Z/J5wiMbSDUUt893KthW+ewLTJi5cMpnEpQUfSUzRdzp
Jp/rx5ftDWV21yuKY5ktpiZIS0td0bxhwxfLb/a54NOfMa0RienpC+TBV2uooEAc
1wSqCjQT3Sif4BN7xWqoN2grMRN3McSzg8H/LfuiIfjtDoIXOadm3L+iGogVGYlo
R9o/Jeak4qadoIEQ+lzpcX9tBnEPTk6BMMdGrlPLGcEGc469e/il/o3L7awNIzOn
ZYfT+dKzC+udoU1kNik6s8cB0chKVrP3r8b/0HbUJorVn+jN5DuQx8TDPcH8d3lN
3zWk7kp+RaT3+kAk311cNm4yCv64vfCzNmpwzuwMfm34p5ro9dPgUBcqldPrDyAW
2pNFywW+18wBZiKcRVtcggAgVr2j0ztBo/IErbL+5qapZBdKS2unE20K1VybN25Z
WtxowFVlmB/yg6oJMd9Nf4mQ+MGc+uIWFuBQ2rKBZbolBN5k50LSQttkEG11X4oM
D7F9ziX9LgNEy8sOS4ddnfxTgVF0tDAW4mQg8nyoYW5zVyJ20JJt//IKYOw+qixO
VAmllUAAcCPk3j2bSCllUG694KzLkg6Br6pafi+BWAnwv1QwPzKu3wWDIX4Kj/zS
IYvOnUj75s+EWfDfNiPNqAhF0JZ1s2tphksfvz1ZV/kOqndLS+iTXHdh7nBECWBF
v84lN0EvpoqsCWpHFMDb6pgkH+U7OT4+lj/FUMkaffaRu6wCix4F40X9kJZ7nq9b
Wp3/fzZtDgcRZr9RRPB3O5PVawEC1GcqnWG595tByKAGBE1KIYoncD+vaPIHbAfP
mWO/R4mT5kZhacKmzH0ozUqe0ZkRanu/tE8F/jPtiHPgpAXavcIGtgIFbmlohYgL
W+1zJ5YsVugd9rYoOJ1f7r6IPmriqyaS3LJVKHNTX+pvXZuFXbsKfjpdHuE//zOh
kKJGFO4B/MfRD8bYwvSi84cKLT2N8I6fGfU2Lt/1i+Rf2X+qSez4ntbBs4Rgubhl
pEouG77eaN5XzxTSBncOPId743R9sqZR/q5vXU6KUmj8S5VApx5bEdqgUz4b+zZW
VHEcCGWTQMdjLi/OWDaj4ovOCj7AGcxYSPEy2CS2k3pY3+zeYOH6VTTuiaAB1WH+
Ldj5ufJaVsB6zo0ZIg4NhhBsDXfdfBkM1NjAxU4NyGw2ULOc7e2lUVllM7kuhBsr
7MbF8w2vgcx6+l2c7V6H/hjD5h48LzZf1TKD38KDnimCd212naSDSJYYhe920mfO
jywO3oha8cVczJ98038y+43AJZPp69niayo5MXO4dVXStWEgtecJ0FQSlK+NzZmO
3ZdjckddWJx9qzHGuIj/7QdEJKTKmzl4UTMY6qj5/owO1OzVdvrosGLpwhupogo4
VLYzwTxHcevxVTE9eAPrsfoEUOoJEINepihgu6GNFNPz3u4SDtyCTUq0U0AY1Qsk
TDDnoA8G1Ps0pSsCDufoMOSnTzQAsUGU/uXGsy3LlxNxvxgn7FXn0Nuy3HSrlJf6
uZfG90/4bfUtN6vdjDkj8U/pHZU9l3Ch5Q6KT+RfpYuvH6f1enkN5e/wigixR6jM
WvO1aiB9rplTI6Au0Wm3oqR6zu2gFL0k0LDdJIB3xH504Pn34PrRbF055eA0dtS0
F9FHJTXlu+qkjzjM1R0W1+UXWzydjERUJbxinnNHkmHJC6jggkW2ezp7q2jdeAiZ
/SfN2lFVkZhYzfCGXZZkpvxLYFpea8QUbrXtfxXDnUuokLAYNLZNUonHntHnVbxF
Zk18bZyG3OoM+cj3IQw6OtSb2knmdyyeN8SAESCCOsigjzd8pmDuBnMrCFrOhNfg
pLNmX+a72zp4stHDaGSqBjdD6lRxkHt1D0Bqj6gf9femkCO2Y0KCn3v97GTNnJ3+
0AQfKeXh+uH8iID1VA7J1JDmfkbPkhtsZ4MpsP0hamWIKEW/f4Ez4HlgZdyRF+o4
nQRxutaYqPdU3fHOPujkMDK5mBjHJb/TOePe8U/QeEK1HheB5t/ULrRhCODYMa3Y
gSTmQqs2J9uo5OzVxgUoT8ck9ky7x93Lgax79T2giM63u7EjP6o0LI2Yqru6s5Sd
zqugJq+U98LMUELQuLhud5oCCpxV4yUoRCy3XDhS73OhcSmKW1kVdlpUQwi2aKap
VKcW1duIaW4jbCQLxAKIQ7k0KDFIacgEQJGjrlxuxu+qtIHveGXPYev66Rj+hETr
AUERrWbd7ZBBXZhQ9rwJ+QxFs/9hyvEVZ2zg9fO51NGKh2TOG7ZemUEj+NBw09lt
HvVvoHBRCuBWt0WwAbAv00lBjV7DsjT4SFdKl7BiQ72JzQnAhXpvzpHL8ALrGiMw
uQcWzIthXW9pLDuuFlIveCPP5S+YhI9Mz5VRpNuf93JTul70Uz0kCp4b1EWwSUWX
K3M+7W4kC4ZbDj4wLCsrkfxYOm5IPRk+Pl6y5FZvdiGKcoKNX9i/GDDiXCG7SSBE
553OjVFSsLo2/i7aBEMOxjK3gDXg5FNXh0qR4n7kZEmDzJ0OYXU9qL0mXUggb2Pt
gyD9kpIyvAyhjupewSYwroTmTtl6BHuToElaUOPvUSl5s8AJXGqQjuYlIQQHhZe5
GBNnSa5gjiAdSmXWOHI8TcsybWKWu8aLetmqW3tEmqgIDOGqcOZvUuzorNdCsOgf
4gMgf/nAmD7sKclDe7Ct0XrLZj0UlWKJFSruXEZK9zNZyjomR8KWCayenI4tUlHx
vupm1BP7v7kbVcVxaoZehqRNz0metOQt3ggjGmeR/xwgpGDcPTkdXMvGsxcnM+lV
HN6nG6x2AVq1lcS3GHUqz6Rh1AfPl+24TdjeGr9FXXaPozs55fYMvtWSpCpgNhVm
3GkUytyV6XVlAvr3SQI3SrI6JgaXTat3Oqy3ktG1OqISpe7azv8I1JVckkaLagMA
AVDpIUHgX6uPyX+PEAf9e+/sGLAH/9/GFsWO8dNcmA/df60Xs6aBjhtiiNLloY2j
AHzLOW53xndW++cg+abbUwpi8E4F4A1kHrvk+fzUlDIW2MSPrR6qr4tSEZILWqHe
DXa/3xfyr8ZpJvuFlTBVlAYAqDTueRSaHJ4NyzYfDlMTXBiosheLxnSmHk1aDfYw
uKrvJSrGiMuvDyU4KwFWIy0tAxeC1LfanS+p3xDIcYsFoUBUJJ9mT9cW332oafa4
QXJT99lsTtrgaisf+OSc3SyopdaGwlxqZLoQcw9R7QIzgAYmHSZIV9VCkzh9b9/K
9/yKRb29g6Q69f9aL/KsO5XnGTpQlX6mO7YGuS3gWjIkTE56Xf03deCGcRCgTljV
r/K2NLW5AMWK1eR8ilZyBm5a4mLIJmskEBcQ8Tlg5Ni2Vi9Xe5KLYeez9U7uOcYT
9SvlrOtYzDV/GiQ3iU/r9wMq+BbArNjzwzzLDrVxYGBSPa/rlzTtYCo+350zyiTb
1yrEubxldGcmGLDGxAoBBB54VOfXgFwAF3Qd31pEqIRXRNcpDChuJdN5Eds2sw/5
IHCcioVOupSZ40KPC5ydlQ9RSGhXFOrMu02h2zbN+9oya5XBqxWqEKagwh5QFHEr
i+YK18LLufKXAGGejyzCJLh+gSndAFOUdB9y47SO6czzFwHi8MCbQwX27HfNR3ZS
LP4Zr5WgYGN/GZkVAXvtXZabwL2528BNHK/SxV8SkU7Mfa7q9tk7XI+hRkp2OtWI
HWF9BHm/hPcPsFNRFLgjnm3oA3tQdSS9kkCtL4Cu3OzjvhOr7/6zIO0e+18ME/tm
shhVRnhdldH5WEukOq/i9B4hwlvhhhtMEHwtAGGnFtxuT8fBslfLu7RovQbmHEDK
e26husHD+OSnZ9qtrEcmVdzRa4L/+ohWuSxjvElSl1F78um/1NiL9yOpMZqhzLXj
cIUBTJ6U2JA6qpQ4XywMe0c4LP05Cm2feKguNkpZj6kWk7OcIXerd6gEVoHBTY4/
XwZtIzypie0u2D0nIjZib4akUCz0lbSPaescX49qodCXHbyIxYouRAes6sosz9I1
ovQ/yT5CBONUf6VH9myt2R6NwlI1NnxEb6JReqRCGq3Sdjq+3jFCS4y14xzvmkfZ
XCBnpq6s1yEZ20wlEOzPZKADfNDaGdEbg8YcgD+iEEkeXFyV0v/BCDGHCzpHpC+7
pxvF36ALYM4xuy7mhLX3T2bijyAKoSAB4FMPoaWgCSD0KxS/1OQ+Sj8xMAmvHrGN
dRQo2m5LydafgQEgF5ByViaivdY2oEZ/acJiHU+XyotW7Wa14ZHhtufKGvJEdlo7
KF3wfQhhmnA7XLCNx4msm+iWsIe1rHxJqmiDgsbGW2q2+UOt9b9SxsJsI/7W9POK
OxL9vvUpQ1esK4DpToKuoPLpJKXdXeQQpN7Dv3sZqMpFGXAtAQJCtLsbHijTDGWq
0rc6fsvLXcN4CqPqtU7odjEet+AFDqtt8Rj1YPGnIQBzeZS0WMc5Hnxx7aGlNTmf
2hrfupSQ7CfpyjVD9XPpXcOtUeY8b/L3Mag46uCs0/Eo6smubok8yz1MTfVb+How
XPY5Q0xc/ggtuUqa9mvaCJYIjF6MN+mzT7+60LMfZQW37X9/YS+WTZDxQVyVO84n
USF1RwcXqFuQsdzNPUH7bM1NtAD5sB9iq2gf3y8qeb3c52ITaP9HNx/B0mzeurH+
yYV9TYxIujV3lSh7R8oeLoDCqOMutnBofjGcP2F+TYQVzspYUOSkcbzzsnGzYa5Y
34vBucMTtq4M78TEZi9GQD5it0xYo2TulniOGiu19JEwf1d3zxEzW4ncrPAPTaY6
W5fzAZb4bysKC5GlvrwxoOa55TKwIMHLlqPca9ZsUlzkEiDL9sfo3vnwEUZtQyiH
e1VZeGE+tihPE/jFJB6oFIHwtwwZzM+L8NtvD0g9If1q9ci2W9Dqg87YC1KBq+WE
+kvpgJn8iKLrpZHdrj9HVGjL+2m+G0/FlmeEbRG71528BsMnW2LinEDBch1XJ+lN
XglKyxeRXW9Ui9OoSPDqivqaf+A7FZ2YancjEjTqaGghZdXQJMaRl6J3QU7ug8Ss
2M9p7xxsQMq6ElJdMU6oq/7MzUw9VWRopU792D6FWZNzMPXJ15fCP0Bt3fxru+GN
HyetlMPgoA+qdgint97eKzGvnKboWNynEQWwlPMIpdVtM2SjADpJdMMVwLe+MVY8
9/z/dQ34z4F9m5jwTroC9/fdUrZ/jT7oJI27zcJJTqURngTJSgRMzl9pQT2ME9aC
aRnwHdrjAKOivvU6iwoJKp3+ae1/7JW/qSwbhtVA7WCkLG7DC21UH4pX/hxmbyzJ
TpntwjVJLnGQYHUo0o3XuL+54TXB927C/HtzwaxBkxAbWyBxP+lfKXxgXQlp5yRX
O55pF2+8SpDmU3x8H10QCZTPVWBj6FaSXIsRCf4dVj5QgtZTGHYht18M088hcmYk
JM31fMKUP0LvauCiR2avnQL+nj5TMOW2UWFulr6VHLYntFCwo4gsNj8ldVsi3J07
HrKpGLwHlWsq2WhwCNF9KvY+7VkYuEqntQfWGL39UM+Jv0Eu1qLbirhHwx4NWuO1
xmbxIDsckGXd87ceP/O7X6FmJAXt4A2/mwr9hGZRbhA0f48oPKvYkgUTAj94LLnG
4IukN34JO/1CZlDHnm9p/xI+0656fn0qDdLOYrx0qvqLPo3a7LO41mIyTfDMQfA1
ZAptb2PoFv28/Dunw65pkfK2AwS9V20KACXZjWeIjXhv7JqrMdBFRlbazvJ36dmW
ryfrvjBAucoMlQ7Z+FV9O0r/zKiy8fJYTJqXUoIn9ihSl/P2rfAJAfTwX3msaHeR
tq0detZBfem2nIjFTE3eE6O9W6vMpPbDUkOSpxRugw0jmL0cvkjcyCU8C1LYtM85
Ngm8pe+48reguWyjQ3ltVPtcBlYqb5veZDHDQ6DiV9PenQrpK1SCxTp57twN0yhb
wwCLMcKfB36WVpnTrhzcSeXM8hijIgKGC5LsLf9NcxnO05GkpdAuAtT2kF7OfyDx
8L2dMGVHzcf87gkUMEB08xmyfioU8Mzs29Lk6G8lzu9U1dqmlqlHntfgHi/qIdQ5
kzy9807oGKdDtOgjcYyAoyJ0jsEaHxer51u+FJ+R+USz0+ysZ0uV6NIplvyaoeDB
fQYi6ECi7WhQ7Sz7BsOuuY5xq5RPPxFaDIO/7nDYdvgU3UIIU4J62S2LtVI3YPpQ
3B4njqNvXtrV3kVFdlH9dsziahKjmo37iXMgxl4H6SRMMuic+uxSSMEhq7OGnqjf
SL4/gF6GtjY3CRN5WhshpFHiipgQNbM6pFckhFa0EbHMg+CVYPejaK1JlObkT8Yl
aJuC2674Jpm4rYkC8eaesi6WrL/S3l4qKfptjeB/fUiIUU+s6kZbnIdn9m7rOgu1
Ed+hx+OvT6QgnrlTE0GUK29YJH+YM0Eny4CY0Qhv4oPmVQklREBN+WmSE2LH3bai
ZuX0QD0Z/UWBJwCU/0m3E5avHkZouYmaW0dF8PFVZfjO+BBpWamMKPY1ZsmWw6pn
tN/9rGq/YWYBbkmveJbAxHM30xUfFgSdPnekgtAlgRzR4GsBbd3ugHwUQLGRyp3K
nhNjXKqLPb2PE2xJz63aBf++yh3BEKHjg2KTC377LVzyC57b5jwY4WaJUNufAho0
+Pxu5k0lVIo7iIPatHIV9EBbkvr8EIIS3bZYvLT+pUAym4bwTC/q/DLP9vexVGPP
Sw3/BxGneREgEdckG0wdlELVShmpGbgaGkbXV2KaaFlSGldYS0jJxSDWKTZmqXJc
zjcCsGqbbX4hbjueRKjNIr9l/dzJNJEjl0jLI+cAcjEXszJtNdDuYWvGvSd55zjU
+7/s86ssvowM+IWkVa4efwYRIqkeSgyPNMpXKdsomSSWXqn3FFkNzD8L4OgXXGMX
JesvoU6lP3iC3AM0YS/WrTtqti3C4dlO4sUBQAhDnReJTa21jRMWVsnBaEIRSZSo
TB3C7K+qmerghpTxRzjDijvztNACyP2RmJav2Fczgi10iD5jKB02K+wdLC1oUlPH
uwSAwXQfpKK+0LP9OFL5BzebWqW57hT1puaB3FTwyi/KJgYOG2R9CJth6DTv/NXb
w+xhN5aw9h/ZiDgVISFW+ODGSmpXFL839RBAZEbly4WA/ufLnfb0VdZnhjuHmOSt
noyApgVQumFSlTl/kvzkUImaxtHvr6RPlq4ZiD9vK6KHQGrc5SNSHJOdw3AYuO7v
zRFJr9I3/FPLDrF73zrfIrUx6uduzWTVCVYeyZ8o92jhH4lfULUhI6Z6Gr6C8Ua3
eg1oVeabDMl+7HIIzoF4VgBM6As1sTcMZmoeJl7J2C9tVfG8cIXeKWT1tGYO/Rwm
DJR/ZD9FF6Je7/18g5jKdKa+3E0UhiSMpbVMO4bGQuIgz/yEN8AAQruWzCx6Zc8D
aZDK51fyROfCk4ZPU12W7LvlEcIXJ1cSBFwgQOpXQxZePjX1l29+CAci4SkMwoJS
Mgww5PRX41oRfQ1xh3GDaGxpOza8EduG01oh8VeGlxxe59GpsVTIerVR5wgiey1H
xjCAcB5HJl+s2V62lmoNsWdaSgsCftjh15mafps1H/w23LSDJUkNp9FORj3YYshK
TiFFvUj8y9lAqCnPCU291EohVijLptaFJ8xMkzJO8vTf8kDTWFO0GMjRiDVJUVz5
tzz7Q6JfV9IgQS0SXiDI/7Tb7mmOm5fZolfPrykl4NPZuz5Xd1m9eMZwLsy4jXcT
7aCxdAeQ2duTmNTrjPf+NtjbEe2jEAf0udKCW//4HVlX3TKo1x5lablkiv+bJ99e
fJ0Da5eg8kW262lJZAQFPDk0/5f3AJy/tppz1e9csXBGti/WzApYSV2Jxbu/N5qy
xnzjw+GE1Gy3mXHbMvW2RwOT63SDkSK2w9i02RnQd8Owoc2DPvIH6dElt3KkJvHj
SMTjj2xRbvbEEJ09CTzNKkfrHDjz5cGvtwZoEY9UVte+YosiyQwL0Tdfoe43dKRS
U3uzXVNUyqxLtDTBWMLHhnF+zHFptw37AggajhfD4ElgVeahxdLx541CbmNqvbFk
bU2JgtV+KIu8D8Et5ReC9dQJlDXfqASmG1FzJZd4IU3YfCLCoYOo9T0RwHS8M3gt
T3saboigDr/Pd0TY0LmFOsLl/U3ZrYxzFvaMmOigVruLXNbM15AGEe22oPYL+Gd+
Hru6L8SYViHhSThpyWdW/gq85sn6dzCr/mONly7w0CQUqQPpQKrjZ9jDvBldoC3k
BAO4K6jWqnZqqFIJOOV+l+1EMX2dp2RLEPIC+FJeGGwL2Y4zbYl/w4OgfRixHiBo
kHjfXd7coz7iRPpsRw8E2mVmQ8hZ+uLffXVhpchKNpY2fRQhgKr7zsEMC2ik3bvR
dPD0M3GZzTpoQczJe2O2cEWWQBwhEu9yEceD2fLPEHWUWOlLw4zsaZd2nTDkLE4s
QJZWWSQkmfgsBsLI1RmVyAGmboAaRQtnbxc02lxDnk+HvK1V9SWMNBhRsLFz3LWr
78jmGAbvh1plf7CBAVqZfPlhP4OwDNtChpV8za91b0+Tj5ZZvFI+HS0kZ+7V8VlH
H4c/9IQ7k3vvpDJRUXKc+jARtYKEaByzU9T3mrXyDLl49gQJqG4hLoDh6/NEMpHR
Zd0JIcB2QU6ayrbq9Ln1m/L9XO4KuPlPPmO2mbeIX96GPr1vkkAQ6vtO78+M9lAd
gxgp4E8lTO8zMv4V68W2wtFtXklj3p5WJGtseEVmjXYVMguKdUH0FF66PKK4cWoG
echdl+3xhTX8KALfI8Eb5pXJfbnwqdnqxR/Zo0lQxKpi8fboRibz1GpucfJUVW13
c9sXrDx2+hrzgz1xJ99Ysz9NCOyaLB1onx0aGIOwxO4SIB583YHwboGT3y/A71o5
arKIL+hTV3tqbdDZTE+zEiVnCODv8mII8xHjvA3yKj59VTfDruZCueoijMHB4tZJ
asCXdqa9FkZd0vBXGuCUNqq8KvF+MWPHpLOLi20SDgxEB/Ew+PQyFlJrZjx7Lxj0
LDs7amSakaUDlzaQcKSSvUU36qG5TWdr1QtrBYS9eg7SEiE2wR2jGz6x25tcJgpZ
byl58vbw0/HXZxNXBklYM1mmQK5KEhGw8otVs9dDftaj5ObuvWIpjiJ3Eh+RTCFQ
LX/m4ZV9wCKssKuvfaqbPKl3HPsj/djrLNcTak/jMnWvsDYGQgV2FaBPj85BaNQ3
bgBE70BgU5UonAeaSpaF5IXkT6L5sVOB+rt2mADKTaELKowle65xzf7IdVP0jjOF
PSQLkiI9u1nQAQaNlsL6KUGZHpgqCcJDNJx1CDYyXINsp97Pq/tc9nLojHqLIb6W
QMFkF72ZNU2HXUjLx4RFnZJKU+DlqIlXmvK5+FPXsEg4k20CJ7CkjLCZBxIYlLLM
AxhDdeFpG/xdKuFWCuIfo381KPt0TBKQ4jEZEshfHp8hH/6Uhi/Yg361E3ru4Pky
2x6AWZWQ5stlug9RGys0bR98fLo/Ov4hZF0JONN3lQQHte5yzEmKvxbKsSsdKFk1
pAsEJAkZh8RPzgRfAgwL61yaNhmssTfI/o/vdYAzIA6joSDwR9eFreXP9BjZW7rX
MZ7vAE5ZHZmtw0Gb/ksGyDJ/JE/Xgeq/mUYGMWstqhtAXMddds1kxNtC/AtXStTm
FcsQCMIrtFkpxphUT64OawIYevGdXlsmcaNmj8VwSF4jUgZpMpT6nQSzx2UldO4r
2dwl3GMdcqxYJ9YO0Q3lqQDK37Y5rVRrXMn/eWSHeKfeJi3reziQdeD7utRSszYc
mWwSoznyMuneo8bIy57v1T+UUVR7ZkySzkd9pLUkvXYMvvs0zo4+saHW0xtrQjXw
/zmdYKqeujfKsdBeJ69aI3ygWEiexzPWX1ol+Op20jS9WrjBnXdUhVe8+Ih7vK50
Vn2txY3OIhNQZK/asPz8oNvQ9zpZ26a0sBd5+Bn9zb737KfkDD95AvyTOmNl8Uu/
4NXihpdiH86MN7ktnykts5K/BvvyaV9Lvg/lBA2cYLlU0942Z08r2GpfVcD9i5KA
nk37x/3M2yXH28nS7rBvWh/JMYusTFql2aZt3IXbb+PPuvkESdcis1k2X57jh7B8
+Ih9MNXUatB/aEWDM7KJNhNQ22aEzeHI3R2exWZTUxLdftwOS6ypHTHIJSWSOVNi
ACmYKja7LGkDq7ImF7S0ERNtDSkBIIEjAaZWwqRJ7a8aZ9hjtWUJBHoD2o9o7XCQ
CLVitJ85ncbV3QMrug1D/eLhu6xgI3EZKo/E7AXJOnim2FZQYhUrVL/71U8yGi2T
i31xo2GFqD2I2MQ3nAPmCyDMt87p/r5NAcfPbTkQBdWCjJEQbK0jHgq39rtYMwoT
Zm3ZVX+rMPP6RZftGRD7jAl32t8GDxy+mKtne+/pIMWJycAulZZxh5gFZlLfBiD1
mHFReCdh5VsJ6MVO2p+/zHzUR//0nW9Z+f52c5Hwx3Ou4vLS6XA7dqsn83AJcuYm
4aFaeSpcpQFtgy9sZDZgADOtVEr8i/Babj3enyU9T/SeCvtELV2CStiY+5xTbh1x
aUwXzeNrLB3ULWjkd6F2YX6NHoceMLI2+Rx6Lv8X9asUCO/n4wpAca3Xj8JbKBil
TanuHQsOq+IkmeCZTK3r8/zPzWQbgh/Jpt0TmY4j4cAdP96fnfEQYtMmMKbH7KUn
9ek9du7UBg8xq/QitXkiRmVXHaKPdgc9asDRlU50xVJLz22SnfExXIRHZmSZLcjG
SXCwYn8XSFXMiUyS+285pXD6wBjMKc3Rox8XuPcVCbBqD4Np8u8MOa48sBSY3MIF
MqHBobroXRLoJ/GBdbHKLgckyeyaWrazVMXdO0plPP25Da6u9zFgyHox53t5r0rE
PKeyfowXMBQLe9+ZglNOZBvZZ8tO3YX1S0NHkyQ+LRAaEu3fequ4fBFdHp9/rAeb
TQOcRAVKAXfDAvzErl0nGiM9ng6pDixM9ygxST94/3mHGzxZ/nqLNQ5QaYfkNf0+
FCVHFf00loKahW1Xx8llA75QDwobmW0RaL+Zsly6elzZwwsZSrc4jVB0RFkaGj9s
6ikf5s5+4x/6vcpLNxd5ISWhX27CGiB1ICfw0PnzNqq0oOqmvZna8a5kizTGHPoN
1zrQkcNwxKItVT6kshdgu6jw9r+o8UDeCB2/cNhSgVdAWVsnQv2etg8yeEt16wv3
0I6jlXgxd3f0yKBq76w+Wut5f3SKNMSsY6z9/IqIusPHs0wcLsUN8OxZ8n06MIfa
5mD7/AtRNlzgdko5QIfRrb35LDdE5s0/Nts/+RLmYRNnCVGqJn5dCJvUek9F7zUp
3Hst0oIUCls6dkiV9SieNP1kKy/d6FuWIusRAbKuGqjUp5IWRZQWlfMeHq3Sto/x
Yi1csgZ/mhkPQ39BBargbUlTrwqn1/l4q4b0K15bnY88Yx8ifoaU9Bj+NRwQQ8zB
TewmOkdIFcBwIkWLSOCdjBGKzJMzWEhHndztBcouSriMDFDMcwnerYvWRftlLRKM
mNwiRnDvcEZf2Pb2siAgcLLqUAkvDjIz5ly9Lcft6bFNHuJO9zT2xrqswl8yYXwT
DC2uDBirtrj2qDyBB2wrV47Oy2Mh82WiLKbyj45v/L9f+FidymNlf/9zrysC2jEI
KpS+HjhxfI8yAUt2XPbp2basPbBdLCY8vBl9ath/mWjzS1UTcZHIo3LVZwfXFDRD
4KS38R5FjkrNUZIVVjSHzck9bmlbkcjn5G4stiSwRpf3bgYzZMjQEoB0MZGNKqTa
Pq5k9LLiXc7k/KfG4QOe3hfAVRrNMeT4x9pNFJHJqOEnuJpMvUyiQZskNlLJxBsd
OdpXc3JHNCLDvv5ZBcfqA4uEQ2zQx8MRaerQ4UqgWDuVthN2uWGLefE3kYrIMIK5
qSbVk2V/xdMZnS+txZHotdy7c2NXhadx88AGMWkaoCnU06cxzsti6/5VAo96dFYP
Rxlw2Oove/ZggOHhzC4zmJnMdmke9KHrTx3KuJxSaz4O4BJztlbL/g+voxoScT0A
GLcU61bBnV3oyVu9yWuQkYXLqDiTQLqLfztbvlZkQpy/cH3LZ+aDyW1MlyDtKgAc
/h8T9LjPB8EirtaIZAYdtDSzPr1RKLY9wbAdY1ziAttRhwgnJ7tgySuDan3I9k5T
tLDcooBRg1tYLtWrhT1/M7cMnY5rPJGNjP1ZwUBg7+XhZHkV6t2E7/TFh51pIaJ2
uJkZIxzZo2wgMZ0Uik51bt5tEfpzaFmfrFlRpe3lM/9HHt6DFixfASR1dYA3dpaG
8/p+gd9nVEZsmf/B3qSIz4dlUD/pwsvED67Bxbw6Q+xyd6gU/gbl6mLlzN15dSbX
5jQr7aQP+sstikom3iuw2RHPBfyeTqkpNlVgDt8hGzOZkvcklSI7daHXrTzi/nu6
KtYx5MOQIrtUrrUQv2chqj6RT/Oja93XAgoI1Gn8TSoL166GpxTGQsHELeAsUU8M
sFL1XuwwLDWjwp59SIc/WraA3uhsKPRaU9H9Wv6A03OL3fI4/mFzB7/9Fg2M5jHH
zPz5pqA//GzuuDcTH3GU28sLr0Fd8G9xy4kuusskHSwJ6ScvzhzRdFTnEP0wgpxD
XbDV4pUjFww8/z2HpA4qpChfv+2snDGg4F33smc1qs5UHqn6tRVyqxtghv3zpJcS
jQU6oQ6UILRhsmtbKBlNcUFAg6IV5rbeoUfv/esei/DmX59mvEjRPSB6vZo8k0fN
FYl3DWKfcnzMMSE8wi0fnAu2E7ZrkNARg/P1TvDXYljCm277by68QMajAkik/6Mv
7CQAQmU54UFb1EUBlBacSZBD0N6bVs69HAG88NGd5f2A1qAA6DkUlKbm2Q7vBzd5
P6SrfKvfvwa+sjwSXc3jXBfoS8ZjEAcDVuTgOfbrKveQ+5CD4KJ3RlI9XnPM56J9
FU5/F5bs5/P5jrOGnGDb+sz//cYpVWtoQ/1zah1GIUZx2qPPkl+46vOx6xPTxHcg
3txXJrq5fLekVz4pB9d5LMyUta7J+ZrpEoMCgnh5XNXVjnFAr6lc0KZ6eWvtupEb
B6oOFqN2zIB59oI1haWkBAZpE/ZOfy5oyP5Bd4JntsgwVTWAeFk8Zy/9fpjE3E/g
YzU0ePyxFyw6UE7R3d36E8kr36NNcKcoiikF5y7GNo74pgZ2SzgKrX+sQoeTd9gv
+GUynQmhRZjcQ3Xw/gmozJ3x6lDmNEx08UmrqhzQqD/tgpuK8ixTQbk1JqXSvvYe
8jqDt5L+6tac7I2S4S3e3B2SZPr2gps28aC0o8tmXLa3ptHkpZdrybyNgKVsVLcc
ugnTiBSg2GH6Sy14XjP4josZFToq976J2mzaMH5vzMItpo8K5Da8fZL4NSDZcH1s
y2VXo+Ntsh5htZ20lAU5yvfkeBcW1pTAivP63rol2+jT3AW5ReIjlXpps5MFfutg
xNLDZc6iiBTI3U7zGnhQQ3R+sy2vfCg09Z3l9VKik0uCyp856/lZwqgfVpCm4WW8
TlVjUXBcthPjB4tx/95JCwxG5NfKha3v8ELvRRLivE7HeiTcaUO6yMB/4ehyE82z
IE9eDi/fn9NY3zJmWpZuYZiyYnxyf/ZaujXnn9lp8BbdCqIOdvkjze+uFlQebedu
M4dwBXYuL40z3+adOQF11kFGGginjrflqpPY4pwadCO7zDGap7RV/5yl6dL/MB8L
m1P/CGKZH6wppXAdx4ESqISv8dLHyeSrFqV7tqv3G+mKr4SFTa3oy5uRs4wWISmq
Ej6+hNZrPLMzlU8x1JMkH1wzJ2bTS1Q12kY4Q2gkQrrK8jVF6oz5ScMqdRtTwzUp
nNEG1psinxGQn1Jq9C4bOfMitRMzqHKNhNa8DAWDG3IqeL+UTmyu8t4rzhmKAKoI
6klgo4vVK/CbJdJB7WUcQzJS503Sxtl1IE71+JZJxUOa5dVai3Fx25rcx123pNo9
c831l4H7LHMPGwk0YEBOT/Fq6W5RBKetPwXZDC6ayWJCLSzKc/cLIkaOxP2JAsIc
2qdMV5Tr/Grp24H69jLiNopQ1LmTHVt3oa+AAN3sJxbGOW+fjLp0ncWb7y3kbTz8
7pO5RPnq0YRpCoYufnMlIIGK8jztahA6e4Cotx1/TJBYL7pEaoIxfmPOrHa7eVf0
mqUd7kg5SmQaV3jFzG1abgJP3q3/+58AmDeWFjsH/K25+10fC2Pjzv5T5ur7GLeL
nF2gd4JB/cTIHIrvhMkt/E1K2e0hNcIHlXaap6OZxS5fjPi/zAHITZHHj4bAkxWx
XEi/yJzsOmp5/i8lZ9QD8eRnCpBfxq/dy+iUpf9G+Gymc3P2Tq9tb+m/c/YvMmR9
z6YINPmNhVXKsPHb6kqpegki1hlIglWIvj28LX70VqDJvvJKb3k8045H7QtCR8BP
/LiArHF6aVX/GmgHx9rA6idoJkWor+xkXQQLWbd7TkoQouw+PT26ouZpOPGpZwLs
R8Wbvy0Q6EYoYf/2x0tgyyZKTR82V6/61JuaQxseQvxUUqSoIWweQ6DzXUIZDpuo
KXxGJh64+ox9IZnivg1eJQxgVUCx+7vs3Ma6DGhlJ7AL/XpfTsHlnAx9MdTKhFQW
2CZkRxJuZx8bkm4xNHFjoiqbBKRQkoKj1G0gC7zelqJyYsvyRpSeJYOmIPt0xdT8
iypS5UBllswfI+LUMIHiTHSoF7KLziBzYIOak2bQ/88WWw2Vunfj0rG0ZQX2av8Y
UVb27PHzUqKWm4pEQRMDQWOw8XzySZ4EqaP3/rUOT7EIWFB8BkJ/Y6EuA2a1GZ/f
OSv0hKHshYlTWmkMFPa0jnRMsKiGbss830n/SCdwutejDTRZVGKTGo2MONP/pMqi
4x15rKWxNE9SXZ/GzgeY7ZQjgfAnepmNGI0bloRkfiDi+MXuUDBdx5b8RFtu1RSx
TD2bsx1ZC6IS32LO+D+QYFZq6BCvubDGAGNVM9rVl9/Qgh+kODnrvAF9k8l4p39Z
D1FU9mx0G3Sr7Qcbf3cltK3480fKhcF5wCGyzq+bIUCF4z5lmPy0wpFNPq1zlfVE
rGvfE6mZSTsc3MHkD3Nq0hnGRFkc+61Ny5lcsLeckq76c+bC07QmqqbbLwgIGisv
fljKrfXYKM470wOw3fuqGDFTm4IEIuxJCDnkN+6khLxP4B0mVGslesII1Al6zd28
QGSwS5oBQMksV0VS0GU84lAqrXfpiXcAtsJVsf6tnUcT9TGnQ95Jhd1ijLPUeYcK
sZ+JJ/MaLW+JIUW7X6kE5d74tUQQb9zIM4d8tNWjeWsFLSPkcBnL24VqBcYWe+SX
ym5+SRByWA9j+tvfwKkjcKvXsLr+sDuHJz9L053SDbfoTYF0/GZdWpjsed36Zwr2
ZhRJCpyezx4Qv3AdIZz2HH2zO8Oy0YuMFEp1buJm/JveHIo+j5NCfsOtV+Iem/go
Bh8vXj6qrw+bXJILeLLeN6EjSDuzKhlUEO0BCO1Tsosux8rS2HbAX/S71gFTIUBx
gZir1QtaWrkQQpfSQ7kjNXB1RaC8V0YGA2R+k7QHiAMvtu2QhcOel4/PKSYzzL8d
HtRXxflvmUAa/vZ47m5SJVceUgdGEbSBADbxr/hB6BRHlhg+3hpufIz3AvDyY/U9
c/D06dhY1KfIzeOm56HuL0B2eqNunNwNJ7Hh01Ifob1jwsUgi56qX2VN0RbKR4t0
8deFgINMc9SnRu5vPTXVMsgaReCHlZxOCcU/Pxij2rRfkDGxIXV9Rbv7p4tZOYWk
dVOjaaPVrPihoij6qtJ1BZe5ADYAB8FGCjuaQLmuB8maad9pCST4KpTL5Gu8lt2E
ohgXR+0BviNRieyLP2Q4swt2/OHUPK8GSCvWB20NWOX9eeSE62WyMnXeaxB9usIn
lyP9RM/LmCarc+9RSvOL1In4/blRqUK1HDCZM6Q6sj9KgRq2TRH0HGRbiEwBuUos
vv/tOJ4HBw0w91Z98xwSgvEElhkHcW6ojcyI7cujX4I/iigw6MFFouNpMVrgypkk
nt4HEkZBXLnAchajsbQWV/2kod9m9v4i1T0BPCpM/D/wt4Uq4Js3HtjBOmNOpU5i
f8dRuhxrBsFeJixDJn1GTLJizcxhNbS/q0wIAofieqgGhzCqjFIgt4NFNUuFiLhb
40UfY4AdeJ9I71ZT6Us90Bv1jldnCsN1hD6VZK+KqaFdqxOghldo9yVbzKrTS/Dw
zSjlKuaNuCgA7Bjb4TyPf2K2H4ZB9Ty45gfXTiETQN66kqYgkqdzm5vehN/sm/eC
+EDnuMWj2KGvyD71XgZKscXD/YCYzlrc3tYD0OxcZ6K2PlmHO6sdRERbG6DaBFTB
EfHKUYLO+gJUinFgKtR4MNiWw68SMGTk/7kvlNkaep8mC63nVHO0heJcWIhiGhjV
hItcj0X8Oe5skpFiC3kWclrlm+QQK2KGXWsDt4kXBWOFLzyObYhsoLeg5PXMzdJn
HRJw+SVTeC+tELPvQBrex0WdklvRQ5DT41AZPBa702DzOqOwh5fzUaSVCFwFI2KB
7MdRpq19C4qNPZdVGqzXCNiZxwRfnZ9bR8sydsPTegVMGVJu5WHSs0XkSJLuRmsh
3tT8MM1imJAqbzog3j4TAKdmXA88y+ypBcm+4gpfuBnySI3hqN90IlQJ0uavTYrB
jX/769I1ym6UhzPLYLErK6EgiRU5clsfAtq6ETg9BAzZQtA9JYFX0Ok+jl6EQbNO
Mfr2qB+/CVkvwystjmJMI/NSrABVEibEfUJJUdm4zhxV71R+ORsiMcUyXFNIOuIy
V3rx0/+7EINiamUXDtpkg+nx1L7MRnyHMqRwqlb7BYmGjhJHApoQ1yrhkXKd2U6K
Z0pO649jR3yBTeqyO/7/xrym8VhwtK99pa+/Rv2DOtF6cI04qg3eoZEp72dUaXsG
2/I0xj948lM+szZXx4SNWBY/TNGbno2qj1ohJS+MZcBNdJ7reLuOOMLOm+sqPm1N
RWk2k57N3ndoi/njZsw0+3lZMoQAOrj2Nx0xTpYMLPAGI+wgyXoj55v4JU1no5qp
QLeUgzVIJxEMm9zbOg3jRMY71pH8ts2GmitIj4Pov6FFOZKVjmrY1mYAIWBW39P8
kKsSdQdsNyaHsiOFJDfBuyZypFMltcwIQHYoOfL+y+Ix8loMXAR0aF9R1pCu20Qk
b8VxEnUv/3k3QV9dtWpNoosqvNkBwn35havu3/ZBC7VeR8N+3ZEPlVdydsALrGpw
DhBJsgJNSX11Ij8MviWgy2mhCg1p2J/5/VO6d5p2uNN8kpSa06DHmPhB1XdTyues
QNvZ3y3ngf/uTmBtEwJMpA8uOlHpPeW0367qoGU+KPOBwZN6mPB5FeCowF4Dsrsu
eW14CxMwwrCVHPA+55uTi2Bne5d9g0NHTw3XsSHz8zM4btoE4QmkUV4TSNdiT3Y4
IfjvZ/+DoPgV7l9Fjez3vGR4DZWe4JwaZcLMfoB1pK0KBTfoPtfM9nub5usjQz2m
a/pVVebuCcmYsNT48diLAVUxgI9jQSuSc0JwPOxVXLP70LEJ/R6G0q0ZLmjpXE4e
V2O0Chd2FzIwBAEse02zU9sRC6c9Iule63/gPH5bg1mjUycNxCFaIkGu7ZucCw4F
bzOB4RY1mmy75fIBJpCxKxMTH2O/UW+KS0xY6M4e0bQAzDvcJb+pyA468SKo6+ED
U+9FoRnm8F2wAIEAKfPyhVzzFhbmJHAB7pLd5Nz0NE3xUfrj3H/FORUpbBApVG3W
XYXN1SLD1fB+JNtWudN2SxR6SZNd5evyDn6f8O5GaZ5ikPl+eukNnh+xCEWjSMp2
+9yPX2mLrvi/ZVQaFf29OrQ0tyN/CzVgqyMcf0x5JhiPf2TtERQpMc1YTfstJ92Y
2/Cn3i6GadPAtsPkxW0Abv2lvNgIdONOfIbQT5LxqH5e091E/cIoK88/RNlxCHCx
rwGGAPsVGkbYGbNO7dFHjifCeALa0xqIMO/XxpeMbVY9m9A4VMFpgrxfV/UKQPVS
aTdWBb0MD1JXKxNY7vXVdFfG7rqkOShzC7W0XhHLMNWK3MbraldcehZ4McNRqMZA
YgCmGk653XuMD2eNwouinfscN73Z+I8A8ckdUfbOzHUvdKALjyC6lfREsOehYRC0
QAlEPSEelkfD5S5fKkm3ezekxFOo4hDclm/wptrGYzWNO9+UT4KWejPwjecq11cB
iEujOpndlikpeVozH8e6cE+6vcw2KImM1dqJF99Z4Ot41GBkEAMOI+PSkxaX+amo
OTQ2lrzsIDkPXzvbeWy8XwbKU27NFuMoCxgZyuGNSPakSLftvvgMAEGpFHbrIywg
3/YYvhD8NeceazxJv58qnr6PnwrUHZqmWW3QkRkLpnUDRwPj8UWtalJuwdptbgmr
J3RgNpFHsOtXwtzYJDjdvONYYJ7983mLKB+l3bi+h1QAskOET/Dr3rjdgtuWUM62
DQa4YD+gKcie9rWPoaf9EOGq8qqxfOVQrH50vM6FjtcOs8tNc+1jbbVuVrFlW7xw
HDKKXryLShlP3000EJPjWLLRNybf87TmsSjZDxOWfUNof8P/cqKucM+p1NLxUORY
jPrOStm+ez7Ar1s6MZtw0V9NFwIa0svDlWaVrqTu/Dyle9nqSqPcdqJAGbgQSXh3
o1FF/c+lWTCSB/2/wfw11AwXEsYRl/zpu3Yl/xKoWeWMB+g91uF+DLx+Gze4QaI8
UWVPPm0UGpx76v+C76mmAKoRJKE+WoxFcdYYY7VvxDCgszKe5CfdyK3M7rLONIbl
0gxRHD575nltbfZQ5uwvq288ViayVcNQ5oPcBjJxktIi0wZbZrGgEm3eV9qy83aN
RHoN0UEZlRAiAdMPj4tW5oH4zrAmc7WdD9RBOlYbr26Haj1GqfgoHHzkQ+oZ2kdY
Wp4TC4In8dIHtzR/02pIprjRwLlHqSnZAiMyC18TF1Z0sKHWhbEJqnu3xRfnL0Dy
7zYttPy5T6IzH21RKMB0u/LhEB7sZaBHRb43C8oaIxqVgN5GKahUcE3Jpka1M6CK
vBrCglMNtLFKsKuAaNSvfdUQwlJiCgN9smWDasMP3qqkCxFJmuFZh5V2+g2R+olg
clduo+nmJgiTeFSzc5rLGz8E98beY3LwcqCPk+mk3c9mG3cIIMwJRoEITSuQ4PT2
yqd7rGIfA6OzEYaNhO9VJA2/2RMCzq8BqWC2UJITLZOE37RG5znfG4n2l+lDnJwe
EwimHzlCGsyRlm0u8qbyRHQSV35/VpHhfXgvJ3KGihZ6ktY0wYv+6MjWPjGvbp3f
9wS+caK6uk7XjJw8lCWlRryloIMfBGNaQF8427vyNO3InwoOWZ5rzDJIB0pxJOs8
kq9vN/9ixX6GU5b/C/znz4/BiUJQZ+ifPFv8OE73+iglpr6dbOK07GIo/sI6LbPl
q0OJRo/u/X5TSeA6Qld+Zk/LbaI7tM6SHkb5f48QIrEvZXXFuooqoEE5nIJH9Swn
VI+iNFW8J67rMgQGNuDuEpxKhTwI24+OzR7wPF6FnFTMCn9p2Lj2xZXXF0TXFgPO
kxwa7iVuIfxurRJWiSxxCseqHTQafEc8zmPNJnGWATz6iFx0wavkGJcSTfZJy3Y3
ZqCcZrNPNB5+9mTIVk5XrhA2iFL2JESSdcS5BltLYSwoGIuTmTCtiHDBSQN4wGJn
eYG2wCHlqmdRmS7fm5xlNnxvUyYc116oyfTecd4Trm4wSyHVfwGAcW9cBcEi8MDd
DXzLCtbhwWKPwrHFTRVBPU62J6L2JN7mgWOyhF0db3Hc0KTnJMyju/evH6jnRbXB
IGneB53jDmzIAU3OzriQIDNaqzPDaC8BrKz3ukHnRCQnX7tXkhx7uuVst+m+cdTc
6nBrF7g+S38jr3IlQP+ewV0OoM9IOeHBhaft0tnK1GMp5v9UnmWyjNcWdBqym81Z
AfqMhO4XDaT7HX8tfnYuhpKZK3zZ3JJEZyvct3ke1rmdwkaM6MTuXzJTebUGmVG6
3gzGSxv497jJMq1HJgDDS33XMBUOfCuWUcmhcORNBBeeF0nNvWLZqXkWP4XCmaqX
FeE8wUkOnrSw9spa+D9ZYoYpz/WUNUgkyuPdqH9eUgmh1uVH4NhDlZDs8wAwusEF
fvNQoFKAfzAjCI5a/dBdWgX8T8Y2jqg3PGVBZewU0TezsJEO8Q5mP/aiMIRvo8Eq
5dTu/R2ULqO4NuiIXLFpDP/6WNNBGImo/4enSy01sXfJx8HJJ02h9fbfgU0VwVMf
dtdbLyLYlNf8i7MfWZu71+NLCsrrCY0oiKOsya4IMo91WhvanPeNIIoOQ8ysa4XG
ROWlHhX2a43XbdHC1LIRLnhSdryl2KrqqhLNcPW3cSaB8zkafOLJcluwdYaNZUgv
3MjNFQNI6d/PBJ1R4AfCvRQk8n1SXFYQSBFUQjAyLhCsHHruvG/KyRbYXccYdf0P
Sg/gz2qqOJ6Unc7VOge61+7123tAGh4t7Y9BpOOlsuoQflhcDPAed2P5528zmLy7
JO8Gvh92oUzcbj55Voo4vKLVA3R+wxF1CCcRPND+JNRu9reFJU4VuI5aBKjmSHET
D6+skxlvNxtHmIGpmU3HxySqUZbJ+gAPXP4hdBdOyoN2vrsM7E4gfT8lY8bmtAFA
zfHDNlDwI5FztrYIM2wSCe1cyJeHwavYgYQ1lA8YldiCAhcWDN0kSi6Txqniisez
BG6xvuIGXKY02EtRhz7rjY64yMDluhbvPm7Pq8XgA8e0KpeFKPmgvkl1JehxjG5d
knQSE+Rx2f9VT79rss6GnkGqi8NEnKPcKtZfC3NPIFnY/dfZG/zpQjPgg6m1AmMz
xGAbdZphd3JyAqSnAJ4pwsjzJP+Ptwtm5JTyv+NfxYJVGL9mBoDCyeOhXM5KTDtd
EKFHhLWf3E1h2qcc6Ntc9kukwTDAfjh5fwjUvHuPx1JDXi4CbohpxZXGfdzMisq/
rmbSf6miPckhnKGIoLta6vExItQjvWUjddvgCxK7jL0Q/t6tu9771Sr4LJ7d8yIj
4tKQm7JRVa2DqdoXbiXFcsGW2pVUud9Y8P17aJpdl9iZMuk/qwaI+Yw9a3oHvqPo
lSDj+l7gx6sazo2VKuyxtKiPoQG1t5ief5fLOnpETO4oAcgMfM6yRx5lZ5NvCcid
O2bt3yYzaaW7tHrmHHavNTQtDvDt2EorKT6qS1EcKYKz1cKe+GQy4C0wwwIwjyUI
2mOEnNZlXIlAHEa88ld8oXRLLoVFk/pefsFOvpXDhzJt4mkxQWpRBC+AqzN8HZBP
77e9HjGj94os+YPz0eN+NljInxjDbfloshvU6l84IBvk6vz3g7lmFiiL3dO3pdTn
2nV17B7jhqD3jL9GsxLa1yjwNk8ruc0T58Mp8jXAP5UW8+mUp43ddfWkRvgeW4V2
i8U1QCpDeN9tWiGdejJeyUEwrYZaVvsNrUWa7gQZlGwXLzxFj+1PKPVofxDdvEYU
H+O1IJTKZWCTw+Uk3q8FZ/xEFEzSmbinF6l5Hli8tl8WDqGZiFTQH2o8rcZqExyt
QWN/k934fDW1KKwYEuUP3ubBQk8sqLv4Lw8XqqDirQUJgwgpoGK/iD9muIX69aoJ
xzHo6/46iL/VCIlLLuZtBEhJMANvhWxp9eeRfAwP0TH9jZOCaqCVpS+W5WnDWLoJ
W7SOZRzsSqo7PWb4524Tgjb4xZj71ltU8amvPT4A0X+Kf7NkGtnwUYFg1oN3NzuS
qVu9oqAxXCkZLMF3aFy0jAFHh/y++jw+ubmlqzFg/dgnyHjSfZ3Yuc2Wzdv8oFZU
X33QZBbUbRTndleTBBfnEAUOWJ6evgIpR0JUvIiY4xXqSXtUz7PMbiWXOtnJUzWV
3AJPhde630WqIuyCFyA1K2O+nXDuWlIm89fRfXmZgPf0xHxJfhr7DSiuWmlj9UyH
4xEtvD+j7E5dWSaS7GtWjl8D6/xCVvBZP2Z7DQUBmkn+kG1e/VsY1IMgvK875UTc
mOeTOvV1qcKWCzwN5E6p2OcjYeVfMsc5NyZvcuBaEBAsqVw/A9QD4MzIXqWzM/Vo
clrOSswTCRUXwLmMsyzNqEiAABGEY0GZHB97eI+jAYNfxuiOIX6dCWIeXRaM7azZ
4E6Ic31q7Gl3auA1ZSWy6QTPnjteeEB8xyswRWE83AmGUsIUYtfJLp4IxnIb2bMb
1m+uS9jw1M7CN9lGqgaYaY2r8hZr+aChlee4QXH5hGnP8vyoCrJeTTd7805QWCIy
hFMxOQz89hf3hHYp3y7+ANMI02et7XyCfAkxFbTdDb+WI4A2tBmRzrC7qav5O/+c
f2e7filiw8Sk/iKKcHxz2NErmTXBALjkcHnO3vlejMyPXiS92pcJBU+B3YnqZo//
b3N85sBrpwPJmbwyozw2hv0XWjovWf87CsAPaqBb3R64TjkPlutLpREuE9avsYVT
NO2GFXjCBUXxGHrxf7ytaINBiIWOHqoXNatlvAZySEJjNoCTkR5WK0kCxQhUlgFY
RxzKNLnUVy0Rsoecgo7bRfmTbejR/qmdN4wMx/n2vL3d8GlMPWuy6cC2PVofymrr
LMmYWXZpR5KEti753/yGQJ3UpEOnJMgeDgqcopLv9ThRrx8cyWnpoNQ2EFqVzhag
4bEKJk4k3JTRHOZkUZ6fDF/YKGX/5U1sTVEKqrwhki7FXdqWAaZCQCPEh7oFBVpI
QEpODlYvKotxRZjKxVQ0PA4JtpNeoDyKw++r0SEf92GnG+dTuQlmBnobq0u5M7ZD
qVjqJhtlxPbshjJC3B6Ecgd9hzdNABrhrsTz9wNoRklR+N+1BR8b2uI1hYp7wmA3
TAIbbyfj3U1oOtK6ViLoQQmNLn21smrjjK9e1pSVcbv01X7hPSwI0XpQp5BSefAY
rXsQsnkkjhog0/VXTDVfCgyIqwgji4dy4H35nwwZLAEc8p86WO4QxcLBmzQKLEYn
+yu4I/bNn1KS80uRgNC6hO3QLtRKfH79gM5JXwze/W59CC3cEgc1yVTeZyM7Qcwd
48l8F7AlRBqdECNuFzXT67rAW1ng9pKhdnDThdOcyJJ4Yiv7FErLfnMt4f5iMAR/
s5BXpI/bIOCZ1Jjbybn/k8hRX75zcL9XIxlURtxoiNGkXqbdFud8fvk0Bn7TZIOc
uFSdqgbJEDWp9VzujhjNRevQujRlz24R7p6WLvvTGHHwTWyr3U/ENj1mYoJ6Ogyk
1ulias4tFHhtkvR7r1kjBtxDLWnKY/h/LIbGmTVW4VSyRplTpnnoCCCZY0crmrAK
3A6zI6kSFcy4kkgybxbbeR2PNjI1cd6bhMUEloYsO01OmocNSTyCYiYWBUdcl3Y6
Cfw5iS9Zji44XI+zHzl2oi9fCMk6bFeE5xn0sCOv1guj6hZBHqBe4rQdQVmcHOG8
4uk7NaPe26vYTGatqai2Dk/ppFDkj1QXI1CEonX0o1xLf7cD4NObKnv1TO6ejKAz
tbq+8NayfW7WnEY5zWG3+gklFr7Us0zR7LJXxyTEGfqV7jKA/ebrxV7n68SP+eBu
d5i68Dcptmlu8Jkq7ETuRChPNlSvl/I6HU/ZMeyiofcSPK/MSadwJdDVJpgzqnz9
GZ7Za5MbqT7Mi0JPa3F1E/a2Z53MDFCjXTYLWj3vCNALWN6g90C4IM2440iZIPHd
kVwnyuBcuJQaRPtkKHde1I1bW3CqgHMwZVfgJ5G3wCpH3herHK1iZ3njmxLx6dZQ
VK287HJoW6TCk1cP5liPoQ5INsSFSrQQjfji8InNbcQpduuaw/4tGFu1EOd0Z9DW
X8OhLbug1aA7wvImjQ0sY6e6xVxvOBlEp+EhvI51uLK1NV5SJWGRvdlJM2Tf5Att
4Xji18FcNKwg6KNwQQXTtwMBSnzBB4ugHIqS5P/WSKQxTMpPsFeI/tVLoUBnXzdV
aFnSIgKYEp4qFreP7Pw7bBs3Y6ydPl2/zCZ7JYEoprpIQL1kBbG7Ha/uhW9vEo7Y
rY7Kcj7NIZAa9ndeshbTAtwgOSr0qZQNVIS6+ICxdGwLmC2m7XBl5psMpLH8mE1z
SYoc5M91v9VVQFYStcDjupFa60T3i0NSxY/o1Rc6MuVwBWDk1EHbvGu9s3JsI0qB
txDulQk6g3ijvTcZUzK0MrVJC5GeJS7izz5SWH26LSjZ9arajlLcDmLgftXdB4t2
jBx6F5iJezF2to+UEqX5GmTLDkkkPn5bTGrH3BNIxQ1Kcebf4HR/3FI8yYkn9zxH
3ryCXIQTiF4y4905ha44JI+5NXO7XiH/h9u4XQo5naYYfVj0KW/2wTwNOQF9B/8a
NW+w2J0NbBtwa3ONSmIH8DqagozqKSvGUBY7guiBeOCYHHhFnG+9wTHmxVAIIKHG
mbLiPZyNoeXYUAPUrLxc/XfzhRQoA0R1ZPwh+HnYMTGFexUOP+YT8bZkXoDdnVNU
TRlfJ+nHElZsdbUQVo/aXrmp56am7T56lN3wMGiTzzNUnYZfopB0rZOa9iSK+AHt
SsHMQFpoIezC0v4EZKDVUgq2lxN1PGwv0dTc2Ohy6WCvpz1TIUIANnDBjwq31rgz
+rYKToF5cvBHgNMXN2CfwkAM/lMz8Xd/R0eNI0xWshCdVdPoFo4rbdLD+7Z0nJNH
Llus8XmdPdiHjDCdWhUHPEJRh6dLBW+hmMJJrn0hA7+DFzSPh7WdK7svdQVLlyWn
aL+hS+4ibAAgoEsvl5rcOovE4iC67jYS3srTptg6B3rBSTfzIh9JRA6xPxvtq6rt
XbiRVbjgS6m0C3/95r0oeZv0kl2EmJCt3sbvQHFuHpgSTQoN/6BH8vvUdFCRFdKF
44uK29DBaZWoStSkAKwtD7L96xQO8Xw71uWJcdlIXoImwxmPIR9KloWOeZbgv2Xw
+sf49HWYuhBecoLRMTIKmcN1D/yncenMH3v526T1Lj3ZbOh4couMhQZvNSmIOpJ1
yeHsXWpolITJy1Fl/RhHxyM83+rEtbMNss3etLdEZzcfbGi5kOMEGbJ3SA3JdnSc
8FSh18cY0L7yLyEhdv+bLrzwrTNbSneHXHDoS1+o/cichzHoYdN8TT1ZbUkf0Ehh
sGVbhfHyhoBBg5nJBxUvCmDcAJGnyM+Unfkp+qe787JShTRjJ8dZNGJPSNUQrDw+
mrJ/iSD6qC9oBkbSpDY47gAN5gcTBs4Y2RJI1Rt4XZItmCgcFbenkNowq+UfHdy4
wRonC5ziJxnAAZX98E9HDV/W5JHKrn6tV2ymUTojambGPA+9IgW2LHy+LFZuCMi/
6w3Yl4b+HqQjFgqP1g79dIrdpZDooPtLZaDrYQdVCY6rC7vJX0KcPwYKZTiOUuns
pse402SUguosJEgUyAI4OF/3TFo+liiwiyR1prFENcOV+fD65t6AV7eJYWXoLekL
ZM31B7Q0dhX0891ilroiTLnkWnzSFsxPj0Xy38wVUJOl9TagkKmaMXal7ylzpeaQ
5A6i0q18b84wDNlV7/FsT5BF20EUtTg+akMx7kI+eiu/GTXPzRP3kV7K+iCoOZ3E
MOA/X26hbHIhtp+Kj6cYPeXqbVViWuDSxfUgtmbBdJxILv0tj6DeoZW67RZEZOP+
Sjh2f7yQ67Si901v3pVgsQDDaAe2PVVHozyI6a+5zlwuFqBD7WC+HmA/+Z8FE2WG
AdXrlJo1OAvT1MFnb2VuhFrH93Jm+NImu6J0MYl0NE1TtMRlxLueOXUXu4OJB1wl
F8+Q4hY1vg5z+qtbPBW2QUH51/ct0ZIAXCFu1O1DgPjVjZJk6uo79B/FiwzOcroY
H5FvpxwGS9jk0NmgtlMgaLS/0Wqa0UWWUqmaREyzRU5IpafulUXU1y4JhWuFRbAc
SgnDAFS4oWjSxwHDBJQU/K2N4I3lm26X3b6zqE+QXCHje4jpRPUMOoC0GLVwXWPe
EBy9hzdLsIJdbY2sxVZIJ3dh3EoVJCcB8e9ymEaDo5KyYDRew9hdu2XXwsKTJB5l
jIsqzz5KXrlA/bmkG1fBpW/7+sRVwNcaTNHqoTDjlRrf/A3bp9wyxXowRWp+JnK0
Ga1/Q9Y/ybFrvwwfPmcU9EhbvAvnGfRJaosHMhpq4rqxJMY4z1gqXsybQxV66mqx
QURPB8VoalPXR/YXts6/ut7yPpbkNwbhpN+f+Ckk/Jc04beHWSqGcd0zcc037ILM
0rSroJAGZHdO+nDQBPbUxpFW5pYduznJg7NbnYHg+f0IMODS3Ud3jlHupUBpWXEb
d2l/X7UjxFfEpA03OZLayePXG4LslLwfFfHhnPlBI/56fgAD88i3vpsfoXR6DRXN
fktd3AffFlw2XB9uaUMZrqgnxF6WUVHEWa9Sbjx/bK6UEqLifYljN/8oMcjZRHsz
rn7NdiDJIknFYF9PUNHLtks4Xr6FlezkvrurwLLzLGvnHz2CU7gOC7enpROm7YGh
odWlK/1GOKL+YWm+jgdro+2y0w76zhJqy2jQNYnwYPsfJheak7fMzI9wQHuHfBYq
SIJCo3QUcC4KHGXIqWuXjvUgKhL7xqDN8kEkaTK3RA+hCezvjrWlg5kiVjC0spBp
ubYPQ5HAGxQsJZiggpVzrnahmDBYRylxEcQSOxW+NjWnDGS0XLvqV7bZp16OS1uu
q6isrDSTZXcUeToLxzX8nA1IuaVyv8Bfdjgji8Fwxa7GO1StpE0r5OdKPRff2kxQ
AzmcMidEE7753KmWo0yRtGnbC7usSvb54yRU9xezINWGD4xtSdeQCBNlQCMh8wzc
o2snst7yWIyJPwZo/g13OrM7vPx3imNiVwhvJ90I/OvH+sUj0IoQ3hFo0NxBw7rl
N009Ed+nIgVtfBSwRj4oGOIImE99zzx/yJ2yHmSC33HHaHXHFbRf9FZqUFpQ0TuS
FIZQ0jY4qagnIPKJWId0NldZY7pJHa5+6NC08Mk1Ocfaqj0UWkTZv1Eq1hVm+g3g
UdcbjdVEk457NWmlFZtM+DCPiceRW5BMVvCIg46pfGLOVIPzYTrRCVz0w/oHY5KA
kE99nw5iiYjAR26JTO4yKP6VnJsffGkgHFyR1faZTbCQZH/UA79yl++ALPAmU+rJ
xSk8ojXg28GJTo7JUBuPZbKZQKjhr+j7YN1e+7NhqSHwxuFiLbxpQ2bJccYwojMY
DUmhEFQP97v0k+j+Vj1ZqqVbTWzrla6jD34p3PTlD3eJW1I/3BvcVvWQbGiaKaBg
Ew77CnnpP9sb9sufg2eo92sjrGQ8cpi3LZKTN7l43Tlb0Aoczpqv1n1uvExV51X/
3yb3Egd+rRyI1lV1do7ltdHqw/vcqjNcAtONmQi10C2EZJC9mmpNxNq4uvLX4iWz
K3ctDD49mUPboy8go2fC6/IABu3gqfzAmRjMDOWraNZ0eyj0zu760oNlOYEf3b6m
blMQV8QVgsl1hQqTcZVNty3ToAVeqxUkiyjfk6gAHY8ihgMQZ6+Ul/cw5MCjLMSF
a4uw8Z6eB5m/wqu8677MDNcEaog1ibZVkuaML28GQULPQLYwulcIWjcgqQ5jXpqu
g3xSkThR89M+6Vf+ejPY2ATY8ifXZO4tJtvxkcLo4pAvTepsTTkdNSdqyqqpSbB6
D/TUZI31o28Axs8/Lii1/ccegXDPKYBR5qj6ZON4pbQ9TufwoGjgBK2Og72eDGew
uCwOku26ZqylFL7DaHbKWexxig0SKsZYEW8ItFpCwZSx8cMZIz5qjYe8Rwq/dHwH
5pm4mJVIDKkddQGhzH259THSuEaD0XJ/NU25KFwYKXkcapmYGvqOFXhaIjYheG/0
j3yKsb+Va+S1cHOrTb4e3dThr4F49Lmle54XljAP947GY78y093h7OXj2TZ4fdWO
13MeW1s9Xl0dpRBmVdewZKJY0JXuT8DH22e42kSGSiHMnD/rOZZiPVjpuGiFWzIm
SOZ9bgYgel3rG168AJqx68fXWOAfGTiczWzHbv/jeB0eE5FgSURTWh0wPFNLb6WZ
jlsVixGCbTJeBq3htyk/UTzBlJx1lAx+JOQQpdImhEbW5IZXgpXY2GOW2BlU1YC3
GHjdytkE+NJv9vZ5hO9t62mFOsjnQV7VRPDHjRgZa2boO+vkr4ozScgihCtKmluu
XOCE8npnvs8TxtG+be/KVNSYkXVFeKlkvd038gTk2VLx07F2cMdvTkUz/zRnfsQm
QvwtNsqXxJi5MGxne+ViQvK9XEyULzPFcvOYyg4rcm/AjpdzkecgbNt8JlFHhGhl
eysJC4QpwHSDGhhOU98TFvNKPAJH1RlhxpJSCQvl9CzGA1ZC92E2Auukb5FZDqHK
Dc1MwCudXP50D60ig8GtrYJY7OTdZ8Euszd1nBtAV0wv+CKCZ0ECB0Mcs3ZXGp52
2cCwxqMdvkmBwobA3cuaXgG1eed6lyYIlomRtMup203GT8aRSMk2kFVjNwrIuOn9
hhc74fkpixmoVC1VMbc44Cn4mnRWalXHPO1Kfry1Elbx13Ub+aMiUh/7rtg77FxK
RoAeC0J2FQzXF49YCPjBT8ygxnRb7EmwOPZ5oQadHGSkACKtjE4GH5Hkud/Xr3wb
uexIxA8WNY5l8smHf13cIxVmEqGF5SwJsu8jV86an8oCRSi7KPjpZL3OJ/KfkEf/
fyL7GYfX/W548fsIaQZnIyVeu8U4WoCmC8K0jmY6AWiVJp6neHsECq7v+xzy22Ml
/R+cY4HnHxpSkjnS/vroGG4512BEajGT9UbuBbQcgQ1PO+4R/314E9oiC1re9nfD
K4Bp7jamg+DhPsIJ8b4z6KISXZ2Ufaaz0BJFk7CZnDkwYfH0VRXmsTI+EWQjPuvG
jWcHEjDxx5PucY6xrwNAGfXFr1pbZzq3NrOkWhbLB6uStPywqKCjpNJWxJ5iI+WC
4/+khgitPsC+ol5AloBHMDvQND2opBdi7qBqW6x0MUPAT8aaHCdsc3/MJ1MGYlTW
dUHCBkan3AmgAECXI2k9f7LN/xBvX9y600mFjGzVURd8vR8VNdFfsE0rZHla87lW
uHxXXfkK6hpX33JmVJI1Bbz1yTdYDKQEwtsGeCWxKg/Z2X0xxfqg90eRurw5x1q4
0kZQ3usQARupGRM19yaFi592dWToblsZGyUhXGT6EkkjLV+/1iw5yoiXbBG18LbA
mUnjBULWmyeG2AHefdiiR7G4KDUx30gb2Nix+e66f3lFIRGVUfvWx/eQJ/DOdYzq
XF2a4XvkWj8x1sEv3jBOG8xbWV8/9kAIgFXJqhdkQrAs1acFiyIXKUUo/HisNmdc
FL3MyluMeJc54XCFq4jWt3iLXaholz6NnUVGv1bQFCFYJb3W0R/1JP3OF9+/4ymn
Cu07CmUtkmrB6DlLNrQnKMlVwuIlaHTA2c4cYpgJ1BbqQlEbT373ALcXEyYvV+2l
7DBV9rcQipKj5X+tz+A8ck+vqcNL4G23HtE/xegcPBxMVomPi11BL3M0nEWDiDUI
f7n5E4mcJFZz+maCQ6UqNzS6jH/ZPDX+fCj3gKKe9m7l/5c5XQ3+T1y7t85nDs1d
k34IeoEXKtfE1LZ2qZ4C/uZTmcw/MfAH2opsxF+Z9Qs3rTUIWIBsUFJWKivVq90c
lIfKYg4e/OjdeTFUt6+vzu7KAb8SXg5d6DUuczKbwrDlXbef7z8y6Udgf9X9200I
NsfX0Pm1f25K7k0OZ5JWlp8Yq/X4k0CHJ+M+2KykoE421xtDnvcUGj9jsQAOgKyK
8YN1fBBrykcNBcifZafepCkM/fWPsJBK3k6u/p3Irag8kFTU3e37/lh4h98B2trw
/NniNGvYAfOKPYrW4Dn2ToS94cXWMmgUCqmmzCSI4XzpAsg6fnrAO0Q2JJGG7hlH
uXe3BqnsljbjP/I3GesBSdcl6bHo++ZvEm7ddHtDROqzgeylIoAJAEWPnChxFl3F
ivppJF8VlL/2yUdZv0I2A4ZJB4A2vLNoAaMbN2scgbo1qE2MynMEYV7XqrNkzAcw
jwPVBCSlEO7vPkiaDY+Y9JaHnTfefWHW8rIF0o8VY/+sJp8+zGexd4/Z1XY4SBkz
qbfxRGnvAm+KyrJ56KuqQXiafCpAH4rgva64iUITXZZUfub6Y1tA6MIDdBPuKPga
eq+n2xMIGdKawwfHhQjQeEA15k7N1VTOeiwRTjnvVhpLE/nyeryb9PO9RJZ5WizC
G+WzATeF27OKg1cT/h/bsdRhB8vZgMCow7aTMwxuQbCG1QXRDswr7AMZcmptb2Dc
PivtTnTpOLq1uGzFiqQtWKvZMO/zzfUG9mrtNDje6V9oQqSPAcjzrXk3c9m9nJnn
Hidxz5GvrTXcGxUzsh1rln2JbceyfsWIELVFWsg4aHZmoRs/17P+ingt3d//DXVE
hpSwJYFPP+bK1tlcQx4HMLU7H27dJozctSKz7oaH9PPAvct/PjPBT5jyYkxCphnC
oKWy/k8Lt7dSsxN15keUIJ97mRxIfsi2sZCO00uaHim2Zl816xkH2htMc9NT4GoJ
SGOKBiDLj8n14F9rnW+87xLN+vRSH2/XZ0TAIoS2/qwW5s7MXwdnLCrUisiJ/7N2
Zj6tgTsLU1JLo8/WUf91CefERQQcTB+TLvdCTI/ldwxoofCTh2U1jeCaWgbIsyt2
UwpKMPCeU/s5cugccYt3gZk1cDKiMmNqrt7BRUysn3exa7lhbZ7/Bybx5o/WCsFt
7Ixwe8ZwDvYnyqL1yla2XmkERzLudiORZ9itLU9t5iiHIE7AYbJQUhjW5XgUy1D6
xP+B7gCsuphfWxCISejNBCjAVGjK936wL1Uvfrb697/iNoo1APbbfX8di8IZm2PM
Qr2VTlFcOXjYVKfPuCL5vVeyuY2NUU+WpN+fhOPm9iAy6CHmOcEaRfm6sfsVfsYI
UXPThB3C/HaTkn2sXRLyWouCwJcxnMEFtxYIPsSU5B3O3uYgPbz5+yxAR2FcZc+p
YQ7jxoE9vGGDkTaOrvYkmFcuTmpC7fgbLnyM/vFi3EFTwD8j1JAhhFM7l3PjsCkn
Q0w/Gt9nhEexWOzcyw80RU+BmbpNkOJMlkSRpL/JTmhdskupQa0Lfd/9c04jzl3i
cC6eD+Tyzpfafi/SVdx1TfPBOh8365lRO9r3DqbOE4/eH00/SAXjyG2p1Ag6OWib
ncjlYurbrQvjn/u6i3MkYCbNi1pBoKTiKqGwwXw3TRwYBcrxMep17U0Yo+cgb2sZ
sEXY1qDp0AppxGQS7X8ViokXrr09lvBEA5pAu2a5h1yRqZ/XH++Hl5/wXLrzN//h
cIyLdrgif/jbSVp9yXfJTciGPjLkhC7IkET7MJItbritb4BGTG+Z5bhCvxTh6UVx
4T3lr5QENkeCUDgzmB8a9LX80/hrisN4HzrLtwutF2pTUqdrkjRsqlC5PXkehXJj
Z2vnbqdtXBJnu2oI58ndraufe/aooDgAsJ0IrINSAmYVkfUcJxNNvUTs6jxvK0Xi
ChctiXzuytKc/lF81d6UxAjWSsL35gcHOalIgez/U/S4QFZ1F3+i0MIk+X7jlU6N
DC8OjG0d8dTtMFE8Zq8jV/b+rsv0VV1ZG6iRUgQPITzkT0MtNKeH7sq7OuPPjJLi
BOG3JnfDKtv4Cgdiy0QFIywMq9hxrz91vdoGRtvZeOEu/dz/wWt1ifjvIn3w9Wlm
HqD2PYGBk2KZ55Q/CCe8HqMDRoBDZsIzxU8AUPVa0cXX0GBKhmAT29MfSJTN0NX3
LM2hjDsHb+N0MBXW0g6gQBtgfS3Qtk7iAaJBfof21kehVaqgRWILR3OCVcN+qpnW
ctv37kaAhuDg6+HbNlccVjdFBfDws0NyBi7xbwjuaCjuZvlfcQ9GicK9wanZ6Rkj
HKjyVIzZBye9Cao0EJFCZ+sTrldxubQCLYNMsftUXto7cyrTrhqtvDrUKFLM1SC1
eXHXOqMIUHyQeb5xEZn6K+HuwEwKtjia8hHNir0N3uCoMnEVQ5r8ZgqcIgInUNNi
uwiLg629MQB7ZSxmCx9/zBVDK7OUXx6yzIhfhoO7M4TeBdGBtbGvc+yMN8MEqhNA
uORYJooLJzjcAVzbOo/UpjsB3b7rMuCa4IuFrllz+imHHDYek5UPCKIt+mIXqHUd
QRTzltBNQ/Om2/w5M6CeOLLXJ2tosFSFMs9uEzcaOmKgbcBWTpPpygXCJufAAaLu
x+VADgk7KS2l99WL16GfZkqsjjnRMsX1FVncxd/h3bSJhtRLE4E15rsxE5vMJeSO
JFGZgqhNhpVDzLlvZs9vxzKBqv4GO538X7OgdcXkmWwzmRK0ja7XMQkUQGycGeBv
gCYYLi07h+CNShU9k9/XGhudWVU13G7GCQrz/GgBLGZ2Is2vHlNJmKevJ7sFmMNI
OcycYi3UlC/yR9zUdUtWZb12noJl7B5N5sk+x8E02T8Vz5+g0EN+B6wAk1lCkFLY
JFtQwprilJbgvt6QunGDqwUQSY+npTAH+B5wlZ1fu+5Fa6qkdllN/WN9Rg9fA9Gy
OeYnP+y4ZdMl6NRVi+UN59KP1pYLCz00mbYx+7l4PZgQnWigTID2x5qJtCf8c61o
VV7P+ZKhbc45SGtqmbDb2xhkdzc77KIOAguVWLBdcGkkbDjHwWxzTLtApsyMYl7r
SU15TDkxHEQ75Q5k/+RTvgROTnXaOA3yGEac9WOamiSW860/qpQFkTU2vMp1NBAB
CHGDDahlCLswT5Pv/tpPX0txakLi7o2Gi7EWyYzA+xRl29w1qAyVwKNTB437tlFJ
3jO+wXx4I4Xx4pC2YGdlAoGjW85WOLeBgiT94E2pW45ZE7uarWVJmV+Sc+rsDJtQ
ZjmeSFtkQAxkQjSMmav/62/qrG2btDaMNz3Rlr8Q/fA86/Du3Ysl2Bl74VgghFhg
ho2bQ6H14qPnXkxo7NhJTwZkaojJNCTDwtWdU/zTZmS0AeDc5jRuBtmDSksz8pmn
Gn6YYdscApuUVYmBd0qKn5pdX3LoLiPvwKvfolc6zFgoteVOu2WCJbpKqd5zum4S
OyzwUw+3t2lRFwhXjBKzAqG6ZMEP2OvVraxMTAJ8ydqnBWlbj+XH72QYJzQShjJd
b7CcxRMm75T3y8M+yfzuJf3PLI55O5zkCyz9wgAeKlnTktEumKqWkCGamqYRPxDG
4sf2wecUCk/PLwm461wEL2SvsWdDK0NuJIeXRo7Xr1i79he1COXPNy7z5IMQ2+hi
8qBVaaTsYAAj8Dv8xRo9c9GuE8/gZ1U5QhD/NFOE/NnLIdS4vpPsWfnth9GXXYJ3
jzWI1AETPzH/OmbS/FIlYO9ZZJhSzwafOLgPf2jzgvAi3e41Wu2wvL2VPqE+ZyP4
pU0mySypI0KvWVs+l2yK0RwJLJFs394yaVzf6VGHTz1F38583fXrN7Pja9Iy7CU2
8+qhM+rfKmrqVnsxqd5KR4PpSe72bnRE8zmvvJmf73dbu/N43wiaMdgKpyHLQhwH
SDtGEO+9FVNczWN+WthvliqreuCozbELXUbE50D2UnVBWmKAxnvPpaygPMAC5WOx
nCi8cAnaWdtwyo5azfIcF5PhIYfJN2pY68eF1RdB3A6WOXrzIBr2k3ELU1VuxTvl
5SmHE0HoXrtr7S7oww+xeqXwpbjNhyrqZAtzPxecjh8EUM1JSkRrwng5TupCPQ0e
FfPLMcrUzCgJ1VINmBMBVJdlKUnHSjHp5Eq0dEUYeCRWuSh6c33Agj44ds8LFpqC
8ERAcivGx5xeth1IQ/jWRRSiz3FTfETB17S21/DDm2uO6fw8NF8Nr5KSFpbIV9t3
3leo2Y93C6znv9Sdo6qygzyUB1V1a2qENC2Avz9FnvQmRZQpPJ+Eu5dmMrFpdjcK
80Hi+xY7KwWMQ01u9kpS55Ykrv2zjZpzPmFonRFTMyTxFJfPlYd5K6ShaSEQ+xNG
IMZ8CPPn3bs7N9XV7VQg0llN35Kkt38DQM2X2hhYVjsRWD+KaTT+xlARZVLdJsdx
g7wSRuaApHKzlWCZKcPwBMGsk39cFAKjkxlAPH1mJOP2EOQU5kMsaaVLwINPB/ro
/WQ5XqBXIDsbuB/C3D1KAuGQ5w7kp+LMRW7VVDbb1IC77NZ/ft2QQlt9Y+RqLjrr
+cvn03eYEpGJ0KZEUHmLALDnDJTOUbf2rn5eRENVQcrLKptnn36k6o8+Mugiffgc
C65s2BiM1iO1p1fohI01MpPA7NYkz+D1jZFOM7yyQ/TpGGFejQNOSS8syPlP51uJ
StQqFA4GXY5xWo1ch8QitbDRlYgwc2BIZxT37CEkP+seRGun2L3jeaVCr24NRHdn
yM7WTCxfGfncOafcvzYXXeBUQtyEZNVqiS3YwMoA6fEGNE5vPzGpEwZboQ0CXIi7
omyTSQfbzrP13ItKVhMxpz9ck+uIPmT+fPOLRzbMBcD/vJ1GBo5bGe4ruIROxzBL
M6dGwP8WLRkbZB7lft/zZRjS5RsclDgr2qT8yHzO3nQiZbWAbZJSoZro3QSMuk8a
fGIkunF7IswBEMdsnwxukzAx6gun+91pXSd6s9CdoY/qwbmGoOgzfN4c0WP0qvTl
8+bylGC6SfY/5/pxzxHgUc80OoxsxWoLd+zDLKy/kFl8+7Fs0a0Hbt3yVMfP42M9
J8uZwqnIgxgsxizPW/mUaCZSHbEy3sMObBh8MAzxe3voFgPFJCGfa0ZUD9QBHVPv
Px7F+m5uyR50DYI+wEu8nNitGGA5Vw+Yp5/VNVgb7zypgF9HGCP3vIV0khBhixjQ
62Qi+JmxzIpnyUBlSnPxfis7W2vo4DcwDTa/IQSfXNV2j/9WLk+I1hVW0GhDz/WF
CKEWt5NCSZYbOszB734PChlSAuuzZBBXT5JK3UKoOS0cpi1YRJOYfPcwNYP7QIdG
/K3wPACAsuvT5NMq4T+Pc8W9EfxvWd7PXZvf202ycKhJ2d35m4ZOA0LG2kwXxDxm
+inYbqLuD7qugOoFBHksuXwqjs5gz79Hrj93tuCYH5JefTuATkj4ZTspMt6ALQJC
m7IAyZF520zBjw6+DcXDgQ1NVqQ4g1dm1mGqGmF/DIAmbv6L8eFMYmp5R/H8+Dly
7mpNMJN3WTNhIVzhO5yZqNKy1/qmPp1LStreSvngaHRF/Y2Rqu4RKL8GE+lv9R+0
xbBODvN3QCH0fiJkGaGckOHI+iHs4VI1uG6ebeZD4t8JyD9BdWww3wy1Abbci4p9
K7B3fwdbTZYq7esTpUNggWwdtZoDXnLC0+h/C2gJEV/XVw9id8D5sfOkDy9+5a9b
N7vVuyRzpYv7IcHywZNw2H58LBFtzcwN4WGzYWeqLIYUBFJ/6H8gfTTaELddb8lV
XmqwvB78RJ2nt9WYn7K/4QA4VQQGXcyA1DmDeRq/Kfuh9+TVyN4J8RULmoFVDxzD
kHEhSkawHrghvWMC6p9w3bfEPwmjJyN47GL6hyypX7z3h4Mi/so60fabdPOcH47a
LqySZJdyWnRII0d9R6QmZos5a+bKVYTr8OdQtYAGkKRYvIV2CC+0g3TaPCcnD88C
Hi9XGmRjHKcebsRL8pX78NwkYIS9/mCaw9Nro04aeM0cDEpGGiqP6I4nrcFjkS9d
WyW82Z53KNZG0aP64pE/Yf/nu6Mks0zCIcPQzkjXR1W8Z7sjPL8l47CmX/DGLyDp
gfZWhpRjJUd3FoEtFftdJQASfBfLTLBbPjynRSlP8sWVg+EdWiGIAXoQq8GbO6du
ku6ESLrWLET6lUaedDb210PrxDFC/QIsSNa4SYCErhQo+GQClcNZV4asO/hCvKQA
5BHsviK7BGupNjCY2d9x3MajxobkS21Vj0kO2b53QIIfvtFutz3FzadbQ4NMH3um
cvrQq4xZFR4YfgUc2Yim5kjbrWVHtQHzKSNMDu+DborG4t22RcjxSJBN1mfLRNE6
M8NuTqIT8SewYJ9+BrF3lI6WOMYlGB4mR9IrBmECTHsFEfZBqoaCa7qmpDm920PC
hNuZaYjp738uAOBFclE0j8mDcd/GdIF/PdktxCHRMGlW/ECJ6gjDdr3kN8MKFWua
l80i3bZHU+e7V8mGyyBfV9Y6cWqdnQwXqvA/Q6d2b9i7wmI50Ok1SbS6VsEkfBd6
1iNAexsxVyzdpqvZdgkg0dMvu0byMnqX2ggyDa3ixG05GzqwxRRrWc/OOYMm/1wE
Ns0IVyLbxnS1NrZIry7T+y+sRiQVOSSL9PxbbXsQ3qmBWcOxaFG7QP08/QZg4sBe
CJKEFD1PPetisotc2W7ZjRcpR6l0Gkck4fw3aiJ3rB/3krtBLmDm9Prn3eenGkV3
+4qE2CmVJ7R8+WnXd8Fo6s6GNt48bjopxgZ37ki33dhhQAYuLb3mCzaHtvO6COsN
c7iqvq2CQYD63AC+mT/QRzrHVjG2iGfkao6gl80UkkWfLV6Gke9pnbEMEjpVVQ/q
eWagEnVVLIDXYZQmmgmtSParNU8ZcahTx7Cfz4u3NYjamwKg0N6d8oZHHjrZoQkn
hyi+bWLCuxr+g+uoKrpEK1/5XTumOuGqb3b4N/+0goojMpVqDjLHKQG/whLzX+Sg
NFAfHZMhRL4y+VQOZTh9VAFLO794Ht+jJ9QmfhqlFQLcon3IojsPXq+NVmf8a7rH
hDfZDBVjFEDCJOqN4bklSdUSuFochukpQCMRm0L0+f27zceSRMc7TtiEtAic/5Fs
fUNUgor2oiJRmGFGZTVGkkC6m5jN1sIrFIo1rVOfmCypTb8WOMCwxo3+QyCZ6Qfv
15K8UR3w0zawN4EhZWPzYNaN9o4x3yUaOP3t/EEf1sF4gK8ft7xTg/yhM3TA6Y9D
I/hgWba/SSb1XB0bYv1DU1gOEyXKk/rLzT937Jd/+zYcsH4cttARC4IGo4M6YjeS
eghD73xRNffRYPnRhFDt9HonKPiHCg36dr4iMg2JIOpfjDvduYPAg3LFHH8XIc9v
c1rKCcVN8Vpf+QDgcRXYmCJfJKC4Zef34WwJCdjwB+JiJ0P8buRidOu5JrKR9Y0R
fIcHP3NQ87e5JspkIIZr/R2TKP57NhC2gkNBTw/zdnCQakBLZ61FgDQ1nlxVeBA5
iwWhrvqBkQ7UY1cSyIpa13V8uNdo8rooIPH5eI2mzeBzTEaV4vWncYm34M7IgCHA
mRN8OSENnJW6Tumw9ZMkN/aT/35L+w1YRqMR3+oJxTfR7M66O5fwAx15RqfYWPdC
ufTpsUqNMGZzR7yy7q3fbl83x0oCImexrtWCUAYeN8p3NntLGD17mVsoILIY6H4G
QwouwHdJND2ctlqDu5nNIOf+0no9s9dLVPPXV0aZiAV/qXsMwqXBayRaXd/jcZ2m
kPUgFZ8F3tu39La1dsZNH7kPYsT9nnzwLXGoiVeR+483JitmiNkmMM39C66zbkQP
0QweSgKa9VeE0L+DER2GjQxy0pPyJXjB3JjlU4nJ2zvj/l3mgg3cRgg0t1hsJkXG
lJLfVUl/kXLYWAAJOae6VSUuC/Z3M6jVXHo3jlVGVQZV7EJ/sx4D//b8Cduq17t7
WE7rgKK2T2c3h7oe3vcIEGBfJ86/B1vqbXlsrrr7+cUC1H5lr+nsgnMKulHF63Lh
dzAiBa7IEvbOJbFchQx0uXatkDZ2QUbD/wABLMOu4E2OokjdqNb8of4jfjSJPMbF
F79zU/KByMksE8IfnLnaFMrzOOeYFsJhTSnP3r952IXSZBeSsMcw2YnZg8HZeCVF
RPOKakvmRIDQ0Dk/ikdCL2sZGO+ypJiCvjDYItK2lMLIIPJeZrTUPRWBrsGPDVrd
fim8iy3h/MgjG8uv9iXe6rXiaYkpr2xBoVUBktPtJ06A3LnbL1jwreMgUmEugvfB
pvgKHCPx68JBkX/nLUxgVQy2PHa1iqNdvDDQb0SVXgf0BdMBHSblapZMvY1xiAih
VQ8pYrz4X3Rk/wUn3wEA50G3hE/Oc6vFQKwshpj3pO7zy2F0BOiao8B4QmUT24Ah
VmkXllG6Hbb2EWk2uSS9H91dD4RIornX0KHc+6SfjS5egP6BBEQ7VJyQGBTPBd0b
TP3awSUCQOSLuv6MlQVP4hhW8aFO48HyZ0Hb4XRv9i+Canh0dARD/fc4MGvLgJiq
1sb8f839qRJIUwIjhHkC4sDsWclP2UVqw8I1OaAgO8aO3ke1/wSE7C4PYHnyom/c
DYYmbZZenxG+lx4eEZhW+rho5BThCmSP4eSsV5kttMk126YqD0TWfVF/FkiN5vi1
Et92SY4QzR6cqwXE+2h+OVlYreAiysSXQ+820nLgjZAR4IlFMbGCKSZnZv8es9em
Zhql4O7t5BcxQc6o41pbGC2ypxfLeulud2oRCBBR7Cqv4t/ghaYxaJy/pb0APqwK
0n0U3ugq7EXScnLe9tf/q9LFGH+QpzXN3yVC5moX0GlqqrOL1rk01AkDJVrdRvQN
wB/qZ8OvkvFRrRnOx2tDidGcugyiRmXI8l+B8wjcTxUbCy+ObcFcs9UBYCW0YOTM
Snad2DhA2dam8sRIgYBdVejrvYpFG6g8XeiFxuPZu/wuRW/d72yIGiTdzpn4rLJc
oe2sM7m2zk8jWipldbe9hyatq9h6reQmxdymJsrgqYg2DCbkxbB+8LhSqiJNCLsP
UyMgBBSjYyfDi+KMxDKhtnxT+jOLO7zpKGvSyhG77/lQFndcHYkqoyl8gUyoD/MO
jnyzdGGc0Ndm64UE19C8EzQ1QMVxccu2QNVagpz6fAiNguA5JLU9xsw/VB9DZ1cA
Th53z8y0cMIQWVAf5cYBMueVTkpPRTON+LwFpkQgG9AE6mBNkfu8j0cH/lHVTAyf
zl3oOatlMKrgZpy8oQ+S+V64cpDzvLVr7Gkd+Mxa6gUYP2Je3GVFOQgEu74ZTxv9
dMTNuvXwk4PMw5Tg22cCUtKqvnZYpg7zIQP9IZOvE/xb11sOUWFE39N0wwuM+h5K
1+zALglnbOxY0OtDqZkcycp55FlExJaIwQljpEjKXPQwyVfKfZsLzOl6CMCy7D3V
AdQUGJY+H0nPKl0rg1e7WWhKU+gPQKDKAWwv+9FE160Mmacdik+aHkR+iSd6t1Kc
APfPEOeUA32MmzvaJtMVREGDaElh6chmxe9TF1ackVcbY0yRr8S7Zr5+L0j3a3FH
piom6WLM3CcCQ08YmAINaf1Cl0l6qh7OTfldoNbmCGfZzVAj73WQ1iHam1RG9x+A
fcPzyexN7BFTM3G3GTu34wxlBzJFu17aaxiWvtpkjvINUhsVaP9osLV7CGCSkERI
DF56sKAFxYXuFZQrs7IlZdXXnyxjn368GJPj47fJvPYhzLFqV/8svlaYeFTTHta0
N/mAW3BRuW0zFOVkPPh3aE17OfSWC/KZyEsYogIlwhiXSvZMHa4C9CAgpSlgHudF
lXVozuLGUqv7X+9IPkdDGheYE+LPlKxbFe21dAtmlI4tDdZ2UnEnlxqfAR5zQi92
TIIY218e6jxM5bYi2TstJ9anrO91Cjqw8h3V7ysq6Y3V/S6syoaVTKZ26Rus0cCs
DdEhP9P5NisX1UxezH23aapnMmbE01TBLQdSA6PxrMK/TJAt6fKgiXJhJRxZJQx7
mOwgFflkqrAG9EF/9R/Y4oc+dYlj95GH1Tp1fSUkExB/ZC8KDUnN5iBsM21W9gYr
ezkC6W5dbEzLSxaF26weHNSOWik5R//xyVV8+AnRiII7fhcprpKPLYhAxjbsDT1H
RpQPfx+TU90sfKMm5YbHLwHWVHb6tRuxmcW1SI21nFOxAf43B+YcM9ZF7TPXioe8
+snobIrQQSbQXkJ6lcfO2V3pCLK5b6EmfLpIxEbcmqScO31FOvqXjVkhotQYmCLg
5ODm8kSZg0GdM72E64FHuEmJOh2PFV4ybVp2Wjm2yNeAp7V+LD0a+JmIqMI6WOJE
pnVGpXC6XTlI6XqbpsB7GxWBkJ8rgCPqhAMaaJwjDnqdRVcKZ0ueZ/ZYXHGBmGGg
HkU962VB6OmLfYWxnxh320wZT7mie3Dw7DePv9db367/fJ6oo8vtUVqDtBpBZvyD
ImdVt9o1B1wtQqzdnECD6LBWQ8C2kPoIxhdRT/U9KAKUxHcfYazCOp8/DRekfLkV
5gCd7m0MF5HJ8g6Qs4Zs97pGfhJnSyO8+3peMecTqfEVx3OHl0ACrPuCTbhzUKK4
ynncGj7TNuvZztOxkJ1QT+x1V3FklvYoz2geQCAyVblnGPdtQaX/KcYZIurj8kCV
4jIBFozg8B6gcGap+FZA9XATMd2B6cErZtF1TDahwhTxDozVnvYOT6zBWCIBVwaF
oklTFq4e6dDTz02wyB4ldAG4w8tvXDqrZVKZa+vwo+24zmRdSKxYd3WnlW4IPzXM
d6YX8UA7eV4v/rm/6Y0RsbdqYN6cjcRD90/DFQtGleC4j6n1rS2O7V+krh1QAKON
JgEzMo59RyWpRHKxj5lwa1Ghb9lHQB1aiL2TflRkXJzuQ0OBj63IrGMIz3OJfxIh
DCcjNqJ7NmQX5YKCgVsXfqAGkVOuaRzt2s8mw++qjPgjLzF3CfEN9hmM6duT9s5c
N46dam1zASgqw++6bI68WNWZm64UDlrQQ3BWXmBs2RWXEnChzr3tDK0EH13aZb6V
ECLaGLeSXccBvpkHtbcP/lMokZJzR+vBHTZogS+q1vz/AfCkUiW/5pXeKG3zR1Ri
7UyWCR69PLI2NVYnV57/MmKslKKIp+XjERfXYOEhDMuRkYmrk4xgAWM4xs/ah3ET
kpaZi/zKsSR9GSXD73aQlKGzs9oYNwGLHMxU0PjP2NpmZ+ir02R6E2qxquGJhjK3
Vi+HMJAvxnORAqkJ4myn7SuWp7hzm7hC2UzsbPVB3CzX/UmpVFwUW+xiWA5j71F5
vZOXyzuP78RIrqQvE9UI7uBISIhz8GqVuckF9Z0XpTDR6v4dlFXqz9tOhQVGEexF
/l6FtfxkLnOTJETDtlBm7QC1nS9PozUNiVKV718ip6MnCgYgK/wZM3WA6QhN+HCg
sFqB6F9k32XzlA6M3h6k8r+sMnEhLxaGGL569IYTQF6OMhlVSWfxFNoYTtMzxsKT
gbEINeRhISxYeCLuU3sjhc3qnDbJ9RA32jM4zQmZJk5LQfCJeFyUJf52MwHg7iSR
+Xxwu+ePBWcf2YGP2BRNQlhFViZ+S5pgydocfIjCKj10KkUXGwu+0yro/5gzJFWa
SjOrPn5jQFzWajifAYtg1XFM/1N8Cj2oI2RfPDyhgiq6NH2gAyr762fZ1MP9gE31
UiOx2BSOiU0QpymLNaKY05MdFtRJQHq00tln3OzJLqa/Ls7L7Qoq8Rfj0s8TZkbm
Tj/X+Kx52lLHOai5wkreMRfBJBHwHqe2/3TsXhPcmiQgdtVHxtXD0cP0k+mACFWh
3KCA2CsMF2qUd3/Spiekm1YjOq8OHLaCQww/ggEuktMQPi5jGmpcNk5NNkWgPS9M
WGtLVFmI1+5+FOFCitAjfJoVNlcEsWExcQ8y3R0NOFHks4ufXVR4elKzyR8MYxjO
rJm6Ku8gaMdKl7+sjmYdvGcZBx9f+h0mQXkC2OmlB1sCKoekHDfdvzHKwsIRyyn/
5ag9uaIQmd5gtnq+fsbdMbfTlPCL8jMnsGfbUVCVLS605jk72vCISzh+SEOHEx4p
hUP5xlnW9iDy3ty0oWBDRyfq708iR23sh9DafWoOmUP5IvioOoPbXMfxkEQqQzvc
8bF0IW494S/Mw47AGqtOME0cq+afNsiUtfa1q6X1lZlXlBWAkqnAQ5ScZPdLIfJ9
gGM7Yk7d0bLI2mU7/EDqrrIchbAZar8TvUdAJmblOAPLSebfY+8uqfYjtF5ZkyCG
a+b6CAAwsDMv5B3bozsFfmTz2pNGn01QA46ukfXt/3d+N4ZoK3i30gS+ClHxdEDW
DrKtU+1fs0H9IFH5cvUSF7CPrBWQEC8NzLjmgBywHsaS9WcazKq43xcsq7XDvyfP
iKjP/RfiPKgPXcw7mDMPp6lu/mUtmvobpiDfhSL20H/ZPGnRV7LHGUakAnaAkt64
nyKieoXJv4baccvXGc/AVy5j9xjR6o+RmwunKYM6yk0BypxSQz6QmC2sFP3I9ZLA
gwgc1I/oJf/TpM882OvXUWJtZ0ZY8qOyYKjDw7rIlA7j2oauYKSIkjiktQoVufLM
sMyzPYjCdg7xDaSnOeTJUs3R9AQiYQPyqQaxIio394RKu/ztdSfpGcLGB+CAaiFV
bXpLlVm4HdeJKHyhRaItCG4oJEa0kKBIyeRkmEyf9fK2m+fCvoWCRhrBei3XBbxN
D7UIr6yKFcfui67sje5Xf4BoXCel8HilIN+JLRvMpMmuJEtu5AD5F6oCnhqZ07U0
IejVnrXW6Zz4nLJdM3lNwWd9LZesdA0o8RWAA+f193ZjorHcWlwNnkm2Bbtulazv
hdlaIUbujhWqCxltroUhfQEc1g8zbwGC9fL4tdnlVd9dnzfCXUgKgw8uCBtwIrN+
L9zjfhHksJY37HtzHvXJgNXG3+a2et/E2YAekM7MwI0jc7Vx7PZrsXqwVMV2jrDD
u0zmYLqcjR7SP+8VslYD6esyG639HuliTsdFx37cX98E3I/Zgb2Z0kq6tcz2JeRN
H7iSnJuR0kl5ydxhIgJonNQp/5+iI77eH8cxOZp034iyj81sr493Gohu2+gLV+LU
Wln5gaQU0yvZ2lzv75PddBjHZ7qbYEn8DDyodDz5tKJ4zX8Y1Fnx84rm3qdkCJRK
jFpMvwjLaOfKn2bpsu4Ri8EOEFCsyJ8lUWOPh36Mv+wLV98Ur2NY6ACQ3rMniW0u
D8hJKaaj72pDMsi2Hc9ugwOWbW9Q5E1Hb5muVYlJ25tcePLhViem/7KXpfI6B3Ij
SuzEEWjzvx5V6SoQyt+2fFd9BIublLKIV6ap4FLllatWE/wmOA1rK5vCjJgsoOx4
PFpNFLBVR1XEf8+C6+MPLgIKQ4XhC0/kkJ3/1HGnAAT8dhw2Lti1mv/zUn1ZfjrW
mGWV/4PSVaOTuR6Qk13FEbG1BMwGwdDyDVgkG7uh44JTMxfqmuOMXNJbZNachnZf
IF0NxUzaXF9PHSpK6gV7HgphaMrWr36BiRmMkQfjCZfeJ+Z2A26XCXzoqMNXqoEF
C7W4D5qdwJaJjCOQj5guLClbwZphZ9rrIjklgXOm35nlCkk40wMWvrLyv+LYurQN
8GAuUJQbNdFb55G/HyeGoF7fkT/OHNMj+u4ui8NwjRiv2DnE9DKD/eLhlm+xKDVF
GnIZOSQ4f3JkHJCFNI/8fLERQ3QsrDswziv/JI7kZu71iarJRaiimacXuwB2BP1w
RcF1HmUzcwuzeEACDEucbQkVDMpkjs8+d0NC2yXRvwIbunYpzYibT8IrOU0hqqDP
1KTQ7EFnwrVjpgiCN2Be7UO3a6md2JZMInK+W5710dbr+CR867PvCC6CCh+hv0Yw
cexSUOmkLy2Fe365sZNxeaclC7SNJmITFphkjilkbuZ4ohuH0KXYnbP8WTuelMI6
YRkB7B/zcfoFe5Xkz+yvlvaRPtKWt7S0fzb2rxRBUmgAp29qZfdhS7L43IFF+Qcd
oCDEHy2axthRA5Aj3i1xwbhuY9f04vkeUk9IQLEEv0bANqLuHrzjqbZBgfq5rBXI
7duqH/sXSse3g1dHyEon4IMvetkDVIFrRJslyV7guh2O4vacGUt+28DgRpQZF2MF
IMQUgCEIKOrX7VXtkpXlMuxcaGv5q45JF1WHEscmCrfGaeA0K1WtEczTaMHFEree
XAUqfdpc2HUTfAObhzdCtX3maX68a8XVNhRWSgVByxn0qKD5Aq8zIqpD4NkAScP1
rjedZoMd7Q/uInclfadVL21tBOsxtxv6mOLUc5j1KciVV6uJ6wODiISXj/9FQo+S
6FbHhW5tF8glDjUVGWB0MQBs6LKjJ19z1Auaif0NUCZaUyKR3OtYn9LRKaS3BnYN
mmt1CMT6+PRgbQg3HWgVi6iqeGeqFTO/5wI6v/kkpummWt27BBIL+63CfqIrYDOw
I8t97n+9jXbphrsBBiXqXuuFWpB50XzWbhmh38Huk5xrUZQBkiPB8zjDug+1+YWb
TO0Ugv1kj3TfYRD4Fxt5zHpDJyvVgpMuTNa4wyTaAi73MZAY4+lZhATy4Rl7lgLI
epuojP/4boPLF7RkwsQKFn4pDhBHD1YHOslm4INedLxUBk015JJkGVZza6VvRt78
FwjLqOZe/MJ3u2vn5kiA41a/gg6NAkLATnsp6eNKVMe/LoOn4CrXhGyLoY4Fm0RR
FkZ2FOn3wEvWuMOPeYiHF7XJQN2r9QqeTq9E1XPZ1AEoeHgBjdIWs09Zwy4DP/dD
Spw4lefvkRIzYS8L3Gyfmhkmd6xfVGLKZJwKUTNaaCrmgEx/MjS32zbSLKXPFcRX
40I3suOvCmds4OWiA3qibRxn3rxvzvWvhQMMbqGrtdJKlN3ADIl1dU1K2D0rHry+
WuW+v+sllrwL1AMaSIXnm0vlKDoT5cZOZCQNedYTweuYe2p2k+kGMFWKXx+kNNT9
JB1cSTHTblRBCGRcgO0/Hbss0tzqVP5mlINy/FMvu0Iqe8Qa0HW21Hi2OXY1pZEs
2wyFv59rrJC2Ek32oCigdsSHwFVgz1WsqMJ7sHo4q2IkYKUou4RDQefq0mPpHiBq
sHymRQ0vgHFjDg3pKTEog5IJ+NoPt03pxBn0aYKWYsq2ZUJ2jA9Aezc7FhfPR1VJ
ZD922EQR7Djm5mZdi1lGyVZuOXHoyCYbSyJwxeu9ziR55c9eTNonsq1ww3HC8HLd
66Gki2MetqHT9LMn4Yr128Xxtsi1+0PqpTGloKBhQ7aWekZ4S4j6Sfny/nKnJeaK
0EgX6t5Z9RMeTKHa2MoYfB9tYV43yhm4BZfLBH/lG9LLYwNCvN/OdeAUuD2NEjyc
3Gst0d3px+DKvq/ohR8V8GwbgsOXEWjQKvngZWpZAnBaymv+tgQFWaPnxRqWfdsU
9u0ZJOGaJJ8fAoyezd0tG+p+WNpZ532y1vRM9S/H9m/2MArq38hyTOHCQt4XxXgI
lqL/NLt4+/ublSgYtC/wkpoC+rAyRsIZhax/fFi5/WZiKb/Ff2L2LDpm7QUQ9xvA
2J9lwOAUuHzCJSJNab3x+L2OKrYL3RQCNh02EA+vq4uabAgsqsAlKEOOncgTgzrb
Fkm8O09i130ptSYqCccaL1USghVVu619dmoiM8+R0Zh868fEyML3C+HD/VdeI6go
L5tCmP8zQvc5HtlwxEdF1NZ07/poFKBg/HYgjfnGLU42YPi/uhDXqPItXrkXgj1w
cqiu6tCEr1KrZL9hJdyJzcJoPj2KWC7rLSRkHZFYukD29L11IAK9hD5zsFbu1e5Y
6EDKPuig7ykT0d0m0sFFzR5dHVmhntFpXsxc/4nMhPVvPk8gCOrDitLkX7KQ5MEZ
F79nGiQUrmmu7s87BeHFcS/woy6XjXGOjRugDiNsq70ckduxz3me7YlThXIphH1S
qNgMQEGBREbjAvz587ZQyCuJAWhLnXjOiC/lnEROQ4fGCyc1nJihtn9UQviKErKU
WawPlVK7Qp6o9yMBpHiRJzberAphHSORy4Z8Pa2goYO0C4VqfMhxXT8h78gveqDX
8GyOiRB70QY90vDRTykNLAI9A3RmByIWntIj/i2bs/l8/oGuzsFGWKVpkN5bjSfy
rcU++k/xVw+Gr4FC74p76uxAemisiPQ0Nc5EGaYb5NXk9mi1oEYMr2FQjmBcAwiR
vieiQCV2ZjzGnd9qCgFRL4RJU9kINWWxgoUhruhSk/PewCHSDj/29tJp6xq/l7kA
Uc87/vuhg4+6zlidWru4tDaOXeylJXHTCPcLWZqrX0r8o702Z/av+rYMqTiFcEai
KuJkBHyH3LH9I2SU+32ZnK6V+Sg2HEsgz7tyxynLaiQPurlmL5yRGzfRDI/SADtV
MsPkaie9xIb/2T+fWfnab6Gtx1Awz7HhNKHarnumYf1Z/1bBBTUpDeVMc0RnOu40
DUxcMhSfdOTcrFWRM/mdaOuqM5RDJn1sQSMeapGn5+syHd8KhVQOg9ot8NI6ZRjc
+ZnyuxNZxG2ClV3ApspL6r2HwuyD+u094ydFxO9HpCAZAQa+YSkSe9sxySnpCJg1
NGoNPYEK229mKmxn8UPdaofetGXfBuQJ1CUqUeJ3hvXq0+BozoGpHl7wewLMHdgE
IHea70acLfZFkEugpVO9ES37VCOACiX2CeaBnnQZsqJpunetn89ChXTBbCVFI9aa
ES1h+OzrVWfQFQ8OmOgiYp5Kw8gCDN4VihDBBYrmYBI4qzyiXbt7e1xlcdydyCLK
11E1VvkGpZM3pfZvfS3tT3x+6WTCgbHMsItS4t/vJtl1dERWifU2gF+ttOqhHCkX
NxeCPFCwBvZqi43qaJfbOoW/Kn2ls54Xhp4rJspZhgBWaysfFz73CUSDAl58u4+b
g//JPF2UC+8G5jApGPH5/+guVJHvFZaYgbb1rdkf0NPO88D1GElgdlfso6PLewjx
5ylvFWLYzbnycG9vTey79i10npaYa0yUi5nnS0QExucEXsSwcsbV45PU5PwVANTA
Gw+U8haQ1GjTHeYNkBQ2T/0T5QLxz0brIzVebdNTBSxkq5q4hcjbr75mjUAtQHTi
1bp9I0TOPZw9Gp8GXgdY6Tzubik3DA6INd3mqDi0wqObYuvMNTSlkUeT+JOOnb6d
YWM0wc5mZUFoBAlzqmrvGGfdRcLP6tQ5X/+JRjZNhw0UD8oD3ZdTHvUWWmCXHVEx
G1Dr73VAU92T5pjg+HQowC1C+K/yIDPKHSXKyWh+RW92cEcRWT56UK9oU9kinDud
j4V8+8ZROok1V5WLU3fdiT0Zahgg0VsWJuKmgZS9PyfZwCmQO/plFT0aNr31vVK1
oz/w1490kIkzgDQ78zAXhQ42sg8UawbdSq+LGphNqkTsfOeB4va/FzfGULKNKvAp
MmEqggoEx3U2Uo72lhRwzS9oTFhUwkjJaxdtIlpvBt49WeC9uuqBfWouWMCVuLyw
X5mSCv7AqayN22dNfYSw21Ril2Iozkk39AGIWY/IgRiLgKCy60qL/o7Mpj92UEjI
GBqH4x10RAjoop7odVGTaf4OAnZbIP6siLaWHEAJs8GWG5H8bQFT0X2IB3yjOmj/
M/tIkkUk8mTXfkrSuf98Qbn/fKTMYmpkGNSA5y72IFjsiCB/x2iBwkMpUpT50Phj
iG2tHdY+zgQLxn1WAI/RGvsemhgqXAF9sUEv4gpREamaEhpTdX9ckgxRD21zZirI
EaZ9QVedYd0/OaR2C88s+jELi7iEwBs9E1Xjt/1RYcgdPyP4s/cnCUTwuwpnKbmG
SBViFZ/hXXf8PmQT6DQriY3YX59oSK2QFmANco8dsEEHMZvfP+6XRq2Z/g8nbq4k
ZcHO4cVC5S7rCJdBlquhdZnUxhZrdVD5L7b8lKO4tYxBIopmhMUwNh1qTwNoYVgP
/PWEii4hcT0cwjJLPi4NInCb71u4Hs7Y0K4l5j7jXyEdAMDLEdd+dY2uU7iwDwJU
fiflnwpGRL3WDuL4EjfDhK7Y35FHHSUka/ACQzNqXIqouBh0y8xC8y1zFcFUPOq5
6JXr4q+JQ3TTRumAr0YrJnsjGz+y1pBRMiAOV03sbWTacmAQGRFnHmRlRGUYZCpE
yd5Jhf9kbHiMo5qWtfSAGx+hCSchA84aeRnjR3W3d5DLp5aUfGxE6jBxZW7gXLRs
LdpIYr5S7saPQl+9yS6eTq3omYHaAB+PUwc9GxVfRFAI433MOv9GTKusFd+387n+
3xT/n070goo4NW2aezE/L18gakA4+wcaETRnPm9NL+G5XMa6CKPBIZQdzKm/qIFK
+PW/qeMy74XVFlgdNPKlZsbaIDrs4mUH/mBQA3Xv4K3eHCDCTOfocl38HN0SVtaK
cyFffXLVn4RiuonenstZqurupWugzUC4la42yQiNNKAb1hS+VBoyOZcSX+6NpiU7
cdGxeHqbt4inPOzszh6LHJMnTjTZCuLpGrxbhaM8CXBJ8Cie5xuEn5xM1sffYten
wvbEnY7j8aoPQWh8D5a2w1Gni/Dm5H0X4Cnh8NATBK+eCtj0njTyP/AIjdl816p8
6RXyY9ucotB0gOO8sGlYjVezXEbPfMf3zPP9eOlQPC/YAnhInP9wH88Q1mPq4OW2
d+6tKohYbNB1M1Tn1WVvwIkxq+eLGygTr533d/mSjZO8566AuTCrXrP7O2+8Ygto
5x29q4TL+GUInhUshByRKmrUJAmEVd3DTyTR8xDzDc+iQUxSGWQqQnfHdXkfU+xS
G+oMGFFCRqos5IqRqVuWNywRGZ/VJCXvGp2FUGS9RoKmhip7o8mvqjoLmIOmpsku
bAnvfdDV/iJ5rOgT+vRYwWUgBLf6ufpU8vweAbFbf06y7lSbRoAodBCYGR/dTEy/
8NcUP9hfkSCszJLxkDsSeHAg11Bc9XQoM5SQNflJQxIfDjrHus7I2VuyyzWDqU3D
wWZM2OLPEdDNMFuwEvZaMR69s0NuzaSsQt9VKumV1euq1ZovT16Y2ajUxVd4VUH3
7qCybFl1G6FjejCP1k2RTT56OL2yLl4DMKy0j62T8FhvKgIN8GkpCIUzCsf5fiaZ
HZe9Ms4DGmIDnWDAzQlITBpXBnW2E8wA0VJbCBCyRVwoUIAoh5JoDNHb7GyYJ+SW
9xjohWhAfoYnYlPImayaCoTkh0LVVdWLSXF2e6TmAKbxsbiiQ/hd2WCS0t4VKM+a
CfObWXzKs+g9EiZV1msbMKHeHCbhePaN8IgzdFoLseceQQ6LoYZ4HDcyFeDficzs
pIeGeRvXJgt3CfnjxoaNQNUkUoi1aw5IND4vPu2k5tCSnvWfu7ib7O3NgGMzY2b2
zIAOxagtYzyMe3dTio1K7Pl73z0Tm5KyKhaQdRjSCU3kAMoz0G0+fE4RVUISYrpd
J2Okldgo3VVNX+l1ODh4VdjSYqZxaMgq1bcojS6e2DXeDuDbewVKeS5Cf1MF3y7a
M7jBXNv/quoU/fRkC2eRWRcnMIyOlHfGxcMBgQV3304UVwOMjzWq2dAqWZIHf1h/
rcrWAtP6IB8tiwH+FWAqiaWctljpNRwvbg7ExQSohw9wPvb/zph5p7AUPFwFY9xX
4iBT/C1K0wrEkQcr72mpk1M3M2V5Lz6obAr+IooJ/VbuMyypjVkM0gct3Sn5EdBc
1FtNHQWt/Qusa8HGt+bX1yNmz1DQ7g9NS+PAM4ALpfnob9Br4cDiwmAmRs675GiC
vnMB72oP6vucEO2a/WNAhbFSvTm+10yItv8u7xyoaFkPDW3k0BlAPYLpCaktcFch
Ldp47VYEWD4jfyBkBylUXvLdGDljIwx3L2oFapTDKm9/R4v15N0wq7BtCSVwaaRW
jcM9I+sJCwhxk1NtPDdMk788CFAr5g0MDcyJE6z/wae98JDblPxenbbhS1zaXVww
FpvybDoNNvwf2Arxkj0oB+lAs5RGOD0v9MpQEeNA4gyN+2y7QO6wFD5sp/yNqZ4e
JOO5OOKHtcZa6eNCMR8SYtTR5fqHV7CZn19HRbVCRiEtRIJiDCPzrLPxGxiR8vFx
hSA3Tj9A+i+yGE3iOFYIiO+qFAoYhdIuDLtpQd2+A8BSYvAaqs8MP6e6YOAfVZW6
byAl423niL8MB4iQiNkLUIT9Crg8lRs4iCdpB34rnTcZI9WYyveDx4va5z45eyqR
Mt7l7JAmDRFC4v4W6QUo9avKLnGQ3EIzdQ+97bUE2Cy/iX9lqWskyn3CsTN6vwJA
r5B2WJmOPoOIrkmIebeP0DUD5Km/BZRS0hogx8sW5siORPPEL+71Dq3RAghcad8z
uvkNF/BEflL+w6g7fPWeB11/vhVE54/sdypEXszt2XGM/kSiiwXhd9rYkOQOuuvS
xpFUN8chw2ETgAicTX33rZ1lTEsbf2y51nsV7ZjcP8by2r2+h5esFPY7sdUgyiNC
0mJSStAnjuzy7PH4TaDKImD667lGKFCxPVk4fcbvKpdM+F+LX5rMPCA8VjijK194
pBtMKIzlyPO3MjH7KKD5kdn7JUWn+ZdNyl/Qks44iuIOBxFPDI0RTt/WwojV0HCv
S/I1LAv64+nHKN3VlT3tePbys+RQlX1KPUO9W+Ytw022F2ZyCqVEu0tBdAs5dCZI
fWMI02p8/M3feVTLElV3OsAxRVNuTFZKxRnW36Y1t1OtXYCVHOrIBhNrkmNqrAxD
ugU86vE+esEw8Phm08ElKnDjkeqUZ8ON3SaARik+Q8uJctdw6bsuWbM9uoHUpg1k
4hQ7OopOCmqFAn8TlS4QFFp9WI4BSKkENaFisx5HQUgFFLMmI7n5lot25VA+T8dU
x6+VwxX/QMm6CH84E2SKx+V+MKIOQNpHfTyfzaWw/C7dajhTiP+OXFxE59ihEtYY
5NNVU7UPAokLDQAy02W2SA8mUO4ANVvC+uIHP8RGflq6zuzpoqP3kvRYKZRu/V09
EttCAhp2ObcsoI5R6qitMTsvH444/a6nvo5+J+OS8H8a1Ax2lpnam0L8sHns3BQB
bgk+xubypN2vl9rKSIfOiYm2guH9aVIEge9/pxcUv+GogSEvgp5GNgkaITDdi+Oq
cBI8O1tDllzngdqkSGRy1XkMeZ2ROXPI0LpHcIrOBBcvsCBx6ASmHdrk1SImn7NW
mk0MOJd4OlccfAD1MEDFrT6cQ4ZMdBA8snpRwNz3MXjk13m0etY6dcKKJTHQpHH5
Nn/sP1nOSSfvF7ffymqRrrM7O6OwDX+/9ObBxw2qed5JseVLxO0Rg5EovsBg1nhX
f9tlIUGkMN482/eEfMBUnkV+Y7jqrj23pAOqNcBB7IJ9DEdWY6X7APJg+cSHdJ0h
cQxPJEjHo5Q6PXcL9p4ryJkIRsQRBSepLwoHdLlvO6s48qrELmLBs/VQu4ZYZRyM
go+LtISZ3B8T78/iw7qjyUaaHm/68u/HNRckw9lt7WxOQ7uF5Sj4YK3ERRcAtGaQ
0u249uISrDUZEp2CBYN6bl9dVXceOdb3cennslCMqi2xqB0NdAqgF2xAm6UaraLA
A60sbpwzdFRVMm0wpCnaneALOaoovllGRg+S0Pb97TWKKErQIrQgVUjbonDHpV70
lzQA910RLrXScHGq/EQhA3YIvHjwKL4tci4ARifj9KQPSZGz7ETm4+7DsJsDRCs9
fgGudhgzqmPTQ0ExAc/xxxZyu+ZZ94jVCYppyr8/sxs2xhqRqDC+IyIryDXU6TsW
0RH4KSc/8pG7MPuQ1qi0KfydGV+jjYwLplcEthznrkQOrAtKQm4O43Hwy4GXiO7f
p3/yUwXtm7DaahXqHzMUnUr0EGudDWDtSS776lL2AyXraa1qONhbuCkpLtEIGejw
qQHI2HV668ggzvYuDIMiUb9yZdnzhxDeTJAvzsOiX4qMi3BkDrExOZPKdrvySSqK
UFocxoFktsRccdg5S70oCMfEzqv3RiNfI4vp/Wva5DqN634E/Rfxvok2XID5M+xk
3+cS5ZnaaX1kR8yyz1FcSoqIgpeeiY1UQBuXBrNu2h81Haw5osE2yKl2BN/i1/vG
DgMj7KQawyKZDfhDoQ7YTjz+dmURZnByMV+SaupS+nWB0Uvlqd4tl315RsGMP1Qm
5ai/p4m6eoytEKdnQ4HJ4bnEQ9lzCDepe+m3rmHnkBT7itKT8LP3T0ButLJVFs29
fNqpMFwnxmUB2SFQJ3y4U/ti+DsfHfdx+DtkPoOaEW3zTnfzEsqsXQw15oxnYiBV
CGt/s+cLxwrKm2cvlU09sum0wMHuwNkX/EJ1kXCGgyybjZ3aIqz+GGjTQQmKshAg
frg/p/bn/+2IldoZ70cBRsAhv6BSl+S+kB+vvyS3KiQJ6fzPZqkBfmILgptGXSbJ
QDUpk8HJAX10QXEG5FJDJfjv9SF/Y895cM1J6EGxycJ6WDI4Zd5lhtafgVQk0Fvq
UdxXIRPIgXqjJllHPxqSI3AcMNReI88uRCZ1jniByfKJcLEs4CXOJ4JhqenC6f6c
/EItb+yZDLKwzfXs3D0hjyHyg6gOI+P705YiwXW+j1IQv7YsDoj+62l3mZeeLDTv
QYwsdhrfmSWpI7SD3y+JMY7JMCfeuGRytX31nHtSZl9eW/ur9IiPf1CD6VqURpD7
UCBLWClNsfHzoxYoVqJBTBw1U/KaOzs//Z+b08PxPFyUGaK6sKE3P13No11YzAP8
lYt0yGz8gGOPHMZULEXVc03XIHo3W3uazuykdXpE4QXgkILvdYZ9m4k0prJqSprb
sduNyrxWbRBOFOsDbEuzcYE5G7WIrZ3PDaxPf366/xLAMDMYWapuO2KgnveSisdI
grImJKX1K8DmnVh8M4vlWRA0QH8oqgxNLhr2H8S3JCkarDzY847uWvQy37IFhW0o
b6gxNYYlR2dK06bPOSTVkt4thTwYBaX+GJG2CA9Bmf9bF+5tRYJB4TE+TRiNKiqs
0W+5V+NHvf1HzBxxQjudGi6ZkhnGxluGtPFIfa4ACYD0p90cWfnFbTWH0H0pYW5w
69V/PKsB4spbU1YUtWIPeHxrwYR4BfYJKRg/XU39Y8Dtvms7qDnzYfKwYPDKmoo7
hlBaolbo6jEIQZ8xduZbMU+mJltnasGnZ4O1KB2AP3BgIvY59rR+4Vr9rphmFq+4
QHNQ0mFT11tEzt7c8gxyz0vpxXaZ/3j34js6beywp1RmpZmj225k3SopnqlYxJOW
O3oN/cipCjW3A/kCqa+AabVl7os/8LhnTRj5WqBNxU7rxezEFIMswhAzDLUF83be
DB6ErGSS36cXDzal2X4ghb99qrfQgz23G+ks5hOBFdTqEut63IA5+DJY/+4Q2+5i
mXlMbs1mURkKFlXszMMJPtbGR75B//2jD2lBP5ERG/xsiCcT42YBOIVijDQn2Xhm
8IIXylQ0z/cL64crS2vz/bCCHmIFRN25AysofSWBHhNc9f1Aqez4hvzv2D9YYZcO
9UuCVVX3a0yeME1Xy2jbhvafDxO2paObqjFMxR6Ly0RiyXY6iayOIdphuJ5IKnSx
jPJYbUeupPMEASRWRtF1sfPiPQFJ7+tbLVJXDl9YeexMD/bqZoU9eP8kMbGWVA5R
2xvHxHINi4BRTYEonSREe910ZzIiXv3p3d4iHaZjO05riGZp0a6W3LYhcwR+7Y5x
GOeiNUIW5Hnc1zXkZIOaPva/5nwYoWm/G353hO8KxBLyYeusj5yb355l+gxKRlk6
POpDAaAEUZDYVWXgoxspqfx/MY3x32kKsPlIJV/8hM5yAdthjLy9aReV1eMgawqh
t7XNWwriM/7V17mUpKj5KO6ACQVkhdXkMX40uwwQ9o1mWfQtuF4H5LPjuBejPoeW
MQn7md5xreHAMHJgpjek3ojhGNjejcS19mrlQxNqxUk/HsL2npTXuR6eUlCtFPYl
iS0uFYAVDASRFJTI0RLa4gl/sS8nZ+/bBbGOhUsV8k9oQ/Ja1BAbPMKKCUbrr+gm
iqLlbzAs9+vPiFX6enC9q7EXJpQyLiMITBEd8Qn+8jQTjQtUFi3qatrYabexB0mR
mwRLrCoM4GvaEnc2FzIIkRxAxUZ1/a40pXbrIeSEu+aHNmS6ZmYO0hjrZurwhs96
Rxy7XwMOxdbggRmzJ/Tq8HMJIx6i+0tI2TPT9zM8klstqb1wFXhyR3WeyOTLeJ2h
mUlvJyiF/LbfKExn4EcsVGi7INrauzJe9ApOwAbo4U+9Df9wEV6yyBiGu0t/sQj8
YGJ/ObtjaB70qmy3b1momn0Hc7hXLjDCGw9Lz9JUEgNboEoQfgQTmGnPgGpdT6AU
XOhOcYezTfLIVkKG6mA7RFQ2tlYp0QrahVKI7H4jgHtlOllAayTptgnLvE4ELhb5
2eoLVyhLo8ymYkqd75okLhiNWoWk2a4BBdKLaeXnFqz+jdSDzaZNGYn7UGpN83EM
ayz4BggXXd5ixl6Rf7Efwt/2OyT5L9gJhaK3e76TrJ9uYd3NInDqr+7Xc11P7zFZ
seJOaDdPxEQqOlOFn7KSEuvD/+FRYegcsX8obzv2qB/g1FGskknNZ6G0JfoGA7F7
tZU/JWVeg/bDAmM8fDHIQ5AnABXAMtMy66tB6Jk29iOjv2bKk4gkEHIrsx+bZo7B
K+qGPKCNWRgdMbkFA3XLL57Ms7lSzcX7cB1cwblc+Q55UnW1tsKSXvZdB9ptlxWN
Nrx7egwgfgqIAk5pQ/Agcd6D9lc5UaH0+OJjmjVpkkfi0ecPO6xJn4BJLdJBeAZT
0qcgayFNzgEk9a8oJmNZH5FMT9/3gmke+0y49x38jTLCb65EQL3WZ70tB8sW5Ftp
rAw4ERHLwgqmgm0Ry1vcvcw5LrncRy3qhZSHAUIdmuhMmyEXg1QIlnvxC1aashQq
edU9Z4dMvSCtXSwpG5+xDlmwLg5wRTA5iHIaPfoCuQwMEEb1CWwNhBWsQtD6jvsO
x3Jw1JCkoB/YvTo5YW+zylULbs8yhgIZM3Msic74S3LPfC9WfNYMkV74g6lqbGBa
hMBswtnLXX1D/Erazy9vA20nUX8/7LMgSucCzB3lrEP3DepWfaldi25OR/PFfDr8
BNgIgpSAzWRFwHf6FHFdHjGXy9Y0fyN5/l9+l4Ug37whOcQ7xkIkzzD5P9IyC21w
yAcDMZoMGNe9Q+B0K4B3ojihc43oNwNG8+Putz4UuKbCmNPN0HgRtSZUb4rExn3u
P59pKII44j766toRUlq56rg7iz/JhIAADZfmBVrpj4P55+D2CdHu8PaSq3JuTkz2
QM9oF0vQkmQZuk5d8UV+E6rempntoMcDP/JCiKzEjwi3h+rshgcT8fv3uJKi9Dlz
i7tL/3EHsrUnqjZ1Ji5d1xrEXzRc9JY2fF9dEtkxFhuM+UGndKGr4SGt2fUJ6Og0
kaDb+9rv8fyo+XU6VuhEt8Gkj523NIe4FqFmX9wNUXkiYaqYZU/P7xLf33llSAcD
jspnSJyAHiZVkTndxsIQzy6UFlmhruvzk7KUlN9SoUW6y1JDrsFVbK8m3Q4aG2Ui
i7RvGXNkgN8OzT8iUkeabNwyE1kDwKZisqX7OGlRZxqobqT9bHPSiIEMn5tKMsI5
eZD2lmWmMnGkYTAN8pSD+Is1rFqOX8Qtnkhuu0Jz+E92OE8Td5FWdOzknPDJgXs/
Ib4sSKDkM5+m8sQ0f1ehGQQVQzjw5EEMxxKLHgS6S1ke48uEiPGXudr0JXsDCc5G
chYzKdK5ew4h5lDRX34FDuWOBBK1VcZBaGOYdCqAU/685s6QUssCr2ILPCQePIOz
vkb5fE/SZKQKUNHHevqm9EebBUOi7V6HWnG/ZAQITPCOUWYvERW9T673L8AvyLtF
3gg9j+NXK2eAhIVoGBUE8KR9NKFcDy2xcE0uNrpTg42yoIdqs/rt0IX6oHjIwH3t
qWgYm9uKedBOzdH9DBs3E/CDTnn8dpwySFyLznOoMe+RthubrtyCy4kXKS0a0sOv
FBlpiDYdu7IfffWIb9MPnHQ1YbM8QKe+0lx4ob5Pb4kJhYSw/S/qRCcIunzZ9eaS
QLVNXCDZs00TBtR2SYm+KEvntUNL0F3C4s5kEwzus5m2NPgbXQmlv5sm2TAxAFfy
IIYvvbJc/k7NiUW+qhpcROoiCxNvp5By2hcJk01mmQoxmwWoaujYkkAYHWITQGET
rcMayoMKswN/Flig72aIfbx20DbvJOs3R5G7L2bafOitUvVRw+c0xJTwO7IuiELM
ZYLfWdGZSPA0JHjMQIErOHiGirYVNzwBGWKCEOkEgsmwtrlQb3fGkg7lnw6KidRK
slBVrBNgDwtopKHySx2b+cr/kvXbM6V5VOq+qZNvwaB0pbiWOfyHRR8tMr6xG9VW
mOLzJNoCFkf1PnoOKtHglZEGQfrDEApG2UhytQtOP5VlqVjq2cv0qVn35as4UgHW
uuqw3KUfFuPP5WqavVpPoEyYc710chioBWcS/OJWCpdFubSEQrXQZ0Nc1RcnCle9
pSIdMGhhFZKIpLAad3keprO2AKmDq6ZtTqWqUQXupMTMcMszfKW+slRM5zdkZMUX
T4nyrAKS15LPunp+YqvXbbC+5UoWxdDOP+K/pRYWeTB+LvDbgR+ylYfom79PApEv
aP/h/uPgD0FxZ7+9tlSme4oEChXBoacok1m66t+di7VB67QT70UmEdlGXHmImVkA
Y0yNtOscdk6hy6F1dqOKZ0vzcsGylnZ0aZxjIKTTVd0cqWxo310tnA67ltvdrvaP
7uVpVbFHb/Woa2jRs/JhBZKC+ORy9/y/3KGyxJdBJ1l+jd3PcQYx7FBO44+7BVev
3nrx74yd0lWYBhnYl6jV8Uh4sAAiKYNnfDijXVEf5hjW9pAxSyczMXJbIWEy+abk
X7tohC1bfWwJf6LIOVuGEaqsO99XoXzdhIbRVTP6hQ6LzEhQTuYUEv0wgZrIOLvf
5hjrizHNSmSOnLfVweGUHXQb0gZDYKLsl1mODWBVJzH9HOV3xRp9vL/urDZtzdky
sZ5LBjaG9nerYUYbCcfIaTepA8IquDpkPB2s924jwqd6+XGKR6gsleZ8Y3q4Z73y
VPwra0hIRKuwnzoDkdMCKbjFCvbFxJy/99wJmXUXQbL6CVoHyMpsbknk62yzzQFy
1liCdGBTAAh4FCyNR944tb5vxoVdcSDKTGJRsK8T8Reiw/UJSQFetAxowzM1jcww
2rKJS1fDyirp671LsdSDlzZcR7xn/KuDtOphLjP8UJKBvZi+Zf1OJ0CSZ5WKruqc
h1WmtndRehSi7BY/fhu22RBMZjgOpWidC0t5A0KokAXkH5WnVbX4B3PG1I+Z/HKx
J4CelARdbNK1TqJUJfYPfjBEErxELvCxn8L10vd9BXkjIPOQTyd2SDPecgHCMY4f
WStUoW1IX/PDuWzhPdY4oY/KVWAW3zz8i56xMyy5PYUiimwnp1wOEI6UM3Um/chn
2w6D3GwrRVsm84gcKAzZ2WhSDJXa1eJPAVh9JqlXBcr4SjasoRp7BqAXqhlEeKHG
KnsDPBcqtMsofhMNYUC6XIF+avbe7tVHEfuBJg1q8jAF2l9iaVvWY8pB6JZ5Nfmu
mi0wCEgplERpIM914YGe5C93zIK9gHtE47JQohobFS1kHA8Y0rrfxe+SdBVTB9sR
HEvvhqv4rtaozLxbf30Rbn3l3XU9SndP1lAOb9dB08fDi1gjoCocETRyiPU7wuKu
ID6vucSyOeFe8XAlW9Fya4BtV5WSWK05Nbg9ozMbhV/xuIqrTLYlfnTUawqdPUhm
28c7fEi6aLaPhzupTlpQr0t1CGaQwo9ZW3DbvAHHCUgo2MWNaBvJuPPMxMlJxFLH
+ev60zX53DgeZOPREsePd8Se2w1VI04DpkAbNq59YyC0oe6VYqKShLjD8R54ypHE
qQxsWOxHf3nV5ILjWW5Kr4ZjxKflK4BZOgJaVyPTD7wGxqHnOWd0OBh5YbAAwZo5
nFJzYoYBFQXrkYmOAxXa1J0MJAXwJui2M1gWh12niY3aWXzBKSMRlBR9omm6G49E
8ThuqaRWCI+3On9SOd9GC2LW4dpMds//g4wcoE68Dqh3RXqx1CSnaU7g9Ahcpm50
VER9nk3yLnDIMNc7Zlfsp968n6Qj2l37Z3jtlg3Y5dGjolXVEUW1ZkWq0fQITgbM
i28gdcTsURgDcrdJ4hr5/U0ZnT2+p+7hVH7xwiAcXPb2udl25zbSaLz5Q1RyeFTO
D83V+WgpwqEW3FzatkTVVnAW1XcXKaYjbntotLaz63qfoLFrq2IBh0UQ688Ld/qD
2L5GB7IZ36mcF+RKfoiRx1yGbfAHZqnhj4bitTq+1ag/5lQmh5S4R43lKQ0JuDtH
M64UIkK0wYZ8RQGMBUvEeup7XFVzD3TO0kTm3USkCN4ESVLToaEZiN46guCoTec/
MZxYQdSNApIeqQgn7shF1gfEVkeVCTFqcfTRDAsW3uE8diKODDNiF1PyGG3F+T8H
lWHCqaYHqScaxkcIpzIW5qH4y2QRBt3vDsNCCKDuPIUxoRqLx86+l/n2kIvlRAK1
1rDXrNuqemQb9SmUbK/+LL7KNJYW/DmUZa6iEITw13PcjVSFU/t5g5e+tpy8knDR
4U2USAXaLFfsSk3Nb8LKvHUamNr9IS0jnSD5NLF4FINWQUSwzBUrVhKVnZP95tZw
N3r2O2di016ADklNgNLc86HQ7q94sN9KeKn3iCrKk3YH/Jkujw/+pAKvK4UmRrUI
3yiXXNVRvRQmiEthyIFiDmsSpAKe2+1he7CHnepluMo12q8s7bbB5ifNonXOpynE
KITyXV746/HAPhPrNfFAVfZ/RuyyZFfqUTbN7H9LC4aLrziWgABfwXiQChIDNewR
87bb6JhJUYa1UJU8L1Ff0wyA3QzE0SfXZCbjjNiQbHemijiMWJjYkwML6vqDxjtc
oMf+tdoBdQotZhPZmAPGOdUbdNbzGk04+T5gHQsu9Pjt5fAnrYHBx8crn62k5y1F
xBpyhJsa/sM7gCgJKDNR2TAQyHoQR7nsjeMq3uowtG5wnhGw1X6e4Fs9pzGoeDHg
IL+1WLBavlCRUdwNJravF77JxKYWHS5qiOoXhE6ILR8c4NY1VzOgLAgbFEjGosEe
hULYZmrr5y1jGgjH8SMHrp3V6m1RSLQYE8Tg/r3N1DVgy4gXQ1U38pFeN+LBQ4TP
+3RX8hE7AZaDEJxKlvaysFrJK54ExmDERUi5ToJ+HgPlddpR3MZdGGATFFmqpg5d
+P3gT5e4KytXSUUoD70etMrjd4BvX3UYSZq7xSm2oRbfywk2+S9HdphIcKUdLjff
IlCT06Kr1QFVQL05nGJYg/2c/0hMZKXUdpA+kNKWsNJJEhZZiR0z501bT9jImPUL
Xh0qwUCkoNydJ72ZKV210lHwgqSI/Sw3RCKaFTSnpmix4Tj+LL3I3V7v9YuQavr9
pjQ+x1NDaqv9v4M6qWrssRqVGo9a/pNjom1OS8H69FLt4shSrfXtiKvvYuY+NYIR
MeE8H7h4p1KsUs0me2W18DO0anEZs1W8/8TsXq5oG6+xTuihW50SYmwHvZ2vOS8p
+Amq1yOww9xZm2Gd76ohHa34Sozy6dg4CiGpbY/xXYIt5yxURT3B6NwbuhT3nAEK
9Ovl0RtuMInLDROkQOoV8zPfo2zlCnSyL8o3lOtgeEsGwJUdxT5/x8cDl0NG/+5/
e71OicvIKtOmQALHeWNDg6Z0zv2rK3rk9b0oEtQK/to1tVGuE+iDjK8Mm63aM3BQ
O3iO17HRY8HoHHrGadz6LsRlGzEwz13R74BC032eYJwkt1fTda8hXdlGyJAz5VNF
Djhvd6/PgSn3Niyx3hxraGIqJ1kMUo6lLuU7ETK9yO4Vfji5HnpzsdVNJi1ULcRk
rPQ/8sIQeB8Ad8N+g/8gi/UnG12ZDpV4OHIbmyb2vD0G6+o6Vt9OK3MBP4SBYo42
NDhR5Kth9QxCS6qZrekkOPfPdCxWnopoojrKPs6KOHQniN4yQ/3wpiSY9pUoGch6
px//cPMgv7ZAaAJWNgEJ/O5RQdx6G+7dAafRSgubvLTlUuPhh/Onh9WUFSiUrb5X
Ig5a3SXOOd/SXE3jMN8Fyqy4bgqj93qZ0u62x0no0ZidELNipW6+eicyCA1ITXx+
GlQ2I2DZTWjNfMYW0QpGb/zCvSDlY+6A6yn3u3HZMuvZBtsripbNm/FLAH8g2aMk
ItUaO0CX6voPXxZEacXtxtFAK7ptQbFw9L8HZtaG8fJt/kLI4TOkKUxGoAYhJf1C
BhFWIvULuyiZvm2UwRTissyBdkmxw6K57etMAy1ttkQHMVfmZjx6qGrmyV96tn5J
1rT59tuG+4B9kqVrNpo3DiDKkTOQ61pfpfcha7FfFdNiCudZXfPqEreFXJm9Bb0P
t0OBjsl8QTT49e1aPNZb3Y5oegWJdz2CIfCk1pMa088aAXJYnSFuWb+p+/nIS8EA
cCOLPWy3zhBva7I3gybmEmdLTFDq7Qmwt1cnDzfqiNP/q6Cf5O2WvhUboen1NLY6
sbiZfjAjUfERdGGHxh7Uum8lIJwTVAbUMWOPZ0pu3agtlC5NwCPH+zw14vh1m4Sx
/rxWeii7IQz/tH1betUh24N622De01TUmZlwxfAp76lCS8/NDgSC25phGN/PojV+
uKdgn/qVKxf5k453h548k1IUz0jYPew5xAOEa128Ct9UPvs9g2YPx/2Ll27jl1t8
6GiMywgx0txxRLR8qBBoBgWb1B9zG1Tp9dFe8B7oF7kC/zq/7n4JVIXUZV42wh4r
Gub1teWZHhnGUzS8E2UZnsovrvoMrhgdabNRw1cqFbuV2Y6Xct31PU7XwkBOe9/P
7DuW+SPh6o/Piyh0q/7B7pzYeYgx9OrjnR3wWUOOzidDKX8naRtjIn+DjVG6rQsj
dacNaHOPkB0goRokuQHnmzjA73r8BKEqn4epqj1r6fxhW/5Tmnvvn+ki/k4Wu5yP
SyY7mWldj/Vgp9Ex90+shVGNZ8Dye4YEoafNgbYZxCPwXLP8G50QRKKO/CsYycAd
xrKFuVrO4ICT2PVnSZUpinj8jeEdQvMp0K/s2iUuHLZwHGEmwnkZ9z0dmlWdjrwQ
xdLuLKkjisvidXOyF82nQWbC/yJpiAUxzDxtOjOLoUtprYpg0m+eTqkFMEAKEMV6
z5pLRBJIDE7HwaEIVmKtA9fitTn9S3Mrsf/riBVfD+M/cS2ZaKJNXi8By7demSS7
3h5eWbUNZez/irhNqsSb1rNMxmimbKZga+lyasTg58gUcorXQNFkOyciIXu1Ae8X
eAOyciltYGkp9LthDk/jz/+zeZFjs3BRYaDOF1y6RMfgH282va+3HRCc8zUIVfNE
0So8YswraTuXXQ1ismuXpCF9ifmDR4j570VmfUtqio50RfbKyvJhdDkF7qOxvemT
Gtgzr1NUWOewYoFi6/BrxWl1YNMzphuSfDs2j6Ro05RJVBy+sopI4doT1oPtcici
2cNhc0ctDmI3awFsM3wqm+7nD3DJhBegOTzvhFjYIJXmTFZDIbhtG5b76+VV2840
D35nSKpzYkNE7CpzxejWXAHEiVfqdDIeRiqF2b+zYRNYbyTdBZUwP60T5UStJ6gT
Nsearr4kJUwnM2hLfywIjsQM0EEhCtDHnPeitvOadOMkLgLR59dGScZYqPRViS0+
I4JhEbp4sQ67i3B3VeYABIQDwOjzgSkh2QDlu1Iz18jqYxNNmdgVjdOruI5dzho9
B5XzEZ32FAfjXj0YYz3ypm13qz+hPUwXFosH/wYfEiElqT+pK8G1TJuV7BTABmvp
742gK5eKLPla+urWBgigbBe319iGYZVgtKJN3ihaKdj//zfUQ3gtl8Rjy07savZj
K9x1AtWMfN5t0QRtaecB/GpRThwl7N7avWTEi5r9qHR3gdxy4XQqPPMeblXOpx9b
Ok/k9Yyc8iQaPr5XbY2x14VoXDyY77NbpC3yhOryvX4hoxCQaNGsC1EnUpflRHkU
GWX3WDSypKYbVs/ektxv/gMHdQpgYpyhHB3pFiVI7FrNUNWs16zRS6en7JWAOsYL
9KQQNfLGW9PvAD026g6grR0EX8azzoY3rgzruLGn80o3q9HUHdDnjCqJXVufMeJ+
i/O1XCvOv96M8Qu7/aqVV17EUgmsqctxcn2EnEv2MRt5v4b5a2rX+mHpb3BMVgk4
/SFQ3luSMAHajirP+qOUo/7j3SeeE1Y0LFb+rg9iW8ZHDj4XU8B9TWeDYaPoyIRk
vIUpU6JcTTiNuNyrsJFBE3ZJQRSJQBdO8/wlgdWhw5yCbQWprFArUq+/sPoOUZ8C
iYrQdeQhROJvAdTKqv90x17aQgZWBdbc9neu+gdo0rhXH8hu7wDUMgj6HGPHKpDf
L/vPBMujdo1FqVkvcI2bhzqj1QWsObBy7fwNWpVSww1VygPN70s+Pl0OQS6fXH4G
4hW1m6tzfZMyhRXvhzNVmKzLfNvjJ3qRnCHIeI50p1Mja7Jq5U7HiBvTy2d+dhw2
5B+66FbZUK7x/pmduB5kKT5eP5Z1vWzr6YXgsqKdmae51zhQo2wbn45pYHU58nns
mM+vpgjgJY+vFi6jGXSZRU9i0YNrfBIZ/C3x7weRhmozyCDF5Xm7iWiXCsDAL9sh
DYox18CuCFHE+s6qLPFvVCWcvtKoMlwG5gR1FE/e43t/K9EWzUc0/YE2DMdxNC9O
Q6+AZAvQFNiPXoHS/IwyFcOTJNt+NJJEeVxCcw5Tj2bOIgGa6ABitVyMWpGeY1GY
Yfi+aGoTzUYqZim3CUT0opd4xnZktejejtbW90x7ulNJXAYHibzT0Cgfsi+pj4+v
KnR9VbcS/BEeL9kpHu/2UT0SZPinE/WBqOz8jtvNAOEBW8EluTe0VAtaj7u9fKoR
hdun4yPLNo/+UV/zLSTc/eNVOS+fOwqSbjaFpZFCMswSH2IVWPJeIrKwA0ykk2UT
i8AJg2UEBxJJPvo9lWwH2KcWP90Vzot1bvWLU6vc0fzrx/99Vkz4xDg3s/4galk7
zAf43Texzt9ZXLA1wOdT4B2T4e7i6m23TO8U1LoVIjTUf7TUZ07GPoQ/99AEa7kT
P5hLOwyXOtKbPo3xyom+AVZ5uN9NO+624J+kVAC8YOKai18TJlNBzaluflRv8ScN
dobMuxaG3JSiCXDtrB7RoRZj6vXfokf77iajXFYiqNdo+Xcv7oWd6k0VJ9/4MsH8
JWLn6ObKfI3RGUEa9/3jmBT1WekRUTpjXCNZ4+cSYWXKOKvLifvTznwxKjC6tHY8
5iBMmCuv5EnPtaBF3HBVGBEcQyuyoQKQ2x7oENWXY06AjE+iQF3qrk1Gl5K57jPa
1YNLl0TbJ03F3cAzomOSs7h8ixFKOu7BrArf0E34a14/4np+0RQTgoo1ud1bTUbD
0fQvWL2p46zNn9Pazql7UhmPU4OMsBMuRQEKn6NyP/ggIShVMdv335yTFDqzbRRJ
zONcx4VKNpysYM2XrwqkaaCbYcVFLAlrg+MIr5yhJ7b00u5x0xyHfartniT7Fk0Z
SI+BxEncvXqj8b7sy9QV4jnwDgtSIe7xN4bmvqEnF/84D2sqbZ3SxRDmbi/KvQ4+
0++5Mf3+yJFXHIg2VY8OpSqxd0H+ICn69ziKWGS9wsshcITfbvlQtIu4gtV2aOF7
6/uTwMw04AAzGB5nXb4Ee17VcXNKvfTIovBJ4ykoKXRwzclZsqpwulXznhVCxB9W
hSTJVBQO4Z5fN8HaPZKEykb7igEx8B7q3fUkSXrdcpYk/RhR0a8Jwd+vbAImRpeo
FNtthp7GHztaQoe16fB+dPvC6Q84E2YPqjJYL3dNE8TCmVMxSN3ZUpEJSPlBugSn
WOmNy6fXEIFXkx9FS+24B3xnLf3TbB5btN35WLTF912fLM4Iw640rMxRXcZY6q0u
TiJEBKBjD4lwtss4C3C7RFdOfjGNJRrseo91V+KtQds+Jg4iV+KL2VZRJK8IXQml
+A4baflav55Nr4mJBOOD0fJwwkFNHIVSlqd6U/6RJFTwUXIf3gtc7RxzmV59rg5K
PC+jxLnSWd5kL5QV7A1/6m0byQQUBsAF8tyeJ3hEueBo/e+5dwhEmuIdn5LZjJCB
S5Y9d2NonthaQoLSEMxeXVE2jjN9g0uyE6lTCi5svy7fyhYVIvA8T+hCFHXzt+vh
lllxorbgj/5jBYxfCKzqyqDSAyDuImkvSzJD0wFjA10cWADuM183iMoSIgI0p+bs
OdYA8Dz8nri29RtugiBfFcTaeotT1I7m14BadtSpDKfTTc9+3g9vzSawuo+83VBY
QTisebzBGAOnyBqf6pqdKMeAdR1+AtrbMuZ2ss7NQdDow43nYCtFgJKucKrdWvvy
3jqGvIo73Q0XYVjC6tdD0zlOH8t5UlHqazzvJyH9aPX76XnLkYiv/W9LkTnCrNNY
Oj9t5RVfovyUyZa72jdRIw0CAYEWwsJUvNX+Y4jHRq9Crut+G3L0uWnIt1zaoKfn
rb9MFAMWc0f98ylhAvyyaNYSA5BwmCHZZn14x3+JQRXm1magT9T5MzKslXNXS7lY
AJjvwXi5bK2ymEjXR5UDcy191ScbnII7WRRxoV5sDS+ETt5dfsOkyolqgUa0zZKM
83QYvOZ+xhUc/FjcSw6EAYHGS/G4s1FloFpI6/OB6Sn+lI2qRei85/Vfu8lh/ZVo
sn8nrNNff08HfqdhgyHz57hbuVZbDoxSzDrgvyafQGzSAu990KClBeSmUJtaNWyS
EKPl/nRlehDcTwQa0JoupGhClnEyoNlZ+3gx+HaHgi6aFe2yDojx31kWGVQ/YqF+
U/s4foIqFyt1n00xfARL9LnPv8z4JNSGS8K6r2xWgDSVUV3svaljV+64G7tnNlSG
c262uomElIOypjZSkSWnH0uZTRA6F5hq6+64utRelZDtENzzVAxWDMX6M6QiX2mx
zyeuqDz2fGS4Jgqeeuj0GXXRAiBoy7cSa4J1vNxLmcKGzsJ9KMgJblQdH8aV4tA2
bJdgllZYluOK7nsu//BOYavcNUGeFBm5OaLesxTFJCmJXeYiyHT7xoBZVHzXXZiQ
F+rH6cjXfZwz/LCnxFK7FEPZaJTiilKoFUM/Lyz9g5XCrXTcvDtRwO2mRHx0gDT7
aolOW/TpiMGx82Opk10Yqh03FjsBdu3Cq7qXZoM4Aphkq9uiP7OcoUTNSemx1UYU
yhbDnY8AhFa0MM67unkq/DAPqQdBayoNpeuBo5Xs7xQrhqHm+FzXmpkgZ1WXrLcc
niWyFIHqKmi6sDc0ppzcqfBxMMAmwN6Is4ZAaTYZKXokuiyIamV5tuxGpNLpgbus
sT49z+tc7mGJ0BGvxmozKyyT+oywOK7h0wvoPMTDfD+/ClZIcSFtoeY+e67dcixB
3z4wizGrcluwqV0kBa/9usZMFBxwTyZwoJVjJiwzwSmp6e9gW8S4GiI8gmaTUaUE
CBL62XdwOuCKO8jXeah3f8bm5cgB9e501w469YuDgAX+YKBj5iMWN+Ls7nmU+WN0
unT09sP9vkdIWNnB3uuEddhVNJv4J93HWg/ZpYvkK17yEd2c2g1UYVi0rGRAKQ2y
U0lyaFtoFTcP/1Zrpc0Dwk1KbI/Sz+EgObZvK0Rc3ztNQPemCsggTA7kMKe5+niW
WsMQLzm4PMOzy1YDxRQ1RJ0gNgbHk4oS77Z3HdFqIf5NWlj9Ftm5GLh+sEbOVHtm
FNdeNRmujdsixMFsI06WHznIm+tL+L97zX9e8AbXQdGU2j9FjADtNJN14mOiKR1V
DzGfDBgZYZsoKbMKO9JnPg81HUvcTXEbuiZKPMpFljVzx8YJJF8PGBnw8MB0UDbn
3I/4ocUn0F4eLCzEEMjcqLOt/ppeAUVrBDhqwxT+8Spc6Jm4yNSeDZkwtKrS+wFd
zP4upLPO3pdPBQakgwdXuRPRiW2wr/KwEkKiTgT4AVNdI8babWjiZq2qQYaW0bc7
MVZn8UN++kJrxUT19lEAr2jW+q8CK4vEVWIqkYsAK9/f5y5pkjLb3Ohesel2B6bR
7RNWcnq7H2fq4UC4x86zV1rwvTdsm8T6eBoEsPJ1gsBsKzEPFvCgydznAuthe3JR
zuTNtCTBwikwsmXWPECTx8zm/baDvlzuOJ73wB1tsgubOxlAgEpsOgdUhU1bfDNa
0Vv2qLJmhos0oJXWRQ4Pfa13EesJSrGUSumBHh/jeRJEZswcm5DEW+2Xi6GWIFIE
S7vTyDETU3TTja8mBpUETw2KxEg9D6jJErb4+8LZJifQ8fWpLO2Menkd1Gzbb34X
zyr92kpMgzCvECk48MGGmBbWUVndDtqXnIo2rfuk8Ik6vgUzV9K9rFXRxJotAQLV
BqrWnPbjtmCNR+X27cAeOuVysE4w+eyijAqExBCjQ+tJfJTpZ5KuMGjtiLbCbloQ
u56C55nJKsJgMZzH2aVyqhNuQKwGPWLCR4/brKji3eyyYPPGMJ4nF7z29NGbYVnC
TdZ5eWgJ9tsMWXx7Ryy3gZcw04gTftQqMz124Ln/taBl60GOHo/2pBurrxh/Y/NR
/KINnBzfLyplMxEfoPKggzNm+TALyoYoiRtHcF/L++gsq80R7MDTs6Uxg3u+J4OG
C4r8P74e+jWarOYiaBuw9nUvowlXBSODn2KHcttm93bA1OMSt80TKQnibzQ1OW+c
dLsFqS8R7OrdRMisSasCq32cfsNnfk7Kmb0bLUvPTILiOQHBRuAVJjmeuWZbnj3q
6RQ4B00qzXV6VQwRtfNXIBiX9Hl1veFnd89ECSwd9pyPsHwmbCl5OMTjg/GZXooS
RdyJs3l7BBub6E20cFR9C3FUl61kHxPRGzJMHpjbRp0SDg16IliLQl5iUkPNS8gt
v+bKiBSWHsDyvYJeiPLbDl1aYnxUSpeT6Ialr3AoGevYvXHsxwxIIsRmCik3c3gG
L0KOb2NdtMMROrkZQYabLIzje2+c3QByol8H3FVjJU34w/H6QoIs0wE649mxnFgt
cTyUm7qlLvWhoKiJflddqVpo3ibHvpVydFw3n5ZZz+p8LNe183fmUSWs74cbTEhG
Qy9tt7iTS1a+lzfB39160XdYJefkwM/2mUMZF02rFz4SsQHJusrLd7VtxT0KOMiW
LSwarPue93FXtzT4RRlkCR890TvreLeukrJdrKTfIdUXTigTY8etSOGQl/NXbY24
fBJT9Q9BVFeiG+whKt96//k+6TGTfhetlUgKT3aylDgPwMDSGBJ9o0LRIR4DYpuJ
fZIHG7U7cBh0ATkATrYggQBoyc3uTImDNvhrKSA5IgF5PeS8X1VtW0RkY9dz4tM+
jdhaWekfSh01TO48BTojosvhQWVb3QdPCyshtLxwcOgykXKHYa3ynqQIaBtdS+bj
0UjiRHN7Mwdgtu3oa2ahF3Iw3OlhbjXIad0+3uUN/8WyU0FjOgC0kYrjvj2sTKCs
I0NJIJtPaCN2dfMc2ZYMSRDoVDm1VWxq0a2X30TrE+7fPfFcBmfOh6+YbA+rOpl3
MIHg04BziZ7SoyF1w1lrSpV71l8EkQUOeK4ZwmYTHxwYgwfFrJol2IjEVm/wEAGO
XajWmXS6jzZ0m5ER1jJSkAnJ6n/Pua64tDIkrxrfuUpHQJWO0ndK9eKdI2hQtBMp
gINAh0ok/sAXAfhtsMJj5xmzKCIaFZbyxvRyxWwkesvl/lFj5tkKL+RPKBeXy9jn
gusqrlpfWjxVt8v9jfW7HbCb2XiMmphSQZZ7z8M5w1cGwxEpW/WYDadesuXhFuh0
6Jzw8neADjSKbNUAm05ZtelWtbTWg9P0dLZ09VvVy3v90QxFy88fS/0ZTMY9s129
WRI3osl2n6UDUrKXKrxl34xJZhDLBhEUPdhJr4gm2ERl2LRHpxuOj4k63oWu3qFo
atxJlZusa4Gg2xmWMaxEh6LO2/fW860gmMYu/Mya6EUXWIVkUm6iqamt0Ib0rj1H
yHV8qFf373b1QudmLFLb/4W73nILIKsoiWfDQ0dtKy8ZhRF297pPFsDcu4GiJjek
GwogjlYgk51NCGpOe/a7xNzDUafi9fVc3E2mDQwBw5ywKSMnj1e2/15G9SVHFJHv
U9GaSGZ2DrHkpy4bRxWB+i1R07vyfhWs47g4IEsDNjghOnTGKlAKihAM9Bm9K4lh
hvyDWBcesbUQkrcu5VsSlTtOI4nUq0dGkCqD7q9KUEa6tdGXJhGYydbdWoqgemPq
xEBdfzC0sss3pPkWwB2ZfvIDkAqshhwBeRINEVYXii6MmHLj+mned2lFJtrPea9M
PJzVhBLgyy2s9noq7opueyOhOwd9exY21DaslIhcLRSPquNDNKHTAdENpzc+Q8dN
g2XypJIpjluJaH5cbooD6ij/+kOKoB8MLfgeHOXj8zR7H0SVHKPDCpHItw+UlbG8
T2fZVd6gr2UAinwnOCJadcJy9MXG3P5sQTLA6ZVeXyM55u6fUNv/sKK9T9oFDaZ7
L0HNWrtNG0ZdQyVkr0lWW0JcESs5fePRMKe7ux+RxwGR8GCyrU70DgMM9W+ftH0Q
KfuP9OF+SSUDc0TIIStJJlPBL21FlZrp/bo6rISenA+ofqqbk3NqfXXk3qU+7qcm
yzAji5TO4X0UQhOVsEQc3zg2II4pEgRp77c4uFnjzoEATdwCRJddR8/4evP6fCFj
GovMG/pWVOsFf5C0+GwKcU8rzync0HhV3qHPPSQo9cUKXIEFg5FrJ8he5x7z2Rju
hGQBU5uKkjW6LGf+YpmBi3vf4pH7Iea3iQYXjrrV5sOC3xyte3l6DTDcMeb83Fvd
9Uwvj9gpeZTz8Qnvu355CzOfI5P5eazYqfD5bTG9KHp6rmSV+57hwP1uB5X7uWMO
V50rtYBLTGz7vdWO+9Ls1d4VgVUfsHxBjXXGABmTv1+xAObE2/1Vru8XCWa/o739
HTMx15SM53NAwVY/YPg3ZWTBXYC/dkJ4ODy8Wk1jzPlTDfRs1h3bEi8rov/ZH+DQ
720hMTiH6FlstqbzTm6x9F0BGedxVtcZ0DmYDmyA2bmAk+oewXYWPlBYwVQPJymX
GlKAFdFXeVmth4dDk6Kww+hbxwLekKtBl0CYXCRnwvZgTZzBTW+79fyR7vSxWugq
UlrXmf+Jv0iXwt769Zr93JSNnPzqL0XPaJ8lAYDw7hVArqVjG3zwy97b8RClm4xy
e98d1V1ouqfBVhbPB5s0jVxZyJfE9U28otEFZfl1Y3mjasU+2ZF7BOVrve4AjSfw
LwXXtQ9H0o5rQIC2ZZINCnImuy1BvcT8Nx9aw24FAlWV+WQz+1zLPl+m/VUtIU4Y
khO2evbz9n9ESbvUvjDGGAQL7CMzDmcpL3kYM8+YZZOhJ2Fn3W3rjBN1MlCu9cOJ
wNrShuPdN5EYFh9rgUaoe8driKLk45kDCpocHxbhEWCdQsbFO/4G6gpoBWDVktrI
1OOyj19xTDr7iHtLYTleA0WerJEIppMMz8i2T743R6zN5p8/MihJ8iT6C0z3LaO5
x0pInudW/f66PbYoofyFP5F012bCI4v2ds78u30F4w9NQmJ/k9K36XPfDgcvBtrQ
C05S79mgwwJWmwqlS/Kg+QC4fhc3ra8TCLr4QSaaV7u6zB27aF9ZPYOXG/gKDuhC
vLOyNxWGn1pmLk7RrP4czBkeB/8qEnS9YCDBrWkD208m9SU8kD+QUXAQFmaw4jE0
ZPoijPGkZM8oqOTWAmiwgJ4By2tKKITjiRar+3UdjMnKaPwo6Nd3rbUciZDZcKoM
4gB4zagLada9RYg7T3sOYSgp3bJdR/MEpQ2Jq1BN1Ur3iN5QjOQig7fjuxfsShfk
GoW1OsdjwQXX619XEh2Ta/pdI4FMQIsHekBmC6b7az2UqImqn/BHYiXw4/spGsOy
xI9oDteVimEjFHe2E7Em45UsgRCz4snd7QDUMLtIgHTL8CU4MMp18NvqHS17H2ao
qpuvleksCX3R3PicJLpCC6fRXIBnKTv+Vz4VYmy8A0rrwfM/3kO0sxSdEnYmaCcU
DL0nLW3bd+v0rtITKyu0oFOjHMxGiD5aldQXs0DCvOXww54xoUnhF0UqAUc1uX4f
BwI0Cc1iqtXgaewydQAXLVw6nv0l4uGWPjz1wAY8nYCoQvBAPIWxYZ/jS0SY1Gey
rHXcGVTUeWLLT4xm9Rkw3u99Mwm7qIArHYiuVs/8yI/xQikEfKRQYMLZkCkLDnBP
53tBOkF34hLDfFgoAX05OBrIxJ+xzB3vc1guYBlJHpBNMYIuSlmZVjtG3VWIzCWN
yllgXRbbeR0t2Z8uiTQh1IsoEHHZcpR+mvyYdKsh0mswouJ07UyzZ4js9pXqaw3Q
Sd/y271+S02pNopFjPy3bQaavPI9gSRe86bb7KJ8cCaFJUGdPEdsaVY5sA579qKy
xH3cYKK/1blNw5ds3uJjUEJbS/2wU6C63hdskRu022/LYvMzO9NPtjbyraT5o/ni
Ya8zwCP5zhQ8Pc56b/Kljz/BiECFcY22H2pnUpAjCozDTTnBhTcmnFQ794LYE09O
/r01LbwK1GRdE2CGf+CalXq4FypJO4PkY6MdUsWEYO389lgHLzl7Ki1D2H30puGa
yMI7m+Y0gxWOQfpRXmsMzoB9+ChSuJVQZv6eQBQU1OJDA4DQ2/V4WzgpwckZIJmQ
aUhahfwg6afIg9EU4Plhunj14Gdm8Vw9+korVafeFcdrokdMhDHkM+/UHN1PB80C
4gW3XQM98PgBlMWx2LrybOSS+tSY5wUZwRwokm2/vW9mXQn1jRiSvPWHx7nkEXy+
NYaPmgzV0bvTMPGG9HJOn2FCXwcRB3HQSm7MxTVQb3PusZz1RHszPk92H3U/9f/l
FFOfmrTyCvy59cRUZQS+K7mzidsbVwnsgteZzp5KHQN5rlSwceY8+6Ci3QxSc1lR
IFojAcDMziIH4S37Yi1r+dEaM1nW3Bvh8xo/Zy9Em+G+5W7YijKy3/oAWhiaC7xF
D/0fnxocePYEuFzE921IcU0Wc0cFSvG0r1u1aJ4I853WDyt3jiic/+TFIZ8T9QGt
i3obmWEJegU0I7Kc6tbl0i+LIxN74HzAKc+N5ik3PEQFOfA+Ggvgy5mjLAzivS9x
p6V9GGjZv+XSISv02OUJCuSnnjJub7A4aeL6mPC/u3QH9AzKQ1DCMr0VjkTUXHjs
nCWQduzOTO2TztsWAXlJQ3SfTCEjMr2r+thW4+0wN18Vo3wNE/QtoXaTxuSk8Y5o
tyIOAgfv+ctzvZWKh2pB4Ja2nqW5IvFt4Y72JbHvntDNWtB8ajSzotHYqyPR1tg5
koNYHK29CI0Yo8b1YEEjr+iL5bVqite2wC2umcjZO2ReGr7JkvkdScba/tsYZ/HT
nd1kw6YsWtDLGSlzChIBm64dUUmp0aMmpCpwU/BC/Z0bXnJL5QO/+1RIk1KjnMf+
nUbBdIycTrgLodHayl+KPjOsJd2Vo+lm1zdDGuwE79uD0m/PvSQu+G2LLRB4KVvs
mXzv7ZRHyk1fwdhmgSufN6yU7x1RjCINVvffisS4kNDsI9rV/zWn6RKOhas6qWLz
6xmHKwJqOACPvui07BZbxTK95UNpJU7YIpk3C3+EAMTjkMyHl2m4WqFp5J9LYsBh
9WQqTdxvpO0XnFC6g6XTUOhtispXUiBFTwBu4sXuGwk4YXb2rB9JuMSxvMU8fnmm
m4YyiB0gS9YXH1o5yYL09lmWbD3Omu1jcj18GkdxdM/n1//stVz6fycb/fsEF7hG
rtTr7e57xjwstXPD7kHYmM8ADiJFNn4P23wZURqCkJ9Ec13hgloEQWCblxPjHz5j
0SZwYGiaKZTZK4UBxseyo4UhzFQ0UZr+QwPEcXUaZ34QNmKnuxHb1ALcT1WYYmhK
MGZjrA5F+QNwBG+ZAC9/lgqdO3Y1vMuAqEZMLBFtrB0+zMzN8GZUKeychDvNFkOD
gHKF6HfPGYuemz9hUuE1jFX1D2tw6Y1j4fnYDxc6bOTpL+bJOAYPIO6sVc5rJvjJ
w3MXrXg0nFDGOsCrvjEelcJmeDPfSH+iPv1h+yR6zQWd2FhEnddeAOzsou7fo0cP
46BXEg2rjfEVmgpnabbbVWNKS4fWgDFu0577KtlDNAnzHWlFcZVTEaaCOBBK3/Ht
7ai9c1Gqgpo/kFf68y0jzG/Tv4Y/HxGklzhe1icn0rNAZlkz5N5em51pdk+NK4kN
Q+wG/tjX3QkOeN6JzoyHndqhatTEByjN87+gHJ4Ium60ON27MYujGRSQs1fnkJgx
XWodU6d9zt9jvlJJf00h9dF6Iw0jE+0VbXdB+8jvFiyxgRmf89fDd7JEmZkNCCzP
7A9DU2WhardS647DiYr0FiWTKnVm4kh36jsvy51U8UMlNXy0xZsUM9MlHAqqzJVz
UBxXqrhsXbbk3IMQic3xD3rJ4BPiBmsaBqbCGyS63E/SeqzAAjnNlX7OsQur9DSz
G/yF1wkl6LdpBfCx5IMPsZo/ay1fohH8kHF4MX7Dy1uetD2D9OiBeUHgG6T/6AOE
N9YBrU0WDN/1MGFsF78IwdmONUhToRhxDsC6mmgdzGzgGFXAZFU8BAMAAtVjwWK+
FpaCWhVEd5490HEJ9Nd0eV3s6Lop2PAwnFNJ98I3zJ2etrwaHkSfLtjhNhl6cSRm
U1jXypF0/Zn19PPcu8Cm+wAzHOpxp0kKwAq7WNc5zcGL0K/SlaNdVRyG99xt7rEc
aO04dKzTLsk2d05sjBY092h5D/KxaYAK5x5RTRmRra5ItJLBTbcaXcYCQxm9Z+lq
2jMiSgQ1XCQ4XaBRY+eDDguTpPpv+ezXfEWB8o5NhSNku52s5dv1WMCzbh9hzj60
hhE6keT6XvDBubXTOKSc8rGnCe1OO0oEtGlftxSC0pLPd2V4QnrXr/GLknQMte1f
0YI0tmsC7CBc/eNt5XnIwuyMqQKDk/kOBfMZmdERIM7o7KRj4alkF5rv4BB2g9eQ
hRudOXVNUAtIBOvECYx9KaQVxJ5JJ8Ssmg6g9XaOoJMTVM4ISMZr1HSMD/N0VUXi
RyhKac1/Yc3ITBZlt+7vfswJE3IdkOL7hnHSXZDPTu7QC7HpcrdhqIV23SZpIuLO
M168X7sd0hXVcvZx/PlJIQKfyiOM3OOQFWH34NtFiYsESwrHgC3XXYP7SFYT9lSn
QfeuagE69zWjpvg/pQtPHNnjKLvevTzhXLV6fUy2d/kqkpkomKYMOpQTVp1dFq2D
DsoVi1J1erOhkNNKaCP3u6k4FQCIkCNf0xOenxUBb4aXsNkf8VpOugpmn/NtzIFV
ba4/aMKSboAmr7/7wwtria3XzLiOWM82spkdwmX3m9NKoRBgSlCGEUBpgF+mUWzk
BYs7pPHpCa79WIMridAdT6lRj7N7K8hrzg6vW/zcOH6ATNeQ1W6pa5lMzss/odYs
Xj2hZSUQ17PV1gVQ6ejDq+CQiHrWpOck8Wsn1G9AvkAgXHquas3bbme3WDtHHhL2
LbGu+hz2KQAWzBn6aLAWzNAjaQXRbvI+x8L3XVy1xmmFgHhzjDte2zB7WU1WlX56
EmVAJOG2JId4UQyEAGkawYB29EdKjkfF23tTdfFxD6r7Ig+lCz2yWZslEur+wZ1j
96pxH+ziNY2Fnn8KW5d9to+3eNH9RxcyCpLQjEI1h7skY7QjLXdP/4evg5LLxaWJ
e6rMW2Tc+Txw5KMA9rhd/9IABD4v1SfylKTLlv35DmGFZa8kyFExcezdD5TC0bwp
F4wXUcP+kIMea1dfBR5eQQ4kad2IyrJ3w5EJboQT5ut8x1HVVHN7c4K9zjDHeim4
squkTfjrrKS7hyVg3PjwcZOkOsKgDXTEN3tfYDc1VpItMd+qBZc2+03cBDB18NXk
l/1nRTr341cOqsekMYDW9LcFwSVsroSvbU0+PXSpb1u6dikYdqGL8jTb51sKuyHk
ZbXqfW9MmXQH/DuIlZ0vFSqi5dO4tvCiDe80ZSJPv7oWOeh4s2bWnfOMOmIvTV4f
aHx4FEv+m0eAbqOQuZ3X+9IrdmNC31Rd5G//KP+KJx62gVXbsno9/E9sWdQS5RnP
/ohABLDK7ayZzKRsTDtkHPeJy9mmDR4rtpIX1NzEuf15EmCLMHT6hNVVgiARMcai
WNFd37XIVIs63Jdx7f23HcxaJyy8xuqIO/KJNdj5F8RY7m7jGlnbCAZoqj6ukBXu
5Osta3l6fUpMTGIDkZusWbWl1M31vk7FXhV0UxfioRmhwOIRstZeFghXCb3cXzBn
gFfbVnPdb1rGCZsiwE4rcAqiN2exIiNbswQQ146ZoPuoYwdLiKvmEPCCpcUIE3U5
itfcfPefWzUPHQW3WniExaznP+9PmR9GhNX7VlqvccmEg8BKtZFcnbWOMe0rOdSY
DmUYgsRYXxJTiZDAmp/G+3cEWdbWItiruI15EdSlmv/ZiWDcObC1J8WSWRwlPmVV
iW8eHTog2iXVY5VUrFhufZQJixTz/viKSu/9uSL7SXpCde/rkoelNWxBldTShGoQ
/baUtNo+HxdQeVNXyxilF2zy7qCOnp+BxqkTZu2RM/MuJT2bA40Qgaru07FIEVca
uONLWtvHa1tqnDwDxKOxD8t6Cn+KLOkQpBBPQjHMiSpBl/wtfR6iZNgQEglPgJlT
zlh9vmw8nQO3x8HrR9+qp4aeZAxdElVLQmUqly7TKlcUgPe9++y7J3DNfEYgZ37R
TpbIbATxbH/Ly6HvL82TbqnZqZeHg43pSwLP+6nW77w23mXl6joUB1IsugspPaQF
dCOIcxZRqpFZmmnvHEOTb6CSuNfWVs7wU/IaVkFOuhx9nz2nKMJZweTabA897fTS
d9ounBh3GGtTutwnJ75tAmgVCmrQc+RTtNSC+0G3pSADVKJ+9NpnqukeoYV8ilnu
ZYA3W45NgQXNoY52ABvR8xgCZKPPCFHcxtP+rFk+jciGxZ4lWDTCSg7pPV4PyE0D
F4PGY7QthgvvnyP9aq5QiJ+/F2F1BXyR2Prp3GvIQHV2OmlK7/nHwz837fT3ruVO
5Cytk/lmTr73w37noDrLPmt4dfFhuO7Hoz+hqcB5S+VKXqFgr1x+w5qgbJwlT9br
ON6cenKWo0lR9Y1CFIBtQ14Q2Mnfr68xjoqmCwE3W78XXARqAZe0sll4GKOJO7KT
ahDl5/vIRy1GDpmJv+DVG89t96i1oH7kMQGTiJGNJEq55TQ/ZtPq+zSfGxsPwhgI
Q3X63f/rwEYRmRWrX+8ICEH+DYKJrEv1IKHluCsik7KFwftABAHgsO1ELBPxDptR
YfvAOLkyjecBVR/rqCO8zjOWmitzAfuQYHtxschSMpP+IxZ+155STa2ja6kEUolN
ZP0CKcYGWgNx19TjbIHwZtXI/wqQSAb1V7kXMgenY24NyGrOtv27YLBvZFWX340S
sxlbzduRWamnspgNqF440qlsrM0GmK+EaWAsTZy06mZxhtzCT7XKqVwiPd1BTwAN
t0YIokKVFt27mNZ8S/byNF9Oe5kAOk5AWJ4bGmBvZ3yOrgecDjXZ2OZk4HR7IwO5
TPMrIVKnzJN2zyPqlpL9azIBniG9ZJNXghOTSKih5qaEtbk6AZuUiezrXiVe5siY
51JoqdHLnmt4gOv4Oqf/LBqSgKLIzTn99uTjxSJe638i6UWnttDev0hvvkJhi+oc
uLzQCFza3fWYR+uYLccGOB8vnXhQuHWKp5RqTlapYf00V71C9MTvzVxCafRfrQHQ
JFvO65IZmiunDmJDOCLcR4o5AchQVK6z2BDJ4D7dvSEbOJFedRcUnpOfBWIuV9oR
9omH01TwTzI8gI/9oINcUmgLW2NBJzL1szWgEPv4GrNnUJoZ7Uet5o7+545W7RUY
Vf00LzmHGAiIhepXMqd+upZgcMefwuSJ/3yc3/3iLL3q8dccNNP59EMXBEQgnmuu
Ay3bf/ux0r73LuM53t7AQefPWaS2fXAIWylQBDGI3o83rD++YGL1qAyo9353RRbE
R2Ze2QByCgIg8nNZRD4ucMtJnqvpBIRj3o95C+C9/kMVO6GhfR0eBXRbVgfApjq2
cu8k5+wzl3Jg5ICjJY+1xOC8JMZIGGs4zhKGtwEAX3UrIS09PAMzY7KQMfJ8VPJC
//MOAyX3JaVgmO/HQkPPvOLh6fBq9ueRiimCpn1TM4YgNwo8ixSm+QLn1VcbeFhP
2+eYvi1euvvwqyqncZAknj3G/xcamNz/QA53yM6xUigaU8mhgnVzyJhf3Bc/DikT
C4qzevtvZppsCJGTjYnnV1floWzFt3KwbkAzVnFuu7zdCo6sBORhhe9o0G/MSPYl
+5z2jj4y7di46mTSxJpnHxbvrUwdQFUIclocK+oB6b9jz0KTZFgHlrqC1m/5AOrn
mNLpMGhrs5rGmZLTI85qZk+bvpB8tzT+nPhzMCQ8AyJxb5/FH1yYqIeA9KteksnZ
q/RYGrMRDUb9BurzyrGuiEXzf/Ge1Y+6wcDZ68uN211YEeq6hss6WEiM75p7w7Bc
a5t0e5gQM2VT1SVbTdLdb0NIFnfrhxEh4TIGyGd3CGO266ndKz0ybFT7da8hAJye
T2sAq37dDkWOWXWnIESBv54C+8ZoQIkYGDtSfkjVgWvO0GPTHZNGtRy/CvQPh/dV
T+1GdO7l0FcAXJUJJudF92dsfP3Q69q5ASsT1Ty+EF9Vr5g0V0cSX63cvSFlJB9x
FnCZggRcHFm5Ktn1a4290sdosw79X6c4yLmxfyysXXgkzSRf9j3xaZhJvHiypWsh
05EzJqpVUt2yBuRTmbEI36brgqAAzWnPKTJlRUZmMJQk3hoGq04Q5HiyBOW0/ht9
ROA7cQ2GIyvUU5xT4yJMtRo4YdIbIiNpmxuPY/iekV5VoPSCCURfjt5Rf2CPCHJX
2ooPoxRh0noFadfBAzOqxeUU4vAfoa94Evgs48/RrhZ//2D85SAXZ2e3YYMc+SHN
Xbu6iQRwmU8X7KoSz55Bv7+zfqrH1ZeWl1j0jQ7pq4J0q5AFSjHUK0P4L7+dtgzH
W1NAm7kf9i/xUEHGxn+IJ/sKQbyemIbdo0OlNvTyNH9ErrUiTa7rfm7FKhV1cmQK
3ev5E8qryWkvmJs5KyprmLKdYHnv9qjo8V8pspi9Xzl5vC2XWEYYJDTBi+6Oq5Nr
+t19Sc3yFjhIvPwNfkDtNQ0fyQryBssCk1wPWnAoYe4m/Sq8RjllPzADUADftrSA
U46ptF5BqTESipKwzPuNbFk//r6+l/sgClUjhGU9e/uG5V94uG0AbJblq3HnOCVc
FPQ+WnX0u1/AsgXymmSMTEFHNiMcWNfukAIUHzh4D3EwYMC74V2Z4cXSCoPNstfK
Mx+mKvzcOmI5pjD7F7vmj03OO4S8BBIsudpeCTZJ7JrNhzmsoi+ieg10o2h/Nziz
oPy9uCEZKT/e/hIf7NjU6K8AA40lzqHyzPk/AoHWLNjDgP4r6IRJ/BivXdkjykWG
OcLzdx7z5unDZ9F27KJ6TQfzQL0tI8onekp2VW0piwPrTQ0efmpWqNNoAvBO6Qlq
5oLK4AHMcO75J95TS2Vq8VWapQqGYvwPU8pO1/GtBoOVWDms5JR1XsINwityUvGz
F5vTcPFfRXZC7RWyYZP918KG5r6LM2gKwG/oQaub+3oU9plzPd/kwcYSPsmR47H3
ZG0Hw9XBeMmbCk+Q1Stmt7F11HlOvbtIAYgg+9FL09rl5ke8o3jvI6q/f9RtV0HL
brLQAZhLFHadNX+Y0ZGl3+YWzP9XIKxxmBH8sb/p77/jN0PCTS4GpdC0XhXL0Xdr
m8IE5zjsk7iiWUtim6At8hoxP0LLezuiFQYhwSq6mu1mi523mPLq6F1VHjMisf5V
zqF3el+WIXDQA3VX5kyZmnK1ZQZPql8TcIHzqYtkCvnxWFqIf/6I8prkeLaH8nmL
gVKzZMzMJOcoOXzCiOZE1HoQCT+iwaT5sa5D/FvnI2CGraNZI4a7MqaA+9HIn9wG
gKQ7uwTHrku/NWW+SKq47Q4V2v71ZGLchu9l2JWEnW1HCyxaTnFBfQvejWXvz5BP
heOb9jThaq9+VdUSDo/YeywDx1ekhD3Kr5XVMusJCqviepji9mV2v8UUafM+bQ9R
Je37XQYS55eQGcKr9V8LuhTVzLI8OlnrRn6UWl/KYqjlWr4v0pr04n+/Vr03mPUj
DRErQPdCBZw3pUFe7h1vMUnGv/vpowIp1O2SCrWHhkCdwyov+/n5yYFecjwuVmLL
SHhqa7frtMUPvaAnHiOSxl6ABwbDKEjA48c3TQNLGmoF4R3GN89vdxYJnF7hyneI
plJQhrfLFCmyWx5T5lyyJPDYnVwt7fzFydoHGR/r4kyVPWitd5+/2QZP/QDU75yf
ZQfLNKvpGEdv0rFu8b+7EQRrSvfjvzMGkk97vA/1MLrz1Zthj2n+TRYtDwNugqE5
pkBqOdpNK28uZyZlRXX3GQqCLp1yBKXbDokefN1HuVBrTDoIW9zvTO1vG1EcvvaZ
nCsCJ2Ef2xU0qMUM6uLlk2NI/DnvGdxeeg52P0q/8t06W0v/e3lclZhLRB1vyngM
n4D4nq97TKdkgCgNcy7Q/j6EmOCwfBh8dUHj3w1ZIWaMDdcFQml3mzh+SU2hPMj6
JKUD697cSHqcXKNryRVJ/e1TV9/0dlW7EKf6XpDI5QEbZ5IrnES7HtQ3oMevjq9C
JN2beb1p+l0oXJQpyAxousajctQmEv9nb5K96ijU/AiQBlvR60W01HDkHT7q280J
WV9bEe8EHoP/Gc0HdtxXh7AVii1PN8uLYSz0atB8NI3R316Va7XDR9uUlrori7jE
cOEL1gLe0W1rlAhaxx9PpCGlJOVZct+bJX4kquXlMgI2sg+E13BimQ+aLes389vG
Uok0I8PFxXJSo73YCFZv7LOko/3JSDPUTUqFL10165ZqopKekq1aj7t5tddOvY1t
nY68oVocjusuKLcuvULZP9Pui46vACkO9uuqodVjdDpnGxUmAP/1K+Ug1xugqwXm
BTZVyLPBC0pIOUg/x3olUj4s/Xj3brniCKYq/gheZXMt5rwt45lWEaA67Z6vz8gS
gcpHhK9K9HTb8n34AdbrpruoO1lqcq3kZ2UNu/WRy6HTpxfHJz+iI3qWUr1pQRd3
d1YTDK+gb8R2xPZ2Mtw2rZKVKVyvId11R880DYRUgEr5aIkogEl4Uyyj98ktmdvN
VJ8cTP2Y0UcclwhBq0uLXBPwtR1QGTbySzjLIR4vC70vEB/zT4XBbndIkmad0Ng0
PKq89SlyDNCXBl8gqodm4lpQS2DwLn4RkFyJZqPCcNhKyW8BbB60lLdi+fJEZixU
VMq+DDu9/kBgkeB5tPpUD56aTovbaHrTRetJH6odezZ4KuTJw6ZZxXYzRUrEOGsd
vPajheBVJvaOSQF1EYfgoW6zu7GlP+lHPEJAd8AP9qNiv0gxKePHqvTvKhrBWmUs
FzNtJoavIv+8FXBMSbLJqeOcBGdiS2d+i/dp+p89seIWpwtVWNOYxWLzaE4pYzGJ
4nJi7oHVeT9SMo9D/aVx47GtDHSSolxvWNsVhbzIxYi2iersYD/5diQXzfOs/yfA
3pxTfz5PeriQx1MA0ieLf06RagqYaIm/G+AV35ScGbyrJYb/aA2i6eRkQhcl4vw4
E4xgCeO6WRUy8lyNB6lfw0i+cTeqbGa+i0TsYVSId8CD9bjDOi2Ccnd8vyIGcmrI
Y9dApPdymOVhto1aUZ55XqDlWAsblO0jgGkFpGuphTXf0XNh1pEgEKTz4W0cfgnD
i1bJUslnRxpBJNZe5na9wP96hMCQQBhTawG46Qz6bMuaFKCtC9uvDbJX6Zk/Huvh
SHSLmtwnkfgbsUBv1qN6KzM7h3RQojEi2T3jy6XRArU/ia/ErWriGFGrT8bKzJnf
ctPjyuZjcl09aTsmxGAq4MCUfejtkrNwuiH/fBM7ujRLC6v9SzyR3ZId/5kdoiC4
X40L8bp2/Hm34BrmTzhrQzydZB6oIOujZh/6SsObOdQlLIcJ6VBRfjB56J0H+CRy
l7tEU3BcAmDPc5RriAyUiQH9PoNStId2Rt57UglvCH2+8Aaq/8ngK52EQCQ/5U/1
k0ga6nCtD5cGx9CsftFoEvRYOlaJu94keSoqIUhTkc4/AwK2Um2KzI87R1pmmZH6
hFXCZ0J0sGwWlTDors8zMmZ2j/XmPtyT4w2SZHWT64JDARJzyyg5JyYMouKLS1yw
1iKgOnn79PYbzU65LoBBDtlX34nVu5hKIwzBjqlsoW5Hs0cEzHr74U47z0Divqn9
S8hQU/Gwimv7QYDBdgRizZwZnIJGRDlmcLuhkGwaTjnnJ/XsF3xdOqRoajX2TDyw
YhTzgr2N9UOWoRnZzdjc3wEa7Vnmb14gTogWKm1k3MzA7a0pPjWQu+cGhrrsmjzx
lAF+s+n0yuat58w8WTuvBBca9mbnMMmxlPIvEW+3rj4/3eNf/NxlFM0TV590XlFy
WWok056ex3CyvAFEx/h97b34f5+gB8APf8MlVWb/DWFROp6wJfVQRuBvyOHjjh+V
iKi16y49x3xqc5/dkoRzILIIyMo9D449pIHtyFWjSIOjwUu898tKI/qN+znEL2Ro
1UNvFRY+KyIN8PNiLdH36W2/sSoGdxdKTqqXl+52kKrsL4FYPIFAkqcc3HX6B/VG
y7pOrEJBYXfCd8U36iKSwy+HdQcxIStCbT6FGIl6zqm1lW5f8MJv7OkqOkaqbdd8
Qr0n/ub8rvN3V3bIaHkSYv2j9bhEsd5svNe9E7IqFnkqL3ssdp2NJtfMpScOXoYc
WBR5VaNqPTpSUh+/FLx/lPJZEp6QbPjwmMcN7PS2q1zJ5aWdkHHQBxwE0PX+vVpS
dRSb0Jmlq3Q8iHrkm3ydkRa/ZPexYd5vTWyRwrI4Baq2fK+dt8OllvL8kumRDT4X
BuVsWtCZxoDC32g8nvigTJw/v4r2jXktR8wRYyf2Bo6ghEzJaiNeVkBz+pAwgY6Y
yqv+QtVZJ9fxoH2UKBdeKfNAW9Z085ltNsNMzl8t351cOB87pvZajpjxUJda1ILK
vvNojnSTC7pW8cE8lSuhjnXJ8wBj1HXBDBx1wgVaV1lb2CIq5j0C/pQ477hMync7
rxrVLH8lr2nPUwAZw/FkTVsPUr9KLviK3KG9n3L28pNKKYviY3xTxpuqd/hFZOnj
h035LcFFdevLqW6PkU7cWgchNpt+YkWq4VLNjwqwTNZquGsfcp+CIFOaBA7Jy9qk
kW0ZcxF2ku09vQEcHYEhcLRMfZA2MxHgTVFcPGsiYaGV1FZMi8xZLo0S/hy2wh4c
2cPLBNuzAwwJjDV2oZS8SWmp+gk+bsDpge32ym0n/QsnhUvtt2TSsqvYS7mWUAQb
ta6LzfiSMqopiHss4k7yETCI/11Y2jclUEemao2Hky68n5FhKHMl/CKtV/P4Cpgt
+eFIXZ19/eCCzMTnRIOukK2rmYeDX7ERSqGKF5a0aEdDTmcG2HhxK7N3IZBHi8V2
LtrcKNtKpM29EOVht4RxdAzBUwIAQbcia+4f726zIWy6B5TAPUEOtoJBLUiFI0zB
xB8gXNi9maK3ORB+3tf5nzFppcG5VnQz35DFy1CsP42lAtjdR3mKFWpRe1Y7pMO4
D1EETHrI9mCwiw9rUGopRu/y52ovq6esb3Rm4H+19MA6E66s4IT4onCfxhW8klbf
amsUDWzEAGfVm2Gkd6ykHzzyGrQgqS5kpYcAjPU0Ii4UmIscfGN2Y3kC9qg8HvhK
Fqrs/u9xHDZTuz6qWnEquQ/C06HqSDgVoVbYcUS4JAtS3sA3GS1YJF1i/YKdCd6r
DndppId+z9Sd/A+ODylTEqiMnP6VdKidP/nezIoHStNMaT79UWIQH0SrriT1DNel
4SqMFnUKuhW9zBLKTU01iQd2p1RvxWJkQdG1WdLIUIRDuKDq6CprYWhK7ZxnWSd9
7okro7TvnjwtGAEIzcCUoKCQCMsdP+1vrX0WnY9atUzCs0u/GM4y9adtkq2XATKW
5LoJTw8eLMZ0t9fyQ32Y91mJDXeR8ECgOa0lTbXAx1LZPBQLQc/opVXv0og0ReuV
PLXERrzhWlr4aSdxezSfNg2VeF/cj5HYu4AQhe82yfLQj0EI9j1AbxNoNDya1sDh
RmzTpOoI4wgXy6g+BtJoHIwDuWmwtaUeeDLGK6cePA5/yshE0y81YoeEkzvEwOWN
8nqYqReKPW5Knp9HXP3MYZ+SnbKYTKFfzfTZGw9N20k5lHI+Y/Et0Fk9z1lw+kD7
RY9qKZ9td/tJjGC4UDGSjnbhyu29XLJ/193sXABUR4GIOntWSkCdREyrIgPh2ZAi
+NVyeDA1VKIvdHSGZoFTude+N+blj895yzdVrUGuZeXFf7D33yVGMmC2FVRJ7wdV
aVmB9t41nLD1S9HU1qC92IVNZIkLv03pA3KL3eNsTR+5UgbAX9JgNvgSDxFpQD8D
XwKC7kQZN+TR06YNW1fbDuDMskROuzjBXjDKma3KABx7+JF6WuCoYKhr1X9TDlZz
nt6p4A3mu35ctm1nw24eiepYlts6YEatykWGO4oCMZ4pcfFaVDYiakhE9mfwm3VI
ac66bVVzBfbChdsb/Ye7f5MG4hu9tl01uzKyrP/R7pLTpOiVpA3enVynKGs0N3Hx
qIMolm7P3JjdLTKaLLJWMvIKwZ1sYQtPsQJ/KJ7HYg29bXkEnshfA+PDLVfXvECl
pylxOzsN8n05FU0BsHapYyubJsfcXHu7+XETpC+iH28dWmoYemzm8uf0EG41HaHz
NvG4TssBh8xFLrqTTJ+jBvL/k2JQTgWcipNw2x9ts1FDn8diTdRniy/VwOxFJ9r0
63YWrY/vtgv8Zn1g/EEAeJOM1he/D8geg6LzXSY9Ix42j+ToGEhJf085JXs2E8st
Bzx4wuU5T87RxKrhNpBwVcKrTPHtFEZ/2cSVEHebFUdb11HMjiMc/PyXsC+w3zhT
xmHkhEwynUKXSgOghkDxME8DMwE0lLIzkKQExPi7puZDcP8cEmi9eGGuiJGJ2pYq
UTV2oBd10hG+slEf+wbi5oWyo2bui1ZfWPTcFp6ljLuaPTDXhd7bpGFg/8GHTFJv
+BH3ylc2wJLa22MIy9hbc09EKh55Eko5TDKmwMd9Eoc4uif3NS2oJMCq5e4sNKV8
F7NA/Izz1AS0VdjmPhBRel77VRbHlvN1pJ5ZdAs30vfwYiqzRBZJPa89idElBOWS
QXf/+d2uVn57MTA3T28rmEX721HzubMrb30bcgZTKvfAsezMmJ61sQ4KkW9qGMYy
TO3xg0G23N3C+2KKGpw7JOWmlTdiFcsC6nHIetXCrPW+kcZz8Mmwfpi6b7PrqT2a
guXfjiUFe0nmUjU58reROULVvjPGEFJov3ZM3kX7O2tuj4ni5onz+92PJspRnFyG
iRQVr8tIrZpuku4NjMN9h/6Mv9YnT1r0kL3NQ6UD7S7bCyPpYPpi0ewqWIqMa1wU
33s++3bDqsMJeH4R2vsjO4IVmnd1fw+JmfrY0pez6Pfsy6CuwhtH1oBhOzowvdOo
dDuTaVJxfnAGH8apa+o3jWpC/IxONbdotNksqawaEfMq3ad5Nj5HtSdxEhsAUexR
0X0uiauEKZoeYYqsgTYAFH6rba5TvPw1RcJb5DKoSRedq8uAfWrOJi5tt270FMaa
YNlRSRycYzQARMZBTIzma+XskU9NKkv92fyWDJki4YK9BpV0YnUj+1xUMD0ElOI/
TGzJH1L/YEFMatjfqFsPGcV0vxEZ7NCruFai+yW1Di4jLP898TxSOANOwTq4AEuN
NTL9DoJYAehNgSxAiPZzvD7YF/p3yOCsgbK28njfXCY/CQO7mFYB/R+1otLe2ZFq
nsKnseUvX8PwSI8FJIQiCSrfJ8zNtl8g/vopn8l0YrYK2NU6faDyFN7Z6ZhIJOY1
ry2IBgIyqQG6Mw9WiJ+AMUjvyBFQulNMcRyPsWK43qTXV4EyCCC7h7pO1YUMy9I6
YIbbhVC2+i7g/vX7Wecsfn12Kv/ft6A5VdmdYo09w5d86Az9WxrSI2H95dNrUg5L
oz1q8LmqAdL3Eye2+nL5cx9hX4sPkyOn6K2iKNb+QMAuqtiq8tPiqy3bzQWNnZq8
iPjHK95S7HMPO9PGhpwA9IflTOPBUQVN4SvwbGg1CVhKbSjgpVy619BslnXzBxWg
unpHjoTuMc1+OcjLpJ+ig+6Rq0YXa1rzr6Ybh0z3an02l6qM+wNdC6ehUfLBi27r
xxCAO9bst7bMgjQNigjdkmJnUEcpEukkGg76IlMa0FnpXVCveLdR9TJRwhkNcuoq
ZILOZKTiMMozluV+yxrylp6vVkVAgA/jUPpZmZJjQHRYxLuX2jKgWXnTJA4yM8Yu
G69ue2QZp/U69N9JYcD4buwgY4Jn5lbuciN1J7TI6blmI7HlQXeL4i9puT33ZILk
e6omrYR2FCMT16OO+khfdjJqsISeDu1bxbIeFmcqdDa1I8OygzBU2RWaKpBjV/Lq
BWy9RxLJM8Htk0fUIGaDEbaXQJzP41P9VtjznE7E3bKqYkoohC3zoU1MFoyI871h
pnFT8702VUgprp8RwqDmbJ+Z1/xH4RYaVV744bSgYdA6J9Y441wZM270BpOnQk2f
u/UJBO54H4ZSJeMbyCQKuHclmvCuhyAOI5r4vutFzwtLTl9MSHdVlPdwuDj3ZtyH
t+z8/xCZAFj1M1XRxbE3TboUslX9pScc8LX428SZ8BtSdXiYbwSZJ7crSUadQPIl
INLZpjS5eur7W/YRgCMweBYYj9uhCMAmgtU6TF0L7zjryZ9mzD8Yh5P/mRQjjRoW
9PPQV05SOZ2fSaeXBmMP900PbmzAvSXwuOU8+kO1BeeSJSiilOEBuw8AjK8CbNBD
P63R59PAoTUoXnkVevKTnzWpR7J/eRamSnGFQLBirOJKi7EF0qXsCnO9XR8fWDFz
3gztTQKyCbQ66rqKWKhMFShIwYrgj2B+sn7a0oZDOfdKqg/qJhjh3VnIk1kOVCRY
1/gTDPjv13iWSa66wcx1GId7UIJATutC0FKJs8sXEsPRpmsT/Y6fnxGIEMFkYd5z
K6rsva34yWuI/BtkUcmOrwaEUqR3r8FcSaAE95TrHIK7LxmAlsKwLw1UwvdItFvS
hSZ3Z5x38wa3sBVmIJtS3rd72ma+urPb1o46jZu6LXrNsINWd1G28iA0qlWDZO5x
dYrTFlaH2lXFgGmsaERbboWbTkEn5Ym2lINBtwun7zba3MEbMFcaDQARFKeZteQJ
LuR86PeNH7fLsEU4cNhadDTTxtkWp+b0pNOoJZxvl5tccjt1MjdKMfpE0f2eftIZ
9QWr0/zdnhbQFab1LJG2Rue/hB/4umaLsZPl+UUJ7omzpD2Bca3RFkoXzsxsDQYp
bSVmPKqiYYx5QadFxeeaDRI3mpxxArG8XpLWi8dYBSNfjymDl6we0G0I2TSJSKIS
eyEMTJAhjJ5A83UfcMVpLbs4X/5zO+j/0ouoN09DkNIob3V8zxBcx8olM2qvRGcx
4a8YUr2PaLuUrSHL4st+98fsKJqQZKOiPUVTBSgpjZ07VgEX26qGAvbCJPpdazGq
IpPRrZFBqyLFZXn7urfUfpK331zNY/+pAjwsheae5Wc5OrGZsjG1UClsxaBfbs5S
nPApxT0APyahkQlMe/VU2Mg5gaORIkGlvGNCKIAJ9em6Uyj+YIkPqfUXRENV0S6s
qT/L/USFUPwweOipAlK5uSrYkJ+O6cBKq/f1eHE5xNmO7HDnsTPsu+jZvFWUIVjC
uk0pQnJxSCkG4F9bCh9rSdXOjcRhGu1xUep6Q5XysGq1J2CFUDT23x9+JU4JyKtB
3zUZqWl9v3Ifm7JG9uGfmBRcGStFq+8Nc5HpdGwxPdBc4d/OF1OEXaVtMq7NVKpL
g14Hp/hiBhO6jifZRQvm4XCel7W16mCTtJ+6VKvkPq1UQApo368yv12k7dh9Ai3m
7QlpMhauR1Czv9RHkM+fY54gcVpvdMUCEm1247/imKtCrczr8wDXsZ7kLzBBc58l
PCOYxhw9aJtPE+nYDHpet9a3+pujRGjOuhDiiJUrVcSaL+wXcnLoiUqpxdVf4Q1R
2nqKGsFMwPGy25lJC6s5pM5nY9IGagLbmNSPn3zESviNx6KRUfIUQMXtlZhmPHhT
jZ7LT5rsagUGgq+T2ythJb4mXgq/5//Io4Tf8Nnoj3MXgwd3d9Ejw9tyhQHvghCh
H0gitM9+yOV6lCTPE54Aj2hEWyKHZ68Ea6hOSiO3h7I0M9ck9wjnRKtBT4ZM/4mi
NI8itXrPSG8W1IAe4BCAuap7yuK34zQmHfaWwNySVFhh6qVCvbDcHsJ/24XyKqr+
mstGc/lvKrVloWivJoJL3QK1yZ7h7S3Fe9lj4X/+vy1CIbELT+oRxkvYCily1n3k
eWlQtDUNkx9BvXSyeTf5XuV4NNUGxQ210TpGhc0r/I6cBEyCGPd+oWjuqhRL38Hb
PxTjleJ7fWmaiaNYxTtu9uEVDKvq6iIz+kX4chSiT0psYIBsdEkM2dYu0s9OOiFI
xOdgXfFidFcQrUZpYHUfetDkOhcI20+ZLUyUT1R+402GLTqaqIDwnmgYIQ52X1WY
tAa6Iv2DzvgA9nCWc838Z2m5/hAMzcJ/YwZQVECngcKUuNrRk3ftw1aYnLJY04YZ
Li3xKmSZW8YLCJkghMM+F+7aAeko+OZGUN+YVHwqDh/NrlDuykGMwI/I/zQvJthT
8kKd9Fk6bHc9Bk0YeIpUjjCYavh6uxUP0SmAvS+rGoE3xHppmmHWWj3CgFvrGrJ2
bzMzPEbsf1hJraqDacJOJydpfOz/KdkxBsv66GEUmZItoRStKyDoP9a6Fsam5wQ+
Rv8cVRliq1tb7/hEK+66DK+su6i/MsX6zUavHJeU4pAKoKKszmogaPLgCd1kgf/E
Yta4Mbq36wBYc6lheYVlcrgj5c0eqfRhnLa4s9bvpi7q4MF1i+ADjCc/KJ+9xi6h
elpc3HfIQ2PUZko9PUz0z9aOSzWz0n/j9+l16236cMvI+rSfa+a5sE5bBbYqCLBs
vuJIS/iXKDwMxrzmekJ45BNIhLvInZBFOrTCm9gM2nITQuTrgLfAWWOjQ7p3Jt+H
dFLhd29pSpGnZ6rqQPW7j2OMW62JfXFz6mcF3HidxtGzODPZPJaxAL4jMkikXIQ4
fQtNk2fDHK8eWEMSU0xQCx/qSgiTdfhHktke2URpcbq5BiASpwFGfn37KDHFrpU4
R48R7uBtHanJHOzrTu1Uqn2LHmlQ7leKjoCuOvWjnX+RAvw75TV3l88BGhSN3gO/
/ZXJbtDX/0imGayeb0v5L3HV1UK0jbPY+FoVa28FogNbD3EUc4U0LJ8WwmmPwRM1
juTNntrwpwbHjchivBc8MgO2mJmL+blr2fKrY4VuFB+u+Ed+6Qr9uD6kSt5T8hPL
4ElA/upF623kY1ugcOHrBtCjGxwsw8OAyuxNDflb9Mfm18gPJyJNcZdBVHJczhRB
Y5MA9uC39dEo83/BsfQ8xDV/M5qj6G/xPT4GMx72gLV/F0QZ0EJPnkPJagZQmh6J
85t0Uvl3dxZMQxHQ5i72Fp8nuZGeW7UVAsr7DsOWE8W2jzcTNPGOzmS1x/WaxHLM
gCxu6MKIBEbMEFTUXvfAXTj5lWnebwu39w4lIMvnJGaPZjOMFTHDL/v4NufWZjCR
80aTZ19SzLIcSYjYdnXeWIQ5Vd30gOHat0seaRzan1tyJotFm7s+Vs8dnmGYOcV8
Et7CtUJdEDejtrnP3ky2auSg35c0mxy/uAInyYtlFeW5C/XF/teghVJRXKuBZbNS
5wrLoNHGN5bsDGsVQnEd+QedV38n5xXxvcESCZ8QxmXiRd50EcTg8X6osr8WdwKL
32eIUKcGiSOr75EKcFqxzy7tEc4QU6FO8vOYjC7e9QZ+9sjS+EBdhwmYCIpjDsbU
Sg2GHA5RGAGrtTQnIKqxPg4A/lBIb6ySkg3CdfqX7zrH82wAivtUSKIv5L6P4y4D
MLO2CY7Bk+gpIulPQ9EMyph/D7OxduunVVZmReNfviuwkocggn7zITOehrvFEtjW
YXkEhn3C52ehs6HdErNWkMDnwWo/lUrvqFzpR9/ihM2kmWKkqHa0W6HtEj0CYbLp
tcslrvVQfdnGHiwLNLeI32aPp1P2/LfpRImcE6BucOJ2C256UJM22e46iKPyxK8F
LXlsFIWd5ENPz7AycHOATUSVF8tQNWsMfkAfH3q5lBkDBMYEkOlvCbAP3pe86Dz0
YSqLFNH4nCKjU18hGEecI62V2myawLswWfABQYWn+tjoR7hENmpsNbzlX/18wlWe
Xz8NJdzPG9yx0Kt7ZjABLkVZLaaHBB8rdieMwdEn0aKpdr3fWeLj8M0g9YIIAoEa
oEOyMncQrhxZ6sBUxFLUD8JbiTapp00zO7lmykpyNojFkzLoE+cb2HeN+W0XAJRu
IkKyQo3JR/NR/WtPUa+dfFg9VtID9Mr37JbTeVHevh8I6kJM7tnQNgq1zJFiDpHv
UB9smvM+7j4xecjDiZgkl0Ilgy9sb3R36Tc1Un3up4AGvjIo5dz4bO9tznZuJIkp
Nh5WEfv3T1K8Au83yM+QtxjG2EWNAYlLor/y+uvVy+9ShiHdHFeYTbl6IWUdK21U
nS/kL2sm3DjcKx4pcodJNE53ImzpL2AY/NbxoGjooqB+lq1ezxHpA/BG/3Mrxn5S
fIiA16/kNPorFlN2HVSxW9dxyJBxClhvPS/FQ4QhbLamA/uR4/OwyFosDN0TA0aQ
JBT1zj8f55Gq88xi1sApmSAn7Y+lhXulWywp+q+qVxyQyn1QC1320XB12qT3mB8F
odpDam/qMBC05nYR5a01cKvucGbpVPWu5JwDffdH3jRXsI1ah6ZbJDPL4sEltmu7
YMLjdHoVhJjlQNcoWwXXkjRVCSjiJwyJZyPGQzgXI+DgeZfsatxA4xhhDxjd05+W
zKG3qClQUbCd7yQr0AA7TTSAnmn3ek6u790OcG+mnXDcdkC7hPIefjkf8HtADKR9
wTJnLJ7Kt4WZ3mLNwRfWE3jIwLwjDF5ExTI0fr+EHae5oOyRoj9W+mcybFXl3rio
dAJX9UGtWNNVM5pBfFOvPVdi06aH3fV8W1JvjETJwGW9yEKG6xMN3G/oMwuYmD3g
QUG/TDbdYVh9RcuXjmIVtgrK2YAC7yGOMUbl+6oaVwMDXsQdwhvffn57vu7VfdPY
+Noijboq6NJjPfuc8dKnIZj84GsXZhbyThUi/jdT3qwv9B/qILZYCgymiWzmPf6W
Ed5mbo3CB3KfXYIy3zaakcDgqKgfSmNm57mRKbHXc1doVhkYI/PDN9RfkDe81y78
6r0ukGI42hnRT8N59QwjAHQRDYjZMI2PWmb+uV/XVyjJo44GjoSHJrq41oKk2MVb
ChNra+3zKCV3l7O4oNzvrWWFMCSaujRYmz3It+PgozLwOGxQoF/u0MBDTVamzV8n
04qButOZ1Fa4lIOrtpcHaViu5RpdQX0DOcGXRUCTB0x/VFGRPovAbZJzUHUgb/oF
hQwdwtF8G+UGofkAPHNa+HcDetWtt/yqdcn3Z7Fl8k/FB5mDoaDYSxFROCW80jiG
wC9O8uPElLhv8GL03nH+9hebQ6dONDGFV/esS5xhaHz//cgs/X8JDHWTiY2sXOdt
1Q6s9p6OBV7nNCPVsiC007OJRI+RHz4EfHJVjH3hjJIOQZEPKxOKUgCL1luTKhaR
h27wLtcV0L6zrMDEEiaxyHduiYLVDUId19sNbjSLg4G1gJZJlcuxbZ0AqkGP8uDk
shF0aqTqQvpkXS5OBL54R+ykMcLi4h7KGOtTtGNtTL/CR7x7pjS47EtAD7xzBO5l
ukDNHaPO3FQ9aFtrnV9o3warPDwTdv9+19K6DcaUqGHgwK85TmJ/Xl3RZbzRIft3
ehelTghZYqUpzNXoz2nlfznl8VbNKj19JvWskX82mOejiSMMelUP0NRUaK5ZdmOv
p+ncrck3z/CEnRxeq2J1o+yFj3jIfy6A9xP37lh/3YhbZRYbEc3EyuKTMTc00CBh
Pbl/maPU3g+IJoMfs3UHOxMivrbGjatcIwt7+KpRak1eApUAWqgpiO8kiivpjMaW
JYKgmn9xOTvkDM2lQzHf2LtgPQ/CnwtdGTdKm75jxA3CU/55syWacJhpfgnm3hhV
19oywog4FYt3ADbU74DAga/evU+f9sT/D19kbJtXAgk9pPhEZ/So8RVkimgHGNIe
+Bt+aIcBWS1BwQEZd1uBcfsV7UfXyEGwk8xSCY4neB8V5avv12pYrYUqsTmsaWKx
KPjCoGvkrx8aWtv9PSYmtt7wtVG9wGZE3rjpC1stdFsh0d4lr11EzC66Q54wOyQY
kIMUR20Kf3qMJpsACGHnUhTGI97YSQ+3gX59Mhjk8LbKG8eDOOww89T7ikkWFYGA
HkE/JTN1HYmzu0Aj7apbXx7xWXo5W7Q/K0zi62rJl/jnBWs34AX5944TneBtbvZx
iJcJT22akeWI7NAbtffoY2lApIp/wd+f8JhtMyWwlLQfIC7AkmPz9IgSDDC9kaI2
JBmDTRb+q6WEt7RF+CunXKi65QvoB0hauqCx0ffXdjlzTdu8pWOdQvq19SIxcOq2
MKTeIIsdphiBqZa+waSvMzNiLG0kcy22eQIs0BC4xWZsERMDse+Kt7aS4zWDLDY+
2vbd3V+GBkKtLP0KFQdnlMkzTmJf8CkBbs1i3iIf9huMk74UHe5lB4KX8VxjYBc7
9YvAcgr//P/CFWf2FfuclwRTg+RwC/pw0DC8xy69FS7r3vtzK7Jf2yVfFnHTRsuW
Y7ir2MRaeKbzobIGFXt+H8D6jtttkqLx4kxxGtSRT1HleX875+X24a7vgsDjzjm1
p+FGlCLhoFiiNH6iwaPt4og1nZuWInyh2lDWwcgpbUu4Kq4wnlxGH86bOFKMTjD1
ci3C01idBB6EGhb3Y4cA/Xoj4cft2sBqgLknstRW9dArKE6vyD+a/lFLmivbTE7o
2WTub03W9GAtTJK0OHP1DBt/5IcB0OyXk2WiQAkrTv74r/Gd5NExx8X6w/KnMRNK
3kQoLWwxMtclM7osov5c1iPHE/sz+BMFqDjQrqb6W8oBUloI+zbMQ55S/B+qbZA8
X4lF3XzeK3VjigRJIbz43TQwfA8xy0k2oL5FFFeETxB/24AJpPmh9bH39sEQPPxt
fCu8hSZHMVNy2qAZXfQzIVV2NdrwSHsB6OPwFul2nZTYO0TpUrfq0PLMJuNAtOCe
O6aEfD77ONhP618J9nEhm/NrvyuBLIi5b0eizPtELzGxxFGXKCR+3E0Vj66orEVv
TouG2QoFFkT9UWP5efyISysExxcanzTz0/Psekhy9gx0ROYwTRM1VEPd//aLrxS4
s15c1y9SoxyXEwT4v0Ap4gAnqPFk3zksjjUlaPyMmPMpsJwtgsSsa5veTraqhRZV
MJVtcbMwcXLaMCTFfMxc1xvN1UftNonipi5jZWl+HrnxR8I8+2sUseAj43nPaAG/
103rGRb+bmKZUCYPVvnjrkblzKql84w1jztJoFFCMd6am7V1wwNhsD8ZAbLysF6f
pNligVmrb/E6n6JKeZCqhYfSmkgcMVTKp8WC8M5xkRGqk6IZOxMjK/b2p70iPwed
hHEEzPdRoWNi16QmaSGB2uojP91V6/LgVmc/XXGvxLDXTRsXn1yfGeMmunkC8WOt
xDqU6cgvSzVbOUFQTpYTdJCnWDITwqyNZBcjH9QeW15kMMPWAUviXzBzAJPbVNbu
JIGvGQG+DUzGuLoHTKDSX7vtUiJdKV7mV16KPLWsOb2v5zAwlmw3dNstbAVAqoG8
Vwe2aj4kzHwdlVwZxREWJBs2vh56luq3t766PgtgYWnZ/pgV18R5CdVXop9CL9xu
yawA3d8/tRP/QGxKBm5odsVZBCiL6hGKKpinxdTu0jJz+29uyzbUIT1lqI8vCdQ9
0QUipCAG/WuxXP53SdbEn8qs+HyXarBJadEn+QLVSGblZtQypmaUPqGX0/+Zmpqu
f526gL/dQa9k5I1Ir7Oiv0ptu9FQBi1z+Sgv9I7XReqnI/jzsqE+xmhYX65zlH67
O11EmgAS5+wyKwXWbyoHQWPCYu5mn0Rc5pAgkWtVA9j+3eKc+SQkgUPY6r8tau56
laiKyMM+UzjcyLAt5gbLnzgNzeYodJm4AH3LkgIAT4Jm0iCxbFiauqlh4urFSeFp
FOFDzkq8GMB2JWuGbmc8jaJpJqMBlX9xbY7Ipb3+ZuDj378K7HUkb3pqZSNlj7Bm
N3Yc7kH2YuzkQ0OqpqX4bcvGLd7lT0VuYWT39MCize9WaYlcGiloDlR4d8BKGt+l
p7DrLPYEPjpvx85n4g1e537xvV0tJd9yivEQyZGjLBrn3slNJghMvumvhs5z9LGM
psT68giQ9wKNCagwsa76jPqtiUQz0W8P6RO5liKeoyY7A5HssyPAKe+PxucubvjB
NtvfJhp7o+umrt+Bu0uuF4ePRwdane7ziL8fhXd3V6mJ51aH3c9Pz+ybtfXQrH2l
GepXFCSVm1X8MeM3iy2PK6UZ2A7AYRDXd6CviuCmcGuZXYo0WuDnM488ymQs46Eu
bl0Mn/B2w/vieCe5EQUydnti1AnRKfRz04gXg1ArY6QRDWv63scOdYCTbekbHc0f
OCPYB9GUOhnEJIslntnqAQoZuznvB6mXwoq1uZl9vSsidd8CES0ILPloayqZnGL3
BxGrn/fYLu3+n6FvBfyJ/D54fS6GS+XIRiGjI/wH3FE7poC0XBBcsk7PVB6O8fgl
hgAAAoiYVnJtU7nZYmkl6FpX6r/55SSSXH/PzG4b7KS4q0sKHP3ctQw/0ODnRN0L
TA5VXToU4kNZkvKNV6+b1r9NNYGdSumBsVjiElTM/Z5rsvkz6KFies6fNA4IMwVv
IEPPdmBDQ8N8UeTkcKA/xU9sA2uSfiG+Hcm/ZqqNChWncameQALWD34RHt3bBeHp
34gudZWZQabOlaby0UlnemjFlKHCMvfeRpp78yjjgr9RZ+8wPVS1n+mH7R4JGrqZ
3nFMUvmKNF+YZqjhk5vlS8DifLJi1iTrQAR7udAyBtH76oR6JXyarvz9o/YD96Ld
1zrJlexSEKsDrCEw+vKUMmGfVmb2eWpN2JuuyDTitJiO6NxherOHYB7/eLobk0c3
5v+mKTlERjr5IbjHVCbbmGIrLtwyVJv04DA8PvX4kdYsLdiw3NGIXi3np2HEUaqm
hC6X6CTgstZhjNBzMgP4mvmbhXBdM+9cauT94wnD4QOgQ68kgi+roiy+NC09h2MF
knKNFnndOXIqyLoBNiORvBmZu/yGzDHRGLIic4OrWD7/OKd1cygeLH10NemF+uzK
eMldQWTlCkW/V7C62YyvnoIUhtffX7VobFRqyNjzLJIC49HDASVDQx/r+QQN4ouC
PAEPsugKMiwYuobAu9U1SU3bMpSX3Sf7TFpB+ZCig8W4Og1HmEfbwZJZMnqKOS0o
tfxFvhkY3lwlbIq64gCOVNgAawe3pln/lhfetEB+fqq0Cr1xenieURM29rXs7nV2
iTyVivDfOph1dnPEP0BJbbLsafF7nfew0Hf0ab9WvrMshy9aQj/qLv7wzxrgjwEw
B/tzhvtHIFCpF4QXrnGSa6jZrHXcAc66Q8fCVqmn+TY+9oCyDTz/GuHCqhdmSBOX
5wCXYSG+i5tYxb7V8NyCZTztBPNPLngaiX6AzZHf3B5/d3fscGWyPgIXnFe5Vdq+
Lj+K3lm1q2MQeMbe3Bwur6vVwUQ7mFGDRiAU62LL8d5JGCM3W566+/sb9wTvo88r
FzlnfQaWh1O+QtYMg/g1KgkLstCUdR2zD+Bz5Ts88hc5rZv91fg4F+nQKz67mhHY
J+Uskup2066xgvOIyiE3ocWMS7EA+hUNKtdw/129zG4DM1rMr+ZTZRuDhRha26tX
CRuMoJ6nb9F5IRUPvg+2YpK0YajZR6jfkAfMfZBWF1y55rpxUGgMRzoDatkJf3bC
3pmg0lCoafZ3lJz3s0MQWflHp6P0qdU1/vt/gFUYmsLb0jhmbgXtPgM8rvbYRZvX
tk+6EoFM0Q7aY7kawCahN2H8o26+HobKxHFRkAvmU/FGa7vrOP1e/RaEwQwyI4AI
EivP8PZtCX1GKq6md60jsiaWGbKuCaKhUKJMlDh6n8RwjQyTh3Uw/UJtV4+wsv5/
304wSXGgzS2a28Bt5kYN/csrDkTwony/QwadmRETlLqDwc0fjW9DA9cN7mAsx4nX
LSgs3KGRC266xI9i9A6qr0yH1iEcIl4wMzIZWJlc5g6IsZePaqXYunh5dFt8fi84
HodaK9iGZO1SJ8kTidAyme9SuFRyv5Kp13xpOZHNAtigy4UX5tRsC/G2teTpb0/P
/LOLfvpriZ9sY9AjbgNT3tzPcgOzgDhvmdqxxuTVtX2Uc9dnRmc+OwMHPOpFmRi3
hBGGL2gcUh+w+pSdDEslUG0PGSuGWlvw4RWIh4ZJOpj8LYMb6DxEvrMYI+ltn3vp
+A6+Xeo0U8ukBbtC9/KRuE3AkUAEj99KRnr2AKZS32+n9cIhFRM9pkffR7UcVbv7
lzRI6/GPDBBNrN5Daz1cR4z5mA6dpIO8SJi96reYKgkr0OweehqdDZUOX2MnqAVy
7mm0La+WWU0O1taPvvN5ByWlEIzp6cD/idn0nwlJ/bBngC2FnMqFEUWg0RmJKXik
WBf3lU8BlG5ialoMQfKUK6dU/VPkSUJldZZ14Q6PYoSY1Iv5ZenN5JfIPRw6f+UY
Wn+V1EtrZPyuJrYMJQPM+RQOroppeWBiN8ElqmCDlTFse4b1AeyCTcihoEzhmVqe
ouFOJts2OjMT3Vt2Hpjqw69gs8MPOLohb82viPqR+S87H4DAsh73JR0usAR7xtUz
Yhuarto+r3GhASA76op5eLlQ9ZEZ7KaSnMMeByQpT/46FVfodECGxMpw/bkR9lUm
dEt2OU6pQQbvaVFIjlR6ibjtMCLuO9srsghircv53dEB5uOJMkAoFgHWO0R898K2
cTU1zxQswVAdfWHkznLSksPlJ1SsfFnQBgKomLGNzOGokF2W1vvOMy9ml9PDuRel
bm45BjdBbA8ManDPfCcNs4xkoHBt2XMlpQk5sGmfojiKgkDc0U7HeUnfHKOBO7/d
f2mV/3NON36y+0yOSNDYxiFj1tfNsXZ9UgPrgkks5M3TLbKjoHqA1nL8rplN9nxE
h1+MoNx0o3L6mStle4RTYXFZdZRUKFnv2g+cm7R+chOeleWA4q5spJyG1h0955Ek
+L/f1pDnuQR9+dj8P70HI7LlAmMshdZeKKt/Fuu/jM+sTrpuLBzAGuZg4wE9GxG6
1zZOjVOX2CiMyZ8PbFxz/fzc1NueUdr/ot0uq/l/Ggu/8/saQWbs0CoaI0So7PtH
/Gg/8Vu08sVIdADmM6dVQSTHYC2b1SWjOwMipk5AwW0Nb/OrHKn85hbTJeSMJF9j
pe2nb458X8BgVODtO4PS4xCqmVInavZmuu7FpjaofJnUo4SuLaS1BftXUoOEcjXe
D+42Ciyinv00uIHflUW0H3iyFm7ZruLH6Rp6VjkS/XgnKPrM+sCEC/cAPFfyv7/4
k5a7+ybZ1zqRzG5smKHWj94KRigbSDOK/8hYcVgDwhInzgPIt6TWTvfiQ3Ih3rO5
DR/W0S05HiO8Mo2JtKv2KJsJm/NYeHm7GUddYfeJ0cRWUGNWTadJSGqEDAxImNaX
DBGL4aiPj8HMd3I0U6tMi45738tjbw34D7P59s7E9ug20O/zwS3Va8vKpnoi1tUt
5rY0A7vFVm7GGsjeKr/4ReP80vwUWZGqYVpkSQ6sUMv2MXcuU68q9z4h43FInwuT
aCF1SoHUz5fqSz5wdi2PLBitOmoIOOPDDN3sZVffWEdANUtANIaGrx7IBcrqKoV2
Th3nwvWsGl76/ANlm1yrBqHzOA6yMuyKeFsruRgXxZCvSD181jAY2BhcQFd3/6YV
6pzr2bHahv6yzdEVicxNoZw1mSd8dA6MsuKMBSEGlMqtiYuRkdjuPuGsMrVOWXMX
TjYFgyHouRbIRtSbeu59A6aAxYF5uph2NueTORVwzMu0drKEUY6SRibXUxeIJfoh
QmJjAatqgD8WJPMvBvMVIaVMRkQyp4cUOPFZoT5trwXAUohy0fW1rqfYadJct+gT
RAKOfM+kIO9UsWLy/gyMzdOEUPXvc2pNThbHt0XlLyDTPBJbiU7EIPOLdFSVYTw2
Yybtmn4PTA2a2Uf6lHntYkxNmyMZZKsep8AqvAZL/FJf4A94jF17BDFWDjq2iHXk
mOt7oq4ub+XLybQpVXwhNuj6jlnP5kx5BrO4Sl0zLnEwJQlr4ujm0u9fyuyC6s+0
TNls3CHQXPcBa2wybpObTkus1ajMyT/hnJiPhUB+BCJQwqsgoJSmszEyKqlW2I9e
2fXJX3aAgayJsD3KtlCS8MHe/iGOz7N3P2xTRfu5WvVaBiOnJNJbWp3OcD9hDcKm
lUQpvnG/lYsDcArvLFZ9tezZlxGKSA9w6SU/RYOewbxJflF+JGy+Pa4AKxupVjlJ
5YMCka57XmdzUaNuX7Q66sIkbmEhqpd0x5+ceNPN3yMy30y6CuLPs+4YYdyEZ3wo
RUjlOlcbSD59oTC4ee1gSa/HHRJgu4jSdlVZ6x+vHZKjWL10rkIw6xbsaQyosU0N
sHcO8wxtdV6eaDQMZMKWCZZBm3vA4ugFFIKnOZiy6gOtJ6lqtVN6ZqJE38bp2dz/
Oh10MZYuSPQULUgWbB+9iSI2MxOR0vZBt07ANOR5iJy04c4Fy5ywXcWU3JWATQUS
pIJqanzP76nSPHBh//q/aD/P8+DSFFF49Bw9z5RGxfbb85HFgLtmZ00jKZ3phifR
t1OPUhXPonAU6U3NEcEWrvd7fknEO3KoZF00zgcviqDRlCGMqbVOHnG7lhMB4GF6
N9xV9SCAp41ZUXbW+IMo6vV/ikPFobKbh5UAtHlZEgAFbEqIgmmKN4m+EC9eMzYl
flqJiEyBt+tA9spbOMl9zTwo0y8JFAz/lJh20JH/wM2mK+g3ZcivBWQhIayWEzkm
WO+nV8okoeT4Al5sYJFky7A+suBaI8ek4t/JfVX8s+gJhGDmy6dCnKR84VU58UAj
PZZVEWXAxpoHsvngV2FJRMGMrK8QKEd8wPzR35Wjz18i0YmuLbla6BHliSr443DD
D9rVnVlTqNj/PpLE2Rd2CLpMgzGXWmZSKkZ/GO/VrhNFbuFx7mfFkpNwanZqGNDp
wq57od1Vk6wL855MnQLqhQOAskp9pwzZlJsid8T0g4ReQlvMzOis96WhFImRZqkZ
CaJRKUlVvnHoLq/6xaYutt7Ir8o7pPkhXSbd/ylKypR7nm7oeTqnD/FmJBoKCHq+
0/f9i0HDuA4rEprascboVhFM7GSWlM1y7cs6YW+zGS7GpGhgOvH1cbMq6WZmRA9a
wbo5ZCfWLtENwy4GvBg8Z3hujN86sKtN4yd8bmm8kvgRVwrWPBOey7q6JRqOMXKd
s66U/S6PAgbf8OFgmMGMtDx98enbMBjVuX239Qe5m+5l+69w+qGEQOEAdCYQ0Z/q
KbBBCXjRuhPS8C7CkdHzgZvKu6/hyvIjrSUzsvvKw9nUNoPdPE7HsH3O2rswsNBw
Lcc5Uc1XmmLL9tdkT2oV0qzNvxgfovZ1KQTzxGDHoEBQnKK7Bl4yTxTTAORGsrI0
1RDUuPiyt+fApmNbsSCYbEDdq0ZX5Ge2gyFRQqIVAfUbJwNn9YOnrGVMTGc9005J
LHVMGyjODA3XpJQFtezhFAF2k7LsrLXk0c/aCIXv0x8L+cOgxvD4/JUhJRP53smy
HRHk1j0ksWHJU7hOx+cPTnip5ldG1f1uUPano4Udf+YVjQ7icZTBifEGBJu7nIiZ
0zkMUJQEz29YTROGholkqQTKudxlY89tUaqiTmtseb4w9uGxmX9n5NzIVicqkBvt
fSotzJ04vyLx/miHdey7XYjJrh7zs1Gqa5pkyT0QTVgDUg8ISfT/yPFPKRFxomZu
D26f1QqBTD+WYiTRQZqRprPzNa+V64CdIntz2x9oPqvN6Hy3CDbL6l4euL68MmSk
NA0WCMN5JdSR2Az25KmGk3O0ZoREPdiyE7yoi2HvRhHkDnpY2H48aNXdmkBrXQfO
tnji0oBtAPwJC7nIXVBG+8EzX0AfSLOnk/R0BQ0/hzdSSC66/wNwIfTcLiYzxjI2
c6Kq2Xo1iyIhpzm/0clkZ3itjL/HJ8++CeRmYD7MF29Z6YOGNCo5cu6IXXol9y1S
3ZMGNwln1YPPM/AJMtLICLY0fwnEKglWZ9gS5qgm/5J19zRa/qE2dTvfU7OKTJSe
69UqRALNk8NY5fPUYHYugS+epEl7TdebNEG4XXNvCudJ3/eUvzElxGhSrTvfoQWG
gJSN0zXV3ME3jGgWv0XrxkDI9JXFL//V1pX/57fyKlAWD0B+5GjQgJpO9SbTRUQL
3yqwSBUaJulNpUFDlqs8R1M4xdV3g8vAT5JN2mMNH6pyENLgZ7sGVtCVud/RTMpl
mUuB/zTkk3vvls3u1PUlAtQu/x7P02NfIf5rHmMW/e7/NNjv4x+5os3VN/LN+sgD
bVbdN3wx9wKoXEJgMu/+KG2Zvweb7vdNEGemWMotaXtEcI3SLMjkLMMUrExEjVe3
eSHcfmEu7KywnwqHju4Pj3hKDAlZGvQE0MPL5QwzkDapfRDJKGyJWigLbGluWEA5
XzdY29D4V5mdNPeBuwdNESsV7NPNbSB2CBbdk5B2EjntwSVv9BR8OsoZ3ZxT04mA
AZ96oiQQXVLVQweff9kimIk69/FtxhF6Z79elwmm/WyHH82569ffBZVU1scZpLGM
Zlv/VfDnx7+R0pTBJQwjny8o/aOFM3rXgLTzeBhStdz7vfGvelNSfjZ59GS+qLZr
DGjbGV3G7VRv0b/rO/hmskZP8HHeqAzVDoJbZoewdZ5/ECqPxm0IAPRolY7EzjvB
nyUmZl6anbJ0qAIZ+/sR0NnpexTnlGVsJT8MqGVgN3ke2se4GAmrgFZ4Tn35+iuz
JzzKUPUQ3tvVlFvJuNYv7dDWKnLe88M0ZZMw7Ffb/VD0ayRsPJukuzXHEQY5bsxn
oEUY/busyp8GgSnpBRMk2BbEta2YNYOm+FggPmfIndO1yNfN1ytEqOmbUdtHoaVl
2Zr4yF5/0//AAWWPCxCpVmPj/B85ZNGtzxAQRhP2bAleXbng8EKoPVSa0v32DwoK
qVbwPiQXPGgJk5L+eZ7QjE8rTL7cAcT8FRuNLgd19M73F+qvyYbPpM5VUMsQKSBt
heKRghuNYvZdpMH3CtZvRfW7WYHJ4P0OmuI4bgr7kkRDJUXQ4P9LcluRmSV7qDH9
ggs9OjZa6DxPYoJF41KrIfUgY1hs+gtktGU1Bgm4+gMr7mHE4Y2SzVAg/7h7YA/Y
m+QGK7LbhIp5H8KxdJPLThPE0ks/ufnrzcIf5SZMqVIdd00DvnvYhNAlrArp7LEg
iuqymR6T9Wp5ZmGgjLFdH/yJK7KJ9sx38wV/+PZXNIQMOey0OloMzeUivc5dIGvu
eGGDYjrNSvGSslAJXpUaJRl0FBJz+mQMCwoO7QsS+3u1/3moldLi7U7ItgvUrB8O
BGICPSl/PfzaQ+aKOLl4d4+8AHVVBWILA7sPZSKnJxDrAuNVRl1KQqxCJxDUf1rK
1cn4a/tYLZ5x43PixPCI5gxNgO78n/tF14opjwK14S6ylYBfhwtvhCmxBvipkVEK
VFEdX6IO+bUAW2Yav1UaFyV/j96IXWIRI1hsnKns8rqpCbBW+6GuwCRBO4Vw+L45
LVodQw3FQ40Iu8PM3FS2x894xcd8vodNpC0ofHOc+KbWk6qqduKzZUQm7NJyyzHh
HkzXDUpjaBdfc+6DESLs/a9wv7EphVfCbUweNKb4y+ZzaEkcSN/gbJRUjYqvjqQF
VPLnJvb/DdYOPlcPxUBPYaABjHwNM+3LQe3hdK/jXQd/Cksp6kdpbP/8VIQUDneL
Fq4JNDp/r0zONL9COMRg+Cqv9c+nv+itQi0QxZgfcs7j0oFiAuMy0W8xcntTf8kc
J+I5805SXXtGGlkt1YWskoeCdXvFun7gbMfZNM+qK8FxewCzAuYmvNI/htdFbjZo
nLT4o62v9z9MvI10qtQm3dfu5O5wnqLNZtlXo2GmBFTisi+4+SlGv0na7kVxDHe6
UkntHF+/qUwKAkDGYgyrIDVwbt8Ddm/7z2AMVyRFIearTIDoshBTFttWufTnlKEu
Al5pKoV83lbw4gx4QELY9IO0qPjaEucLcyOv0DzTYOUwYU5pzSThp/IiVFSYrLls
r/8lbdH0t0nItggiT4XoBhBvhEAIyo4uW13ZlOu/OStzPRuB5zD8YmlpbFruqDM0
p+uEJbJvsv74jqZBnXe8qD7sNUOLs2PvS12/KiWnWi5SwRN8NUwUnYxgPm5tan8b
+VOdZoRe1HmjK5sgyl0e08IPQc1eObOUYZaZv+VE2bi0sYe8/6dsKFL5sbhj4rtt
Wyc8IcG4vn84quLi251CSokBO1yniVrta1hkz2NFBguvcMHwIqeha5qPgw6QMDjR
5yHiKQJsUnj0y/8a+SgrArXKyipcuRamu2dzRAmUoo2dHlqDWEDLh6SAsAx3hb2r
Y3BUtoy1FIVepaw1LNaxQmho2F/K/76BIIOvF1Ld06G5GMwaxAWbESedWfRs1i9h
IreVeis0zCKOOyCcIBR9rHV6IQKQLDofgZFiJqQhdgBG2RpeXjpINEU1UlCzMLtF
Bdz61l4fK35n6M56Rz4r8YRz6O7O7+PtMw+fc9xomZ5XF+vsDFYn9fzsc7ehRuF0
QSWaTK+GwOGiqnV33X+Srg+DOQ155vtN6zMT1b1mNQ8LdpNK9SXoGter6h+KTkpm
VftAH+CJo9JKzfsABNKoTc2ereewGYnGlHeAGbfKncUtod0XJjUcycs/faA4hYL0
/EWyRVlMjJBWbIrENoOLW6h3/smxrkKMjdSfL/TziTG+8XvtuzDwBBU6s9vBXGET
PbAIs6mbR7UN8hCkMy3A130QgCihtAQ79YOh6NKp84VM11izi2u8PhK5jrEUKTSa
PuVQTaOvouuHf3kytEB2pGno2/zJv05yYvpQ3U4afWPwz+KBhFpg1hszY3kF2acR
NYocoZDuvhjU28JQbMRzSpv+V0yNiDqTUZEDmR/kiD7tdUa49oBVrG1jNk1Ru58N
Xldds7m2HEPs2HGaAzL029lZCwwVvggW6knid7S3Fo7odvPjeu+0db/2Pi+eA1kB
Lx0jifNGpRwX4oUxHd7KCQohze+Eeh9Mv72dYXP5yxvh38Zha8iG4J0L35HL5wzV
j7xu+A6l9sYHaobNh2xHX9NDwhn3bEKnO8cXKlBCYhmv2gb1W+3r5gbLTbeP5oAw
IE1sUWYMNNJREYAAcn2xpI6YFJvKgovFQQqLi8mJ2a2AuMOzryf1gwauLC08CZiD
l4NDMEX4lyj1ymtKqvaXC3wYhaFR1QW+jd0c5eAGIDOxpnBUvi1uGL0lKvP9asIp
DBftpvy7IS+v+1SYNjt/krBWY0+iU/P4JaWiwQhwVhqtuBp50KeRjZqY6YkOi3YL
jzJwU8kwbtQeMRX9OaOb1Hqw7rsyrBV6QM399bd5K+hjFkQF8BIaXShmW5ahd7i6
/5pJ0pROKjrnoUL0Rfl0AYyAD4uAE2oWgjKOYgHMF07QiG62OAZ6D+UndBVIdMaE
hxIaxFXXVRK2OjMKTHvSFSGJlr8wMGqNKtg79AmT/sq/ekcmZiVQvGGm/yykUIR4
6m2lXNB30G+kOk6yNqPspOvaiYWX9buitPMrDPbYJ5BvjizWFvCY2UARWGb3GgLo
pGgmOCjsYYmmCaxObDkRDCd5ZyCSakzHfoShMQ+twJTb3yXFlkJf4jS5cuExqA12
/BXMF2hZ5P/PqDSYBgmYOSsUOgoH8cVRy4rX+t6angA04XMx8trCGWJu8j/iVZaZ
g/EMARGiq0lU/yLbiwpWkBdISAUT4bDBKrFsDaLxAfAhJMmudDFK5kfR/hBKlfXU
YZW+kgPIwZb7evCNrRJdHo4GoGt6N5GhA4ZcIiLEsgsC04mrsblwCoyIK4GfFYOj
Y8C5a1fasA09Jfn+6Li9dFZBfdnY6gIdoexn8HGVz72ii9ANQZZO147QjtzlD31A
ZkZfuQLnnchSm/bIAKHzMabmd0S4gl4tt1VFl7bZtxaniSbJ26FLGby6g6aTLfM+
ZdNcqGgydZDZycPohg4TKPejx09K3oezumDQ77cM7mZuq95HHNyO0kENtD2XotMk
5awQwRYxYh9mR+KOTgTz6qg6wMtjcrsWBSH5ilHpCFgFYCNj2VfEvP0IL/CMH/iC
hTHgAlmTUSezur4sUs3lmGg+3DcvY/o+t5MkkTdLcM+xW+Vakk9Ym1ONnqZCL/4W
VX/jDAOsIuOh8Z80gK0A4c8lnMYI/sTB91Nmsafx+ah88yo08gbi61TeMZRwawpu
en9FWrPl8uRHlPIceermYtRn0/gzCFc+oBQBF61hzrZN6nak+l1C4+T9iiltYvRx
GJxunf7Kx1rPCHPEd8VA0MTPVSJQFbr9gDKw129bURWGUuLv7lEuiOfw+4SM09aN
ELUyEiEPtRFTUOQNUq/YA8Lsh7RAClPuLH8TLmlBgmlzk04YaP9wY92g23Q58x07
eSH+9aRuD7wXEwI7tol1SVJib0V6MgtISJggpLBR/IgjmSC2bp7Xs8gHyURKx4Xs
HkmYDKoYXWwtl2+kY0pBlIXwh5HbtyFzN6Uc1e6GDSSZjY6TjC4RHmRnjWblZ8gA
mR6Qh5L4qxGkj+mpfTqv3DQpslQ46HvwzqSoRHy+gLW6sgTBDixwfzPsG/o0CfqJ
xBJQ/N3aTPOsGDf1NAakO22gYr7QM25g2tNgjMnODaVZ1RRzlYIqzktz7sQmu2tS
RmfacpvnUE8NtdvJlIQJhjq82BubA+HeVbiWi7y9kZvbtDJ+2OtVEzlb97T8HW4v
PbUs9CEp/1CRxLOzuP7gZNawM3HoM0fQxxrc0dc4CoJkjtO/y2VhWvOhAsfJsprR
r9MrDVB5dSzsWwjVoD0mMQE9avJGOmZumpJCKKwuMD4ScAOBdO6PHrbkRJ7/f6xF
9B145lvN7TtPl5lfC+njpVH9Pxrv4as/HWHeAroAey9isQzPtSsAWDVRnf85tMK1
edEB3Giqc85sYVC4E8chLurRa2ifTs/k6FO7pLtyo0SnJWx7zLaLES5iU4kXY+PZ
/PkRiThX/XsbDhznv4rEjlywO/8GjM4xC3ylNnPf3a00JIeXORYzGZjHyHCGGU/3
i3pCnk8k+C4V07pFO2ZihDyUctuFPqLv6uFg0Rk00sGMV38Cs50daq0x/i66XLs7
TcOu+BWfVtTmf6RNXr9Y0gyAw/CDqVcpBa8Lgv2pXHc361fs1R15trk6uzw21HBS
drRwCKl1Uc2qAvaAtFWkH8EtULCAgUnGzSvVytlvinm/TsRIuvc5ZCtlDCTV0L4g
Aa//eG3/FmASIEh0czCgd+MxcIYHLLg3/AeXToMIfMYQgsbHFsk8t0+fsT1gtyEK
oVKZ6rILKsa5w2KqySXs/N/cajJKePY3Nvjsn13om7c9xANUdGfvZsgUa01YL0Gq
6EPH/ZC2dFB6sjD8NgY1uehsv67SAzN9S5+kpjMjlXXNdKdqzMspzXHCq/8VJsU3
Vv7h1WoS/V32kQuBtwpAvh+ZxRyQZKXQd+b5wgI0eUC+6xNOTDC/P7g5WsqWYiPr
HUyz4pOF710jSoJIaHdpUXqYECKUbZ5/Atb0pkLyAc9QgKH2x0nU3sWTJIq3tw7V
s2BEfOqgERI1x+mDvDaHxy/RVjn1zlfs62HCOtHclrDkem3nWmfhKQ+ZTh5fFaoa
3cnKyDpyVE28U4z2vx6Ib+rGVjUEtzw6nrIbbvTR+IQ0LolrEIrfBLF3mWMG2fPj
BjhohLndliGjqkCOZ4UseQCoBEzRgGeWkfxSIM6HMM2/N3NpO0HVxCpf2DIxKQ7m
gx/jYm6/iEXsM43QH2M9LohU7TbC7fZBOuXlgJfUKLR0RSINY74c+UcrXa5icsJq
cZvPqUn2UGk7zaLgsvWjTuw9FLtQILDM16mmX76nm/P0FYrN3NVgwr8NkUzzQMnt
SuPu0b5YJmUwYy4hih7ixKqVpY4xRxWXQrdybxVmtD/VbAIaVOtB8kmzOiGJGWen
oxV97V3vu3hWXNttrTus8qZJrzch8w4BODkI8P/i/Y2R2h5EIlqGPPBhJsoQtXuF
Vjejj7WgOM65wgyRv6jUXows/GCZYITEKXHZlvWDm2nGGtCQ31NQux0fzkiBoJLh
Z/upa/2exWcHKPhqu5hsL4wUqovwmgD1SlVUEYDrOlu/7yazkc6o6ssxHzHhnQ6m
FYq9zvO52G0F/v81BZ+RXb9KyZsXBLrl0/LUpKfgKq1aXgCxD/M2RRm657p9aGIU
7xS6fTdh+Gg2TBvIGZu2JY7hzixxF32NLjXGAFLCDu7ChjDUX/zKNk1wTmTBNdlx
WZy30hZwCcFU7m1hGWz1bDr7ITBfZ0MRVNgfFUTpOAK6UWhUWBInoA2mt9gdb+fS
Qb13E+vcrN+M59/pEcluvaQOB+L98LdsGatNaqaWdq67ZsvTilNzs2tuxFaXHzh1
QuJNJi5DWSqQ0+mgL3f6IXNX5DqUJ6kSXOCPt8FivIUM/vPPwYP9qNL07mREdAXc
aZOut4RWGzhDUxgG6FqHyLLAeQAj6yl+vRx9h3h/CBtMqaEfU0hQ8s/RnGOF23Ct
kD0ofzdb/oPdhA4gL/srv/3c/RwCacYfQlx5QEkcnzUAWeIr95lHhHFQ6sAdEae2
M6Mv3SsRsYNYZ0+qnEk4U616phzcgf+2vDvYr0eyP+soxFBZi8MmXEkU1zbVo8pV
AnWfsRXOsWnbVFthhV2mFl0VnB0PsDNcjkQc2QZnXEaK+HkWBT1k2ve208NqDIpj
I4tMNMJ3p7y3buwtPFSa2SvClx8crxxQ0Em1N2WNPOGVLDz1L3Tkax+l6bzwyONe
tUdETtgrrXBLFhA5UZn0eShn56e/34MELfHDCoG5s8R5RuyiNQ7PDuXsgtdGKwUS
Ysi0e8lYS07HmOommTQ027LwmOub5/iEYnv5uE7ar0SY5y80ZUGfK7RSqgkuNySx
zWWT6qn/J0kZw4xCREyBQylDzsPSETDAEO4D5qtnMTLyhVXzxKpteYjwrcr6CvfD
KqXMstzmL03s1rRAM+/Mlt1DLOkbSKlpvulcY7yhEk+HS9A+1daPl2br0hhXHPFO
eWuBcdVUvv38JnVwJbnDaExk5BQUS1doqxf8KNZkJwavhqtK0Br5PCuVmV+8ypek
FOkfvlRN5Hu+UNDPHFJQ8jcdHTVN5NcePaCis/6zG0WAOzs/TxL8rQJMeJuPFrku
eRhEjwRARnFCOTijDxnNhQWBCvM0vFtPYajikyNe3mks0mIPqju9upYwY6qhk/Kf
djLhZpqFbkCZDFc0F7Vcj+Hg8gnTM6imPoPjpyI6STqQni4Oi+tKYSfz1yxFc2vh
E5HHUc8GYij7BkOJOnjBRFPbARw+ePL2iN3P5sbcZ+bXqj8yaifoE+tX2MMI832K
5rZRsSRp+re6MSvqOWPwSCUlyJ9SVuHuWENJ6i2FHcylPhgLotrPKaWvDpoqvLcC
jkjUeEjCG1L/giDlr+B3f2NMExjaRxM26gZpfg10ATrCIuXvzLdr7fvK8OjcGvAN
Rv8FTWD+BJ5pKNnl96mAmQ2tRjiVoTdE3f2rWf3AXNpIgJ2Nt+p5r5E1vqLupnqV
u8jVsdogX8CijPwSgVTVclC15S3r/DQuEccXsvR3HE6jXsxYznppyA+ZtRoiGmw6
X9TxhajGGQgtrmwPC+5P0jLRrKHO9W96SNcw6vYB5rCXcUSkP04dRNfy86u51o3s
S62isQcjMhTeSPPU9pL+5OkRzzTdEWKIcAbrwRlSVzDgDiDforJVUEiNXjlEEikx
WBoaMUqovEHls6nW/Y8hxCiphoCm6u+O0X69P0FTITPziwuyUf1pxoz6Aicg75XD
j1Zd9TeGr+Cm+cbvUced67tUrcUQzW6pm3XBW1Sng43FuKlJ4mtBMKndFG+U3Prc
GCu1bPyYRXpAdmw7ckGLpiYVEQmbYwhqfbEMnXL2VLFwgKaOnu8oVgrpd+0lquVn
EKvKJQ3Vd9Jj5mDA1ReSDR6kvWzhs+565jdcgXz+1lgUAhe/G4CrYjy0xHAEtEF6
YededxRqvp2pFsoWBkaZHC8kr51dZsU/276sTWfGulR1iHDZmzrUIsbUoQM1NTAs
Wf7VnPzbWp4w5q9pLHsY3KnRXjHkPu/uof/sjq7O/hqCNDfRIv40ZtPTRAmU20vo
knlFF70uAXDCfQvn9Zb2hH819aHvpps+1typT3tg7j89rKh+7pURCOKxO9bNUakD
Ce+/Wq9WZ9L+JLQH8SqQvp5voIRTK2u0NgSZI93mZvWHgOf/Q0dzCjyt3EbRS4mw
EZq5u/bISsgAiJzPlJnKwwbT5wgrMMpuVhZ5/Np4HFKe+2ksqFIKqLwcQ886Ol9Y
0+ZCe/kYP84NHzYh0qVMHbfRgp+VIQriGyV6m0NHPDlouk1J04AxWrzrQx8vXFza
1eMQoNOqT3gschEy+7KE8XKvX4xvHC8si8o4lcKXK5bjkPaHRy1wIvL8Ajn8FYe+
kd4jjLt5Urk4e8zx7jUp/lBSuvLn6rfbQHFLpbDoD63dP5EnLqtU7I2hgEcBoo/i
duR05SsriPz4nY1WAg1znOWFQDpLYrVbRDh2VapVw8pVtSRQgBCMIA69N1LJNEHe
K2huGGBQ+g9y2i6oX8EF56SyDKGZiXpdSaaPLqoPNbnocYPjaf+Xl97vXVDF1e/o
F5CbgA6+8CrDGbtrislZfhiFQHGY5Y7B8KxpCjINSXPGpwDsZPNHJq7EMkqK1B6C
tV2OIydRInAXwi0gv2WhtEsL8UB7YwyZOxZe2ocB2FU4Hewr0YCX3+SFQ7w96H8c
x1xztYPcPLCIvIoN2gIy2Ny7WeISDrvstZHCXXSNTdq79vQZfJ7FHrRe9wesKxoR
FObUMDnYug8Q76MAFxOhbL4V+Gdp5L2ySy4sW5xrAQ5TsYALtpWpi5Jfz76ywnCV
JkjJ/ymHGhpk2s/BmcNtEwkfPdk2sDWAAnmV+CDgW3wRxsFSZA4NCEZyxsp2uEPs
SuYtZktSDEBLzUPdVm/xqnnqSZzkfP45OWoBKhM5jmcP60esQL0xdZl2Gj5H8SI2
HIkJz/+waAV5hdh3sP372fD729efTzKZt72f2PdJQs270wTx9nHw34+EegIiD8vO
88CD23B5KTwdfejkpp6jwgH5M4nryPIMzW08SaMoXuOaSgDfrQi0HlQvyA2NkaHj
RTGqcKqjiTT8ELLvE6uzg0hACeanGwnIyKtnAuCry3btmHpF4H3xyjK/3SJ/sOWA
AzgdrYqpWn4PtWkOwgANKH+Mh1Shb0GLDQ2xbFn8CZqdHT/+0+kOXBOSE3EOIs8R
duopf0qifJmk4JRVm8of7KOYxF7cVvkH+SumO4lFfwhRk95Mu6CO1PCulCJnnrKa
g5kLsLhvrt4zrtrZMhrciWscRVyGB2f66P2IS20ISAL36K3EjXjbDIYUzt4+OxeN
d2/Eb5WU6ADL3ioTwdfD55kz1dJF/WVeUeFwhQIjNc3EgsTSQq5fqOMH+dhA6FP6
obbJiE6igITXZr2Z5z9YZy9JZ7994fvuBANpkAxGrvVW0BAc7/Hsoo9rSjZHIxqC
Wds8J3Bd7SG4ye/JOzv1LNlv6GTkQtiTICC12vZyx82kkBH/6VxQO13As2H5NvWO
qzvGldPiXu/dC9GroUrDOsuAHDlw6mFhsREqzQ17mv0NrRpGWfoQR3E5rZMRlG9b
Wevsq02QdbvDWjoOjsPghGnkHNjFsj+Y7b3RifRQYS/Disuhd0xhOH4sfOBZ26PR
bDcIU80hxVEvHDZ3TurACA/TIR6wSvK7hFi3+0ABNJS+UlZ7/WAJ+KtXhhg3bODu
THN1Mm8m+llHVkEfHm412Pyp0AECFA71osDWcVvabZo+/mwIASGwUWy7OdKBd4DP
s6Ni5iIbaE69l3+Fh4TcgWpW4YZ/XufzymLNRRpGVQdEK5xMS4lkPymQ74oV2I8U
JQWez2SiRls9PPI888bRDjFhucUB2/WscK5Ix73PjyP8Hq17FWJTDHNL5V0guIZy
gsaseO79Ewjzar3hMjVZKobUj7JZ67Ol3HTbgFFivrOT0whXmaKSYkCwBfvoSF+A
Wantj0z9ll+ilaQmK3CUI8yDrhYM5jyIDgOaUsia0RjuzteYXKwJOTUy73ar5FG/
srSiJSHozGgllsCfSqiFBKdLV+foX1gIO6RWo3VdCEUjrmVSvsh1AZ/zw6BaZe7z
kI+yTn64RkL+2OoW2limfmPEPSZCkK57fYmcVk57q4XjTICrVdpX2aSpL2hwtpWC
6fx1zm9OBlEyp5cMp+1e7R+CXextCXpVgsVtfpDVV778kaRRnBqXmsv3AtCSeDvG
EMQTaDJ38L3uypsEc1jvJA7ebk7lAx+V1yMKxd2eZKHtkCdigubsnM36znmwh7hT
TlSGLicpeiXDAgF8jJRO1Ydcn6jDK4vijQzdfcUrzGuK0AWzbXsEo2OHL4VoDq2o
pxW8zkJO9QDaW2VUZWwalijfI7X+vgrTW5xI82jwK9PfgGShKoJ1oZ8nAI2MIhLN
bc7wIgCmDWvbMaWfa1rlH/omHg8UMSwvvbW13LZfCBaHaceC2cRTvIWQmtzt7KdE
o9WfAcskv+i/cZEsX46OaFKsD5gR4f2038RLShzs6giMaaKntVB0RxymGQ1vAnWs
5GX6OTyUPAgpkIMIFjkelamXK+5v4Q/q7umRuth+SwPwLjMQ8BRjvXlTeazykb1i
50UN4JtHWAEJEfWcIT6YOgRtBKoqMVYUNjaRBcGbi3fYmgD6p7OkQdzygYGNmX0X
o4iaFvAjKKsNHYYbZxfoH3h54+JL8CKnDyoaNHJ+x1dpKLbb5GqioTJxUybiES5b
RwLISh2+UUmsWQzLkaB105acKNC8z3xKBTKkSny+GiYXmyPLcoKdOQJ9L6/msQG8
ZymXDDPzkUoQuPeJWbQA1//HaiKEGn3XEt1lMQ4ji50a/TJPXKw8ct8cj2z3j7T6
JuT7xYFnqhj7oQH8y3WKAtfinx2cvPHiTpb4y1aXaPjyD096e1QP4NwovkmLZQ/P
GiCyFebQBQP5VPrwjfmaqq6XqNaMyDJSuP3FTu470bzP92vSCGqEm9OYOEynhgMm
Vq8WkuOZUHFV3AfpxqI25T5VpPORcksiyHa5zVWyCfeAAGdFPi97fFrkAqb0e9FZ
TrBBVqKpfhSecT5z6/tecIsRteDhhsRdcTyz6b/7OAIPIQGFwC5h2b/bV8TKHn4f
OO6+QD4yh+EgMIVLNCN72wmV28Gbo3W4MSyh3fSSXcFv4MdCmJItGEqhfJudmahe
xPAOPBe+WASAPdPjwaey4sVbQTbokRzvI+RI4T/bzetwAviUXFpYEkYAvGBA5sSD
dssSZVQJ7EfE0sJjHG7GpY35eYtiRfK25Mn2uv6/Z/inb3XuNlzP4KnV0PEt9FAv
hyQuVfezipHHXFOdesnNh3J9hqqRO3+J43U7yyS0QNDc4QIgz0eG57sre+k1hDkL
kHCUSENTshx3/CaSrET1AGVXZGDmLGjNjk1Eh+m62F3Ub7a103GNe9bX2abHgOz6
vMaGZhx5skHR/e5+KgvuUlGxpaEaU/ikrgnU8RxMi1MlV5w91zaBuouUT2qspoBp
thI6VrYdNYNqP6wpKKvK2LZiOOWRlYZjXTdNo3qU/lWI/KcAoI5pUjdRtkmyxrIx
ZIJJ7eU5oSbv7LdgAuj2CEFSc1q3pRYMjtML9PoNYR0Cd6wE/skiMYqYxx4ZazyH
yc4gilBNlscnz0BbDbKfKuXIkIMap4j65rxWf9GV5RlUCVxQXEmWWfqA5k0rAy0/
I8rY5urftjTmffSMuVncN/k49yLj1x0UURVMGAGa5aEr7qUecvctVrejZ45j6cq6
YLecf9FnAYo/LNNHvqqEyI2vpypsfBcXdmWxXTSVBJnS9LwszXQSSFKTjRlSEe0l
7UCYhrLRB1dzST2A9bnCdX5szHqGLk35s7aIclWL/c6RdoFC2RiKZ73cNjTvNE8F
WHtTYRy0f3oGPo9iadaQuqxSRJTMQj7BcFVlziMgVsyDOL6PWTGo9FkIn/SCunmP
RlKLFMwCtfEBZdsXwa6YrhIrfy7r1/ozO6BNRz2q3iRxcqJwZIIOkNmGvTcTiy56
CT/XENOtI2kub6b6lchFrO1GPWWWnLBLhMVZpNea4kCwA0n+dtu5rmEc2WKQ++To
CNV6icvk90SLh5JWl3nX0okzafHQYNvck4s5FL7McrBWcI/wxkZnZNCqG6QcH4OI
gqJdEuJQWYrpeebIHNQ/0CkLbjbc8GCR07nDyfRh8X0+fVf8ke7QT/ZNbMyMtJ1R
ElZUNnsC2LTPkuSKz1FK1Tb2o4XeYP6CKsLTnnDoLF6SSn8lIxhqgIloUmO4yaYD
XvPzcEDbtO8ZgtCPYORFBrvYDJyNFCGb6hRZVe58zPkQHxwNvRt0KtC/x1UHiNSN
HF6BkosXLRLllfr1neGAYDo1X8QG+In41023X0pwPWNqvDOcXo6XnySwocYNMbT6
mXoHe60By0EIO41o7lddoYrouXDEhLqP3Sr9Rxxdrz3MfoeKsCPbVh2ganUHMyXV
6VYUAOugRiSwbXvnHdyh+XrbQEDDawjYYVWiiBWEWWEnXMEKJVfVrxL//QHDVC89
2iiftl6xfkdex+2vS4p06wDGuTAKDOENaGUAgn3yE/ITcn9lapeZ1oDDSoyZSlN1
mygvLy1hwg2JEn3KdtimuEkCUBt6SKx1tGDEuFsElovg09h6CDrqw5Nhc7o7A0Ew
Dr4+1nDld25wl2NQ0qtoX6UEy3WeXK0Z/EFBRh1StuNgYtB/1GIQUC43Xl95Kibu
+bGZ29C2L6XhgcDA5XLqlhOR+0p2MLEtBAlMwtrDqKsW1rcGH35qkLBToJQ2hyqY
wO7CgBe4rosdJsifZNmsTKa7dQtAVLd2551o6QFfdepkBCX0bX/+LiRuLYWpPit5
luh1lTgxSe7vPSgS8eB9zcaz4vUDb4Kk+sQDtna517uRje2jwcpU8C9V+8bLPqBO
2+PxwNtKjfKepQWzjbZcr4K9tqDP1X3LHtaAHhc2uDObnXHaA7DC2Brnz2CQPy9H
SlHk4QCif5kCgB9rk9xL4vg/q/t+81KNgv2ncnTNJcOZUqoWO4xkdu/VaV9o+Phg
Slxbl4HiaWgNQWUl/GsNxdJEsMcW+YON3X7v4WyNXW1egs3BrFX8m7z83g1uZ8Gn
LYQPsjyHeXQ62lh0baDbWDLqrIVpLDg2JIvFeuq0SXgDci6s0IINZub+iN03Rwy7
4i5ugA7hfJVtvdZvmHAD8iFggBhq4IjgnsYQktXiOp6BGGCFZdVfEaMbLbhCxS+F
1XO74EtNl5+cOWpucpm21BV3u96U/md0RyWfzUYTNdjkpVPKwUXRXXD7Xb4PbbI3
B/bN+F0k8BC7jLFPEoMG5ZJLrHACO2O63al6Gik/gg0F8Ku4rHTu0ZHXVN7hA1fE
wJVTUDalq7Uj7W6C1kdMVqWl8hfCs4XGBGl2k2IpsJj+VtEbMXyIaGzbN2EEBqbP
90L0JAVycgx5tPFFEpsXTXegCv2ZC/fYDnADNBcd30B2a9wExmIsnWX0jPg0oT0A
3denLBrm+phXOwzFV5pRwGWXoEr3D0D0RB3N7Ny7Zgy7CrWRrJ/eUFsk1YaVXBuw
uGDXuwJnA3M48DKH+dTgBNpXeDy9fCcv6ih9b3hgvKlavSOjeJF5I/gyhGXokK9C
X3UmaYgQWg2D+jryFKwVU3uZmQyCFUQn5MDdM1u5xZ5Co4eFq6LWb7tJqtkAJt0o
iukwwYV4Jd3SfQ55RGLylz27li4TryVQfkfOP1ER0FCFRu9cOoIGLr2R0tof1Dt3
bVCXAOClSqygRzEOnfu+KYAQ6wqtwfE1R9+WQS2VX/3EO2gag9AX+v3KfG/aDEGG
wQCfPjW443Q+lKvPsDJr/zSB9VRpRkzNLF8kDVjd9dAMbWi684VxVDWWqqkhqPA5
rvYsnH3R6/ZtHN8AfY5g2cQuI1FGlOVZZ7VjsDlqkfjvM5LZ6Jn8iEP0GWkA2GhF
7vAWZzDrImvAnMzm64Qu82bYHFI/v6se0q4IlpjZid9v+D+/wjwcqppayVKsOHdK
t/1SxhUTYn2ZPhGP6INZ743XAWkHdsqlYFCHILh8LnuY14j6TIKOPuMirmKdFmej
GKbRW26bPgVVqjeU1VmmAhoSP88N38DmFPvlcC5vZXlx3FPfzXx2LI8ys75PlDBI
N/AOhipkRVD9gCRtVL+6kKHvzL/WzRMYH+LPxomyI3szB328iIreRd2jS7KZpTsz
CC/tI5gtuHnFxuTr6wE9tuQbOaIODgPoQ7cP+15Z3tbJG82gACbXQyYSR7NJC7N1
RFDesoizxOS9bDJ7FLg4jYRz+77152XmeCo0Iu7PIi4929R68jbPd5XpPjtzYTR9
9LfQSjNrDrqbKraelf67jx1+ji6Wr1xr9YbXK2BqbTaTvcPfDqMGB0YdNKGbSKlQ
UNAS93sGKOf0JpTGW220fxAIdr1VM+gWVplvdWz+jGKFm9pJgkqNfJ0PyPZzNmTp
ANEGQI5VRdKdatWULxSXwyzTdgO9iI+KyYFU4xZ0oVFV1zCe0xozYaJkH6zLDzpq
5QSOF3/BIidOX8Jawsj5EC2D0XBljwUXCZO3OxzR46N+Nbmd4kJJOgZLdFUYH2Fv
vQXNNM+U/+yYy/Q1r+c/6D6COLA0mC8I3BMqrrcScww2VEr8tkQy2hrMXQTtxUxt
wNDr/23g8zHyRc7m9Xt+2+cj9615Wo0TFrWEngtn5qXSbfLRWUi8T02y+bJSohc9
Jky0q7LY7MtNYsALusa8imIi/ORc++DFoAsm04CRE/lWloYtuylgRs54SdOcrkkJ
dtSa1OCflRhKdFROo+cJV0pRJBut9nWRZXXE/BpHPd40befE+53jmrIrU2EqQAe+
wmO6GOgrXMBeRLsdvlNtzYshMmviOIahv6iv5NNUScSactmqJCvHjDlavQVfdoY7
2jZD1I0MTcpzSIzLdK7GU3Fs6SLTGkihRu5S2lfAZUudBcYzTGIWY8wX8a1bZ3lr
02DdNBSWBJiKPo7UW8Gf8ZRdQ8oC9fc9lqZcjfb0jAjbUDN/0La+wP8swnkGGHCR
IkqsoPu1nLY1y7B9+HX0kZtMwE/ZFAy5eBybGYXn3seS3+pUNPpuSvKNvgXKpIZy
klIcE+0yqqkMNbwcFefceGkJKyKDIvD4l8L/O0bedBxA0+ZIfW1qAIBzQ0Z1A7RG
4m85QY5/JIFmIBaSwtJOVQkJ6m/SnWGYHJuD9xaPHakOozzcVQ/SoNOeu7FDSHuA
kgTneF/9cmEGRrBbRuCAK/9dudVjB6GB5FWpoeSyukuVw0BeUFF7wx6BKJlEi7qq
Dt0YaRjZcuw1dFjCISBe4vjJMY3muoRzXvMujEM+bUgzRG7bEE0ovpIi/WRYpo+j
Acj4FXJbZB5yhYdKDjTqrEvN+TGta9RD70Q17hIEy8eOZXiQaUgB3ueIcQeaCdzs
ILjLwbqdBN8ptmsYRzOwAZuQgiXbntU8mQyFx0U3SwPKGZUNB35x7B4HVxdLJ3aX
aKc0b91Dn8Ghc0mVY6TNEVjjj5IbubeGjmYbnP2gbQUkVYyq0avd2zgW1B6ELzMM
ui4buaAeM4YkF0Ljorvk06w3chE92FpgfK7bCr2C03Ezu/y00V4KThq3wK7GuxF4
+pjOh7P0OgPv8Arx7Fn5CY2ZRRJC/odzhyRNzRCtOcRdolAuJNQkZfP58ePDZEVz
TKjQspbUgeEHZYYBvx8yDh3ErjK8JaEXy+utuBzHa2cCAN2EQRJDRNs14MWG5j9/
LyoBnwbyQb2M4g85cGBr1CDWiwcQD+iWtiKkh9UO//FsMFHwjZ2ghF/KQOmSpMmx
+45b0HFTgG4eSNGklkgujHguFRWLr8LHPXD3hfK1W/KKicIZ6iBAGFoeLZCsfijW
XbY0Xkdil/Cc8GfWYOW+IK9ykdNrA/Ur6dGwCUpJqXvwmBJv/tBw1QuB8TT9w2NG
tF07/6KJXa9TzgMAyLh17ltdHsQhKKq/vvSmHzhWW/fSYpQ4Fis1iL9Ictz9T6A5
N6vJFLJOO1xRNgz/uFOBpeQJ02CL5ipRgBYEr4vdqFQtKzFg5Iabje8LcXjjLJk2
T3rgcZGOYX5z2v12ieo9csIOSijexIhkz5parTx6o0JU7OQSsCBS/9w0Yzh0Undi
dyY9/PSYhnrU2De2xOqkDb1RSg8iZt6w7KWIa266KOnh8M6NvPEGmIckt6UNQai8
E27yiELV0dw0V/NrtE9H495lf3xOLIbgqZkEzI1Ciqwrankh0+VWI4fMTVD82W4M
UkGw9MBRv46BTgyRZU2buj64mOmSAhHmFrSjRdnryfQqlDF0t1yO+OxPAHaiy145
Jop8JGD3BEc1nBn21uAZ8Xm+VbK22pEkaVbmVbLITSUAl1HdmbeP50IoPxUslVTf
slObpkSeunL2VCvKb/GKnb3M66uPVukClzMY7P4ahhN9A7TOxKPMYDBunHNRYolG
nEn+4781kqATY57k/8BEXBfhBJqeEGutM4zLcM1xZ2GJ84neanOP/zYHnuR38Yjh
IJ9yfJKonA72sNREFhwvTBVZCWlxKaWy6d9mCCUY0AopylpQYtnfZ5+3ZiyI3HJd
3qm4D9p+up48LUVeV0sV+I8v2Dx4lOcKR/JLwdp0zqk+SF2D2XMrSb6FYqL//ntW
t5I93IC77JxYmMOR7aZ6JvlJRQOOF6P9Xn2rLmoKxB/luHRHEKG05W2r/Q6ghuhW
nxvSQyMBfeYc3/yDnFXUYperxnasmkcCiqR9EKg7tGf5u07IFWsFmbmxxrbpTv37
/aS9wKvo0fxmxlz+FzAqNSONE+ctjSH8ECnARx3glxCzFwCbjIm3CxNzYkFhwtjK
NNRu/dvXYtIn13uNocxnDV271SP6C3UvCKu8gXwhqIRJsH8oPObY2n0JU8qjoFJ5
E1RfwHV88yJwiATzIqUoD2qmhgHn+rNoM1ed9fBXZtWBTAr/0lE3/qxEdAv0YApD
TSZcSaYwMzCWq5sXkrvqsVTr0iiir58Tld2+UuKTabXtKaxceW+pajcNqGIl/33q
NbZQa+oZfYTUVaBmFjbBDNv8kDLK94S5U6fp8EG2Di2rM6KIgZOXnUa3iSSgy7v7
IXGQHcase7NZSPAWw++BfU7oWNzV20HKxFYeIBKUU639eI6dntaCruoWFEe1470s
3lAqHMr1azVv8mgdoscEZOZfNDDvY/wpz0n8JUst4ixCbogLvnOtQLev67oUi60b
8OjbMNs0Tb1OQRMaDf/6rH1L0UmYvKqTF45dbr3ujmD6MPa/kIsTLvdOGp2tfrgD
X22V2p27Td74HSP5FROwd3hYACzraDd/+iRc+65CvV8TtayvbXtXNM440aButtwg
tCB7VnibGx/3WgsutvfhtlVGjAdmsmXN0M2eBjp1InGci3EbQhaay7j1WFFYkv7d
e9O4NfhG1U4PJynkDJ35nmxb28LeZykKJ2jm766MXp+u7BJ98oUAewuJKEzsHTHe
gdz2iB7s+9dTJrwrUbN0AxoZEkzc4y9umrZory9CXAVnM1eer3pk0Q09mgQdBntH
uNDpeyAKgXgXTKBLwpbPOPXrmmBYoKwuuZS9Vil3IKblduMB+cFiMPJw6L8fCr9t
qzBbnXuxFDpN6WHJwamvvCh4rPwoWwHYkq8HHMUOPiFbWGP6gTEmzfn65FchM+Z+
6MUlLym9Qm7F9c98S38k59x8QtGeNUnrzUYR4eqlGbJetO/AWIw4AcBSMR2ewKMr
GXqHJpg0U8uwHe/pmpQDlC7rgr4LDRPjUEqwlK/5hsoD7ro5tPARJqrShC3TN974
fjmfp5JRciHm6lWweNjNdxQkmSMATxcZd2V0b6JdCs2B2Wgvt1UzBIUpLIpbzMO5
i1dDGxVh7vKRo0ZC08pO4Pol0IEb+UOaez21ju3GUHjJ+zEhovliK75SVA/P/cg5
FEJYKtJWFHHB2hC7Eypj9pnDBCfB67yNHw2nZ56loYKKksuZGnoOu+1rPYtOWKKY
aFRWB0YJSf1osiXdKcISubU1MTs31/acRZbJRI6nkA7uisVSDKDSNZgGQnDAuBX3
bAmdgixq+jVkCM3Sgtk8iryjf95rjMxO5/rtCftr7PHqcy3PSfqMODKIZunxkvip
t/QGc2bxw0DwzeVWtzwA5jsnr+vp0Y5710AcPjyGZGi1Iezo0S4/8r7oqNY0jhbX
UyM1Uv9ztHm2CvSHsrdeqKnGMDyTaBZsI4Uf4E0AQtxawG69iGe3I42a03vZ4xBV
eTe7CJYlvvJ+nH1biquyd/mXyowQ2dBXzgv6lQWQEttb1nTfTnNc0DeWgZ95iBWz
T5V6OnvFiLd4byQ5WPRwinprBlu07+98QsW7dP0pDPSoozFI+9LOJBvEWp/nZIqA
hy6E2Kz1GvYj2aGOhMoxJU9hwRgIQqT8Xs6LQ58M4OVfexW5WUTPDInqArl3qpGz
5FyyOPuMilSAursg5ULYdrUC9IGgi3473zh+jw/kr2PVF1OU9pIKTzVva16lgAqp
Ua0CtKYzQiiesAkf4ovGQhidq6OeZ3QoMo3EU0Rul0u4KLY3P18767BdSrx78jL2
3NTAlAccUBNq36+LLkMHeMQroScKLXjB9RzXFUMIPlPApk/j5xGs9X/h3EcxcXis
O9cAn8aEKbi1uXCG/5UfkFDM9rpVnKk0wwlliW+5QxG3P2+vsr3qkngIzd5bm6Rx
ur4t77+xfQyPAj8LHU/L2fhHG8Dy0c6DaPpoYSCaYPgu/G46j9UNU4b3dHkCYr2D
hQ7rFZ87bvGnLbMHie79T9/sOD72HfiWmxqWIZ+JSJzS7e0JaC0+DDhn+BDLuFrB
5tFhlRFaWudB98Dz9lbeP7afGueCY1ihH3QDjl1Jyl2zlO/84JXUXK1yQwJ1rElB
95l66vQK1N8ZO1VAXNC2ngUHfBiawfPm9C56d7Rn7pxJxxNmpgW/cw2o71y4LY7e
+FVmE3HNErS5qut/DxP//31zwCpVx8ujiGQhyRhsExawKYiNpyRlZzULt1w0bhQs
zLA3OfFi4Q6wIyVwxN8Pt0q9xyAcyrN1c/GrzEuwXgpntF0/w/wo3Pb4H1TyIHyd
r7PXRJVkOLi0eW1wwKNlN0lkvCVyvW2NJe1fedXPwfocWQgIvJD7tZwYLrrNArAR
rp/ip+3roDCGGAusBqml1DjWY+o3luqB0IVoT5AficaxQsLyJIriOt+Xx5yGNoA9
soh8p+IbKpUhHYxitYGKHEfKw6WVfq6rSmoD+z/3zxo5xd7BhmNYogcF+SP5XmOu
+ADWL20q7CzWbQ7Jtk3PJJWHq7Kpk7Fv5ob8mr2Z5E+I52shAq39174rrUFziI7A
rtNh+38xtsy9s9f5q0GyNyxBSR8IC4pGzqWxLZB5xRWmY8qyt/sUFz3QUgW8fmRJ
+v/UhDk7wTO1/Uf1h3vGPxLhMr4GXnIr8QG8iW9/xEPlTRgGnaDi6cdi5vap1qL4
b3W8P3agxAFIJ7onCFCdMSwazB3jpcfRnsrbh2PuPUU8krsPxd5VM2fLIzoP7EFo
yLlcGp2kCllT86UBVoEPx9VdYSAEnf1J4cmCp4670WjoJmlgb078mXhCI6UyQcP2
x6mD6LFk5paRCo6Nl9F2i5ZLBzSTP11oq1Fzhn8FKst1upehmljD4XqqCj75x8dU
X6b09p7A19e1upAcPj7VmbbiZXXj2FD0ssfysNT53hIrJG/u08omdgbH5fo7RSOZ
nkqOPUMEhpzqzjqysDSUPdomBSBgoS+bNUdfyBsRJVnDDwdNn7pBGt6HH/SBNi+4
8QGZMI6acrbsSNcXMaeH2RKAUo8MzCMeFdWa/3B10zVZyrBIaNlUnT9QVLG0rCb6
t7IR6aqUPRd/AsUBe908Rye3skDh+mDWd5m0pGLkTtVq7YA+2nszNAhlwxTUEKv9
dOVPg+d5QIhOu3JEXoYBC0yk5P9epK05Uk2zAq8n+USOcDdO3d6KpmUbbVgIRGWg
m2hHNJpRydhrVs5Az4g5Nzuqnc2BVdVqknqbrrVeAUwrXCxLoGPLVsGvtQGUoBu9
dY90mVYsoSHSbajxa9wVd56VH99Dw+0ikQCGCOGVgtCg4I6DRXlZeqhluN3MNeju
+FE/roFjaMLij1aXGe2RLmUzNcuRgu1/FtmcEuph2nJwBgoC/KEqDwZmSGfo/Qf1
52R+DVU8PsLIna3CE3KnKL7jbzIJQAYN5CtnSURMuI6/vD2emqGFO8cULndtOuF7
GK0P+7wF9/L58SUfRUSddvlvT9YhSqS91b01ridSeszErI3b6AFhIX/eLkCIC0ih
p9a/NJRO3J8F1LVj81UyzJN09fy42aVKNFduUX6MYgQwrLHPe+GPhY+7FPxDB/MT
aFogwB+2sNwKBR8AF+sTvCkQ19Tm4lSgyht9pC9PUUlovaOmGvPbHhU4y9dzro0v
vS9PtDM6zTAbXWHpsFk7RC29EVrLlQ1Mc7vPVnzOAqGZW9okyiX9e1kZaLCXcbFA
pWds9sdTEIrMmlqGRH1Hvn1djoDRoW2/Bl+8h4sgAMPYfMyz0m/3IvAn5iMCb0P3
aJDs0FWRHPfe2+UHUfDg8yBcQs6SmrF8aTrIkL4AicCcnXGxcbiz5oxB1l1+zNiB
PLn8kVuBZ6oJ3DVESK03M3lQiEUpaGBBW97o0jtN7NsSpNwbKYhhtdn2sVylycTq
fjSqzbbeb5gKVF84rSRYpRRh8q5ZRNsZR8wcnhCryNvlNnN12P0NLOnAaCByIO8m
krdB+QYgDZ3JyM9N7ELIj1et5aDFLyKpHDMfHZbQh3K7sW9V8ivdR33Yb+sdTGPa
FOQZk9HXXLGIMXeMpKcHztUBswLUwHUtZam0cuxvr2stGUMs3V1TIhqhdNvb2+qz
DdaKpuQsa4GuQlprEAWdvrj+9LLRtCbb4Ffjw9+Pr8kx1Jx9VIB3Z9ywbiFfB9Nf
ECjF+CNZTDtUXw15+BMXF4GFEsoAvx5SJ1kkTyNNI0PFqAKdfwkKUg4TGZN7Di/W
pS2sw5iyNmsbpo7zYEGUjYpxVgBxC8sNSSyZ8YJ5Oh2w3mnQ3etFjYE8FGjzUNA4
hnuSIDlABTku3topFiyadGdmVuMrVc9r7tDMD+yVza8FQsai2l2d75gf4C0QtazD
TmS+PY1tv2TZPZgSdDbH3dLsZivCAfIk2VFHyaQcYdCgLQX9WqeyKcJGVYf52bas
GSv4Qz32mu/Hqf73cOvGY/5HUIvh6Ea280JXZ28KumYj7lmLp/tw8VnFkbemY2kD
m7YK2gH0GeM3U6MhzHiqJv/eetzTSr3Y4dlVgT05Usjeo5nFsPt+Ba23IOnh0ghq
shfL12dTp4dacpdgXWS1vwmy/mTcoqNyyg8AT0H9W5dVSTXNTtrNa7brdQW77ltr
oN4u0vlyMiEBr3eNq5yX6OHhtLEDEaJhTBooebyVvTumbLXncR+vrjKA6Pgbk/sT
xnOLyF528lEFYrlZIdVIaIuoQyyt0SAQjV9GGxY0JHWH+gUrvkhWB5tQuvxSbyCq
a9X+Sg2f1fWVF+fQH6IMXsnIcugnaILhY4Zdy/AH/s4W/cHki/KayUTaUD+Sec8q
hRCHyp461+EvjtZyGyM8NeB58//dAPPTEl07P0cfWaHcTjQA+SUBxMdZ9sXjdTpB
s8FOXh1IDRq8TIhr9obT4cUmnbNMHxhzeRiDtSWtKX2b47ODWAMChlfk4W262PJJ
zRmtodHRXC/k8G+lts76R/IQk2s+ooFoBl+UFzjLx02/2r/g8NnY1sX1gprg5Zsh
frHCTIXFw7RRMyhVMc07YgnHyekSuAxybv/DOkbmrRjILqZwX5db1fRDb5wbLh/z
kaYlhikSo6njxlVaR7ehSmqoREKjiJNWiyzy89TaJDpo+hSqrtSnAvdldvuIq8B8
jAps9UIgL0G+MHeaHneRKjui8w8Mt6E4j+nkNmpielcooyx2IHG4S+9duCnt3aHL
xQCaZdTcoLjeztDsQetjati0G+6+Fd9czgHRkp88iz4sUZZOSDin3B++AEq6eN+I
2Q8HudqgVVhZw4bdcEr3ljd5LwZxV5ptHMN+ZVoERDWNkRcahCevlWD8Nbn37+w0
cpwqm8rRtrCeINAWtA+a4/E6V3iHf4DRud9zLKazFZeuAjflQ8KwuvoE9uSUdWz+
flkLVN+JqaJuErfxw6UhYrV8Kianh7wvLWY43808eqgdZv+XDTzM5q3NSwjQ60ju
1EfJ1FFKzU+tZKkyLHSYvkfMNNkRf2Zjqyp/+4NHhVO7MJICtqNOCkx0wv9Zs8y5
5/zMcNDsY+ThwPxNvT0TEbZnPkbSlszsYkCA6Z2j4i9eQZticR7zGo7278yivNZN
hlqJ5YZ8AC+wUH3leo7TWmR68K6KmdqnnFhVXKiR/X1IScdwOJYgSEvpCpsXEtz4
0ui6mN3v/imJHN8PK9b9qxWjztcchWWJFQWHwF+g7mFsm0E3OjBRIliSVX3mwNzA
nJG5DoO2K6vmNG7yd4WnWp44KADE/vY3grhfnDwH0bTnz+0P4xhp2FlpWrznQAzP
M6wpUYi/tDnjJeO0kK1Reavk4yRw551gx+jYQ06exzKj6tXgkaJplAEEKmtcQ/or
TbHLiTVJY1WSRz6hNykpMeZr6m1S5EqPPYZe1gr3TAzUaaKt4tEtApDjG9+wy9BN
KoAoukA7T9AUiZLZFPs64xqO0vVDM97SLSM+eM/vQGdUWJyHzJX2Q1BsLqISwcsP
0/lRL/yj0PrVXFkHNCUFs1gwsIg7pjcbBd0YE1s9k0NPIfS8/vDSur50N0GFtxNZ
DCSn8T8AieWVYWwHbGfmfLVsLZyHD0Q96bTNvvyBF5DBy0Zo/V29FWsnt5RmImA0
XlzCmdrhtpieV5M3AB4ISUp4Ub36vyLWFs3MM4GyncC0KGx8qOOFJZQuF3pF1ZOb
hcbCHTquyUNUmq7pTL96iOxafShediFXtCZf1OHreL3Wp7DPrStOc7L/Bm4f0KZM
yO4u+VprHtUS5+0nINwaQ2cHyXmqzMB8bfuTxfTEE1BWfh97hWm5Xzoh78o5acy7
/TNT7ZzCvEKlaBNAK2ytCZh/mZn+Y6ncX6W33hg4VrrZNByGoC13jVX+kj7UXbGD
WxsdTxCuscKuxMG/LVmuKdNvF8FkiqUo1q4o1wsvErJGOJee/PxVsNUOPeA6CQv2
Ia9TsIml0YFSNZJmyCUrHRqlz4K2UIUSbGGpbikXiHpUSp4pXq28rEeoahM+2hfV
ph0eJNYv7nh1kqh6m8vQzS7nGXr9uCNXj+ZO4/LoA9HP2k1SOUEfjRpdb2k8m6YQ
HAXkK51ClEjn1CIMXcGWUkdU1Z7J8SVMf3l1+sIXHW3P/gQw1h2jrOK2P6iolCDV
q+Uhu3WuXWxJucW1ag5EeAiNo5ulBr5202Pi3vbY503shKCE2J+z9TWAj4bycjjo
4ZVC5jsNLuSzhqpSafWdAqQLrnHMBvbe68bILQUggJTD8jtBPXNMJhfLGxdwfxrC
9NWOfWjXR/kz9jBPqHiv3LUCJC6xLSj1e+6C6nOSYGqdnc7zaSQ8QcJPbKxv25fO
pwjG0Lxz9LtR0Ul1icqLBeEcIcgMvLGYNN6DPMdxahuy+2EugWo00yuZaN3n3eg8
mXGOgzHw0v/IGdRiXdIEtwyX1k0NxhodfR1gFSnURiBI40pBOiSP0k9lBYJxC51C
d1RkK4aX+eL/fcUlCWy1mrGsOugFrwJZa44xAZ5HgmaWdAzRM2JLrzQRFYqjroQu
AYuyrY21td6xznJMRuypHxKgVMf2XZw58TQwTsbPIy5nWh6SxxPDcjh0ryKsetLV
7Yr8kbZdrTqLOav2lKo88VHPTmzf/PRlKOyicGNA5Z9423mA/uVuEx19Da114A4O
P8a2x9CNS+n0O3oDruzAU2zkbvNGiQqR4UxZEqYxRsx11e0pxiBMafgjt03BMBPB
zmHmuRxsJkvuJqKyfnPRZMAiYD8Rat8DHqPRMAQpqjiuCBhyxvE1nn+L/hp27gBC
mswOXJdOIUN5yf3TpkeHWoyDf8PElUP4pTiCTZHNpcX3lwgRJcKEgWH7TjCOfiej
P6X14FkIQ2+T9yrmwFT6ch9MIUnBYz4jAwr34Xr7pxOrTYjjfpprjfrBOp2prA67
rvqJEyQUoHIBfTiyhmgVmygZnjfd8ohBxts1LvXRS7djBmwdvbZB/rPDpm9rKoIS
M3iBiRMSwTAMphNsDaPkofBuBxrQ3qkKwnmeh8Ob9Wct0itRVwU2owz8/aD96lMP
qkbB/VPYTrMQ3rCZ4NoDUIHZKBis4uhTrWfNW7al6TLNzwT4J66IyuE5EAbCs480
J+YvBzbEslrhElZV9ODsimlopwNEBo8CO7SKHO3NXACpj42woZcNZ0cNbfOIM91o
0RsI5XI9R8zNEtJ8Zh2PnrUUvSnXNFU9Q68h22Fy5W/3jrQRHZbbnnlZ9jETmehz
/K+CJLGCJQl636nIiu+rFgJJr3doSRoG/9sDjmFm2zsr8bse42RejRRfAYQ+e+tG
X0Z9CDrKrVUoPsUc8UZHZ/wcRHvnHDaF2UDaIZHpMX958m2VveUWZFhNS/YOLy/8
sciiRp65B3ymdWvIVQ8cAqm1l56DzaDpZei51f3N/SUXqaSATyvrSdp+iRa6Dw87
SEzjjdX+La7sDXIGxXj69mWC0+oQmJ2Ad5H97pdWtqq1Lvg/f25IQ1aNV3HofNVI
12yre54HbwZ+Ce4g5HjLSyXsB4L/VrPQfbxyqM6P+9OwOSvqeOquKHUzhfleycDm
ikLmB7XGpbqXmTtmDQm7xT5LuIdY28+OdeMhX2K5SxTFX3JlV0oDZfZXDdlrWx3b
WNt7vpVZdvd9akFUfCsRnpaBw4Wcr3o0cfWCGRjqTqWzRrWD3Ls4jLupdUeUC63H
WItmjAz8mh2R/G3QnWZScJvMR852M/mHQt0uteVfqoXNazm5MR9l5XPOSRzTrbSt
iUNRlvW0F97enRB20NHUOw4TQi20FBKNFkLg83VjSWvRDUBAa4ihU/EqO6ftHEFD
xCnINqB+jwQmEuCIyzaUQCn8jkp4K04oA3YpZeh205eLkW7H+xJJBAbkN6TyWTtf
wBrpzk+ZZYnw610IVpmxpxWlFbvFQ1HSYKV/NDsbzYWd/O9qYGz7TlT03Gc6mSPT
gc1v4vHGWxhX/1WpjyTpDFpxJsnBgBSBpxUPfdyKLWmAD03YPZ3/uBNwakYJnob3
JyXByThu6fyN/1W0S43n6aGuxC4Br67QNBZwkZeWCcBnwm+cGu7dfgjQHTcYY442
xn28+WZ7Yxkkx+xakHqh0qFE0ueSZO504QyN91P24ay7ozmE4+YdY5UedIQK2xJb
e6BGIE6WP732K9G04lXZyuGYz3MXtVZnRoGJtdg2zeV9ipUV7ihTvT9RFp95chaM
bKcN1QIIr12RznXsKMJXB4AG/Kx8kDdvE5tSVw0gWFqmvdiulMsYpiV3N0YR/bAb
nSx2HkD/FfdvmSuHZceOKK/dDeiuJy7bqpgrWKNDonYsdM6M6tH3dlJd6V+/BYgE
UlhnCSYVJQBrRvHhcLiiakcBGOBJvQ1eOsJoSCBPvYRwmW75oweQeIuf1Wux+dgB
3+5N+EHMsNcNFYes8Kgh8ddZjUOPpEAMdPMWEW8AxFqa29UFZD3ZXAvKUq7BKID7
maHNC+3rjjcNG8wbHHqNxBpaKZXoSK+UPwdiSEmRHO1Y4Otnvt8zXmvo4vjzRwQp
r/w4JbsFzRZXmfsU1Z3/mRGxzDyp8qRE5ZTt2+3GW7pM9riajTUuII8qbidIqjxv
8mPdpSONICkamFO/Md7VaJbi/ZZD1ZxXlzGa6r75rHEGvHAHgdSsM8pAb51IoM1X
tdaqSJBOx5UyRWWM3rNxSRcb0gJ/G4HdbBFGudOLsUGEo55AiNOpcxzHJNxh1pxY
wykiyohMDDsiick6YW+hrzhp9JKJmk8AaiTEEcSS58QoWozvsgOOASJJaK+cV72p
735buSOzhC+3Oy4We7nUtOBqHejCEYtcP+nrWdFfs20NrAwM+YF8UxEVSPriryjt
MwWqFrnxUBWQm5FK0h/pw+4t1bbV5XPHEmGMlIv1e65raL9McsOZqtPOJKLGH5N3
jfaPnlpSaXaoJN1GsakVs4ivqI7GMR+BmC3ZIgs9mTWMnd493nNOj3hCAfVOK5EW
0uKx4ANsTXJu4g2WNe3kBt+pozpke0oZ9AbIjW0XMt7aUeZ8o2ixngIVAkDsP24X
yooIe0wSmoWc8yJjmrxzcY+O6oZtqAHW9BWZLO7Zyh6hzJJlubnoT6ZAVwqmNAGW
W4rJkoPyZs4AezySuvcWUEgFZh5gyA2GW0NfC+ZEIQ1vEzkCMPtB90T64x4UFSN9
yuphLShiv5dk06c1gZ4Uq8o8RXiqCPIaMMVr8Or8iXPBwU5IGKnl6ifbNjAvp+Ad
DTKAlDi0+cPyu4qGcmrYIJzNGuDFaKOeVoycmbllt9FNwJ53aik8PSdaSr4WewSV
84koZlLOfCnbWbs4FX+BFk/B++fP661UMYA34j+w3RwVSnpl6P8K0qDB0a5HtsUL
E0bAs4SfNpJVpI/fMr1t63bMIs4jvoHD15dyQ16GGdo+HhYRZlcqjL0hK7xpE95j
MGN8xJN8lFiO+IHKi3XZ0/l6Ps5goXK7Kf/wnI68xKWzLcacQqbnkOUfOREwH/uM
38YeBcl9DCKDv+yfKOzSB956tYohbYZ/Cy2VkEa1435gelr8Ot9B6BE/geXT0xH0
51cP1gn13Nb3gmECDw5dC9O/ITdTzbNI+EBuvwio7phCkOK/yqY1Q5kQnUC+59TU
oRTaN7OSO8IupuGT1M0SFInO9u8PA6B+PlDPf6Sd/NXWfv/3PXwq875tgZf1zEUO
8Bw+sjqcud6Lyh5pWWU6Mt6kptp25q67H9zdciG59KxsZEGV5lA+lefT8WfnX3Jy
Tl85PojEUrRtVgfokmfPPeYG3FT+G2uIDp4BpOg9u1ZfF0ZlJdXk9If0ZxRv0cwn
QGpvqq5/kyeweH4c+RT8nG2W70pmx7nStMItPhBdXnVO+J2Avr/sDN0b7u7AVAQw
iezvIv8qKnfamFURDFVTWBHHEm3hCUGZ+dep60I2xtAEOlJfaPTBTkXF5IX5LO06
q4RtwZU8jLHUpOYs4f6HZFHAFbOvTCwYTQSdPD1YFYQ6H+2vdgHSOL5b+b/Cgu7E
qdSAmqvaKff6cDFs7hlp/k+Q0fs5VYNV+Oy2aiFR+qZzQpGirJeaCPfD8fQgfxfc
HagdXvvUDwUHSZSwSTt2jRoICJeOcpdW+EAWtIv7RO/srvgOC7bqbFRi4XeyQFtU
jIUHyi+BP/AYJ2wQYk1RUWB/z20ysyxYuemUM++H5mswa6gHB/6XBcC4LOy4Dvrq
rmEKXStYoZP8/drP56tIZF93OfntOl47EaQlYdVKRbYhDOaVOQrEzGB861QspWN7
zJ5WRb+otlkw6HuUGtc4Pc92kmdXA7P0woEVUXETZ1V/TZ0xBbVortjrYqYfCUw3
PMnzAxjDrj1YbhIpnIr7C8UJygW7yWSBeacQhn54aGIonSoizw2YrOnoimbC+s9i
SDii7Z7vKqawEFd/WEgEqowvTRHByq9YUwAms4anZXgkLt27usE8hK3sEdbfoeVN
Of+AN081+I/fPqVkn2EdZEotD8PFuVOt5pl/psT0Wbs0lc95PoXUNyNxxCQhutn8
iFzgGY9UosTqswOkHTrgLkZTJFE865n/Juy6Iivrq0iOIGil9vAaW7Q/MWYyEbuN
ZfhjVsw99G+/3W8/203aBaRYwER8AeKrD3be+Fkt+yKfpcUbimvxwRAlpuxfi2o5
cBieZyG7wWsGiMqtvu5w1zA/XRanqFPDkFO03PPag0KM7uoQwlk861c0BoQ0BSqM
5tKI5hHx7fr9BsH40rSJKTa4S+H64oyevwGStMGiYLMs+75WxzjEL6mdHQat2+BM
wXKY7Tbsq0W/Jb8JpsVoVgfGeQMyJNjh2v8rpCm6bDLigZI+UNo+7Fl1p9trmOzR
2QyP6Z2kl3mkt4EH8NcDpKiQCxysAHVyFMbpX8ZGgG6pRSZgj37YFLmaMXwxcpIp
vvVwB43nHGXIBpXQgAHLiALgqKHXu3jY1hTLj7qlJT9jeNUAA78+G80P0yhVyaML
tkl1mCD90HtNBnuiEFz8alJTcXYQElG5v3wKrOlmk9BNMbavLbF0wMi592az5l8p
5HJ6v2KueCOhCljygOJcgz1HIQi/90LEbOlzqPMwvvBjvv/8SCls/3cG2H9iagEl
RWGeDSayYcTFl/l5WNu5Mk+SpqdNZnPkNclYu2xGNbasWmg+ayF6Xj79i/NBq/93
bC7SaB1oElcN3xGy9ytEbYheg6aebbCNXWwpIQJiEmIWGNliJsEs3l1K53U3vl5w
PKMjL1XI3ju45P0++D95mpf5Vgym/c2e3Ksx4Tupu8G8lqh4OKsDrPedw5Do9itv
dKEH+GUuVH7/5O64jsuxbwtDotMMQMWWhsuFAkWhsr0sLbgZvO/3ThXIoC1Q1pTF
c/zHBk9TuC0CVMzW/MOmG/fqa0Fexn4hCTjE7oPVBkiRiXJ7zn16exn3mmDGy+af
M8BMpYS2jW2xCsRLGmDYzWoOLmXp6mSjfb9FLMRCAAQOSFyyDe3jF5heeelNs9EE
rJ+BHjrEKqkFWJrzTm12DRUIVCoLABELgn8Nm8aexdi3FTIxBbA8y3zkai4DUybG
/yluwi9Y7wEHK/jYWpgjDP5SSrMY2wH+sajkN1Yd/x/pBqF10fopWCv8MJwnb0gb
bbYeFpT6+j+p2DmTsg8Amz1DypZcOYM+UNPTkZ9FOgxOHSkQ/IxnX5tgqn9GcSPa
8Z3/PMMPnnh22NDO2ZI1w5k6oauoLqQawrvE0EUEEq8y6C2LVCadhkqJuiFBkocN
u2iqKkomCi8C4Ks6G+lVQWCwvN6qfxoeTiWN2p6S/PpnZmyyjZu8PHhg0V6y0yyj
vMP9Q8sylx0tAHuN9T0gNzpsPmKqbBRyu7gBHgA4QDmBBplGAJtiz0KcfMfkqCSy
/C/QG170N49tIIG0vRpdBPXJH1fGw3ABKydWx/dJ3lFMusBKjs+dzOFzVSz7wIbH
9xdqQ2zE/G0ulGrPe6a13RQLb9aeNfVsXxDH/EA5ne9SN0NW36P25JkdUVDzKQ66
2CtaRvIGSjoI4PMyJpitSqNdumX4J1jE75VTlBMJ7FFiqXG/RdL1Gr9yGfomqJJC
XQYGJIcPHeuxFYoR2CZ+Lkq4uxm54K+/veRPA2P6BfGMOHgxcJcHFijLUN79IrlV
lsYPRA8iyrTSFqmMxQ7x12iz5S5ntrd4pq2GxzS27Sl8O5IHESVKsQ9w6jrWqLk+
a4Kb9DKzqNaxgSZ7gK/BZoEZp/Ad28aJaER7RAanpHBjeWaHb4JWkH/VMK8kT0IJ
eBvigZkYApeU58c0Kzfiyit9qn+N3Z69OljsnkvZFDeg7FHFjESwOnqFqu3vLIoY
qa+ZBZ7uFzjCJAgdXSaKsEgr3St2yi+oQqN/CYyRpWq2VcUUNkqwRyVke5DQMTTK
IA2GQNkINCCPT6yVHmZYgNdgVrF0FPLy06+39E3okxYKcILfPeTvCnenWz0x13nL
kyl5DIfG81NsbhNcs0Cga4RF4XOV83cgMfi7Zv3eWgzvZ04z4yQC1C2XWQOQcvn3
ITPWN24C9Mg2gV6Zssfn5rFO1Gr9eT5lECftEQf0/+mAlhfFNdAwinGu/HDMKI65
jH8W1I5KcuYWjzN25FNME/Cg8UWsXYPX6RZZJIF7b3ygrW4xlaKSezD9XxQv8/Eb
bKzSrbh4tnwVGboVoef3G+Ns3GGtx3vWovcdjBND82PwwmHx4+GaLHZ/5b74NYzR
u7rmdzvhsvK2L6UJs77n4K59idHxCwtFb0Po0WB5inqAzldGzKW3vbOfvthQdKNx
3LXna3Aw+pqqgdl3Dv2y+G0Re3xPKHzKj5tvPt2wmcfM8dLiiWLuGDde3yiQnCQP
QQwfC1w2/Im+O7vPK4/8RxDlvuSAteYUuJDOaGyXiuMVmVyeYSr2yLn0Cc6ZwuOv
pfRENLZDDMOLtZlhFPKkIz5dCQqtR90mYJeHfDlSmGo4x7h6vRcP7lJKY5Ls8ADv
M2ju2hhkPqfgpr9K3sMDsVFETUwga/L2uwPogxpKPfzveUDZlEBM4ggUmkEwlFq9
Z/i/ZYHZcTUSrE6PLuAqvMN1SqCu5cs65GNVb9kMA0+XTOqgfqcVx4dm0QHnp54w
85nYMaT3dSkkKnbdQNuF78DtFKuNIwzmXnGM/eXoQb//PItDCjZvncLnAm/sKORe
pOzV19aQSEazcVAGNb9E52id2fwrbkTxH4733ZfkIFT7bV3qL5Biq8ohn04wJ/fW
2Xq0PjshT+ztrFq3/ErwsRKStz+493DcO1hx5zh9DwaTyGBqhuyCy7MZvjRA5RGo
tjTJUQFrxdxH1npWKYzTYSiltGJXfglKKWkZfoeBzY8YW8U9ZmDktZNa7z6DLpz4
ClaToemCFwY3JMUchGNWLLMKC8M8g2RXxU3qmKUmHM2WxYXY0PRF5bCnRgDqtt8n
g1j8H/M/NloPAPHT7xTgSQgANHsv3/Z8CkBYY76Q/yTaDy6vBVQtNlJ45yKwhtbg
WGwzT+Fgzod8Vah13m6LbkzhmVVDQ5prBFdKDWToEZGNCpNUcL3LyladOMnrLjY4
aUVxgswqPRQH4yeqZGxVjbDUxMNjw50XRRdsMW6EYaRpx31pPwC4kovGa6+2Xjd3
6NBU6MDg75+gfgSm6EnQbGoF0V6MwNlls1L+HvvH2f+TA5hnV2Iz7bG4JazKOGl0
zV4KodcqoZYbt/btERDcAKa97vR09xIw1B29el0rC6r4Sx3rhsJ464viB5Q0Xijn
2LKAqsL2ba/d5G+Z1mHvPI8wvt6bcff8GA31UUiQpJduqynEO8aFF89ksEzhlS1L
z/Ace+R58n+hyP0zNeSZz3PpkTgr/y0T6s5qTb+kfOPgkL5fo1rEF8a9XJDOHjr7
WBc1T5RqG2v2KClEtWCW+Lihnd17yAM31UbrkqH9g8I0/MgvxI68VRl4rHiQpimq
Ag/Gf28OJxSSF8XdD4yaynCTY2hR6vR/jsowXe2AwwXHKUq5PsnM9tnv8Sv2tVEW
GWe5qkHA0GwJtM92L1Km6Q8Ud5LXmk9TUXMT3sryO2jurS0KF/d8+v7FrLkvx6Qx
01O5M7rQ0KcihbO5ZzQuoDaz5Hp6EdFCaB8lUQNaHoWDCgh7VnzGqmkImLPM+y/U
fJQY9hAmpNOBnL+9ZHk5ei4ngv5QZ36tR6VWFV0qE2LlE14o6N2wHv3P3CJ1nG18
FnocT+BMevNLEK/TlggXU7j8+qYW5eV6aK+ErUdi7RX+T9uhTpcOGGd7TgVOnLyH
m0nZoHQ6Pu5wuS+JueffOwokuW7PK3LXaM3SEMZVwoSYIMAxHl3RZFGkoY/P9Iwf
MXlrBfZgN12EYB+C/gsJ9X7iNjt9dh0SQPYZ+00CARuekuwdR/l6YVy44Nq09kfh
cKE3bhsD5YwaE82S8gVWPgnL6+VWdLwbBLFzjDimYbWa9qdMsm1aROdKEdeB2bS7
SclEON/mDF4LLRiFBfL5rBnQ/0wiCtWLirUcm+CeF4C1z4ugHXGVdTEj5FafX7YD
l/tpRSmcSthXsNrqIRa7BjZj8A33TiUl/lSWAxb7zCyEbULzxarB3yF8eT8feELz
uiVf5wl7+tKIH0lBHQrMsWThcPxu0yFUigkK76Hb+pAZFcylkG72WiALN3nGvNnh
G1jEX81NXOKzeg4X4ltCzfZigMo4srWNDtiwDa/xAMgqNRmdWkRgQpRFmECO7zSV
DI1WxEZfTuJTJOBhxrVi9P51uZamw56IpqURCFxCyBlDFHbvOyR6LYgfrmBVoZ67
dMV7wQ0gUmJU24Hjz1RWlzEJX5byXWs7D9n0V2NgpbaesGIypcMGmWIeWizdgc1i
F4QOtWat1kaVLT5YtdEeGvpgPdJ7x9ePo6FqGtunl69HkoI6vHrJ7vbh7KkUS45g
xDqUZiiwTp52GAqCBonCBMeCA9Q96dDZI2MO+43x232EcvZHezq7OC/9i9Zumbew
Nn3DeukyaHioPATfCWmUwhsD1X0TIG7CcqZgzS7ObfAIFBPMYNmq9t0azFQx4X4S
6YitJ9aIjtOazQ01wpuhOdF6XC02F/qfu2yaOQDhLJ4JVSJTuzbcuUeeL2d5XY1e
NldgLUruPlyE1KFwAImTx/ThY3/QcFyph7eBKc6iQy125A1uVt+HX8LXo67w7flC
qJBqR4U1XdK7/bBziaEJYKJ7LYVu7r4UxWE9qUwWNAYhxzgjNGG647kreV7z8MUe
7YewMpPTLbZqMzO67tx0h0QOCIJxPk2xgqqSBj1InwJLLU2cfOokyT4t0+WfHLni
PvYp0033Xi6AFaZR4MOzmbtYAnya2w0hIG2wMNNIyYwuL74c+p/dHh0Lzrwcx4yE
55nhYSHz5CSougUO88jiWIxh8oeDduJ1aTBPzQP+Qi0gBTv6ub09tpr3H+Ay4VSI
9lJQKbq6CHYAeqi0rVZvY6Mlfe7FUAAD+mYUgBHvpoB+i7zFAGOCPoO+rphr8AA9
p+EounjCP8rvDOXMtVg3SucFv4xjcbisOORDTQFzF3yRyh0hZM2ebu3wALCyJ72u
Crq18Lsn2LNdjrHM7Zg5w9CiPGRu4xlRW17p2AvrBSwjCjn0/XGhfiFK1dEjG1WP
Kq+b+Fpb5+OGkuuVZs+4RFS5lWe1HEwPFHedLqcsMExn6TeMg5Ypc7kT0CA4P7LE
2PlzuQizMjlo5/llaxIeIPW298NWoyveWsHCknzFbzMwbAQCs6xsM/sRT+xQDM9j
flTZ4sdASGPzWEK/imKGddx4egvq6K7rni/rcb7f6nmSMJjW+WWtR1FzquBgMmSk
ZCz38yECHK0JVted6CiXajfKG5rOxc6ui7OeZ1z6rLcIF5QzV7UsYiA83oeOUt90
tzrI79pfvh0jgzo3Cbabs0OxQWpokFQchF642gZ65Td3wIc+Ujuk5YxnctlX7oTj
UGImWujAhqwUj/NP1X+8rZfufvwFzcPv2piVIUmejIKB176yoJ9rH9HG6rcn7LPy
eRW1fbuoXU/z4vAKfO146OLpf9YY+UYgxABsHM1G0p2fEkOC1EUyduHr31stBZny
UXHNHMJQeERHxAiwiN6Q98rI5++BnxF1cRoCY9D8oSjFAr/ZGs7yEpfxoYvLqexo
YPj2TleGrjIHpxrrWjFbyIvp4NJ7VS6C7J9S0PaxNAmUqW75vxMeY8ojOENQrawm
I41v5M24VUPR++1Qj9rl8uC2Xa2XsnCVm6686MzdA9FtrNo6xHGhOPVJUQhJKgOZ
SqRO+984vH8mSlzoa5YaZN4QuVymCPBIY1DhT7KqcIEGyKEmX7daCM57OJu8Wpra
ua5KbRFty1LcQQtaBTkOmxR+NugQQN9ZtWZnXKR2fr9b8nqjTyHXXReihhyAOaUn
URb8VIx/PAru+VxE+6zssPKIQ/xfOTc3uDioi8qeYcZ8O0P6h4fe7sjYPP2bDC9q
IzXMaLp92BlhQMqD1ZdbpP0tSTMcHDgPVW5GAOLxxNbfmXLDD3gDHGXSS4QerdKu
T+T8XQdYcIavRNRq/P9pjV0QnhLH+hC5OTDLahaE5g6CcLF7H744xGLs0vnHAFiY
YuekBJYFNkBsBdRfHwvaS5f9Ec+nh6Hx3Hg5v0R/oHZ3vOlCImX9sZ+bs30GKgxe
xocDBQf546TOLxOojDVLZfPCZqx2yjdOsdp9WRpbHX+NB2VH2Zzw0h1EY3Papdsg
CA+Qm7WwPpYAz8NK2uvQLhPY+Y8nji9v75CRLSMBeyOAyrwaO5lA2eYKA3NXrwIl
AL88Btxlw/go38nQMwrnHJ0x8GtPWuMxK971RyCiElD3QHHS0yjtO+RfXCuL2Pn4
HBQPxZvzFCVpbs2YxthWl2SzlP14sBH4T1Hy83jARKtEguNPavD12AXyfEKRVs7a
mJT4xfjUOheu/nFpKTZoNQ8p708C7tIyiXfr0j4yUBOejxwoAe2Iae3iRQwnL9GL
BXMSPNN5d31RsT8RDt0LlgXEXRs8ziz0Oit6uMlaHvn2NROnQuL6eu3uFqnHTwmN
3aPbnPY4Y/q0X0h95QoqtNOUcBouxpIR/g4ayo5//Apb5MOQ4BDEQ+Pcme6pMd96
FOGv77EeMoShhCD/YNXF5MdE4eTm7ZGN1UJg1kdj7hi5mkH4M9axFFQ/5LQZwZx8
wwmx00/BGYBL8OXrWf7fmzIrFYWtj2KX/bVcH3hvlbvcl2Du697p20OinRG9IreS
8mFFMMDnJN3idJhIyREJ//x6L6FllfiKIN1cxJqTwK+khomqJJn47Vb2Xv89kSYm
W7aOhxPPfRZgmoXVHlTqqC4oJ6fGJ+HQMCP02SdwWpaAZyqKZp8ScFJx86jiFQV9
AM/08JdzJI/2iP2oi8NFstDvG2vzg0yJXZRWGB9Kv1zmdvpr5RqNgUbA50EtOXcO
Fz8gnSD2D9dUrtlcVr06/tapm7SFzclZtJmSpZsXZkxZFUM2VGq/1kB85XnNspsS
7Dg6mgb95slBDI18EbNmRMVnVkI+PLk7Jpx/ufG+gvq/JNiwEG0lu3SVf+jvaUwP
qEz59u1zFaMVKapLIY6ladv/wG1Hcv34VC1M5/7/XiFcfrzUI8jDj4q0U627N8wb
lMVOvjiomaJhYwt4F7197hOnx9vXsJas9y8G1HykMPVsJFTbovEcPFQwUchMCBqz
Yl5C3OVXAvYPQ37CxDnMiAEkNEltjLiwN8okSNzpw0Eo0KYVMNfXiO7PNNJr+zaq
P0dSQaQogIn/UTmbOdEPHa3n+w8cr4UloQf1kzvVo8B5VueXwbKzFJk9H84lP9Ok
YFQSJkobjJ5CXyhWGQ9G7fCWLwW/z3Qg6rX9P54SjB8KQ2uk1y1yomYjH94YG0hc
RrkbJgCQ8Ll9fXrQk6lYUV/B3bfHuYafL3Z3D3oYAYlO5mBwn17W3oSoYKIo4h/K
XTSIFKSXnfPUroKSLVpfoQxh9ABbc0rV6Ki67dVXbj7Cm794f/LunoZGFea5hPb6
fyvLLn8JH2FUxvUoql0qGNBfn9X5wuk1+Owm/16TFvoJz1RPoLNl1cXtEZ8NtORp
g55nEjLu+9yDa5BHnLdU5Z1CLoCWcTSo9574XOuywSuzJ0WmlaUfsuhxV4Z6mkgW
FJVhIZuuiUqT9cDuqI9EiaBUwjUuS9nv7M2u7GGA7sLjR25HHvhhjpEcju6dvDP3
5PdMXZir3USG8XQiI09hMMrSPH8yY38NNYitwVVzurTJBrXw4ppmyYF1rAyWT+Ai
gvFLz99aCyg2NfFHQGN7KdbcXmFsg0+OOz+3Z7DnyQac0z4KXyBRKp7Ji/VJN+B4
et2fac+Hm7U/hKro1gRnZk5NDjIQaaO1SpKRBjJggRErLNhyMWgFnxR/W5rbANRA
JGWAYO+8G5viDa0JyUFXvUvnuL8G3A/YiFXLpxE0NPSkQDhap6ZenMtyXJdqRDTJ
OkxAsYGTKCTzcIcc/ury6h8nlOuAsPYDuY7kjlaBxo3+H9MTOotLrD+QAzGN1ht3
cJGYoidY1j5NZCN9GZGGpUFl/6RCWKzfPjp1ZYbBJM/PlnOTPVxfDT8ynxZPwMqb
wbZrASB9oQf33PM+cAEa/CpHNuHQfP4aoaW53c877Qw8dr87lnpz0/uBA0PJt3j1
CVSsuY15e/uN9W9sGUNrosv2jLoXrd8SE42O6MipxAfBfQXMjSYEJwEcc7ZCv82k
3Q3jjoiKL4c/RbXWpXKtHEl6Iw0AHLQmXiYQs/ZiqYF0lAeLdi6MHFwlEFG0vqW9
0i04IK9sz4VsX3YzqBSuNBLbqfZxzMqwLoXIQ6TfN+PHyOt7iYQvp5VWwywsFJqz
ysvgRp5oKC3VbFhjIsyLKpAvpuEmZG1S0NeIDgFtU/a7hr3Qmc2/HKC3CL9OkE6k
zMHtZLTf7TmTdcK4pXUHUzJBUSRGGVGmoT2nqysa0+mA8qL1OrVFri1YRwtKoVUX
6G7kPeZeg/ObLUvfV0DrcSRQn/pSArxM9s4blQWYNOxI5Iw7JiS+ZUYtkHgYUtdi
JLuZ7ujjKA9y9vpyENcdrLl8t7i8tti1+PC2jkRkWMBJxoSJ6pNoc4JPFiZS31i4
MW+k1O0e4rhJ8cvM7REIKQ52X8anLO8h1KcRNyuW8VFMHDG6YTvdSCqWzd2ivPlP
C54pbdmS872Yi0GPJE1ghRqQi8E5Drpb1+1v9HNmEWJF2ZPgfp15utvDUM0SMaAV
az1/3abdL2FZo55f5lOJ00dDhkWC1dB7thpeRJecSUp5IkTqvXhyasbuVWAmq3qv
OiENJKiDX4OXN2PITEpk3Rpo9VSR/kmGorAYcWLXn2p2cn+ck5JxRYo6v8yM9q7B
DZeoOjTRjxpbLx049LC4npcyLTp91dcO+6t2sGBa0yvLtaHhO/i/gfYjDQDaWGAt
wvfP336sBnY7KxY/QUUA16kuieu2t/DqH5GO3gmeH8DArK8i9K/Cq3hRHUdDGCZc
5pIh1LWiWQMCqHn6i5UQUwwr+GvWgadVuZwVIQQoJHKuWqgI4vj8Vbf8/SXrLodk
hfthe65A2sN//dIcYr5Spbj7+mGqVO+Ep9kaCVjeg5gh1yrQhMBSC9bWjBE3tVKb
/2+0ABx5Xrqe6zSSpcIeeGQ3uM5N2vhlBUz7+8hXHitQdNTyhUfILBW5DwQmKmTD
zTxcbigh5lRfOP6Lvcby2EeWw9rgi+l1e61gn7ATOBBK/mU1kTAPEh98n02TFiPC
/S7keby+KWAaBVBcai38cgw7D/mj64AmXdh8huK4y140YzazIqzHI2Z5k5EiGU0M
UrXj6nFqJHKWqWOnTA/ns35DrIwKf3WBgl7A3u9wYzp+unZ1IkM1J39C6YbM5LA4
nmdgYnnSJLuha/mqrzNprd6FQFFJSiIEDo20mfhr38ch/xcu8/ds/TalfZvO2l5Z
8+T0OMNtztfhICX0Dl69DyybAdr9N741mq8XwNdWp6ziVXTe4baxYudFJiVklr5l
9zPQ15Vj2/A5mkdbKywVp4rAid+i3MmVkr+K8kUOK9lHQf5Mfr8I69RDci3+OyhT
dWFvFNzJaU8TLUXPvxPc2/UbIPjdHp7HqKr5AhWOiY1q9nRC/KkTijERVh2R46Gz
DPgOIwqYjaREglWUaD84QdBoCZW8ekTMT1SVqkCelww3y5r07oqT6UwkihwbQ9rl
GLpIX0B1jlWJN+xaGP0kwkYj3+JtcvKPGv0O+5qFZzItdqJJ8JjeUmZCgIIEiA5L
jxDSncbXFaBk8sWkmJ5WPNh18HCoyeYRJzV62cIqR2zO7nODnn9g2h6CA6cCfXcj
7i1u6+2zB3ySLiLlM9hVFMm1dglwBRs5AmTJNVKKJMKoJb+FdNbsRAN7v8v4aZDr
xmrCWajGISMzKVa9Cm4a4jSS/ozRfhhGjEShzIHRv7iBa8JAAhr8b/2ZipTc2dcT
fxEvQKNBIybdnVMRDIv3GsZRPo8lGRGwekgE1eGJRLJBXfelY6H83c0hhYCltfms
WCyyYBCBM6bxA+w5qlAuVN4Jmw2jX/+Na6nWvQgamYbA2nTLJyDKw9eaRWP5OOa7
vK0+AVS3GaR6L176se+aps2/0XjtgOp980lLcR8n27Iu50/6hbnXOBaihSpfto16
Up92wcJAHCLGiJq0d4ZyRg1Gr0n6wexb5FvE9unwB6pFC1XqFxM14SVHmblz6tLH
dsMOBTb3JAKc80Mtfrn0PjWNUlve3F1lGJXBCWuoqx2GI52KPPx/mL/C6HtZiRE9
B5yCYtBXnb2yZZ15CLoJN5wXThpuxSg8uECtDZnekma4uShD7wHpfLX2eoHPuVJ1
TXVPoCoq5Xiig5D1TbpHfab7HAvw0eYhJM2sh5pck/SMMp0vPH9/8nnU/YY6oGzU
kDCGZBKBT+Ukjg+ubms53ysrxaowKpCIFMywXCSpenCw246GexHHvdJlGYBJ5jxG
hUyU3SxasZ9iLxEBLpgGYPzjrdRQjwquaHFJ3rQtlIkWu9mGiBlzm7kjQXJAbBkR
PBrhHv0drMrORO8eQIFEHIHISZQrutO0ImHGhfsO0fDjHfNgV2aAQ5Ikux8ulP6L
zvYo0LIHBYPCrhhzj4GNQbYYgApyZo8QDL9FdlGffnMNyZprZFeXgij6hCA0LGV9
D3k3bQCE6oy0aPiie4nCieDHhguNx06NW3fD95R1cRhfFSU72+9SwVZ+hxyR1F4r
QWKIIPIHwX2cndqSnxoClBdiPUVlIECTAL4PMnFvqmrJSdAScS/ysEEXDroCMLYf
d6OnuwCNS3C46fBzpeh4QpdxZD/HpR3GzqwWb0dmatAIAE0dA1o5307mcXHmXZeD
C2dHXYeWylrOb83N2rjkne6CXxx2SupvXwWRDgZBnlCDBioURW4PAMenMXK6kQVv
qq2YDlX4bju7J4PKFAuzikD7eB+IHkehsOGXFdKML4nKG4147K2BHrjfuU4rhS+G
c6ojjfmcBHSXZINP9rNftQQirJzIqjHSlmmt9OoWYKYnXt4eH916WUeNYWOQ9Xdm
04OklOuqe6IpdUXN9DF6P6LhvSLY8xdPaEt+1tvLe5MQO+FQHHXGLyflA56o+z3y
ox6ES8GPVMm+9ss6LYh6MDIpqUOnIXpPBb2fqvB82Hjbdq+n/u58wS3o9/wB3SJd
lMBVchgr290shaJ35ep4zGG92SYl3maufdM2u+H5P412C5Y9Eho5krL0AFE6vHua
t9RGwJELiKgoDVtkIg2dbk0t+5DBT5xlSalVhtzS9vyzVx6xiWmFXWLCNSkAk2ya
FLet29XdAOYkKzMARNaN8l/GgMduVd2wV1Hwm444C2YZu918LfHpkK3zY82hARBF
NXFbxRdPt1iPouvGFqimho1kCSVITm86/44Fice5apS3NdcPcN747P2MKJwe5u3w
wUwSXAq066alPcIDrZ4Z+9syGqoR3qIMEZQ7pVh1SZgWmO0HdEMigEqJz6dqUYV4
swMtbnri6yqk97bO8z9ZllPcYfK0scDKbSTHzqxoSvZa78+84AtIv//kQCnCwF8X
0OVFHqte77bXlVJOQwD533Zs/+BFEVwoElv/yR01Wla/e7+42aCs1x73S1EeTXqZ
EoGvR4nl0Odso8/23ehoGGZDopWBahE0uZKPrKsCDhaxIpyC7efsYdMWZwBl6WCc
PfwpvYr1/1e9Ua8qP4NqXFEWkoS9NQbA3tPbQ2548fnGx8k62Kai1ujanLltSMWJ
zk9Wsq23GIuq59AJxkx3w83SQvKqnIflBb55NE5dYczXWDKYb8tCTuRKeZcYZAHi
IMRICla7xJhgSol3aCxRFy8ApZemrYMk7dq3+xnSXoi1fUYy6oezptmoCzc9dnEQ
HaF7spvXmX9NQeX93TSPYNnBIyuPHzvxKfiEqOL8WpXEXI+74L3ZlFky5pKiIuCr
+58Pe0BORUsfX/vW2mzM0JZ8Gvqpd16uY/p75DUwbSJn5KtyLacBRKFcYz/fROBz
27olNe7KElp4g4htaZMAt4DuH85XzDRMqnBaGRsoXRaY5fmTSXc0gk6LVPtZ7MLF
SshS5Eq6zQa4YvgUbgQHYrtwkS6P0IZW4W54DHTsa902iOckDoPVzKt2VHqE0Lyh
kT3CqDMQt06iblYHRsjjcltit1Z8xD5aP4Qel4wTVZowYXtxnhHu4xsqxiYDzVYj
MUjLBy9VlGQojmCP3vwi2FPHOxp7ehlnuBLgwDsiuhID04sD/sk8XuvhBHBXgdi5
Rj+CXxIwo7+L2k155Y/EIcaW53E2OshHZOkX5wUgEnHsgl/ExaGz8l4vQEyIRBPB
yrfuJy04Xh4xXn/6TasnoDp3kAJOyLURl+Y2ZuVXobDJV7zbMZR2UdW4yRcP/MNz
IgV1AHXy8VBSJGeT/bOuGHS3A4m44mxvzePvo7G//Gr6lc7htQyyM6AQl8guOWiw
WL8yeiz0yV859tmI1oHnrrRrgzHzA9ZFQHQKGdFWF5saUAVQn7bPUSLXAflZ7Fhy
gvhUKws5RaXYAnHta4fU+BWcB/b+/Qb+jQ5evBUpVAnTk+pRahEzNmuCP2ylIIP1
3bo68g+7Ouj6qkr4eCX5XoVtXY8y7g924pQ1+qYlSNOVE/n6rOu1Dv4tQs1111sk
ywoC91s8ziy/S2/ORc3T5jWF2zJ+WAURPiGo+qR3yAmSpRNaE3ro2Wk1dQ2nCw2F
EqLxguAWKIXLan/osKITJOvcV/cLkBsDSH7iq44IQ5+pPvmoo1UW1LUNMib0pA4a
U4Hh61+ltZ/sp5ITtntXe//X0jfESYbgVTsZO4lcPmyTx16zvdVbsuK13W1UjCov
FxB1WwkszChjJr22eOANXhTDdxlRSDsL4+8tUBqceoRqj34CxZNjKn9EMlqowJBJ
/wutOPqBs4ncrB69sxN01h+buamMpvWaXxRMpJ2p8qZD8REVE+UnBXJRfsKzdXs3
UbRX2Qaczu1Jy8MVpYQgRMmIUKIJ7Aen5tnzwOxb78D4MkKqw0+WVy/b0PP/LseS
1ubmBWqsS4pCMVFutpffkver4z7ge78+8N6Qwb6gxp8ivIwOwZj/C0Pmt+8NC7Bm
UyO9M/Gttb7Xfu47ijs1EVMTORvIEPsohMmaeyTpBf5Yv0POnOd1EmnzZ6iet3ox
hdyABQE84Izj9iVn8hxR/2//hhgnTjd+EeYoMqTtFV31Ewr4lAkNilb46Jcte+Xd
AdPSEP7lPGKk8/wbflL21NO5upYfzASmozWHiiycX2pjaddHcXAhQWhk0yX8iPMR
JC+KCYtgT1mKchC+rsbCwdtNx+MVh5tL7qEIDtEJhywdEjjvh0IFqKX24ehMb7iK
VyFa6DfnMgwQdPhU8mj4oYg5q++vCYEMdV/l2lEhfyOk7fy2WP0ITBNKFp7Pnaox
hyVPkTjodZcDslLS4TwVuWj7i9KXBjqsUKUANHapsUe2OLccogS8BW6JGXrhQkGU
kLXWhtN3avIlqQaupuqEWrjhiLhGv4lPB1J4NppO6VCv9fYD7HC4W6M8S2iLkbPQ
9bsEGyvP0sAQJ9GoVjqiIUcMsYS6L5ntesNQUYVPhtKSTXvkW7iCpgunPqoV7tgO
g5IXEbih/poSj7RiYn24qLMBpooU2KkkApliseqnVS9YTQb/6UFkEEr6XJUQfb1X
Sg+8eiccTVzEMlTT4+XCrT7x7kDAGf+rbYKcKppH0D13qX30EGqkwKdQtVIpiiSf
iLXGLt/jgTWNs62hItRx9Rou27eWeGInuoEPm+lvfIXFHpQ8eGTEiu8z8zI/Uol0
bIIzD0zJsBePWJ3Ui+4J1NYFh/YCdZxOW1pO2kVZomCxIqYsmt4sadIBd0TdLwHy
d+RFUy8BeKLhH60/cIAS2zwGk5kzucnVmCoyLEs2Bdwk19Dp3jhRVqlfhZ2+QbvD
4hnV/FyARZtyz+3pVK68h2ASAjDG0eAXXhTpG/NJwqsA9i7Yj1HzkHl68/32eMl2
c2/yCbcjO5AGpy5EhwBg6FsUNuTWomh3pg/FxkJW7kNf0R5qmRf7YKfKxcVX7Asr
wmGOZF0tV6fvMsjBTbmuKn+AnIKK6MM7P/J6FZHoRmt0mYapIaCU1PKz5bPYtqpd
XSEYCG+LjgOtjFZ2yTTKE7+V9BDX80CwhgJgji3Zpp0uRQh4rSD95npIvy2JZHWR
Urn6gJF3E9m/niSJeR5QOw86bLB19w5Zqh19tzHQZb9o48S+ONjhxXb5wESNMihX
7yP8iHDztyx+yRW5c0p/8QoKUffvuXyhA7V8f1UZ1SdR+dqJjzvCFLv7L6wR1k3q
Js5yehEZps/0ltHShXi406rovJZ/L6XLoblj5HOctRolc9/D6y9r3xmYGg0/2IWP
gbfBeum6lDaWopO3nQT7qURLibGpfXVwA8ip/dFJVvWtPwvFRGPPcoEvtz9hfZXp
FqWu0JYO8IMZjsK/CqfhpNAfBIh8K1GE1t3mb45CoI+gYAvPoZnsKeon+E6QBh8Z
n1SdmPIrc9V5fJKSdLEWnPoLuR+oD8fgsx3STeUEFhEvMN4gxgyRnYkaBppLpoSS
5NW6PwxVhrcAI2nva0YfJzf3CXEorsnhDDBinNbFa4CribP9sBjO7z730dIcGX6O
soX1UJ0Fr0koCGhNLKL8BgfDwT4qE7v2Xt4MENqd/sQyOXSsgLuoxs/oWo3tW4i/
Usjuxc0/jolzCQF4OWJYkqfIB7xsbbaENZp41Ocd/cYATDC9BMCijdW2lTZLbeq0
5bLiowmi6Q9jrFbOCCO8x/83SyYlQIVDac/3JE2m9HP4Kq8xDIJv+hGaEtm9ashv
kIRxwO3GeUptAfXcfa++OOQsELng3QWlufqtLyu9fZLvV1m1N5mrJBt4iAzwytjU
lGdS1bUrPmvDYGUIdaPz6EmPMeQQxdo+W/Vzbm1os5ccaNRKDHdX3mlk3U9ExNCI
jp57hDCyqFaXNZvRo25m3byqRvrKNa/Dn87nx4WTFCeTs6QuHKhlEGsO5Vwqozwo
wH0pHCh4zRCLzQVk9Ct656pjr+K/eh3bJGa1IUCK+AVjIjIPd57rsFQBCDSIQNmT
sZtAfx/wCDBvAq1fIMdRFYcq0uelcwLI0+TJ2xgyEKRnzIxdFMw57pfXjY5gy7hh
OC9/sz9igivAPactNcn2V9CWBAz2Yt/+ryQJc/dUmLuDmrtW7gsVxId1ukvmEJOD
1yyg1G9j3d3MqCpF1F6fMeL0m6Rfxrv1N7IRzZQGNyH6cWFqs4w6ZEXY7+wiqtsu
5O1cV1CaibRZ+my+gr3OB7fjdaJb2sK42gizCM2sA1IqaoeWmR0fi4uw40Ib9pMI
VJmgKYtcQjaBh51oppNkq/5Hjqkx8Tj62hpzvibcIpeiogjqCdyOgE92MM7e7KXu
YOXm4yuikgJznGDwBydpAXfhWsp86I7503z8TOhShtapwIVBZwHF24apijQv2WVh
y8Z72HOwNeIeJ6qk24UrJWynHR0F6ISHFxLunK4XU8DbTn3syRYt61704Q5G0h7q
hhBZ+0Ex8KDqvfSFCKYWQb2DrCn5vpzwa6BW9EIje3pIPpbfganmio9RP3spyuUA
fS7YpjFMZWFcDiQJARuke86UlvoGiUXNw7Lft0K/iUwcFl6E5MVUqIh11rYEyPUZ
QJcuNSlfCeD68+ySDycxFJzfLdW80bShRskgSKp0JkYeuR1UIzn4TPx9KffoHWbA
tI8SaShj83CR8RVXVV/pD7faeYW4G10ZaY0UAm+hKB6TqFVCqUtUDk1MlPAzM4b/
QynJpGrMVcPWTO6iYdgt2udzqjtSuXmUBfId1IorrXdS+EHDmwddp1mKH1oZN00p
Ho1ViHZ5lrq2RA74ZMcZOisxYGPPzNahTaaEDcsp8P9r9j0NTzoeItR9SeL0R3DM
2mS2vXjbT6tlacCt79C52KjSsTpyY0dwszB+aQ6YNQPy8Kim7LBjPmYAWKbLdm0D
mHtjNZXiPnK7ywIKkZQr7L4khQQBpgVd4diAmLwMy2fU09Hx1zqt1BYxfZ0qsjFi
qNQrcpc4djk8LgrjQK618rGFlH4T4HbhWM4roBaS9pH/GDz8n1hH74YQbHI5sv++
whOLOO3THr/PE5xiy6FJtfpUzfX9phDpSZqm4Nke9inqEVOvD+OXjk4Q+iTFV/60
ofraR3J+KPKaKJJ3Er3mtjG7FwYaTd64NzR1OWLW6c5AklEfR1PGqW/GUkszFOYC
5/UYUwboL7dntggkFu/gFXs3dVf31dU3tvpI8cYkahRs3M3xPmsK2QKDDjhFmr13
gLtAVn1Mh8zTTHPsS602vVTjK5xZ83tR5vyQoWOqxrE5bRIKOm9SEJI4EUQA9Uy2
odICpaeclAt75pg7yhTZ6+V+FGnbDANe/x976y/RvT+6fhe0q6pfa/E0z4aQIxZh
MeaGEBnubc2xUAfkTkQ90MEZleITzkan0RXOaNZ21uUHzEcvd6L6aCoVKOpy1Q7v
0c0JNHoZ8n2upgs8fXXSH0kWsJSNn3AwUeyhrE7+lj/uqrYUeRINPxSt/h04uEsD
k+LEb1o2e0bfqLPo4YT6EaGRcW32IFrHO+LxwJ0XZKLmr3YTr8FNQ/Mhla41tuwd
+5ZuYCn/eaCjJ5Ls7C50RDT5FjaYW27D4bb6MLGIQmI/XAn0+hkpwT7SF0SdwnZ7
ZBsYjJezn6gQ/nTNhQu+pCuhzJMu4j0eoFb+LRqCZYAhoB19x4CTFgZDqUMov5Sr
OoZ1mNrBnq1xxDvGYNUb4xOEFQkImH6BglwdlCHOsHAlngNaxk2tOEje2M8UHYVG
3cvjBgBEbXoFz0y4P0lEgV205oRLaMx5hxaRI/72Or3poaEC510iJKgUsaDMV85d
WQpdPDEwutj9IeWZdOyfNk28tzXxr/ZT9xP0Yxci/TczK4CEV3UL4jQ0DtdADKRC
FFP9Ojy5Sk2AFV4Ut56GqpfJhvZ+jjF1CH21nd9gQWjxP946wtXWgS+fbe0AENN9
nxQnS6nsKcBA/ucbwumDNC+G7PfuuBAcsez+5wT82q9dVH7YPDt3Z+JG+Diy/1a6
Lel8KH+Z+W+BiGBI1I59LLcgvvTJOK4sOWVQVRgU02fjT/NRv/dGBOLTDl5voOCV
JZj18LZb5iMrpfSwUFPSgWCEHMUr40syL7Q1yGko+pUk9h019B3lmrYE/7iSNmZi
PQjjxUYCCxEyHJuyJ+oSj2wol/rbkvaKI7wJGCwjhB1MEzb+37dSFFthMMPocPqK
AH256ntig/t5OTY1OMVYy7B/jrIFlt1M8VgxQWq/9yTCu43Ydg72MqEC9tZTUsKG
ptDXjev5bNrjs4l5tcqj5iObKCOkERQ8DauhWyDzVqBVi3RIo7FbRhaPr1f3vSsX
soxlZnRW97iEB3C622vXZIEYbfXCCh9s9Q73O4xU6DL/3d1XyWSdfcbQdySwtFy9
SEA2YdcgPfmADgyUjLfsTAh4EaL/mvDeXaPOdmuNffdwxs9nMWW8vYeQCdL24l0R
jtj8ekuUOSDqzIH854PBPaXOjjan2mG5Ocz9HFPrTYVKqmu+LDHs9KdDF8mmPs03
kU2amXlt4sROqNnEvR9kit+VjhnBWxMmts8V551NvIfytNvfis9cuD+MwRC61Zg6
Fol1rGOp4Mybhfl5DfIPQKH4e9nURdFbfLrngmA++4dN+XAcEaJJRLDmnSvNV8F/
2VpQiD7ua0J1SKq4yhauw1MGYLctP3ut/xmOBUVZIncO4TAKMdZKZsHcRfk8NxQ0
9ya6s4wZzzI0HuhUJVmIETCfye0CKEtUEyAQiv89J+uvGYUsKSlCxps8/sfHq2or
2HgKxn33zK1hbCS33rARpV+jIsQI58r4l7ptL1PQFQWS5oY428LQRsY+ntdsV/mM
U7p6UpyznY1/RNwwkpJIP1z/c50zvzJgCaLI26swWNBjSXHN6IOn78KQIoBJW9+L
2mH+hV9tix+yQsGRlAKoJQy0O1usvcTUqAGpN8smQVESVh66GaGN+cSeGILWw0nI
SWF0/6RIjJ//sv1atplt3ixkk13hHXxNkcTevgnW3e3FmR0UDdGVZBY1fP8GEP8Y
ZgA5OnSmVv1EcrRTAItN3SHFg6cje+9Fa5I6PEc0ViSE5LnVA9tsX+uDJTIotc5B
keMOz1GYCen0PR/Z2zAjcmCxxKEZ+RkuvXTbi2fNw7pk1QLt4o0o5qdrTyrCwXFo
THuWfvar/UCQCruP9Qso4XUcWOzY9WKOsDAjHgdlnzb7Bf2O/cQRioG9AWMQCLFc
xnMw2edKWPbF7gwlenyGGH+p0z426QqrX5bpr8JznA9oxlBGFaziTXhcAnBaIE3S
O5ki9df1Ous4DpyT9dMltxcVZM+avzCs1ivsYHULrLSqxxQ3dgtoqFStSlQWZJLd
5S8uAei8DHaAtL/Mc/cJT7M6yyPcfDMrk2vDwHxKgSNqUpGfTAi88dpowsSZfO01
AqiJ04fYpGK0dr13VRrkVvdFL5ZPpyFrx84Q4Mvd7Y7jVYv+sgEQpd8Xiar1aKdE
sY1gtkopf7p7nf2Gs3fpumA6FOevAbJGrmsn2iGVaWaGNv1PDhjjEcNkkyx0u4xy
p/ecqQ4hqgPzp5LvMsQr4BopOolX1P6Yls0xffPsprhnrBT4oydHfiiWqMappa4q
mc6LpfYsH9wXfPvhXxM1khkG+U6lKRa76OHhSX3/9/FhTRQB5DNYhOZ19xu2ByKP
uegLFZhN8Tg0MM8Jtbzk+qJY8p/QBxf9kI57vN4yaqvAFje2yKbPBmL26t9FhC8Q
+3dQVifzCeV1dpmFXsm3LCbaSIKLihv80xB7cVq/MyDBSpQsa0xkxDi/EsbFbbLn
/G4iCCWQH8NcZLQCUC67rnzIOT9y5VxHUePA51PF4kGT9UWMcTiRyY6R4Wg2W16x
uMFuY8URixsgQnfqi5bBYIoutefXtq6/XzjWa0gZcyzThCsNHXSCb80K4bHBYVpL
ixNFdka5sTqerc/oxx72TsxRBkWhzhfL/8U9iYNcA4eohI9mImHlopiEOiszrXaw
KA6MpTZPNMxT8zfykqL1mGLiY+sGWqsjT6NWE4ZvelpfswZejL0cvFk++gezMIme
72Y0U278GhNXhjpHlrZvtD8FwuT3Cpp9MvbABdVqrdaGv2+3+RvXwy/anG7qg+NU
k4KwSAxQyODSVmRSOfBmxSJaHLo3nzWDCz9iMvw1jnJ1WP31cuTSpAhQg3cl2QqY
pMMZb/3DDBPX5enOpV7V9oM70VdKCo1AWDNaKaKQSqSih8/k10Frb9fGTnUAAQ2U
LL7C29r/6FhAfpRwaxGtHeDqW6k9TmO46F5XDzJWuo3KEHeqTPGDaDHWLFVxksDo
qoopHQzfl4gOPCoBA1solV3vp46jpDQD/ncx7DEsnrzPLOPg1c29D1Nah0fKxhJo
9S88S38vwAFBBNwfqC25TJ7QNpXk8ZAhSxjCHJjZ/E/RPuOKbWKEBSvHzNhULmuO
nej6/FMw8ogCVhu6cSzIE5MDvF1cty9CE0CSlW/2SIeWwgi+qNxFRyY/BYyHQQUF
fJMqMIssmIYejc1s6wLs9DBvM9MVccKlxp/15okhmESUfFg5H7Aa7p2CdwBiZdG3
jfhcw1Bm5FIU52EPILtg2qNx0b7tp7k6FX9J2QTXzLMoo/3pP43V8dmWiKdWRnWO
xO5lJvsYQpfyuzlMOomeWu5GlYGqD56Mx5o04Mb83/1VGmtODGW399CGiruLSVMA
Ullw/uKEyGAYnnWOC7rX4b2+IytVAQepXnoOWU7Z9jwbqMz6FRGxf60zX2z0+VX/
Ulc1jnzR+8VHOvA0l6C4hjboHDN2t8Dgn8Kv+V9sNIJ4dNPEW/hT3121Sfo3vc0x
jodRqopYnEMuihNTo2iYsNXC0tkA0jhnkZZ474keqtacCL1F6HJ9unrQWhaSXxo2
K8CB4AN0k0YPg7aRVP2ISufDcWImgqm+ihVxilCkykl6pfHeeX1XfKEvSpsLRviq
tBnPM2Ix7YPvn6vBz6AXJvdkozzqdEE+tLRMxnIiGQLGCf6zi74EO2DQDurCIlzk
DTvZeWYSR5kch8SfsBhV9wjOca4625m92IFbkDlr+Jnqo36ymhx4FtuSPxfsQAja
ssCdTk20Y1mDgy7DecVLWDEucekQaBPuhgpX6h1A+cJDHxTgBIk5142jJ6L08XZG
T+ECb8tMy8awiiwKZO95DwTpVpzdmfwaym+2G73gJyu2qvM2ekGaDcM3HcXC52SD
Dq7JTL6ND0/SiWD4npy38+PMH0vXcnghEzoJZaWSAT3P/ofvjMk61+H90ny9GISQ
62rs4jlIX1JXbZc2R+wY1XRNKsRdIrsu3oT2Va6qgC3yogW9k18rUdHiOQ9RDSnc
9T8Wnj/9+I7+Nct0HWXPQYxO7brXGWqy+f0dY3PtTk7YdvZz45GcJ4spmECjRtbs
IF8ewObmFenkGrVSP9s3jpycGGs+0nsM91bqyb2VQUgnGepwqnsC9MIFE25USDNZ
fxhysLBAaTxB2W2d1SBVlg0/if6ycowvtpr+p3V/p3cwHYI15JzK2/Wv2Bmy/pJ/
A6c2fIOVUhKPNzBvODyk8DfS0ieryYdGcaG8aqgENTPq34KLCNBRw90gcDuGVldz
O5iilFqgBcx9WVKpCdFimcj1Ikc9CsHqXKo2d2XB8dEmF8bkK1OQq/mj2lZpew1b
CkASjXDjL6pNbLv0A1t2Q5FEXmuuk79j+j+xPV2MZddDmPmPEKARm33T+2eo/LOY
n7Dz4JU5/xwhrh4dqJ26YnkmbMkBCUKOohuA+SI6Y1EHXWm98LnujKgIFvH5gqef
PHmk+ynkprDzjLdBJvAiqAO9OhVNA+9DlGTGpaofTLKsiXFpLkmUEM+VP+vonH2o
5v7i6h32a18Rst3FiJRuZkSiR/+61fdDGKkboFRres5Iug6dtKn49mh+QknOWdtC
avOgyuojujZBqS+sV+ye9hc1AoOHAZtJhKks5unV7APlQisssOLOYI57+IKgFH+6
lgt4P9ejCE930r6++8ZLjI7ItO3c6+5/98r4m8qbd908vS4E3eGfE5/ZoPxRTB7k
rz3411iYfRgP49jAOLmbdBp4z4Yu8jCF7/Msny6TghxwBFYkiFi4V1dsTkocGkav
BouFX6eOtgy6Yvpbb0C7XThdx/LX+GO/VRq/b76AxaDNiDE/+QMlFDEYMrLscLyA
OTCUY0JZgymo6W0fEthJa0tNq9hgvq+Skt3eNdF+Q8vQVCSHAAjbGRl/kuFx6UoM
7NywWeWx86SXGsNpe5lM2veGbc7fxE6i1a4aosHkitpU25QmgLHcfza68lLrztw/
maQyVU09pherkvLpx6xNUPGHW7IVErsVRiyeHG4vMprVrxSrxQnXyTwj2rc6UcSF
VqPXMnbLmsgBUYM15S3MdwSZzd02lQwTMgX/8pmCFFV7nVk0rktNxVKxgx9Q7e1B
6XRkyeV+EUUrBBAHMzjkFGK+QZLSmUFO1INQelWty5JFXsIMw9f6cCA+WmRscLdy
9bMDUkoocukBHaVn3Zv6qw1MY2XlGB2IXMRe5Z4jumeZyuajJZOo5eiUH/lj0Efu
sNtPwWLOx+qWh6doU5IUwuMe8uEOunkk+VTup6DUEJxVVu4SJr1+kzGHqmhvUJ9T
ay++PvEuikXnigY3hRiyYYJziQa+Il7/ZsZ5F6Rc5/xoZCKcIMYKGuURcex2dc9e
7WcQikq1lY++grVq0vg1GWGhcf+8kt62M7vP91kepqlqzrjEvnQiTjeGwyUjpCHU
QehRqhU3fpL4ZAfPMQsOMUrNRlZF8icWCIGpVYrCxL1mf115WRpzoogTYevoGtfU
H/rVDS+BpFhXfyooOfOMugukpLL+P5DXrQe26KE2Vru9ZiKonj6Ai1agpvM0cOBy
24i+iVgwChfMsgpxsjFJE3iHUK8dESG2y5YfuHZxbrTX2FOBP6eqUCxWyaUWH9qc
n2v2qxS1svjtclT/cij5LTJ+tfSwiIKLkY/Y4q703NbXkHoxaivd5jRRbTs2qZu8
J15nqkpnJk2HVnRDd4Ve46wKBYA6P2tip9hX39zqkbUH3WRsYTgZWCPOj94eZxfS
vGACyZ9GH2C8lwrJJaaf0c0IkR2dBYkwMEZLKooRpM8uVZC/sEhuIAl0/310Xkba
mZKqaa5Zq7uAbaGfV4c87pBq3NvQKTx4FadkvCHMTo4WaORl5wZklfzjVQNw+hip
VouglPitbjvoaRE0l9vyBHhORydmceeS4KmeVuuU0GTZwV5s0inVMrSw0djis2hg
QQQF+ijGclCnMENSW0DsDFfWVmOk6mLVIcNVg4OYim4ZoqGCgTnaTbpZRzPtzBiN
UlNLyOtNT05OuuuX1X8Up2KOECJJulid2k1ntSSpFeTHEHvo2L4e/RIN2BrCArYm
XjWqNTzCnukpdIxYCyksRh7+ANt0PnKB/NN3dTqDvPeccjR/ENYtmLyz+UguxCuj
d/aUTxNKH+XvZHY0wUsYvA+Iz6HJTwjbixsO3p3bMWLVhYiMbPaTOqCtqcGwnxpd
fCZxGKHXXRpkk5SGAAhVhCEgXRmAo7OvnL0nz++2RxepqJdzm73hjqEmRQ2D4vS7
lK7TcrL+l/YntB4Y7XkSZ6fpgelwbY5oIQeAcjHlwft0mTqHhXRIm4P2XSNNE8g1
GB2qwvtKQprkdC14xsUuaqyUAakd5ornn0Z3NyrFKK/SUkGMv65c0rK/MyLhtKub
54Ar3RDYjciqSKIbNDt4rLXBYJKA9skI8sFbSlENdkEIlk6nH5SAv7XDSkiwv4SF
LVlFnuqrivgrU3zqUbUgicErpZhb9mVL047rxbTjgdxQn5dF5D2dxM+zYlIDh6sC
FmVhTtsLWRRLhJ2k26HJkvQq30TMsEQiF5rxvr0vGzOpqiEXCICSXTIFuhrdpVQV
zfNs5qMLFc+p50Njl6enhg0wm5VGjW5k2UaVMZmtkBwNsj5JHT50zgkScw2qObrc
0J5fRgsnCmfNUwyK4hSmdKLKXORTNxVP5zmXNMpkiys9J7ihqx8Cv3+rHZAFPuUd
nIXTT5Yhg/fiYvp74zkdlWqolm5PMzwUsAtSlNjYQt7pRdBbInSVOpQCDo3qQzNQ
jhBQWxjT92/OTdaW6/xmqYOkAklxl/DVtJBrkLp6AZ370bKAmoVYNBU8IQkjwH9h
vK+4C3uRvgx6UNqglCJijmfVQ19jMjFXq820Zjd0Q3Fl/6szfAPnwMBXyPep6812
hmicZ9O0BvtFUYSe8mwZJmzkBgjRYlPPW9n65528RNBwiEySrzWzkCXrauqdVlHj
Quuasv/4gXllkXOj1pMGaHTIAzMt7MoQpEURa9GTQjMpCXJbKDd5LHtR3rUeX+eN
80VaU9lydcdVe1CaNdx4hKOLeXe0+9qZHdWQZKTwWhOyJVnLXwJPn7xASoHNpAA6
u2WA8abT00I7ivyGDB4LYT9/d/2SACGC27prhMcJNrDc97Dcfvb+Ju3+6gpB4vHL
dX5MqHPlRRHrF0EJLA1n2mm961+3YwfyzKKDM2pNHVqHQdtw7K6YnNXsjQABpzCn
xqG4P7CEf4OoMF/dNfnVDpCvO2eBySY4jPaQSNpEsBBFbFA3bhFMiD2JRa3r3Kno
wnGE7SRfA2Xj2ChV4h8AAspSrWaBOCpk3DJZBnI7fktzWt7VHKbJa2YAuJ1WzBYT
IHef5Z4bxFo5Dko9HxQfh4KpcyVWL1vyTkyOy6mmZw8YU5tjV6GS6xjuoyCp+YeU
Zbq2SfOX4iTsErNzbpLrgQGjQF8Rj4b2Er8mjZuoNjvN6C3q5llw89NgR95+4Pbr
DdK6mrFiPaczApKFwN3XNmlDvbnVBSwaBuFLX7kVeDgqZJbGs6n1VfBSzu2dUlWf
EVVF+I/zHNisluKxIlpy8UJcqddaXGVoe+fm/m+Kwzs9p8eKis0TPiPFS3LaR58c
oqUHfPSrx8siBg/FION7qyZGiGDnBY8s3mNqK3mrLCM8Gi3xFWc8hoUIcC4YbfRE
IFlz0owPopLAgM/VzTaFtwceHYHjRn/6L/nMQ1B2kVLQoQ81UEmRSHAoOt9kcpyM
GGjJ0fQhu2DP2y1YuDtx48LjGxMgUMir4M10S7VKdBz4IS/BlzRi6zxTmp3ZnyrA
tNxbnA5hq1/lWjdue02X1QlGKLousY/elKdjX/NNn785A+imEvpBNISmpbuqk6Mf
SizLetZB+Obxjxs3CppUfar0fc6LvHibTf19CtKMG7olwoIFP79TBiWff5YOQbf/
CARdL0wMW2+1lOA885Fl7Xk/Z8C1HaRawdrxjiHPRc0R5bJPwIVvy6wCkSTnx6L3
+0EJ1mllN7dCmMFnBdndt8kOtzl3VdyvXuPZNytN6rCLjM7pE5la2GsVH6biNZau
vtHVCcYxjpW0VI1i85Zm7jQbf7cdDwF/AxVhYIyE5YAXnKT6/l5L3JEs/2owWf53
iZ9fFoG8iF7tuGiJGU9fObggx93kKgzedQrBuOiqDvMjq7v6Mc7ReCb8DD60gidU
HQHDQs47jkooJ8iUmI9hV7iZGpTf3R//ryoXyc1siCMAvwG6aR+J5LmeEWO5xcxb
KA0c27dlje+DmocGn9KbKGzHcxBVvxHuNeN/Vk7CHv6zKTgLhVO37RSTJm5hCSV+
rrsjthpg5AwkQdNa+EDfU0K/en2lTgO1dRV+EXUN6M+y+YAxHsNxuezeNwubV86t
+/JzHCzwhPfooYpAa2KGcK+6hxMRZ64zUqoWjkAZivQPzXWpaSDrCfg3H2ptGuHq
Svj7HaOv+PFBC0b9/aa75GEiMjvtUTf/pu7D9W5S73sEJ6dCU5f1C74QkgWsqyWL
GnRH7pgka0QyLkr1YwekMhim1UFoLMT8aPDdzUhKm0o23nIPW/YZiArYPjpGRiIb
kda1DCbwZkcj84ISLQel6OBhSJdH1sbCZN7y2F3phep8RnAOau9kzCMicwRAafaz
QsiiU48x4Qp9FJ+WDUv+pJbGyeEMKUfKHJ6gpZssryEShQqsi1MVWCmnzS8N6eb6
oBclSHWMil4vuTulbCkhwEcjOqGHgjN3zyXeK7ycMs8pDoov87rMOgpCHHo3ztZ+
VxUPRfyhSGWsuvz0osHJdntjPo/A5rasqt/O5tqBInsMvfhqd9364Yd96ExgTsHg
kV6FFq2CREYWIrKp41+iS2GfIM43pDXXgQ4tUigxq50pp1r+bwCZESHO4uhAzvsh
YfDkFLkjg2dj2l6JYEhTI0hXKFxeU+BQpqfreaa9+sZHRupHvayoqYomTRqX5wAg
fBw3nu1heQJ353w79+8V5laW+ACHfS9zlvO9V73xJLKZCSauAQF+qox4X7p1PGbn
vZGeQjQztgRX3acd8LI5urXANmCB2KeZXO+CW6+xXb0/hQMKw+kGc49vSw7L+5ww
xN9BMNiENmhfsAZDWgBxQb/aObhR4d8pluCLCSOqMcP+KmCnBCjJ1PdIM5DKbMhN
+kU0BXDM60wpG1fTgTmXUuHj4BJj8oYEbA7HCni4zz/m2QVBE0wVq/kQbLOcuffm
+MV/jz2YsYQDNYsZ/Sv7cDdzvesy2PEODdAIEzsD5YiX1PpRcsXYXScJAoXjwm04
ko0soTzrPDQ2lb85j3Q/WfCwobFW9j7/8W9JUpCyIt1aQdrajeG4QGjsIaMhvlPw
vzyGYIstz+4HZMpS2tHSTejeC1ltj/ZuGc0Ry6SYuMlttVTPu8u+XbK6cpOYLkF+
nEUKHMOTMAqkVFSKdUrjRt90v4u34NlmV8Y4a++ITDCcME1fbt3fIys4AU7wyIQ6
3p0kcGxOloo1WDGIROJPVtoiGZGLubsV/LSfg7DbkajA7XxI9MlcCgU9nSF1SQPc
mDeTF9tkgUcXbfhFWcDwpvv1avrtPGars853y9X8bdxS+4emUGNmtumz0+UCnSqE
9H9Z3sdqchmqHtO1y1oQpwCo2vhJmCs0TruN1YZFhGmINB0zRCiPl2K7St2XqtQz
xaJKIybYM43IAgPYvlUkFOP4sbZljbuyg7T8CHCzUBB4fO3LSVxhrOcx2WgOp4R5
Vtvl+Xb9BswfeCs5bIMHgPQ13iXXY8MxxvXcYin+53yrt2sjXSyqAhf0dyoHxLZS
SzxFULtjo0I4Pew92KLcN/l0GfrqWKpyNnFIo9FqV1Oy9w0uVWxTgI8Sds2mSgGp
Ann/BK8yO9LAz+R52rfM5nLCLaQcmB3g0UcVMkVADVawPMzjWE4XCAXDi6fA2XjI
WDVwCNifdG0ef9oX/tkNielbFIiMckRj31N4+esoBf8jUT0EtJUGBsdmAt7gfdFB
QkLGCe5JAhzQbZMlCLkTnPPyMYaLD9xD/MQcmpU17Uxj4SQUbmPnff0qU5MnX5P+
1yiHKWZeM8jbxBah06kpoSSdq5lemjXs3VfT9dJEp8rYXlY5s4do7MMMfAgJbDQJ
04S6+3BTnZa/dK1b9R5gKizfqtgv1X9ZW0nep3E7naZDdyPm3einToasgGig0jHu
bw/q+SbhEOZblIb7A6okW3bO9HsTP0h3o1ZQ1x814c8ZTHq0WbvVRqY3TZFrpr8L
1vA3gRpwGehqEcVEVo0CQKHlHiZibWzyFStmauSlMZMkBnY5eAX9i54vBDXRq8kj
1JDcqSnh5OvP6IbbaG4e2cwq2F3toGf0rhRxI7B/dyho0WUEMcuvryQyllG6IcN/
0ioS7s/JSM1nRezOaRn3N1DONvhhxn0BkRged2PuDyt4G47sI9+set+DPGKap7XB
d1CV8XX/6H9WD0Pi5Ek73SAeemNu6UQfAgY66Qf29ROOfJTmotT04Qrt6nBcxalE
/VgQD47AFcyHI0UtzYykGHUifsEt4nS3lqwfx3d4ny0LxZbsPp6bDz8/ZnUzeOY2
We6P2Yhrh0xksKT6WrEm3AjG8Vx996fTPWbXo1hH+aBYD1V0/CmjCDhQUU+iyoaQ
OsTrBR3oVH8nsdjzYIrKAQi4wqirjPvXL5oTgiaqUbx+V+Dl4afV+nVWFjWcwUER
MdKraidNcRCYZk4UadkhE8b4RBm0vl2abU8o6mHtFaMj57Vv8VjFAtx9b7G0QpiG
c1A5xEshLk+8Bw3mkh6V/P4BQucQjaZR1xmqCUNHmczeNAiUToHp+bBLDgXybFEn
T7kQ4M+3REIPTeIvLFAr3zQixVoGIcSDpwDcJ26XaKAV+chphBYh+p8XtXmxtxjX
eROfrKCdNRMTnLtYrL2zgrCmEi1SuZlV/+VmvNuLHjO27lwtkBevGHqpQ3aPrfLu
tQ1WTv4Bl4Tl+nqpuSGHrVZhlbg3IB9ZB49YO8fYkGlqF/XoXYBf18Z0oHhmMtBg
3hB1cctmse1mNf0EaHzi0Uy+AYQuyqof4oggGGsuQMZ6Xxl1b6CwWMonavhzHlY4
mWXsh97soYWfN1Dkh2xOdN/rbSdEDEJLtRQzpoNOMhBIKOGwZ41mk+3auYROFAPe
wlamVjN7yUGnB0WEWDomB8rKEuwKkkSpLXBQTOT+D3HzSFufnugVZPKgrsBF0adX
yq7LPIAUTRVpk8YKoLdDvpgf9vAGA8YhpDhOByia/OXuqmQTO6k7F4PAV6jaItET
HU6w08j/WR8IqfOKC6hRzQNu1vtY5f/OhRcSzsKQuFZyIlvKHo91vr8wFoY4oIRg
CcL21y9CwkjWgbD/F4xlq457nYHN0NOSPto3SAcdf758X6Sh2AXfxRtnbE1biA2D
VdtIpCxkhRQD5G0VJ7dQXG87nGc9LWlqWN6T65oO7fXHNw2SqG6NCsuPJGXcrCaU
wbVI39A06LXnaSI3UXFP0Cd0f5/PHNtGxNU6NvvQkRfL0HXUH2b3F15bRRL9wcSR
FszUaP/+MO6JU2hZ/3K2snVhpuXqsWqnh+Z+gw3Ypk7uzqYKnluuRGte/7Z9E3X8
Xo7SD6WGXiFFkdWx5Dk/BBpFBI9N9dEjU6tmogPfoEIuKzUjDKs++vE82OIPEJKZ
OX7u4GdV3+EJ0S2jOx8EknQ5GJsLJnvTmPZzdxpOR135l8LWyf1UgMTlPIOyDy0t
vyIKNw2iFy8bY3GZb0qIbxoV1Ou8iQnca1llwYexFlnxWcVxiHLfdbsWXaRFJOVh
Pmk3gIvHGHbHDGntd5Vjvo8QprDA/HXO0g+R+w2RMtTNgVz63tke3iL8G2IkOWBH
BYmBsEm4niGIwWhCqawXZw5t6O6ETQQ6jUrsvUWDv8UTts0TNgAy847LWE2K76hi
emsvG0lLD/ai8+9bfa/4fLWg8OUOgwVkLLqjKtyx/VJgbrXzSd8whWwnuJug5/tu
uIl2/Ikz4yeUWJsjKcCLdawz5ix5cZt/uxd8w0VTMm7ww4FnNnsrT7mx8JAwKQD5
bh3Wqvx+VZVboYxmyYqVLjwTzkLiuh/V+ZzTjM9p5LKqqSLg6NMSmKfYWXbU9Lrh
6BvLMgFwUl0kzckYihSOyvucIzta0/YzX0XXpLvSj2zMCAjThL5v4YtOSn4aCknH
IMp7gMFZtD+6W1vuYHuAiW2K6oa8wnWw1ybNJeh1hxWCt7xMl8WSvlVGPtufRxvH
Ju7M6PKR5TfDdaCxRmFNfbpeYFhuph+DvVhog/yGfZ4yy3rYyvdgvEa+0BrBuAB+
uXuVVtrk2nRmEp16jJiXohylldW6ruiCo1wYs0KIcvCoKwXVC9gTAsxCeD5lFtII
uhXPLVyRms5BgDL02EPmEjAlszqMV/pahmI5vD7fKP1H+zGyb22cRyPCjUX6rY43
wbAS+ZL7vjMX7jSFCNaXS+XTT61Yys/kjNqZKNDVf8Q+ZFAXIUFiTDrb9nBNMimI
W2Y6Bt4IshQ0F2l4Q+I1MZXBn2HpDWHSV0f16ABiM5A5PqhMRHuf88zXGWYEOi8c
YrG8Nqk3pAdOb3FeHdjuihn8BsSuZIZCWj0fzSO9m7eiw5el5T/oZtkymd6ErFcm
+xTSkL6WscS5nKeJD1hoMsyCVpwebZ4RWribhop+Uqm+Nk7cqOk9TIX2w+N+9Gn8
YNbtHql28ATWXD9QiNGXslI5KIW+JXkCdhkcsdi1wqtshPUuJckcWtlHWwGl1Qxa
Xgs9v3iAhT7FnGDZrSW1zpwkvprgv6tl4xWa7MQtuDPXLdAoyfPtr5n8WCTc3amf
MQgyglptqQ8TYDyJLyvBfXxB1sRKLp35s0ziN2w7Gs/8AmMDR5/PiPq0oHWb45Uz
yNHIbyx8NhWscxjNajrL8ebPYxLv1HKtH6oG5m94V6QTRj+HUX/K43r9lKeSnlPH
rQa5BJQSUyNKSJrrPRmCgCQbXWudrH1bvb/rHecpsR0+gEOhfO1GeDP+cVrzkRIB
d+rDlS0yUPDUiH/ZhJ1s9StuuNmTiXUx26hr8yjsRzurbACvWFEWm0Z6qgs47iiW
B35G7ytxLty2YeRqslSqGNFQpRRRX5l1MXJ5IWzBk2sVHhUxARibVYvORv8PNp3n
k8w0gnM5IqEh6s6Espy4tldh+og9odYzYPsUXQmGiDtocKMZ0PzcC+SKTNjySz4R
DrSMPHTZpIADO0HgtBCzN/Yg6w2vLPo89opB14jWvx4oae08wJlQHUEAQVRbkPLe
YqbfiTnTOrvA8RKs1ba/4JcZoqFf5rTC5e8fCY0dEbLCvjP96HP/es6PICJSPjbF
8CdMuL466N6gzMtTeVF7O7qtTFCgb5oym+TjI3dKaHIdWAns6tWHqI3ihcRLBaG0
ElMzsG8SSP/21kNbPbyY0x16O4Z+vO/8jegyYFCvaRdy7jRWLPhlaideVjP7x8do
0C0oufkd3O1lDDNRdQ8TmVGr91zyz4Nj2jr/QEVJn+urcotCHZwDjxhwf6hIUfL5
HKp8uS4BSZrr/z6vlC8BJqjoWbAe3b3C9tH0lsfO10FByA4rGnVY8Ssajmh/ebSb
E+SqKgFePSq4OC0tpmn5pg4Ov0SWhGcIuA5wWhDA0oFk8od22lE35CYmpgrqZi4A
I+IafFJg44n7W+qFiHIs8n0iDWpnz/e9R2B2AIHlS/F7C+egUhi4+HAMj5GaNzFY
6utRB0YxYDL0/pkOZVesGyTYWFvBk/de0rubqkBGvwo8CKC0/fip6Ev3YxYhcDz+
W7ymE60uFJ+agC4xhFqSPfxv6wDoUJkKFUVHqXvLwGhIMRq7xCbgixAiI6z1Suh3
ioxaraxdBmZczJhYwZ19RclsE76iXiyh+jAWtGZ7uHw3XnzVIhjv/jnwHvmk2VrM
o5+c+oDDIitCtkENyLbfOlavaN8OL6r122JxJqENTtNwfg/2FqvlTIfdMUPHzshs
4coLQ/dt/Q/rCesZLrCF/uf47DeEDFqYijhbLgOtSz7n6+v4uwWaW/gJ1mae3BZU
95xUqv9iYZBggJVZKW4ubWQsY12Qsyv+DMzXTzr4EJsVjKuFPpf4VbaysSsZA2If
3ljqOTNh16AmjZyIjlwFK4LGsR5UlRGqJHGjzJ6geSFTM+eu4q9eoHxh74o7KeCs
cb6FC4EFnx8Dv0Nu0c4sE/H8Uiejul6GsVPi+KEnCqxuPjMv9Rxityaln8n4veRZ
lImI1YDnM5xVf1sjeyQ+mK6GXORJqRi2oLOTn7NI5OOiDaZcgmmWEHG1qEP5rm5u
3arkbUPE3AqpMn3v8KypEjTjzfCYWHV4+cFJ4MwuqnGqBU7n/tspQfeVz7ILfrvy
JzQh2ekHaBU/wBgUaMK10LUp16eDARDN5OGMkmyafYMvrd++N9tAm7NQ81Jffgf+
BrJkYe2WPeczDFs42H/wXZmnClrpG1y1DtBUtQ3lxHyl0FB1N8/khop7fEXO5PUY
h4ZYD5ZZzHDUUPz0Em0QZs2ULK1eObPnJHVut8DO1vCOJZKTgQqOTT0D+sSRZDqF
MG1uiFACIBVn5C0DvSM+eb5dQuo/cU7itSsC1fTYadg9IfQk0FpKhOsaGqnCYCvp
j6w+AWVN+X2sinNZiAYOzdazfsCKsu0qj3hom93qujKhSHCFWUEm0yC+Zqmt+x4P
k+/Qz7ZfjdrLTDIzzkIl7js06LARq7pM2zxEPDcG2BnFpJidLE9cKVPK5t0rMN9m
5H2dLzFooGsKoxT+GnPq/KJlF7zn7q1+Ze+0X5XDM8/JZC2zdEzPNpDZed1L4OVT
Vv5kTPuLpI2aY36hbLITD/18MJ7d0sWwHFAWE4zzn3m0UqLmO7Rm3TXPgS6L/n4F
/bmr0ZC+8F3StG6BiKG3DOMncQ29KibX5ym1yJwBIsi/ZbF+cIv2iV5J/hjZHtjM
1mL2RccI+Mk0ajJRkXMdfmMjudiNmHmERIo9GIMG7u6INvFPmI+K7D3Z2X+DsWDq
6N3fojxlowvoQe63i3Vg+V3dH24L46CTKruY2SDgRQB8QzUHbS2Xg7pCYRI9BHFn
w09sVeO2MbJrVWW+L42egK2+cIWaaXx7CVSXP2vEY9O1XCiznbSMgoq9bF96Irhk
2/MDlIpGlbRfsdxrLCEFPG39Z9gVeY77Vm1EylGlEFQbP7Jztm6UEYMyaCtfdgmL
3mOutjY52tSXCmcCcgwaKsgLyBCzz/U2QPTTQ14fB7UCJFrTaeHRA2e8CqLkfsvY
l4x9L7ikKKg4B+T9kJcRIuHWM3W7G4xdM7q9b4SSWX5YPKKhJXreNfv4K7Jnmob/
RSyGQxNFKcCx9L6Xh7Bc5pZEf3sDg6ISheJCotJ7jn100zJvEWIUuyzlbEp9/Bki
nXZqLR0oBrTdNL72cBTTKPrNTcK1YBsZHkdxAD5oO12wkbmZ59eoauLpVWu62Obx
Jsi5jshNxKbjXVrQp8+p/SD2HXUbCB24CWBH4xkYA+oR80WU2nqbEYamTasC3mWA
NfwdXZBrn83O7wSpY30sA2kXAyzbqLGNy+r3D91PrFK3RyU3rEAVXtlkdgKocQx2
eGlgh2/YorFmHxD4izDID/UQ2lPYl+OOlqFPYayDXaehCIC0sqG/TTotF87/Ww1X
RgggReGa2nmbPgHa6kwiM1kEb2BmwTpAvpONaC1VoOsiwc5OossVR4bY1/iE3HwO
JSP0x7k7ZB2gmQPU23NF6nz39XJZ5Y27cIZHj58Dbn/CdiYX7SSpoio0BYDbRzyQ
j6TvxKD86KhQIbozdUzUBvmQvFt37mhDXkvoq1DxGMQho/nkNt5RR32STESI1mV+
WK8FxYUE9JhCarqC10uozh08g262Xnp+RUgnlVHlDA6hSCs03Uj5XgMsmAGQMmEY
Dk/TIpNk565vQLBAXcMMRdMwehHLvO8+jkVFSNhbtr/wTXCilVleik/iO9ihQsp7
1v3WfYAn0Zcuv5/V92X6Tvw02nGugSDJ3KowplN7Zwhmzm7y/bU6nMOclonTIzVr
9i/iQ54hXyUzSXgHOjcddbQWO09dxv2PWFEh8DvPUGS76lLzp/LJtKcQ7KXSVIAZ
Yhn8EkTrEIcFz/ToeD+DtMV3LzMLBMVYoefIl4E8RC3MB1exbFwelEfPoKAZqLsd
Ok+nW6Ap090/TxMmPNTGIFqy3hEyzcCdDGzABq2rpZyJcub9L2P97xQwokwk5juu
u10lkSmnL2NVITTEMyybDNTUhpDJJDd5E40R2Sxd+r3rdG0W1tZdrAkwI3dkOw0Q
5kU7uvCM29lYwn0d+cmPAGlr4dVZjxF9K3QV8zvDIov2Wa+GhFjgDaIzED4dVJzX
K3Qqg0pG6vqsqU5oWRjNVSHsOTfLYRCSufjbNplVR10DUGWMGSdAvhOlVfkMEhhz
VUZHwGDB5BFVUXLOzcenXlv0+NMsczaYcZFlDXXWJ/qm4DfRee6pfk9Hg9oApItg
JS/ZQYAIApXytgfsI/Q+aYdTDxpPx36RqiMQe24FpBafaZcg8e7Cebil/P2uV/Q9
rinVOnheSnUsWB2+rrud/4GrLgHiNzlWmETEkS7mWF+wcaayVNoPn57dYQw4ywQJ
26rna5sM7b52aYop/iLONyAH4fmIhBzvc5sZIHnBMfmYm0hoOC2akYxsMhUt4QDX
VxBRSsFa7hoZsrF2IfDl7gYM1TvD40yyOdlW0yRzRD+wSWfoK3kMn2aHrDt37Z+1
RJ1UT/eBce/G/rmy2cVGIUutKI9Ld1DirQaTD5x+4chPAw1q8V3AGxXOSoLnoyRF
Rk4kBKChtsAzK43q3Z6eoeVEqWcJgDW34KUHVx+cmtXRMGfaL5lDXosdzD5c3JKC
X6AQyMxCjS/JZELx32+ZzmI0pE+zPMMI6SE8SH7q/GE1jCB5irzNt97Tbw8gXnnj
3/zluhDQHtNPm8af9ypHzqvo+3JVqvPHMMs3oxJ3z6zFny8GtJgdtIlnguZLZUhy
xlvVCRByry07Qo2KLqctK2vRISugkb9+5fx/8LmDGDoezNL+v20UeqftKmTwsmhh
ovZk4dqoZQ5BfCuKHuGZin+3Uw9GsTVgdMJCX8CNWszoiBrcacOzqmUra4fyzjD4
7k+nNkfGa+tsdo3Fj3+LOwk1ULTMA9DzFXfSFZArgdg6Mdha5+Mq7R7invTgC9E2
qg9hMfnsKadY3bhTXxeo3tP1u0NO1Y6MQF6Dsj+4+U1upYTn44Aqt9+JC3QyXlMr
vr482lZBGsbopBMpTpR1wg7i73vGSaHn7BNq+thB2peSj+b3bXiw7Bxbh+XMjx8v
kURZlmEQnDh4PRHh5elKJP2Q4GAb59igTgFE0tWOXZlcZYNns1/4PjCSzXU4+ncV
ZTZd8QKYx+no6s8JWTPAoDsgQD4RC0F084TeFvOmDORW4NdNGvzWl6RK3tqV+b0z
jWN7y/hMXnb+tirWslMyjdhLS0Bp7qbKAfFwEvwcc25YSqMmiizUfMXcNQEHlfrc
xgz36W7ziINeHRhi1DTSkqoRwptfk4gSnefuAsSFj7s00DWb4/ZerPTN5uqMkWD9
njzX2iDTp9m1D2HDvUtAdckk9oJwDYpwvdfqjFUt1hY+E5PCUE6qZcWWLfc2ViP7
gZV6p8Djosqy/nrOtPVJRkh2KC8yrdx8RqKPzMZORtkm1qaF1Msm1IrMS13fEe/R
H15B3AKhXSE2RXVSMaGa4aLvD5Hxp9Oan1oDm06iysp59p1KCwLoIX//nR1juCKF
vnCEDcSQVr89jftysdqbdjYGvozWEi4mGc2xKyjpqG14nehEw+gzEI7RSPs/V5Zm
XEHWxrTaRY/MaO6qb+0AjCo7HpL0gkxm0TPshbjSn2M1d2z05NvypxNMPEPRpDJz
WE3CS4GkCyM4IwlOKF2qSdDArp9bzkjO1XipQp20HYdaGTlL2JMDgVDalrOZZ2zl
JYLTKgjGZcjxEXeXWSBhYb1jigVdiaBWnH+aTYZ9erWE2l6CtTAu+LCh3dmiQx1e
83Ze4vYkn1NfROcqBKl7C0/dZUU40YqHajciEXRECaH2dWFcJ4TXhfkAQ6IyDrhR
kUpYjyruZqp4k63amainBQnC60ivncYuIgK5ACoGYbNBzF5wILimn1GfluZI1Ps0
7CkUyIZ3BUjZmXsjCkJxc2BrlzN7LMTAEee/lyQHr4/NAtf0i9ErVHVm+hXR5ypr
GgZSrXJZC8GfnklLZvvySEUX74VEHw3Cjt6YafhhbH3EH8z5Hr5mV7oHzr828DXM
RwLicyFHWvY8bDzFo7nzJzwosHWv7jjqQDlxcrp+aGZwJ8B0yidSIjfqT9BoHVbu
3jM4knnPt7MY0vYfhMOb9jvEPLKRkqxtvtFzekyqeMI91idLhPJ5nR1olxDdFkRZ
oPwSkmzamns+qdgfZFaHgbMOp8l6QCgIsa4MRcQGhHXiroDhDJZhG2hIRXZLEyF5
o/OPcKaaVUDreQyPnLYGfDN5SiwJTXYdCTZ/VBu6yVZVFaVlu8zgzaScUiAstleZ
vEzPVYT4ClqttSxRke9uvlx7IfAZySmC3oHm6SOImLVpZOLWU9U54tcXQ5X8XvWK
EOXKBAAI8ctxh6ZnVKvDsuctKD+ISGZXkzLTnsWScHS2rjGvsjPUUDUgSHEsQUBb
GsDMxVFomvhxmeF6jJNT6WrUWmkCLZqe0naiAepwIuKFc00tSAJpI1Jr26FEpZFW
qT8mbUnrQKGkF9bjuPh0VQ3oRHv3b09gcGypmFUuGU4o8YluCecmHGj8w62htQYz
Dq9E+l9wYnMgDV2FhiuMQU1Lx1Cxyf8gK5wXx+qYKZdjwYqNX0RmNO/4Kk5iuzIX
FY/d3+Ew/0AwrkRdIdVQch8YJ/xeUEYw6xaQDyAySigqv3qj2LY35SRC811JGMeZ
qT8tR2P4mWki12UDAhw6DZK3wt4Drypp+4hoDItYwtWXRM9gBDuVCeYQYa1yGV9V
7PkDwGyfTci+1DXkAK+lw/JqqQnVKKwL/6dcTICtOsVLErj5e5yyNNf0EtASkTyr
MByBcV2dKX22bZrwPOpDBBH1dio9l2vm2xyTMhNcFWtA3S828Mhngt8tJ/W5KIXH
IKcHCv6WbmF0brYcA+to3YVYrxHcqUGg1waT/Lcs3oVVbEeaj5nIHxHStAr/coQJ
P9YMoilMcLJ65M68Vt2A8anHi171KBVAlVT7zXEOppp72K8ovej361GFpcxkPwZc
l4uoBcnCAOQLi4YJvn2gJ65POsrfho7TXgTU02KC3gQNTBwmYZwRv1mMI5uA1Yw6
qsgrhfiBFcTM5/rEocDeiTWEPsptlHS52qhbDvSFVpKOOcnVlv9sZ4WBlR+fketM
Aom0cDlg1UfKIjbk0H+IYRcrsQXjqAYYJja3eAumGrLw1G4E57+ch4gMlD/sTUMe
Pl1dmgqYzuDm6+VFZDQkNtNh1Is0+bO5uks0TQTcYDuLxxIBcrvKUVvvD3omnirW
UKst6JLxDFxgxvzaiyz3lVqiKeNaR/SmV4i2PXLxAU64bsRMhrPXSkpWKBzwNvLb
FHVod53JijFmYe8SPw1494KLmBMa8IorWGidt71VOPNgoA3y0CXcDYqLu17/xeZ9
zF1JSSGhjHw8QEJ82YbGcRkgoYqJSwF6HK+FeUIN0kjLg6Qfay99zQjgPfzFywYz
WuMqgp0VZO0d5Oa1QZQSUo6MZCtTXz+eO1iCC1qrPAYqJkpcy/TRbx2zXSf4avAa
jvP7J4c+b4DNwDbE/GVO3TD0uQXpP+z9lYAxvCwwkoMfGoa91yJZfC9wiOOIih4c
Qt3LSVqmDWWVvP4eMGrFWJKmt/ZsDJ8TZeBDiNG08Rd/SvKB8YNXTwTowDJbiQ1h
iK+PNA0TabeTHxd1k8vir+5BVDbniwrH+fst+5qnvNmZjNYRN0ZzgzPjObdnlylt
avvvhnEcItmTLCPPNzWzVLRTmcwwaw6TQcEA0R3evdoaOWwUqJ6cQ/sAeOZXuOOd
ppp1kFeB9YLzOTR2quF/oFi7FHGmJM1zDCC8TPOfT9tFxi1s7KTS8Jdyu64tMN3I
G0I2N7zyxW4qo/rnGYIPjarwJRrOQuJig9oeB1f5TGxJ9Ajht4JnLs17jAZJ7miB
CCRmm58M3BpUaquTz+nOUPIifX1CnLiN2BUDMjU2nGGoleRsrkSWwkRsFvmCkOQa
TcPaWuxuvI8WeF7U0ikU6vsU2NmvMiIWmNjzSeu32rz8EnyYZtdgSVO+grI0tlbp
IxeP4EZQO3U7E4WOpKGgFUWBfjEttJ6FcWGyGa3EtSuE41ZjcjiU1EmyJ+BAET47
ZaO8ojVeJvX38NM/iHBlrKgB5Rq9jNVt2DkckFLT77tevquJHKcmj+69bsDer3a1
J69UzvmVD8PR6UFh/ffVLz45R0HHJd/YPrAuA9GoGu+62vLEuFnuKz0XYCea6JVD
T6Qkjg716CPIyXDWVOS+YdCK7H1i40doe5FxfTGMbQGX02PXAZLiUhPHwqyNJGSg
NBJOnzQ/UU9YRAK7QX2Cy2XUMv12gIVGXoLQXt9hDBZEDucji4KAgHbzgtdz4WTK
JXj9+m7qfhPGxPHcvdD1fUazk/MrefmiJ+NH2HHvxyjUxHo4F/i6yONWh9ud8zzG
wo+DD3SJlJeGXqViu15+wK7zBna7/iBhJadJmt/e2Fx9fHpwLRosKojhud/ZOX24
EYaZ5VYY6Qcy/gfyfOQEwX4p2HZaHMfZUJrAGnQJK11214IhfGUSPlnA+xMT00zc
cfoqL/gElwbyH+oiXJoze8Btc4X17sQoCiERRp31TI7COAOdE7lH8u0AbcYXegts
RPkikfGfwBfBw81bxzekiixOxGO4lb5nXQ8LN8+d+qepiCynBr/edYCa1x/m9IDr
zeSKG6dVZWroDA3lS6EAa+XYAp6INoME8O9Iz3aBXxypdkhx8ieLUFViYzngXfI9
VMeDFzOiV10uMy5F4Prz/kQ339lCKSbIXZrQJ2X5yQR06CGNS+rmtsGh4xtZ/yY0
b6n7kgRmPDa4B75cQXpI41X1gSWdWNm5lNFDEsUCVcPpIzl+WzvB8BDrc5fk8NQT
jCmwdug3mRdAqFh1mSghrNoBfc9zYEZxwxYIwFB5V8BZQ/efikAEJCySrucnai8o
3qas3Nsa5zD/M3wmJ4GuTdp9WAP6z48ZM/fP05R6+JnoNvMjoT13iFXpPlkb2AR+
A26Em1K7kuCfjYyxJ1wENq3P4+AHyaK0cTcnWRIo5nIjXXuwIDVtglEnBeJcFNqK
5q8vxuGjz6bCtxVwTbXtUrX1EG8Fh/kFE3JbzjCX+qvmlJL+3qISwEyia5jvm0TH
Gr1WWUWIVZlzdFOK0RlIFoAyEmhfCita+EJ/z5PMh0F9/Gxeu/o/CAYm9jcqz9Ca
ziDPCf7fCv2WKyoE2HldNUhfg5zp2yTxn+aMX/lgTrDautCSi6tY33z8g6S+vs97
mCeD3aYhxXSiMLF6OhAXjBCMC63eZB56VHCAclwFRVAvs9uMiaPIM9PEIMhY4Jqg
ii6U73SkwkMTT2iSY7C72Ox1Hl+3sfYszr0F8x0o29XDJoMTlCSTU01YEKDS5rAM
b8JIoxhpIpmJZ0nPjTrliReYu7Lv69hH/ZBJd09FKHM/iqcSuAAVddYXHQdL7YMt
6VGNOFIpVXFISKKdKqQ3xu3OpJTYKg+f7UaSTd14buIpsm41H2phdqdWYLdu+h0u
Citaaj1YswFmFMWcARa7dBTXJAdFOwgeqmsevWGmomwBcjj3KX0+B8UahQUyUi+j
k3XUwYrxGkK7yXtvrQOt8wbYdT62neTbLaKpCw9u6IiCYDBcvtheTftibqks3I5Z
C0i11H2CQ443TEZCfvDObJOAo9oLgmaShRQcQ2pRQ79aPonVL7VUJVW4ifOZNNy3
GIzGHpMQq3unEYnEcZgm483fIMmcktf06RMP2Q47WcOMTSVelG+iBCEPPaHYydxs
uIY9UMA1P3j/O0jPgxZ9PaNkRQeUNoQEEvT8nxtpGYcMekQioYDvSBd+LOu2GJOo
riNOoEb9gAQoI0wBjYKcnG/XpY0EcDjcdvIScQ7Ttv1c4pMJBDFDmGuxwElTRMev
+CcBFoy4lPw1ZTBISL86+wVIYCOeSCz87yihCXixummQNuTZ5Ot7yqMw5RHRcFwo
qjaZA5C0BdckaNK1lnnbu2nDsFhHPlje/4eq6LJ0tpngD5nK3YsaPBatgefYVACN
ov/nQ6Te2SMLuMSJOapczSMDBscoRg8J3UCztNZrRIOrg+HsKyHjXu0UF0Rbm4pl
PFhtaxSBRwi7u4+766hVKLl4VJxHNXqiaY2/G1Kv7kx11FNDRhFY5f6klmTyN2Ht
SLpjac5ixF6zX904iQxxuEjuQuPCW70oNKycdq+UnDgBlQOvgVp9dBYmEVKHawHC
7sL1lDuEJ12aIev+XlndIb8JUJXewFJCeibbn7B/kpde135xwAyEzPhNHLqRNorc
JWa7W8Kv1z7AJp6+fQ1SVmQk47ADzfHeUnJfemQicCtz0GRvtdwQq5rbWqFQw9nx
QHxIS5WXt9kkJXFEASH785sghYtYhz7O6TVwOoimCP4jCiIvXaq7oe4DKE8Va4Ov
sw9Ux2sgvtorEAVP06ar/BabxfCvSU4UCe9Pm0KBGXdxlhQQHUBpcGiGNvzpY6ed
k0iIg89DqBWlEckRaEJK4WM7E9EBkjsya+Tn9GwGk+n0+5CBZ1nb637TEmS8urq1
Fu0VwL9DeyxKyQuj3WlQTq7OSU8XPfDKOHgrVrtljW7g1OXL7CJLQCtmbH2ey6Z/
hR38K8WVY4jSCWs7qu58Rv5U95Dg1ftLT8wDdPNqRkWlF8pzGTM2YxW6PXus2Zs4
kXSjy0dmuSxUZu/hNtWMGF4T9Rvo4ko7aRJsoW/LilmqhsVGOXomyGeezWMsROEf
XGQ936Nzheauw6bw/KA3QhZYx0r5g0EJgnDa/ZGpllvU5jKadDDCUciRpnKQcFYT
OKCHtXp+2tfKCw3AOcSOgHfkXtCyarTrqYt6wHVkDo+HA0f9vn0RXjVpT/5wZAw3
U/s1Q9NNk0aTdRYynfKQoiZiyBkEnuexF52WiyCLO12O8e+yPLpjeEwkB7ndsfCq
b0eHsdf8nBV2qyiCAsXTCERFi36mWOJuQU087kqqz5QzWIrJLtL+wMt2FDweCWCP
dC+qP5TnUqYjL60yMHcs3Okl5IIx27he1elj424FYqWKuah7PiegQlnUVMOS6TDh
QpYUVLuWoN9lChgl5gWsbzK15ef33QqNzt/GS9rkL8b6IqXmotjVFpICxoJ7wgeg
B8JtIVLxuYsWyOMN77UAKJwxRSPTTgMwzX4n9nORsGj3LGT3szAnMOCvkxApo7+4
PRpc+4SNqP44g2YgS4XHRTWxVdA96Vedj6KTcopyy6YnSQojg4/gxmYvVz4HF9ol
r4oQQik91T6Uu02e4DCVwPEOKMphmjaKvMSU5JRQl4DjjMkzOpXlhrRwBDGPodfF
NM4DAiyQeeIHdDCIAdTsvzRzOQqMG02dHYF1i5aZHJwv1MBKGdKAImREv2C0iy/P
xeoM47aL16i7B0S2oKC3jdxfTotI9b7yAX+VIg7vzdXheWQggN7xej+AiTRJVd1U
hZNtdwFs8jMAlTF0MjK0Sw7SJUOTjcDxup+9Ua4XtaTguPN+z+68ZZNbD6SsuFh5
78hKmWy2/sZCWpv+ZGZ7BbTSdxpouZe5BNl5EvfOkTcnNImnwt7dYg9/Cp1XeWdm
TwHEde5QvWiaS6S8vgNMWPCknslHCG+5fnp7/4J8sp4G/lkSbwX+nCFZBLM3iJkP
IOwTjPY9Y/4f0KZ2/7+lD5vY95Bnkm1bobgycle3+U4CY2MBWk15yMRvlUO7jMk2
4M6pqVc77H01hyHOmSaA2JoKr60Eikg/eqLgeYzG5Y188IIMvYKCbOS+IQwIC/0w
0xgaiJfxti9LEXxcM/ShhyAifPt6UxZnNnpa5BHIMpmdXQ8mQd/2PtG/ckxcauTG
K9cKyg2OyzozfbLpofLtTDF5dC+kEoMd2hN5FtHb7/WePkeCKr7OBpYegDjdQR6z
VqXc5M4sqtx+VByvjyVFUIoamMs970TozLbNOqyxXZ6Nk60R2U/m62EjOJ1gkayi
+2JRVs2R4aPw+6KuXZz+JmvYizPIRAByma0T+4XqJYy2nMdaIELbKYSSKl6UUNV5
RuuUZGRPFpLzbpccOl63rnv3tIjZm6RemTA5yU7lx+BzksptX9TZSWzLi4rNphUn
ZFHvsIWZvse23BcFeW82fzsQMSdfsI+iPMQs5bPsDAxRCz+H3cn9jt+JRajQp7Dq
Kar4kiw2zH/0twE2sVbnc6WGov3vrimXrVTjWECpLq5idEG9NEyMjPiGwbDyjIGt
BhuQyxXeDeAbkzy5yqp59IJZDgJ+LgjSxOZWgPV/H+vwmdLZ7LsGmvKvDLl/d4gP
F+EByVdNNiJjC35u8qfdMc3p+Q3RiUrKqo6TTRhPK9pRvHUDNWZSK0+e5GM9DMAU
L1mrpw07rIoQBP74GoTZZbkRTFzMmmb4KRB3d+hTVJSFqnr6DWWbkB2f48paZWJ1
qCiAMf23lqVFJnbW5ncozvlXnVYZY8hXOTmFl5tYEjN8YDbe9z4nCfex5towcLCS
MxRwkkCSHuuD3OKcemiM0FVEhTjICEYY8y7BMxXVyUo67/2lrR4SGQGWDDorkAKK
8x5af/nGTCNnwduCbGBzH15V4Ww+GGh0M7NhPfXZsih1O2a5XVMxv7zwNs7+/CKf
wHI5YIjQqxqpYtX7Po0RqsHqmdxe94rwBxZt+QLIVystoyXAZ1hOcBKnvC1V9U8A
PcaKWfLfJ0aD1RSLaD3Uz7MfHwM56wG2PWFXprXkc4gXm+4YkxTeKDM+H+PYCSjk
mnxJG3SHe/3PgyVoBobd+b+u7Dw8C+2MOfNdcBjQxrWdz/bkSBIpZQZxgaYsyqMj
blGcNf4/eXuK8kxMTYoRB6w2ez8S46HzqHswov7Vlee57RqDJ7BQv7I+7pfClhty
mbqufqs/ZJRl5K+mF90dHdV36O0qrVMKqZcPNNDGWqzMfMP6J3607u8YAgZP/YDB
zOYDrdp7RUTMemNJSyM1ixkdho9S9tMBf7JQz4BQ4Ukqy8koVqANnZQLyO80Jtof
tyh+M13eOTtVrE1kHsJpqIyiTFL3X/lQ6Ent1vxpXqsYOPBb68njmMX+HITNLiQT
j9on08cLT16EuQ20+sccusimXcMrTqYRKncPEOTrFwytvdR/RAPz4Hdb5QPVK3vX
aUeIj3RKQ3dV3P0FBdtSbObetFcAPC0FFmR3J66tTV4b8REwKp9p2ZTUgjE1eW6t
EdMEImjbCvvnLhcMQkQwWSKbTlVTNppZPsAb8+aePEYQZtcPfOD+DX3qXZiV3IUz
oUtvmRJ+r0GFHVcquQUzjlI0zIxxYbI1RBg4dbDJ5FLbH078TSTwFgJLDPqqqFpK
LUPyJ3CJTpecfb82Axd5sEJuVykoBaKyv72VPa6NSjrmZ8KMpFZbjsv57zCzsJW+
x2zU8q2McwsQar4H0N4+RdANTZBMxp9f7H3fA13jCE8tlR0R7bkBzdIYIhWyY3Kt
3Ah6rS1M+m46Ih636uDl0CK/twkE+f5MjBfWpeTxC1/vq+o54pjeRU3RIjlzwhfW
TWxkLG8jq+cKeGOfrVjCaed4X8v6Jr5gpaBXFX1f2Fxc5aFtYmAVykO3Ml18zHxI
PWpQ8Ug3YiYN1zryaar3r7GRiBaHj1G85pEzptkHN0ViW/N/O1O+OXBm8W7RQy9s
xcBtP5TIiyZGTbcsx0mq5UXx0AMBJW912IUjwJJ2sXQJId12ag+pUG8bpkiwObAF
RQKwnhdLguuzGc4wnl1Ur/zahRcVT0AbRMyjxUPCAR/vpkLmjQzEDYy4M3PaU5B2
+ptYi2bw0A3h4fkBqhS8RDET+d9K4V5IDPPqXE+Bjj2D2KtNjnGBXZb/3T4DvIeo
xomXEVAQu4fEr28livF5UZoZsRLiVmVWgenvs6vmyqZRGjV9ZjUpqOLiI/9FyOFT
bVmqpnF22YucYkECa6ncyRoSHFhxIj1OkUmesocY2SN//EL4sBl/hBg8D5kI360H
RuLgEyhGDbCmln7fVrbvi1VX++86maEQweOVZSMG25ASApQOzYcHjCOXfvPaH0Us
XTxSLxLNROrLT/3FAu8JlTThNjrm3SIg/XwYlRN5w0W9u0ZL+qVvnEQdAa39jBli
gg20pysbLfus85+HugYSDDDCcyyBvZTwGPx5AIvjK4hVNliuXhOUqoOxkwVRejhW
RuyuLgzLk8dNHbyrpUNTSmISFTZDpcb61MEeJJY9CftbgF5ZBPb11b6ah+TkX1iU
fhkhZAzba8WhX9YoF0iEMfwQQDlv3OKEuUmkpKaPhuyELo96rZvQLOGekTziiILy
Aewmw4a3GvQx0mfYIHXhXJ0WgxdT6Vnu0kHS/KUZkhyjKmAnqs+cB6SasDAjEJNE
tG1mh/Rgwi8qEm4RslPlsR+oGUZw+eAGayh/uHSVTDN1GpPRSeQKSqL6VSBvXKqz
fXxZz7GiXmytGugF93xQDLkxT3FClkSScB+Ts35xfpnFq6wcIlyDb/l2rIDi59ps
XHfP4th1bJDHwQwcoyB6i3wMo3qUzjEgesj+phEdfkqRici1B8TnVnMecJZGsRHd
LRp1OKT3c7i3lOsQOQZkdQUoZIMUD+iH3vSnr0Vf50FkBqUJh0z8f9gJo5W/tAs4
Z7Zjn9XLkRVq6TCgcCHtnth6bAb1ByYcvM/XO00r49m3aPGX3b/+VMGg50ld6DDA
PG2LyN5DWcGeyCQJ3Ml8C2S/vT+yoR011donCTFlYw7bn6/Zx5MQ9CZgl5R8VTle
yDNemwX6crX1IDGVwkvDTj+uhWrRmqe16qTvwA1XZqCSSa4DrUbAf8IRi4fSKZgq
RvJ/DZ9ZIuHed3mklsHrL1MVLUl6ACBWFVGhNQNBGyPHAzcZ7cGQbhNeRQdFhNLu
AQDRxzLviVtgSHZd4U5Dn7/QLrHagq/OEX/EUwk8ch5dpZMp/gKoaQuRMC6fOiNN
bIjDqb0D5SIVUFviU3tSGKbCK5niJdLQTZScuEJzieYYYaqKoseimGHC7f9VnsxQ
ywxlStzOWUBRwTTbB0a9AXMCGLPk2E8ei+WKHN1kFmGXlqiocsVx+hJB6vI4hhpL
FW7r2S3cFFDA4pPUF1EatMAAL1f2Vut9pB/QnbPWywe6PHl1tnNuxFmmgbZ8kq2X
mmjgFOCpJKTtewh/wD+eUfuvMjOj77nO1eGYEVBPml3etx4+0iXXhlhJpxrcr+6o
+0GUFA//52FXMkjRt+wM9FjoYaCAhm1HDtv90UyC2OsNzS+G8iQ8d7TRYsRwv79D
+PlyuxuTkV/bHhA1u1+sRMq4yxtov1G+T/NWPrEe9wWElSn8za3Un7aPh5NhCTjL
GAoTkjDD0RONdwlvd0OBd+Bl/o10i42/Hdbdy45PKj0Tn0+xgkcV54X5PtLp/MX6
cCJSPLVKkmUkLMRUEf79L5zOaKi0Qp0Igmtr1VvO93mET9hUrBLb5UTcYcS6R80d
eTRhn+eNRNf+c1xTs5S3XCLSDqKgj7RmBKKShYyoOKv9MMNlxx42kr+27JAGF0dj
gsPeCYrZiWTa01tIfS330OrxVwiHZ6Em5+hZtdOnV3HdvY7u2lfaxP8wSm4gPfzs
tikHwW28XDdC42lESdEnL6Ie6TP+4ET6ZWoNLLkhmp3kdXLfwMkZ2Twgvr5Icb0x
Rbl7F0UaIokvw4t0d+CU5mIyCfjqrI9/lEuIGz2n8tVC1DFw77MlYTQKxVBTnnki
AKS0Lmk7Of6YZDVYnQsZA1c9ttRkVWKIFQzElRyYzCyIIXUqhMl4skt4O437Nvfi
uInDihGBbfbX8OFEpuH/WxoyCegJotIIyyivjFPhlh0iFs8X5C9/5EL18Xd+LiPh
meVG2fkKwEK5btQtUTJCN9RQ3r6mTkqZP2GNOm6AOe9yMsIGUfO9EtQW0YK5r4oq
hkyJ2FhTEUIjV5erAqR9AHfXjCk6S1zCZhJuR+9ogVX4hmt6a2iQGsDe3RypB6/x
j0b091vV3Z7IK8tRXCD7/wjQwiIRGCfsShrgOFRklGfVK0+VRIln/F0o8Jj4sMK5
w80iG3GnOXfkkGlsbGMPf+KQ6Y8NmGMWrRRbPnJZD4ZRJ73v1rvWDDiYrbDoVdDC
90E22PYbli2vC5lHZni6p+Al4aAh4BT4opza4G6seK65ecjHWqBXP9VM/KoH57oC
UY4qzGB11I3U+DddqrfuHcfHMUGOfjJ3kp6S+tktFk91vJZap45zAE9JNxbIn2ww
C2iienmqd0n79TR8GVlLIkkbTsUTEJGsFr0/ZRhqHDHiz0lxLs6ttnFqauRd+nuX
t+tUByZ/ob9BIvBUB59nDZfxlp5k30k4H7giUQwADqlmW8/MmZby9YE6UFUEbXsv
7yLMAoVv0rDthmoizB8yxlR5VWlIqhyud8ja25Vb/6emNNUpfswhjFV6SOFWe+iE
lBOfyv4JuRFtzfmTiXZ+irQV1MzFug8iOK01fFIedhahdp8koXru2oHsyz2Rh+wM
KKKLSJGY10tZRLUbAefxVv1cupW6PT4iaSAPLQP5FQeT15EWdCuHB6Y0gK0o7gDL
1w8aquvo0+FcDFRgaxphcltASYIEdgGKNCwY92Xcrth8YzbGMv4qrrrkpdat45iM
1S03dzWsNx8VrKNsUt/dBHCLHFgw63L078DB/dF957TuygUlITmjIKUTJ+pwa9xJ
xRANNOvDFGNq1xHaZHLQ771wNwm6Wqmm3hYigqn1Iqx3bQYK3VGoZxOL54516b0r
GQZjin59UgoGfutSoF7R1UmcQsOZ+0pfDLtueSOg2yWoF+yKYeBXakZ/teh66CJl
1JbNRChRTaoJruqmduj/OACW9QNIdVi2T0HUlhT6ciFtvatgn9zXv53W9IVxw3VG
HsLz4cceqBYvHZN3VykiC2m9kiCxqaevxzAKIztgt2wxgHPH4Mq9JKDItKpI2JrO
DdVZeZMGLZYrVvcMv4RxfhvvEGdcnFedq1qQZlTcJfDdMxRqmQ/irFOYQ9iOUY37
8k6ge7d9N2ERhFHHh8erUeDGzve83JlwG01vk8bYvUjmCB7sTYQVwj4+Ey+tMIU6
luvXNwIFina8pHQoCUGrNBNbIvfqzsAOn8IU7q1hduXSowxfWU7fPxrVt7+aLwJo
CicBm4xRN78Rj/fqJs+Iw8QLlzIy6kujz/Ne2uepfKxnYSgxgOGuDwClAjpw3fB2
CvlqyXOQmqCcUFZO3aaaanaX18kwfPbuTDJK0ejRHFLffHhWPABAY9uRaebmmicc
GO7Dj5HxjGfoTHcP2+b29umHJ7qUvH4EjL0goQK3XnU9zq7mf4Le4llPUn5QpdYF
xWjWBmwI7LdcfgAicr0ouGkLapMuZpgldoPDtkeBtl/irXLyDGaanBmm+EH4KKsP
L8hGl4nlCy+X02r4ZpAS2dqh4RVlrToDjpiALFzfsJg708AUCBJk6iX9Xf5fi4P7
qOgbmeHEduC/XEyw0aqCsy2FueDAQ/UJSmf3oC/sVApXwu4pjqJZK+kFPZq8xRh3
EQZSrczEeBPWuyLM644HjzlWvsLPLy+CcjcSRo2L7xez3I3vHD4Njg++IiaZhr2g
eH8dM6v9DxKqO7TB2B4t9X3EF9Q1x28imCBHnORNwXc2qg9ikPd6qRqTOAXRUUJU
gOO9I4/nuIno11lbDRVd2d7G8Qp1Tp94T4BtqQ3W2eOfG3ySgcc2rXqgJd93lROL
Xl7tXe4EV0AP2ywvssquakPyeIxLwubKJXpvI/+9vXRZqCFFcqeomokY1ogQbMbT
CYc/UGsn11EVBTHToYpMe1dnk0V8V/0f84jlj7yw1JzB/h8NihdHEdGHBRdBoE7k
+MKj/miwzJq4zjmmdpVNhyRv7jB8XdbwVhxPuca1s+rXHa0twBwAKbs71EvMyGua
R1x7JvjUjK8bGICTNZ2/6fn2V2+jx4oQrK5a/cPX6cSfyxvhgx+Dp9/ccdx86nD4
tgxHCUO3aI0uu/k6ab3ExzcWDFG4qD8wpCo6Y0HbORYnPwHybvBfsePNU6OOkpVh
obCtiqLS1r98zEe0glvHhZV9LFBTLoZfRHa7TZ3+jpIV3OB04LvinhZ4pQrP5X/x
ikWwgA4TjC9V5OfptfmHootmQXBFbPQTaUEZZIPgbwIPA/RNUu1CZV6ZUsdl27Mo
KQivQRFn+hChXghpH+zIULKqdFB/m9mPwOp+xiN3ib1YuS9jF0sFZTS2LdyLgEuU
mNKr7mYQ2Jf7U1pNP+STWZ0VOtoZw7RumyYUkH1rVNfwK+3SPEKFsu0J88KdJVXe
EH6PPyYOTHNMXJTzCXYh9UKvlVvUU2mu9QIek548SNmas25IzWzjsli8POvuasIL
r9COn1OnEr5IDi/KDcNFwt7bIUfnlYJ6d6zPTuTgs54kI1vQ0YdZoUboc/6DdtkC
CpeqF8fybLFIH2uct1IgdmxQP2rwd3z5viXixlBAr5qpXOn9onHWG9ZjaRF7DFcI
qeBCwMOu+SPUn8JJnnzKm/20fAVo/yxEM796JoOzL9bWjWANqmm7Q2MLsUyNVm88
+9oosSLf01Ncj3QmAACH3fOiNwEswcFluDCooNN+NG7VQj9xFo0AXaD1jlkW0kEY
uM3FVk8N8hsJowprDWBaro/gsCxnvCAjAqYiXXnZZXJTtt01y6i+3lUO5300aKrD
OzI85PDQEi2QXErDX6t4kkrMwFxfm4reYCrzxJYJvxaIYYE85vBNjcL2cBaIKjoY
rzNZAhGb0evImxEk3KoKAIwBS13kpZswd+pZ+wFW+2y+1Ttkhoh47+wH4PKTDfxE
e+wRJrxqrG8Zp6GeKTas30keqBt8SnKdmiKk8Xbq3Whlj9jd5iL+COzeTw5fybUQ
l/dkLq/BLfiwnCnMzmgdJMDwEih931yVN0iGMjmb4Q7M0fT41vGVfCOPQAQMpLVU
pgCu7KcvjA2swPZ3O3IiZTmsXZA9b/Tv9CmaZSBzkMDBmRL4pyS0Tr4QOO1c2CZW
5CgLxsS5lpx5vx+gwgrPZjXjzoBww32kB6aWqNyJxOI+BOWh82ZCku2mjiGxN59B
gEYjUz+MUsKWvGnltu9VrWb5Hf3Q8CZjyGYpDWvufk3etqO9K7xF/w5QS6ny3mog
0S0iluz95FSSMzIu+3k1009oauRHEgx4Ehe3Cj3quUf4C+IF3sOhtlGH5q6Vxihg
D/tkyWlw/AB7mUz4dqWA7jND0a7mkACXoGSR/xLfNZfTQfX/GWmU3jKGbdwPnVmT
qQLYDGT7JuKE8gLb/M08FAn4XceAryDVMVmzYt+17bMOTV374jMLbWTauxVfG1jS
hAgn1D/4GqNYRjil9LRLGBAHQJMzwGe2khtUeKDnfSvf3NTuRc8dbGhUCtdoLtHv
JhKolPoFHETdXjskjn8dPBO6dC4aZagKV1iKAWl3TwRLPyFoy9XGk4xWQ+p6eg+C
iFnih9xcIHZtteZ4BkOXlSFzxNd/t716J8fD76ZltwO6Ty6E0wnLSQx1c2lQUNSt
V5ptCgV9T14xL603v3uBzpefq6ELo0cJK24KUYSfJw1XodOm1K7i6xocbifyPH//
W1puPNnX0jGUAp0fYoSd/1us6WbMxF4St+/KFnqaNkarc5Wgcqe5yU9Hool5IKGy
Pu8mty2GUUNLkRYn4KFbANEvnV+lFAG51jGnffImPd7U1eITSz+MzWtYFyHth0an
QQq0aIYLIKCeg8cInmT5t4jbAX3WNQ5701a9v7+6kC/t86wA6PCtu+78MicAdyy7
8cAulFYeAgVni0dXrkuIuAFXpvf4Wt8PjQcFNDDcaJEFEk3JA09I0O4LOKpF3Q0O
mwHdBPxuV51Ti3rcbiydeOQA6JERaXQgMJfN2jX6CYlbskvvMrzoqwnErKo6VsKI
cebmYufusyETDgZOoAl3P2Plv7dBb+0FcHOS53TdKLAVu+MmyMB6L1onOxLHz8NO
LFd0zKPUZisjiYqew+0W+ozz2bbbw2TChm0O1KgWTmTKwP7/jI98HNXGBBn/FL26
Lx9c+eR2lpR3KH4Bp6Uol6mQDq3276HprFSfPgL2Lolhc8KVCyfEY9eLFK5BijQK
lHzl6WZ/K16Meu9llnP5dy4pIPW3wK5qg8mYy7iS2su3iHn0SbPkAgGnErJgUR2Y
3XWwYBRr8xWXRpxneDmacTG4I9JPMOs1KxPOeKS7Kh4cpQXY5QLThUl7DgTcfpLr
ohEuB7B0lK4tB1/EihzhoWfgNvjS7MBZ8tpDvAedhLw8Bqw3WKmotxzsSppOgaHh
09pNErHV9y7IfVwy50Xnysrm62TaLeyu/MiW9cKzA0HhCHygPkmIXfbQJXBwmOWb
AH73iKaEYqSQsPNJhQJJmsSSH6NcT44C7kyIBBPAis80n/fwov2lfEvfhdihSIBv
KJXGes3uhsyGLCmeZh8Vs0Y2l8QiU5qj2vhyQMb+BoaBY78j6zHoCO8VAclK9YTh
cqjpZ06roKj3C2C/CQ1zAjpCjo5b3911Bic9J9y5w3tn/u7/a+CTyu4XWqX9WekM
22ZB2oLT/LIGlkXFZTQJTH8O57/gPI2Ra4XR0MIgTVqrN1E28Nf2Bm4u9CVNqFaM
GhIOTuPeU2Lm4lOx+lP/pAFPxfUizL66x78b73ZEv+QrzhIpQf7EG8p5iuFiJdVB
8HV1dM2A2KE+74lmmJCwN0awc/ko4lSKteMoZRIAkVpUvN+wKC6zWXj79gW14+os
j+O3uFW+QyqWGz880n6LFv5GLAfFRVWBExAhiFVUqn/u5l8zSMmL/vrZwOBnUyeL
wxw9CTHUoQ4d1uLHeDdZgIaUnL/TvWKekf2M1YmJvBquuuSRX/1MftldQOdeBtvJ
10+GLPzoV72CWa/J7IfPvz0GsUlrf3/hCFV1XRNxPlGNZthj+vDOPt52Lgtb32t4
xVs7HDHFxO2ItlZ+soIeNRzTHTFp9LGHlnubXdPANzZlyMnVWhpKlz/QkVuWWxEb
a3XeTajllcqEVvEoH2Ji9xiMF7tjObrsfALKBSg8Q8JEqjkXe+mSDgioebDtC2G5
H/8oDa8e5vZKsAnbNsreNU8+KSaXBN4PaOtvwYQUDE4kUNSzex0M+tjTA8OnwoEH
776jSO1bQME4Nh+dCzotDNU+maOxbCJ/lIsw/S6WlQpOsVaqEaDnTL5czenUz/1q
8rIiC6allTOY5RIgoXT8Vudzdesj/k18h88fl03LKeLpyn4erPBFh3vpHNrmbpiD
0iTqn2jsnoI/hBxPIl6rrCUDfZNcKGsPrOEuOtj3TMCZ/igvPaKoY1xYEnUyVEQB
qzXm/wtedfIYcNKTno/uoe0gOfRa1qL3GRdjCYWe3bjm6AJo5acMpqEv0seyW/zu
6dH3QvvU9HfI6GN5EzGMc+DM+1hXGW0Hx8cSsw5VBQ/unsTjzZtHVv4zoPtLRqkq
qYfjKzk0W8rrn2Mkvj6HKk1xbgVidTcQsvDDG6KM5Twd2Q7dMQwxfHAhOJvUW0g6
k7uXmy6pY2kZdFMmbvIGMMrFatFIoWCe3p4b7hVKpJMSfBY2sGEkNP904TIMmaoz
BeDfbAJ+5rQupnW9sT2iz2V23TLPs4XWH28qaUf189yU+kmw6CcPvfm+P921vdbb
pbhO24UOcW4AkBYrEFZpH7CulxZPeMe4zybHglszuQmPPLM16jYpi5sZO7vvyiJ2
jJH5bKDHl4dzD9xBl44wd98ZJg0XoJDYhaVbmnxRO9JXYtgu/qrDtaGFbPYuc5RI
RHfs/YA63tzSbVFH3sHL/fVe7VI23cliC44UKcElzle1Ex2kGODhwQgjHUhrbTKC
BwN4AFI4iKvlbcLeNek5HzY/D1WAR7Z+Uzm4pWiGhuzlutIJZLN+5+8IU954RoGQ
aCGPE5SSz0B4JFHsojmlPOvrRt6S1RGUGbRF8fyCgk32cyKAJyaepiJA2HlgFmlG
b0Yzye/IvVLeBkhk2Wzw4aJ73Bz5XFnv5+sozfoYvRHsPnfLCIGRW8WV6QpVilAW
E4ZOmV77FTMVGHI7Qa/b+OEsq6mm2KZ5N/oUpY3qANDxBiUOzYlAJxkZAyYlGJwE
FCj8N/YE1qT9VV3ufVrnO4jKiAtgGcuEL9FXpnXYpypZmzmH5IrkJiV4goEeW2wZ
eziUvQTftw7TLJRyHigPwR3PXXL8jcLfwymM2uZejg4RE6xJ4/ibUvSd5W6sEMQI
rggdAb1OdR6n8LgjutOg2HYzAI2sEgSxQefyQA74KqqAfDxeRVJ8l4jb0H8vJNvk
BsJt7LG0FV3jALVNuXdIAdRmjDJ16X4P+M4oLMhjimQRploFWRUTX4fLL671Cw7Q
OyiJrQtQDE3ZzwWtBn0O4+r6h9FQRceKkn6/ljgsb6m2praiNQ43XTLrmOS/WENN
abpJcc13uODAjVqD4vAzulEiqDAd4oBMQBxfWgnIEIHBdKPjY1s5g61QI1JgS/1l
OrlvB7sIzZIUzLj43hxncMmv1IyB+F5eicEuAmtEVc2qWit/TZwBrzU2iOZBIkT5
cwk84fyD8sXpCQ+DpmPA7fSsAYUuPSTWBRtC+lFufFmARyPXXvM7L/HNe9U1qQsF
cphY+6IY5LT9Jcn32Rm6gKlLp2G3hOgQHBS1KjIDj3+7Zqu2f7EsXyrC1dC6hpjM
uVrkHkaG3JLaLz354pruut+2o6CjfkDTPv5PMtaD2wpSS0rqKp46n0HOMreoSw/L
KMOxMVAgm0uJqJBfxAa/qbfTPAizm3uUP+O3V38O26QcUrCIwupCffdoVCbPABur
2obQrVqbN884TJWJe8s3RmbcsxLwj7ZOVl2DRZF9H6+iO90jGlLNHvZ/AmZIUXgQ
aiHee+W2240GWiZr9KoqrU1sRkrw1l7JiEbhyBwStJDByAErPO7uORSPSnVtF9Gq
HSuLXzUTNBVqXjaBnz2UTpfn9R6eeTicVBEUXaGK8dfiCY41EnBL2qyPFo7TYKn9
lAG/+rZdf1CfInhBXewe158JALARTsBbTEGkg3iNRiN/EsbiQe8Tj/BlmZeXu0l5
YCLRKT3U36ZsvAGOKcM+b+2Hwa7vnscpN4gl12e4gkOSgY2GqaUeVo27+RYGFNiN
JdxAVOH156hahrLdka14rqjbk2dR0niFmxWn/mwD85ok/Wj/5MLf+Fmju75uEEdx
Mlv4aV2ZDJjqzjU+tjFgGQtl/HwIxatz+QEa7ac+vl3vu0jaU7bHYzbbBod+R4Iv
OW1ZKl9ZqVuTahIvXisI/Z39byNoGS2H9PmWNsadOu200yffO3AOnkESOhbUG5Dr
/BbCggzoHN9rfvIKUVbncixmNikvkrAyZ7ceLyoXs6OLK+6U+hocL0yXKVoTiCLf
hPLMPm+iJzsyL3Z2O10PPlYVB5qytgu0hjTSoDOOTV60P4YKfF9zRs8wkNScu3LN
/zigajs+f0UtiiXyDVddcX04Bn7mWufXc9tfOzKe6JX8IVQ0vTNUcaQ0uJ4xdhk/
YUtFRkmrtGaks+G+6mcSkr6+xKSGMJNgBUT4S/h30w3qfqzvUFcpDdPyHnDHVIJV
AnTjSuIuKnho2YZitxN96IiIS6BkICRUmmz+j7IBkXekWZMYThWvqQyqDsjD+5Xn
vXrC0mt0daBG4LLGnIFzyemcE+heLOxJeihcQEwMVkMa0Yvjnql4fhDqgcZoxe5I
ebOLbQunJOe/rZ0lYtlrjTHFgqlW4od1FL0aN1DgxeI2WgG4Yz5UofTrgpvdZ8Vd
IljXlw4GDC5jOnqQTKm252gDF0Qo4rJUgGoaZT9sT13SI6dTqXwbXS3j2gTLhlq9
wBYuz9oRK50032+oHA5S83vBg1lkCxUtPD/wQ3Q+EoPMdrZYE4fE3TLiapIgZwiL
yS1CLbm0FJnYELZLKMWTMvQod/nwotBRrSrD1FPpK7dbvKCFeY7nmvbg4u99LCfb
6M1kIgM3QXTqIM8JwezpEdsHGVs3VteY3sCY0A0+8szkfEOxG5o1nAnUij5MEJM+
KY1KxokFHH9y5bbtG4bM2zghKaYwbevRp+haAPldkIfJqBhmTR7phJZTX/NNogm+
HP7Ie71woZh+cPvrS2tW37JQ7Ql3HJjOPp668R9TyFtIcBZOjoJsDyG8hM13D+88
hmwS/BYnA5bHnEK77AtLI7Fk8d+2DIxKx1aPWQvItnfwCTZz7rN+L5Kq1qHfZfAB
nCCEWRwccBhdxjLKy2hMuS26yb7ygtql37C4usI9kSeBP29r6KAJxHOAU7XXNcDp
tfquqalsdyVYCA1wzuZOB0rRQ/hgvoX4HOaCf/ncB81i008cUOQrtWdzjbfcxXev
/1xmBXfMjYxzSiaN0MuWF8589MeBTlqIuYyvrQ99ff1Bi5EMJaXGdpfYV74CFsLu
0VHh3YV7VVcjqXzZSLjFag8oKthyGlarredz0gPnobR1ogxxxQJAp45GTwt2uhQk
+uGAPAn36EpS7xUTYJvLpkiLR+Pb/aheQW+gCpXgggHxT0eTnglfeA1FK0EcCfra
7gHxX7rpxKS32P6PxilwDt6hcEcdzjsRjcPK2sHfLurCMsWMGGVVLHeTzvhShrH3
6wYExQe6KOv/qwaMzaRGj6X+Q4aahyo09vL3jOq27uHAPd9qw8smT4AV5+1QH+qe
rX5h3UE/mS61bcHH4N/UxufXheEaqXCY1qFOiGEVTYeiE1AMiiouv0GylDBOOCPO
RBE5dFQJTz/fQjnrmxh9el5oi0mplc0u2kDPm2sTnImaYndZnniIa7aot+vWb0XB
91cCsc26d78L9YY+048GG8o0XKyzKaeoOtbbRXsASABAh+mk/xuy0uulNheel9ga
jf2mT+36ZyCizxegNa4LY+073dx/snVbusZDLTR/44esfQij0jADdBDTDiXp6aTQ
mETBT0nTEBLSJLy8/OQjMGPcbixioJVEjqtQkW0YIpbr5E35mt4rqhVlDdl0A777
+Oo6sTMATH9S7YW7Lhufnw8FYhP+ZaA82linF+6ERoHcpNDaq7Ek61t73zB1AjyB
slznm1NgpewVy64PF7Y4vXxXCNMwKVcmo6OdSmOcevS/+BC+gBQoAg/K6eHqORHt
KzZCar9kM63l004qaC+KN73taCJ2qgNSZ0ATDlSeAevYCV1OcFnuZCnUmjMPjrFd
biNDCKACzdVKLGHval8ayHcbMglStyv6Ngn/61TMXTm9rV3ObZzw5tFlyomCpJ5o
J8zIGQTp1qQW6+EHDl1Q0LtiHb9omCp5WJPiyJs5fWVDXMUY956z7Zq/wQop6z3V
Ep0iKDgcBtjMNF4Cv7Hclr62F/jfjg3KzqfK7ATWw7HCmfGhNiv6eLmPENjMrB5W
Uvbkbmg09+q2g0GO/uJ9c5IDrbCQr+0bedmzf3CrI7u321HGFgrBr+tkW+LZ+INq
nv1saEYxSW3PxtRMypojyaWvsVSgNr6IlAT9AjPtHQ/3NbDBVSUYWWZHnrlWegia
xRrwAPHD7IU6SGpAy6YatQSmji2xLm+rESwCNkU3sSjo04/5HtwsZfYx+O21fiza
hH7FTwagAx4yJH5ZliF7SOXCiDHvZRe+QKjBrqcsfGvkvCR8lG3rVfL2n5E6xBJk
2nPf0hWj4k4jpOsdo2ftaCtISLTFeNeb0Z8Cb2zncE4+FLy7IEoLEE+Qb4RxNclA
Ky2Odpfcc4Pz3VYGJUs1RpsTBjuoxidQ1vSVMQhrMMb6Wwf0y3PAL8kOnhT5jzpN
IlinP+BE03OL7JmLyRLGDM/n1TgBKnVWZy+XTSDP4P584G6x853YgHx9kZD8x3MF
JqBtcJyiVEq1lZ9EvyTblkEbNpJHdlggomARmLYxkF3jjr1s73Kiy29d5tCiDZvX
hGLdyS/TMzt4GhKUl9e93EpeeitQ6u4ziSvgKz040Ex21tsPMbrt4bQgqy1npl1E
3SPRBCVMmpFPh7FVt4PzBsT2tHtP3kmddOKjUAP97xfVo07LFJLnyxIwr4XRaqmI
N9XSKI6GRl20fe6wHTBJRh4X+DYvbCXJ7PH8kumhKBWI1jNi6QCG/CRoOO/MHMjT
kiJ70u1VwZp/G5/KoweCjpGsuqvRfmiGTkYcJMLVf1k1I8j/qgBS7r1Fety+oWQj
hMrOrDQivxUPjC6mlh6HCT42JRDSMU3XbtKQRk4HQl8SndrGk1Dm0h5lRQRYlp9K
plWBBhBT0PmFhgsmxGT1/cEJoWRxEcscigNNa9Sv313DgncsplwFxc444Gm+bS7Q
nns7ThHUkGgyDyqoRGQWzbc41DKmdyaG4VvVfz1Sf82x+lOcRqxzK7c2bxWlwzo1
9pHv3MyHTDRjIoVzJyhdxKCg+RXnHRb3Nic6PY7lACfKw+nW2W1eI+kWS1ap+Ned
Euo7qEIZ5vZVgbrvKGzByDa0cgs22qafljboGzi40Med1J0OZl9KXKXFc27kGmaq
1EKP+t8jnTenoAvpQsBpsUBOKHQ0CMe55U5lHl4ZIPfxeXFCFxmrVFACk0RNn0gg
NOq8IHnQQWkxoNAb8EibC7ZWinIObCBNxNrq05yoZtH/+uoxbrYlGOLArELJjdFZ
lWSvDxSQDpjjbb/ShdCq0hZm8rJCdiNNw0Eo8NzBXaV7d/X8esnoBkAl5sd+2Mwj
LjFYOJblmK5qYFlp8EiIh0CZqgf6sAuQ6NmIuJJItoVu7s1h8nBKxFoEJLLNICfd
6Sig3j3/sTdgjOcUy+yv2DkixA4Y87qh604eECoWcJ9zx52QxHexZOPeB9RfoZmH
IVFwEQJjT8sy9GN02xg+kHXI9kU05AI2FCaa0QgDp+XxwcRzE6Q7usGPDS+aeZEB
o/545vy3t6C5HpJaGyw5joOXgOE3mmhPvkOybUczw4/JyO1rzZ+N70mmvqS0F0qM
BY0zLTh55YcZg9OGc4YHDsXOCtuU+i1mIUifQsbABNSdNbD2CD5PMnhVC7R/46AP
lEwzFjOo/29FDelyjfoU7WuwigfKuSJbWNdfMbOWfSvmv6g/gkpjFFOb/Bnxlicx
6vZOKRm8CdxVQ+9gbhtckNmPaDycMhzVLeVlMlYsBPbCp6x15JjsEN1oBn045lVC
lTIv/lw0oIgSd4l3/T8DKMXIoLVlpaaqiO36uFydnORlYmTe0AdMnlHM7rL4Qyhw
NcNzGyk8u+1gJAW9rF0W8ve3MyAxc3Va2ZNmNs1gM7xOnx4/85YyhAQV4QtV8Hti
OjBqlsuf9iXtRVjOfJgFPHh7LT40zPWh9/kTHgIrUGlQiowaH9CniaEntZp21FwP
T1pv3W9T5DQftf910gF7VTtlmShisTJ2+PJVaG/LjZ6eaDDVxUV8161qB+jiFhHg
EyiHwHUWCk42ARH8mRLCjU980qRKh94JJ3/7JU1kQJaiXHhqwQe119Ddlb7jOt2z
PsbUkzkEhkN1gfMgYlfw0pJSDTjG1LbYdEyxyU1vEMxsxkQYrYm7zBiE24ztie0c
9yX4oGcYSG6KM7kyvQ6hiqXwtttronIPphinAnu0jkr+Rqp4NlI95Z7L6+Tw5eo7
mFoVmc1xarrzkGtETQb1V/QyRnD/5RI/OfonDtzEFDh74LnUc9IUP8lCnEyJcNXD
/f0X2mIN0jZ8FIn7KI+l8l1s/cp8vXnYeNkflA5CObzSzRaUUoR+Kmo2onQeswCl
9qldBwqleM/IbKM8UC0z2BeHvB9nYIhSp3pfj5DsegrgcFAOJJ78PWSwjNZ5jZ6p
n+AG2CWeg6cZ2K0R8E61ttqjoF+xgEsUaz7EDacAld1thZgbkWtUc7FMslpyV/4D
yddNSQRuIyJC3nuVq/ZGZ7wRI+uCOv4zcFK5OJ1LwzLmgCKSnZOc5vR/RksVl7ES
XObx/6qWhCM2mP7T9qKYMmyLOkoptgX63625wppKhHUN7RDpkpJooVfEWF0hZ9sq
6nKwD9GmMFlro3esK5ef0cWYOB5dB2ngTE67hj8vHqIFtxyINbOz0FPqB16/xvn+
ei4UBSSk2bLrmxed+7APUw+I4+Mr2MLceOtn1TApQ0j/cpD70AQkSSrvIFLlgyL6
PEhfHY4gKwQH4ITl7BjV0BDymdZWY6YtYskHv0RFzpSKzJC7960+WfFO4LRmRtTt
DHZHZf+MXCMvsaMJ3hoWbrvaGotcNO9ZDbMaAWz3/Ze857x14ES/HhCHPjHEQ5nO
6EMySCOG2zfhUVG86VqlXU5P5iYLKNK7eAEUJrbxRlW46p+f8DqmJR60C8RwUzUo
aKjwZy+LY4+Gr1d82KqLemN4G0PdOD3wyH35qnZ4o+kUADkDvh7OYzXEyGJnmBlT
BvbKw3lV8juAhSJmIKXAD+16fCFFFjfwpgz1sjZdjTgu3I53/0rSB0DDHjsmacZX
R635Tcoz2oFOgE4qxLufSL1lkYQ3nKkytjP88zghmQf2mYj6QOzioleVQY0Y8HEB
ZAEnB/jOOi+K1yfJMoekVt0JWQkbCIquaHxKTYNKTzHpJkrHgEIV5GJPCIh9xLiw
onBVtRaiIqM8sVgvwLK3XQXWBJdCPEiu6BS29lDkqQvI0U7+/a/I/pvgfbyhliHn
GBq2cqOL4lWZyheZkO5vm9qjufZR1DbV0Ndx+ob9Cz7bko60aMJ5evV+9GLmbZC0
E5zUlyBybFl3bOU8VLDYKOVWDRMnj8Z+W9IMnOyAWnjDooqB2SomVXzgn9qpMy3C
dsaqJVqVWh2/+5XAEo+Mk05UbVEe96mCCDgQIcnso/qMAnPXzuTBzbt/4UmYP82S
9Oo/EB6IjzvZnrEnbYjoDP8UVH39EOhHct6QT/mpixufyJo87xtWDxKGoVe3duhU
IWKzx3pWgNeFZbyKZ6eot9lxbkBG26Fm57igzufv2kMgiDWoN+hByeJ4gIXY5rIT
B4INp+maFE3nL/ZyxFrqt3D6R4lDdHwwif/QtR+94nnc9+7+6PpvEyjV39wu1Y8/
JsNLZFgymSGKAOASaL2Ys13IcRz5D1UCg/2WZ08GXtJNI4VVIhSfh+lrowodJx1J
AfoVGxjjNeZ5TC4BLcIB5nHZs4xiceHYzhz7N8/eirbZ1pJaqVImkXrw5isVPa3D
hfC7GAf50rGQB441SqlMeTCsMFdzdtMLO7Zr+Q2H2is77NmBsJh5l7ycrXuY5ydP
n/2CDLCzbrRWhFPZlbCffyvm7KNvwEKPPl68DDjhOs3pnYY16yr8f8MYDLZ1Vx8y
YHOZEFGEG2WodUYY95AdPnMdCLyv+cQOfq8u/5aV3wwTw2jCbwTyy6kFfr+pPp6x
V+9Ze7wc1ZRkECHBCNNgGJKsZBsjuZxLX8Zvx1xBMbXTE555xWAEfUK6QKxSZv8j
hUAhuBk4mikuruIqO6Ailb6Sj1JqJn18uWaoih0DSQEDaG5RLwPjGys7yrLPeO9g
o9qKT9inYfsMzBS5ZxiAoIU7Y/QpkOn6GPNEal1IrIRdaE+MGZzawtVmI32Twpth
MMUpi+2C4fwPdZxavVv1DvNCPKL0oHV1slCAHRcJiMY9JVdTlF6M1/6Ow2bhwNah
oCMQ/5UT34rmqbX7NqeWFeMtLEhvDjEgs65TScS48RifRWedk6xhsr/dBaGUN33x
5n74LgNhK7rI12wjPB9TESbLr8lmozreL6wOYcxePPOKO8GJSQ5wnHs7HZTrLGRN
PLHPSsKMlAqOaVK3+omXfv148BGXz+Xi7+km0dQQaHKm6ezit+LeTY0Sp0FFsb1G
Tnz0KOV+be8+6tiHiVJjDItDi/RS8vuAVdC9zUiY+Kmp530OOFyaKlPB9iLvF6YW
KW3rs6FMzKV76fB3Z/50lgRKDOus9yGfhzZyaN6QR8/DVwmhvJp2XIqP3LaAn0cI
SaWrQRBxjs13unqUfamF060SnRFuzfX0cOSBHuf/BZWDSdxfc+6kSEUKmQBtjVIV
nm9TESu9gNqj5gLImQjCTS9k5OGGmEi/pONhCG/0+RUO+WKogWzxf1SQ2gpjxjDb
Eaflg1ypiAj3nu3tbAikxTqisVBD1mCOXpOe3e/s8vVawN2cHCmsdnhHTJwctqFk
lQ152fhhEj255OSvhXk6NnYXRvPOWlnSCLy+AVoVVoHPBD0ECgMf2TFD38/n/wlr
yELyOGoBV+amjYDHs+V6h0kL3wozSjnabwLtSlC02JCHH+OqJXDz0pNkA5BUhHmJ
jzxOIRv26CMBip09pmG0uHWuLghxgYcG2428rGf65bJY2G64Ynkyfr5I8V9h5vEn
Wynsw7Xt/2mbj3G1o8KB10GWxDv48e5hMNyzZbv45vl3ID9512bTLFJQRdmcutnu
Nci/LvG5Pad72HuW16U1FGgvSH4vzDCRnge7s/kmqgIaYb+dlqsJTSQ4aiDzkAXi
eR8COtpmAK0FnTO/ssJRY2TBMr/9BCvIv/acIavEvnt/7RUCMNRLb9OI3N87atFi
IeAqdKoww+21TVG+y2Gw3GvWGE3KhIQCOVauo6uq8MfOU/iHFlnk4xfl4vC1+Kv+
l/Yi3Kpfd+9iRmnWdPKIGI18yCSXLc082Dg0+fhHLBq6XA1oPnQi8f1MPtnqkjGv
0j90o6QlkDuGM6N38xnn26XgU4FRige76BlDXpA6zCF+AJ6OHCT3xzq5TaLcn55k
MN92mXVqH4eCq03entwio5tUiWKTo4kFGarnBuN4XZIa1hIPNSXXE/ejTR7zxfq2
EYlszLgcwIQiV22joF6/bw/O/Inz0HU7w+X3dexgw7j3Zt52RsHRwt5O6NH3IU2A
f1SQjjVD7vZaPEPoQVImzVV412nLMaMkrj/qGqPYuZindLLnVtFlbM8MfHcOVxys
zlfIusQKEMe9XpPeb0YimKfo1cMH7uD/GMTHd+TwDuUXtf3Tx2HVNhF7yK2t5r8Z
FBI2wU24wD5AUIxmAS7n56/Z2ph3L+75Dj3moSVFCWVOgF2vr1M7xl6ZAjTKeIA4
nCgWSiZJ0PCLx8GS9BqaVS3KOTS8S95whsuXhQfKM+PTzTw5Mt4hsDA+N7bct3md
67o89LolymlU39xENi3iaMQDUDrojwhgg7JEokdFRXbbRnq2MAzRFSajWF4HrcN7
TJxD852XHzI5rP3Ckq1RqgM49xSDEXxYNF1vV8ORGAeIcygbrlL//A58tViyD0Aq
52nGL2mIVNDVPu5GcnGeJICTM1CqDCfK3d35eW99QgOmhZ1zDbe4gKCPOwlt0NdO
YKbNAxVv5oNyQ+IZ7Xk6m3doW2A0nG6kOEoP27NvwikYNkd69P6FVlqgKG7C+FQn
/AoyyGy1d8UGB57lv9s2Cms3WlM39BDev4LQqtI+jIqgZ/kAH1d7WlWtWuBdX/6I
vnJwVlEqtNTXpuSxvuvs39+rtKX4jG13G4u5JQbE0ufMJY2gs1PXho44pXnrhStW
i7uk3UrO102o1/CWMEOzrUmftbHtz+fHmv6kmfhjG0O3zEyEwmj7IqH7Sqt6ZNmz
JJZTelR6La5O27pAm+fweQQz3b74EKIwxJoIkcmexdrEqYbK2KDF28tjZQRMcl3s
Wcj4pX0D+L7NqLY3m5k9a7U1Qppn6m18xT7ZmpucYJu76m8DZ+CxfIb+mG0/KVrP
XtrZOiuebqJ9MAbCz3BdpefGkROUHbIarL80nH8r9aAZ6qj5sSiDnQ6YZ2Q+YeTt
y7Zho8yo1o2Qx7VqG+ocIG6x3MwEQ19xjys9UBZwM1GbP8yO06p6+iJNVry2CGti
Ecp5DrZHdyv/hqNoA21LRWPkjzR1bIwfI29RL84+pwZP0U0mtC+AomJpZwO2+4/F
sDRY5/RLNJ0fzp+UjDi05yPHiiF3Z3AoffHERcerRLW/KrKnAGfIPOqJGkXIaWMt
WIHVP41HZTRylQ2K72kAxTK7soFXzAT82OOSo0ZZ42iHIj5eyppcrn3QO6mWqPie
26AHEV+D9j/cr9Aa7WxH8jofKOZHeRDNDTOQdKk5aNIGRGApIrtZUWMNoyq5OZe1
sKs3/4AdPaN7C9vnq2U0YB/OIAv9v947SktC0aWIXLiZhperq9EJ558awzU1wx/M
mQcD3QljqPF+6DFoXMG3HP5Som4Dg+5osRmRY7PP0WwgmocqpeTabY+NF4k3WG8U
eDxX+IrUPWHar/Qx5YTMCxsy1QR6WdMf5trnL846P17BPX5ZCCJj8pi0YdPkPTKC
mG4nDS3cFQOFg4aHI9D8QSI5oPyhpngb9WXh8Huhj9AbwEYnWAxP225Ehu6qlliE
H1WRU1eKZqbz5cxb+MLKO0pFTiGBgL3Yl+VTpz2pglMj9IAGqBGtkQmq290txHx0
2+9aG1mOHsf96QrrQbBaUJeY7Y6e7B2RDTRsE6AbWwj8OWMrWTT47sx9TcU4xzyN
fKZGJkGci7J4+aI35Yq2UXcxqn+wxOeTotC9yL5veaBVc6opLBEKGnjoxl5HIJof
l60gyp0OrrrSFN/RVbL9yfrOdOcIr39JY6JGdQvt9nyIlYDRlb9X7xLNuQ1ZLaoB
ZTONn7r60Y4KwWhJvscFs3xdCO2uRGnhY7fj47E0RyWB9MqnE3muHmCt8Ncj4GGE
EcLgBUlJcZSey/ut9yAhbNpbJgqchltwa1GLI4b3bEjvj5N3u3NorzhSy69McEY0
VR5jl73c1CH5vQveUK7I67uxX7+ZW6c+0cOQ4GJtyA9G8w5DAE4OK0iCe1Ur1CKQ
OYQMk3H8Adbe0QFLifS5QSXmsk/onjc0jpe8h+ecvhGz9sLSjoJjFyOHR6ThNqIR
ORigtkbwWiTBSCD7dCUy1gpc5Tz+3JWEa8anEHt9wdXfuFsih+dL2kNA0hPeGck+
4kWv/fz4WUYgpaGBIsWswU81u9Qsbr6KCIjEjAwA1y3uUunI/xZzpOAqVyw9O7QF
KzDzYfR/8MNLZLyEzOtQUPemGUKa5Ttqz8IsxV6sXLurHDBBUi+p2HoG6x3X3RqY
HU7QTnWA1OXbQuB/RNV+0vT3Q2B5TYu/8e957e68ElY4ICtoAsIxZ36DKAGSBO7A
2n5K0t4jvtFvO8u3IF/4LM9E1FCXIJbQc/MNn0rLe6fkIjzYRhl08QbJ91Pzn5Kp
7x8ID5YeBrZaNjGQDNszLVpHPhnojIvyeak/s1oSavH7/PygUN787kNSXfKav84V
vKgsj0u2EWnWQoYDtlx57D9S5WP6yJnzjHDk2hICdIWZ7WaMyH4K8vKo8neaTWGj
jk894AoWTDJmd0hUZ/uSDzKx0Lt4U/9I0ppHkz7shy1xYFRUA34L6R7JeWFM0Ooa
9UdyLKuWPhJL5nN1wnem6AUndLGyKs5BH/eUF3YOigFyy4V0Sa3stqdUbtfqP1tP
nVOBnewRs0AGRPRwpiZSNN8/sWA0vtRujVy7/PNlzftAqCDgavsar/Pf5pN+2kXl
wtwzYv3MJCuKdtA1DgGB2MRtd4RnmX6jQeshqbIgwnbdNd4Kcf5WO9MRg2MlX9oJ
9SRXSYLLFoMcgcN/1PYcfk9USkZvIrPuG28uhesQ92pOLv0AnxjiG2GS1xqnCp6A
dq307xBOaCC4nxZkgUKtnZ34ZdvqATcSe/mk0jOunAdWcc4kmDOuJcbAfuYSQhFw
iYoqKyvkq9FI4FVDl2J1TcBTWCRpWcK0/R/WBEIFenghajoolZP9Z0eKQpTt/PfF
S2dGWDBpzHdxbh7ZoBx0LeBBl3o8McEK9oM/vYZcixOguPaNVcRKtiu6oc+irYCT
XY/GOWLK56rQNXwWRS/yIKBpZ3PhD9g3KKdcmzVc6JdIBtRvCspUa+lA2HdHG0Lc
hyHpbf7+PN/BDf9r2wtgvft2CY/jxW9jns0zTvDW9W1s8t3MWdi3L50LqREC/gO/
9s0gX5vluawON+DU9uyRn9HyGo+IfDA2ul6Bbc72S50oJWWB5aRmvG4ElQGU1Fix
R5f+BRkvZhi9CFI9cGkVtuHSFqTzA3x+ezxqG+gUg5cZ3A4LbQjONtIalCpTm/Zn
h+oNBy3SrzhFBq9hA9YoAF0pyroofkkbgf4Cm6u+zFm7I8vttMcsDOKfD/Nwq+cs
rlYCfz3Bk+6ikdGlYap9PuQGwjf7nWpP+cP5f6JWsChYYx/bV3yB+oWpyK/Nn7tc
DFvv2LyCBmisIDC2bIfP9qqnlVroOiVSCRYj8vfOv12bdcD/l0tCXKdduFBBfmf5
UsCzv2sHHvK5dz73ILaQsiYoQ8EfnaI+UYSPkxmEoaMZvw4oKA1AjgowDADKrRo8
SJjQFPLBd3RN+VgKUi+DElZ4IpmWpW7QYRnAidOzwovuRhjiX6QpWwZhx/OEiVxG
BKRiZ0qg5WUMRXz1QvyeONJ+tHDsrC7nGcuMBtREiUwyl4VCyblgQbrLp5bCK27d
+5+QNaZjRDcA4Z9UBZLUqXsaEGJb2hZsbefIpqcQWPLiKcmWhLOHmrDBVbzhAV7s
1U4rbaNtFB0GFlAxR2FGmUARbBijZbwPKaXq9PYDtWC+vBcpvez6eBv6XEJ3xAvj
5EFOxsWuL+jJzT5paoHMyUTnbUh4+s/eV8l+7NHXXRSelspPECp7Lp+U1JMGlfSQ
AVrMoLAu0oNdcJ9XdRinzwUa9KYLPwQkgOTfZijROp0pRUTo4yZGsjmFEGYHiduD
DVb+hcnnAJFAccnRx4GLJH+vSCdTb0Bi2IcNoVtH9/pCSHMZVSMMQA6KUtE9rg2N
jq0XwzFeAy0wUsHiB4apPAtmg5RnI5XUo1yBupDyIEmtebSgWKzuF3DJf08pTc9h
q/XtbZ8bi83Yj8mKGvafQ80n9oTjWJs1aOA/6+Wnu5nfO0n5LBIttbkhwymKQJdL
+w6oFS0iEO6Pu8kuQpir378pzA0Th1miyGizd2JoRNQPcz5QAyslV+UW6h2oC9Os
KXYg0l1/GdIH1M7Yp+yGwxP3IFYJhbJGxwF191HEmVMGmR8O6f8SfXu9f0Xl3tCK
hHRzMpaC35DrPqG25N8ZcyE8jfRwXxBspnNX2OqXiBmJYj0PAHKxyQWTw9u4U17B
P/URFxtp5wjOoFtjdLPUQgNBYZ5z1AkZTa9DBzcQcbzVtoRufNEpQm6iI53d3m8L
Yu3ILVf6PFDKtvo5XQ3P8ITOpqawi9tDZQfHFp/Wk2xGJH/dr9HghwLEx+o7ZW9X
sZsBl8vh4zJRczQz6E2/TwyPKoVxfRjznqtazDF2WgQl27HeXdonH0DWxPAaaHWQ
ENUte4QSHSzv4TiMwdYqYJoRUz/E2nM9eO55vHUAI0L5R6McN3d86dChVJnYEiR2
xJzN2GvLqgFobVq4++mu67I5yvMR8TqHgts1vfUAA0r8Ssa3BfHyvj4ciMmoIs+I
oYFtAY7hEXVXQ0Skg2jQ+WKNqdBbIlOTqK2zzRO06DcxeNsE+z90Q5xsyFoxrgwU
a9AHC/wjviTlEPsaEAF3b0YgEkPUKwJ8+kfFfED3FpR4oi6TUMkPfu9yMpWoS11c
IzF/JKl8NfYZG2QpWzbcNQwOPrkNtIlg1Jsff3gypUKRdVifnaL/DsHUYRrqJRiT
6hp0D8CUasxK61QlnrCCQUrSIAhRhDxUcE7hclqVamKaQWyiE+TCaUCZmvH5RNwW
HTOyLEpSTFEPiOwmUUNk++0LTRZcX0zgQUjYDnLoflM53srl3VStDWU0ld8kvZzM
Oj3z7NszhEI38xTbPBjJJmpB5UVaAUQMNXzFkGLKoyEbT7bvIAorBItb1nAabrdc
amGOUHlWc22U2Kajmm702PyxuWWmbhlTvackyfaP7pBI3n43/Up+CXp7p1u43YBv
bihfY6pD/nfAJ1ag+Z+tVsk81yr4hOxPa1N0w8Ogk5rstH5klhHJ1vgsKR2XQ2Fm
X1lBS5i48iPJ67A9rpRj1Ys1YRq5xYIyWHk9j5zznVZmojAh5ea4BeuiUrBAqFRM
2oNaTr7kZvS9XskGyRhzjEqns4v69c9VvBafqlCjr8f85qJWn8NHTTE/glWmINet
m5MtrjMIFze+D0w1ZOq2z892xsWEnFYeuGqMqfzdAcbW27kZ/IiDdyD1UBAqcwAT
52u8k/0cwtEdwZjyU/ljDpYrT/XBLOg9bKXFcnhfb9NnnVJo1BAZQybSNIy+TiX6
om0Z7AgU2s4v4apYiYKf5r4mY2E+hhcMh1Hsgint6mt18Ik2acXC2n8D/JzHg0vU
5PGzDdand2IB5snlC2RC0PjQdS1es8oPN901nyf2jKqaf4UNeTShs2ly6WHXsuHw
1Aqbf/T+3qzyjZBfy6vPOwys+/MfqHPafjzWR8QzgUdEhpLFThbXeKse0UwnA05T
npnfFXd9SsRzZFxtqUkt5ZZD0QpkCipz5GIJ7QZnl8zsA3D0ONvieMXZy0OfUAVM
kQt+Tpg6oYqXo1BMtCu6xjHSYP3ECMnqW/vQMFld+LqXOWMQKmPua2RJN7gS4W6W
K27QHztdU0Nbh8aaiBjKZrvsC0F2jNL6JedxDfCW4ui1NkXXbGX3eedZpQ9cRcEe
U8jJiohSzqHYbFQ9GS66CpnSb9kW2fDm2pi3rn0+dx3FhSHVDhc78ZfFvfklJy2x
e7xGRvW6VhhGdsDhNOUdC8Vg/DJEWz269gON++Zmh9dLFsGg8v5JIiozXPkYeMu3
nGdXT+/9H/9/fu3vS83SaspCBvjLFVW0ou3pqtQNA2Qd9efePuNUjRzgfg7Ku+Vu
6fQOeeZdR5dW/WtNfKLUh9mNLfp881HzzADlt4NVuC5hAf+QWfwkJFmXQopI9jBD
IrZydZpGJYbXo3ZKUuyXb+1yQSGu2sNxDhtM/cp6IprH7LaUgdC7AlIdPEf7gtXI
wBbmZS557Kbx0kvK0wdGkD1JWMH7mFClZe9tAux5p6bRQRbPkcW8LbPZXP+82tOb
2h4cj2SibtoiahCvIiDPBmTiBIR96RGGTLTbivwrMD7JHPyxbJSEIfUfOgenUCxc
ozBst9cWNvpEH7N30XydY/yjxB5AZpVEAQPxpMQL9qH2I6Pz/HcN86ZNh9fHVscJ
1WINC7rvTTY+OXYn6sKvMfyBBaiQCJYwqMLR3qeYNnyEDqRC4bxpgRQUcKZE4zL7
zI/3dYyAM2Ey2kwBX7eonfGj+3xltbZnJA0FRaj4Q6jY7hsIF1/QbXN3KtB0NWmg
swfYZtM4nu8mkwbP0V/t7tz8KWJJYXtScwvLyhGv3OsxyzmtVtCTYWxV4D9s1ilq
hvg2c0rRuVqG64DMlfRSwIYiJtpx9mBc9wE3lOot2Ca1eMdq3t5SWQqrN+M8skrB
iA/am7lxokRoLR79TFbLgTksKmKNSTZ+L2EgZOlKewpvFtKT7JUkzfdevDxPL4ER
lNn7k00QMn1hDuqPoogr1PrfK3u83c/13wplt91wyq6nkX0/Is1blLvmDLgD+Rih
oDZjO4NiQPvvGObMFddcUAlCJTjrPFHsleJgqpJOdIGgBSkhxACTfDkzAGuPAFQL
ZR2O0gLvCWSONYt6A+8YAhdIQ4qUL8KHSRVH7I43mv7UiEhU5aktPFvqWJ4QcBUS
aBf69STWiHtNko4aOhi2rTsUZ025h33p3gyp6VtL1jXOxA50+K4aUC4/prkqbr41
Pbfq+z82xI4d2yTdvbV8kEmRJUXkrNAectW0/Rcn2TOtRruiAgjj+oIjJRsZiO6p
LW8l9cU0UhMOGH5c2H8npQFn4boXnD6jUPfFyShOuDuYeYstCc4O9tXAwdKXQ5+8
D67AYgQGeqa2Gej43jGsCll/kVKhMspBQsbLYyUKofrXZvr0ZuiRw/ThElbNDX8I
oBSFDoK7p3FuSNnu06ubGmoYkCMCalnMl1NgwCGRKubThF9s3fgpA7ySKMdv0+kz
fNInS6KGD49sI+cTxq0sb8afS/WPf3cenh7wHrGzJA9+Uf/olhW7P/7e964DXLk2
Bn7p3avP3vatGd+SCL/g36ZRI6d27Qnkbo43dtQg93ayeltIUU0LaX8RLELWilQR
HRBujsGX0ADlT3E00OjAxHEPY6gLW1+z4bObn3JYnSYy/QfKHjCD7XiUZ/VErv8Q
Mn+24eQqxOg6fXLxo2g9nDC29PO94f09k7XFqXT9fDVRg52Sm/oxfAbCT1bVjV5t
IaWR7QcwA59Ufcl2aJCzOg4HJBDFfVBglnIw+qxqgeHZznOzKii8/N2mwwujhPZ4
DXZ1v3NQwcM1X9bY/Ehv0WYiHJSH/2M5H0XQlTPjpRy9e8h9Ibtlg8n/kardKixF
LyedIenRbPAp7ANNDST3dPS8KVi1FtDIPPneZ4tM+GzMk5YGZyWYpXGv5JgqkU6N
+T+ra3VM4aEcX9iPaLVScX4ITjLhXNGjTRmhfvVgL7ZBK/DUhf6uLz8KWa63jVJU
V9BqTco1p38FNvAl+vEOhMVgfiFaDn7JKej+98BIucbxSSVjspG/JgC9qlwRbgZz
hLxuUuRdOXUeDUPFT4XGjb0kLGMs5XRHl1N1SKKmqcEFWBvmk4xrDLpu7rE95FM3
f/tj4eVUCIkCZoKiou4gh8TOdxzK7HrSv928DSTUJAF/7SSpQgLv415SE5bC1/zC
z9dXBsxSX9nexHaC8N7ClbFwpn2keH9uBNlsch9+XEf9RXYg4YNFlCMiJWEMTyLC
bT6aVLy6mi2+1Mln/+pnOAopmHdhfphIdFULLhE7unnGurUb5Rj2mNgq5VtujXQd
Jod+nuIx7+fyCVM3DUvnmiLhUSmiF7nIJ3Q1lph/qPACYqBQbunva0ZQypwGnQTp
b66iyjPF03cdUGeitWfI9/wjADQ6ikywgQPx4/SrST0ODzIqxawDK4MtCUuJw/YA
aG6yLQwi9koyrILO0vyIo5mTYU67f1JS94WtLhMz/yQGylCGohegFRdmHqYxw8Un
AAHXzRy/bRkiwJ1NMLsnBs9HlcgLpPItK9gjEraNggvqLjCWmmEYNJ7eoSwavNJd
BuFsF+nAusj3nUUBh4KIJe9U0AvZiB/vuWIF52WUgw5jTma8BBm2WgYhei8/SPxO
sZjT5jyh5S80E9eFKBGK3FX3LwyiUNy1Whlya7Tm/UXHzbCTrTBfEhKI/Jjnz3wE
3xCKYy6NFrnWQvXLfjSx0WVaXlXSi60hb2qizA6QCP6KZdk0rQT1uE1PQuhU4Cdg
UH5dQrZVMUWapdPVuh7lF8eE9rV3j0mMAFba0qfSQHSaR3+CPDc5QNDqEMi1elav
G/OjIsfFAPlfd19ZhM1vQeEUXXOYmuneDboFzevAw953vwziBGllmUSfD2Wsimbl
94nedHzj1JK1lc25xDZI9KheI13WVbStZJPE9wfkWQeDZyaQWGHBGBkqkyLSLbyz
nRh7BawYLGRlS0ifhNJZuhNznfKOtMc/LWE2u8XK3odm3epQSu46/g1W45rdyAE2
GeJ0x0cBQCaJK0CEFvspc0wD7WkfsBiPuqMzOuM9traNAzVfwSX9eG8qsw+hFyd0
quXlOL7Y/vLoQMolm2wUbede2DRtUkZGUHAU1pRot0uW9IFcaVbDEyQO1TAwnxp7
F5bwz/a/2HR9e98HGWUcI2X+Nciqpk4jZy0sPPi4wxauedsZUm8ebcaas+53X78r
VKweRMbuCZLj5zzuqLy3au3II9NbmtmnpqoL8vdoB1s2xIVRY9EjAVfLEFBpX+/t
/BK3u7UzqpfCVqUq2KV5C2Sp4Oo9JQ0Wqg+FvgFQ9/2oYBY4gUHUkVMwUGyxSzTT
ql+scCc2AjBKutZ+ZxmZ+HkvW5eFOlMiAK12CP+eoT2UXJUVJJQCEhAyYYfQpDVL
GxweQ2w+nuW8WEfmOrF6XFp5TqUr+e9QNvq4tXMeZeIj5zCGYZz5+CHB93R2dCha
ri/fonft7Y0RtyCgoO/7rKrvlwmblZc4izsf6KZnVJZu6sFaQCm8FHpuUPqbr4bi
1QYiGnaiB/ax6x5LwJART3FGGicJ+4Cx4P3AcKjYxEKMXLLFXqfm/x/9UT0SX2HW
Ytnm4CRbfWoh/x96+fZxkLtXwOyI7qKLteJ6GdR+ft1I/YZYVCxOnqMFHJMLSkuY
/Hjn2qq2vIt47WkXy+EEQGxJjiaYD+Mx083scPwGyeaCFX/1ykq8HmWunEZNPx0F
AVn7M+g0i3bhsZCfHD1/GeHr9kMd8Kc0YeMW8khSs4f0Dn0/SnJ1PEtlCYJWVmdI
8sAkpcawoVipN2HGDXlzA6uzIl5kPwKWlCcG2srshlYm7FQkUknP5E2KG6XNieUu
iuv2tg6ZfM8+mXp/XTISJUrBU8ZwUZj/qHUfNQ/C0CMqJrh/wDFAYdzoe6nzraJI
w9Pw7htBmk/nWO3isRYhJudRLzkcJV7YXLkAr1QDBhj4aa2HOwTTz1N3/JZsMde9
P/nACwCCAM1wMd6lV1yWPomDJ7AsOsjwUADTFPXeuLTzHcpvDY/ZLFXCTsLLpnv3
HFNJBUnS6SOqInrKmEP5usk/bfQGSwI2RNkMwHDJLXipFsGIAUdVX69HSZS2gCrv
4PrFPM13XpgLAaKAhZ+SxMKqSZDVrnLUqeD+clyFj14s77KPQK4Jf0T4ji3Qj7T0
KZMYw6KIRTbIoGXfXWxl7MwAPEG20RmpkVQ94kb1esptOnadeeom5RakISkQRHw4
mDfiIY6DHgQD5A+MkjgD8IfTcyBaOD9Hto6Nfc9JNzq/wmntGgJft2P7a4urL26s
ezd3V3oFWOh27TUBrCi280qPbJS/BJK/5WRHZMHxVhAssh7ECboSaF+wwJsXSInR
OqLpDIb2rOtL3L2ydh8ioif3qBghsDgc5Jmk18U40dzx7N/rvkCr7V1XXkvVy6hh
EnzmNkwGiIFxV9YskoeGfEKG35ucf1CrTo2Vfi4jIHrbsmEB7hOXVJZ2houmI/7L
m307lhfaZS4ov5T14mDRoiaOgXyo6Mx3vf0uaBFYwI5h2/KojMXUG3PVMBuUXJjc
AULXyHfbwV5Be/mTrTuvsAEhPBu6ElXjgpNFgcCQ/NxZxJaiefd0BV7T4LBUH7dZ
L2w9XSYr2OhZais6WYbAFus7xNCHCLwNqe5dba8A5enb5G7KJUW1Ois8fovPnWS/
6Q3MnY6JYUWVNe1ca1Hgc3+ZrX1pnKbuQVw3swgKBB3wOOEiMijtP3B9MH44R4U1
snqjHaoDZgRuBXwqiGa9borrT/uRLhqh3zI7PqzjUXfZXPIZdx43QC0ZcvsotvaW
O0FMbOxH2rKKpB9LlDO9gBPLK5rs6W1ztSvlVvD5pvFVEC2JIZkNneK2WqXVRHuL
wgYdnAoupvsysZgGnQlqjYUKN+01veUf/+T30IkXFdJ9VvZMKZxXHYFCOsVI3gsX
iMEblxi5dD5Y/T47hcTWKkMucZfTNcEKuZjmrojm3SVnWjwItRF5pFl0dOAI/kyK
7wJhl6HM/eNPWgZARbTXPccDF3fablNAo/cF6BmKTLGi1QCcWI33HPTMerAHXPEc
bBFGagum+ZAjkqn2d8teOAhT4j6ywUHnomjE/BPrFLkyEjTrpU+EIYsH6UCfchch
1f5GWU2HbJ2Zb4NemlsFJI2RLA2//B3h20wP3xyAqojq4zRGMI6DF3x2bfxZIl5O
4DFHEI9yxrrjpbQWOS7F0CpuRoR9xB4dz6/0aLxeUO6okv5SHQE9ON/Py1nl9K4o
j/SAtCJMsrqG1/HA5EFM3UzikJFI1Bn25+Ts7QbNTmw2c4uAptFQZnZPvwu8n6W8
kBb3aCmkuQKYZdEjKdTTS48dsMK2RiDlPVgD1FU9JOyznuszjy/YTRrogpwDWIqJ
11mibr9pOHEJnHhNQ6AnZ8taBtIv466qaF2fDR5p40ODYB8+CHn2YvgMKvv4hLRV
X/r5WxIIWLD/hV5fgBbjp0WnR28R0jiJRfGWBBH0fBocwyTjKrmOsiiLGYJzbIC0
GriM89F2vQvJlXtEoABfYLAfQxoly2SRlYSTgF9PARbLPGaiZT2U/jYNRSXEjOeu
0delgQsLAN4Q3cINe2+20TRYnPTwv6jdmp9kpS+aD8loG4poDaLEW6yuc27oR7nu
kb2II0bHMtwL7Y/BVyrTO23UKQBAQjO5AfbAuOb7PxLbLUf8phXiy0Hckhl8znXR
aht5Hq3kdBpyka4mm6sHz0QuFw+gUXnY+FHw48JkKth6hKMWJaljNuoUc2EM83+g
puuvhDBMjPIWI1dWHjGzFhGurUn9CxMJ8mYoAqW0GiISxT3RiJMVt5CsHjrCB6b9
ImzBNM5Q178QZ7wy/Cc+mKsB7lILn88JYzh1sY0ygsx/DcRH2jOdO8eM5Lxy6kBj
G2Ku5O3j+cgI0dDEgWzDUi13TVzkVanXp0G1JRT2lfjfysVXPoPJ+6b2QGHA9Dmm
tVNL81jj4Jua03JhIN869Q7TYhquT+dc/8HV7vMAPRl39MUojSYyI5k1xhrExyNg
CGUcYXO41UpL940Ry9F0pjwFSHZAB34JhPVBv/g+IckwJyjtZYbkQ3mnZRenlNYZ
NBO6fcO88DE8auFMmVCkndliQHbcWX7Pe1221m47Dqyzg3ZTKMGfeHKPSPp+IqBT
5mC/YO8nD092bnQbhIbKQySafnJq1L9RjMpvQ2q1t2PE8zSiucfRL5+RP75WI4sL
t0OpStULoC4ibQFLLPJeOSieKM2iJwZ7Tu3IoabCNNczvPTFmii9g+bFWPUqr0UB
EDmwpI4w0yNWME+1ZPvTfK25aCBxRzEV/A2xtbjCHmGizaU04JlvbaYJ9eXYtTMl
TTkySueaqMSJjtZ70/326fZNF2hNuvh27FNTKF9GFgI/x6eox2O9iYQ+xo1OnP6h
feIfxITG3hwXsRdZkgdnGRh9gdPAWfH0AXCBg3bmzf0OOOnNy2ei/8YLPrTIQABD
IAYikXmqX5J+NHXJDVC4akwVqlDarUM7Og8e/thJDTMnFuAOqSF+eWxC/wGbzA0H
4Jy1WCcAldchUvlF5rHc3X2iyomp8e3DM23HmYFLchBa+QBPfOsjN1Ah61gizYWI
1n640pH3cgmqicko05j1Ot8xxPl3PFCfzm4L3CkUrFt8oROXxAajfR5+bdWBsEjs
axZJFF+HzM6pmH76QMbyiSH1FnnpBgpoMYnYxTkzp4Z0n4qsJElk9tYq8FHQtbbB
Ks3j+fVS7t10OA1drTJ1c0VWA+E0pulpwUXz1KAp2NdI7gfEjrioK7SHsCxb9d58
OckEnDPrHCjkkmVKQDTFLqMF+9vOXPJfykNyTPyZJzh44QonxuZl7IjxaG1SLW1c
6h76OhtIjbeWfnU6VwgL5rkW3k3U2Rh/Iek5rSL8l8lEVV/uXKyqTtSDEb/dresj
dut+5x9yKjb1hEqsfojC2Uz0CS9hYcYXOubbQylnTOUKKgqcJgXvqwiqGCP6Jdum
uKjNUGDB9Ny6j1cfj/91fe/gry5Okxreo8vhTZpgEzEe2IaiC6kt8YDT6ObuC8MC
/cNj5WP8zCyrmGoA39D+fIpUWEtqjY+DR1uRPhbCrOdsvcQJwaZv49hbRDmQabfX
U7BbSMHDSuSXXAgWAcWtcYDWFQaaGIBF2QbqsdDHxggPf+4N3XxTuSpNjdFl+Z4c
dG3y6n9b2daHdtgIXT+gCG93rur65iyqXuEe8bI0MLOFahn74yqq2EWWbTbOG9Ng
opBDSQ4UJ/B9OjBq4x/pYhLypI5XiIpMwff2RTznQQvEKxjcJqkjSElsX25NjZex
AVegs2yw4fABWGDE2T0kQV08zAWgM8boX4v8ORGl7QatYR5sljOsqVaJf5RGiKC/
sHvXq4O9HwEsvFLw+goDNKG4GM3fh+KyJaeZxqB0Zf0tG6+glwGeg0A+X8HyZWHu
tVQ+yb686oJ3OFtgOxbQD/8McJtYs8dKDIGYFiuSYB3zz7zjz0Z5xjbCf/bcwLlN
Vh05qBkegLG2KhfntPl+xH1lxP8R4ax30MiK0LqGQgoYQCM25XDR1woGzHQ2MoYt
bJoyAax7WWETx/0PmcFW2RKZRfrCfiymURkrbfFgxv/MWYRrdixvv0JPGlIOIdcH
0fighZSBZ9iIRoy3ABX/F00CDO72Ob/iiAYPRlCwQzgfZ9xgDxu34yKY9Kulipzn
eWPpPOSeVRZWTyYNvZRJ0SlrqYqVyDR6kLYWQTdvIXGZkorTdRaJqFzDhgAE5CBV
qphUcuxUg6NBMJQOpVSVp9C9mU4Jials0W4/DOmNVew7zD8T9BtEctcmJApSbDhL
t7zQmQcEM8Yksi+/f/COD6LA7nEfNDgRkPi32o0BX/EsgvWXJRPe/MRmaJt8Bqbq
vpcnFOM6dJphnMd339ygKF0ubEquYPRQdy27wuzjm2TTF4ZmFYUcb7iWkDcC0fE9
RvNJH48JWOPaqJeqBsKHira54Lsbx4bhQP3R43trhYQawUk0K9WbSqpHd9raA1J8
LzhN9GnBKG5pst/jvxUGrKLg6iipcLOCgeUxkUd1hrB2bkfFS/aJOFEdVmmNMn3S
V7mA/NqNFwMV5UVSr32Siuk8/veOGduOVt48w/TB18kaNA14o/8lG3WEwVBhwK8u
vuc8bs6xX9nWp0/A4PGVDHnkJWMOQ/QzNXaN+1m+bCr7mEIPfSYP5YP5Aq8AaQ2z
PM+DPkYd/sDZjkFDV1NXBe10TFibo5+kMGG63ZdalgIPxlr14b0SRrkaY05zYGeX
mT9YLLxE0g1RJ4ojFCjIRhqPNsUnm5yak/G5Ik+k4OptabhaGykcWD5WXYeC6UqI
+XB+wikRE5/qODrUkZ37Q9W3gkqkCNtUGVE4Ktghy+HRWksv59l+eEXf6iJDXXJ5
fNhUyAThtAqooyqiuqEXfIebkPof7NipE/wj3MDbYey0SXQ6socyF4P1Q6Vn9Gq1
gSF82kJZJFAOupe3C/aY8cm3S//wCAqBKSq+QBPqzoH19sam8Z49vAwwTT12s+/O
iEt9ZcslIMEtO1+ZIBmm22Ys/gTHxFKWDbKO8jPr9fWog/QpcNnUypevdeXcdETB
U59VVJ5epdQQiQsQAv7BfwjyzpZ3ogA3nyP+d7A4l4Nyfhk+ygHkciCHU3VKjmNI
CilCNMUJhX/rKejYp3pAkrkqiTlDkmGIxDD5wJ+E86jpiSMU2fN2t/6pp9RjH37v
+RoEZ2QnzMnwRxkAUf6UwMYHhFqzc66LHWsoGr7rZOm1O+ArKhsYkXXN8RbSOW5+
3TF6FOR4YHVJgGgxymUE8xb+39edF93mzOl8xO7h7pXnvI31RXbbRhy3JpvVw4T3
I2mWIXP7C/2OvCvupjiJtjfCVu2e9q6Nr9ovtatyK9+voXpuqCHSUbgHXSoAobLB
Z9qcLuhHWL/Ub+fzoALLWlLBkcUce9BM5EfB3rFLxmXELkY4ahxuTXaa3wtK1EaB
/8696YHYhvaRg1pVndQlRWoMs/2+3PsO0no1eEyDXYt/K31FjMjbnvEmE3IyRPri
UieG6CoSFrY97U7M1vxhbmhESvf/BIsXoYoYtRxHGfBCJ4szE8t3h5GqeoYt6U/P
4FJQTj1QVafmPtE82eN9QnLs5D6CA5znth+YKiutVBced2MlJWmXBo3YgU56CKF1
HMZS9qIxa2CWmzYx8TjsZXcLyypd45FVxBRAJYtei/qR4hRRt9mX/e4YEKz+gyBi
cDDi9obn1wyq0YEKPd2nsQpVzpNFFeyaPDV+fafZPrR6lDyn2N9tsEVMjAgIgo3Z
FiEKXDls8cw1LPrWumUYmiTUbaIbTKR4lmFYhbHf0ImpM58/23/IDF/FzNH9eubX
y4Zglh3G6pmQ1EqCxHetXuXn6uZhaJlDKoWLFZ3yE3hFyiltyN6LWHvJSJdW0fOv
X2cAUU0wop90sIu25KzcvPYhM43ttGBvTjxFLk0sQvtk/RiRZShiKy0nSXF4J2P1
uUNhqxEqSlSdj4P/g3Igbrp4RlxpJPEUJ7kDjO7J4qJ5aS0Qm7D54/m/Hj1ZWEAg
TJbZbC+NtqA7fuzL8YqiI737bI0EL65KuQtTMoHyRe5KVHVChH2ceO4xKq6LdjYw
f5GGE8pZxxNr52QPL9IPJsjmjhP0bB/IQ8TpeMLZRmH3tebXcdvy3Xc0s++kpO+H
QLTUvElBIzD/KOp9FwUmBTr04HDetpuFIw3tigrEXCoEipFv92pQbuEKxVC7E6yR
mQBtrAbXz4OSZbrlR1U3YZGvTAbWeokthdJSolTqKUgbHDHgvlm/kgLouzCccigb
/EvjilQ1lhPQ2dp7wTKNohuTURQuDqpiG9/btRULjDVwcjG5XAaveQuvYAtDo5c3
eehRkVbkwhWYLfNWC+h4UTDQY2JgX+4px8/msIUhHO/c3Cmp7R6qb1uQQf/wqriX
EqEQnnIJotfMARnb5Pvumxqx4dq8K5AFhwjfV5iKfnKKa76xPC5qNd1yq0Cmvs/M
L3ue1y+uvIOxltcte+C4dGtLb/Fu3EN/aZDMj8ei0fOILaeA0vJ00h+T77Uw6Blg
LY8lsLjTjPUDP6RNoPQiSeCsH2uYGPGdGfmPqzLnx+tiLoRTfn05mp0hk50NUtpC
XRX76vLvmCQtFDUe6frKw8E+u53ZPZ4ZRfXCdEO6BA3PHoqlVVVn4BCE7J9U3uvG
Ms+vtHhO6pJ8KP/suMQqadBliF9WMG8t40QoX0izR+WTaQ3v8RLpcY0UzOGpyj53
5HZxitJOn8XpHhLRw+x61NcXLHrBwnS4as2lsncVhVqSar6OKZ9CS1NYjF+/vOJl
VAMplVXwwJkguSXk1acPPHqyhQCveeO1cENRC4+y3lBwtm30sb+2qjkgb/kbBYgP
MUG5JDen4mTcaA8k74M+xeOroN4GrL3P6l6pH5N4Y7fbDPXdZy73QLHIXFOCFbdC
lSb450iOE/JG8fyU5tsR8M6NuT1UemxiIZ1Mtrdr3QzZLCxkEVzd4lnQA9OtF6AM
c2iXhSxCNe7F4j7rouZSyaEXp7mf+Odjb44PbDTUEfE6pFKbIVSxAtu6Z73doEkA
ZN1tW42Nmm6vRZvOYoUiUkFbubfhfLzFVhUSZ9OnGKBbVo/hsSsU2NbYq2QAaFuN
wOwaZv1uyXt+/YioiKpLxn9nWxKX+AynGB/rTL6Xh3NAWmrAuWnJ0s61Ji/6lvXX
+acZqdKausexA4ZT28bERTLNyQKvrPSKwrajqdrChn7T7hPF0JXPsTtm955DSWRm
nKqYy3gKxReoH86h0TzuYZOlo2wowvvPZ3EWvlRQFE9ULVR4c24dub3K7hau1gVZ
D5+Ar/ds0mimhymallWWNgBdJ62ZKBFq7R5ITk7byr9yLLcjQX1LNWyEmEBgjuUr
cm8ih8oNvMrQWfD9wqAp8DVgfqCMuA4uFKZyw5kCt510K7I9yEWYrM3sZ4KD8ruK
V6kuhZnQh16bmmT7ZYAJGXI00xAk06eXG9cZJXlhxQFUXJmG5l1DDFGRldNcEWkX
TtT40WMZxS47kwEMycX1IcfU7/Op7S2zKuFBGDJZpgSyT6Fvcygqe0GFT4eDLbTK
vUvYsVPZet6xPo8cHxSZJS8FaM00gbu2r+MkExt3SMzVCOJgV5cO/U3RpdNp3GOv
TDblvzmj+zXq3zJmNOqukVkLDgQz3HOBsfDPiEOSdE9iNtz3WI3Ee5TTBQt4Ou7g
aLleAQw1mx49R2s7Os/xZHdOUwCsjLYLK4SuoH6Endvnu/oG1z75mg6b47nHlMkX
wCGBCMciE91/wXQDja0Eu8OuoKbWPWj2/mfOee14ZL0YI9XiFRYfKHlEU5xz4iBQ
3sCKTJg7xVHM5Z8zWn8gdnB5elCS8qK3+LT6Huy44uEm5q52DlSXWot7l3f5yJMi
Ec+8EwrqVO+XFhI2RYA/X4x6FffjJk+AvBB6D5UOtvf5IaLji7bG4nOz+KuGGt56
yD0dQSddMHuQPuW8ewl4/JVMLW9GWgE644wsvTbhDpkIX/Lwn7boVOwRYwtdbZNu
kakBwYosXm/+X/X/oHegaVTTZo4Dlhab8m06dpMSdT1xKR6qm/2HWrRSvipN/WID
JjomxTPQhothg4Fym4MII+vE6bwSunq0sAzJ1gySybfop+Q+iUSGkvBFwthW7VTe
3+w4Ni1Vy+E5511khe8YtBi23PQ9vZtWzVicAJR6TGv7zSswN354reFw28wK99pJ
14mzEXmc50LZ568LdlBzF00u9/OBIgcOVbSLX/1EFHOJ/+uQBpyoNhZrvXHE+AmC
rfps3e4pdQ1jyaA5T6cX/gPoixtaA01bUe+KPvSwQwKwdvfQkEvCWEGDyIkswsPj
S1Pth5FE/HwqHz/oUS6tlYpQAzudaUsi9M257kANSTFYRkh82Qwb6TUoB2pM2RiD
rchoT5gDuoovuJT8zWEEiQdqLfw0r761yoz5L4v7VtokgWWPFUZIYgEsEtM/DR0Z
4A1iFc2DFj3ix2tV9ThsHWe3KBysYTALtY/mXWgQBp6ojC5fgCzCXhg+hbRJIIOw
5mUbcDs8iXjIvjzo2fSJumtJorIBXE3k7oHhxMF26iXBOFDSHZGKfK61HA5QXLVH
b/jgB70xoq6TNzeUjzA2EupET9XStZzhYnBn0kNBxUn45qshfnRnQcnXRpQ/Ci5g
68PusYLRdJbdwilVmhmce+e+bpG1JX3qHMbRmzosgq66vfRxc/78adP0ubmGBCzf
mdeAR2y/H6+f0eNSqvJGphAys/2TK+fhSxEVuV9dBRhYM0FseOe/ml7dECUWy13Z
7h1vOojq71pEOppk0KDgKPhyc6otBbOgW9UFGQM8Zm9LB1Zz0Gn/48vJ8YqVe9wq
bqA1Amk0WhtFd0D6m7asbnOqp+tQ6JP7DrQMjdfMyIgUHeFymEGbU+adzkoqhpzs
irASDfolnkeMeCPdVcFsYVW1xpTl4UA1YP1vZMRhSSOPiVvosmtkmSDJ2s+jLrJU
nXuUimAHfPlA9qRVvCmbindT1oj83mXG1PXLf4vHj98G1FicvvBowXW/uvZLZHnm
Q2mPBtNd1FTJvNlJ2mvu8BdFjYaDy33idS2TGGiUFG0RriSHTpUK77yyUrjx1LNW
lstFPZaiBCaYr3B6TzTXvnQjY1jONzbCv6ytKzm12lP4yg/rgfbu836XwshymqyT
zdoR0mDZe05GkvmInJT6uYNS/9OlmBipP/IDyRNyvUWi7E6+FpNiDm6BoOk3brrk
R7ACp/aUP0xFC75Ym/bFERzaid51dMpwS4IuxkO1ek1q/vjAW3tiEuThwpQc+34V
mFiZ4AThLJYYW+MNGD0cUP/s0cYnQaaEdlkFUGSnepVgEnrRyWw+pFnYKdUChepH
OyK+MtS5oj4sVXYsR2kWM0V4uHQEGHHTiASRjPxITWE3GaFC/YAw/uNcmoAaRBMp
RF4UwA0QUBnEQKkDNrfHy79jbr1IPUxhojv2OgIKwF2H4nO2xOWXIbD1tSgvxzof
IurfxDYQwTeUeFMriYpbn18XC6NI2ww3IK81nazXRFe77TZ3xNNE4aM97STKuEAI
+REOm6NcEJKM2RGCO7eB/g49TQiwXyXjSHgQtv3sUQQ7gPwkrULqbNL2MNpQfbty
zLTXBJgh69OIg1/fYPELGvrT5ouqo4reGYqSJTY5KMeMGGjK4RJ7ObT+Mjd+kr1l
iLXoTUlrHEGPgkJ8Pr0eiyhkLMwgKeA/RHgjZhJx3w3+Al0MOFpjKEF0WSNuRqYS
UDuTuNzvDzGueyuQIHPKBLics7mQa72GLAHz76pfQwKy7LapB9K18OE5pXZYkHaX
7frVcm3Xf+kC+yR0fe/HT5V9QdZhNpps5PlRDhQHKto4mz4I+kmYqJ+mhXA7DB02
+L9sThlcRL1kOSMPhZ1Mrg/v/LMe5qc4f71SEl64JLTSY2iSu0o9xih4DvHQgDj8
l3firF06/hxn6O37gKDpFi1kiQ8RAzEW6sE0AGu/YRGg1tU0MA/IrdIgSUXmEoGn
LrRxr0T3UW32yN6mPY0oxtRzkiF928cFpMPSsiOYXSn/lkU+If2OP82hmhZaek6y
gUKMYm/A5JFCVFNl/lJ08cnuPKvUHW0fqU/NZOWOckG7pbNWtpTZsiZKBuiUfb8s
GQb/QE+nqM8Q8RWJQulx8LEGrKKSOU3xPnfvgPBkXtQuNBw63ts/AU+v61U42+mj
rZdpHKd4HZiNG2r5pRECNvXuGlXaeLPcmpCBfx6z0b3xjVossfHGX09BuwuA+iLk
ffUg1pDBW/Em/Axm+Y4Hh84ty43lfGV1c/U6tp9Qje7RqEh7WMmEyC9gGYN+y6Zf
KA0W3AN7l5oXQFBzTOgHVRKUgApMKsPoF9S4ugOHVF/Ih+wqJ11AHyn7y/pVSG2Z
EZHxea0KBbcVAA8Zs7c+4bZ7b3okPT0oTl/vs8gLNGEPG513PmS9hHH54gkddWEk
VGlpC34rYmRI9jNEVIb5Cnnx9io+/49I1dIHvRgugbjpQ0sJRhQWzeF2/7c0GHYJ
rLbW98KwaEIRKn4A/4DmVfR+AGB6Bxy1LRuj0g/T/njfgfOB8uKSZmUEbFjU2Gzz
6P/B4/HlK7qwtcW/03tz+2xYAvitPDfWD6/APYvRq6OHDRpPRAniUESsbzc/V7pK
Ni/kPAhLD/dYUCOxyRf+H00vN72YvZhBAj2RggsPiBEwPBjTdHBqUug6FcxNQIhb
wMj+ABLfK9yDzaVy8TUwYwsv+Y+BF5MM+sXydgH6PGznsOawCegkxm8nDD3pvePR
nTcInT53bfq7hzbr7fW75q44h2bJEdoxj3eTePGerNVg1O11cp+Mzk9tdOyr6Fpx
YfNWVsj5XSMv1ulVEeLsWjp+xL4yGdlbyncChPffxNJhcfGRCTYYu6KVyjy2caRc
5MwHNnm4onHwgZfqoIixDAV3Sa30dCIzybB7H3xfUy9O9rEYP8TrZWOklax3SDHZ
0s3axzi7nQo4ih8Mh0fP2ZBR3zPtgccdbAMOMFz7MlodNG8yXD5fMzzpZV/c2uE/
DR8PkMIfxh8qghKTHzYtNRkkU+SSUCPWzEUw2Wf6kYrlJ+stX2rlCv8d7njPA4Uu
pQwCjY8fNiScyRyGPWI8iwISIqjow6vFG3HU+Z5CvX+Faw1u9aKYM0ThMlFPBAvp
sRfrrA3gluy4e41mrOLLeGCsOn66nXauY8+tJTF0OjVRXqfLrCEO9YruwcyzRHhd
yvfNcLNTowLSK1v4MCwGnh/teqfmWLqweL4zR7jd29whEB4FqBbH+LxO+15enChL
y8I3GojHPDFpKAamuhyvzTXnHT9wbbQ4LEruDOlH7S7WhJzJq3rEGscKFH1T1VUc
huJZlAsuWzAJq+Zfr82PUL4bBLXFOQtO+fShVZ4rSETPSwHrncZ2fc8VUMT8dyTT
+oVzknqQHlWVCWKJO1zSQekrYMsL9zX2Q7nsXamv2IIKWaYjv5eK//s/w9sGJe2B
+TCM0uN2MnYcSSR0NyJsdwql98iYA6X1SFLcpTAaNxwbZDt9S1iq6V5I8VrlUAAd
xqyYgBWJp5RIx/Uz051useuuQ7kKu5gmx1aGELfRrKRLMXQNF+AnXCsV39b1Sk+3
/ZP/iYMx5OtP34BAHmVmUALp63JD8vibEx8d/r3tKnSfdeKSci6MsgvJIA6KFSbt
co+H3QmaPxhxhSdblAPnu6+CP5EC7HOadxwgs1asx6dkJPjbvtWdw0nsKN7hy+9p
R50Vpp5uYRICBycaKBYGqeZgIuKhEc22R+k2tdIf5gwPr9jMtQb3p2pfWzwAK1m5
Z90pAURYJFuK0xlCwrfFNPC6XWWwTWqReheQL6r91bbx9oNP5550wGNARBS2Zc4o
PTZjw4Z2g/z7l6l2GM0xL3jt1L8Y/UNQOg3bLLBQEe1IXFT5zOYoHkwACrqO9HGU
wMOnAhq4BqGxWxucvP/lwT5gQRFwjF2ayw+LcE9UMwD1nGNMKgVomYYSyFAJNIwL
wM3eMtGwYwh5yjr5Kpgz5XT51TUGCUC3Xrm2AZPpHuIgeThqnF5RW0cJeXqe8L6s
lPYqtVRUoyhrmnrZKtJJZy9dqqzttUZyC3uiaRhmtbeNR8KnMb6dMCXIopX/EYJb
gpLGou6HAA6vTtMPrkBrfQs0Ae27V1UIeUKS5Gz8aYsa4FcmXmni/4/cMghY8LWC
qkHoxMUkUbdHgIyTT8TZlcDVcfp52Igq/agG9Qb+QP3soZGFX9AhvfKBGN0iB8cH
gBpTlQebi85byZmPZE8a4zHfOlWdwU04JF69qBDmPlfL6Py9AOwq+fYEnjnNWERI
PMdQtM3mqv4LLZb9BXGd76A+1oFttn3ruP+BhPWIfqHLJ49JpslY6/dAJVDLbD5q
LzdCc1aJoaVTtTzpvGpOyd+VC71hRTtpqmcFiIZUmgzjcbijuRmidXUAW6SB/81E
NNazCqiA3j3JFAqU6CsSK/ZMGSfY409ZPXG4KmKDCfSXKnTeiJKb4FS3MuxTrLTC
NAQWpzxW1TvfMYMY19qv5XE5rGZRk3mt7n7nfOpNKX6RW7+89uuzDYL/y8WNq1Vz
AFoqCzelPf7VG39iB5HfY29a17XdcuIp4+dtJszc3AXGgbvmjjl59+0x1mAVsQxx
FbJ6yqhG90UFQpl+XoFVICNKyRn4ff43Sar2kwj7/JIEaFqEJay8/0SLqlv5w+U5
6k/HPsmavtpNoG7ogVqp2utS+8/Iq4hmRNKXsa28krLkIft+TRipayK6cXIryelV
b4jIwupGJDKM2CN6DPjEDIv+Ah3adx2gPKgDB/QxwIl0t/8v0sPd3Cv+yWoku+xu
xP7I2cqWUWhDkYwVJvrZ8+8boDdYNF/BsNBQ+p7GkOw7EwVDRBLQKfKASLKXBahP
ICA4qxbh8PoPnvqfR9PWRFdPApjroYbLscUnWHlOyh6AM0hDcgY8QRRJjCLCN6oW
tkwtbU+C9C6DWJLhbITLrMnMZXAGLz9Td1qH+yV9JKu7f3vMdsvebLVGzp227ucE
65057gspjsCcDo1UlK1bamt2r63lZXhjauJlD2DNjY09aZBr99B9jTGzbvn2LzOY
7CPTOdgsJ+gk6IEoF6a/qnpDtdd/+xy6ul+QnV1DNgXZjHHxV/MQgFZvUVbMCFyh
XQNVv5bZ4A0kik2Rxa46P4/av+O3YP6nDQFyHdUNhJW2u9S160RWelHVwpa+sDZr
9yR7jOYZOITiQ+fBSbJnZKtAGcTfzG2rs0w1kpo9YnpiHMrJuS/TCPi2ccPf+Az/
ImcM8Wd5jmZdeR+ypqZPME7tqQUy6a7c0e2vrkLn4PsTZavDv6IXWRhPDjnJdFHf
sXc+rw5ToqQZo720vuCKd8KFXEZQmNjPK6GEkMwO9u7ylRQ/1p5ZM3O0mVqM7B9s
q2AlumOz6oT3N4jwA4EobLmud168tAukfQ0tq3sTNOP+nu4d2Klr0G4yc382vHWA
b1YiVOTNdMseWtSiCzpUSeHAJZYy6d54kZ2IkGYgHWVkq0w7hM3PKDy0sGXMGHwL
qnmyjGciwOPZr91AJbfHdkqzFq2AC7Ob/M2mJvwUi0sLN6V/5hFiHMQJVmhIGVWZ
yFcR3H3zuPyXLVQvcfd4GGft+wHqdQRnwfotn6Qf9pn8PO2Urc9TvDmpYUyIO9Bx
EFmJyzNydbkspyB4lvwIkU0zbCFtSBOLdaRPkjP/nnGDW6v+Pu3CrlRgkWePWfe7
lVahKmhE9h18HO7S7p+BJwKHUFvVbnXuDAqwyqQGXB4T1cWPlhIQ1PBudz4MEeDt
RSeBjU615SjbJetE7NftJr9hKH/z8ElSejG7zT7Wzw1MhTIxkac4NU15RGLok+g6
LtIep9yigUbCRtxhXpoYCtCbXI+Lt3IRvqEthnby8hHSkH06mCJc513q//E0DPs5
GMuTOWO+Pq9prJfg802CUKfjkrSbkMja6Zmbd8pLkr6CWt/Vz5qBAjUrpicz0MWa
ZzXGSy9JuXhOrDSTMS49eGJgZNgu9BWaPE/VzJQfBCIGG40tHLlMXUCNBru/h91b
NFPgxYAgbJOn0JOFC0d6OptvG/mleagLNgXRMlwWDOiajWwei23lHRzuEpw8fLbi
blwJn4PzU5t0HMmMPR87740FeL887tpOHFX8V4yDRNmp8/hU4WCJwPQBvH5NnZXV
ni2HBd2Phngkd5V0Y1JKTIjHe/iXmdE8YaS0mjFH0z3m+HeN3rQJDy8I6F520vY/
FefkpbbqaxThtgZHOCsnnyXRjHR0nP+RCXOvRNqcrIFfTOPn02MkYvVpm8gNRMjE
tT0adcAAHfNj/9s9+kVNhY6NKvFlu8hm41O0mN+XfHvUvJ3wn8FwVi/VkkL4ClI0
UwPRmZwXwnGssa9TKK4UhKLf4EOCu/Fv/Um6IPdCdzp+AXY80ZaOozdrHMSK3M0U
/qUKEIvChLpwH9QfvsQXOZSJz6Iux2R0GxlpUk0dy1te771OeCr8z9DwCrnMNNko
EwNf0jlL1cuLbQzTb+nqe/KRCSuE+w5DzPLNPT7Pkr0rbqVlqlVygv7YnxnYbROD
0SLl9eNvDdknl6F6l/I7oVhNm8wzuuy8VChZxOrEKZW9c471tJNO4PDduL1fLSv8
RETKS/VbHmV6e0MNmtBuS7RxErWoUNubSbl6tBi4f+XAbmFn+3zvan3/0ODU2zVY
p0jPxVX7ymRaxq0eFevXNoLR/UwccjGbU1S1eCFtJx3I2diWEN4pvhjM1iY8auRV
360wnByPFOBhbjbDIn4LDJdLtVE4aDdvBlpoPdlCsLtQYwguq4s6cUIuQGTtxPs8
lq/X4gj3fLIYTIQ7MZtuZiCEYU7cfCyMl1mDlk/d2lysB66KcV358Bm7rveaQUh4
tfrGrakQl09EhCICjNvsDDkgvxULhodSNGZ4YXmrNtORB1xRkPV6rU3bwZ9bZ7El
hav98XKObCBLjhCJVq0Li/0ggSUHs0W2aB7PImKvSbhtieru2ttDmKfxwgCrshNy
riNTiwdSodP5yxVJawRccfqrM5CqtgQpwwXqpvt/Nwn4YqD0+9/7lLKJoW2sIMlw
EcHWEictXiJurwAs3yzUeNof920EVGACOkwXis6hqzrNO2BUUNFxCaACtqck9XkC
fqOi0gIDYPUQx6qkNPqjeRP9c1Uoq/dDym1opDE+ACjSWp6U4j7xNUSF+QIWHNyw
qBN0VWHThhlQmQKDRIlbf3OJdHsHKr00l+jK4SFxCc8xUnB6JvtNKshNi9jRBwMF
fSxs5U86xrp++nxi/OJjnic4S6YHy3DdFwA/inteGuDhDAUdHlfcqQTl7OHbFT6j
awLYktaM01dIHP5KOr1cDOJ6RQm6BDWS08MPyDuFC0oCujSsa/ypirropBFS003r
YQn5sSGkG1bjuMRjfoMVtA7KMueBAnfRcW2fBzuIsfH9Ve+zG5eTcpH8bUv1gGR/
VpFKqrg8lsMrCIIFqui8E3v/4xMlSYA56//NVWup5wEqM2TXj4wdkdhUBqdneRLl
tEnPXyBg8nDMl9O776OF2hNaURHHcc3KH/Hk0Uh56swRIgy6vaG8I5GaZgChl3yk
wv2kkKyAnfCCfXjr+87kfUy9v3/iDGbzH+o1enzo1qWECtCp74dY2WXh1AKYrl4j
knwOhPYjSsC/vWH/etN0iUiUkQDvYAuRNfeHrHUt0KYCwaIZFMsc7cdAgQhLkm/C
fhqxQOYLwc8IW9kllCwgeW7+qFNZlzae+0hoDTG/S6CrXwCCAP4Xlf43TUpaEJ2S
brLrwxJ3kto6J9uZ5WzVZktMqv1Dy8qCR2IanBZ5RYX+BRmeOwxF3PzsqNNFtb8a
iVlm0ON06K/2evBKgXU3J+QNvfgON8lDtENHIMVpH0DoXh92obM2THW/gS2FO/qN
9G6Mj/DIxMMJnHRcNnLw1eLAaQIjlW9whcIFaLtsNrm6HxTPAc/djn8mlD3vwwXF
XyFmzxLtOo7D5Of9aOW+ZztkxywgqlYdNqTkKOVod2G47NzLA2CxNwbkEP5JcT6P
DIyyvFLyFEZJEu/N7TpKXgbKv02MDr9piEGO5FKmkJhExXytkh7CRbKXBFvbP+dR
2BTzmZBQIWZYmwWDZE/a3XVXPlsDpq65pHiMwtbWdJ8eEFA+rsH7IW4AmIKIbzDM
xaxYEavW6Ck/EC1Ho+PwZOPA+6M2kfEiHC27CvSNwF3pRoMwCEp/6+22qMrx8aIk
rlUdqXW/vzb5ZCvogg9g0bomgF3fKVZmvycScAFFD2HTVqYzb6ufl3fn5cFgitbn
U/lioiIoH2ghoncUiiioNHOVrxLQ+1Imrp5MK8vWNZHLiT/kmI78MvVJxGixaxkB
gSdVr3LJW4oI6p2EFWPaoVHLIVlvEXIrA6pbYu5naLojKLoNxf4m9N1SzwPfHi+G
pEKQFIrcBC/ABGbOUdBbZiY6DzYi0Ry1HaQt+JiSFBX3j0KUm97hRJw/gMil7Lch
F1ox0VEZ5ggrJlOqoZPmYu1epmvEcK5EHa7ZO9yHXGrwVHjH71bx7Nd6ePOTrMrD
j6MDSGm3XAK5bROc4Xn+V4Jhym3Ep0irFHewJ+3jEJ1KppRoyQiYkWMPTNAampb3
S6Vq9nCA5y2y3nyfEtOOWL7C3k6QDVM35yocDjHcba8rBumLzYMzlR8h86lCjpkI
xVJyDYb0ilyGFMr2cFZvtgmO8wHMb0Pyd+dl9gJ2CjwWQg5qy31pGzDSwGYQeBv8
j+38zE5B2wSzsA6u2A39kGLahEyt55JkXRIkVgxtgL8u4DaGIgr58D27RPJm+Ogc
2oyQ8pmihvMSxPQgYKiKZOiFsUrC2sfgO9LGiru6+Zn7E/IX0VaaKKcsttJrmhzB
CYwojRg9G4Woo3eMJLi4IlZV++8w+YyKorf6njFWPo82a9KVPX6IioBpyCemSNUO
IoTKTFwMg4w35QnPsYR74E2IE7Jyf5pPTwdzQk6daTci4EQKYlbjJ40r5SZO0A3M
SfjUMkNM0QfLqRS2Wvo6FEd/dtiMC595IdGza5Cj2EbqGE103GzVKVKPDRfoPBty
MpRR8Y8oJAf9bjjcVhm266WG/ds7MlEYommZYXrPKkQZRSk702cmDYrxlLMqCtGJ
g0Ggv9qncrDij2hy5v3RhAf4vAjb4KWZadgU6Xj/sJauMwR/C0tck8DiIi1bzD2I
oyJfyRns+H9WH/MQrfGqcmqyQapAy0Zup/vJmtLutiwUleNDW8p3TldxvzZ9atmu
+qem9sEVDRAonRkUgmp5huPM8AveqM0WyIezFYJqzdNAEUXgRQHVAF6HHOHYed02
5Y1dzPoToy5DkRmhfKzYZPtWk3cyjuR/2Z1lGMBR+X/XhS2tnYIxDJXnkPEJzPnX
JDromG71J/jxWwurfeqNW6pzc0zXCn0bCL97t8wKsT2F+f3cCA5rahHyL58imO5f
Q9fL4gqICQdRFXLu6hAm5VStSL6SIdCxcpa86jvEpkjT4VB97phHC4ChSCIcZyxc
A+uobNsSfs9HaMAKf6DpZZhNE4HdaJI21Y0oTewOs0L3KLEdpczHmaa+80p6SVOq
STX4KG10f3ETwotsycJJnTLRqjbkG6HRDqSsSzoHhAWpeq1J8p6LyXKrjq+TXe1v
zQY+kbmGJQcN332gZ46oB+TFBuOCxbutSF3fzud3fAvKjTmZmMeX4c4I2z3ye869
c48J9QBOyF4lApZMd+DYzwqIjKRD8sUjUerJt+QbVHzBziWa725r0uUvFYQwpVv0
ExSmnHL+DRjzeEulHafkjFHlON9690EtQnxqF5o7ckn8OzKm53kz2I3wPrk2bn6F
4NEtas/3vF/E6YL/UyPmofpusF1mqhKuOndce9KVclO9hwUolhfSX3Lrsp+5pJDL
rwLBJIImrdLpZtfqHQMW7oMEBBvh5Rarvb3AmAUuFpupJduZab4680NC9DYsgrz+
TElMV5Dv8KGKdezOwaSVWtYCgr4/Z4QR2/KbSMuycfNVB+zIJFFzKJqIvbCno7PW
N/sN8bMOt5JiI0QLmwHBqvD/cOBLRsAyzTcS8T3PYbAQfwB2UoPY6jQ4MBnKghIZ
0MM7Z0m3s76/a5ZTG2Gk1+/vxA/Mr61HEdL9ALpcxAioWPRYlqUVh9UKkmGhrHP4
GczkX+oUQ0nj1SCiyDFAoIxfQjEVoRLm04QzYY/dy8F32jPLvp6PDMIAxtfzbYnu
MEoq+9v0m5pMlyk8iprAnAzcHFdUl5Dk0ISXzGi1GHpna6NFZKNwPD6PnIW7aiSV
DPdfPSrql/0GtqBBHPo2+q26xUziq+ZZRwIJsCYsRc3JwsKIvOvANpMjlA38WBMZ
7q1TD76U5VlLg5H7tLJtNa8q82Skx2YImC+A8zrF0NmZFeD/qUyQLbkTCBQbhtPn
g+U6n3dlP1nqWsF2pIuORcEvIEYemkAPISRUMdR8Vfw2rMVUDyMiioPcU5OePzwn
d/tLLK+mVCr2/L1mALnlGEt6XM8uAipbXJctDAerzTnIzRAQ++wTQd+Ina+gbI5b
ie9nCwrzmBpwpXMc6RdGsCzE5bfgASPxL+l0AG1Ftm/1eqkVo0xRSaxZ8WSpCu+n
dDX5CFAY3FBygFBApnAS2yyIzcpyJqOkLLnnHY7jporwpvJkuPhMzy0QOsdOFm1P
had0IjSKQZ167lwTxy/pncz5U+gTN/TRhXxNcPX61rguCUN1KFrKHOo2dv17VaUf
dRYbi5M/g7k0bLRPMoQN7AaCyx+hHXUn3xS3PWCFVloZC99+rnoXLZOZb0iROmsI
KnB/wE5oGuqArGxdUxwzw+mbIfe37W8aEPpJjma3MjvVxh4QSGcEEHwIUtBx1Wvh
CvwjO4kOPUb2xmc1jrseb7F1SFXdarOCR7HZXIQfG3ONuWj0+c0Aina5CUInAEVk
l726rwVco6jZPP/GHsySK3O4/FZ2RsAT7mZ9539NtQXUv2mp/zRQflSDixgfZeK4
5xwpFUF/+ikdpRS7SjsYHzgbh4+KSJjTZU+xVnjOLmWID5FZpc0w0BXsrbj1Zuyl
OEDLCwHy3zkQIh9bn2QXPR0O1BjcNWy9vguZtwGnzi5ND3wDX2Bf7jmwerbJYqoO
VWhYwdrw18TPyhwjMk6VfTKnnVeUvRqZHWvWD6Jorbjt+SSU+nRK4lX0z6GWj1wD
CIzUnaOBkdt5sSVJV9f3tPFIAhjTUjPunvflD57Ggcag5vNSh9tnW45xyAfOzPcY
k1xG0pKtmObLqBCf4SB7wn2oQmVNt5ilqbUq2H5u9fZZIGfWR89Z+C3MTnQg7V4K
BrIrBo8tvskH7MZUr1yQFbh3lqtSIszHMkwhuQW1Op2sx5Klvv9EBEotxR15QN2M
vtMfNEy/jnvsekH3WTHJvFPZXOtjQZnwaYlL9dSV30KH37/fNykrlBIfp19wZe/A
Fud1i4p+4SUrqaINAfJS3xuRhkbDFy8aT3jnteH0kdeAXKmlbtLXpv1jcFSqND17
dJzV2KWL2wVTe4EreK4qIA3cBeB/mKfXB2+Okdhw1RChxZ0dsrJdw+gBBp3dPHlb
BEQjPSz3wlkUUXpjcHUa2aMhu+sNkoPjgwGPNissS47w4mOSOTOAD23cewRHsTz8
L9FSbTiF4yoIw0z+vnguw0GEmCIkggZZvfDxsiSq5rLIPJkWdkY2v5GKjk5+yNmi
WwlJLv8mcEA7GkWvN1vSEJ/vK605E3S4s6GANbBm6N5xB2X08rZzBQsf+Sah+Ejf
XF3aM62v5yoMmvUCNhsZ2uGQ0QKHDpBm1rjNekLNy+BE9lxjD9rvhFzIvYTkPDZU
h/n75QmhabFKaxw8MFnHWMdyG6Wqfqd4Om3U6Z1ArPfQxcBDcKWPzSFTFK6oRVor
u1La5fOH9WpOy/Ds6rd/QOwiS58u+siBtEXW0w5E/CV9hmAf3HA2pxvNuh6lX8M+
xh1mbgyTYHr4m+s1aNxW7zISXgdAGMwjJTbxfUO+WJfZ+2P58f9IIYMCcIpICdjk
p36edkj6BZ+BfQzXBxnV4UdDP3vo45iht4oHkAPO2t+kwh0vSEFVpN482xLWHlgX
hvpAIYBNHWRKCmgwzm0UrXiyvCEFoynNe/60mpYJJTEr1ARm0fzUlm0fjkgpwKDK
26UWw3DCl4SvbvzLgfb7E4EtDbHR/YkTCu7Aim6ImL6smgmcvZUZqF99Ae+BHYwE
kJKQcfkxa+/VlvRlrxjl7SNsx63vCfOWqcqEsNN87HWg1uKzkPUSgTlL+6JRvvIk
QjDhK8oSLcUTiNggGBWoSK8oHCXKXX1alnr4Meq38NE7sUo11lmeVduxEfPqo2Yh
ZfSIia7iEU7Nye7rR+EcfIEd0etxp5PyTPYjJOeed9v+xBigR4co2xCK6RdiABia
plZMVJhVhQGLNezYP9+cUvXtDJ47M+X559U5FmzUz2y9ZihME7Lg2LvR01xDMlc4
KVgxfD8ka52SosgRZ25NxGZwYoMbwXDxfkJI2xVAkGagze7swkt5vO8XkdRpO3ec
U0N9VLl+qzB/bZ0iNsUngc3HTiIMVgIdOEAOos1DjiNLlzv7HfEpUbs6EnV3sIlU
jTpuG8PB8pyDLYCyHl7Z4e43l1fEx0hic4Rd2Hc4h7VWlOznYgU1zeF9uYDJI0qR
wHSwijLLQ1pu+P0u4F6zpOBAEcuRWG/nDJFztJBO/1HpBktds7emtPuhWu8kr2sU
SnYxpbYIo9/+9TAQbZ0/RBigc2POhPVY6j0wTyRs4DDixrNmPlf1j5L89i2OY/Vv
6UJoW8/SLf9X4tfpsULGXzFkFNEKG7RDgS03yLCwam7kTV7UhU3k73R0VcilK9vg
Z7MNzfvU+X+EpxS5BfPU+BU22iaWJimZDrhviVfBm67vXq3/IDAhMK2JlzD+F8sS
kIPuNRkaXPJQd8rjoIYHig4m1bT9G7dO1cfJOvQjoT7xxsmmNtyEMQIpLTZE9LPU
lla4kXytNL92QYpcuQB92xLf+NS4P1PzLOfgDv6+aj/b+Dzv8n6rLtW0AOuQ0PI/
sT28ejhDuqIKhjBhh3Igu+ZEiLRe/Nnthv9asdR1mzavytr3v6DQ4DA986zTLiv5
DYQ+OgE063qUx3f41BJyXYGYQ/Yh+oCkV5dSZVhZflOy17tzW36IXz3PDXYMN0yA
W1Gf0lxs/D1TP2U968+B5fRxkbjKY7bU+PdgxDlt5rK2L5mBze7Rp0Xl4EVjIa+r
isyiWFkQv02CCBsf5xtPZtqN4vyPydIlFq3VJhFwiWCxuDtaUBwb0M9ZlLLY46F8
dO1UX/gZvE3gkqd/lDN64wHknVhxTRx6hfpOhJl9g7ROwdB3HMXB1tbfyfgPdnaV
ufuL7TEjtxP/CVVI2STn71bxAh+JaAWWBZiy4a1Op5w4SHzqUtxr49O3gm8Imcqr
CEbVn6/I+dn6qKOdcn8vgg2zr86QKOPv11Ysf6PMKYkz9+j5nF6MuaOU1MwOgtHW
SUYQyTaNyqmCfCd6jiOKwCHJNPS1oH0/wQuevrQV7Fvm+rF2wCw5SipPg4gmW14W
Eb0xE7eto2ocKrO49FXoO45n6owcOusBksvTTBGPScoTmDmntb0FLINskpUqXwKQ
wdbDF0X2jCR0DmopCBFbO+nMHP85qt8CX59m3UF8qEJN4CTJpf3hG3gcvze9h+Eh
YSMFGTTWe82JF94McyZ/gmHinB1nkN2hUQNuZq05xrll4dK6l6QiUzu46f/G0gDg
i3C2eK91qjvWgpm84NGmYpetW6Q/GIjzGu6GUNB2XdK8ecwxVt1decS62/umMmtm
PErQieu5xy1ytn7eyImf1fGel7XjlCa63CXLRME6OIsd/EWYGu7mlPYWJccNJyA6
Uo/NINkYO4PeIK2z2kTu5uCXKQPsyTATkIKxsZfetXLc34pqhJubn5jtSMWj9tIQ
gA8ZECgnxLDeX1RUlQw9nDWtAcxzNWVCfv3EtzuNWgZyriU8FV+VM83cy7OLCVyL
AVyIAg+amwOmfAr+lpkx6xb/hmX5OgPvaXYF4yMSUthkuhgedl5Em1ig872MA2NE
+KWEhV76n3g2hzJc9GipBcwFZfT73qxgPqWXiKoHgdOl9vthWy5AbgsqZrvP/eFc
kNrlpbYQBnzO+mo9drvdRKxqu3zah+/Tvg9FFT64xB3ekzFPetiDtXICfgH03lBD
Dn5sNVhXUDt5Wl353G2N26TVdf8H5s6dRt9dsjNtRnWVaUb0oFLQnVTYintQh7vp
/H7yNmC6fP4ow2ClEVe1B/0STz+DyR/05td5wVDxu3e78hli1ogtjP/0SYaomNmW
jo4lWlJP2fF3uFre2BHUvYAbV6NwCXkNLAflJeZkLRB70/lLQX+5fnkcflTkSEP0
EUpf9DKZvcrdxRW3L6JKA+EUJwuZ5k09qGTpwX83U1Lv4glfSeGDK0OoKWfI1yI7
LvjZXD1IiG8v7LJPJUJL20qm1xyEj0U7vOybBuuLwgifBUrQHtVDDuBq8MGJ6Dzt
rtZQlEIHqWAgmH3rBMipaDz+ZezZLyYWTxy7puNwQqJEi7DEFS3WeiPHAPJ38MzL
Ac6IV4qtbQPp6kzQA4/Xncj26QreZU5Lq4Fv8ishfcQTDhXw9Ma6ctXfQLccvMrN
sFDKZMQ9hptNdkE1r1ucznOCdiLs67FbPYzVOjaE3ol/G4IadWbzVPXLrorSMEyQ
fsVeUUfWzX+rNIDKDNmfuEmwJyofUr7iIlJoclgxj5Ma3WmXq6vuRZjlPTE/bSUV
E5kcM180AMJw8cYPNQ+OKykQO9ZBgBsRb0wPeKyCEfcVRgoan2isPUnCics78zYV
6WRe4/EochdWE8Bx2PMzLjBVBCBKmNLIYUyz8YnVvqHBvs4ZuE/MfHNuEm6O4dHU
hZ0piyM8j5MnMeZZTEGnv3FLjLHq56mkYjCtqYZPxw6CFHl7INnpUz3xjK9KRNJG
xMDGobPHmvfKwymSvwhlhQZlPpQfQ0gKTSdkulWCrlVFiC+CoZZxor0p4V+L41v3
YTsy6b6NZLJjC2nIQlA7DDEBnKwBEslbaINQdgXHWdNskXO5+5XgL5qz26iPB7Kv
LeiI7ysmyz42dntsI6/9F5JONzkdcbDsIUU0to5QaQjm+eQRmY67g+L687NiuDJQ
/nUlfPt0HRbwwaCg2ToNqFhHX+PvZOG/lK39rFv7OIXbXR2bdjcAtMRw6hRqto7t
1xDO9DlrqylaPWlt1jPxD/W5mgmFfb9em1OIznltowVwSw6HMSZ0vo/Jrp1JWcE1
FAoTRFm7Ag5+Xl2B24+D7v7wD72cEPvafYYmXjXWK9TUkZ0yEX+5I2L9SNTTiR8d
sRPnfKWmxmY4X9jlvV5MrQxtOQJue453k5q4Fb4RLXyRvfJJRka0ivNrq8wcUggF
9/wYbrVvDEdTCtv+bJJNHec6K+a32vOlNc/nNZ3SXgJgnIY4Fnda8kNLQxBdY+s6
PsmbgwGA0Nkjuw/hPxg1yLbsvyjoZyKw/SRA1Hkogjl4xTbfFQlDKD/uyktydaFV
fbLysE/Uif+eOcUq+5wQeQs522UOU64FM6ynCLTes9mGItd7JJg0JNNDc2dQAgy7
pYO+A/d7i3KbecG6I/9i8IwKrLwbwGtaxviBaQW0G2EzIeVjasZxaZE93KcEWXKV
RomGVag9F3ekrMF52i0Ysex+E5RUUCgnW9QtSJ8yjK1wVW/SCE1rZG7tVoPFYpSb
bcTn482Upk024Y1dXLg7uy3P8Xa9XGRo6QiQzY9U0qKbyl731hf89JJEPZh31j5v
UM3DyoAcRlgf+yjph9DfyOF6y7oWZQD6SPqpiN64FwKGDppSHkzXS44JRR0GQYsQ
H445SUNlnsZ5jSn9i+Gp3OIfd6610xUOgGI2xt6/gpjbjAn8dKqIj9AzxAdxGfyB
+T8hJfJGt4N/DDsGz6/0BfyUiQhYeiisMPOOzkhY8ac2kCN6Tozx7dgDUTWLv9gL
kz9xAYQGnxW2FSGWncU6yQGM3yczNn/I6FJWAjsPBQV6dTGUio/N/BPhiab9lCIh
mU8W/Io39E2M4+ahdKUzdZ1iFB4MNsmuFtw9r5UF33vqxErtnGDUnHuhFU4bgtAz
A+dIMbtM258QP9K9gfRfgRN8GUiDvH4i8W/7Fe8fYSu8rahst6ytAdNamYTTfvQ4
b/TGTqbitVa/VxOOSNeqfdv4ipUJr7hknwMVJA9LQVcY1wfRDa4gIo4rO5STjyec
LbdgAAr/BrD7qgZYnwxFgMAHX2eGSP+F/RSJ51a+K1VZeuXBScC3K26R3OyN+edv
9lWIqEOwuFnjAulv9hr+eU4dbPEecYyq/fmlRPnhBm88Vzz7/FAenQGykWGuujj+
lVkrOMxsHr9jCV1C2xw1SL/8SCMVVqZhOtBb6+TXpY/r6IkOuogmSBUbskms5QMU
uEwsedV5QTy1FGtmqNJlej0WVGMSwI/dTIYeGfmYhg7gnt6aZEuyW/+L/v6QyaGx
DEaPjx/wvTcN4dxRrEdUPbfEQdDxCp6X/NQYt680X3DRCFKSCOb+ORs/LSHwmc6u
IliMnXROQlhPMrXm/I8SWllxdlRJAjZ1VSkIgoFs0lEVFYghD7Q2WH1yfaOmgK+I
UC9Y1Gg6KYhEmqfoXXbnSySW5bqxAqTw/v+amH9T64WI+VPquo4ezXGnOR/QyVij
MAC6+uhBNPfAtfODUiNzUOiK4Li4F4YFHcwB85ORmIL31RsK9VbqNJT48ucso/lJ
Wn0oSsf6aFsODNdOEU1Hksi3oRztvIyvkHDVhkOLowYVhLoAaiVJS0TC4f2QAJB9
XND++QYu94c913eRRLwDhsZcbFUJYsOGzV0lSPt9msfXshLAMeWHdXqdLD5Rcf+K
hlB2JTeDJ3BNwGeBy9lflkOb39Rp5XH1+P4zRTxpWwtSJfWwNhdc4H6C/skLeHcv
TWJLRfIxpIaB6/IHaNsgX8S7JwG2oQJDqkplkJgmcqbYq7dRnaBALZYWDpb5vnvW
CPh5ThbNMdkgRNMRnmiKPaRcGs7Ty/bdlhlCF7NWlweFbDVxlZi8ctNDywQXrwTN
oMnFt+V4Sq2mN07xwX6Ng+Wtn6YMBBqL0qR66pBWmoAl+Iwxj0v/33bBIzq7MVbM
ZbF+ujcRktcGH2WHA1jku4GyY8QiZzt2JA+Hna74g1P4h+nTQglYf6SPprSKEWZ/
2UgSC2mGCF9HzUOp6k3LQ2FsFzAGfHRwDxpoz8sEl9tWRau/SUAXkg/jSfHfuPHI
M3QUbhRmeNb5fhJSIzxBWA5l8jmuwGj/pat45oxvPezsx9OhtAlxR2lfjYCSf1b6
Q6Fl9jBnQHJsWCNXOQZKFwXUCo9bKrZMd8AukY3y1Ql/Rbpg9o7SomyCd+PiUral
NGIhtt04EwAjQkRIN6pVYw2sz36OIEPBJ+CDSf0dAzZCjSriLAr510mckQT78xjw
2uWm1IHplkaZa0tt02eBEFpkyTlKmoe3BClwajw1TOa7njGEi6o8ZBAekdbMikXg
8OKk4byeQ4y9C+wHfqI5gce3HU2sLtHYteoIH65BC1uH0plNdjPbQRQEYYNryq8c
PkOFeohwxpKI/4auE69G9/5qHTmj93D7IPPD9ZVf/PX9CVAzw1MvDfsoZQka5oci
+3BJGo1ZxRomd/2MeOp/LZ8VVFblvoue7odZjOqPNOWFD9GS4jinl+nVLwtwxxya
gMtsxhDKTBC7tezkcc+LZUwSPFN3eF8bWZcDcDeFQqzHKDdiU3846acXEaNd7bdw
s5rs6F6OYHWKZVyh9wPsPu3CC9ZI6jAxgeyp7XQVnM86NbF5YzUmKHPI+VjxSO8T
3bvZcFKqh2IUrrvBTdTYQKgEnJDOtDXy+3jjZl3iheIadpws0rR4PsfyfKWL5RFm
YzaDDeENXIz/nDQLPqxJKvCsMhudaAcgL3EFHu2S9kTZsTNlSW3OseGBECQex41F
Keno9pZMcVm54qoH9xAn2AIo+hVHb4etNd4H4s2adGqEWSN4vtoRkhdIm7xVlE4P
Mg2AcVqnE9jhzFrFOsP0zDExO3PlOoHvzCB28E6vcT5h3FwDufPj8wr9rSmK/CiL
CQ5XKHcH68CQCuQdQly3s2dEljEKibYifyiKlkfvaY5A1RYW55s6dzDSX8vZ5fNT
l06PjybMfwPHPFpgT35GePQ0mRCwT9ike9ZM3D2KGYFILR7y/3VktNihIPo14D/o
hzFgPXpsAymt8Xv67FRWoUuVsWyHZqnP+667cveGUWQpXPU1/vOVKweGsKqCaDvM
69tfIvum0IGPQZmad9WL6+Yvs3tcc8QGMu/EQgW5fYlCBXW6DPneqb0snTs+gJj5
FHe9Y3ejF4CM5E4pvDc4G1ENCds9yqT2y+Cb8BSXoi52j5SFEJz9xRgeQ9ace6RB
mdp5aXjmHmxspHDuYmtc5RFMVGoZlAE/7ArAj9GQc2gRtJ0Igt1mGiYiU6BGOXfS
PwFrHpf+nZB+N1q1HAK46ZwrpsLhETYudv94f2I5A76X2A+y8w7I14T3Rn4BsYkR
7C7STWJXAGd6MMw6iLco+bnZTY4/ilg0qNKhIXBTOzFrhyXMU2USjG/dpYslN5yx
B5oDZ2bzIvweHGW2PAqNCkB61CIQBz0hGJMT6fZ58fagBZ/JCSUk5Wv90DhJLOpQ
JJcXSdHxq+tlKMdbjflsBbVqbOamiZegKdKbgzgU2RQ4grzB4adwV1Pav+UfW4HE
SOzstfnviYa/vxDN3bXOsf9R91u17Z3MKzvHO4hLp6IoytPvzCHlFVBJv9n8Hh7x
VomExkmtMVqHuPwaGuED6Y/h6QOovT/HRdH+zBmh2W5t/t5bpd+NS4snsBxXqGW1
bhqtl3+IdAIKDu8dDC+sHlNm2JV2fshv2vV5k/frKfCkhFi6NK3TKf0Kw9bvVqmB
Hg++skcU1/hlKiWh2Ah3HoiWGtRnXZgxHRvO/N1IytM0bli3XZtJ/LgHa5HNiGQX
OxtDb/CYsh/ZsrQ9ccZ2M2K02UFihbCwrilerHNhlqNBbYpksVUJkKapF1ikTVWf
cFIkXU025Zi0O9vwVpj6ue4vGlF+mOIfcvcstMyonl1Jff+ASRyT2yJTI/IzM6ny
yND6+4+5mxe3tJFMkt1+koGnQ8HwfR1M29PO9pGqyyViYJYQSrq4ce2jLslaJmiO
SIcsXG077oklD9ub3KFO+qthpCZ3kL8WorllYq0jH8AD2UrgDrVgrt9xcCBJMNGH
vNMr+RFnoBvcyZrefGNjGlBCRNwuyc6lTYdN+I8nLupcghhTRhAgrpsMbF03NKY/
AXYZL4XIZfPjiiKueFA2MzVINNoCf3IICAx9J9I2tlSiQSo4O46pZ4yhO00N7DQ2
NSo+eoNsuze5SDIKTfINFrHks/HTS9oPiBR8WNHD1WBLqOMbf0I1gBjrn3Hh9Vw+
UaLOVECpU1ZlBSvPS6g6aQw8ke0l84UsD36geXTX5eG1jC23UCHfQI55VW1/xVCd
0f8VwJTPQuYXxUPzOfkSaShlUzGcOOe8+H+mu0AEjjv5S1EvQJT3LRMwC0HbFNV0
zw3112lIX1rAbQfXB+gKlDpYXCNAyRPHEwp01K8/nUuawXlXJAWLfrStElVQfhDd
HXQijLQibv/QRqHorPYMswZDmVHqMDF4pSgoafz3dTlSYBmDKfcuwDs9jwBD3TQb
1m5rGx3qSTdBRJG5THBo80zrVeQ9K/28R4LcSINhmVpZaTIX0ERN1EPg6sArBjdR
wZQgtfvW5rlt09gjOh2VmzLPO1P4i89mp7XJ+DclxkuH720d+rEjxO/vDzkTH6mD
Cr8sT4grsrR6U8KPrw5Cjus78Cee5PU9Z4Up9rtH/3wQ2lFoZXvEgc0P/uR2XNtf
XoK6AC0A9NnCBzMEQ0WZyoz8LOYnJe4m3NRsP/XFNFd9p6oj/yMpL8Wdzpg3Vksm
vABvmK0jmFmqne/qXBDU5xHAMvGOc9bv2ucXGrp1f+Wdt+FiIN6uSyWWZGPTnUeG
BVR1DFIER2U+Gy/JKlZi2rwIysfucLug1ZHMn9MnY4xli/ir48S9bcH1aI1ni0Ix
UJ0yioi2onVxU9vvIApsiBhGjfojj3WLsakcBurPWbjFsXy1YGAL4EtwI75beGf8
2pvRf+8hFh/7hg0bMNlrI1lxB5ZYjkvn2ss/m+moHBEuqZmjBXBPiCQkJwyM8gMT
bUrvgGqgEHCJmRSMvAdaGiQw9O3hMEqT7RWWElS7ynJYXUfw8A2MIwGh+0q2+pF/
RGp37htaxDz0B4O9DVMIdLVPhdiLacU2fESyz2BLbOjH6GrlyoBQpTHoeK0NND/T
7EfSIDR1PCEOuRgK/7XYtFbBQ7Skq/0kHIAw8FN1UwbUCHOL399CYxULjxRluqaW
5nTy5BvnkJV+02DGB5twguwK4mtkW/7F0LRMJQ22lf3I9FWHuDX3mTjHPKohTsNI
9jo+/i8ovMb2OST8uP1vhIOs8wxZMHKHBEJseurq/fyhdCKc+lTjSLJU4Wy5hIrx
LBUAyhoBE9dqzCRutydvH+0LXCfo+g7E7nbTVLzN9+uyAJrNFKylllxh5aDlgX9/
nLAo6NA/2WW9RrbI34xYr9Bm4uCWM5KKntn/MU8uAsZmhFfwY+oMcmFPxdVae+m1
2dnVyGvlMSHzYQXDFgc/YX0YNlPGjgOQ/kTE4t9qwIiTBJGHfJSCJFWzKQYnskW5
W5YyNzZSiJslmvXZZI6f1pexdhwoq8qhgnlqrr7nyErzHvQwwrXc2jNt0iWlOKcF
vALmBxOa9Jgdfw5XyQJcyvILlef4X1LF9XthJiKW5nU3eBmNtlZgdQmLfcEr0oTx
zaWzQ3wLdKP711Ri9+JJkVnraVouW5e+ywwhqA+rSj1p8wCYgaLUyTU/tPUbeLl+
+JF5GM0A1J46K9lidIqC2PPxSJwrcCi3BPR1P3Y2fQIhSZ/ft9AWic0xVCAn5zoh
/ppPASbWujj2u4ndXV+qPOvR/3jonC6zUF+xEwe1QPj16/HJ7HV9nfdf8OUP7KfP
Q7Ho7O/V+suvpqky40RK1Jt5yc9Py4RyWC1dj3+bJPzswO4pmEzfUhzXSAy9Je6H
iq2uL7kLAwjqi/PnJKfceyoeyh8rHukRi+aWB79aQQykGNBZ1QGctPtkPyIQ6Wv9
n9q2wAewJx1Qh9Y5TFX8n9LNQZ8y+ydP4lXdXLaZvaa44A+7/g9ZpkbHdwj1Wofu
LpNdbf2IU1ZHC8BO2/Wra0XuZTqAS2cBoSgEibOz1xHwgQ8hXMqJvoIaCr88LXxg
JkLWsnW9i23BoUX38bZgl5dIg6RVzUo9gZeriGwtnlfPWK+H1KU5YWm4riRKsx8S
F4j5aKpyB4LSXA6Kidqg8cmGj3DCB7DhyK1naKo5jU6L5gW2Cimxzbwkn23uHxE2
RgHpyEJZAzL96PlBP3fL/v9QjCQZgwc4pcCKckvqYeGWTRvijZ+uJPHR8h94C1HL
E+TnOp2+5W5At57SuEXJ99Ts/MuGYMGWJ3C3pEOB1vus6SvNiUQLwqiOUOiUUNVI
0Hz3GO0BQP0dq9Bc8KOnzOl5KY2HVBtK/sGRt9G67dXwa1v+94nqtscBTS709UI0
BtC/Pl1Dk7MF27sni4Tg/B1Q5tccYFyCXA1rROk43b5/ZQR/hFTluEdve+y7Pggc
BrrNA2eK7heupapdHaXZcafeP+J4zuhuHPmuOjUijNiCDpGMq+4BpobvNZS4mr3d
gE/+HVHjT3OywJ1K1epV0uGSNNzA+XFO3LUz6KQWRlkQoEsOeFIuQzm9vcu2XDjM
KWMd/onHJ4+e4Y3qLOS8AztFUp1EL43/T8euQVFa26z7zqmq6pnwtr19+kIjPhLk
HPDW6rnbouMqlf1nfsW2KVz8zgAqyA7e4dJuoyjZJFGerHJoBg+yepWZR8UdNeav
87UhaRoYbApUF6IjQyQs1x49RQ29NtVwG70ZMz3yHw/J1yGQRSPv5jh1u39lt8YS
zdEPjtCJoZK9ZRowqssm3LD2KC2QP1GmD0peJsTO6/iQaAEePMVZfn7FoydD6V4q
VMWwZGVbrLv/qc2G1U8o/esTa7BNq9kMpKwgIxf+9x3sbHG86Bh6owzVn/BVMU3S
IpCDt5wnskLzdFTQMXkCK2tyRsXSSAcv3Cju3ZceHPrgjTuLbgKQulhGlRVBAo93
GWg/seIfXGMjM4hghIUa4nDYSZ6owKBFIRcu+P7uwyi1b+ZMkyzyFCtwUQAAJRQc
4oMdWS7TEF5bYcngQvbOIEcymSDbE1luuQjH95xCzQoFMN7N7QY/8aDNftISH0jV
K/LqX3Ri05z01vwm/9nj4cUVnnghXfslDRs6oIOaJ3iqJeffIFCj8VlZz2zNzvq9
fAxJdGHC9Re1K5Z/55c1G23hLCV70xj81acbaaErIBLN4qE3Im5+4X58KHEyY0cl
K4kwOXIoPBjrYbzPWncF0d0s2BGuu10O9MvaMRTrp19FuBZWw14cqempPuOfug8j
BMpfqbAf4ImHh3WfmD3n+pfZzexDomM4DOkgiC3fZ2kF4plofRohipB+sJtv0/8b
JiM83dMJm+7ZOlHA7Vny7LvKZyrEJWczoFYtsPk0v36x524TsZxXm1/1ChH40DPl
ZoDe51wMAZ+VfCXF1/kaHSM5/egTkSFVWWa5n0tQ+Tz/79kFxQpw7n+q/4Ld9JrE
9mEPKj6wm8ujnMrznzLUW6/uwx3MK7V9Fo8J18aFKBsstEsszVUVwaHHlTInnujf
BSqzEFhxj0ly9916MEKD1jELQVv901tIyUPtKnVTpwK6kmtNjpnTYwp5/onhOUty
zcVEOiXlupaYNgtqFKnOcAp/OGnXXzkZ0mZ1a3Kr3T+ZVgZLb5hkKgs8MZclGDZe
nr2ESFAXudch94cH8Gc5GgxbkrMJaPVurWdyC7U5d/yoxv262NyD+fKgdzeaazSR
XWa0ZdevMovjs/NTa1ezStVYi3LaG6zEBZSY9G6e62rp0ojWeUkgk30cVSr4bK2s
mZL0pSlStKjMdaGQ3Lw2HcsjjL49vVgE6mVCrMDODdVOLoLL0wJQy1MssbMItBWQ
/gXKZeHKLUnj5Jtk6j95wKHKmiV2HAjoidD4MeTb07Z9xS4YgLve8FrdkC4xU6H3
egEEBYN/bmk+qDhY7Aevk9+HGJM4Bl+p0C/kll3orDZfrmAOTrngBeUe1z79f9mb
AmodAM4uDOXFOiPlDYFnJxIpapZ6eoidzFXIdUzuWdfHBUCrOZwxxYD8i1tXm4+j
XkxNx48+ab9GR38QVf+jotwZeT0S/ZCHteXkNonjnjd0NVljEv7NV0fMx/1GJXy7
lTcwWCRqSDuSXMn01W1KvNMtPIOfDWhQKmdFik/IqTveKhB/Ycx79NX91G9buan6
9tlxnCYbZf1P/I6hW0xGvz0GQZD6AxmdI5/7+ofexefGRdvSLEraKy4X+HbEjlNf
+N4UcEyyzGJ13dQEtrFQUyT93Q5LGLJsjbaiURR506zGr/E5vPDx6d1yPWd+oO4V
3XO3zg29jnJHCphOZ61Sksp39bwbj6nLCJWDSqDFAvWuzlhZVgkD0dRJmP3OA3BY
a2L06v9BRObU1aUtyojddK2LQe+1avYs3K6xEE7Qb6EZLlsRDbn7TIEobrwfe/BL
xdsExaVS5uiaahu7J47T9QbXIvqKietaJmFAeBp75qqKxJTDn9DsLcQ5tETPl2qb
skO4RlzlkDlcKM/0Z3zz6Kou/39cdLNh6wQlg/NzFymZ7/BrhiMpkyPcOVHlQd4Q
eYaiM5IsOuxkOS93OCDsZnYNgmx0ZS7UON/WmtPNvE2f1g7y0mXXBP7BJ9m+ak/B
LrXrYs+Ea0osRGlrnfR0pUSsVxYSqIIr3A+kPO9SQPFCRBezuzSqt9S7N9ZfR7v8
OjuBcNnlk5nuCHXvYRJpFC/o6lI3PT642ES5KL6T+Ma803y1kZAwBMDxi9Kt1rAE
D5kigN83AkcOl92zT76AN1NJLQiJ/S9VvYFVHtccCDnDjkmryw4ZzEEkGUaonz/R
0QabdFWFoxsxb5iXspGyXdMBtxaOI9NGU0LF1oBTT/NW7faJKH5bwjO6fUyGbLFs
evRudk1uXqgQRDj/vqxfslm4RqfzQ1OrZZQwvYuF5UIBAtccarw99VFKY1r2+OQj
MkKzYv5cjPTTTAdmi3Dym0+5Qc0vzfYM/VtdIGU2JKypwtrgFHJrc1U/v8NH/BOu
x2+2BNL4p3/P7mKHtBnPvgcIuceZal6XOCaH8KvaKxdNP24UtecSEnIrclcT57Ya
okRuG9IBmNUN+VVuf6ctct/upvJqFixI2D454DkfZLse0Pz6N/0m03mDmKUqwRE8
5H/QdzF6xQMKIiCixaAkEUfApnoNQAZmX7BWotERasAxzy4vFetueambvb/OUFfB
cVIDNvMm1BFACPfzUM5uEBtJJtjxLhfjzldMGSvx8YCS064O11jwPDfBL467yhQK
Mqu4SPzBDefg96cssKWxiB/hJO4Hilz+3o5ShGSuMrTkydwA7T29sIZ3SPVL2eGF
DRs0yGZeMHnwDFBVKtjIl9U+cUOC5a8r8F97HruWqnjn8g0X+5H2MmFGWnIaaWj1
oumlc4Lt+zfVTmCoemMsIQtbO+DLTzhDJu2RFCzR2vn+ruRpGOGy3mVr4WgfWH1p
FTtQoZ6S5U/Cgggp1qKOZN02pUcIKaaFymgW6FCNGAaTc22KO6rP6rsXu1gUAGJH
E8DY+4SqRNIUe5kUXJhXDIkRpAGLrdMB+ljGd6oQtMXoIvT6n+SWgIhuCkg6qdIs
z5TCphiOzwOzJgHk8hrCINCQmj6z27TvnZErb5GTDk2/NO6FG7k37oREPwGyIBvW
clMXvQEjLA/wOpn1JJIfVFARf2AZU2Ks8DqqJmoJ/bEyL4Y8C4M+MvI3OUD/uzoN
cRpIdSWAbVyxCni5cNvD2rGE/iyrffu87lE+MuYmjbcN9bZ6T2hpSCyoOVk0I7lF
Nih+3FIUEk9N1jBwyDj7BqQ/BnzU9T00GN+uNdZW0zOnfhzHB0gOByDBx1oBbde8
/xeHM6hGB5aPIjv0oUsHQjoRCip/EKnCmDE2uhOO7UB8Cb74mv7yUMugVMCtJfz6
FxZGk/y1eNQ1/Op/5YqXV5OpXW1oGzHcX9F0lP6s7CvXrklC1LtNAlGzDV/OiW2W
NduZqtcbUdfpyFPuKn+jbYazxRyzIr5q/W51lBvdduohkIf+dV8qxFnJzdBE8LJ8
K5RFW2mcG2hHqAZv8o+sskWzgAA0aqVb2hz612RkMsFCwo8+ykhJSOoWGnNRSYv1
nlGwIIDBPTKxck3NhFVTTxGrB/LBzkcr/mF/7a2XW+1q9nlxN2FQMPLAAbhIIi8I
xt6gx/W0rvE8IrMPEH5aIo9iAJ1JmDqWvfyiKqWLcHj5FOz/Bwwbbq02GFfmuYWj
sEGEitWQboDZoGwhchaP3MHe8e04CMFNs5N/W1RBkl9h0UORE5ASrVBjPD7PAWPH
wpzu4vIgd/xEb9Fmx6xGMUiACvyAwgPXBksD3WVPADnt7Syqs2Jf3RlEujhlOBmh
sY5OoDrtL/PRhoizNNn8t7Gwerw7fklWEMykTSpBlX3U+GL2cJZRXq7FkmJE2aos
OBCht1bLiFA0kViSTPGiaNhGNMbv7GHid6B9yjiXO5jaUqWostMsfxpl46Xz/QJa
wsSya3BuRuC/8K749NCCnfz2FofW7nHq8LLFBT82GWpbRsnywTgdCp6hvcMXhpUF
c2SY81q8HTPnGHEjmKs73uGghbCWX93Q/Hfgg9cSkk0RBmeL0dIshAHYxIIHEN2C
/emtROL774fwSUgcYxQ4UmcEi+N4lxdMlezTK1Jzhhr374eIGiurBV7IK9AWD8h5
b3oYJV3v9FAx2pKBcoIiQ6XzGKW3/j0J1fn8k2J2Dks4060HMBJhqjNHjkvuWDbs
Q6ucg9Sy2DCXn71BVTnBQWAyERsooLn4MY+B7xY6oP2Aoqmo/zHcd6r5X5WZxqXg
JOlildbxLiQNW2qpUTu8LO3O8nbIOoglYBJptE7TSmEeaC+eVKN4Uw+1OeXd0JF/
590VjxxBF92spc0r+Bjui8VtAqRsOJe0mbWzNwGIbusiGBUFL4TqL7M5GdsHcaNt
bLOOGSsx1bPwHzjBLG2dChtw/3mTJLk/j/BIKg3tiN4h1YPK/Y9C6snTdatu6RnV
a/bXfHljDAyN0zseGE2Yoa7DIIo0S06lkvQzzioZQg6qtgfvGffkN+jqngy4QQb1
19xkM2mQiOHSlofz0HeNOGQWRNLU3A/xvDFD49nlHfAXyrEs/I1nh5fU5nnGSBk8
qCmhwt49Mq5759Sz0QG6L9IaqSQTS7+KGGG7FvCOK69vjorCUZWCy4j3oPvN7xL8
holqu+1q1Ztytu2cUUrVTAFPtp/6jytLLu+H42iDORc7tamKygqYzew+jPiHti2b
nhZF3HTRsHMtZIia6hC56r1AN3sNFnzjcwR0Axq/Pmi+PNyoWvDHwS0KOneItRPa
ZMcmioysDkiMHfaFfvkQpymB35wFonO9v33PT13t9f5MyKo7zLhGmy9DxMyz4zil
XHjYYoeOnrXzQA5d4HFkWjs3CmxIPgle1zAzTwlnMyYRNz6qfHCI9+F1AJhlrjgi
22hgjvMzh7ZML3sDUszfXRnnvdozPI5MmJ/cnoILLIJHOvfqhTExg7qEdAnOySLU
sl8++ed5A47+UMdX5ARe+WaMM9yBqXc8VvtZhcMFF10GlQMK7D/gqwRt+dMllOAM
UkCFwHWOFOaVOVtYH4e0bL1zoKMR1wK/bfTj77k3Kgdy6iLwpIdybGtb3fHXw1sH
YoYcDcTqOIslUkPHvahSWuDnQLmEIt50Lr26zq5A9AFKgICxiCvw41rrqJ0KcAU0
ZKeSApRb8AnFQM2JTkO2CmLPab+Kn9T3pPRJQRGz5Zzj18OR4BLb/tJhzlGWwRb1
d70oy/v5K7Py7EcO/OWZcAbzFh+qcwwLruWY9Mt56nQSuBvMpYKDscYjCdoXfGcu
j0hcdI+dz1XNLpn5DUY/4KsgMBqYipVBlvfcJW2dXdm4qmnaAwtbL9f6VKRR7EYv
FfRV8qBVom0lAebzrARdPqJnK8PVdT+3lePc1+RpaicY0uUo2CywsW+E5mSqIpjR
TiQPF8ue5IOq5hpycY4rlytvR26oOLBOhJzPPwunScJqjgHEQMcWPP2HtH+CJ5VS
tZORYz5n4wpzmVFIhRfLhWR8MmdEg5sR5uHNaCe9DuS6FGExMZcGyCkQkywFgruv
IhukoYKimLw3ipbmRF9DRieV179NSfvwOVsdhUsoV2h807SoyPlQPOZ/NFs+MfLH
9x+udV+WchPD7okRAGI0ny/6PN8HKQIWYWidpllKcx/v3syfHU7KjqkG3OglMKaZ
gGZU6eMMitrMZQjEtEpKHa2sPRDapeli8dd7esIeoo6DQVwBuVmj0gARfqC1xZjD
PVYQIchLiiDJ5AJ0YofjxMAa0o9IsPdGFQf6y9tHRPmhlCB7vs6/yi9bvrnUoSuX
+t2shAZ/RquLFMVvZSFchpFNjv1YYf/Y1bgppEItyVTc2wCGMbxJnDBTMHAuQg21
g4JQvbYotIU8lvxkkSU0N1kKB3QZuGf6PzpSJ3ivrnvGz9T0+KT8hYkk2PqfHmLl
MllgBpZEsYaRM121uGo4SWPp2JqrxfhwvS48MreJGMsFc8JPU2lctg7MKGTnGWkJ
jYXH89BwuQEUVUNe3AlyJAvmDdKjpVjpDIzCdB4wkNux06/vlmRU0FkUz51vXz+b
9YUy+3PGsazAdQEpI/voitSCtxIbaL75L6qPSB3aNHB+Sn/5x+DyPdKa6f1GlUT1
C2CFiVirvcKWc36uEvGD96zWPErz1Bp2ULa2iJ/X571iUvkbZbxJiFdNjRwGdK8h
NmimK1897XoH9a3e66o41t+7lpQoBnhoBfrtODzy2GyW3zOCc7CSt9BpP5k5I59y
gFXeIBX95/bzxixhCXsYqCRKXB1SiAt5iiBHlPL01JllT243WF2n39gsT+VoMUw/
tqaYQOV2K/MV2yuyw3dZE22rg07Cl+svbCoYidsfuKZeaDGHfQ78K2y843BuCl+S
auPDg7CxfWCrhRYFcb2pf2FdiAKEY0xXoUJ/UuXiNyTVnrYSyVomYddmurQbajRd
u4Yh6HKmW8/cSr8i0ZWbsJqc3DaXqrvKV3FOLc4aRh80KXRanaEUiJ1L9DQf+MES
XbHtqRn6TfX7kimBG7q+sLFCCCVDCsZG+VPkxqI317db237DMQCemO4WZQ6JIvfU
dD11+Kx4mVIwY29WgNa3GJzjwUfx49eRbU45vi9YXZaennOaINbxAEfJhlQqMMKE
qnlAGmkNUBPLOMJk5cZPNvucutMknxC8ZeWXw8JZyWlMNK/wnYaI9Yv08CQmmgNq
yly4eD5aMYCDwPI+/egOiyX6ANud1ByMEwcsJvq+qpwnSD8MYzyN03Kv3rEbdeGr
n9pMJB+GA4ASXpYJrxTox4jD/gst0Ivl55AIsHFtA4aLceDyHAxh+Z308R6zsRy7
2QPwKnFtTEnA+xMkkWlBfkKeTHbg25A/WqOmqwsRDVXjC4wLhLv7XKaSeQVBZygG
t4QtoGC5ZX8/PbhOUMpcqGH9LyksC2t0D7HA4y5iRDGTXeKmVrDyIkTk/WQGERef
9cPsvo7J7iODSxOEXEbBIEvqwlVyWGuktF6xs5ui4Rcn8uaV6oPceoIaXLgkWL0L
w5Ry0bxdu7DC1r3yyi4nu//Q6tOfBPm0NFaFLrU4FWm1fEi/6qI2vDUklTqhXLGs
/5839HJdKldKI8UgxEwhuWJzUjIgbJoCSesAMVvnzvTXSlERPSe1FwkGQj+vi1LM
E98jpp2C/VtHoT7KI3Lsd4xAziKjTZLDVWbieM3PnZmXGS67XQ74kj4NFwqzCuKU
IaaijJMb9mHE/J6Nv7gypQeHwnAjMFU0hdrFXUsPi6nfeWCwEekP+pYQvJ9PrelD
ce+2WiPMQLQgWJwjZzWRYUsdEncrB3UrKL0GQErQ86mljt3Ik5mmMuozfjTBSFpH
Zxv4j2EtKCCJD6guKlhpFMJ+2qsH37yhnEwyimro14IjjuAMhndqDHcQnQwFiv+l
R4ip1PjvwKvPXEPO2j8W3EnLjQ5NIuiJV8HGb1Yazc8Wbdnb1Q4KDMRXEsOFZj/H
FrE0WxvdnoFD5VucTwlE48ypVBAdkGNz3uYDgI840MhTatNmpOBzweDNz3iDLyAQ
b/lpDh3fc3efTNYIs1WeXN3xzQNFRf/dCcZsHpcyr04LpToVohscI68/pLhfZA0E
WkKQkKfvBjnWstbNTgx4yawaSF6HPEL+aNC//hFLhtvA//1E+d1Dv0i7DVj+5oto
7u6Xiwvqc5ZZ1Ze6/Fxhm/jf29Rrcuj5e0YEzIdl7Vj511vHwJX5I2GycugowGoz
YADX172s7+ohXoczflvV8pb1Wt4jEAQbkLW8Kk8ksfBCZiSR+aTvlX/tc9Fl8nzg
nblTD8hdtZMRvR0K6xHXo3FibsCHDU+w9dhuEL11Hije3qxDo+BSSsJAaIAh/7Of
YVwJ69wmJ2OF2mFDjaLRF+PoFKDlk8b8cO+z4TIZW0xi1XXimx1ea9hURwCH8Gfg
eZw9Ha7pnh7DQDrg31vEUIKf2z1oQ2u4LgQxzsoc62W/muulRFBa1uOmezSb4R9g
Js5in1X45BAxrw5w+6DU5XP6UmaJXohXM5VKIhe+8aJabLsBru3uLfIADotNBTXP
3bAe8J/ceAocxzfkIfdo6mfLedsnjeWv6qZQCx7bGexmMojLw7PVIbdZO8y9l7hT
kt0n/l04Wi2LinuQh3Bm42z3mZkOfc86P0kD+72GtR4nNXjd0V6nmANqTlTCa8tI
hVOOtIQ1tYPo+e73RW+27bde3wwMr1YbIc3DofJWrVaIP3CjSK4iIWG8von93LTp
CtVGDhUFgv5IQzFilChWpRiq0GFJJmF5eYYTbV9AWOj2VSNdsZBfyJ0+o0IKwVIT
Cg4Cer0THm5Dhbais5Ge1XT0AGu7Q7D5xjNVqRjBgJm6w2P9LTTCkRb0FLNqFWbP
OfOOBc+yGpAba4yRdFLg7/0Ut6QOz7ddOvLOpRKunbKoYqXpf9yN4RxmBRUQjNBd
UuKztwCafkYunvhnOq8tgZVymapZXiqsaVCp2CxGLxwf1fCf11fTLU9oyFg8bO0z
7m3KqruDuNLrbPDJDijwARVGNVxO0/A5E4ImaNQlusOLhwl9TRGm6eg4Uom/Dd52
6noOf7MPWuZcwvNTs9axX1/RdYGfklREAwb7ObN7uxvgmY48724ytJ1S1PsP91CU
rS31QVLoO4/y2lOatkzsqmhdgvkRMQncvHJHhCXO6zmXvmYDc7MNkyRYYdeKgTWu
JVJqI23ux6GUB6FKehi9g8kXVbybS1Ag09oZq05popHtJ2acuFldOYLFsZLuloKU
INSPJExalS05kn2kdip0cLh/Db7xQkFWJI8JnA/spLkwYhHCG1Ju8Fln1rIj/XA2
9AsYAb0qAobg0dKw90jvuvjOXvcFMCOYTUlj2nAfy96zCHRY+zQvIFZG4pJ6UgJh
MN6KZY4Zpd1n/KszUof/9ZlwOuvSZgDijFsal8H4dbQCkFHtWvzADCM5pecotNp0
BBvwyYO6Vy/vgr5GLKv/khmNNzgLyUAya58up6TNmciYXE5b6Pmq+mFHqX/keYrI
sQ+K5L2Yt/vSBIA3VP0e4Nq+E+W4f0uLm337Hk5mOtlmN3LmyThkJw/cof4XirF1
4NQD+5iP+H/E1npdrs1wJH5dly4/2ucpWBi3Q9HuijqcHsfvHeON4jUg52fWSooA
05oRxEMWCslg2r9MtZftlHCdQY7QEtJkn/+H+AqltfdDVSm1+K33sVjm8jx6ZZCm
YfB0swey/pWxNxGWKSBi03+ue7fkVwDoRf8F61VxWypH9Jn89ye9f+4wQInXRdhG
5MBb/RbBjoUBD6v7Ghci2ANaJOBZO8vmKovCglEXsZuoBTYpP1CH1kyYoWC/KIlw
a+MwTA2sg5H0Z25xIdLRe178SR5jDtPRoCZlOexrPYUSN+Tu92P7BN5ys013iAfb
RW+9igX7QT5qEd3vi1c3u9ZTMU99k7LKfmkvw1KEh3m5IWmkVVIyGsR6HTDs2nPR
qCMjWmnAV3l190DeehYPLgBObTL+ZqcrwkuAaRJxzkz9XiQs4Oo/3/b8IBXnhN+W
OlV3xirlEaYrf3rUqwJTPYc1Db9l57GXym4V7OP9+gDzSXBef+0waHgR6ps+GloV
W6ZXuQSdhjLgo99MFMUUqnxyvyG9sNpH851UcAaTy2zcO93pWjl8Ktsw/GQWcxiS
OYbwmQZB0kin/0llsXGlx+7ICLS48B1+wN/1Yjj3LcNoqTpmLfUDnhKeKeGTYbJk
P/PUUDuXsYhOMM3iLno6nR7bisFUPR5CIw6kyOnLvH/GSa+AXpwBdlo9/cbfJfAF
GNwG7OA8wamPlQlvj6hAAM/NvAqU37HJgE44aUWFG/P8jEiuXeXMx/FWS0WT5Yl+
2Afav4v0iUKSUzpLn+C0EpsgHMtqcr6vF8NTxytuUumY5iirqiab2kxL9+kvz/1i
KS/HcbxxoBVNIF5x+tm36x9Oa3LJB05CSl/ErtvrqxZ/31GZyR9vCVtc3Ged6oGE
e+jy2+CSas0+/KqD0zzOvsZHjHroK2f7bOiLfqIAEbvEWpWrtZl0OBD2woBrp74b
PDtbdb04VwZhXTWJJd5yTKlMfoGf7aA93JY5Sak3rUcGP3fHmy25ugzc88TNADZE
k0oyf9i/ADZITphcZ+HrfmmEsh2Xj6wy2jaaDjNhklnPdZB5DLKPmFmtX+VULsh2
39TLj4K25kmpOuCKZ83micGLuNpwTbu2X/IORAYPTRKA9llXsstR4ar5eYDdoqft
0Udary18aFy5hFQ+qJ26EdrZXcEGycc4TRoEsZVwSbFOZoE9ie1+vXMWCL6R3TRx
eDgkv2iYHEDVOxPIKd2iUI1MdmCh5AQFfPRhgvkAEF7HP1Gen/PyYEyiZycEarZ8
YdT4nSKytr9kyseAQ8Wo2TdbHYBdpsoRKQ8bYvySLtZ+C04GF2mEaI3wQXlB0peX
Xhgqz/zVebBayHRr2xMih56WNRTRnYUMn7ZmlKKfP/yOFDGuMcdKN+fhvB8fhidv
FCIWg5lKxjv6ozLW/qbS6BTC5wPRx/34YuueV/m81UFhHEIH9QNozWv1R4jmMXVx
db6oivo1Bts6moCJLhGa8XssivD0N4uHQ2maLnxSpOZEPSKPnHwehXqLUpJLXHkc
cdHxjxK0QSZCKmT3dTFQsbW8tA7D35PH4017DYSCjtjt+cG7lg6vd3ACIwh+QmKW
mp6sYew+Ma4gxur2s8h+b2E8evr1sbf+w9aFo/Y7PlgoxCQbYycEVcVDqUexhsXb
vGBldlBN4jDzF8odCsofMRWNudT33pnrQIRcdzocnxUKrd4xkPnONpXLaq18dFJj
Ht0w3uNOkrZZSAe9qla+/w0A7t8+AcWyXJYuEzOmzJCZ4rPUFn+Ex5i2Roj6vX/3
WxCr3+95osbIfcDJw1sde4/0I7GuK91J4SsGyCypJU7e7LfgvoCMjxGRDXv4dkHP
7UyqwRIsTNV1+BUUKCMXvG9AItTcfy5W8BObdzHM9vYHsjlHCTxVzITldGRhDo5q
IvcngeeNzDzdgis49TWZIL3QnOYLTgBP0eVhtRDL/chxpUA3sDb7MNMBvK0D2G5W
Z8Oqwtq6xcU59Ur6RnBu+YkGJegLYsOfD9BMbsa/pMrvrQSB2uwb7pLnT/wNCdW7
fMtEKMKalf34nf/JQWCvsYqgnZ/wMswyuOH24CpKQSNGd34b0FNdGW5gbOv4C6EJ
5qMlywCescypY/ZWdtQr5Gk0omtHtNVjxYHjpJDE0WbtVongncr1Otbtlqfu89nN
XADsaTPoLbrpiuFAH8JgINe2+xu46RJgrkM1aLOIKbee7ghKwQ0yboP7nUeLPHJr
jOps437IPn2lXEFy7peNg/KBGg3vzuOXDVPry6xKNzfdr2HltuVKN1pRykeddeo2
FpSoue5splzVo7ZMX8n1GH5P511SXfIHsfXP7ZYUCvqfMQkuBEOUnBWqKXOuA210
yZmuVsCHKWReQyq2TvnUxKNQdDi3V3cnPiioJL5keADcmbOSYzJ3ekZMFR9aJpBS
cGekf0SZPQbG9ascEFsLnqtabSrd+jCXbd8ChWmsxJf5pW4s0mDZM6d7/LamVC2B
Q/QlLD3pAC8Gk4bO8jWai1VDW+I2IYDHDuxeAYQRSy0jCwIY/AbVHJdraT8+820J
R1YE8LKwu1ieAOqnW9qHhKZufV8fB1gTS3j6C9O7XMAA3JQWXk/T7HG3F7IgiTJ0
mYcjQnESjQqnIRGkVlRqh7ESVfmdQetHlVmd5tjI5AqNbrRkVv+XPUUxgtrIVXI7
du+pmDgb06mBQPROTFtXSXYEFqBFdF9tyTmsJC1PHKTKl6sj3kWzuhFyhis84Bgc
vRfBNtfU5ZJTR3A/HHQygfEVgQfH5C3IwGfKECjsw2oZRj2nvTSob3ueZjKbUZi0
l801tghHAcxhpDwBar5AAuK1T2C1f6liSh123Wrztps/xt02rVxKBxzwAC3gG2lM
V0FT0Kwk5rkkYn81UQ6YEw+fbouOJrOqUIEsNHH0/xVDV/wk+AVRLbt7346Dl9oU
BOdYO9npQlnmJWpXGJI0WbKxfTvD3nOEJ0TAOe7kpPkz+/cuklWgKNcOfSw5Pkgh
51LNOye3Y6wlkhCsiOUR2wUBxfwUNcf9KZJf4NYw+B8RJm/Nu7Nq0aAlLtPBC7/p
uubyVtJsF5pSxXozQb1lN94spYpltD4meaAYd8HPNOEEvc7gEvsZMGFoYtswydEB
CEAZ5/mPwrhVpcq9IOWofu2X7Ih2mKMSeHbPsC3b6NeRV0NfT5ZTWMjnMVvw12OX
LPiRf1pkOqLAQBpoZzu57w5R58CqCX3jEDVpkjlWlp9AHsavFxe9sJAB3sh8/Vjz
L1o7H3oKpkGXCAHQoWkejVGzbUlQSKxnY6DHdOvqvSzD60BcO5I6xDYFFtprpJCf
0Fnc6VYD78KKqE4vZXIJQu0eMjmRamfm9pXlgvByIGTQz37X7nLvnQsD2G00x4ng
zOumt2tbBfRtIp1Nwcp8pSuo1se6S4GEs6cbRUa67UI3idUc176ORIW8IvaWyonT
DUviup8fAmi/fZCH35IHAwuCKd8piObVJrahFKHUAhzsHWse90b3iOFLYhvT5fdB
x3VS936eOHu76atGObuphYltNuwABqXRqBg9Ym6nxBtxjfShRFqtsniwihSAFiGL
5jH18tNdPwSWulck/xCT2jqdBaJDzzOWhPZwrAHB7LqJDvaAavX6soanWK55vay0
7K7bV4omQ78LofWT1xL0+Ocxr899YZkNppfIaA7PtXL/f9LXVdnc2gJAvm//SoKe
BT7xUppKJePJh2Xyp1Y2D7GlGEw2Vl9eJRkHsGEZ4CGr+qiHReenxnWWMmSXxcWA
3XPgHvdhNaRd7g3gQVRPZbylejWu2sh69CKw22BbF7I2g8gU+vKA8foER7o392t5
lJAIeQarRSAA6GKfLKjct/Q7oIPySmnx51PHlRtfoWg6l/Q5mQx5OVdYkCZuyE1m
oTMrWJ/kzTOQaIAq6bny78ZKlxUm/y354HZiVveCkQigo0K9f8I5gzE1pUEeXclq
jKXX/7beHsLQe4f3Oe7PltBCepiybWHbCs0fEBIzRz6umInu2oxRHqr697m1EYc+
Lmo09MvCNED11q9YSTNFzD08Kuuu6KvAYpLk7EG4jzh0p38hSonk8P+CJhfl/YWc
5oUSh6DAYn0SA6KZLXzNqBEl3zUjotlaLoeH2WH04JyWLOXRqw0AFtfIPtBq8Ebs
g0vLCqPRPSC6hWucHT9scpaTXU3eBuAEpY5zj9PA6Pazvxhqy6w/reTnQai4iYDd
AgijrhfTluLfCEMZNk+zHBhEyLQV4HSt1IXmfv4WjU78UY9TJusuA1A4M6iKGxTc
b/5d3Y0DC2ILHflyt4sz7k90G3Fb0CHoqktLYkz4D0Cjdvgr7cOAQjIRrORrRNDP
cePYjlRYZx5lF4llKKi9IzlX1BqDeKcPn2Xiz6kni89fIhZfdRjP4clKvf+FrJMY
9Ae0KREShKRVw2UdhzPcK8/czeB0WnhTDf+8Z0B2ord/PwUKBUlJC21ZWxSsAW1F
kpoqcqGmP8l5a3E1PFtUhBp7dCuCbsa1S7+dWnFK/7/hmWcdDZtPOvz7CBz/++2K
+0B0DrcKARPfE+yTL6MyXQjb9nNd1eSAcAv2ajeI+qNIoKLzQWy21IsWEqng1oxK
VvBxNj15gLmUYoiHyV4ZV912c//2C70bkBX8T2NJOm4Xm3exWG3+ndjUskVq7B8t
ADfF8oIdqmcbPVXvQUTTg9Eunn8jWKEVB74kCWib1MsA8NdaSkPs9suVSQ17Gt3z
sn5zvbFystXZYQP2CVoiJwyI06rTIgyNxJIpKI9kbHPwIiX7ValnApHaB4KC+A8M
2aqIHSDqCKX0amVm+8BRwUxIOi7vLDV9wFvb92rdZxvyrVqRcc892RxdWVa7+JoI
+ZgFGJieIbdIPGA/QEc5FP6bFnL+JhGzEMEzXgznJKtdBmrgtog3biT/f20VoSoK
OL/69JiAuGizdekLqE5X0Bv0s4O8QDcEQaLJoCvso2eZWrpIbb/D99mMVH3xVmTE
S5tnAZUYcM4DHNv6PqRl57sJGUXSvE31E0x2KZItz6D/rkR3TG8C+nfFRoFkbkf1
fcw7tMK419QqlB1wjf2Qx6KE2G1y5unbxAv5Kxvhdy5Da3sTgE0ZmFtobwwS5Hzn
306Ums4eeCh2MvNWCEJnpFf+HAVmG+jTGPtzV2D/p1H+ZwthSg8JGXbeUVI8NWmJ
coNcQc5td4kJrk3IVVFitQjxNuytcDtxhFhA7vvNPzA3KvEzveCn67sbwhNYQZif
AggrXFktZDrT8fvG9mRPIAKYV5DIeDPnT48KxRuh1Fxm/96Dm/SlbnQXoU3UQLjU
qKO3aWmLJjhQjZoQy9NAqy0Hz+83EIwYJLeEPavY8D7jPR0VqvpyzkCCiuEqb4e6
hce7K+n4jvU5rqEcWQ5N5ujK/TeZRXOX/DdpMXR8s8fa7hmF6NhGbBKdlIh+JjWi
igXr9qeGmBWTg4NKilOOiJZW7ady7zYMeYF7+rqgTXzcxAekbpjXr6qMv0ZkmVYz
xcAo9HJSIMfrLI/Hg7tvtYE8CagM+1ZQg///jbK3JXod7Ii+7/zienqBZ4gcg0YU
axmWKtEarTqCDj1RVtVepNmXFSqIRfuM5Cm8w53gRixIhDBa5XcJd+41HimbDnJl
WJMj3WM5RACDk6IyT1UBJKYR+Y7+PpcgiHCP4Vf1CCymF5xXsLokA529rCldAG05
Ssm+ARI5lsIsQkfhCX+pXhEnR5DsQ8+PLkGhMgctwmzHufp3yrMSebuW0xV0zHlB
PD8VSdiH3P8AvPEb7eIJ04KUWfdcsuxTnWKVh4OeFOhEdAR1f7T381e4DcuUdWg8
wFByFsPNtdUQ8xljJjR9ZjzJTBdtNQfBp7XexUsW+8e5M8C0tjhLSXLLyU+Gg2fX
Q5Za5VO3oct0ybrfMZYjGkfBxIy3Yvq1hNj7uxDxLtL2zbLSO00oKH14d/YG2EV0
PnezUW1YfY7apBMuoSALk6m7nQbWk6d9lbNMo0z8KojKqBD/F2BMGv7y//QpcPzl
SXL1lW9m+2ir9iBK3K9/J+5NPoWIi6mQwrjdozPGrVa33xBNUFQ5cSNAcLn9F5p2
J8fIxKDYi86gOZCQKrqnhfv4N7fOnin6uddsJSd5icm/faLfvib4zJF4aVQwxNdS
V1oxEwKWBO2J8PWyHELyjJVwhywHUpdfNYZeSj86zLnwDdkckYIXTVjgIt9BKOxE
Cel6InoNYjhdrJ9PdsUHgeTPpUjWGz/ujppZ7u8Q0m7D2pr6NdSmLc5E/BUmOnDi
Fc5P15/Wp403ztmsWB4ErdF/o+Q0uff9qsSN6zVx74UVl1//VRVlSmluqPAznJvz
7ZKSAdeTHY2Hg5y6UGf0GuOjgJOmh1ckM+ZRxcz3x+trHEPUuKHg3GTlVDqmWq2z
aeR87vnRWQuBKi0wklhs3RVumALX632B8/Qg41F7ebYUShAe565BP9WOSlF32mM4
QanPdqAo6TmM+KE3LgiVgbO6/+vE3ao8AQu1LDgYn96y6jiigRzVJ/9C2ZPSlY51
hH/80ixXLtjuoOxLcyjDpvrjxKurfY6yHKlQdtzDQk67ogQvppmJP8SG+P07wZNc
8s/HQ5stOyx8ECsbHtVcg/KBUyeSgAh9WmFosCWLla2ptJXipfOA/mw8vIKTXb4G
CHk7yQe4f9vAcOMZVL6s9TULF4rF6QXTpUWl3C+a2eYpoPCq/FI8ZeDZa2euLyK/
0OF+BvbvBDrJVVb1DV1hJi6jIyUronUGcLZFD5Dn56UGbchFIYKQWBkxSI6FypLs
GcGDm0M/FszB0rX/G7R+GaxPi/0uSXEDlv4hRjNmS28bXJm0OYB8y5twYojwL/B7
+Fod81NjpAiAvSkMAWk33ex1xqty7xasfZdHmqlBRpnl3vWlXQC7l+Vsw40B9crd
g3NUnNQo8uql9Or12Vzp1lcK8nkfiqugKRz85yb9dbaKvMexFtLHTswbKNJQM3f+
CuDkmTpEqgAy8d6j2/AKPSa3SDy0w9bbaiCRkRcz5yKf1HPfTbhgGMZuuTH0XYi7
XYaahbuunUC6qOgtuwc2chO7V2wnR+j6GbBF5lsWkT1esk1VzS6ziNGLK8PxfMub
eyaXR7K7ZuGa5Ua1+JgkMKe0oR18NYvbVzT09nzjuhJ+LQ8q0S4shjmf9SkM7p8y
uovCDKWkkRlgJPxqmL+iaLobzcfT2TGGJzXd08htSpoZjXdxWvJfB17Ux0bsCJ4K
n/ANZvK/hPI57gkkJWTPZHqallb4n22FwsqLzQDIlTnTt+v0ijTUzKmDtx1+ieHG
tE3lf3IkJh7V+tlhXoChGtLpf81SPPoVYkpZhttCjg5ePQgz39LwKIlN5zoQ4W9h
snqxxy4Zorw+M/xnKoBeD+bof8KF7mpDRg0mSyyONoCNBiXrze0u7EvNyauXGpLL
UpznpwN4cB5Gbb5lV3pcBctXyWB6p/d6mvg/IvKlinRSMu3ZNzfS7/0wqScLpbL2
4si68W4w80wOhvpxyzn37X7KDTkrsmH+FDuK2QRLYS+VIB4ZjV41FqCVJsSwQoii
P3ohCCyI89B7XUpylnqPQBRhXKho8phUTS+TC63G+VH3cgYngI4AxSoVV2slMUrg
ogwZASnDdDLWJkUdvlvWU73Z/8O1GfM5IIHdnbWrAOb7FDMEAMbo95U12mrrmZCD
z6r3h709lWmpodmmI5e8ZsByS2kWujYA71gfPRv9aHZbGkG3oeC7QqWC9jqExaG2
ZH/OzwjGT1kLl0PUilFo3Xf1VvG1jn98/2yvhvzNZATyhPYvI25tfIy2zeGuSn96
ybwQhuDry0VPirx8K2fGjo93alyUmUHM0an07bG99lEwZosoVj30tieY/kvbB+bu
ov4YpYnIrYYeWVtPUTe/Q76QRLdrFn9bjWgb1mq/YEeD8F43gZrn9Z4JUfC0MuQN
deuxeZLuh8ovKbLBnEwmKz1ZHepkhbDO/li9Iq/jI2toM5Nz905J98MWhd3L75xD
/aShcOKE2sVw/CIckPbZMGY3WhWidlpunArLeFcEB8kRPO37o/ok4Xda5qnOiy65
7OkdkFTQNUWEAMzT5XDnPTbSMGzHgZxuNHd13/4WVCbPksf4uOVabRCVplVclDuj
a7cQRCmEwfTCjSVXyPBo1YXb/A8dxGq2mur+56QiGWLjBBK+L+D3alLc5UGGmN07
eeNd4V1bqV2DhUGUSB2o7q9q+QARWwVZtXlaTkgkAJ6Pi9YdiQH1pN8RhZyRfReu
rNXk7e2ZcP1OpKWSxb1hmRm0huuv9wq3CapHxJMMYsFp09iRYHOC+rB+IR32/Zf/
rpO5uAXHQ0g/d5TEO2RMrX2oIZzVaRCAajc5cmjU7HiBv21OxH+qA+to+Iyc3sxy
jWU8Dx2ZvnpoBO+3Q3OXFwJ3zwfrRGJHHiGJMqJt6iCGb0wX7jhWloHwOGc24RLD
2XdQ7+z8430nSI7+/ZOR8cg8fImoWG44CcpfHwfVbfDZ7a2tPiyi8r3Nvy8LoGiP
o9hH0FRj+I1qtAjy8TgcSSZbFXn60GbH8KH3ZESjVf9kP7BbqWy04LXo9hEgiiYB
07AyIwE9mBweSfQHaUbo2NHc8ikoWGceXpEPm6z1NdmZ3Z0alnb/i0kFFN3d6JVt
lIYt6nvfnl/f7rabzoyCQSKB/uq3NjDuiYCuThTtTSUrZOhZAMZqSe9zuDSzz+0W
V2JeaNDlBZM4X++u7dmqWhC3x/3omJEeBMkUBnwJLHH2lSPAORA9rhtNpjatblCj
W2EPfES5++wqdNzKSR1tRo6xmRwlkHnipgRsi8mMukzVMRNUe2SY66z4TWaSCpTu
zLwy4hUeBJNM/YcbXmkomNggkF/vz0uoR3mNjUiGhzKSbZMcTNHJpbGjO90N0I5B
2bJ8Hi29KZHgQYaT9aiHQ+MknsKUtQTHZ6Q02UEsJfLQuuP9qy7/ou+v6+DEcBGY
d/YgSTo8eXuJ7w+CMbIs7WUkHZl/FuMXa70/qaED0g/oamHDNOrpzYnuCRb1xp+K
XlSRh387J4pCwrAh0Xc/L8noPOHnnNYZRrCOKPLwX6KE6u7Cy3fuKzY75mIwtz5v
ymCHZprDAamUEahrWk9z4tVx06NTtlWrjLIfLKmOzmaOIumk0s1W2oubMt2xF1Qg
gK4kzgVdTQlrOlqaepsUrCYOFeL+a8Mm4/+S/yWnXQgj5If7EI69pAPtF0erDLY0
uSSXuanWI4N+UDw3DWHbTf8vIuB+mG0bPWIJls97Ycj1azyAYxfe1R3evcon1lkW
9oWcwsiigB2MZldFXj/m5Pfus2iehm1Ojr2Jpj2BALOVEP36xjmhFhL+iK9tWPA/
DpJ52XZvbsR94a69MDJ9hcSKNveoSEqgqyKstYK7YSnZEW74n3JfpZWP499QJTm0
AsHIu8FyLAD/V97QMi80VHr8byUczjVsdFkkJ/GP/p0WHysdKIIieknCbMVX461t
M040zPApeOtYHoUENPsITXSG9GhGI2k11IrmD2Hj8erxOPBwVejp1plJnlxySSa6
XXxN40dptiJNdmIqMb7aCLev+WFBoE4V0U3HNNCicvJCMEaOhm1UXzTy0ue2QMl2
DwCG1jwQ1DdcSnLG4ap4tMPkoj3zT7rs6S6HXKatUR/cML7BWvdgsghfy6P9FNgW
tPZEUeUBGbV9GE9/eRauJYh4Lq83Wv9yTbFdD24ll5MyQVwnR6MAMNLluPaDVDRf
aXUBRiF0MwHtHGrhjht0ZwSE06BfzIX+Y8VHTmU67Cdihpn2IVMTuPeJix20iGWI
SEb8mzRon2XQZs2yEyDhJg04C3S527e573mkldKbykYve1/aIqvKElu5bYPmbhUb
auetryzDrW4sZxTac1DjoatqQRbcAq6S3xB7g/fpnbiBI7eJgaXB6FGah3iv0y6A
tvaNKxlcqoVYKqlsw05Mlx16DCt1zAappnozNsH3QGumL2mfN/9LBBxeaGvpwroa
kE4NlyD2JmVnzzEVTC4VmL52jPhQkWakkxu5HsLkinwCPIZ/7kIfda5DT7Uucyzn
Aae9Gs1PYztT+cOPP2GMvekTnas25xr+Vl4hQf0oaMAjsxWGekuw7OnlQOrZZUww
HcvrmtEyP8pLrhaPT4qSPD4CmJCV9EeN90rnSjCe3g45RNrrl05uO4eJKnjzGT++
NCwdtnkX/7JRomPI43eLwjE3Meg3ADB1vGdv3tJyxDZEe4+yKGtSdk4zfGZ7hHUc
pvg5H3PqHpbeKpzkzUS/ihvlKhn5bwEZNfFj8RFBB0gDSu9ouLJQw1pbYjSGPtC/
j6hqMR28HtxWZRfmITrqigmDbwpAVJa5oYvikuu8PsocyjoKxqqBlvc4nWbazoDZ
mIlDdv78DP1oRvfvuRQY1pujAmn1kOgLh6sLY+P0uBKVo6YDvyWEJXSE74YZ12eq
PNiXUYMLxFpdm62261NrTBXyfjMl8HNB0rURvHAUIX+7u2zR2A2K84jHP8AG9zVS
xYUWV69+ORGo4RKObx1GPatrfpPVsl8dUwQsU0p2OyGpWrlQ0VuL2lGWWAeWYoye
iVkr558hhSWHNTtQr3JBPr/Cy7Sxy4xZnowGjv+fq1XR5sHZ0DOYeoelFNVldbbj
BBXTxwdr9F7A1VEuCwK/ej1dbPTX2yo3+BLuyzO9ebmfaXFBh1jTbhlLF8Qwhcik
zXTJSYhNDtUgnfxtSk+3Z3XWicfxR0dLpQc2Y8DGutOUd9hAkZ/X4TxDOugrUrP8
hHMNyLaqsedQ+0qC5vPW7g7ErTTa33uNYzsWvFSnWezz6M92CLtUzfJMXjTzjUX7
7FT5sflE9WoSUxQ5/0i17fjJYCnFdToxFUv93ngfea0nv0fDc3NO2kCFnT8PNn/H
9RbwgCrnVAZZWZ6cwhpE/GS2QeSrD4umzSA2Mouf9C4LYZoAbt+nghoWN5Yq0gNy
eAbKMqqR+DdyU5MX/sogFq1HimenT17HoqXXqp31rz4VeBU2dtQ6c4rNeo06w8fp
vJbe+SmC0BgQtcoj7M4yusbHdkPaXb81IXFAqw1nFFgMGnIHUSSvWXnfJVADyELM
Wthqkit8RPGA+/tZcEbMS4r/YhxS8vYGG4iCPvbf7rgPsxIAN/16TlEWeQapwxNg
GVnFTSrKSH2EGAtkNLpL2V2rXhSWdN7hwx9O7goOcJHSQJPXn+Ag/giEuX3fnKfn
XZ8CuALOrIYOYy0ziO0KVeYSXdMCUY0Useqr5RJ4i0zklPJxNA4BuMgaUZPmimzY
+HDmQ44fO6pQsJnqGurnZbQsL8dx9Q4Huhv1Xc8dnCq5X6fTulFBC0K/2Z5Fxjdi
Eu9KO9ZGsipVqOHyxjMCcwC2DeKv1FA+4V9Arh00PNwaX4w4xenIfuRXbH37K4vv
0akTnAMoNhigL0/UBbHoXPJYzzcnGxt4ykYyIgdQzxHDFHIevtlryH3Bp6OVgnOD
w4KF+cS/cnBJir2xhw9kaKS759PHiJD/2Hk3vHURmj6aA6wghDupDqD8Qj8ENvcW
idXxKZQ/ixyyQu3hwFKU4EStOvaJo0GsYxr6tpPDqm1tv3CGCUhwq4nDJmbwcump
dmXzKvbcksH65L6B2CoxkKm7xzmW/lSE01g/e810GwPbjsjGVPwcpvSX8HwB0gOr
skBoXTiRXoMxhx3IJz6T9OYOWhU/p8vEWHPdr94PzV3Dq3+JUyKhXMkelQsO13An
KBf+hEwkHw5umN0+UbJ82ksH11KwfFqjgBwCxmDrREkWsjsDlZk4+FkEmUhgJbPW
8zog0qUqcXTtv/RtZVYInYHCmPFR5VlcOCNdUBj4v6TOAuX0VZVT4XNcu0F94u09
FpQSVdS8mQ19pLYDofws8YLc9wL2mJO5B3u4nN5HxVG+YBXtVh7UdLxUi/eqUo6z
mlkVXfeT0cKseOFLf+2ZAsGs2bYtGNB6inYsgkWXXKzwdJKf8vsXZKa/YXIrsQ+D
GDkdQZnFlkkUM03cI9qL9PVTLX0PSnbUY5NtoRn2rC4KNExdNAEpahbUOrW0E8uB
eLL1jVlPNFQzpdlBYlEv+Pw8KeOMcuRS2QSAgC3ycuo0cDHiITFmDR2tm14y48lm
b6vmvD3vt65UCssuhOwORU6nc9YmphaCoH7p6H92/OETZz51n7aLd4sjn6g8Xvzb
RH4XF9NIGIeRCMPvLNSLg0IX2G8beyuy/7+KIkUeYKyPbXE0aO/NrJnvh2GYaUjY
F57G5thjk+lKDyeKw+SBn2WxNVZbdXK2MqngzLgc4f7xiHCPqb7BST1TWHJ+Mmjx
1fto+XpXtFB5eXcx6ojhafFpAPr5HfGbaGoYIcHjMcjTmcfzfjZtKtKRSaFquX3O
wZN1upLTs8pS/867QXpPv1ecOhQY2xKC6w2VJxKciEPhfHu6NTYzx+VZz/CryHuz
uU6xIBwq9gRZz980MyRmRMIfZjI5mjP+hAobSK+5bN9JX5QmH+hFax9FjpYCzt/g
vDMOGYY9pR9Xw08rVrsXLp7q6nmi+FodM9tz+2MCj3QlqEBy+TVBVmPEJhbShRO2
ltwcRAYlfljX8kM9j4SQ5VkbfNTzP1qi+gDnEKrUA0iVpM2GthVABwY4HFZ0GkrV
nVLEqm/CYCH9WDAwQxWyMRpxJvTNqYOX5mS4oRfmFsl6z0Wz14J+0Kl2h6vKms6V
sO0oSfFULRstAWlHtC0kK7JmmsL4KUMbs9BnXBVn83aOUrfCHBZMDsOovkxFhN+f
tESbQrddxkkNYmKy2rBkDCzcOwmZwfKS/ljW9TX5oH7t3BYXnCWjgML8fHjx1HHH
Ff47jLk2H1U+jV18wNaFcmeCKq03m6XXtFy/P6krsv+jv37LwXlhrVRuvZkeunkS
wOuBHwn82c6kx0UxpDOsgs1vg41VukwTdmWarWDe7cdxvc4kUeOHAJ6MMYveHuuk
a1tQYN68+QS6gDthECPWU8jAw+P9lG+oKw2bEXHVoThyuk9bhCTap1lnF91fmkLO
xoOoQuxPzQpDnMEPZLxiFx/eZh1RnhTM2aiSy2LHnMkb2oT7NVparMq+QQUaTTWs
FvitTnRJsY6TpFjE/TD7HdbYmNA81HtFz/h1k+efPJ1/Aqzs1ynXW3BDWw1g11I/
4wON8ljrX0NlsPq9euYTeEceZu5QWxp3KzV4N+74H+k4JeXjAIxvuCuEpmHvZv+y
wz1Zgxf1z5VSKHUMxUJhBfi7dIWTUoDNTndTUm2J/N+DQOhjEhtDlLMjYBXgmasm
TqBvKHONSwuW5eAl/ZzldQ1aHnYJb7JiWYqvNfTCgKXhSLpjVxqsyTyfELW5mLUf
rasJWqcf7DEuKsMFmj6hOY1sLVJ6F8WkSIIm/T+0nNmAudwkxzacCqUlYIkAQ7PR
iO9eG3SxLlN03pfLg43gXgsUmDmHwB5m9hbXcjlsNBbPitoWSsn7/doKbJeyMpVz
mjkUThNL0y4KxHs5EyFaqfp2V5HCNIo8I7lDdKx6Ki7v82fGKWxZutcKTmZCk7BX
Ynom5Sja8s17//oLwBs+yJgjWOsCDZrSYzWtLvgln/Aa4r5VK6BWeM3uDclgnV7H
RMzgZOndlFUJaZmBvT4+lOdHI4SiMMWt4lzSKilux9ZoQSwsqOccEA6ZyzEe7RDP
k9ujR2AkCCSNVDFV4CafZ8U20XZCJeVcjeZJzauLywx7NSAukomKKtsycbZ9CLFP
m7dfD+Xq9HjdtZ3+r6gGTdsNeR+HwV1XpKodjlMD+rI4pVTYt6ujmNz8w6Xcvvhy
hv53kESAD8QY2yp6d9snK2eS6fLb4+02lhVbyOuL1yIN5m7/nNJob4dCYPvj3us/
7cD2OqwVbdHRIPd7N6BZSsEhhRl83m2A0w2dMbwfJy73ERVwJEpJ/Ed8Vmcjoymm
JCbGpSbFVSjTkbDKJZJcy7dkWZz0h6ZKgH5j0+o7NcYIasJUfgCLYicsA004hr2J
w9xjvz8ws8xrxR5tewiqk13yoZkQzJzozzKK8lTZFlbWL4hPVRWq3JyZT9Q3H4Wl
ld394jllT1iUgw3LfUr8fjXAj3SWBiR5c7wijpdS+vhpfjMxkMR80IMYSZJxe6fI
weEXmtTLnczhNNoJoaN0su2Qow8zCoGdoLGtjZ0X5AzGsQlGKTf/GpcwYx1tcZtR
noWNTJ9Ff3l7bIAy2AFhq+JE4CZPSkhA89ggJZmfQ1/61nrGMszpBA/51qTOU3m3
5o3Sz7PTbdlp/DPqCMw+o3V6nVCEyKLRtoRncKkgtobD+XW56PtCX12RSeEPVEjG
rr4sevi5IJac1YZTc3rXGHOs3FtgC3g+cHVVUA0Vz3QiENQ1iaEF67YWtEQt5kzw
hvran+dwsgs3wTaNq38PxDzGNWG8xndmSb+jXbXFeSGUd3Q+IJspX9/lnXJVu8oa
53wsf1GNDAY2RXtBjMrHl0ArxCgC5APQu1jH+iAe1ctLM2I+P1BwhEbbuvPAdb2C
Bya1NisUaph/E1lzLDoqAUhZdDBprIBmpi/qOBXnQUuJVgHnTycFtGVmBqdcopLz
E2mVGirqGn+FKb6EuojYKiXoxddmMl37zYNfPkyH0z9ux2iduoJVLSg0Kf2Tw0BL
aa+rOZWXtu3cvcK4SQQlW1xg1dKCzHprs8c7N6MRMCLNgwU7eme+AfNT+5zUE/8A
BvU3NvWVee8Xv0904Q8hke+cHzvXBCu6yFt4oDSyxgeHJfwl8h/6k8Ov/GJsKR+m
bqC5icTIJ/IsEI5cHtImXzalY0PmOFDyphU9VOZS8g1Tyf+rY0JjCArUZjh48n/l
m8kZ5onQVUqWtQQh1YY0zbiGG9WJ24d6MQCoworvxgWbbnNqai/Y2bv637Zlwa8H
7yinj9umBFrOF8cEuayNfxqjAf/VkyU1zm5ptHxpGLM601yBpe7JNlIyajRt28KV
sA5CA7V4Syh0lb+qZ3hkSF1bO4wi5woAP0PvwQuFCILaL4D9K1qa3etkd8qP39St
g3FCeAe5VnTQ2XrDlrdvoHAwBtz4gDO1jf3xVpb36+JVI32BiLzFqwhP8VE7SsKi
3qcozJIlQeid8dq5AKsLHvLEXc0JxP9THcETBZGo60NsP8b1dbou7Ap4Oekx2EVt
g/w5meDYiaj6hXBDmVXsLmeJDUrZPfhIW0AryaWPYXCanHphPNgxH8xQUjKCZ1gn
iiMmTvAYGKRZtzXOzzEz4/2/YVQt6k/psgLnTI+OfnaC0HU3yxJVn3HfHW1KqUQu
ZEC+cE6tpYjAUs6FE9ZucCbshApaOZkk8gKZNzoxO/uCYBehJgsZlwrpj5LwNMFU
pdt0P13Avbal81afHgMJQjkR49xbE8JjvAEPq0UWnWhiqkI8dH07KgxoeV+Jvipk
HgFOCtiYXFpAgyjb7034ooZPkiuMeCzQZeMaivMw7WfiISY6LGqxp/vtwE+0ZINS
U9qqLqXpxazrZGRgiU1O5GbT3kDhVRFs/HRlgfu2QEHYSIvHISrlIDR8kIWeXYwJ
Mzko66mgTAIUc5AqCKwcuSzBtNAfaWdD2idOAVK2YZiTbW3yzfAm7QfKJ5dTjmQI
3dJqUEs3HaOhX1FsbbovLAZSVM9PyaLsZcIblOnm/WKnBSd/b1p8lTzqY1WuCRFh
i1R3vKStgB8XjV6v34uiMdVkCvTFq9I0quwnh7gpfwaM5hhKz8jgQuzThDvzpwtI
Opf/O+25xVcLR+msLhJabm67Z4zfXKf5jzo3EjmV3OGkH2pswTQEYhdfE0BAXWLi
ys1u3DQvAhY9qsap2Gi4YeyF/5xhgn3W0uaeLSCuGOq7PNmap4u+9Sn0vg9g1GGe
IVqHEtX1gmAM/CmRCkfPOPyjzPvVrYbKRU2CJcJcrNxj4oh2cb0QqG7yDkfthieM
WaGzUu0aURtQ97vArwXg0XcCkOk1TUQymPVMG/ysIApAYfmh5BGQZyxeDpDf5WnW
hPEGOJsQRHz1vpDHxk8YGzvHXaOQUr9LN1YnaRJKCy+AXzwFSP73qhsXFRuyqWUj
/TuzyRgQrhoz5B79Ub9mIxd9Ytxz2ZZ0uLMY04+nsstFwfhzogEP27rPgqIc7l4y
DwR4H96jJmztxEjs8iwHncp96g72Vlw6dWoghNqe9AwqBju2jrGGlXkuP23MuZ42
FtIceSnJJdTxCbDGepAKkvKlwlrDONAQn6RtwmkSsC1A/B+reQP02e4u6pL0uw+O
zZfWAXZ+O+87AHoic/oMrVMyOXwPLCyS1bWEBBh6WgKaho6nffuq6X9rSn4y9fSn
db8MxOeEQXEGsLUieLnhzqXzC3NWDlTvuBaWbR482NONXM53LXsFs081qV7wgrFc
mgyxgu8zbhOIzFZFjpcPmUOIWNCIdZHOFjeb9tRlFkwH6kpjaV+HUyDp02ES9Uan
Z6yslEh9j7su8SHOJQrhkAeBGrMsipay6+JElclox1yHW4poIo3oU9TCiQR1rPV4
WImrF98fopWxxqMf7NnuZt+2X7PgkWqTiqRE+Gp1P0zk7LUN8Lha6lLMtCxv4LfB
vp2CJ4jwnGVLVZMwuqyMz3s97T9PrFSkdxb+g6RJwV4XVdWSa+CMIo3JeOFJy08F
Ho1YdqKoNCZuNFR/tUvUmIEMNqLCAWOsj4/LdZ9Dydl3yhqqmNS4DCwt9RL35cAh
yCxnuXEJaG25Lr9UP+t/UjJThOT7NErrdzxBxzefTIZhhVRL1/W5GAEice1d/r6o
o6sAXIbSxkatouaffOUya5gcP1uxG7L3sLcyzdtPb6i2Dp3wfI76liQrNPpJETBg
XZhmbeh8lU7g+6f+481DSoxQMlJiGsfuXnQ3mS/YtYqgqEz3JEKiGRuTe7RpBOf9
4w61c9rOkwaGc0I3Li3X6OkFQXKxipOk1/255J1WX3rHuPQoQQfEx/sqU4sy3v/A
ZPDPTuP+MmROwP5ISK3JfnUy8R3+Saw67TWUcSPQ+z4wQLn8oNK3ViTWn/N3/alR
9T1BvkM3ngYInZA3sSKDjOOWfe8+sWSPnw61sjegAMvLgyc7boe3a6l/y9bQrKNJ
JWyIjfVsgjhmAD7CWRbc3l96CnvTUpWo4/DMHMB7HahmMU8T5Eg1+3AZHh1khXVf
o7kk8nRVXpZHaZHrs15axY7EzY/PudupfD918ntj7HqfHXdVCYXkXgq4vEJ7iT1S
guHO8BBiLXxwi/ztEZW6Qk1QorTcnVPXdq35l/eUZZqCx0gtxcgL2pEg75CquK33
vbk9geCRu/R0GqbxUo3dFxf1Hx80njtmvNDMBeVGGNu4TQKjg2pLDeXc8FgjJIpE
xBkpwBdKmPu3XjpzLG/mlVucYW0K1Yhp8uElbICqmdzGoT+kViiUZdQoxEwF7vLi
mAjtfCOqklehzMnGiHcWrHjV2UpR/0zSja/SdBSCPVQjzO64395R4/GMqwi3l+jn
BZckH7zfJM7zDVwep35B9wkI+pqz0fgX7ycXPKDyKd6VHatWZKDxThZ4STMrPRZ1
mPQQSpo4r2t8/WTNngAHSKPAYCjR3MdKGZlCoPqbNf/xgIs5CajW55wM397BG5lm
YR9d4OpD8AKKTDiWqpK4iK9iXh3438ZFZEMyWN2GD5jLez3/wLt0bTKdmOCkWjeb
PSuDxhxg7fMOw5uC/LH1yZtww5Wd1SGspUw+7RrONadt51fa67YZyPqZleJSE0nb
UE55P/8eW25KW58wyqNCxdF/hsOOfGNL+fV+CXbN2ewzVPvqIjIxbGyy7sBP/5v7
9g0avGuHDU96ofeZ8b/1TaVzbh3BsN7VqtUbz8UTY7b9fnJdEMCpyxf/psRcFyC8
NnCNYYBK6K+gV3VGib0YeiYwGrH0j6rLn5zlKRHQWebAisjcnShJMkZn3Mwa7Ti/
68f24rdOBJP+07DQyaP/2kh7zEf/k3mh3qXSmZv1S94iMKsI8yLAZlMFmPAdDMRV
4l3EziOA8tcx5yWBYIkBp0VgKTgre2fQX3XBRVOHPp0zXqijX23N00f4cIz7pI3H
+DhNJbyMa8VfFn/IGsOVVZvOMct6wX0cPW/kwwPJnI/o7I8YoYikercxRuA41jUX
5z5Y1JTzB/nM4W15rA9YazBy1TsoFsxHkBuv0C+df8zXSye68pUXN/ljf1qW3+pw
4nXjRDuo7frf8/C27lCM2f8GZPfQWoPC0EvSFoPKRMEscpZJrsBa2yF4Nl8DM2CH
mDC+PN5p+JD7x2Ln+vENEOiofper4tChuhHxO4uiciGv9BTtYyvXi6Zc+2IdEnNS
0XDpC4lNl6L57vNqMXRIrG0jDUiiU8UuECQhY1itymwAUwxvPsBmLkxWHHJQS70X
fzyWIxYHp4uyZp8guRKW3E5SuVLcxP0g98nWodZ1zYQ9qyun1TcsqCp/AYSGjV0c
EfWbHtqIElk+T9P8WLRY+gL6NhAiPhgxzmbcCG9C5b8L6M56QRph9V/0aN2WkoU+
PostOfVvuRMFLWQdAhD3/NXIfuzA2Qrpr4mctwup47Vb0ooJVa6HwR9+x3g4A+re
XmvMBIZzgUdeUbLzVinYf6iHqYpq2TZagNO4RCXH+D0/t6PRN2uGn08rhtjJ1Wbn
MCuB446LdYaFhMsHTg8fj6E6wwTs5E0Fw7LkToewK/o68iXOuW9DCqDEZlBcRJlh
3foRChQef0+Hz8gVIbH7fK7zNBFN1TC/nvGfnzw4LDZkyeN6FVxAaEk7J2uBztJx
a2bUDeNO4039NX6u7wDSRBjAA5HYFVlnWByWfNnKBGUpFsLpEoXQ98+F4fQq1C28
8fN0Ezht9U+mh9p25aQK5mLyo+NBNj4uda1W1Sq2gGc0g2gGxBgS9SQJoUof3+OO
/j1tlqzhxuu4qP6u+CKnPKuGhvG1n4vz8mUT9pCm4coF5nscQI1l0Wxezk2SMcZr
o4SSu5qWNALSMbEKoQ8T/rUemxqfG0L4fpoBuF/PqSX6HsW8KL6Id/eaov6mXBux
12gUBan7sH4a5hXNKcwC/hP6Y0TiYNh16XvMBZQbUi+RVS+dXc151dSinVzaT5U8
hul+/IEX8t4DWhpKv1BIuLg6iye8TTrOwX9B85TkFbyfBM6ezt2Srun5sauFn4Zd
F5KrDd+SLwOWee3ZO4wYioEHog+5D7v8+jTFiOvVtArSlRcfitlj41s4p/SLOCMW
ogm/1WYuA6YyPDieFFtO8m6z9b5+bUP23GLz1i2gBXZHHFNFJxTE4qTmfjr8cvE8
P8IgbsTJLx9j14yiTqeN3RAh5PEKqIzEnRs56Wc3Y2XZQzC8Wh3CBUqyArjSXAqk
7K0f6qWjTEiNybJqV+DB4YxQTBCHeVlVDdKALcGF02TXhODe9gG56CHKEfQz87tM
YCYHROAmCwePT2dSZbwY11atZhDqPNRCZevM1w6gGx/01uJCXO/jtxytmfI6Gflj
VVk4fd5ejXXFjt2124HJwdUcaGs/abGaaPUVAEwh1nQQN1J/d1z9vwpubG6TLNyf
ofwiawwCCzLO09PuvssMRVrKIFdDT0G7VROUElNS4scp+sqIrD79x/SETvB5PFZ1
WzmY3bUb3cbVaYrK5GK2zWmp7MNGCBVRli3TS5hi6T8hgne3SdbSKkVP6WCnl+gV
RVPqiaVaB39HjHaSs2sIqRgyC9/aM6UUzUKvJ+hnNDJFS8HgyEWy/j867OkEoFuT
YeVFRbCkMSW8kG7TCipvJdO3jkI2f+IsVnmocSrevYcbq9qN5fOsj71vTFYx3mos
eZ1MTqHI7CqHxfH01kiLfbNnO/+E5KdiULFokTd+lBcLITgXt/pn5AbUhQGfLDak
D0IPZEzsT0a9zxL+NfP/SV+u9rr0E97AtfnlUsvtMt41L3bfZiXZ8UcigA2p3a68
Xw2/dPDN5Y9NGxsqLagLDF+jEB37TCATokJXCcps5yjSR+WBSZlc/e/z7xlLc3CF
2GbSLHbcS0A11K7adk8tIS64rNL98vyppFiTwbCTadhD9dQvMTxYDz9mppeNed0g
gyoysZAK/0UksTHrHwpg0UcCNpzeHi27F7t0VSVMmkFxD8jivo9lnB3LqyaZ/X7T
7jKJtd0Ui9nOOLfeW+wKscgeUtbwJJT4S2XNvPGhaxUQO3tZvIIQntAHZxQOs2mB
u2fkN+MFwmWYLbIvwoCgfkr6IgADDVjR9zlQCmVvO8j5MtqK22Gzyy/npxZ4lcD6
HbfHq8AlHTzV7LqrUUQZeZfXFhRn2sbqK0A8k+7FPAc8jRKLMFvvkftgmrhZPpQo
WdQTCGBpxWGhu1n8hnzkgEwF8Gztrlv0nssVGECtGL7G5pE3sA6BVuE6vKPi66Rb
pDjfo88yyqrBFXdGwaSagyn5dD/d8ekwBvyVUGOmsqT3XhUu3aaOOkMjRYlomeuM
Sc0Nv77BEMTGkOHTC7n+h4Y2h5dHd5AYjID1OA8/wwSCJubYEawVDfSHbLjdo6yr
OlDcp9trUWleyGUl6NYuqrX8FMtE4Z/v/TbHnBYv8ydLla7LFMjSLiMDub113k5h
TNt4BHDfqARi9mJP0/Xe3GwVEDj/6ymeOUJauCiG8YN9vc4tuYw0xOp/e0BBx9bS
1yZsgx4VeyvERYAt5iiersuT6f/Reef5byfjac6MsOJFv6EoP8ibfs6uC53MUR7f
VRxY0ADPKO2+fy46M9kJb2Bjs2qammq6+IwkLWk2L2JumISPGeqXVh2lAiVQPg2q
Q7kSl5BR9c/M86OkcoQOrmLxlIOrNxEn5KOPgjrERzMsid39zpA9KsXIUUq4afa4
HxxxIPrqOHz5rWW/OD1LH+Vv3i3ljSi1DpVGIEe4qkmNu2OeNbUkzLXtP1FmloWs
XD4w15CvT+Z5c6WbfGfGrpO8+RUfP084LkRAcn8osukQVFIW0HQMWDYUmwy14Is+
znRbw7XARNCk1O2Fkp2su3OITZy3pAfxzhBkzracwm4Wr5kPhj+7YUd5+a81fbAs
MG0HGnVUcNrNBryMmGRQ7QmOxSgWm2SXkSd1XRWJXh4YTJeMkoOyrf6fZUa5hVZ6
uUyWha6Gnx4rih89I8XTd2r6oCw8VMHxjSyByn1iimY3/uaJogWIOeg7dWVCDYGD
VUHqr2w05P+o35ZEewNAd6oYgFZ8Be7Wvql3gcj1b+59DmDFmoqJgm+UlusN+E8F
q42v4+tEwAMYucyM++uNIWbXqErDIOkah183M1Ps5Xl7QjV5P+MRYUIkC5NMwKhS
lHpjFNX0SG0na6uloZfLdIzQkkIxrculA916M/Ns5X2LbsFV4ayeozrYOiSy/ssl
s9hj9s1ni6IiMOdPFifY1FpMPv+/idRGPRnJyHWk3rRyNEikQMrD93l6FM52D7dp
Kedk9kCCzpruL5IoWkF9PsIO+AB+EiCyz7w82gAw1FZfT151Af0jwVmnNj2FeJLA
caRaHDerLbuDCt+YHVMCLZCCW0yryFPRwj13OGdq6biQnSBuExoY6VJfzwoOFZHO
APkwGQL8ocdDUGvwUWQ5Xi9+BpFq/iLD8pYwZGAJk8He8OUy/mMVfsfFD1Gy3j1m
H/wlb+ubldoOdoeRRBb9ye7Q4TkWH25Y6rhjoNIB0DjiGZqAbpXkyfBMx14MibKB
boU7cAt5r2No7GFv4PIsd364S5cLuWxv0jJzuBrQyKdbmZnsoltOhHwCyoJxqhz3
7v30go/NsQWOpokTI+EKLuiAiyF7TUQ0yxSbod1Km5yGfDEjHWZJflMNbn8+L5Fz
bde09fmoFU/hJR3p519Ri5FAv8zSMTtWKAuyQlMz/giUu+tTUY+9YVmGhUTVu+PH
cwx+DI4QZfbueMQk8eILiKGD2O6+erbfFbTbSVcUTXBGFyFnd4ojZ025CHwQOJDu
pN8zJrD9UHsDrv8MDDa6RKCmC7kWq7V/6VwxuUGkHQlruxM+bGoU/geYbmSMYuXB
dLQG+EUVLFU2XV7f05+6bmXPYudlOkOLTZEjHgnc81LAeMBNsO0IvQHyoDq2LLlQ
mS7Rs11Jaqd6tQ7MCBqKiGC3EgulEq8xOSWZvAU1Z+bYloWmtuq1QgdN9ufyGOB4
grHWuXud4eyNSbFNqkiMZ/w9uvmjwWVoD2kSQpkiJ8Pjic6wOfvMre9ZLZ//z2XQ
AqrzTWpLUgTvOOi5F19HobHocys+haBYoTQGoEBhO877B+2Gn5+4aVZmctV3y+1C
MQMmyH0Ks91KtvahVXl0R4T0NIRTYEPC9L3N3yi2WK2j0TjQMCune5nB7FW4SBmf
WV8HC2QZq1ekUN0ny9+MlJTf3tI10fGaIRuzHYV4sJ8G40lzcA08iFJrYLk17/wy
BmY99IWYZhSSxfuiNxaBT6d3+9DCF/vb0TfLqEacgd+Ylj1q6BtIk/EKrWiIcVGw
zFE8jLPyCxS4RMfkxd8F/eEJbzfjclXE3myWwSBqyVRZ/yl+bQPRVVH093w9/id4
gYoHZDWkwzQ52wDwgvdbe6hzZFCMbYLceauvpS94buzsZmIVzqyt/aqCYUf0AeNe
fpmVMkKos90qHe+Q8gu48eYv1Ezc5+U7L4R7yUHPqDd3FmLV0m1uI5q4CT8Jnmuo
CFRCTB/6DNLHtan1Otk15sMMyz6CddQdAJ//Yu6XKZBLZtqJiy04Z1a9MtcGRHf2
FAbfKjt2xH0HDn3oBb0jjXEvbC/siBKsYxRUYw/VtJgovuNwnFfU7wQVjtSZVNUg
nKQWvDs67aklqH5xHIQjxUyw367B//X731fuHoAuLPkY8WOn9cpCmuRE1P1Ay0eB
FO/oLISB9rtsWgz+Xv8yGDWMNJ4623SZ9PVHmaKE5JryLrQ81GWr2Ni4W3aBhNX4
2IEKZhvRVzhl19F3boS3F+5Ty55cPO0sKnbkl/sU/YTBeRoZ071MnJVH0D49fQlB
2cGxhQKyYroEw9g1o7CyzvLgCWFbRSEZIh41bz+ghESVT9J1xbb6U9Nsv5ZwNlF/
rkdeeWxODnvKQJIyj+WTn4xvcOZp5/ea0razXkQDzaXDIspzAJ3IKEKyPPCPDAzi
hYEqD5oQpHgZueuy45V/C/MXUQwmuiioRyKFL8X67Md30olfyWQQTQELgejV2dwX
FuNSe5K7ACmXuZ09BvpIDrAUJjDseRGjO2FdcXko1YZiTh67nr2pImOI/qAzT15S
utaC4ITY0Ab3Abi6SfzmFiGc2pu4O/BFuE7RcnTCVj/wwvsnkTq2htg3U9XbyFpT
vYrmOq9novXcjqJJVmOTo+2OpVMxyvKSmJk9EbXvT9Xw8YCFUUPHMvvePmGGFS+k
PYONSno04znp+AE0xW7HDWDeIOqbnm4suLjW70WHL79UDKSbAzOt48N38unq9d6m
8umfmZYJKl2sT2nzDtdOF/o4nnz+sWyL3rYROayUKgTgZ1817ItcHVIcmq+3Vc7W
fR7vPc9l3FB9nE9GoC2WEvmZq0X5245N0/N3SOVS61vDY0WhjlJuPK9Ef+qfuZyS
HNSizkgiWsH9GlwhBsDcds+BwFiaEKuQysPJ4Tc5jO0WW+DeHLM2x9tzYHkTPxWV
jRANKAFRBvEaOY8H05P8Tk9dLWuTgbzYd7aS5UEV5kD6h/z0J02f831qw21UqQ4L
dVl5B/nDwkZ9qo0LbXyCP3OwVWvimWvYcNb2LDOb1VnrvZNZLrIKrNPDy09Jg7Kl
Zt5vPPKSoB0pCkWt95Kk2CPS8KkPQfIP/mtKCBzgfXqnCTdfGsvQizphbH6eckoi
BdveaLl0rjTGvwezb4JtzDUXDTO6+tQgtw3HjQTUEnzpZO0ZLPl9RqoKElRH7fiL
ngyem8YLiUREEyHG2jPGsC70muxPNBhFlDamyA7S7WmbvChxQ01FyvaOWyUH56Ik
Cot0Yr9snxdiQkHRpM8903FhwxdDXKyILYrQmxkpo7MRq+py/mWwzBArIN+0R2NW
LFXmtwjqSswdt6bZf+6o1VsuCMr39z6f3x0+w4Ldmz5s9qiTad4ORCjvwjLsGfvQ
9DTtmyOHCbjlqywQysfz/ujMs6Pah0J66KfTFrNK6lwR8e+Dqu+z0kkRxKUYpd44
YvkUxpEq3YB0GUUgKV+cLH6kQjQE7PnPuVZVjfBQRODNzOzA3urMqvyV/Gm23mQ2
mh8SjQk/RQRgiFh4EBeiuo+zMHdsKk01T/0yhAJpNwCtz1jZ0dK0ncD8MGYpGgWC
vrQSe0ITU9cCT2QYgB5Ra89/Ynz1METxZAp8pDOLeGFc7oNl4rYZCUAsPqasNTaT
VKvz/tl91tx+3EIMptmYtLeFU0UfPeMDQe4UNvNoQfR6/ZqPXOw0sIblT/c1lkHu
qvj0WvSnqaHNvaOt8E4e1pLaCnF2kobN6dxO2D+WfKUm6mAb3QWj0vb1dwU7HVe7
1uggJHPYnjtzFSb23diSGJfbEixll4F+zAmM37qDYZNgWUv9Tf1ZmaoqZ9kga/m1
G/QZdTe01FtBS/wihlLhRszcA6aZEMG86ShczCZIC7V1V/mKAUxodIvtwgVi1gKu
5g2dy2DIP0HBMu+gjV9sBTEZg5+EMLAiAC8Jd/B4wYJhO6YXgxy1CHPOcA0hGrFs
VOm4OWQwJMtgo5MlSyHAZz2jVjwyPec9ZPUPkA6iBfKPzlxioEgDle4zLSAjyfxE
aEPnQvf8aVkZSa8vOIWUSjAa1p+JFNcHh4M//pX3ex/xhS8e268UG2xmCybAEy0L
m97EHFYtQ5DyPgFRjZGXfNrXSZQrg4skHcEmtNlBhmqjT72SXm7Cy4pis/CWUvb2
axkfXLoWzvylFSZtecgSCVNM2doO3HWCL5GVyOMWUmculAmOkrlVHdi3z2VZQbFy
cSMrYzvSbZKe5aTxbfgRX/fFctWpUzar7WYHyni7OvxV2IyQk39V0aQfa80IpDSP
/U1gz5o7CtHYIGKYVN/KGbBE2+7ryRKBGSEXzopVKEsFNzfL+ur/jU0dY5T/gbsI
Bqt8r/hICvchYEbBsljVTHQUO1K6cb2uePMaeYOz3t+/6NY5xLeXB3HmATJ4UyWa
+lvJ0Dwc8tGWHGhxlStl4Ji9VTG2d+rMwo+jEBXVXzQjTkAUj60qNMsNJg9K/OkH
jcURBAGd722ui6LEpCHgjMPDQfjCr5CPC9EYz3b8C+KSYl87tM3RsW4wgzP5ePMh
sY33y+G6G4zL37a5hM4KNAn7LHOe3l2y9w+tbfaHVdxETKA98Ge4+khaZZLJdKg4
imU2EPmtDYcJzzvGTBTgCStYLWo2o1dD4Ct2aE3ECr7Ua5jNBqLHIf7aNxgXjN5c
IercJzCvrtbma1vzNPVsVWe8j2HTQ77yHgqe+aTCvqfOllGfR3yBNcJ7B+zzrhBv
ObPPYLPGXPw+s+n67BwMEaXOk2zfoPwRvoVbORoVBWc7zCnZjCFn9nBcp6d/7PEt
MAhj5vsQEE3B1kg+wvBWQrjfhGQaoiN2qkp+M6K/6C1qF7nmmU6TzNkseCjC0jfY
EqUYddO+c7HeE6Wz0fj0AetrRT9t4eO+y/rvYTKPslYSnVtXTZwYyUrn35VR6437
dYpUFpnrhlqI0H/3cXuN+z06hXCsB7sgp2ZNqXyt0W7fvjSFKE5lpNSZRcUxYCBT
pTFTKe8UGb0j4YJKr4m1hZE8kIFt9oTM8kb38R6SFI0ZUDitVOFgi3XGE2iBIr8s
mjXMiGxz6aoBNfGPzCn3RD95Bg9Z+7BMeBwP8QWNipAF5iLs/RCrgEuO8mwxczr6
meNGg25T6cpudDqpJfATnEtO8w3IN1GWWqi1DQRYpZ81RdGVpF9FHQWfXnx6cbHH
YxopZ3RheYjWc8CFknaXit9Qrjfo1FTZBzD+wj5Ju7XKkzF1AnnkEm4ak0HXqjaa
AL6XAzwWwdrBPuf4p8axddNes0ZerD8SAQNGqed7v4aQzlaxhHaVumHZ9morGNlt
KVgHpllfpN2qNqGQ3C6WUBH9QL7ygMf6ggVvHF48+tyI89mvMPEDt1pEH1cEleE+
inKZq4hIBY27AWXoD+P/Uqa8idPOafSSwMcn3EnRrr0vbq+yY7jSsTiBXyiKEhfK
knKqzn5N1/Ur9v+9h6FiZErBOD+AOyJnbgbVVsGzntEfclt8FexFSpUrOY34Jyzm
fvmNIZT8SW+DzKA6bB50Ggr6x3qH4znpHf1oG6Io2KpoQKojTRvY1pRzF0grYGMS
MIPSUXTfSZwvUChJiFOr1P1IQg8CBcN86rAhS7BO5yWZJHK5r+IeTefhjsFz3T+9
djIKbvbsEYxMUL32GO6UO4i28PlUkKLbjItMw5UjNJ9VGNcyzm//1Ti6xAtMe1Yf
NWTCwIsWX/ftTFcjIPSxSpQa3g2XFGQxnvNBBl62Tmdm17hrf9Mg63UeUuMAnHru
AFVgLRAxvu05TSDn+KY1A7JCkU/ag/AFzjvf/rAsfTXxqcP3EG4YZlXrsVbus3vA
5INSt0utPmdfVzkN2b4h9NGerb16IoLQqqvSjt6Jpi+HU+HhVmp6ebIMBXGSp/AJ
2enVqs50EFaR/AKmLhAonUJgNE7bIyoodVcpWSkKlB12cS1+bn/0pmxIJkui9AOB
/KXxxLeB6hpApbIx1i7LVM+uGBKehA+CO70hcpn23/184QYc7TnvwH5Nt2Jw+VrO
7rvC+1XH08kxcEOjZQx4aAwOkrjZmAJUIfX3S6yI9+aKqiVAox4aONij8VaL/hr4
AiWb58Q1AxBH1qDzvgPgpxVi57YEsMbfwdHma/rLhm/cL6WZTdRuALni7dNU/V1D
H79xwDw132jXvcAF/Osnsq3DtdI419FO6Oz8ZfWM6lGdjNlTP+UAWiDCE7LBAWK2
7L5Cw/oQUTwdVogMzzzAwII+ax3bgyiuECiMZ3wVk3LqjpS2ocU36Dqc2XMGNCaA
Yy8XrvmagBu4NS2UFl6KK8zKp7rUWhJMvc8INP6M0VtpUUc4rE6hgPoVEzIoxMgY
jRMxxsRUxm/ZlqgnaUS6qPT7Wyv09gRg/8hJG155Lo/2AQFftejeHqtLQlphektd
sC+3+JbOewk1SoBkW2d6/NyLUuOnE4rXylBO/75gU8I0nsGPz/C6oi0zvSCWGiMX
1GUvOqhvcN7BpCsZxWsJYhT9K5yjPgA7AYuXqw9nyOmnVYQU5t8P4P9zd5p7CS7z
kTNU157LQsjAcdUyhG4JZ8j/gMIcLTUu1C/7sWxFss56hccQR3YCOh7ICjcPOtEe
jsD1zqRP0x+9Qdbyxoi92o0KmKWciyI1fv5qVpK8D+L2ix4GGBwiQRkAZDKQWCtR
Xjy3J79QtnKIwLBS1eW4CoHV6NIApGoqVL5BEWFIJx7Mo5Y1cJWUqJl2kgeK9ytd
PY2+dKfMJVVSHEx5QT3RLUVuc8Wae4DxPOFZ6hxIGDcUCgFe1/oyqCeoId6Hf3tJ
pc1XDO8ZFAp7wmDN2uy1c2GLDv1/dwWrAveAuQS+e9+8JCnGLFurUyuLr6eAwoWK
Y26tFprz97Qsm4FUrSJaytGaM/lHxWq+lNLUJwltlJ8AUOKkqP1ug8sVoymZn/Qg
ZMTH810bLNMSg1jnINDhJHbgDjKMd6IOL4KMsrqi6SqfhxI0iV5pPg1nqtSjdlCI
OcurDfS1Rxx26jNb7Ku6F1jMDD+gCD2SnFt8HfkmXPLK3WIN72JTe8ZFMNTfFx98
wIscGmYkTwsC8BcorVJIheKA1spQedsiDGKxTOvmkwioLPb7VeKArBjuGzLKfpx/
RmL7Pdl8lPHnlicv8xsxRx8aJqHgYKKVI9sJ9nAbljAfDuPE+/tWLfIElHp9O451
Igb/PZkqQoigbXx0OlKq+ZtJtD5BVgXFcNxAql17Nk8TfJFBUXAz/J4OgBKpPYY4
eo3CR3ciHGoUzvhiQEohyU6l8MSFq9azy3FrL8NalFhZKlH9Qrx5YDsWzmcWFb50
mQo2rLC8RwTZwDcRveW6JnxOzwLLTeQYMU6QjBHgQR09iZoFrgcDEdn52QftrPoK
CI+XF9XohqtbgrJiVLaWjd6VOTKt0Os6AFnXSdDYOD0LUsNC2Rmpl4m5XzGmVQhM
AdXpqYdVmYSIHyRuxlMKYiJFUqNxkKAfVm6qDKFYe6lIdsDOAJhYP9BJCCnkL1Iz
qb5tDYTeCqGCkDN11cfwwYVkALi0GwrgIINDo4RVfrc6Txcm5iKK+lKiSIhyQ9AJ
SuG9QK2qr6Mg/cCw038a1di1qjDA2yzvY5RQ+dv60oiHSY+hFNGoL7fhY9lPKt/0
zQYIsclgGNKw3H0tbK2a+diXvroPlTiLLgIp+UCIKuCMYr43tPlhT3ceWs+u7mIw
4Pna8c9PS0h6w0hMr8DSY4eFeii8dwkwp63XBxj/vh+t53ExfA7O+Xpisrcqx8AC
7E9O4ELOoX7iH+KwsLGwcQ7OXhmNrccVUeUXk85XTy12yzO3HVeSKsDCTaIV+3l8
SYEOXZTvMAmEcx/pF+RytysWD7CHMRQump0phtpfxDiqyf8Hg7bWSWBn4Y4+XWFK
gMJdiYnjjXf49xbsy74VwcaScOT/VtIGY/s9znE7HS7//aTP7RA8MdI+PcsuoNUP
YXVEr7GzhX2qC3ZKJqRO4qPsBCw5WAH3E9GCn7fTaF//ac+vtJGMGGDByhDLXc4G
f+zG5vhhmxGlVcYi6MRbJ6x+asKZF1O+6C5290McGshwc26JJ7YEC/vmlJ9me0U+
Bmd+KV4WcoMcfS1nRzXHMnH8CUP9EEmr5JR+bJBVEbM+x/sYPl1WHZpF6FEwS/r9
t9Tb2n44RUMdNLSofuwLuTuT9r47PkMa3kROsBYOgaajQb7jHbV4OPrVERBThpNB
TcKI8yvSDeBCX6P4BAYBPoNBgCgXRxzR+4mx4bGMvrqLYlAe60LyOWC2kYfEa+dw
Wf47gTKztJTB6DYJNA/s6jm5PQ/1/LB4Rc9jcrDQEKRkxb1yr/J1bbvmwN8yy6KO
Grwo1ZnMH/eHUrmvgltIB6Hv+A2Rl8XcO3AQ32oh0TwxL1lQo1hSZzEQfEp+Zln+
L9Gnkh2/nkwcvP58JruOIwDQnU5hW/j/0B+iKxIQ433IdsPCYW0kpFnBx3Q1WYKs
FFa54vShSVdpwR7xYmxRTSo2yzToIefqgIZK6g0AQnl4IaDHGGprri8Zj7ongdjC
07jcGT3ZolseITTtiAtdVASuk/WIVjPlBZuyx3saWx+NL0rc7u6MIiWY+2l3o2ia
EbSdKMmTYn59iee946tT1BnAeTj4Gloiouv/Tow0EYhO8tGfHSavGxS52274zZCd
Yzh0hqd7Eq/BsHtyRj2dqHAgdCZ59jOnH8wAJziU/S8dDv2qxEG5YI52sKU/8zxE
up1sKXqKr0cmD4jbke2JwKtzaozHk9N4hNkbfvPasBgPLAfOOOIRueEZFHUmfuoa
JugXKOwfWcrKWI6hlQGp5vBihCH3rWA7Wk/mgOV83x+dJRx3Y87BiRBeaS8ixKnu
L3nAbYRO0ygFa2xDQh+dfBXSkU2+ZaOe6746SSpa3MyCTi2BWLP1aZu3Adxv7tUw
WuOBe4j6gZbOhDNfq/S1YH0GCas8clEzBqMXaODINPTChmTXaCX8S0uAaZEdmQKV
3yVFG9Mc/RO4NmIEefaK5DVaWxH4NtiprwFaONu2zgBBuk3X4hKmBSAKYUqxRhWr
uI4YA7hb7QMBW/wqzXTD7poZtX6zUNziGLq+/ZlD8apfrywxmm28tJa7S1bfNbg8
qdeHFrs+VTf5lvGndZ02OKgSjr4x9UDymX7wDkJxNRrOMfbQRkiKBsQW2/ddtX5N
ID2I+WCOGNLi+HQiM4Jbj4nXnfn169mFDm9iVQCqXMNoIqkys1gIZhdSjPvebyoV
iuNSCqN3cQ4sqyI6ocRe0MWMAIY7oS+G18s8coE6M1MF/KlvkYSUqaR/1PIJGjVP
ke47XE+BZ/okM7E618eZ+G6TTQLGbCe57moy01YEq2KkpTXlLXtu4pMmT983GBB0
iCsvFrMknbw04FIBUPSZ7VYpFf1tfJ05EYg1YyyAe0NSsf+m++ILtJjC1lyXbsEv
g7KTXF0/SWYhRcNSadBgM9d9aXoQzfnPH0/BH8rZgL2HwzYYGfPLhHo968qKBolU
huHEWuEE5TGzOY833wwVd/NkRbGY9JSapoV6Dr0p6nAvncjMzduyA3PMnv+/yRdX
Lz+If5HgGQHu1h0kuBHGosa4/uhrej0YBVOjXPkfEZs6K0ke+fUx9RjUn1SvYYjM
FPIMlNCLBbcliWhRTpgdMRG6f5ozIzXcxmNBq0JtJjooPLDCkXqu4wl+wwlbde3E
Idq543prTBflvFuumPsvpQtd+tSN1z7KyB2JDCB51/iHaSGmQ3vk8/V5vAj1e2CQ
RuyTp3+9n7dWsp3lv0pGWTP0zGgQ4nUpD2dJhrEg4Fe6KYQq33PKrQr1S7BjSOcM
kHHVLC+eQJvGeJUgREfH3tZx6S4WvFgUGICT2O7kxSpzSgFMblWt9P5j+DJysPbN
RPL+XraXSfTqb+jaFyyPcsVY5IdAzLkjFeze5tNONBDJbZhlglZy5EBi2/eZDf9t
yqBu9Clu4MjUV1iNmdmxW6Mi5BjEarnF8E/PsNpFlTPAf2JJM9w5RX12PbtOjY8m
taI+ajCU1vd3AAbvxjK4R8VwUeNKQHAda9R+GNqSE7esExJytW7qnoX0oKJN2w87
ZGU+16m/qVGhzmIT6A4J0crrByK6zScCwufyuQUURc1OGc/e4H+i7jqjWxTA0rKH
4RBfGCy4CQ6CfCvE+MXGl0YMPy2IFcz0EmBbFhYPwRg9Bq7hRBaJbEcC+9AaDWes
6ZOdUKOmVsqBYO2u6f9BokkA1SpEJF3Vutg1YDtkguWT0HHYMSHuwfEIoNx+DsyV
QMUVBbgcV3TmGgaBtFhfs5m6W4F3R14Pr+JUxL6xXYZ90JOPHS9WxeQx6QerPBz6
HCZURVg4VgqFaE3byC1c2dgnRX79Z6MnSa5WG3utwX2eyKt7xQsnfnFrkwrYNJIj
TR/CUrkMQsYVa8xdDAZJB/R1U1qSYWe8NrNDMJgChiZmmxXAXp02ZcuUZgCL3vUa
4kLOW8PQ3jyanU/gFMw83upXE9rZXvIRDkx6OE2CClIu9BILK+w3y/ytelErRI1X
gZyCYlM5FgsweklN8g79eRYYUEqw/g54Su5xRxuisDXraxss12+rcgKfMyTbEA2j
L8BnrFelYaPADSjKjJXXekbQ1C8KwA0tWaVYz0z2GPldR7CFUDkGdebmMDfGdFr7
lAPk44VpyoDU25isH4Dq5U+AN+VIDCwoKmYojtFtpSsW1CVZPRMV8z1Dyu9p/1Sz
R8naWcnoaw0ZSI29DBCG74rZriDU7mbdjlfkgR/6ItwpyMdbHg6KLCdZCcVdHwZH
CfxkACrUxJ+ZiyyEnf9v0ZmFtLTMl+dUcBRNQwjy6KTumjHTJsw8de9ehRIZvfaO
A0Xhi8aXuVcjq8q9DCKvVdwpcsD9jdLrFI4eptmJx5KhUcTnDaWPdAhV+LsSrsjO
IP0p7clQARpeNr0NDe8XqR1Y/kcyQsnyU/7yCGTZ94fFrfO+iL/6TpFbps3BCTj4
Kugeuo+7p2LisqRz9p8JQmUx56z4LzxwZQBVda7/zkMd1dtz2cqQejXRHU6UVIEx
oPeYHODmdFo9fxKKtZWKNn4hwR6hIPT2IJmj1GfeLlN7sB8/wpgTR8td4RDrWkQe
E2UfRDORHDtJcyf4Uyxi03G29VNyEaC43FLZmsEMcoSw/zZvt56xs2k77blK66C9
Dmt5vl4YnZLe1SG561aEFeivVMUOooyFPxGOaBvaSf3zvafJcb+QnaIOs6VRrSEd
b4Pxxl1H22aSTgzyK+hkt0qwCEYVsrUyzf5SwZj593lqtuEejGJm0EOxzsENEkY0
ISP/A59+ECzUOn8c5qmddoDDJhxYN81aXz/YNQRBz+qlxtAn/wBWrak7AphqJHlr
akYhSQYJ21U21zJefGo3jPvKoDS+phP6GCJOkDZyyEXyMNlOvR04xWHDU+XwDaCF
60C2wG3IGbV+qo2AGJPZH15h0fXzSgJWGmGCkLiIa3qGjfjaSbUIO+J8BHS6CVxN
2yWY5N+fFlAtvVXDA+IyHfhTlDh3TOeO6NKudRXaVC+c2ry8iCh3u+Pr+/NQ47nA
foIcnSSzuPoIh4d7QGGnppDOua5cYMQnWEnVGfoeO9jYulcW3L1561JukPJFZqXC
pi+9Iy6dIQOcJCtmz5/m582xpTRguI+z2ZDQBDIpKS2hrO1EQHU5hgiKtEDKqtg7
eYFT66njgTFoabIWOmTygZ4OVpXoLiIr3boNH4fJmcBokbhAR6zSYzPvgPyGElPN
Bb/wNXRHCxbdhlpEAjyBgvtHg/6VBKvMRQpSfzYj+tJRlMqhu9RXK3LibpKKrZNt
Y2m1O8OIlwHXbc6eTlmB+xDfJ2zag8vDLDwqwscD5LhtLtANHtyQ3tkTbdPQXcPy
krCg9Zd9yMyVmhw+IGg6svbmp9QwywS+J6vDscTAqcgFUTojRJgjsRDQyLdVNt9q
KkzdayjH7bLT9GFOchv/bl1X2FEd4gdFwBFIJmfzGPXT9N0VScz9me84cA1E9MEj
Nr6NSzzUO104xwB6Hch9cEuhJSiffJoKm3E482F6UseVt/fyL/SjKOpFxNEs0Krb
gojEPH1nocc+boyoJ8R7qaxl9+7Lg5FUG3BLKRq/pXJjy19akY4jU3cZG5P25Jw5
HeQ8QrbSilwYnCbWJWIi6p7KKUqmuVzTjhfNlhtvSa2uwC1zTJ4SAxZ6fJIWTUYY
4PG9sLZvbqmBpkNO/QvRkBlPzOHd7P7qGgO4NDAq/CUJpB6raEZYyMi/KmrSNqa7
Hy49RF6NvsiEFe+jN2xYABGCwPY72xRaBad0tNsQEboHcuhtnGsdNfPB0iJx09VX
QhTpqEN5Mqzy/X8+Alpew2qk69/PneacfspDL4MOCm4iW+anXxZKxsEX9DBL+wEe
BRcZE/Bd7ncfPPPJ4tDqKrhixLWQy+kpJRQ2dn2YTPpyC3eqrRhKQpqtpkC2RUnN
82tNUU3GbRX7KnkWRoj5MyIU7K/tfrkMrXJ4GPQf/uOvly4+cGXH+R8PHVA95Neh
n4H/eAclwym78KKFLG9FPrhsaTNFJSz3v/2X/rpJDTXP3I5MeaHcvjJLy+GyRS5D
H7XfUk4pLfvRqV77l3J7MWA2A81T39/ODGWWBy3ykYAB7U1jEGEExFmc4JLz7b8G
DxCDcbYfkt3+g1IHtOs1hbVybbY6Sv2HeC/nr7lpAsajnPfdCyd0JtKLFIuqknZa
67cRyd9jYJAgjdufmhOROXdRQA50sXnqY0w8Qqj3ZsTH4fDblL2WBQCjQ80itNRY
k3bcWQtwUQYbBUKwiwkrCifE+Ff9GgL0njymvC8G54uyGzgOPBcmYpAb+T1tOmHz
zhkruktkPG/V4qs+aImIxjy41nOdPEE9jR/4eWkMyHGhPT4cVYwTOOpOLmY75Iqa
H8HPcMEdAR2zvDHHBLeALuKVUMiBzBPgbuL9mZDyhFWPhjkTknfZaa6y7O3qvNgT
0ELrpVovP207qohs4PJkj8f9sEejOeta7YYMF1hivb5IwpA907WW123j57RhuUP0
ED2SiBv3bi7pEQslOjbP/spBYp0KkPzRH3WgtC7xH7VEp6i6WPz+ew3ddKqHIphD
GDQ7PnP+qo/dfCEzyTl9Qmery+H0k/LzXTaSFqoBhz2iHxqE5kadPlDf7aJYDKHS
1rAR82htMW3TX3I0fcxjiCaVrdGZZpKSfLsw5FNveMutrCCYwE7gU20794a90Css
Tmt4hY9JJMI97QGZqfqpTPMg2S9fHNiaP/P/BvQc3JQ+PXX7lc+qTaQw4m+o4fs4
ayh1fwXhJAOhhyILOuC498mGLA1kTzyzjItvjU8guaqKZVGBRq5EtXnICs3BN6rt
WzYMuZFCLJM1D0cAau8ca6KVziwi2xD/hhSDh+LwtruSSaDfsHP7n0j3ky3BaxTT
khM671B6NiRabqql6jJyCizc1AvOS0f3MXbc9/k4eC28J3aZzzleqpWG5RmGEQwy
HXgDKcKcXrvE41T7o4dk2RbdKg2Ld0k6/ltiEpfNQA4xLie5LfIzY4R9nuZCqCyi
AzMbIuarUZ58Ywbyz5nJOKo7nuNZhmCUBZDXl+11Qzb6NlaRjcOYumyDXgV1umBL
xeVjpaiSN8DmAj2S/6dgAI/+z8iDPeeTGvqxsvvGwiowiW22twbRfRKN3TBuJFuY
siC0xqTY7hnQ01c89lz6fgSZNEGyhRHKCve1i6/Q69HOWwrF1XneqOS9fIX89rnn
OVkjRO/RbntZVSpxyGL6c6qVE/iKJikCwyOJO409uBSzf/tJDWCqpNpmL6c4c/M7
bEwF2L5paPqVEpNETj3J6iKvHTtKnV0+0Yi8HMfzh7o9GWZ+AtjXJPc4qP5ONVa0
YZc7ZBhSzDQnEtOg2LLqYhkx5GxfheHsULQwc6HCi4hfgABkLvCu6kc/qDkWD4m+
FB+h6UXpT5bXMN0gpdsaQUgjh+vrCDDVDdys8hFrO+IcugfwZtffZbcjOLUttMdV
cDzR5MhiqN7oCB7m031WAtLk9OVF4HFR3MM6VRyL+xWxOPqNQEuzCnGLenReR5YG
12odyrL4eiPACP0n70KcM/Hp2wPxv0n7I/exWtcaD9Z59dprzF1vSkFFns0QylLB
3igfhvFOV4oHrLqCTP9JDCLNhrWow+4kPVDYsW6N5rrhtsXKAY5yr+IGZyREnLLQ
ut2NpgrvJbWvg687P5COnH3P4rSLeyqjkHx7MyjCA4xRSKzKesiBItP0uwNLrhLh
so+aVsC7Om+j/OV/kRkrxUCK5qspUpRXzIB+9dyvL5o0ppXRGpazwBEwOYEHkgm1
hx39eaAHLsokv9Cu9i8SyXr059obm1I0TP4oLKYhjgY0qsqhwO4X/0LUHbHoxuBr
/10QhqVq3COvNGlWM9fXxSc5wtPVLEZkhHgiXQQ7TLoKskE0lsKhJPtW8GCjagV4
BfkDUc1hHX8EH4f53ZXVw9iU9bJE31fHUmkdELGI07bnBwxDGtOZZ0v+3StyGgZP
AecnDYugHuhVTZsb1Hg3Vl/nHwAD+S8s5uBl236IIg92v2BIm2X8cCKgutMX/GJq
Q1RND/44aKpTr+FWE/5gtinzKokwi3XWGtQn0pOE4glzVFwQNXMHpd1dJC60DSgQ
FND9VPS9qQCvI9kv3jXc0CHc4BNMuBfoFqCQSYIn9WW0+kjyUVbhaxzjeXLTOZg+
YfQnXZZP7fyewTwuZ5JXfiVpfVRuITaAFD1uqJaMsNdAO4zs+dwOObNC7eVb9xFh
RhJnxl7Vg5T/5uGqGUTwWHftCjVBAfIRYScHbB9oeZp361bLrewYZPrIlxGf5G+V
UOz0pnkNiFOO6S5AbH7TwnpNcg36ZL07KmO2FiU1w07zLyX28NsZFSlEaBgoZk+2
m7A0BkfSUGzFBVO1jQRAS/ta1xXWTdcz6W0fXXXqCiWEA8J5lcGGfRD6FrKJYbhm
spRRpzYxbfEPVcao+fd+AZjwFhc8HFXe0WX3oQCQtQXqpOXeHJMz6Q1tx6wpG4cC
/RgRLmh+WmnYoSwW8FYMlK6ZPP+kRM/kz1VT7aaqmVM7dXt1YGGTIvJ5HseFeYkv
53BVdpPxGXh7nzal14lOgZedFw47myr/dOQMRSDIAqO9D4vnvX751w6+JDjs9FJC
nhwQWX28P3yE+L6kNQgaod9OVTNkmOT3ccha3vI4EccqCFlXmSQ/2nooGCfDvLdu
GTkpX7GCTUKmmTk9oqA/IRdDe0EPlWDa+xzLMVY/pDI5CParEV8Fj6ARhjCQXPYf
xY3KWuEAlFAqbi2jp7Z6O6xGMRxwwzZ9kujdpBPgfsc7x/9Ul9PPa5GR0gFF7D2v
N3H8AEe8XNEAtUA/DZST1gyX/J3UPDqvE6vRKdS+XOFARuvS0w6VO2jJPpDbPcWZ
rFPw8YSFQ8cxcUBedxDsceA8vmR4ykRG2bvpzv6wPbqGwij5bbJaoMuqdfz21A/W
4vD70HNvz92NI8RdX5Cz7HMrT4/f2cFPkaG6QJ8f/XimWcNOfGohzswayWTWNwdk
HdYAonsv103+swF5c0o/BghXZQX4i+3sjhYywygPUMPzWBC7Aza91Bsagqw6Sv6/
osqFb5rtgCQEWC+HhvhHHGVWG0bxNAhkhAAMuMPCyQ2cflZc2WnWlCMPmJEYrSVN
3liCgR25Y+M3HEFo7lJPzDRvThNH0z5bui5EHkFoKDwqpATJkMpOejMtUl5/6abf
2iYWVq3nCIsNwBHuVknm7x2JfkBI2lZOu6+aR4r45UWyfoUHgHPproK4XpzHyWsc
zSDfb3wzthXxQDKjssBI/jA31gIPoN+q5bYqmB27al3fH3dhNgePdIcZ6ZYuk0ob
yivVK78wrEFoGjq2OuJNQWHBvTQKU21kcr2cOOuAOQt4m/9LtnfCIje1U9uBnxD4
M0rg9Obn8KAelAlR3N6tyZYDJ1JT8xTh+pRHqpKG3GPxkoG78VrfKI7XOJydF/IB
Kf2o62hzyfiTL7SRAgAczZmXkGpqiXfS615Bd7C3O1kJLgr+UMfHBp3s4nCjsxeL
TSnI7PtWondeFoaXuQof4VLWjr3TakO956GiwZSrCBGH+wZAerrXUacne7RSBDWT
8r7o9mILdeKinfKqyn/dggobgnfOvFW0PdJ/0QESLsfp++GN56Y3VfC6d87W0OO7
O6oyidO2JxCR7aol5HzYclrcl3Q1rPzXyGnaCUl3xS5TSVIf1jsGLiUYjwXQ+z/w
BN86Gw4f06I2vjIoXMuauepR152kIbpoKP3niSPsgzkoxuJbR6wjbmiq9OZ0VG89
4nZ0y0u7mlMlITzBE8eQIJVbIRh9bRwAyYYC7pbIF6vaILZ+w9oKbXLNicU48UUA
NLfj0FlM2Ws1DWQ2TOt+Q39w+y9jgJZ5lQ/NIt7cuQKPJr/mx/QDDcLU4QXGHNyH
6wwEjYwtCW6ixhy71ixn5nlfXZP+9J7X8aBi5+R6IKHlJskEzpaUykt0lneq0mkq
/WN/FxIOaB1yUGwjxEgx2TRd3mLhCqbjxJf4aJFs2nTrRHnOyRiVK4KBKLXiTH+k
guV4rIhEDo7SZpiEczLmX2cxnHObdreatOIRB84b/LdqYz7WCxTTHI6n9nr0he0v
RhSU3UdLYIstEpjgOLVDHVpDYj9w5loY0FN9tSCHgfkNAvv/Kmu+evB7t9J5gOuI
jE/o/Ah4NTmLI/g/elw4tCEWXUVa1TqongrRj3GWhL+2ntLOmHQ1BX590CcItDVT
p6Cism3n8kx3CCwYuhlhbttJneBxgpN0tQhvlwwalu+SYkvmJ9tG8mgRRKGp/4/y
nJ5cPWnfKEkgTxe+72uID1srYNbVLRQbkzbzR+sxMbqd1KCMf2/qDkUEGXLoi+NZ
Ldqet3OgOCY8rsiydmIgPS6mWaiAg0a8v6OwrfImr7rxywvdo38vnDQt1QxoQZlY
cYndzQaFIYNP8aJMj5QYMCDMuaEP+MTda5WBJtOk2ZUx/4JgLHxgUtMhVIvVBnlj
U0+5Yi15DP3GX9LAXPhg6n5ucsheJ014w12txkLFhLKuTR0+Buu5bEkTUTvrzyMW
LlIRuCMSDQgyuUHFddxkwjmBEPjFESWpL0icdkJUksU3OKZvLlgbViG1NLLaxVwf
+vIbseBdte8CTBkDobl/Otoyfbpu6S14FD8P6CwsIFbSUwAODYwm6Mt3anbKaorI
Mk4WvgjYRHAFjXAp1PXPK/pyQgTsjJnpxJ28O9o41q+DnE7822ylzkGTO4eh5Ri6
oQ21KmvKA0PJlZsIt+s+b679ETht6w4DPKZIjl9uPvxgU3wm7dmjShGb6uXGtOja
6Ia3IfMhHuak3WVtt06hEp/cZNIg4kRLSL6tvxdx89WUNwK0dN0rj1rWY0KaW4Jk
i8Mm0uT6HreAdyUzzCbzcWv2JTmTS14hl3YphaJskvH3p+baugcLB3dfFUduZrGM
BnnDmQ4lquVsvHgMeLWowJOEWWaBHTPW3L5NmNNksmpTZVCtXcgAZGIT73GaYUnz
qdN+N8YcfOlYBJsTkZ1WN3QVSgQWd0ZJNPKK3PZCxlH4kQ/oyOFqrNINMPutLZUS
5mSgNek9pfsstcqsdT3tzKupy25vKOc2RF6C62prILR99CWgZCGuPC1wej563DW4
81pV5T4wQ/eegbxMYRSfddgdKDyHA8ZVvsqIzob72NROCKzlcqxfJPFvrSGpw8bD
Of83I9+s2eg8uIB6bMKykXFi9Zx2D3tn7hmIuFfpDOnzvsMxU9q4Y4tnQ4o92/mS
kn54YouoCB7dZD9piKuBS7ebzXYipPUm8zABOzWnN141vFy5CAWBFsjt4/akBRI0
JhXswTT45ZlN3zaQsskdrnh53GVkaEned3z+igzv4pHMSP1CzH/pHL+vBElA4nzC
cIxO/OInWx1WCzGcOuIc9YErO/rzMXiYaR3b4KSqJ9arR7NfxdyyODx6crH4a3bd
SvUcxaUpVGgerBEXrmemTqCE+SdaLZd2Q0vY/mx0/9mLCt6vR9UmIqzFZJl/V/bx
uXCPrD9QJfXgoqcrvBwIARJ5secFagshe6xT1G98ltJf7hi2OKGgdf/iSdixD3Qh
ZFoOhSOoldrcZxKPqB1/xvsr71zOWz5OV6zWF2wZ8yqt2G1GLvU6ndiFfxWXLJ4C
BX7xH7U21l8FYu1S3TFQ2l9u00Cftv8mpLjksW3IRz2DQvsBBb+xESyIOdFBN2yk
6N+HwaV2OXRQagRxFdfIvbIuQx+0MrKF6sxlzakPFQHTyxZqKwgxB6jR2rLmKVAV
vsXnFYRVLf/UmQaxQ13l6y+e3TPIBrZ7wIgmpiJJp4Sm0jfrT6zuIfaz7uGcQ1A6
dDOogXznq1NhHklNT96yDS9WUXdqXs2FmJeS+MgKGpY3E6qTAB/jb9uw1t+fa2xk
YR96ariPN14O3t9sv5FfUJxPlF0Dt6P+1ZojSp5pQm9DcQkyDLVyyv+bAcE9cSXU
6CfLX2JlsINEkO6S1JRi9MOfCXLhzOxMrt5YY9v6AYvFUl9DBN7/14eHB5zRqSeV
0V6vGPpENjqT2D+f7V9lzhIk8YW5jkuHl5cQjReN+CvQKuroicV/ts+hiYA7S/DK
7JHO8zSkgT1C3t0W7XEIX4KQQhUwECuMOUH+P96LjuWjCfISIA/ePeOlj5uc5O17
saKZfHGo5z70bvHYWzTJhMiBcT6pdaqhnboIbRsIttmCc/ZzXN93I3CJUHNNqv4o
EeAnG3yHaM26pTnVqNK39PDiJsaXtd+mJZT6AA31uM9NQeGqh5LrFVEnjDmRa0p8
Pw14qfzb0AAtdxghV8iqLSDAbYlVsIhvxP0H0wMbypSiTDR7HUYK819cYrlw+LsR
/p8vioZ06qCbvW2tcRNzHzD0MFFef9zJOtmSlk3lwyyoepEjd+n041EylfLEqNPe
HGnMTUvABleEKXAO/awcD9Ru8UunjVfgGN0Cr+x0/v+U0Wm+3YFeY2PuNUCL+L6x
cyEop616NOcnFJO66ua2maPfp+w14DKqtWuo+L9D2usZkkrJrwkQAjrxsWDQ5BXs
wJ/bkk7gVLR0N5UL/aWyksZWrByB5FjewFp/XFcEE9FDv/M158e6lqJ/1w8s8JFd
5q9R6hQZAqK7hbZRIK+BTuZ0UCkRDWdAeiIA8NhAxL29+tR+ZpJqpma9bUEpqTcm
/hF9gBZNaBVQvwX3Zbq5tFBP57DeW8OmAP9RrcZXKP/mhqLD5Ikysuxkz/WtGqAL
8yku/mub733Ov/5MiNc2Dr0nJVfzkkG3wLwvqTq9NJhDUmf+kWmHomyZUxmaLj8c
tfGa6rDvN8SluS3pm07CHy/PYhBONgiNCJO19tgpUnls2KAViodlrsWKy9bl7eIh
9V5Dth5UywI0b5jFbtV416asMfN8PMeVinuoLCABHMowrsGNiP3ysfGhE/Ue4ANJ
ROVQhGdAU+ZUTdvL01h5e4v6SXahqMVwavtnZK1IZeTGh06OQrufbpsHD/LHbtSL
8iJhDfBd/6smAqd7aP8ci4lhmMAeBj0kFN9tRvpYTmz82n3EpnOL2BWpNVkgqfP2
Fr18s8yP2T0yA4Bf9RiXdacs57N3/7QGbI5phMyd6vJrTs1Lrx+ySha5Cv0kgRFi
0Ux0egciyosz8WcR7SCGNG5tCbnAUjoLt/LayhB/2M6LI27d9DtFFrc13Srg4jJK
cDpPj8uOGL6SWF4JUEAtsx9Q/k1949K8OahedXE45M2GH+w0P/0H7Un7ykcsGnjC
E/RJ9nXKIAOYPXPrqNcpfKb8c8JLxz+7tBiGkP3lmsWNGAbuYdT//4m+It8GcB3c
jY5grnkI2AQ70Xp06bYyRIyLFX23XJ/CXFXGdok6Rw7UBYnRWWYUglAq0jHfIN2K
cEEDrVsIePcKhFtx/76EKZcf8I2eQPcj9yvbZZUqjDdYXOvvuXPVkmQs/X7KXikJ
i96Q96EHAV9N7fWFh8iRz7Z1IarX1F8N0ozCfFI6CHoYLznzEyvnYZ+iU2xuvPw9
SOTIdgEDwo8sJpN5nzZ/FgSG+XJQ9vs2YeBXg95BAwRcmJygzFCVxlUN5qe3oHo7
zRjAWbVTEzAhwqtaydtYW6e8iYNQf9xRF+aFAkA3vNFIvLkp4BcHrR/DUUcZVzid
kjMIUWqTPWJMOm7OPgwjBjlp6jB0jqLilCk9IHsFGqHgQOgMJWqKk5e4CtjYXoY6
M07eguNRJxFGGc4j7IsC5s/x37ODA00k0LiQkXjnhoo+xd992dB/OY1RibCINAH8
+KWD/agY54Mc7kqRXzDAmH5TVEKu2kXqeTrS8sJBICi42v/0ZOQaFo7J0HJ9ctlw
APo7sgyUAAuSVGbsJMnbFV44ilDABVq8akOA8HTKZKX1CnjtDMOG1hfk2R1Cm3jJ
AQS6ebjjmrtJ8iIT6/LntnvL0+rkSUza/uXRhXtdm/hzPkGCcIBEonSea6gmjA0z
+gkqNTxl9gaU+WgYepR5YowYAEmvt3k77k4BtHbmPTOycvBMrE0vwQrS5CjWWHGm
x8So510QOyE68Zsm8sbBOssQTlT+j3RhOQpGgTOvLbDnfarX0qaCT6E7QXeNqfib
lyfaBe/8QaYbXvvIhfAof7q7DtItEkKMyD3nmWjiRDEguyc3VLTOXe0wCHldHHzh
uYx5+gjCXdsuioeVD5WJkV1h8U0ccnYHzB4aPq3RfXVHf+bAsMf4feOrQEI8fGfM
s8YOvWRl/969QGQr2JotAMqY/ukIC8xTQcLzZArvg/DDpymOJKb4OsX8FIrbsK58
eNgSq1Fz5+LRI+lEkzh3Ul8cDSABe69ACyHMhlsmY79RFSn8RXKRoGzW5a89JIeO
E1J9b2Ju/y64Cj/xA7X9Ow6WrtvAGi0I7DiYeXoRl+gI6TgJ8hF4xhEWA2q2AceN
ekBi/i+JCfIrhVedJsKGmolNET5LAivCr8pJf3ANI+XoPw1gw6j/oJUUAj20M2MK
TH+jWM5xM60MGqk6U5HGaGonIoHCJ5ZfPw5zdBGhFyZT3rUgbvJ7MKrCX6LIU5uo
OIONEubm5HjqPpiOvcXcAm1uzbHvazYJYpoAolpRIwzLtoMRpVgtE8vKrY1f4SEg
zHQkFd1l/uUO8g8IZiJwPBQUGjTD3f5tQEvDobhuxPcnsJEWAw3keM1GSfFEdnJp
vj80fSJcbVe7FBPuNEFzmw8uqB7f6wnBhM1dzdj/TvzWk40muPqBtMw3ODKhTpIf
7TKE0vwgLNhrWLPKV7fKy8H2wIVavC+ZsytuT3c6lAYqepq3J+X1WlaPtzyJpkT0
SCvKxw9hblaZZlHO7DRXQ3CtBJ13itjZBfwWktqEpcGeaTBzYz0do86/RWGT0NrY
yxnFK3KDTgAmu7vDWAEd3XWF8Dcf0zGyuOxs6PEO5sfictaDhdmcADZzM0vw1stb
uQsuZRFrpLdDbUibFyCLVLjwHM4OzHnzWiNir2ztby7bSe/Z/2R5aOQPkEo8vMyc
yxWCJic4aJRuWzepscZfdRU0Ef+VgGR6TpnvDbnEX4buwdWcikVrAJCjpOUiRWT0
jnDjRNOiwtKrMoF3UqNpNvwc+OqAedqYF7BTiyCNbd/1869AA98mdtH1T6MkTPpV
HN+V2Y4BXShTsrgDEZWJCmQE0r1L3vAc+FFYZCtwQrSaEGKl0rzfRb7d6C8NN8ZT
6lZ5f7MuXTzQs5nfaaBpia5trbO7yTBfNInqePR7wKmKRavEcJdqHaakIcWrcDBO
vkEOCf9tU4xpbN9CWkF3sGuWQYl4HSHnxD7aYedh/Ruo7nLD6Lpo2SlMyIEINd3M
v0qcJt0YGzpA9OiqzYR3V/Jc6g3cMDMZ/Mt2+TRn2gN16EDfbufia5V29dmmviQt
G2fQ9xIx8CMvFqR640Pqn7ZNB19Gw6VG4WmhAYTUkvRfyHG+QO4lfAtIEs0CyIU0
y6b8ogMsdt/xkKBa1OnDcJo+2fLQtFILtRQBK/oIVcWSfJob4GmyPQ3GyYbMd4u3
qZ3PhdtpfG73vShQ68GSeAogrA+bu9sut2mD6NrEdn/2a3mt2yAYAxD2c+HL6idE
6YUJI9wSCV00iT8BRNEkZVKx747QwpkjbunhEttRn/BL8eros5YJIGkhq3uHpmOY
hxXAt7mHuPEifPLYEsm4EX5KKqa/8gQ/7h1HyPX2tGb8rpOWPMRdvRagcESUJwlQ
LLdDP5DRxKcTpIHWUmH9DVmWzPTZJMBouDDR8WDjkCp+kuYL5Tw3ua+QugcT7ACR
oUjXG6BWIqFdXn/GPkRhpnvQU07NbNASuklkxDKQAeUnwfVePlHeZNe3LpQ6pkoV
fRN4YV27xxOPafthhbbOHEI6bxyKOpYsKCtIIB/0Apg4kqzLTFb9mzDuZRDAQphy
MbY0uc6i6kQNC52/gV75fxuFpTzGX2niMr+qZwCvrErYtrbiP4DtKDlkziXd0+lS
qJMXFbI0pF/mWVmQLcKmsL6LyqC/UPWoxYQiyTPUT3RPaN4kgzX+WlFY++rx9fQX
kdUPBim0ModGQs4rNzE5IoHe8/9tObhHXu3L0Uhql5eXxuhy+MYDwtI9Aq+Buwqr
jdEWaOgfu1QlMIKdQ5T+fRw55yY77ikZ23Fw7L41cC666Y4YWd7zxJYrw+R+gZkl
pcVILUj+4tu7L7cIiaBR+xJ9SLsdLLe/eXfvKO+rqOAuv7AfPbmBYla6A9wdit8j
BCq6oaqa8y7U3AmvbeUtg8t8VB9P8H3v5BhGvt2+WUJdl/3Nqq/+A/BKihAwtLgY
4AhHklBbhZix7WNtJOvSYKbVKZxFJa/Glo/9WKwQQ5ZDPpssH4YM4daPJIppYzi9
zSfIXHCw0Sr/RL7BmrpmHf5/kjVwx4Y8Ec9yeHErLekMA0kiE2l50EDYcXO+rcxf
ureo8JX6jmm3aJddkVWAtjixhVikgKcb7jMIvRJFOn92yzfJhPPJ636qTJlgomhS
ou5JQrNBiE5fU8mi1TRyO8q8QIjs2WKTcX83oakqeQMykDRWcdi+cYgOvywjp5wc
325+ilOx7a8ovCZV/Gt+oAka8zMCZJ9R0sqxsDWPQaubqkhuUdcRzBitpUKq4x79
BuVbeqeDk0zdEJyqOZ5PvbrYJGGdjECcHo18Vj39JLP0BM3/Xw0dgsj+eWJutUZR
QQen/qV5tv5Cr2kHYL2A/psWMo+zvYFPk7t0mFC9YKYwQZdV2sfGV2Pa1LautkZV
0xd6RfhUrvYt+LnfJwVXsFM1fo0CaK1JbA5UkEqhQEf0IQxKGp51bgCnzjKDwWnk
9xwUaE3EHi9Jsfs3Zy0477E/nBpDluArpdCmrLl/YwdUwOVTj5qJj3nzwcmugxeF
7yl5pUJQBA2TB1fGCcoknkSmGLwPXsi2fuITLv07j7iegwKN4yTBpHiUFGyZ4hvx
U5PIxlViG9W1cNeKLvt+Mr0J6oM2f+GY2jKayj9pCEpKGA1xl6S2nSur8Q+N5Ila
AterAiErYKPZa/g/2AkESEShpPp2UvfsCkHgo+AFl7S/on1hgsANM9HGfG17p3eW
3VfHKYC7AE/KLmXljPvBPLPHYgYLw3M760pdAUWwhR3F2uFTazrWem2I6QtMHpjr
ASifXhWnEyXK/3JROn/nwbD9qG4EwupUBzjD6h8MSqDjMSbZ5ZyemHZMsyFtQ180
5fIXfZ8NDaL8aUgasavkBQhy3Fb6l3l4ZInade5LkpglgTy/4lrB0izEnCBL+f/f
auvqqQGK3hC8GD8AvJGj4i4LsAQP2BmBwgZoFLS1zC84bFodsWTIHjKhn5Gsc2zS
t4wFIe7xdKA0zHk7vH0AB0IsE4PKc+QgsBrQWHY958dwzvosqUNB8sPBUdlsD5IV
cjDydZ8FxJ5LvSvflh6tpRJq0J3xyP4RMJVpZxVBOaqfouEDm8cObMVeLvGkjQz2
QZAarLYSdKfRfEjhIKn2FtxpkeLVCgBPC8tBMXG43USLIR6o65Y8N1Hk5c9J/cmn
Ue+g5KERWthwZVdZBbHOnPbLL2gvIGirDDuInV4yRoZFeT6yDq3MYnRN3ALeED4e
e3upmNLkpJErK5lcY1Opxlqga7vqXyLs6CgmbOwASy18pk81uA2Ovj24IQacvkuQ
fTZgBGhIeSbrEEpqIqf3gsii/0+FmRmnOnSFZkZmgMglnhSiUGO5gUCDCpKcGAJn
QuhtGdkX3X+5hsgKYcze1bwE1D6SkwTAjHYyO3H+63KBuB9G+ukycbekThBWr+u8
QV9iR96RsUs1E4TDhob+2TFtQMwl6UAb48qx4WDNi47re7Hd87l31NH3Plk7HTZy
b1c7u9je3+naED7fAv9p8ziMhvBt/iDU2qd7BuTabUj9/bippGolBtJ1bu06Eh0I
BmLnqKxSWFReC1/ipGeO2LjcXnDtAiAuKAABlssJBk/y31+JQAk2nAZoPjGgAC5/
m2Rgc5FlCFQ3LfZkiQbDZbQ48Me48hw1RI55Xag03FVxh41UlINfl5HumT0sOfEh
xSV5/ciMQLlfFxqgoiYMQDelg3iL5L4uaV7OysoPp3lhSi+pst53ySc7rT1diG2c
GL5NPFr57KMKlHkhcE08H7r0nLa8kUTm7DxENqw2TK4w2p4EnN2eIFEekdPTsNn2
jAKSAJyEsoCLxhXB44h2OlWGo3sI6/62FT0F0F/zDW1feJcry0ay4UxvsIDuwewd
hdcd7MCBjhg5xaOJQc3ua6hIjrCahWB/yiGOYytby0sN7cyxzclH5MokfjjTghFm
UpAABPc/scnnXGDLfOSES/izcmgp9UnoweD5fqNqQO/uE+9HlNl3iEd8zshh72YT
OPJtgUNwJMN/jh5MujG03deAqPni6nH0FycM2EAuo2Ch4fCU7Msd/YkaakeTZYSV
wjj0fYJ3e2om9h1pnaq/NsUenFWirTg0/uZs2JvsrnlYUTtreFybjMcp0HRFw6I9
O1hG6Rj7CTxhBLkMHqUmoYUA1RmyXIkkKFCwHXyjn4FW6BDtWqLFNuwUjrPojsPm
/8/FyiPQ8ynAlxKIpJt2+w3k3ZtJHoXTZuP5tnml+DmLGZHfWFnjDW+N7H441tUa
ODVidhw8INXwzQM+6bQjwCMY/IjYM0pt5+i6W9RK68Yvdsdc6DoaPtNIeRJR1j4W
zWQ24LmmwUnoLIXVsiijUzxROklYZUNt7lhYSD8M1fyc50URS3pGm4yDLHCniRhm
fd9PRqfv/Mb9FKjcD/xPzuSuSq77m4g/+xMh0lTBjW7We9M8RTex8IhreT3fH09d
5ZIX0dzYPIm/VJ0NEiC4fQsjZklRyBTianM2uc1sOR5mCiZP/arHwedizXktQoxF
/ZeZijxgft9lC5mH0K/GOas3yW5yZR5znueS0kO5RIFnybiFzCxaRuOtPQaxCrTZ
LmoTxEabkqclLpUgZvnRhAYKSBfXSW0kZKT411hmtJUlPQehPQkQ0QgOAjoJVIZ4
Q2+kpDH5FpO8RfL7q+JwVmnXi7dQA7VVTvd3Y7ftbWFVx0ny6nOJJ27vZ9aHNMYK
BkCeeR+MsEUDqH9g1miqmnyNvyP7fgg6cH2PVaQDZow3chXfbErJC+scDT0CWKLQ
dfwzGyq6TUFcqYP4XGWRjXrPtEQQvArwKgCykfnDMrtMb1sIKKnOcdb3qUqOBJ61
iAjc04swgoaTxmkRHZSdqt1T50yonHofUs61qFgIRaF5s6QZHWhCPxD+/B/OD0iC
ifpa0Aw0Si5Rs0/+jAysocISUH34X+1wZIuytIIB+uwav45DbSoz3SfN/u+XX6oJ
yDPZoK2CjvEM3OMl5618m6Ohl4i37Ok3VaDkkttqeXNni33vDzT0wdwL4CdB7qfN
l5LnY5jCydYQ9wJS5Zc6dkNkRHO7l0s900MKRRTP9gKegnn3GY+7QXaR6XiVTmMa
sIvea1lPSuemBviN9rudLWJN9t5AOorIQBxjiyCx3sQOU2nsujGVFeCeNZsGivhV
jUG+qzWwX31dchQ6Csa5dtQjTIVEcdXx2nFyP7xcN8CVBs3bsLZWRa3tfyEx/qfU
Y55Ygva70odY3GU3Av1e1iQDTRe335wqFFbZYUrJzBAjCTcdAvC8+uAPDyD2mtup
TmtwuvQbdzG+C96lbzdiXSJtwuMq6aE+IIX50sdXJO90QxEkR+fzu3C30DHNyb3+
KU2hZOVq2iWuJY+DZevT5VY3vMFFMXuh6iZT9Y4oqrojFrqrAoKtoApN6M4MB3Hu
RymHrjlTDK9PKHbFbzy6Xgy7DEdqPTbQ2qqbUB1jwc1Y3USqOaOy/KfMXk7M0yXQ
LM+j9tm1t6O+poeS7tSz7CTxX5LqXe6nhJp47UpQ/VxB1PkV3JcYC7CsTNbkqSdP
sp7ZEE1fQyz8xkwSeGb+m///a0yStKnkCsjxf+8xdjy3tj27TDgGO2/OGSx9ESPW
0eiEKV1lIVEnwdc7w+qwfs2j9Kk1QLulfjPEDrK74xLjZeXfYsmoMDqdxK0lKhik
iObjRDTR0/rSa3ObcgWgZvMp4qEB/lRdNEXXr/vtL/HxPd7e9zIUkrTm0adaV7zM
eHd6CNVQJwOAdwnrxnFbXjFmdRpjckDg/OOrAG9exiQ3Xn0bkmpVXF1ipKPLj5KG
GlRO95nyL8MSlxSgCD90OGiUptqyxLoA/+YkTYWtE+RqFuWGcwtYa/SQKPY/qJc8
jYb3MLb20yRUxZWuLCXkm4+qnMWiRw9K2RF5KOqrmJLrTJgq1KPnuWdoQ5PXJSy7
1MORLXwIe33b/kaohj/d4rMZ9JotIly0ZLflaSTu6Om+ZtlszwTXaBy/b12sGV6S
mbxsJz9J8XU1VvQpw8xKk6D0Ud1gMPjjhD+gYji6dJTdDXozUAiDPhamxzXT3xWw
/Obmc5myRxbcauByQ8tn+zIafeEDdNRqB3hLtLhmosZGrG9bYumNmaGR0lfXptGH
YM3cNfkIog2jZqJBHFEHy69ISHcde9poZwolpk/nGCr2RDrG3CeiuD7TbPnJJJWb
YSdxsBgXqKJTJKilkNZ90RfLzk0r+OOG5SZZSzxmbA2zXeqXxplfulhmuyynopI7
/VZfbRUcfH2aUz0iz/bw8rz48J8mXPMoVUdbLD3st4iSJKlO1EzgU3UaBULSKbAg
ApyyrG/+++07n3xyFDLLlU04AbCFWM4WFQh+IBZ0iUgxRLQtsVX12C2MDLoxq8EM
Ovw4ktsF0OWM+ZbxPfPEir217/vJAgCP3GEfr/4iFrtXwLUbbprUyMA5DpNWKKFn
huI4HmCggZGfb+RGO7OBVIfx47+2E33Vsjs9TpyzLZrBOXpG7SLB63ShlfEdEKiC
INvfnEd/wXGAzxaohmIDgcoz6KPtb3hT/YsoVc0Hzl+Pa69nu9P53m81tBpvrTCQ
DY7MBNTv3BgxCb1hfrlDvqNABG3dtSw3V0fJO0FG4bncmq/UWyMms8y/M+LieHvI
0ZjeHrgh/uCd/co2BC7XZkSwvCmYeruP9cCu2meEoBFZG0W1c7zZ4MMLTSa8zVRz
uxSEoQ6dgwhWhHkjGifW94Wzykrd5Cbsu/zgrxjnexdgLs1quf+LdP1iVyva8qI9
zCmz7aIKgz9EWkIWsTqjMBj61NSZWsL64j9X8fzdusWEBBGbBl0zlDxAfqnamQsp
/iuQDRPajBi3iUhOeHrAImiNRn0gEd7y0zWTGX/xoc1VLWwNDj83FSHZf6sDrfWy
ZU7koC1vsvVFOuQLfEY1WUjV/KLGSGzxgaVmYkgIS8wuLPoOufb9puuDk+cUrMvT
QvcgBJI6PVb8kkynmshi5silBATreX6sQmyscOrpmrJ+e/RDtRcif2R9oTd6pGfk
xuxRcxZNQwHvEVQElPBFu7OejtioIGeU799he2pP7h/rL3CPLJUfX4l6b9OrIuK8
aJ/QJnuoNbmvg0omgOig5uuCXVdUi0ENZxMPLieHdQTqpPtbXQ/IuuI1PW9CiG5M
JrqqS1sV/kXwfxGoupmo4B4EeQklnV/kC6jRW9vIMBMp4eBvj00vgevdWKo+bbyY
3bVJM43IOTZ67rmY8vBFGejb8SjmZwrOQB7AmccLHPb6PLlRtLAMCQMWSWLhxstT
GOHkPiDqn1U8k9aAEIAyesyu3jR6aNt9u+w8vRJnyeCze/CKC/ekFMiGIZZDPQZk
AapnQGpKAtjEF/xFlgHTM1GLJJcpZYa1mFIjxsl9MGQortdgVKkKev5xp/IDJEoH
6pTt19i2ufLZxQUyL8by58AsNnMuIWMxaKlXKSgdIWZc3M/vnwlKrff1zTZZChIA
yEwcoXPDu9sLAk9t029fvGujohM7qlZTMetRbMhevF1Zx2/Eylvq5i5Gp8jIbqBE
rNzpOB24qNS0hnUQoU5tUyk1q54JMd106hP7FYFda57kDegjI9OKkNrxEWk04De9
vqKX02xDUFY+gX95a2aiesEszL3qlWWGdtc+W9SDoLnW6n5SmUdjpyXHLCPiqMX3
dCmTyigrvicM7PM0uc6DN2O0ip5CfqvD0r1mWaNNlKK6Gy+oiuL/iunqMvtPeWAl
60Cu2pZJZ8OoYU+DkZ+e41TiWBUs8HX8sHXCbbstqqfbeNMxoyLdSqVKIDnGjH5y
HTzpNS3AsjIJKnmCmya+LnL/+WhWaap+9P+uN6gTE5czSGYBVD9Hh5C1/xtPjUGZ
ifKB14QhxoxL+p942ujPgVEhCk1BxRIO69GAs1+/ugFPfVlMG2bSXhTRTSSCqsQz
XxWngRJx7UJawiVimHsWK+OlMea86o4HKDqqvy+pCmA8ADic1s3Sm9znecS41igF
zzk6OR5faQDTAZgQru8z9Eb0Zxj5PQK+jbT+/iYaDuCoRiQsDDbdfnciVo/nGo7x
Kdpu+fTqd8wu99qEkdP8DZ7ytRYj3FlYNGFWh7tVPOjWodOhgDZqqH73bR09j98R
UvLKYtGC+e/YSR+o5KunhwU3qqOUvri5t+4r33UcshiusIk+7Pa7GPYlw+bmNvzL
tBusZTn4jPNJjb01ipQKDLBTsZjCGUjlesX1doMx0JzueW+qn464lgxu5rbqww1w
502A+owU/xNzzBGRjMRVA5XDR/gwLP/cNuLqs1IukBDkmm0Q7JRI0ncIoXqTyQ8T
76OeS3NXzyc3eOBCFeazstfVazmGQUbCQ2l2Ek/1qA8fzrWut1KKeZj/X7TzKZXU
F2HDbYT2Mz7DALuMrHRjpNwurdHAc/6xXGNzifBwsW4tTNVFNYUvLdgbPp6AHaEr
Prq1f+ywtMEel+FzfkPY6kxFi/JGIL4QUdc28Y0v6PGy8HY3J4k28KjyiRmNOCVv
+naLNzEWq4s+1pCyyEYcpjM0EwBPtrMM4Ph4qzutn/7tBxd5/Awr70UBAis8PfpO
7fG3cCNisECSUYCFSU2D7V7lzWGhb0INzFxePcx0uXaaWjBTFbd68thRJE3TrpN0
NfuRSBEob4C1Fzi4FetcaWyzrYCchd6InG7wBxZzooMUVz+ZHL3Ks9kCORFC77Lp
h9cyg57Mq4ehwL+pjWvpjxkK8FQeU7MxqFXGjJXjNA2+rJQchh8eAvOC9HVDMN5P
WkDVDrslpkdnKlvWwVYIlxV+mY3EByrg0DV1p0bWUcfHfoQ1TETCWT+fpvgwk6Ut
S3Zs9gSFTozfyjtyFCQXqdXqpL8gaP1dO/EZihQWHoSCmMblWDzKcdhgGHxPgoX9
T0If1fn+a9nCYGSGdn9v/T7w70YGbgCAqxKJEPMB/uvsgHUOnQOvslrqzMDC5qEt
S8qPVIvfl7kd+ESOCPVRGbPThr65D7Z9+Xe1BCU2D0sCqC+mTGsyZQr0LvQq+RW6
WZi5l2duUDWyfXgLcW+OwQmUzLPG/+U6TMs7It23I4g4qIMiVwAy3I/zYIUqQgxv
/BJEHmTC3KnhsHap3vTVbJ9Qm+a5Skp3+6ejfscOSxaTvDRDmkBarcIkeo0S3zBN
zgG3h9F3WAFsvHNzWjMsZpF8tGh1ZEorxPwPvz9MDzSXX8SjRpBdBiCIkhcqD0dP
qGfA0GPIUSzSwAAtCaL0ju/3w2QyLHoq1oy7INUoR6UGOqJWFjiOMatshXy65T8+
0vRvlZrApSI21PcSpfWRPL5vIlK92Txvx8LmIAZ7Sp5Mw+p6Bj/7W5WW0oEeMUmu
ekrOIPxxZIreqVmvxa206EiDJvaBlEQW4Ll5jo1wD+DN1CqxS2ERt8tUQg5SbCMt
gACP8PYiHJATwMWrEerBwbdfPbYTgZpiJdpLjY8ubxPGWwjeHuxsV23DP8Qo9O4G
rY/8mzpIp/DlafyR0OGdpnbM/L6H6zr2dcWUDFQQnHtHvBsZo+4WtAreVtmMiM1N
q4br8oq5G/332xGpBpGQu1ftBeR6rZyZ4GprpcnjlgSQzOsaybCtQnvJixVuR+Hd
31TPw2XMfE1mr+YWQVEUaDZRdZeneZqf1EihiJvYqSterbwQ2n3Ci7NONpoupknn
A5CFyvmxIBNS0qWQK7V+KKrwYVTj0oAzB8FRB91FaUXPmRjNWe+NrfoYjyHdJYbX
8CuNbFMTmYdVJtT8/AujD8825yGSK9xVDorGaRNb/VjvEjnuJ73NrdmLD2Xl5Bp8
g34ID1vwTcPcGMnX7aHRW+aFR5STSCBWClQTUTYT1OCo9zDO395hrc5voL4X6NcZ
2EaPts5TDUc4MSgjtTexhD1u6QgOaeBMNn6j1XUTxfEjFfued4pnwOwVdPrAlAaF
X9ZBDrm7tOQFeqo60AB683BdARVs5bgsYU7fiWl/a2WcPpyPwhUwdgFA7gfQWfn5
EiLsmenTx9aJIyueJCvziEyUs/RcOt3faDR5l7HO353oZPV49812YQxgO2jFUCDb
WQu12/4XhTa4wNjNo4VXuXTsflvwChrfxvY6GT08wiSBDsaUDjpHx7ZlOWxuOS1H
MAvNsNT5VYP17yq5zon5MopKNvPMH0NC/WWn7b8JcXeXWcRtA0ExXjC0PKdXVn/Q
TOnCKlg+AggRRNG7I313hhA53ydoWGAKfqhdsGaZQkRVYqaTFi+MsY4y4Lw9z3bF
idmUQK6HT7zQC5doDl3NLuk1qX7fFkCMuR4LkgjuHXGJZz1ost7U7VIJGPceiCEa
mqbohujojTJ+3pMbHI+ddQI8PpIlnSX1pFo0X/+EVk8SR7PAk8Cn6wyhYLceERhT
WE3SdwU0nj8BosISxRrjjPGaKE76JhZG2ekuE+VkFWal9IQfqRw3TI0NUW5Kidcs
LSy7QvuVo8KNxPYxMyffoFv7w705onyCMLOL6ES13x2z+NObD+0W16km9V0CGiyJ
MP2cVS21GGrVCpAjnvn2lpQgW20UNrtTp06hBddozIcT6DcyNGFgQnigLW+GeWFz
2IKUJBwGsPP6yUP52XrCLTtZMIrPex10QFRjNAssIfGro/BSp4NZa8f5c3D2+eXC
iBHiVD4/GuILmHWCJg+pJsG/uKiXuc1GF4RBYvV8QQCz+CtwWKuC6QXqhJsy1+zP
H/VV4GcQhNSJs/i9E4134sL9o4IgLK/jtS1DrTne+lssrF5nN9dh0cTSPKU6AGWC
l6nhML3MvZiKt8PlBkIcQjmSSSWDNuLnLuRr3DoHMrSbaviJ0MP0bFa8ccfJVvLW
TkkBBZAljPDg46E5iXcDA6TS9htqpTy32eIFMjstxCzEBjSt+nCaHDdRQGcl7YCW
Z7UQ/GnDoinV59pdcU8ne9p6UVQDf+d1NiPjp5lVA55BJBVVhMVX3pZPkvoWnRhI
LIzG6is6AqMBKhtwE2leP8V+tiKu4/vqse7yo0kLgmlJdcR7SYDIOyO/acegQQw8
T+TXAV0nWtA+PK4ycjDyxC8TsDw+J9N7Pu0nzZhRdvn4y9IgJBM8l011SH/luopd
gEw20vayJWSQ7eIoWJsaEinFXWdnjfjns6YW7QG9nNmuWO/gtDVmDLE/68wEhZgf
CMpBbXwmAWoRG+wWOFu0SCAQtPoPsVwuwwzJqmiVlucF4z9NlJ23qcCIFvLzWwau
X2YoamD3n3TZb8JR6sOcygH8RbIqTO+393RrAeo2lE/BCXCA/p5TnTyF15XSCDdA
GNwYGqVVdYcj9yEtjfJwYrsWoRsh4GbDbCQTf5T4nIqRQeUkLFTNHXLOkPy8fUCI
oceTGJWqoL+UYVMf3nSZyroVfeaMGHdQsyG68i8zEGpQxrNA6E+NNCqzkT9MGBZT
R1p+kVrzr02hrqujJqmTghFp7wyjmEh7dx4+VTEyngHtWDMTeF5r7ugDxJN2xqUh
HGaWhGV/YgIq+EUpR5JSGzRt5g6Pkm/fbTQG9VS1HseQ5Phm0KUJcZNHZzIRiF1i
j8nc8RJqFzLhZU76+W7BBx15u1mxnMA9JHTjS5ioySEYCnk+iRafABHw625clfn2
IfIYSWQrkXTnyfxehtWDaQdgdIwkS8zSeFzgR6R92oE1ulR6HSZb58ua02ShRIHZ
MGngvgAHdK8iogUbf/H+cJnvmrWVdvKjYYmNYNGFaAFf9ij+KptT/q+9nE8HT1yw
Vo6yy7DrPgozWb0O/obO8v8s/Ae5fA1FXHh5qvrRuLVwDngjNYpIDARyNK0T55Lc
/dIAmTa6Vn+jliI/4qM7+oP58EnSK7VkGklbX3rS70i46/LKGKj3AlzzakDS+NSI
DdYlrkBSThCp88Hnkr2dFoBQEozJVWFgEW51+08LNpD8H/Fg6R8+i32Re7l1fxm7
TkFD3yUOaabZFBW8StCUyr4cR1iQMc56tjdZw6Mweeoi5rXMFRl/2X4BoAVbak50
918ftr6LD6SRzBXHU1Y1HsFFtPmEOKEZbd8b8Dt7ehPReSZLHB9LPFYHwKGRPofI
MGxLmxNigx8DtMnYS4cxq3XnaMt++S0LEByyEAnIJUE/FW2aAxPhd2YAA8Izxe7b
8WE82qAILEgEWP5hw/ufj9H8rOCgFnJeQlyV9Qosn1XRFXH628h4H3B1b5hElrzt
QTKAsjeURjTAgtRNRoTMN8jQRkxSBeOCtOtRVz8Bbx7OrKlXSm5dysxLwLFF3AGn
Miyb7wjB4BzB5rvp5GD+QKUN1B/g1FWNGXpVpZnmAPJ7kZnjf7tN5HPVMNTKWpTV
9/kx31NOGr5BfFenCnvwA7ZFLXDVCyCdfFI+76WBrC2oaTL04+e2fHquh65GwwYf
WKrnnKemvDTwc3+2fHPfvfpxKQvtWVstMURocsobNxoD9MO1ULswoZt75YTuOSfQ
J3gJBJ/Ei9cPAALqA98IOFD7h8T2jld3V7sNsyCVUkKprB6nZAuW4x0hVglSVopT
iB6rQRe0P+y39pqn1A/F/mavuHSUIJpW3Jg+hEjRR5SMqYupBdFPtEWE7R/Wh7D4
krMXJ0stHmNTVxNZYjl/w14nszpF1XRgwmZs8Ob0WGQ4W6NKkgzp2xKaM1AF0TOX
NLGtDDGc6gPX/EJALRUefoV7M09NPFTQA4N/Kwfc3DBfNirykybP6958NxUPLkWK
X3Te8yKT//WQ+29hVlEPzq18MkTnj+cAL9EpEsmRCMuF0BqrGtVi2ObQPIrwdXG+
3JnWVrtP4SwS9N42LJcwr8gYQsNapHAShQD7OIxq5MS5/op0cZ8ge+yM6LbZjJkC
0AUsABkqzCOJW0ZHYvPXR9jUuc70wKVBjqA9SEGis+GG19SZz6koh8zgHeyDPY3M
t1itVBJvtU3edGwkln2+i0LPbyt3WNAUeyo7m9TVzAsXcCYUWD1rG4yYWxB0tVJs
0MHvzBV2zaUhoGCNHLb9pcVkHjYIGzgxp3swvJWNlRnrAFDIIaBc1J0GTf8HjhQv
zaBLiAhvbyKBrmn6VO4MrDhmMEaK32teOwc2ijYwC+6flEIoD0gunL6mJ0FHTpnq
clY5qhekpCQ9OMEuM/B7++x8vncKIKIh5iWCUSAG5rF/9h/bVVCaJ8tUla+XSVwS
84HhM3guAALjrJ1ZiLqKCpYyOJz9Uc3m2aynQaq2gjyMjZ0r+WS8Z0QyCWGsY3g+
Vs5R+M+RbTcRBJJY/wmPfl6xjrEWb/bHI7Oi4gQkRmhZdGj0K6GLg1o4I8JnNpfc
0W27/jNmQW90piUl40i3VDM6dRoZdyucAfymcfA+A7kcSlpxATrCZT9pK+HZ0apR
af+GlGATsjzle/0kJ8wzxf8+jnMQVRwAEdAcIkB+th3d/kUQY6wZSOwmuYE2OjVz
qdZ68Zly9y5tf4b7j9YMwSHEIr2sERzqHEPcWSwUTFnjZIPlbmmynsj94ZDj3qIE
zkhvBF4OhEaXvatrSfax039jgJ5cCDEag2bgjtmVp9VqDuqqwnL6T1i5rxeRwErm
vhHlZxKqFRW/5GIRMpe1ydhuvPin3m4IV/B4jzRunhVT8ZTteC+LgoCTLwXpQL6k
BvSxEdO2Cq3SqnTEFDYft7brSgVrfNPLrr9iAssyEXTS6CEDN97t0izYSlzr/Ro5
r9ND3E69W4To5qCHH+Nrw4FfQCAPXnA0GLaE/HQsqrUM5vvzndZCfYNn3QVbgOsm
268tZLarjhNB1CNrmzQpTNndWRaDGXDgtTsDyYRNKhxxukJrldIpMVYdLoeqPEqs
zxhBWv1PWUxZAxzDWozyJbYxmN1cFlhbsv6+DT/auwilZ5NLfReJYphFufyM2dSc
ibhkwuYZD2MY01KzXW21D3aNOADn4IS5UiSC9wzZ1gqv+s5hJ4my3bhPIKfOFXH9
8MJbmLfi2+HBD7uoyFZsxRSpEkpbbTZtmPZO2H/4bq9GeRZ9cYKysDvZrjSrGUEi
Kbc3EKMLFvOpq7F6N8oQoxaXrz6ZKG2SJJgla0ELcmVcNlpTuQpz02q/YhPmVPOT
ZjXAsGy0c2J+zAJFYSDtdXErwdGkv1L29YdfPDUV0qCJyKaW2nqQ8WUkxEkBaTZH
hpsNz300IUbugKae2Lx3uujzHwY6agjTeewi9ibaKEahffqTKVFP2tA/iLxlPYl9
OfcQgD+zjBl44Xb06KIqiG/QKr5ca1k21JwvqwNZ+3QwmN78EO3jpVWaiC4tfL9x
L4BE3FnMNM++Jh93sgrXS5IXS4H8lzx+xK0K6/QgNyEc8lRM7Pc2vcj26K+gb1/o
lysx/IznMawnxDxCw7M7Mh4RtOuZtYauvTrH+IO8K0ZoIbz+p/7KgN0X/QBhJtcE
SEciOO598CA7/Aoo6TW+0ls4X9je2824hjb0SFFd1ZIOwoFiYSvpi38MUsdv+rRL
CkGtCVUZHBBp+5msrW1TYLhSVc/kl8U7CL5GdNZ1DP5SZ+4J4QNmX+P7hCrasfvz
Rb1cCbmfQyZnwrrMTktK2WrqNb0Z4Cc7v0WxgMm66YUWTx0lxWaMlsXm63MIeOhJ
6rew5S0x5PmC3vqA7Lk3mvRHKTKHndNUv+4TeiEhc2LldgmWr3uXUgFaAtIjIMVf
5cITAhl0RNlJPcE48BGxImPV0Eya4ttRSJy1GiDTnxVgezRqtE6dU1sQmdPzudsm
mpZT8ZZUGMAwOPp1gG6EILyIliHf38i8L1qCJC1V5EiNHwIwCg3sXDOk7+8YwB4L
fnHzgZciJ/LX/us3Zh3k7PVV9uwNwPBl+aBiXxKRX9IBCQVmhTaLMA/vIBRoQxNH
emy/idNZFll+f56W3rK5eAQrXoFG/uT6UQjNx4PQxXXTaxbYX35LD3e2js7kIP1x
9avUL5eDVxeRIP7VcF/VtvvMXPJP9XHpM/3rHhqsBnJz3Netf3s9K5a4TqE4atEm
W2YFiiig3SPQwUV/MSl2B158dJvGTdzFG0NnKPyhDA4F4mLkLx9g3rVvCuNbibFA
vI3/t/Tw6h3wpo7Hj/0OHuqLgRadkTzw5QjbVAnmY9Vd1OQFqZCqHw6ubgFfFmvl
GfKaXC83rWO0wRhnhlHc7NMHCqKfPKd9M/jDEUf9NSQNxSmKPOVPXlJm6skbFTEL
ULHbPa/Ah52bEHfeIOAwyrDSjqUg88jNFVqgx/6xalOeEmd7AK34OKfPV/1eYwkX
MDiYFOsoSZVBwgPqMiQNaVsH0CpFgYGML96RheKVqN+jn1IgIjV5L1biwfcaggDP
J4NLOOzFjkdFpqd2/Dlm6KBifhtwp6yZSGHYDmplG8nMyfSFIkJoN6yQGZ80kn03
95Z1Gm/jnKleGw1/QG0l15Sop8ydENU6iBZr2cyLsRM1O36yNI061BSqpptRwANd
GT44uroDZ9G3RfUgmBrAWiFYeUyl+e4HryrEQiC1McnwyHjdR1lMSBbLaj6UCKrJ
rDHOPUuZYnRA/jglBfzbnXPJFGqypSNn2rh77AK/l9BASmI5cEsfQ+XXSZP4Z5Qp
Ga+WAdBR1taEszWv22QLiBe6HJD2Nn7GVeIWOB13OgFjN87ZLXzUYsjWXmoh2/8m
kA7xM6k43DwXmsSSxkrg3IgwoOlmRoCAFexFAUQgiUkQxuGjpi5eLyN6vogaz4S9
w/y7fYhRTWLC/UKyiD9HuXKG8S0K0mZUFm1vYWx4fFltXfycF3XD/wET4K6m2HrI
XIIasPi/O8xyl7TOSahmsgKLjHXF82XTGRqDu3NpSlPeQ9gNlcoR2K2oa+lsc6gJ
7k6FngNlNlZ1QL69z0cyYGSKio1GiQWO405r02XI7eExTIstkxwyS6aOMrnRWZYo
XoiRUgg/QMqVSSF479/PxqMJ8W00MgyAg0MWZVULF7dE1cUBI3CsQRNLB9VyEOci
zp3OMUrD/Hg0wpwvw4TdWMayhCsdsTzi0zOZjlxfeB8/ZytzGQRLWg7+idJ3X5FU
eKO4ClcFLambqj93pKbeYO9nHralcx2mquPZOaDtJImvfSLAk7RkV7iME9lj5Cs8
iWGq83Dqxmjb5dvNflSlJwsrutdyXGjrA4wAU7gJTNH1BSw+B/9XO0mgi65OWKP5
J/k5rSyE6CWctp8XTd4Vv2EQTbHkPKPZYnmaW3DbLH9etauwNyxWqMXBZwuvDc83
tHw7Y8VcVGy5x8ZOc3ciQgZe3P/wo3Nezz67VbhmOWRvVpmPIl1HROQmFRC5PiYV
fp30Fufwq1OYu6Kp1R/wAiXXQ0dFhM7Z0/aOOw7uSktBwOWGcEMXAkAUTIScELhv
lJmraU9rIy7sX8IeGQ26Jy8AFhI85jNa/1mjdGIrJKIydY+/GaNytsuYfqRPyTGK
qElFeF0S0Ztl8j5lZl1GNXtfq5OuUCsn2/MGYUPKaPmLq+wzza9z6w3D8fL7vGv8
KKRA3X60ceaGjIJm5hGXsWU9HTnxQJTgEKHuqmh0cdRRTQnGnro3o2xFEHC7SR84
/efsQjUrvEvs/PxzxOPV/sZHID14apuq8tPGnkev5NS6iLFUHD3oGBgXx32Eg1h3
ImjjOcB0m6BmPENI3rhFOgaFWOAL/fCO3qemOPsi9Be9KFvgRWKUvo0vKPgoNIph
rKwZrIOnchAsn0cV5/2X66zpVJeWozZ1/JyUeWN/OSYSNgDCTHwneWkBHo4+T/Qf
rfU3U5bgcvAF/1ZjN7sjL6+JZ7owkD9nmfAGH8aIIFSoZ7brBbE9ctTe22TgJeNL
tqcLRPojywJ0QZy/gS2W6V1JW8lTJxX3l77C8oJpCLfoZji64eRy4FbbErS09qGj
DAQHnZPVFpjlW2wug2EUlbHl0N3+NEDeO+NjT4MaCN90rp5YDgjM/hugNQ6qbw+k
Z3QEQO+G4ubpOSbGsQi00+dIrmOb6X2GV92Pi03erwDW+ddvxl+PxuCdjE+1CwRu
JIAJmo8j6SUpGO+vfsdcWN24MjrKVgrKtFFCinmcwWt7m/lEgiB6dFNjC1tMJRUv
2gdxzH+MwzE9n9IwVUz/B0B5SYvrXLPAbRiYCIxkyrKdDI0UVIib4nkLWCRZum+r
dBZjjtSmhzghlRmR4FE/82jjLwfPgE2S9znOUqni/14+Eel7vycRuwd3sh6QBXp2
K4yvQcewWCYDVfvH90VbLEkQpEMebmHF/M0RW4B66NQxHRCxLl7oH9HAleDUWk/4
hjruBtQ3jHXo2eKTGz1rJy67EVL1aVEr/y2u+/03F3+zzAX+h/Ei29541cEsCbVY
CghzU2ynxpc2+haCtUdPbAbtFCsZHo4F/9+8LYrPFIUfGzp8+T7Cr+INOCQdZmwb
k2JgO0FlcnawXhO42rfFw04N2Zpy0re0XotCzjvFmlnbk/Ay5VcGxWXtnkHMCxXa
iJMIfnG7VK0wUr1UzjpykYQjPN1oCbOom4zl9b8uGl6NZtBOL7mod+fIsXDcxD5t
X/hf+OjM6hU1Dkl9FEBqHi5UJn2LLH+rmy/ofoWsl0b3dSgOSN1G7nXGgeAzRUO7
+raWJ/RhOB24PAKse6yuNamwkkP/TXWOyr12bkd3cghLhfahY0enQ+mWiSuf20y8
R788QfoBsM/2yqfuU9ROAskaYGa/4dmAEAcTOPZt8nfqBat1bpZEMerGb15FPchv
rvE54/AzKA+wptITZ44NLO9HNzK2MbQuJ2PRlW1tRLnRjblX4IoDHbXy++5KSTjf
C5/l7BnxY6Fn5pWTbLldyZLp51BmfOTZvjEoDf4PAmGvWLKGhNh6o4/LC0cF67DM
wbcMe5ort71NNRwTUn3bBXj+NhxX6mbu4e+tCbNUuh41SdwcWXLke8IW1JrOmZBX
FkLdwaj90tfO+DIhJGGEDm6b4YZqHfhdegF+Ey4r92/y0Zok1T1nDz7eor3CNbBq
WCIVEjGKOCwFkuhNVph8XQmrspcvbzQtRE/Wkk4/9evNVsYnflrvJ44oLkjRvyBq
qNOXMhvAxVYCa3TUcaRjhfz9IfiuC9Gss4KruD0C/CRWscK3PpEBIpm2Z0aEoYOB
EwiqqXl2WLQ/sjDhL+GEesl8TFceKkI65TIrAtB0JeHjAd48wjGQLrJeK61b/xSY
B8IhWXL4ZgWoQveE4u+v9l6EWcTZDJx20ezXmoyR4C/r89Iulg8QGqZ+n6iF8QSr
Z0GDUXyLokQ6ZvsTJUvSJEyyvygnShNyO1cqz4/Yfazq6JkAVWM654MMH2QXyUir
XnhXgLcGDsDtPnWVgwZXRsydi7g018Sk6CKOe/pH6QyTrDqMOczxJ2cC6fVDbECK
rvMvvL+NHzGlRGpgCvONq32qDvOB6rjv4r5vyK/Vig8RhJiEhH/G01NePVaPooQz
2xM9EE41mGRuGsV25186Na76h0M85O1ZUZ9/pl4Nqd5Q2DxM0E56Dja87lZ3vYFT
aQf0xwTVecyrCsc8Jndx031oCKekbBtd6NO3AACoJDW8dSvTry1B2/drD93I0tBP
sBrRFN5Fn4ROlgASRBxPkV5wfztFgrBI0B8rz5MBxkX4RyMZNGSfl/7pMswqc2zB
OpMQBmxmjOeMichYu5mOO09tu71A/h1VDhtj7XJRSnJCPvydm5OlL9cPCz/M5bFb
8xxTSPzWCq0CEZpd5A4bnQWyPtS4gC2J4CMTZY0eZ9W78dwcnTTJM/BTX+RkjYk1
PNTsZBal+Uth4rTB5CR5uN/fDwrLzzDtgwzZN0chlUM+irzMy9dp0nPB3PvhRtRM
qNjuIo2679cCV9WkM/muK+pzUUdcCLKV9nsbnmvSjh7J6oYPKJ57pgvg97WQPEik
55sTVtsKsecqPlwvMNrFavIHiRgiTJqWhte38q/k0sNqxbGZLXnjzjS6Uma2sX2k
2nv2lztO7azFtFcyXkYOJabWuRB4DTiUtLEKdyF3NO4ids6jKKnx01RPhfWmQ3nK
0YQkCVTrRsl8ZnNCD7Z0OorWQENZFR7oLtDU/KJQmyijPTQBdAapb+aPSuMw9IgW
JPLDClnLV9btyXf08rPYLMbs9XHpKXYSE/apc081XlUGkj3Jl4hDSg9WfJtcxwj4
yDoGPqS2cvf7UYext+qiWw3kIzOqPEliWxIKDAj1BYLkc5vt/jR3RFVTOEiaHZoj
PNUtUPNnkPfkXMw6ZCIT8ZYe7pAgPS0higJiJHnOSLRVZ2FMF7ARqiY6rkc/BfN7
GBkRYZM7QtGilNaqhYEluPBvDmBQ3lruySBEIyWJ/laKPu5Nzo9i6sIFaIX2tbIT
rdsbBq2o8iGJPrfMYV8W6G48nwjB7v1uz0owQ5qjIQJ/+8Ipf1r6hLu2LAZ5x0DN
FA+h4tuWXYKGFo+ODy7lxqAkSKubgAhlrnt18yDru5zbSvL9Xnqqe+ifOE/JhxsJ
ZPfbO+T1o9PJ0EE3qO93c64/Pmc4N95tZhduAGLp2vXoRqnJ8CFNotIwVmWMG6If
HRqx6DOzGWk8aehbsKK5HhWwtIqcdQtPGZKTJ6VwiRhYGOSZODxcSJN74jfBNIyB
DIRfOrkesz82fFqcLvQYjUQZi0CG9XRhKCspKylQZFJi3Fac2wh52sOWxlHqHKvc
eUf59BMjTRqxwP7RUcAE1slWmAAcAiwYVfX8PiG5dzvyuHQNBdYMP1wfTSneoIW7
aNtyiJ0nmDfbJA8ZaEhzer6EAQO8NpN79n4OFJqaeg9hAKiSjBWRE7AFMyPKCtek
tU7ts6XkapjWfds3SUnjSI5/aWZLjbv8pIgoloNL8loDdi2dpA/sirX980bV+ZoM
GRibF4u6gj6byam7dq0WtxdBYlPC3iukIothTylm4pd+B9zLg/uBaJ/QBpMQIeMZ
T+5vfIALrc5NOShVO5awSBbMF1WLZebnZPK7EXGDB1Bp0iNCdNSqcw8gzBylNWaN
WqYv3Or2mK8UEmFXbn+3EBE8pXoGYuazmgj0Ec62Xvs9CbaPsfWnST6LGb5ZNg1F
aR926leInK3r65/OfXfpHKpzzmfW1zYZEhnqLW+2occvAJ8XEUYaet7ui3fNneZz
vGsu5v7zKJckVyrTcjb4vOtasoBLKJyTxSDaAwumakpnw1qPvelEsFWq1uI+OvIC
0Sq+N3M/EzcSHk7zV9ZOwwoRewkD6GLbuTmzx3cIL7JPo/a7ZR4tWguSLPO339+N
opJz4Gk3WZvsDYeF9jSSX42vDT6jnkxJ83yNoWtaDjYD87tMxg1LM5xwHU+z3xLt
/K8FB0zJgHRipzpR3z4qOdaXBej5wnwb/Livi2M0U8jSVCHQQvPIKFXT4+0s2a01
3xD6vjQFiaEqsJwI6FrLVjHHPffG8Fn8AnDHgmUpZC+DfG8p3DA/Qm4Rgw+V8avV
Wu1zBcSiEV2wyqPi14Qd3pc93jFxXj410ykrFv2jPrNQfXDySiBXvsU2SXki4wnf
i6G9EAvnDorCyt7GpvuroN77P0LvbB+Nb4J4dzev+6+ZQlZFWk0t+ILTFy7OaAGp
8DeUx5wNFgbEqSQfQwgOWsoN0dnGXfvdjJMsNspcRQCKeC+hy4P50AgNaKyBepiA
kiFaIUd9lcHa5lC89Pxldynvdhk4nKJD+xHmyh0DfIVNnOaqStO98Iq1gVh/1eeW
+Oq43CDcHWHIwDzt/eoZLt9Qxsf7l//Y8/ywX62Q+bO5j9++DgHzKpzPzlowYuzW
TVoetNGByl+2AN6/IStqUUxhG0uzDhTYi6WE93QjvjiYphfyz1AAcWlkUYWw1+Bv
CF6ucMuc3f6EFZYrB484+OKQw7gcYmHGF55lSEcyRwfelekaifu4Irw/SYuaG03k
ovDUhuHGLU8VpwHQpbq1qvZhYM4K+ZMLikGIcgQ4dvoeTSDFVS5BmW9+0BaZPPBN
3idpuywd/N+8RSJ6qhIXFfibolUGJo8PBq/iFI1l1N2R0jvxlyVw0Gjb9uTrAiFU
JyDgUQGkiz28T8wJGYfVkGcRHqnB9LYisuUTMevIImbHPQZFTduF7nIzrKoyV9uh
q9EljPkFNmtEo5XFiuuuPa042buIUOjXTtvQNuZX+U49fRKGxp1FiKmok5FWEGG+
+Zx09Ct9MY2l95aifGqn7daQ/ItanPW78RTWh6MpDqksr9vBB0nNpGSAmx9/+kCG
H2lqFBXmiberDpJbYuzNuuJUTj+1MztOi0JhjZbFxsnD2MUBZfoHOQlFg8ISMLbP
GxdLYhjJlMxjZ+ze1h3Q+ibx7asoT9Y+9uNa0cxt3OSxhENYYqZEyKnJMWjTPVCp
lVBOCWtaZZ+kFoq192+bQP+VWeZvaOPjxuEHXlS+U3jJpbNgXuvQAv4Jsu0czqyk
g+JJgMJrw+9tOxqYpL4dEbOijrgzoi8YbDy26jeoQZx6w9zjcvrEwe2ocVP5ZwtK
J0JIHcj3Ooq8csDGWBBUmL9Cm2W1QW61FE2va+NN9n+kZYTFbEbeQyXubEOKuTFT
d7rxco1RYRWaI/KSP6+burqB837rwb/pPFAaBQ/lr5Ihws2xPyQjt+fk7Citxixe
qpQQ4CrR+CaNRn9ZI7cM/a4rN5Ez9BNNyE9bJTrdDtzWDJoEb6tA3n7RQhsOrF5B
PJCmbL2Dj07mmS3438cmxzAp9W4Us/x5CbC5StgDgZ7I0LxC2fwhmTqZh1kgFtik
+DARkZnj7/52e/hQz4fQN6Kc1euIQZ8mjA7aVgez9NAMz1+SN8q+B2WGDVpJTf3H
fuOiiqkRWUe3srYkjpZq3K269uAKGa1sll8qssiql7MOQlXGFyBVk3PIcij9Jwe1
JUEOJq1IEEWvIeJkFQth+aw0nRop2mHAggDzanMOEjBLEflFhrGo+rYiq7sLi5d/
uWPMQPbL0KI9XISTshF7WqfVjIuQeM+69MZcFcNNpB5KLb0kIHv5W6u/ZxY4YEqy
jfgFjNoNw3b4KT2mkDfQf1hSaZ99mtWOYIMwM/wkYyjLjaeGdjpjWEk6nHaH7RA8
Hm9lpxwD9z4hMn/jbROggS6+tuVrRqqicc2ADBPx3jY7LcyRYAF365mVBvopf4PH
MDlMIue2G/LeyJATqEpum3ruTmgQwRVj/56JGhXeM2aKdfZmc7BgFvwRYVKSp9rc
pb1J8psgQGrKRRgEDXkdr0Goa1LTSkjnzgjutPsGT/DO0sU9kRNZF1w7yM5nUHE4
QWVuEhWuOxSFglQu8SZQtb3nVaGJcsiVgUM66Jk0JpD6qoGGzKQCIheWY1GeAmrx
KqjohT475EYH7fa0NSx6ridXd4cK5QkOZeAS338AWmvuG6ByVQX3P3tmDVsq1szA
y6YSI2fZz38WTNA0IGbnHmccMcfooty5oZzCncoCsdNg/evOqAS6JBnwMeO0UsQ3
TmLTL/eqNHgV3dDK19/ycE3xDr+5EeT+HjVCEqZ8cxX+Ulp/LMRnUMHOHmLu9uW5
v6gDGA/TnoeAZZTBEsIVFqkkLBW99/iy5UGu3DOmW55r5oEYdyb2xwsXPMs8myGM
LZWpbg0IgLHVp59WZlcnez3xoZd2D8BLf0Hu4Ah4X+ILmp5D5JRLZBUeJ2dOEiJR
j58myuvQ83xo/8+bp6SdBwWKVfO5Wwh5hUEd0kWrWSVnBdQ7XbUr8rQO7Xe4jYtj
EXC5l1CrNctKcqKuFHwwo1RtRM/uqCkN7MZhkg56CwBPr5j/4L23adFsiMwJLPnN
/+ZjBFU+Hfspis/JXVhjTRZwClIqX6pMwhNU5khjomFONpdgQ2AeKcKCS6rnWAux
DZUr9toY+mJhMC+ftEIfCfuH/lYgKJhzCQ9E2N4ciZOlaIMUqszznZsxfDU7c9TM
1IaRVCmC9EE7UKn7iDpjfNh2h5qcZ41k2mcrzy0YC3Vl02U2jLNCqUPOhsMw+lKR
KYMxEj4CplPW4Lrx3/qGt0iBmLHBdfpkiyny2Zp1gGdDc9o7n3ril4Vtr+zDf9D1
LXix3q3SdAnuKSmme9L9qoRDEiAHKTG4nuU84w0jUkhRHXqo2isxQfDYPxKq+Y4P
GO789GJKPIgyigDBBhycP7uEmanL6E++kHe+Uz6OWBfWr/C2FF4GpgsMHciOU5FE
sT2FTyEoFQia+h3DyMI3OMK8WKWBTgUeoMU3qhL3+686XM3CpubrJuA7fmfYafn7
q0jvCMPrq5fOzPxQpOD1dMDxH0FPtHUZnhNbwkKLFNjHWRBMv15TIY9uFDgu+XeY
Zs1fhgRIQXIa/o+p8RVzyaA6QFauccibRi2CZ2jlgE6WRj2XO+SUsl0sOksjXcG1
TfvLmgnx0bZ3++WSJTc2v22RNWh+tZgBwfNlB0ov10pw8/didrblcpJ/lIP77s3C
e6L+1JCAemZVUf3/kOgfKwY3YLumxJexAzHGEn9WWIZDY7xOVXncwBbca5l91905
QOd/DtRbLItorW/kcRYN1Ad0WiK6iq5yRyH/lsyKIuY70pFyRexSoOF38UuByMHP
Jpy0OiAlU3p+0A4TP72ItYLrZan9ckquYWkPmMpRgVTyndERQDEPCMa2BQTjhQ7r
IYt+kz16h8fZCg+mjU7/8TtXOXW2cafejssnruFwSWnobiVMLFTjAeLz6YR0X713
Hxa16qK74aucwNwQ1a3J6I9cM+e+CTpsQAdnLdDWH+e6mFF4p65eOyBRAb9c2CBt
kNgsuOt+IgpuYCIlLX4E2us8M6uXYW6kclKoEDI6tKpOQCcBBjFW4xsKol41vg2G
jrte+Mo0vrkP/zdZZLLwOjudpRkMPBw436/SgW6q5mca4ouUn2pr3Ax8LM0QC88L
Xt2NFPKXgt9254XA8ZHv30JyOtVAJogR+uqezSo7NWA7RDX/5D4adXpKtClZw0OK
/QPO6vxb4F/DlMARTmHw++GDpu/3BleSFOx+rtRP/b+CygcZo59IBlPswXXUVbVQ
LucqeJJQMuiDAdgo6t6E6tDKhDgJP99nUPHBl2nRrdeEzox6k2qsJesqTrstpWVz
E011IS6EQWjWggjGpEnn63SE/gc7nISkE+udQVbTUsi+E+uynRguwQ3xsTL57Ouu
wNGDvHk+43du/jeFkezzvbbNyaEbbGwYY8sfKvgDdKLVkDneAlfBhpylILaJB39D
I70RVmVHW7z01GrIrKluAuz45gYeGsGEnki+B2WiCyFluTF1UZmvS6ZwAJP+Okn/
rEfeN8hHlVcGFb3pUW1vLGwkGZW/0VNdDjY7XSCPuIuPJZ3NECbQyNlAY8pLSsqz
LOWQ5VrI7WFC9fA2mUeydkKFTN7WkhhXdNggT6B/Awn8RlJRrT1o3nvLaayD2uev
bDsMKr1QO14T3/GvI2tuF/sa4/5iplKHHe0XxknyisFrC5e2A+lojmIs6hiijuC8
U2ZiJsdgfuuK/8vVqOoLvva4aczOMntvWLA7FwDWMMazPSUhm2/1ouj4StUTx81O
tgIOqP6LziUPlV8gsTCWlqjsptSaTX7sIiMSn025PqwM0sViMXXN2Bfjqxr/VwQS
423lLGb/ZxuUjSxUtmnawZHj743IYql00/ib/h3IGhyfuneFnz7OfYqHPdYwD+Sk
eNFh34mlml5TSFkjNuSyAanm9dieVWZx6HhQeJ7NuzibETIGmqNnwm3Udw3TMW8d
ysd/xtiY+akJx+jNp9wFMWFb/FEHQ50yDN/JD9D/q+bc7TJnrWw2ife0C6Qv32bE
WIyg7+eNEHLhC7qgBPZZRwl1B9HIYcTi7FIwjFTZSgI/MLEOlND6et5WplCCwybd
6SpqPT7rCmBDBAJFsjpJrbTw4cHmD2XccYDYCpNZeMzXT8vXQ6cWGJebGrW503Kb
pWj36GbvxAevpSCaT41CFFIkP3GlnZPUxMpjyualNvEFvWtzpmjUGONFd8I/XVxS
jqWuKe7f7e13bBd52xCzNkbhlinR+02mzc/MtwC8k08UgPr0Tte4fg6dJUeJrG1w
FIg79Zeui8d7D1CfkkDZgVgaeVhi+wIllCnph85fBf5G9JwOtwnxAMlwhOxfZQxv
o9j7B4P6ymUQTnGleDjCMa/T3P1eM8eVleIq/mgAeTlOMZLzI9j/pF8j973xONYP
jQgRg1da+y+4YP3CjxpvXMoemqXzdytBY2nswOeXElVDJKzLEjtEsnBKcZNCAprL
ciIkL7PpAfOQBA8WFMvu8Pt8Q/4WNDbucLO6Tp0kGriAdnPIc9P5/OH+rEtXClBl
jLU3P3iryl7Rpb91z7uHHRrFHDRGWuWwJvd9Bka05Jhmm0vbRVQ8OvarfhEktuUM
Rvy/XR7BNUlGMnMpGUs78UuXo1PCPC7zHWeRHVLKYlmceaDadfuZslHuV8kSzIYY
Foom+iHEd71yyCBKYC3X44mSH0etrLOQCGexB1wJuJg8j4xb94LS0uMZr1uPkoit
aLc2lIm/UbGXd61Iw18M+rSCElo1TyRaMCKfzq5mdz8oMYmQr+dVm+LxP04SbHZt
kdur0V58oRAbSSn0HPr8HRv2tNeUvc/02Rt6Py3FM2gh9agLRkR17s7a5jBuhcig
vU9ZGjPewI440ATMENqVjI0qPHpNWy8GlXZbsykXd+nIh/88aSuJSTUyAjbU9vWk
cGuYO+jcq8Gygygc9eOgMKNgYHrOhJ7xHG9ryyBPrMby3MwvVtoKQeCKwjyipY/6
tR0EAQwH7pT0VssLcEXctGBp3Oxe3x5HXmI79OGqIWWU8IlfWmEi9+T7r2kcVm83
BnAOI6yr/r8kCsPZLva9T3D+l3l74ach/HeJoU8PIsiC9utVFeW/urQgIv6Sf+9g
rCYr3HkW8dFd/E9y7FhAznTaEjYUYYAVO8/GjdhuX1twiNqDgJqtkfp1d5WAFgpj
NAjNmGRKGYdkaVofL2DlT+9XxNn7WtIGM1HLsmbNxxvmr8Bd7097qy0ybIan3beW
r0HihovGIqV5kYLEa3L8RYgy4d/wU+pY1/uqR2EvDqAS+DOQVBbIk4f41/68BYrV
/DMGB/9vGsTjoRKbGMa27i+BcRAl7mFBhQYj3oz0lccvwcIMo3d2V+sJ23OAvnvO
2AnYVdf1WRtjI+JyBeAqxGFBUi5cK9Y3mJRLTk9BJIJGkZ4URq2TfXlgY2x6laFJ
YVpNg8mp9jbu62cVE3hFPKHl6UYmWtaulHnovqnSFT9vItNTzXvMxapa48naS/tm
vmvkuySHuxA17CKvMoO4U5NONDxBsC4xYbLeEYNRQjuVmG5Wpn5flKOVIxlI7SZj
NSqJOZgmCDhYIoGGG//PriVHfxaxWcOOs/YEgUQzbSbXtCR1mpRrfV5uEKfgFcz4
0WVZOmz259PN7HmSZ3EMweFbnSARmvjcj07WwVNJ1XRfzerCgUJcKu+HbTCbvjv9
nDuc/FVXAA4v66OqUTAX84jRUqc27uUHSo2Jbrp+L8FG0WbC3ORkFYbdidua1TiF
jYiItrIntUMTNpc1s/P40fa7Vn7gZXJ7UbSpTUukqRH9kEkaqzDc4CZFy4QoFbN9
+rl1D0z3t83MhdvmAnByyXJBRtt0vFzpsREWhGIoitH8AsuywSOhfgV2zpl2i1WZ
Ib5Gf/2W3FXziPpgiOxcYbUfE/L1RxlF0svBiP3Ru9pIMgsxp+wtD3F0Jsba6h9E
ZHtiW8rVnezKZATXqNJJP/kfkFbIGhEkhPx4ilcP1DSEzRqnmoAhgo+VVEnCNlY4
BMEzuj0HJJ3Itwiqj4WVdIkluV/9PBTNDHZx+WK+rvOQxFoBb+/cNOSco0tSJm/7
Hgfa7O2z3HRQs+fYyUpZVDZS8YAdnjEYA0COXMD+N30rt0gQUE56I9eBcb/PuSjW
TkLLq7x8MkIiy23qdS4uW6FD7xjrDri16zf2ksUD79UeLcoqGJIc9CTkq0bvz5Nq
AejFmn29ikOZjO6gJ7X8MwpWutqdI2UV0cGNQw7RaZAkWJVAQYKqTxGXQ0Qp8jzf
mMuqBMVTBZ+1DlGin/LOd9SM/ymFINjn6g+eI/FIsbWIC/xRXTuqHrxEsWctAiYG
9rxpX4iH2jDqS43Uc5SSIKeGM0LyIlSKzEjsynPZeMw2RB+WT3C5/QxnveDV55n7
JRhgrqFxOJ9bNE1CaP60NG5Ush9F05xveuuOElBqYxKEkGHUtSdEOS0NZEEDGvLk
eNtScqIcFTkwKDaOv48kMrpZgMIijVkKIqutFMFl6PBxAOX0pSShpgtZ9KkdudQk
9v4LMkqRrMUCF91Nixru6Pz1cGVgxjOifzmqoLSBsPPCSYQX3IoR+PuHuzUpNrzl
/XVx/NNX+w5dFk8LTMHoNgpJm7VnJRsiHg59sKRrQl+kXbLF/55NrWtbM1ehf/tq
bN3bfPtdxQYdcCn6RUNRycm72J7to/eDkMDhZTSRYkdBwHp0pTkuolS4rwUetXCq
UnYoh96r0V9Ti+EqtyfRyXa3K/kpvnU3YPyZAKenjSBXseGGL5Ny58wDfKbJaEBR
3RCUxUOCzlhrdWoEpyK3BwFxPZHdn84GCT1gXYXib5mBT3Vnjyl2O060nmlt8h5P
y03QuHpYO1c7dbzhqYRs7u0oJ73I4gTMxxEAL418JE8WIF7efVL/4bdel1CAfmXx
G1j2m5lO896AukUrESb5X2lgxSBQ3W62JLu10AbrD+g0jvtV+aZvI+M3P5LtXowb
E5x/wxFlgW469ALNXwTAD2HTe01ogZm4KhwIDTMB1jQvZKIRdUmL6vruvdp/GRjY
3N/i4rmHQHVJt8e+AIWiqSCxk+Zj/ea+bb9YQX89C0MJpz2umRtoKkeStb1gO2NY
w5YoBsD8YEuldbPM/u0vJNTI3M/C84KKxSTBjEJWNWbGhbCebHj+IVYUJwfuas0M
9NcNANWNZEi9CFhcdmqyAF/d1l/XxDxTUT1Mxn+qwH3fGWv2ZnNpvMw7vca+NfnR
qBppyx9Gc8VnlBLbDDqS86g7wRPIAtDAKbKPpxfHCZNCFbdidCatlLuMP1EdK/kZ
ia1Eu/3SIapnswGMsIx7lI/LSHwz501LVcUDWmvarZAv3miESxvrRig3F3SibVc2
5/saxquLlsaRfc72cJHAVqmliZlPtcdz9JITPkxoHDKMjbuHSCxp1phEipc3aX30
6J8qWGf1eUFhuB5e9tuPImzPi0wPBsGC81g0VOwmyTvbC/f2iG7YCfA39fzfrKa6
dINrq7enqqH/QFrkgGMMGqzGxqy/6Vn9CpjF586jRCX36UUFro/Lijz/4zbPcoHL
9MYmDCIHFBkcL7ZPIPZRvFKWdCLtXZuqxpOsaSElT5goZA96RHB114Wfcl/Z7kdN
wRsajeighr0eQrSFTtxPMMQI86UBIYScH0QSSK8k3E7TOTmBrz9tuNhdBJPiuIzV
yiSNu5S7cZvzcySgyr8WKEH84Cm1rOw35In7iJ60sX9s7vTSXEsVB5ZBcwbBZM6u
i4snJFPnnJPQL/6m2pm41ZQ45zlyaD1p46NkMcrbhMogjn0unftszL9TNvvxAYYx
iqzuYTH/W0mndHcXbFm8vBLZy+sCytg2ZX354iyCmNIsAAEuk+Yzgb3fWxENz266
aijvxPnKMe5FsQewHuyvQEmCF07x2/CCSxxQ4lFE+C6zzUk+n8wYk+Dboa6CUKZL
0l20GQ2g+JFeN3l+0BipuaxOMP6Iowbjm7bT0nCOeD/QcRn1Y/aWbDE8SG70NEXy
BhgUt5EkBUomwT62gx2pEogm0bsM3WnMCcXpqePRgwJxOZGVxJVT5KkRShO3gAZ0
bgzZz3HFcHWod/069L0lvX/e/iq/C8gUj8JqAlL/9ZWJnOz3fAYmP27QkeIQiQAm
9sHJ2BQRewYKB/R2Zf68JmwG++7AMK281GWHooZC49M6gWlptdutqv2piBdLbpYV
yT4Yb7OrZy6wYihzeD+vwvgwQRskBXz7s3sP2yxJA0aFqUqAgrAvEHoLC67mE2Pb
24/eIlPvAwSWXNcNKjgV/dJxnUkT7kGdZcNnwKiaSjh3qpYQtgQ8TFRsJuKz8Hr1
ljAWOk7Lun1lxVoDF/CRdxC3FxZYuBExc2owVUnfXHhpSErDLuFkg8/tWvg9SII+
6bbWXg+Ricc9WY/bgBbOiv48Bmt1vMDx8nXX9B7gTw7xCzqOOmHYbYzp2uO/01y8
1vnyvm1av39WR71o52h2dvxwuiRMwd5j/OjN8eijjL8zP4TvLbW4wm3NkN6UYR+z
pE5in32qoXwaKBWSRWVafMrqpKH+C2bv0v1FerpEpc8349p8OXjEUOEufSd9ssA9
kxRQhBTHnzz6qv8RYioKT9SvD5YL/bdJHu5No955WST/uYxFhfh8U8QzWp/PXrW7
XGNPltLCP8qp/MbCVbmDlil64oCx1tNINkyB6n84fIHDvmAz3O90N87F/G3xa20Y
h5TtUI2fezdnigMlWOePJpQj70D+IZibp20yHYjm7TEfWDXap/akwGaol96rcV5K
+7TpjkLTHFTcoXxV2sXKIp0ZZC29HGVD7QPMijqQmpdAfpN7Xe7/bB63/LYauxJb
n2dOMoshK7Y0LbQRkOF3qQrYQW7JW63g3KZ0gImijcxomljx8xK8kHdh7lQK2Qjn
2PHGPrhgXzoo+Cxls3hGnPAA3k8alUN64MOLG2eL97JrRk9exNZzjPK+JRJXyPZ+
qNtlIdOtCNQrtnRar8c/h1TtUDcnhNcs+Ph6xgcenbCcnko6eJT38nqkKKo/R6Sp
8k1w5r5BzRnxbYigSvRQFdkI6n2qhNJQCVpkqgMOJXMdyNHz7eK8hqIidp9/VhyK
dwziTnyrm7+58HEwk7ZHqcWMbKGb2D3v806vs+Wj2OFNVadN+u8n4MeIEDabXHZa
/0LBmYOAAy4YLUHmS6m2eoA3dRwj/AInCyT2SuHFYM6As0u9nRwn7ql2l+1e1+9v
qqUULYf/5HxvtOUyIF3ZM1pG71pSmMSk7OQWWQ7qLVsVNx+UOH/h1bMYTANlgbs0
rBweEM5m4WVwfJ2rGqVDti/XYcW2/7cNIgGov2XXrKAFNVxspxpEkAlPF/4X/Erz
fkRnvFwtr9hv0LhM2MBV9OAYBHayNxNRZvBG7cOyPK8L9BvOvD/5fOdTb/QQ3v+T
neYaSkv0O5gcWOWkRF0Y/RtqjSdDO/YiAO1EGnsOl+lGAHg3FTqJx29gPuDXGpUR
coRJ36QJwC7mqroNiZODhE/pP0GIVpwBMdiefdmBQwBjM6xwAdWC1jvQkpHlf6vE
bvE+CgrJTLVJrv/p8V7Tdrwk2E4rFKlNXGB+eev0Fxll4T924Iz98XJ7PmGGFA0+
P6/nCyOQCPtNjfzsfLBS2LxdSIUZC0VWI3M9mcNravFLixrKvipT4IXSa08w0xCK
Sn23ejiKfOcZJXQZ0ryKcjEP3rsTrgCsKFpWwmF9Debn3KaYU0dNgKeyN3FVFqEJ
mURoKOum9RTXp7K8XMhAIVYDFyuT8bYuAygIvj2eV4F0CKCQYUPgzMi6XdZt2PKy
P3H9JGhvZ/r6UR4dkKQOwZe4ufG4+OFH9/7nGhl/P4Nz2PA9jriupp7qpiiJJ6ij
UfTXFiGtHFsj3n7BLBjAWId/EULdrNBoz+i6ZFPc8pdLtaO7OtJVsSg6UOUh3E36
TnYink2Xe2qGFhHhbPFuna1XCHDMYuG4qCIA09YRVqLo86COWuL6AYDJu0QBsVDA
WlZ6q95wLJ4BBrx7qZpur+pixuLYnBbIDFttWkTTWESctoQHj3dBx1bAuM4C8nVm
NDkpU5EXhkPhxXPYQ17Kkzw2pIlOTWrET7UTVbj406ZL0C+i1EaYQDGS0V36LlAl
aMLh+3tsaZ3W0KFbsDAzb65UGrlpLTAEdbhWgnEhyQeW4xVXysSZkqP+y2ystgeX
txD7PGWmi88etWAggd+VJGTAcBn/2mSEy5DIXtARh3JPRkyTTYmcSjjwWQPGIdCh
+klXyOlg2LYdDy6dDySzs4DeoMXxTrJwI2gCi/PMybG9uVOe8x/2qUNUK4cAv9Kt
12/buFZFY7oVtTyjNH+onmf+YzUpvv9f2I2wIjgONcF2+gjmQnTiYTGqYO1d5vLt
GNBbUEpJWq7wEVxno7fT+mVBl+1MmC52Xo9Gp2fBXcYZwecPbgfu3zHWTxwD0nqI
1tdmD4FtaPTgY3nWjPuMy1LyFQaTeSD4xSI8KE03R+JpPyQqNhErIK7IKqz5AE1j
i7fF5bVytYz5EcsUkfEc/bPfTun84eR81Ziyb0CP6HzGGrnAIk2tdwtoPl46/DC5
k9ANN1OtMBXmUq8paCzmZaDeoPvwp8eg1sFZkV+ynY+udtOOk7S9cxex600jJpMM
8CRiHGhljS0or5jh/w2lTVs4te4lqo6yPZtUkobVMo2g2HT1jI50clCnsOne7h6P
715ps2HRgI/Ljq5Gll6u2mA2TgFEp7xKiiLJ6CIAQw0KK049S3sawxVUy2ZnftCL
O/AI0mdyfYuCNNR2kzmAmVMayRTikWjYpPLfMbdBO4g9guBHh1GywNucj73c7myG
2fjPKd1UE9OhXF+Djox/D8D5fh/ZU4B2svZCU6Hg4p9RtJ9SRo8WrGHax3EakzMR
aDk8c69xh3F3+P5P1bq6Hgvilb3zcwDudyHkefKeySgGCZ/3RwaaZbrEFxHFIT+d
ve33rjq8qOghQbHG2wyV9V1sOfcKO1+5yvGTsxA5DmhcY7rQOlvaJkxf4CqTMm8u
lh+wo3bJFGhZ56L8L+S4XH+1TaMPZIel3OZ5MN6c8MR1GPmZJk1pQgS8hb1IS+eS
/recLfaAbAN/4wAicrOJwfSRdfpB5AeBpUUI5huHXJeMoPrTDVa7nDdKZQF6/zL5
ZdatYPtmFU9ON4+LHPjfloy+CnnREb1cvUI6TJomED6UfG2suEzeWwB6nibZArWH
BOPCwLX8s6RFDjpN0c0jZn7FnFJovPyGbdzQjeTXE3nHk3tZRdcc1q0YSH3iWPFv
Aqwn00SrXKoK3iB/LRgc03KtwrvW92f2Ug4nZcoW9a8DGgUDqtXchm1GhXs+bRTW
8oWBiDwzuMeO5PrBlisLopjACloV4RvUiZQfKN2fgEtgq8TpDg4+1iC5+Ufm3j55
4+pjLdQUSk+j13GrLa9i9ipk0jjxfUGHdpL4+TwZQO0QoMv8PaccG196Bg5kk3sH
uYrpNLShdLXYaRQXRKUM4fEdZ9Rm7hweyj/gS6DsQCJoWYzzfPZHHSrJycoEl285
CFj4fj9EMltggsmlq4SEA+L39mu5nrP2YRygsmWfUB9SWcKvVU0VRcKMSOxw0Gp5
XqqcQlHGzqyoZ4cYHWDf0I1c2CxXa9k9vUHHj68GO1h9uyWdX85GbVIL6waPWCzW
7j8Vpcged8Lgp7sMTtyTPRIojjuxC0C87su6vLSWitFhDyShaYSkk5QBgF2BPDA6
M1FGuyD04J2YvncKFg4k5ttcLsrPpKb6Q7Mr+pqL8pOMxBfMfdmg/BI2y1kfw/Lh
XmZLaaPgw7NbLbk62OAVwTQnb4gUW9lk3HVK6zTd13LzzElWIFux/8isDmLMHVHI
ngLHa52lGU7Rv00H1Lk5XfS/MqzBEmlKpLAj5I6nVEirzhhKhJcPJyuLT3m8PG5b
K9VD64zKxOCDlnTpwRnsnNJY+xzbJhCW4nDceHPWDCfwBfRvJkZbK95PMxLgVetS
dRpuR8dG8xRYS1CcWIhTa/biXzA1s+tNSCOrYsKjRBJHHi2GadoIH+xoe1kYX8Y8
H0VCZU4BsKBhFIz8N2E67SXoA9vhEllLPvI9k23hsLUMX9GWpYG0Y7gGezE9sIwI
RVa57YF1RfR59YKKZTTxSJUykgrZO2YyV1lJ10LpdTe0OxJI5hWi6aJRmUG1GJPM
u1m93UEuDIYC2ccV8wZhUIC/vNj7y4wTkVT4KWejGA9FUvli697SkFkGnUwtXCeY
C54pWV4ppJ1g0TsCDlKT8/ogfqZk8uBHRE5hUMB1WBA/x8IS/sh4l+pbGc2lvNgU
cTpf8DQKQ4ewhw8FysDoA7thGOaIua0jaCYEVmEdGnHWnCIDrZCspLHzDyryYHtK
2EDKCzXXFwnHdySRtQ+C3jh3dmBeWmRZM0Uu3ddxu7+V9goVhCvLAH+PqmzMF7uT
rpwiBnv8jqo/+4eg2voCgeaj7X25NigMo/483hVkkJV3LL4eVrccxKdFTqSOswaJ
VLzMRKmGwX8K6Wd1Mf85jIl208X1R4/veYq6e/dPvt2ZULk6Cfcc6c+RSY/nd8qL
zseOKb57VPDcDC1tTMPaCgqAhwau/+4L1eGMTkS1Bs2g8soEVfxR/L5pFvEtBOaY
woy3GjY4crk+t99bngE6jhkBw79aIBDVPQyFgMV/meKZiS4hqi2z/aobZc5ydlVZ
RqH1O8nTNzEI/5RS5jhxrcZdARpzaU+Sth5AkHAGsBbKHeXjWEeU5nFHhDZasr2Z
SGx7WFp189RbZ1yj4W+8bMOOvx+qIJzj7LsASyZtJwZuRT/uuTyRpIF7tAtcrgWU
oadnnz8z7BYjnme1wArt3s7mi30ywCQgHzb1bmBUSzopfhELFJJ8u7XScBYRctzM
oxE9Nw/Hn8vetshxwZEbrQbmBTw5uFYu7v3GeFyDxfwVGgRJFypf2tu6Q+b+1qA6
xpNA2EjW7f6d8/uSIhmh4j/7UCzutkcN93XboiFru4Sit7k2QqS2SDwnSBhMx+3T
x5FahhxgMbU6kczqK6b2/fK4k7ca9CO/9aHZrIdXWz6VtQOnYvzzeyQ08sIuwsDZ
K/e7ZOHh0XhR3iDk6CjO2DepPqPon04CnsHtQspNvDP4/GQvL2zGy1QH6HOUS8wJ
e/aeraymEt4phtawrDfoI0z4Ui0ks3x8IwSFHt3fp23hQyjkzHglAcHNSlsY6pOS
AaUerpHUxa4vTx1BuhopctVmorLnNiE2H10qtDsBDSHiiHAU3Lvhb47Rz5oot3IX
d7K7H6Hg1nS/N6Qw9FSGrBDCjvYbseQccp2NMVBqLw93k0rI7JDy2WQuG6KnH7Jv
ivR7kjuxPIKw/W7RZEzVPQXPAHclxppWCEmlMZTw1QjdfpnOI2YrJ7XwI8rdO+LZ
T8zeva3ivAFiv+RWtkTfbyZCJf2rJM3IMPBlnJveaYlFaMYhPwAY5oWedHii7wB1
wxNvVxwotQKGfZefjq0zeRv8yIDOFNbro0kF6sFfSBxkpF7mao0rncO6DsJFkbHQ
iLcNHhVKWqQPsVm0iLf6yZOMnvEXlHONz8KJpKag1n1kseUr6hAiRQjXahyDAOOQ
DvGtDAkp5Jl2Lq8f+R8LozoYkYE4focX9jza0yUMo0pkd4kdqb9B/IsCSEuqSUF6
o+L9U90SKuKjmY8Gj8AHSw7QxBYO02bGKyJvU1rHtPqK8BC00y/T3DYtnijP3FjK
QzB1MCxhiM2fqYBLJu38/1h7ozIiDawiY5rQ320tZAO+kDnBn0IQ9IgF1pCJSdVy
0CcJ/QgRkpXRV4mIpZBZR7B6aC4hRVT7eZwbXUyLslRAbds2vlXGhqxQn8iYTdbb
C8VV6rUmGNmNgOG+n4HTPjX1H90uHFoMJmq5Ua3RWbGLtjTW+xff7UW0OPadGGGq
d+HGMJk5+0kqzEldElbxg7CrCWByfgmFZ3HAuPRZ2RFQbsvIwhHA3OMyGOiR7MJV
oOeso+WLRZllv1Ib9GOwj20ooQIVXHuuO0ZXl2A7M05QdWeRYWpKEPt+hGQYCmnf
YHWk3UeovLtdEoTbP6YnxlaD8Jn9x1ku8osyUtv4yski9rV7gTiwvzNRoiaczzDA
iXFlXoWq3MxIisuW2OhfvSJ0SptKHJpxiMC5CjeVIdw+jtaO7AUae2GXReZv+gks
YNKT3fY6e8YEbcmxx224e9//ibq0husdVyifKmsw/kYkI4H2biSIC9czuDqnvmIs
PDGPLA32td4qRWTC1YAHEYfhCP2HxnTuhwsepoyAL7u6fQzWfpveVQEB09vSSZY+
sc0X2BekgDQGWxosq2f8HWSIAHWqcqKQSsRX4G7hEE+HnR8v9v7ZNoCeHkj8V0Zz
7zHePfyDCLxz8KKf+Da5vrJIrAYZIrZvSoey03ce3Ar+Tn/Tup+V0kPkh6W7XB2Z
2Z5eVVa1VuJvVUn6gr487IuCcB+Dtv+wdxLFFdAUl6OhOdNrOPCOWkJw0mOuV8qj
HxScatajild2zQEPZGbu1GBJFmOA1788Pmorhe6+pLdwg824vYIFE38UKEKUyA8K
aCaOoGN1yTMFcXJLSBs6znz9bbtBjrv0B31CoOFkoTRe5RblgdINZ6uIb29Tvb8g
hLzYQFLK8JV2TkEWi5ePq2n2snWbKp/WZT3jHYJAtgh8msUJcnlHeUi4WdImnmcX
MG3IJepqATZo79qxRIJ6nIvTS7iB+jVI7PN8CQQU81ahlL11v30jdGo1lJ2KN2n7
tg10ynI1pzhQ0xzMkZASWV3MMOxDNp68AL/FbdBeQ4CSZQWmUh3QWqteJzwZXoCu
lGQFGBTSK8TBxUkNT14v4PQoWO/Pt+foUc/wKT64kLLWjiwGyE6HZ6UeqwRXk1uN
kxRiyP8nPSG8jW/CzwIzT5jpnZw1zS8DPiD1HKG3Roip9UyF0/E4FbPEWk+Y4rL4
QpvfGWJnk2C/YFAiDT4e1P0HKcLbyal43yUIaZ52D0lHDxpm9rkQiHEvtstVp3X2
PlC5oW5cfqrkUAnQUUgdGHtm2Q5OubVfjoyHznupjhGF2nllx4IeC3qBX5I7iLLh
DnKxQWZxNK/mF+mXnBtOLHN+GqMAwVOqgxGdc9KANoiHXyKbi82JBzboZaqlL8Bf
asJL+QgqQ7YPc+h8UOcNcPulJJPijZE88OUCP22N9JEkiE8Pey7Rs9dRJKPRRjdN
xxbDTkKmjC2zdrHNQXtvsuyesAy7yZnZktAgdxdKI3aOh9L+Z3ZW+f40YL0hOKxS
Cipx/ZpCohi9tCHB7uTxBlD+cIHPLcwMyBjHYFTc2Ra/Pqy4RPp/irp1f2dcZvxM
N59Cbb8gm3QjAvlZUp/bTx+3Jfa1/XrrAXAfVGF3zDAinR3kgoFsXyMfFqHFK/nS
sQ60RBxDld/UHxBAomk8go/9Xgyf+VJGV1pakU3bzkvp5lyRQoFPbZAuDtNv0BxF
IacAKC8/XpwDvOf6KMFVMk+d1W+lx0Lmhaj1vx5VWXQGo3VcwJT4w60m3R2bEzIK
kEJ0ghJ31McGDlnRHUb2Jnlx78KmQ24exvfmqjPhaEi/viiI9h1mBItHWWl2vCD1
C3oDFldaS0TQP3aSgwW6sLC/gmmKDz4f7DV34H+Yz/qf8E9MhyZHfOH/Yjc3SFtW
NXpqglEsYep+L+sthSuHL+m6aPSZ0MPPayTg9mC7POxOslihn/HiN/tjOgiNXhmz
sfmauu/rmVq/mQe7TDpFM/lrnbjiM0c/WXYC+al+JITtZinSQvvAQ4GKr0Vdevk3
z88se2u7ZGehIxvCnP9EwI9VJIB7ifCgSBSDRl0knYPUj00SuYoenovB203awF7S
jBom4AusZpJ8RbLliB1szfzJnMhu2OVyg22/L7GGfTqZEXvV1dJQaVvKZTUcqbBG
HDCUJzo9tfQ/Op1iHbHaHShwHbM9MJxdXvcYHzF5ODgcddYE7SvlMbTf7oCsfqol
pIkSSnQPvDtoiWvzmFBJ2L8AMrmESRgLgJRfpbaTuWCovl72rO/qJkHd3wMj4v/Q
ODNHy8Ytd/lS9MHb7J52+eYF7oqu7KxVDvBi+0/8pXWe3IHj8f5E7ekVQUwzYnHC
9uSOESlmiYj8ElSTOg5irgc3T/v40NLtZsJ7wgJN7QzBekggKG96t72A1PVSuyY4
qZ7wRscamltO4h46koEVBF0kq05tAMyPUFTe7Y2cEgF8XnOQpYpeiRCBb+pFUh8o
m2DlgHq8deJ65eWeeGJASyMn9Znhc5+0OzPWqlC50SIDO10hUO9KBpWmL8icqARV
qQiEUqbVw6jwN+tvP8HO8nMGoEyVRf03LuYWxGuJjQ49sEUM8BKIxJfc4RZfWdkU
VzLM2mlCjJ/8SDhQJcEQgM8Df7Cj1HLztgGCvj4rqctEB8VU+P7K3wDikiX6cBiZ
+NdZlgVa49CHlauBiesOZvynqlTEvPH7IL+WfyOCNAiJq97N5yv+CYQbsdTo2sPV
f9nHsDDTTkGMJQs7UpOfmcGeycjKOLh6jQK+UUZsF77od+ft7B+yIyK5Amskuk+A
UcZRnFPb977cbz/lk6EqAjL1EJ4GBVZAP7LA1VF3v+0LPEF8JcpsnlVIWcG/duZ1
enrxfQ3Qs1Lwt3C0XmZRLIQrWhhhXTTehnG2rpyTfTPCG0OO8XhM0ZO1I93URSAh
iN36fmerISZ8xzcu8qkKaQtsLv3OZw2jYeB/vLSbPZQ8sy3Db99Fq8O5iS9gl7JP
Ye4ZEODX0N0qThLUCX8qS6CIz/tfV2DjZ+T2x2rZqCAlv2ubgP8fFNIQkWnFKm0y
VyJ7kGiHSw7P++Yz4auMhR01iBN2+kOS0CqF75dlA/2hVYvQCuLd4audf/gaPL6a
IRJ42D+ngY1d9fDty+4swokRHnhN6qMIo9F3NxxS+u1JTGFplXFLMNaI1FnbC4FV
U3DSMRfKCuD/VYMOQa2zvBo1tKR2XejDir+7GFtA1SJWyUuHk3QFkl2GN6De4t81
LsuM59oUGuCSikc6SfQhMQ+XhhqZYgM5hiROlg0Gq3oVpy7qGDnKIMb+eNj7ju+W
KHPV1wgXV6Ae/XrPeE+lbghvogbT52fWKWjowElPMfxolSRGw1sHevKcoSg5Hgal
rrVLF5QPulf5w92CHm2Cb410L+9RkACE1Jw0YutUis5SxeAp33Ui0OaGn7VFNJeo
B/BgqjNkXPjFJju6Ru8bpLglXuyN4X1dKV1zwFuGA0hQ1e6aTf5V+V3hJLTpzULM
9QEwLckWoKTZGdA3m43msoy1O6VwxBrHZGDtLfWSomoXa6hyc+5MWPtkNKMDksFg
zclNVqfRuNqew29a8aq43ygdOusQH5DD1GMfRGAFG8vGDPDWA8hg7e6xjKAqg97+
GwcCyy3MSA88RVdE74q1BFhdm2qo59jEtsoAFrYGTMr9Ii0Rffa/CeIt/sDIrfg9
C1hk6N+5kZk7Gz7kHQuW+0y/9HGJw9+k6Ngs3XQ/XdbKF73B6PZBv/alywDF5Nsq
Ps55/2h+ZM56SMU+fVrIpCKrbWz6TX5DUnbR5TRieJvxUjwe6eKWCRwp2eiFPoqg
AonCk4GJjBd4pavdGqVGePHL6Ystv/CQgkWfPOSkuj/hDiZZp5uBqB3X4BG9VPFn
QQB9maFPJypz1pGzR32Fx/CwLwb3mH9OZWbKmbet8aDPWvx4zXuBKvGlgStg/iv7
Z4KtyWEgHA76FuYGdUS0sZcSTpEdiTkdSVGuBtBPXZsIGGQgiF59oPTDSmKNR2YC
Prv2jYgTz9XD92q+CAtJ1QzcKuhIfablU9vRBDw8DJa31xoc8RDNSFek9YfxQy9R
Gpugb9+iczdyHyM1sCmi3pHPFsU0slJUE8ESanhZRHvMa13aA0h5xJCNRzxzhcIw
PIYg77IX8hjLeCwzbGjQ8xglSyjAxGnubpcVWAtVHP8W2T/twd1mXv72lObnvdIo
4OaLuHYQhqPsUv0/XdPjC6UjGhWbvqMX2Bi+whyrYQcw00FeKimfrDr7nXqGoTPg
AxtGk09+ImhzVkErrY6wEytJ66aM0uyEc5clA2WYw3dHOCNMrM13ItLhrEEqntAI
M16dPFbK0l2p8Av4+UgYs0OXTr5RUp3RQQ6rgDgxcAzM1m6aXSm5oz0meaOcjlgD
FLy+DqUfi7aNO5qJYG6ElMut/QkmNV5ss3yc3ChKUcIomiQlcZ/m32NRih13LQU9
4aT1GCWyaL6eOC+FWcei3dgYVWjrGRxZP0oU/MloejFL4pRktS8CaOk4xlDt3fJP
s+6L9jIWNUdtN9vGlKBMX7Tbv2Z6TP2rNl+FqwbF5uJe0PgpZ8AySGbNhJ4TkKkt
yd+TVlUzDMo4QnuUss6R1hdfuysm+OssH8AXhpPxLooWoVksL6bOmsQRV9APK6ue
9ZTQnUm00Zan6hmP/ST9gRXEHlO3TDUHO8ct/E8AQKBx+/hVRIzTRnkxHWMOOr5A
o2xmZMrOV4+BkqgtkoDgB/UKzBVhbN3plhFf0VioVO8CgyAbWAp5X0Ot1XBuahXE
hIlR3KT+XMluMuM85yWJ5bTFVxYjd2WuqhDFSNaSN5loMEvf08qZgBqc/GEQOG/x
IgC7Fl8uKjV65Rscb3P9hD0s7lNYEGVb+WaaFwE6pVDizy/ukJY0qSQWMUYexmqw
EmXhuXwfxvS/jajy/ZIhKG3a6KisLes1wG8W1WSsmsrx6gHrJRbPfewX5vIhntxS
GjYjG/UhMnnIsLtTbiG3yK6f0hUFHEisXwDcUY1fv6vBGiwKQwclG1dfWtbbImkS
/7//dEPWimolc5ClhHpcZ6osmh/vwiio9tFB9N8zLPHYCLZnujsym0qpx2zS169u
2VswQ/JGY/KSQ4PNtxTf9aBDNJIeLxNKzVAWkjLr7paHLSdIS+urBEg+QyHQKSM1
M3hruD5aNY/9ZOimxv+/nJXPMx5H/e5jbpYra2vW3MhqY45hCqVnokBv55c7iJ87
zZPXKn2gEMLWYBze5n1/JDEb1CNEYqWEz5ywP7D/d51VLdRk9GOSUc6fJbKdVLnp
l14aeUUQhizn4/QSVLJv8OUKiMp/9TH1UgKLbFxNa5yUWVD+H3qG6KSsP+3kcyfZ
UtWFKsllC7ntyxj2ULAUzd1yTBepNmD5EJ4cpaAy9vYULF13uYKQ0rnkxRhaVZBc
2rag2n2jf5OhlwSE74BIaI8+RaX8b9HSqmaBJZYwHDeBo9lbexEIm9e+dwlQo8AV
mgorG7zlefdaCUZwbQEZRpB46WioGzbAkeCKYj7wpa5B0pViLFdtaPWzr9V3kOe0
qbKVXmF2/JcVek19p6WPLY5AYsQBXSdZ8f6skJ354HtqogmbnDnKjyLXsizBKvWA
10/n6ny4gfdvUy6ZRCH7kpa/KHmt1ur9VfAMA66HE80as5bjOU5UandnDOZFsJQ7
LXjAX/KNxTx8Fz66UlvoAuIJzRINpOJ31E22dMFybGzjSS1tXNn6TEEu4nM7+t78
YI4o5fwiHy/1nXbherJKqU6AVyLD0x5MFxuzkjC4aohXpvdtfy6lDg4HIaWnkXo3
dL0BpKUDBrU76fZphq0xF8kuJKp1+tXYsl6PjSzK5GcB2MpA8wWFFc9S4q6oHYVx
d8B97LXWJwcxtwW3CUpfDuVlpZC0MGWxjP7uKNnXdLHlfYEPK/BHVaQGPJcQ94uA
gx+ir5cKHKp35ON1L2UfLRoUZ1MI6Z9cms7CiSPXpiBGr3ngyoqKQ0VqE6AxhNPc
kZWi7d93h8gQprOEpGzHhFyTZSBi97cnWBCOGBOn3PW+GIo5+M8u7uZ3MwvxDBf1
Qrccp4PHedCGg1mbkgiHY+9FcCQWwhAlPtyFqJ/SM1d2G8CPMTaU1ghY5vBPNKzx
sL9M6rd3Ium8tcqouMgUqAduz1Je7UDTXhW4tHd2pPk32FYVbsiVxth//o7YjtWF
X1tcGAoqu6JvlYXmynxNuMDlpEkUlCm0SU2G+jHHn8paYvaPz5BC/7/USSJbouy5
rvhoO/EONcHM6j/UGVwA/mhMlxZ7RjT2iDh2UbIjA53U8Bs8t/hPRHrnp+bAyf5N
P8vOKPU/nHAnrChWnoMCxi1WPVFnFcRoud5N8DIn6qAQN97/yrYI5/IQJmaJ5CQP
ISWE46obtnQ4lLBQCq/pgiQysEDhp0KrzyG5rqlH2PMBnqeujTGWQb+n7KuB+SWY
wzmvXuH8zqFOmVHB2Ue4lCxqkdkbjsCqLfxXsgC7ihqYdrme9dIsBjxSgVV7pnL3
l+iWrkBkFwAqyA8h2dWBM21am3GMZcXcWJ94rDtkRb8bpQ0w+hdQxpJkvYTZ7cA9
ebEOiOfRvgyFTGeBLOqCFG8jkKBqQOAT98bb28ZFxYKt+5PF/XDnra/v3Yd03rcQ
yXs5nvSwnjgw6QnODKYH8LRhu4MZ4ukrr7kQxYNx48+pw5DpN/ZPPFHD/ByaEfDw
56hC8wNokqfKTQrSYePtjA71I93fYgLTl8rjNWW/686rkF25CRzlQLzFTlEOLmOg
i1XofvoOwjqjC27ERyvmk8woXF5tF1Am6pR5dpLAdCYCke/b0DkjcH9LxLbvQw1s
pzgXqZlrfkKW5h0EUGDBdwzEEqhsDpVR+50BmFUB/oIGfKD9rOvesE8/q3WCtgwg
OEWcxnpikATQLWeBEJ4++cSCtUU1iV2wDer3XZpXo7Agn++EVmP0ePSpIjCEtP30
KpkpEmi2W9s8tGi5QIbtTGO5/TKLhGISRJ0XF5L3q4M8k60yktii9uJZBG2hRO4W
UPUJgzUY46I8snvPzmdgkw/6IPBMMdvdpuYjfnnryXl6Rassttc/jKQQDonp/42B
eVZfX65NKLs8sBRGMLf6PA+4dS3FlUI33EVv1lHjD5vzZHNL8qQsDGV1xiaTOqxW
3fXnsCEj6/sZJlANnSDE0HYT4rflqIxaVw5CdPYJIH5ThFyV9oFUSWUFvOl9V/8C
jJ/0rXdhwzjIxMlmuwiHeDRR2kbmdIk7asE4GlDz2BYb5jKITUoZ6RUm6/XIvGUb
p01hL6XwQLrSSRB1D77jvDsqWgVbQ2iCDHDyrr1Zv88kcz35aOkhiX7VPBcwdmza
gyhVo+ESODl0ZDlVcafov4HVdlq/ZgZwOrNFy2G7Xj/OnwGCnnO0Zgw8WwV0PauD
QyOvLBHqzBTSjed0tnVl4hqiJeWKCnz2ead265a1v9nBA/Whe5xbP+UieEV5oDm8
gf6k5CgmN5mUxd2Y+A3Py1IahSKrJt/SBomFiQGbVpe3q8uI+P3PAPlxIR/v4JJE
Igrg8BNYt+GT06CDKoJmH6ofpStKQAUmrpvHrtsmCPcud3hYP4250h/wa+ztpbwN
jG5GCbVYucXz7BKcrw6DzrMgxgMACXEiRcDyxB3iidDeeUezWOIj9BngxowQhp/r
/u/1bg4bcAYulp2fOhhEGljzgrTfUj51S7VmszETVBy4fMDZNa/Y+qUfaz95gLJh
Yvspr4H6sP30U0MMRdS/LJJkbzRbwlQ/t+notG7k6+0lrG3yFZArpEqRDUWRgoNm
tm1p3yphBJegqGuVdQoU/mEpNP8GQBOTb5s8c9c68StnLNvuI9EGgIo0q0NMe796
Pox7YMSqaWDg10oRyZdHeqvJ1azgqz6RUhCW0TKSwRL+B9BcL5SZl0GGYNIO5/Wa
Lilvd84Mosf0HSRvHfvaoWWFoE/50lzBdvonLJeQkp2JxJI1UcBQW3kCGpzOxfPG
Ff/i1bcQPLEE6By7u0xmxpoRoPU6tyZBUfyRdatwG72m7IZS23KWVEr+LSH6xBnz
RmVUvFL0cGNM2ERi/n1/6zOMshPNzvxh8sq/oCH3pmNuXROl4YnorSFWCaUcVo0i
huBSYXahXcz38PFgoR4rU0hkh/yFapuUs7S0DGySvqBgGTmxT3jMmvKNagmSazlu
2fTRC+y4HFsTKgjmaBDihejkv7OX5TSKhrpUFvIsD90d1KhRWNIjFFBeK7zf14ls
XLf8TAmDgB8NjwH7lgLqotUN8ek/P410bGux/2u/5y6wWPN1VgspoFQ7BlDqG19+
k0z+tgZDiO3RBYKICJj/+ZhpiZR7rxkHhG+8+k6eIcYYwdb/RZWDfqF1y0az/oY4
2yX28lhHmJEo1+4yOHyvrgme+Ha8gpacpEWoJD8VycAALh2Be0QJGq7Y29VSpjiW
hxz8tNecsb8iV1+iIsBPEZEaaqjDwxmXSVmGTclI64syIe060C2/wtj6P8i47xfs
GXiNvhuX3upjcr7Evjluk915hG99a4FkSVbAv6BUi1EbHMxwyEcrqAtw1Sb1o7Nw
z1qBYIWfGMf2IZqbKCh0rOkCEGk9rxsztMuopuSJenDhvUcl/AxpwPpAIaFdULT8
uqmB3DxqjDD/JfwPhgi6b9boxYCOoiPjlFBKf1vbowSG6ZtrSurV/GuCwmd5jfLD
dRd9Rw3rMML4LEbHcmiMsDN0jWqjn93XRWsffCJjKdhR3qWhDA4e8vWa49gvyGeS
l0g4A051CYYBfkpxJ4iuG/+0s40tVTCsdJenVKCPvU7CLJzTQy1EEutQ7BmeH2gr
6QO8Zqh4n11B7jDAJ6gK/Y5YjkoJXqpDTYQCYqlC7dgxxQ+inKi7uEnVQkW/idua
RFqRXc2Ddy6F9g+2N+Y2qac0nrNYc6kGjFgK8JdCGZkPhxaVZEmP/vct80BgoqSH
KXOP3NfkExWcxgcEUzIeaJCVDrTtPlGbxisTGX/aLHitt40duBXUgMgoiKXc4X+l
TQHpQHDwnRmj7VCZB2PacZ6WaZR0ebzXqJ2YpEWfkfnT7fQZa8qfrI8m4gcJvHvN
sf9Xn/if0LuzN90vDvVBRnf5WH4hgjP69cFQoOfdL741YWtXdnxw0CC4TuxrAO5G
rgFlILaTB6Yt6PBhaFZdJCkkguZ5hEfotucCfUYyBDMbQ3Af2V8n85YQmyZtLTXv
Ws1ml6/aOQwFVIkdjjJY6LFl2WbWROIu3+8EOMixOE4BRmbSXxiAkkCIijg7n8Py
K3IWCE7j/GWCDP9Z9Y9+0C1px6LEzQtH1MnCHZMHtxYhui2HdLgbNBMrLlrmREmL
EAZjvub36s7OrWYdA7H/UU4wsq0xgSbzpBMCU67e8ZqEMW+sQEk1osHn5zMqk50Y
DyX8+NWwLEnqDIgV3102S8LcwDOI00pXKwJuYnpT16n7bYCvzC+14b6T2nZN4J/i
we8eUFd1QiFp9+DziY2vTrI4smX+0SGcJXCGmGn1A/sSMc6M5ioauCaAQdcBxorM
T4qE4BEDVP1K6F/+uV8jQGPctRm83y2OA+L9VCTR1KCMa42evTNjPydmW8JU2WdA
yJHGp83GGVQPjT7i+6uB38DGb0nCzalyE+mCI3/MU2KyW3dF+C5PR57Erw8MWfzW
XgfgxDVLX1IsDvYBIpCkjhzNV2BfImxdLty+ie9LxNb4E2rPoxlWOwdpUbg+qrOD
nAWjI9WoM5a2yXKPLIPAZEaF4qBDmvCKcNpL1t+5FKCvsT/0v3TpVlgML1KHskYx
7svQCFcXSonBPZMLkkQO8l1Y+myQERKaP/xnR+2GYmcj7GxXyMGZJ8YTs6XdJVWf
hlE4PQO/h+6pDs1zncEMbYg6q6aXKxXUckVWMJPbyJeazzMMi40DXY78g6BjVpGx
FCAPOUd7IOt2yK8jEUFDN/3dFng8MOi6DipL7/1B6TeT8ecoIZAfRoUCGV7LZD9Z
rigYnyyfISHrmTmd9X6aCSoAz3Ybz0tne46tsIjXuQWgrEgg5HIq+B/jST/DUcTV
fCiilZiajp/Yxe/INrs3sQypBGkXkfrU5ApJJb6LdqWVmiE0JNT0IQzzVnHyRLKB
90s27pOR/NzZ9GZ4cMTZin3s2TCPlvD+34WXX4rqHj/mw/tHwlHA78ZmXpacwqeP
nzLS8o958HQv5nEELz1UlP4o+BVc2U7ZECzsbfX60ZdXHPY/fQXmgYwl6vGs86FU
4MIVSQo75qWkboR7pgmqgu06icqB3vHB+FZ0mCGn+g3hEs/r1a5o1IN0RA34l+9X
AD833RpEdsZ6NcEf5wqV9KMenPWxMpv/ZnOyQbrsldy59fQeljV/0usMJRlgbUFK
RcExlseQYwMNm1fQPEFZfmCxADZYQqDXpt/3Y7iKlOZk6A9DdszN7QdJVTfQifNT
2nZ4IY79OAg8vKPmn8qLp7faubsHt9fBn+7W1GI3RhbPQqpMQeA7l7ZxzRBoMVL1
M9XPI+oyUisQxy0NbMcBJMeqOadx/gyTFiMfmnUcKwHFtIeJVkfLQLiTYxDOUcWk
VcZc32B67ROJxn1RKCHzTCc5UlfjyTZ7Y7rwSiofZrqKTDw+SQ+DZ9j/ZesEmvDm
UWF0z252JYhlkIimjen29IxOnXiV8pHiHnhAJqVsnW0JyLuMQCfUUwzyRURsGb6t
hKNb1X3zJ3JDqtT+WfKcjQifbg7qsynw29HDe7WH6V5qOEE0ahkKDCC1HvZn2+rj
xMQmotPe+a6N3R064/QCOaA+amGPcfkU/+zGbthqGs9XH7cQ2vIXRcXzvBrR2iNL
xj6LpyB6Rf/XfLgk6hsqJZuf+ZQbOMbaigB1NGQchpKzESLWSW80+QJPszRc5Muy
4l5gUorkAOLHgdhT4flkaED0OrmrbSRgN50Q/5cE57YboYkE+8BUcqD7XilrLPh5
5mcI9cp+0Zk30nkiQubcQezk7sHi2XE1U+lKDr5Su7ULP0Td9QVleYfmP+/9kGWR
JK4FJkie3YFJjUrxvDD/OAnQfED/l2eGJBaitc7hCdmJzZ4XbSW9eD129MkAa+JJ
F3UcVV7lKU4YbekRyQdcQC26Tbd+Ewsa6GHbg1nVee6xuPbrv+TO8w2SCDoo/AM4
qG6MdJQ511mnDBzvSTxbEO/Hh+slnd2wIzYQ4Rk3vyWMJikm+j1GaMxb9s44muFb
tB6h2nFHQex0jdkmoxo+BasXmgXrBjqWtTrtcbMtLgGX3+NCe6MXrrJ+yZoOT7Ix
b8BYDEZhGcD0EAiuvqW9miibnGcWKVihVy52vPHsCs62ORSI/ubJ2E6LrFjOJHx4
ITxFg2VirHDc2PZ+dvqxHCLOrzQMXnVuCMfcYufIKwi6X9CZFrCiRuWQObRF6KsL
BSCe+OoKp9lP5Bmpi1SdEe/VQt/dP1J+Vt8XFm70mJIUXJYRkM11vwrO00/Dd3fj
PiM+t+jHdkF4GyxvrB4vxp/XoPvfItlkf6XiwKtjgzX4wHYcHbSdJCVSYpJMMOJc
gv5tziBtp0UlQczoInadMNfCNa2vRueqAgsSBwk5VTm+6jAbpbdsOffFlVhJjwIX
NflGJHwp6LGOaRGuoqF84gaap3W1OILL9s7M09jxCskskLa5irMEWpnR+wFAJnyb
h+h4iFDs/FbzYzN/mH++ddBEft83JF1sZH7KtoEpqZUxqD8pxQtoxZhvMCmBJ4kZ
tE02xEZc7CKxGPv+iRFSTXhb3xZkafp3ue+oRvXgX3x07KHBKqURMHqPeyemEWhy
uonlWy+CzBxaN3MYT9tPncKs+pJlifUdW+aiwg9Ejf3kGVsdG1UaxHI0j84Q3pvr
tvC7q1Dpq+JxR5jZY8DTNl9+qaxgaamBeKfqOEXdNBfHVCgvkwOK+5ZdkYa/zw9b
Uhdt4xE+wwnrBDXlKPKrDTK3s8M2krQnQpKGXU43OyvDbOuBBiyQNRZN0Wk+xtOr
fGh6gMpe8Z0guzxWZq8M65fe7zu744ivG+JOaZZ/C//FReHnpuARmmOXjCzs8PZr
yYPO8iGA2y9Sp2ZPjgGk+SXah/q/ceFyewvU8qgs9ItZ3PlbX6ryZp72FcaPIhah
bg/xpdoPnuOlrKjKnSOA6n1Ir6orTTrS+9gQwTcJAsqA01tpAeHGKuJjzk+5iBjU
sVywzufvIJWzpNqKiSCjpaWlLLYxE2Sy2XLrxXXNjOYbv1ziM8pJbcrn6WnGlKRP
EkhDvX1xFBWoCAUlIrbHZgVRRprDLMIWOEgoRPfuFZ3UcaSP8SCfN/JYjPjQRBah
r2G2rrUScxgAiPVzsXGZ3k9M4k69q3+fSOCim15YnxmVFvTuUXsssK5vzSQs8W1V
dvSrMub4qEgdrsvIQl9PWrIP5d4hCP30eHW9olRbMHJA7aEKldUqMvtdBR6DE3VX
nj/eoUMjVnHz2lLVeT6tJy662jm7dNYMJTXzAYF3R17MQjtcHdGnK64dBfwCKZg2
/lj2toAMZ6Ze0yGRJNILF6GvKrFdghW2lIO8qXT8GZzN0k2m0wvbrPhS0hVboPx3
Mp65k9MbVJp6pRgLvAPsG/ZHiKKZzEJ3sFzwqB2ZvT5D5GGpPdha/QS01hbMdzME
JYuabS3eGSNr1nNCJ9Fmzyx+ft5tSVKy5xADYMpKIkuYtGDcRPdp9hoQiTaiIE4K
UWof3PPFyYI8quR4QkjLHMO1Erp5zwHQjGdyLga/kIEMyORjyizaW1AT7jgTPBtE
Ym4cwVMNKs7osCmbgf72v9WfALiYUAPRyoCLq2QWrnMXcWEHidIL5MQrWS4mAkyT
3iGEXyGlJ4pS54D09R0sEVlQJPeCJ6mAU6JbeZGehI0bu/1JB+vBei4jZK/pUYMP
cjx56geeWPvhCswSjRFOSAh+UM7lApf9evjTRtbZkS/QVzOEveUf9awG7yxWj1DP
VcQqB4Daq9jVZLsizmzlNU29tbJogVONueV2v2UixfZyFPeu6RAfa9N0x93xKFZm
j8hm+VLkjJ/4wWMdtETa7LEVj4xtmmwrVj/cezez3mAF7eEQEU43WccWJuOIk3qx
B0iewUV1kML0H9MgNcGQw/bQC20rd5yRHRvy7+QzAN1nA+WyPepCA1PUZIiZp9qn
MG1iH7vfZaclSp3pncaynYV/Lg+9NQMFuNiZkuJfLo/30T3tEbWt+hsnuqTChx+m
POMRz94XrE8mX6dbKO3+tzKkTT188yb6NbSYoMUdRMrSe1qtF8Ys8OGiRKDjfA+q
WVdKPQYkB00ftkMPAiqZhxerOySQOzgasOCf96z6AvdM+PnpY8GFdeA7JezM+d0X
2tF0c7gsZzmIYKVjHtLWThTQ/VPzH7N/AGkwzPgJG3vpvfxDzE59ZWtB86sNkOGK
wYg5QmUPkLAxQi3HKyF1b9bAi25ebvcOf0f+iOfP992ox9e/o1vQmMiioqnjJxaC
qitHZT81BGJviEfpzzX741YDMYbgzLzLKeI0kkEuDLRuJvs37R+lhIXoMqbBvl6A
TbUtuv871izecSUocDMPdNFLXxBtKfKL4gcV0300LQtsGhlY4uU03VcYkajsyNnO
PVW9voSfLpq9A+mbqawpPSB1jCP+yeWX8Vd84iMU/f8bjR4yuJIHmmNpOwwJSnHk
ddElTMG6QJrtJRG3WMRR4Rb4f11u9nJoYCvBAitJ22FQsY6mshmqCuUgz+NSRUwZ
jlc47kQ43ZYM+KhzqWwW1J50MGfHrZADTXPwW7Z46hOfHp/fv+vJvcyMYOvya4cb
YD5B0LCmvVoERSjgBZB2V3JWb/0CjxqCM5/mrPrjZ91c3Z9BVQ5a2esSEyS3Hbp2
g2IIDt9UsMRGN6eODV4WN3BizRcggqA5Pc+k4dvbtjTRJ7t2n1W5J2TKB4apMMui
j239MK7A8MGnbXMcjg1EWC3ScyfuBTUBte2v24tmcGmgsv/Eusw3t5HljCVNf3+L
13DqICxgdOIyTBKZG/ZYGBTnNgmShegSwoGBx30WRhOSsILWwO7KG2TnKcpEBheO
x+qd9dazpRY5V8NTBaLHKdo8nWm+byEMlAadypD4mx3JGH5rxerIZb6G1TeK4B4r
/YKfZKVBMFBqEg0R6LoED6q45UAenu3F0bVRRC7b8HdzSdnYU+d9CE2E1joG9BeI
3Ai3Yp3XdFS3OEMiZpqgfFWy8CJqPUS8d+Ryc/kbbnNJGhB72PONg9T9D2iqE3DX
m5Ei2URPnh0Zg6zR2VI7U1Nl7D9J7y9GEK81qepk1b+Ia3FQ7dTWencmtYDHOQfp
iugGU4Iozh62/2qFuiiHDgMKHJ0Uf/Wm5XhP75srSw/3JE7bQpGcU6TMnJa7ELPZ
Ijby3FRLhTqFHdtwGHMznoQt88Sd3sukdnTtHCLyHir9Z7jeqELG9p9Z687E9tOi
i6/8BFkiucygBg3tdstEdS0c86czkwbK/pbxTePYtGq5Dltd0XubEbcrIu5RPf+R
qgPPqSWIfY/dIdBXevwAEnMLLsn5BsaNMEkZmpmxfI1okGcuw/d0EcDE+315ftx0
YoSA82FH1CC5k91I6/cUzTyWPvy4dK8w2+3R6FjhZt0HdXPx3mySaojDuEg6ZAAa
/ad9FumhCGzAq153Pe/IaxJCOBy+oMc2rerUkNYMowVD2oM6j2ya10S28Fkv+7cq
M1uCZArrBZil6ThvYvwJiscDi6yucVt42Or4J0/JQyxycxd+YlWvLNAZJ+RPab+B
x+CNOjKHqCyXVHHCGYWAdLnn4g33DAccAyZQ8epUaDuQZImXUC/FkLAiFHaQxrkW
xPFZF8GJwCMY8XRBL+dwvAYjSYaaVrsGyfM78IENiDSJaTCsO1Rclmf6d7KyToTb
5542SHO5eJOWYIx8FGcMco/6Hn81USZyyac86Ot83meYGK5cqb3IEJuKNqgettXD
/IgOfwojMgQc19EwLbYKmgBpweKngJFsZyPn4Elrd6rEiAO8E56eNG0gcANPr+vj
WSQQoU7HDjyC/BcJMCf4bhGUafSpeAvxlYiUxpQddktlbOT6FAtpQHJMy37P90ZE
NpEnNuXIYj1MiVEoH5QJ5zIn+6ewBoZZSMoaFO//ISubBM/Toh30IPbbgtOEWT0j
5W7yAeAveF6V4AnVsRPu2hXA92GA98cypPSvgacD3zHkGK8qfKnpA3Quh6FJ43oI
tGnp/rlUfi5UyiXjOtVSnh0Dazc2uaD0Um+567cT+BQMGqn16xYuirl/LvCOQzrM
xjGdYy/c1CzFYZfSRm79T37ZD1E1EUhyH9eItcd3kWv7h7dkHHh0jeMBP8/NpCct
EqcNaKVxnfzZOaK+qiHCUAclrm21+YG90MtnxYJCQ1/IQqCAfBrHCm//laB2iDPV
u/cr+tpU02EJqPNTcCesLTPtdz5KZMA2trl7x6jbtRQ35tHu+DXS/LOBslpF4ns1
yerpGruo/jSLIJrZaXgJXXH7RcdqPhvnNXhpf01QBX5aqaJLBVjvASP90umDfzE8
xo7AqO1aXYRe7rRInIrgxGITB/ZS5+annI5OZQJODNNIPz6lzGX97QOQn9U95v50
iSOt+WFekVhe5xvxQEAj4a0JNaimqrIT3sVwZwk8vS9fiXhu1MuYv2H7ARAgcEj0
NRUwUJHOvz9cDq7oWd2iQiCCoPifJpUqU/pQ6uPoA6HVY+dReYEewY+z5ni6/jSi
6aa8gUuYRfJDdbnWJL8qaDCB8p6jmRMItIy9JguLF03Z+1Wz6Y9GUplneyZ0NAtV
ed71gJ3gsI8sj/w3D0Dr6M2vWiLAC1fWMVp5kHUbsUCzentjMA5JNW89dbofDO38
gczuuor6Ap3z6y9pGsQ6hLdTv3oD1FFr8Uf2cTuje9qlB7iAfJn3aj2Eo+COHrp0
orgwl4NPnqss4CE1/mrrLy/vQ5z/S5QAJ7+2OWwruX/MOE1VrYDOjBQ9mXJGDSHC
jQ5oG5wjvGPu35f+jwwFvXIIhKtWRvpWhi6xWwl8L1DT/6covzgUAQwIs5EtObQK
FHW/qFpQ3BYmigwFam6o/NH8cd+6OmPUVCuGWVEaY1ygRXmKrOwfB56s22/Jg3cK
QeySEn3v2gciV9PtPabpwNxdRnfKWt4pv5KRQW2yGKLKkA32i5exO0h2Vk3/Z+rA
P2NVMzPtnZcIqsxZWTdQYvaTZ2BsFk6LyfdIhTKTGr1aSAFM5wSImVjNe+ZMCIe2
o/MBfyX2sPXKPjj0cpOcQjnpZ38bR/loWTY7q3KWNjFh33sJ9OxpP6gtR8in+FN4
N0hifga1wolyCkqcNBq5Gg8xSDyfU0vJO0tNd3FcM3qMSVKCDm2AJFyywfhLEgOM
DchjiMlPmzX27/LbJkCAgQMf3uvOfeNHPKoD/lXkpWqQu7WUx/vOL7AMtSp0DQhL
VDwpC6bIDKx4cF+vEUkaDmxCT9VHLTSkK9ypCbe+ET2I1d5LHskmvKNgW+QR+Eif
se/cd1k/zm1qGijliauRBivZBGcibNpXO98J3hL2R4TjfG7K3GlW+TdGrq+QijWS
vpkZAAyC3KDaPfF8/tDcX8RLhWeCneRDOcex4EEOri9DWiIIsj6cXAv0glWFxME1
fT4IoJMdpA8/XVy6lhZgrceBUF5AlJnwIjr0aUkzRNhrwXP8Exk6zxNzlFxIuhh3
KkotI0Gl/Fvk+XK6CzS/Hh3Vdhv0gIPCEWkwEJLBywkKEFdZ+Cw34bo4QmZaJjGA
DXQHjCx7/mklnJpCtuRpErmUP1xu5rAxAARtMpneXwrs4pPs0IBL3lTYMqVW9uGz
Ryt+7oEjpLjuiSg35yLTZa/0cR5SesE4V7kTQklIy8TxqDWzCIGHEWq3KOMXYYlg
MXT+ffNawBCV83otEgsv/voe67aP2XEYiJIxqwmJQzQ31SkBMtlkFXyT0OOH/3YG
sbeGM1gS5e92IzFLCYPime4EBC8rxe4OABOZcc3VGSatLDSKb2lDbXfH5izUHu6v
lULuu/2geyeu7prOUHisoilsy3VWyCd/hyJkKHhg9WLwnOq5xqgUJvM12+79AWL7
Lna0g6X7tWfjo4ccmm8SV/swEucNNJn3rj2KQF83TkkzA02PTDIDBG8KmMuZ3Ayd
3crRCUbuX+HvjUsnQduaJcBkg8xk8f/Kk04fRk9ble5prhiO5giDxIbbfrBanC30
Jg3TP9gSihuK4aisxfSR3LHNe2PdqSyZXiuQzakXNJzwp2qSKNaZNB8aAAlhalqv
6OUjbY4TmVTOxuM8oqF1w3TPu020ZeK9D5wRr+DFjqYraKmxL6puzvI8x8jOnSnt
suEaLNSOXcA3kZ70nfF4wqHQ/THbUeQAG/tvC3nHoKPnKyZDFFJyWaJ4CPlNZ0Wg
8HUoNkhR58HgnI/z84wZ2JddKzPCVThf77p/XF9WHaGR4uqEgD1bydL2Ib6F3Vyp
+Lwfii+RZuOvrVWCnx7nqdZRo3RsJtmkZJ8FQAYnCJiVQVa2+sMGtuTUqcWZjdwc
NPdQTxCFXq9FYBzjy4+b41h8lyqJNVBSvtqpwAIQvhoPyppmgSWtF5Y3XvTnjS4I
ZbdEhg26TquxhidO7TVXm3YAdOV7O0VjKE+aqR/coYEJe4IIdfkIKYCS79hkFUVI
wkYJNEanqPhlF8AQiefpjrbWWAJHjGU6Vy7ao0ODsYukG3vpLPp8ipeIzpCaJOyQ
DTx7Vxe684Ewe2ASaFsgvOmjvR1VbCo/m2NX200qvrFuFnrHvpfmX3pw4S76ghAG
v6Rls40q5Xvz+eZcHkBCvAnotqwE841btAhFVOp3TlS4ry966Bo0NQ0Zh5UE7xsl
7XDT5NsTVmGnNjwbHyQ5RWSjuTWSE8t/vLc0EnYUuf8pqd2hxyZK/6cQCSUHR6az
Uhb7xlmKT96reS5ZlXfcUGXbV3E0jtr4As6l1kOIp4TfhLW1dRF/p1GgSMyFrO7i
iVm9a/hvz7RJma+y1FqR1QSoLtG267GjXVbDN8ohzyLMtIiN0vkUTJeTBxkU7cqz
eZwhF1SbUzjVGT+hzw91TRUs4qV8ju9I06jgiwVxY7pDmYBjXrDHugFllrtfbNeX
KL4ITMTQGJixOFeNVGIIdXiJHY4bjFfXSOYzygR65kNMi55A6fyLgoIczRlw0JPO
5N5qLrHQ3efAVspyymQU/HdrbXkyaH2rMjKsyGEI6NAzRJPV10vbY1heSKJb1CEu
VtlrZThgryxD4ShpaQNQHQ42nBtFKwY5jn+O1rB/tslu6DYjM1QycpcePP9YFqNz
3SXt805U/8Z4xGEJEiaq9JJqyLUKKsQlxa7KEhaU0fHisI19ppGlgFxzePV4n6LU
RgEOFzMs7CDUudkCX2oVeIs1D50klGANy6OCPEaOoWX1VO14lbUkG9+h9ePw2OAR
zgpZhROhOiPTYmTCqYXG5R5UTP1yzqseuhJtMeet7L3ljrMJCNjLjm18j86X94Rk
s6oqVNv2OfHNjLuyyp/knvbszpeaJMacD+XVy4og8GtR7D5JxeXZvwnv1y5euLw2
hyoye3HymLkqdMCoNuA9lUeki1QjK6/6UaYuCe1SWZoDFtjBwO5OGG9Ml/sdwoqO
MlZkrFiRWRmRJYTtQMP4sbNbPsudjfwW+hpaREFCjCBiGhUW+0yZpWzGc0mOLuk5
xZI9N4bGitvSezcqJ79p7y9ydqwAViQrAKFrHU4+cMYBuO4SWE0SG7FQZw/oBzcr
c7JffaAlmpxfZYppLa3T1OFRaVB+DZfXGoCUOyFXSr+AmIUKMky6AgVRFgU45lXi
/wf9crC30iQBC7XGuIuhGn92kgrR1I536pIWGyA4ZTDpYD6gsK2kXANhDUqD1lEU
ij7ZSVX5xsp4k4dlzDDvIqu06fKdXbszEaCtyeW+u1FIhO/kIecxWNbaMjoa1nkW
MsKyjBaNKtyfg12tVnuAigztSzbR17MHpNEYXxM6x81Gfy9E8N/iO4018EMILth3
k19sQfZipqRLu3mFOCqoWk6M/OEtewi6Vx2FSGL9jqqca8e+z0xdDbQXYS60dWZp
OV2DKbVvb1FlE7wFMGuAG/+7vgREkuEzfW7i4zh/HaxWUHDYeNKjKWZB5kv4s3tF
zYEAHKOoCLtUhjva/rpo/EQI2jAZ/EyajmqkVM96HcMlileCQQf1B9/PCX8Hb/YP
SH6x9eFC8NxqtdGGyr8Bx6l+lJqFEDdOH2n+iBLRoK8LM6/MZf4oop9OTNxUE+9j
shchzrJPy2QaOjv6OoR0PIm3gLaOghToW4CiBtikUc/dTgDOvNKPL06xvaeWKzMV
tNVuC68oYcaggrt+jCnfAI1To6OGyEf3/TmL99DrJELtmMng03YDPKbM2H/ZCWSX
Ghr4K2KWv0NbBjAscJZezdpMa4esaxrh9dL1Pu7plWyClUo6/GIGDctfXzgjMC74
GxmwwV+ij2DAEIjo8I7aLZFHrXQK3K9G9WxN9a9AdcyqQ9fJvfF7iursF/w1PeHp
nkPIexJSBh+TMLpufmytddWHH0KkZvGRf/4AVHk+E3NGuMwS+rjKwMcrVX4LM0Ba
Dn56LKjQo0fNW9GDzt6XALzaft9h4x/ENlSg67OGi7Dy7eRKm93Vj+a69LSUZrxa
ZZLZNkrMsr+Z5OuvFps8diI7RRk/FTRkMNFRSKArWd+oUonmUOg7twQ5ORXEWU2u
0j3ITiQ1tNeyzPHUXKSqJxgPzSj4yRwyWG1yDKyVCSDnhYdQfZgxyXmBVkSLF9g0
GELQR0HUJx2uUyMsQdQz20VKzRiRoyAjtWLfV4faNjjRHTMZ38TRnjfPsbbZx3+l
CzbRvWBo0jc149dCZaW3Wovg9OE31XGGXLL63cmNmF07EC0unSEqStJHWxJCTH0Z
ZH0AZWypwurSUyUDTdGcKj1/6FHJDlFZPU8/u4unHEGX9/8WsAtjVtAgSimAllrT
FWrxLONh9oQu2b1IqEgf3xKip8KTAQV3PyZbsrIQPQCZFT6gYWi2uYdgXwW/TzqW
dtmozZDUQFFQ0NIGbXRHv+AXDp/Zeqx+a2RrDqLGr+yDCKKqFDueh9R29TRQCoTi
+bPqljCNQv3ckAdOqBth01WY3f+AlPhrco/o7/z07Y+N3bJYNslXSbZy9DYUe09i
JqKn/fO7EQD0t1ZhCjx/Hil89Mk4TKY/hSmpVDEgYwRh2OHg5+7GUxV2Hl8J3Fyt
xvnTZeBzq/oGoPe+jH7+4iHns/d/DVPpUpRa3RxxN1p702o29/A8y8dlsxKgSHCj
6WdRz3THmDdSvMNuf59fHQdsfiXcCS22rsut4LHhcc4kD+6S1CjjrOG2etJXvYT/
VWy2mLtNihm0doJf6J/jlFvtLbLf22Vp5veQgidmW6LsclIRK6aQA/R9SqhMnJuU
Wb8T9iS95Eii/VU9HbXkJ4rK05Djn/sxOu7U/Gb9LYEeB/8kIP88qN8YoBRV8F7A
/qEm+tbAentmyz5Wse9Wct+PTyvYhdPVfbThmC0yPgnCnSLuuIcPKIdLhOTxdF/8
Qa3z9UyO/qp2tX0qywkoRUmGHKgalQ4iGLcVpmBd66+LQ1px4ciNyommDg4ecy7Q
NO/1+gnpWGulcMImy7X9hYViEowUlEM9HElfTxNoyBg2CMH7aOArUXOKBacj366G
f/1pL4PwaxHZbh33elE5PXE8OC0t+WLYffxYsktnb9iGdMhlLGNZpc4rIUhVYxvF
s08/IGVIt+1w/7Zhk/tdynFiYZH7fv0xby9NgsdzwsHvYiNhxkDLnRPcowvFaH7F
V4BJ2ADCdARjBjWyuiYRWxOXAzlrdoGHbIsxIfSou7xWigWvcnK3HHcnZVRx4nOq
/vffyR9MBEZf7rQCBmKhGTde8EVC99+LSMaydp2K3QEFRGai/Lxz9un1Uwv7NNCv
P7aw0O5jdBfNx4V2f3okaedVGXDKuvbHzF10OnONeEV9j2BEsE3ZtxuDMcWl1+Lq
oRkmDHmrU9reIH+aDe7x5ZrkqDItXb6MTBRVPvyq1IbKVmPPrsnrApcAL+uTVjBa
em+iqmI7Rx01grPjs0NQ61jvJWuVIb3c59NedokUeZFnRv8O0jONV9/1zO9jWyOi
YzJI9afycRRoA1BoJkQaEjiskIbQy3y/yn61J85T63ez+4zPh0sY5wv6yzfTVwct
3JFn6hGIml+UkgNEKieA0ZRYM3h8fJNWkDYqsTFm8lVxCQVfgRa054MxWvXr0J51
SIYRV3ncK5IoUsHUzZAfVUlfrLMD6s7pqYkhUlEAMIjlaQMGfg24XAbG9nmAvHlb
uA5KVvcUNNMSprU2wcwiIsu+knesoCUbF/9Cx7o+vY5gDBeTgiNtRvaTNIXjMMNc
YvpTrtWkrcCrfrv2aOqbfom7aB1JA6vdicCz3/1+pPI/OalUQqzz9GgGSyzUaUgh
57mxpZ5VJz4Nw0CDPhbbS2/48gwmPhvwp0OuZ/Pa1YKOBe7h9AlE8+wSJRvSXN8E
0BJKvPTdCEfYJHy6h18VCnjMQUQUkzZaehBEZBfF+selwITFEQJ5jUjzEk1aLbq5
bX2qRHctNsxukT3FxaQbSwU6LSi5Ko5r04EsrwHRXs/FMgGg8SPWSdBmfwtXJpHk
oK+Lu+WpuCj7lRYkTB6FC9PP1xbRh7aF0mZevT2neU+AwhtkIXAL/Jj//16DZMXG
6xw7RgMaW5S/CvPftg9fb8++swnLtxpPZsjgp9T77yTPS3KxlBxMo/Z3zksq6mSC
RgVzpw0q1G1+v4Vwna2uojVC9K8cH5P8/VAEt0UzTr5Nm8MvQlI+aen6zdbgMSEk
Ek9QtAx4opmyxMeUXWS9cmd+tGHGBUlcQZF+E+1wd1f2teTnx6zuSsaODvEB2CtF
HWAX5oM7wyfH+B70ClwhPJA0AcfDalGky0P6CDc46Tlksr9hfvnCV1+CzCVnU/5S
8nlKlU6lVuuXWJMj8fs/nVHNPw86R+VLCGXKzUgtE72NUzU8kBESN/cONzA+nl36
kTloehubOhJMCUTHDD7iXN3v7VW/8iZM4ZL0liwWYpii+7lYC2xtfiXI58OfRep3
tJcsgmVhWvCuWov7/g6hGFRFyyQQ5o1RwzbXDlaPSLNTu3fiy0662sSJimPgL8Eo
kE0YH27sjU0NlzYCqpcIc54Ay/ZntXZ11z1tcMWSqQvCel6WDBqcT2bk9uApTSAO
m5Dw5c0nptQGUdKBp5kHtdFbTfFfaJ96Yv9+k9w2345+/aujRIRN/zObcIVQLxYW
OpndxwoGFeQnWge9TdO67IBuvjUdUT1S/q+TueEkKf4YR3HfkYLQm6G/JHxSXRCq
UyowYw5hKQdda2JQel255VfloKReTB15wgC+nYdhnom/9/A0byRQwiluUlWhzdoX
dq8/OoHhWWsKo7tdO0U+Xq5BjEh+PqCEfQItC3w7MSaG7XdVSLd8dv/1hjT8bNKS
O+EfUGVZyaMFPxIEqjTRZFWvzWLjsoHK6rQWrHzte9OceHZOox7yhugMIGOFO17y
cbzKwGWELQE/fnS/4J63dPg1c0PTTNJTx9DGJvVQllSMThF8vkxClBrcNc2XpFyK
1jHtJDpze81FFrDZDfx7C4Si7vVL+p58KYkwfhSholuIXSqQ5ZfI9tymWHkSrpaO
D9nP+qWdQ+6IU864zkHTCuAauqFo4puSlYvI2TInvm1yQVNkK5kT98ocCuHf4pp7
icWzthPIjqbYdM2l721FuSgeORSBVNSnwI5cvLtB6Fn74pNsi7R8BMiSnXQYgZta
XM67iQ9CUQ4pALuyFNPWqQ4v0ryXCfX80s/R6/W20OvCFY72QNUyWclpAPEn1+xP
1eszMapAJ7RrmFrc5/caYAt2lQgD0TNfQYca/qrWAliTfU73EqPRaWqzc9uVVHoe
pGsMdK4FFN5hilXHFgcooEusDN/dLFmmia7zqHkyYuLGlBLOxeVcsxA0HesNKNQV
9K8rSzDyjujtA9KWatGsI2k27EvhamuKboYic8Jg/QbB+ged3otJFJr/M9vWO8XB
GXJbXOuriODMekqeNTQwg8nMy/mFvqFMb3pCcAAGSzMBEKk/sGbqWfa3EW23XNkA
svQwRawe1auJNgN9HG0BJ6hiJx8eLoGipeFP+t2keLo/y16POPE+8Y93svmB2USE
K04xO4XstmGUJRAcGPnhBmdrTm6qCA/nUU4fZtrBIZhk9auw0aKee1ws9GxAa6It
bOntuLYbyYLrK0B4msYeUYiISI7pwBqPv8MG7eEi4BYems2iPWAu7/DekvhdnerO
A6jx/jrHHobqHpkLuLtvtCbMYziMw/4gWmqvbfIXjW3hLAdDQCClAdeviHUxxF9w
pVQjE7fJzT3AMhKSx87Ue8pMqFaY/GKZQ8JJJdL/DeFsAO2iH/4DT6ozeNYYG7UJ
chN3O5EejFkr8feqJqoWLba8XkJnsbsBMJCOYgHm/0ja7I5ROrSqvuAL5KwxuAdl
/0+dDTFM1czI1LgBesAOd8X/MVb8dVwb7i/2PJx9lYJKV1WdhpacdVggX6f40Bso
OBJ+Gl2hThiS7SzhPn0o0WbAitVnO/yQYwKYfliq9V7AbqPil4D8nq7eh63s724H
LwtO5h5WuZgNouGoOVOd2EbHMsZ+nmXUbHAY95DVJE3eWb/WfotMu3tslXA9eThG
SwKm1lkIi5LS8Zdo1xoc8EhPzqCLVgMspRLxCQovLphxEEsbM3RuF56SY4D6AFtK
ms7k4CnaJSnaR53ly8em/dTtODxkyoi5u/rn2MmV4Rql76p08bDHLt72+jlPi0VD
9rF18eI3/QLwIrpOxOj82YpPZjnnHAsao+YUdx8os4mbNtbSju8STMmY9X5MA+dI
H1to/kTnsaSwH20hPj4pVdTeUcIsnZj4D/wYt0Kj669GYFKZnqfPdd0MDL6WMp51
8j+lCY9WBTHawoEQfObCzKaQbI/enOufhfA/EacDXpX0HlcYtw9kUjIcb6slhqmZ
+8JCBtTt0GQwF95xz3gae4e+2jkaetH7Gj6Y4vcNW9X4vlewjxFOJBp9h9ExfAh3
rFspGO6cAErhvBd2V9nEnUecgMIZOYqvxAzqBEYhX3Az3QpiQ0Ry9W8jPiq5lD02
KG+LEyyCnun5QmFPSljbv3GT2ODRThyPlmeQJ4yIKbv49U+06Gv3YlNEPYVCwRp+
qhd2XZCL2FJW4TranxO/cDJyTsAjs2eeaGbQYa3qx+at7MS6ikiU14/Ab5Ol3KB3
TFY8B7UPonGaUOBiydAcktuDx9AjIxqkvfRML3aAvSFNF/pE1WDcMyFnKV7Zfa+q
iqETAyl2DCIyFZMvIdQW5yZ813LorAw0cz8mgb3IUSllH3ozuRS2D6+QUnVt98j/
R+HDVrvZFGxiOIixTG26/qN9X5+Twt3lGw6vpBox2LrefCAqx3kth3jqglaxb+4a
k8/NXr3WA/5yNPuQWcs/LQjuwkw4dSX2vnacjSPNZ/vP4DFdDKp01GMf+AfDNgKS
ACZuEQIDh4B8c0vhutZpw5NTjEnO8R9crd76aSJP/Fyeqx4kLyNRLccj52bSDsVG
CWX8lfT6iRTc9C6ERb9ut8quaTbQPvdyPYQjpjSF1vkkKpLCnhogedlEtXoppAdV
7zgC1Tqa1OkMm974FAr+Tq1ea/TJfOhiAXHk7/AHFQaAMfGIw4AI/J1duWCwNhcs
5xPRLG97hHMJWX5vbUGeDS9zCWy78RPKadCyNf1gNPT+vlvFpgGg0UwccDDSqFfw
Dw+XpUCnr7Mqj7/j//Qwh6oKhuLIJoJ1cA+42Hur3ebrrdzBPs9bMmpnFKRnOkQ9
lM//XNyXl26A5sF3Z5reP4qH5Tgr0zuV3mQpMX3weFO0h+tGvsgplx+l2JLkGuKh
bUaiFmWLOGQwN6cIvbq005CvRJ655Md1IPDxBdonpJDn90/VWb2pOdkh9GWI5NcG
fx/uYE7JKzNjTE9J3mwr31CCZlWq4ZtWTbqe/pZgJBzSKmyYyQJnzgDajoTKwUxL
y8wBNcu7MjXU1fsfRs25nIYRF/QLFas3KfxjkcTJHUxN6NPR+TbLcc8+nfwfCkvi
qqGsQf0G4cERMnNYmYkycq79oOZFNL67u8W6Z+VJTpc6GKCiSZjBpG+vbV5hE0FQ
DUNFZNcRMQZH2dojNvmnz1qgvR3pH2CXuJglXTZg0y+fUECOuPgEvzerRJ1wFaWp
Zz6hh1Dd01ua+UmRo7BfNshVilkpPrgYBaSM607hGRk88dXfqk/BK2xGaENy4MU6
91fHuCiNQRzVEM3CZiHbOs+KP3tIRXfm5FW0GTXoPELN8HC0VzL2lZMzqa4EMDFV
TzE+ZI79DIO0INu2K0DIcYrE4CXvvsjJY7Sd1TGaSgZSwjkJ0IlEFXTUSsvL/61L
7L9bWYMC8QX/D6W2NDYsOVKlW2UIy9V4eCKU4RrTpkRi2o9/rGM0jBPbFhafgE7q
6Rp6GDzxdYlaao9373etylO2O5BgbkworhLMDy1A6GLQjRLbSY53AWQ031/cQUe5
B80fWm3pqPfLJVqEWnxHSC/LxrBic2DfGYC7w7QWN+4hRnBlzGVdf2POod9MKAy1
+7Un0B7zMaDJE4LTJV04JFhEhRku1b0fiwZtDtdXigyHKwDVIa0Jb0g3nYjPNqTe
LUrKr6kkfE3aNk5YBGzSw7FJxmoVK+1eVLI1tZcixElkrRPYur671GWkPxeVeK2s
COrd7KXswhpw/lzBOT9pRhkcuXiGt7e/LQo1D3MybGGSJ2F7nnxBUbKnr84uFjnA
T4hkFdaEcklTkPk30rMefvbRKJfn8E4hTJRdDRne4LfxKnnxhqMpXdpjHB59uJNc
21DXTFkZYoJkFEacwMlPpqjsfhP8q+IIb5D09psCBeQ9pEMZ1k71tfHYL5w1SgwR
iEsQ5v8+TyFmc4toGkUEkbDz59hSJ8xdfM8VHNGLXpF+Gx6JrKdX6f4ySZMxhgYx
U7UF4t9hx7NZrquVRG0+nMH9HCucoiotGxAX63fGzUT2T/b6/WpR07Fk22YJaKWV
T7ndVXfY+VxJjGxhEmijLni5FQw47dN2wAIi3k+9qXhQLBPLHsHAIMtZRlpLZp1W
vVDxShetUYcQGPyDfabNSfr/QTsPnDz0X7XqlRE9MBAA+yMifHhUT9oLYJlmS3WT
YMsnzqF0uq0+QZGyjN03K92FmMrkY+k5Zq96zjw35zepPXFdpmqcFY/QrJwAO7ND
5mc5KH3O0Rbv/8fBP1MFG0JuS06LsTPoF1Kwm3VbwUjDpL5oi5S14fYohbgJ2ozg
q71iB7keMEymu+7gnaBZ68pNtMnvbz94xgMtG0G+yCSRHv/2Y36L9h72dovPnr4X
MpM2vEStgCp/TsIzuY0drad0tVYTApChxgah70u2YbaTa2Tfpzl9Nq44B3inz9j/
CU+lbGYeSfqSyxmB3DISEDUPZQo8M3zaWrD0R8+F1VXNQrh9ijrsyBS0fW13CzqT
Tu9HI7/7b9Zh6OC8fhIynZ4i5DIq3TaBeR7fYeUXJS7bdnChXmYyRcp8uYVbWblB
qJtwx9+Ogwtroq2YrR/6I1RV8BcJSXIR73YLw38nJHsD8E/WKEjrdQqKhYRDsIlp
IpZl/x7EI57GMLrCH8H6SJ8rkNjiLG76dpV4BVltgPLI24rXZXc78wDWLKps+WdN
waplJuLAEW5/IYdiI8oGDFFnUUQq9I7RJmWar/IAKVweX/jxrJFHGDLpUNFw53Mh
opTRuDo29VZXyxWWwP2YFiIQxZmADUWDZya6gPbj+NB76RYMQND3X6ULhZC0r1Vr
WGiTbICqfR9MbkN05smNJjBx5m/UCUe1R9PCSaPt/IAn+2r6YOHs9woce1eCU/I/
gn/r3Hyd2rG4ba6e6Fmb9UWFKJ59KMKUXGhUmRy4YKw3Q8ZJblxL1mqvdBqcs/J8
Xfl5gaie8LQ80Gf6WEzlG6cZEbZcZKCxYjGVynDYkUGic7JLU6E1UylQnh0GskaS
sRGhE73XcnNmg3G4SBYMpCBPDk454Uqr7T6PF9pn/HJJGWmjuKULtwD9DVQmcU41
vqqyBRj0qtRdLizxmvgeqoIOzW4tDhuk3y2fHuHDSVJ9FXlqwAKSi45Z45yEUgds
Hnll/5BtomC7WAcMJeSbXphwm3Z7D7+3Tq8R1Zs/61haRtbb03ps46bLHspQzjMj
VgcpLVeQhT2rFSAeOMl12qojANLqbYWnHK3YNvKpqclgcdrSaReve8PjtGeTmJzQ
m/JY3X7xtVSXGBEnjmRFHsHv8dNRfgDN3ggRPWktA0KAUzUcju/l1FgFqLV56FAx
ak0zCWOaY5QHSQoFll48kQKkVv2iKUCGYUjeFO8A+myPVV3z69rCvEYqn2aVRAO7
+B/WZzIeu6HW4azs/DJyu3CwL/nK1R+sVbBvFaSkGapQ/iQv99g5srN9lA7kxgPh
ghrQosYbvdFyWmgNdN8w//MvPMeGLZ+3aOm+cwZoj/Iw2m3Ru6JeEIFBRGorJzKg
Zz6NVZ56PJejkDCr0usMbIx4N1ZAzPD9ETwjuSCecLruScQ4mqr7K8xLF1vVd/oR
YWxpiCHxfQBqenSwXlLqi3qvpEyhL+MnH4ZNzg3qW0oUygh+lB37usTvBjpZkRT3
wf1qBsaqjSwG+U3U0tibJH1dWfgoeKqtBB/o/WnBzMCmiogqjR7JCTwDztvJ6vd3
XNV9JB8EZMi0M1c62LYOdjGcW+CyanxexoQlxoC5fRwp6d8Kh2ZRMRA79XjL4ukR
Jj96NWaoe0KZoyZMmUkf4aZHkRHbTOFi7cGH6lBhckdwJWcDqTm4nozCNUhT1G+y
8q3tyqRPr27rW9yf9FN5mM2Rg2EVakWVmJijbIA+kMSsP4BfiU09LupnBS9H+zTA
XDf6awMDoXRVHLhP7RkomotRuJM/SxvlVMLGPcE7Hs8t2A67zVAE5YRRCVvZW4Z/
AU0MvBuKU2EGTwGMYJK+SGow8YOs8eJwiVdKU2mCuEMBN8yZsUHgMf/aHNjAEkeu
jQ4VNW4n5AkcbB9FKpjz9Z0HDmr53Ew5EgiUdE8opeJTnrnyteJ7/+/exF9nzL6W
p8ITBZl1C8oLTtGZACDqnwsLQ9duwU7ntIvamga19LasUB+S8FHflVBElNdTbRM+
voIN+h+NQ3ckj48CCSv9n01dxVeihps56cs3Ocv2YAyY+ExuPKLhxufZLTzyBHz0
NwDPsYt4IbDu2dL4ZmNkEu79TIN1gHZ49etyAb94ZMRNF1PtAtdcmIBh2xHxFAKH
9JKKq7NJHwdAp1XLGcc2c3YXvMZ3YwHBcMZy4/TqDoBv5/CjRDvv2IUs4uUOsj/q
09djj0h5MtYbSswUaO95lMj86AILmJiUVHQBKFzlO2hCg1dwl9xjl6vtCD9t1aIf
hrRYChHoFMe3DGanC8kVG7bx1hSb8X38/UDbXgJLGJAARdfZai8GSZ9dahp647b/
XKVR/hO01Iqq5HB2zvuVRtBl4R3Y8ycA3bI06sbicbdyrZZORD+P7CCAzyDuvj3V
VRvDw3njf93zF3HPGmXim8xM59G375j46oEmC1r7lpFIRItyz+mzjX1CGicRECrz
X9hvcta7BpYru7tT/a3hOfZPjnKXQfLFh3Xn5o49xRmYLVdEhhA3jIP1uYFR92Zk
xXgFNWozKpPdQMT/QSA3xMlS46huQNMWUtu2tccFaISLfl3H/TCrvEJQuk77V7Td
nRrNx0d400kOxBXHsAZ1l5LnS42k+9opTqEAHygCyqSvy0H5TimIh2oiWwK6m946
Ghcfg7Unr+WtSUSUk3SnVOzcG/K0vjRX1vMqvXaXwL1w/wyBuR2bA4j5p7/fskVJ
ZfIF1mfSGyazCUvpohWM6EblTayHsFC8rbJIpuO9KcsldO1myXc1iuLXma8nHFUZ
XTfLuTBwZcOddYzvmtA1B7gRDGyXy3DNPI4yrhY1v+jw/ZjfKCk0bDwQOXXJMkau
2tVtkmge1jV5SRo0+r9iwt+9EW+6rC+AdAEa7MbSM7Tvki3LyXxNh2uvpy7YFtqv
9O+04hdJ76qMOGpgHzUILPNcCp8kWKf4fIkxw63pBkFTvUunJVojbllBPvaqTA6l
TvMpRoTPqNqVftwEyuiG+QTFHhYTuG3a2eqjOYR9m7O724wvzi3uZoYOP/XZQWtE
gnzWNtU9XyxyPzhtofqG1FvD3+mznCrbqzp1/0yk+5v7RuDQVbNArGMuzOHXkulN
xMKfyVm1BzaEew4+47PMOksmAM2pEr1eNxHCObQ8+u0/HTO4KSVCr71Sg1kx47QW
I2W4Oz4lMnOcdXkohrJStjIm2pJ5EReKkHIJ1CqNaUAiOMbAKVGRNbuNmz/pLYh6
HaMaLdJvsy1HdBIZI7Spp88hACZ1zR6qV73Sl/R0mszqkz1iOnwUkxX+9Y/woBQk
G8+wfzo9GfiCDXDwu5I3MsSAlmxOLVeT2cuDRMAXTcEC+P8t4QqHPNQFK4kS0oNO
SdC7vGrdNLU2XSyGED8iHb4Te2qeRa5S5xsDTfMCvxqsv/kuP2TZ30ngkTmyLDM3
mm9x6AXx03gy3t9jrWBw/ncBPkmkoWpME9TtqrKJJauCFok/8Z7yH/cx37k9AMs7
6y9F341bHrcxoHHrvzt3som5DcvBm0CxabHNF5F6yxk6coGsnMfuaZh3oycjvC64
QJSSGaIbpahKI4WM/vZqGlTnUdte2MkuOix0RvqXEOfUNKNif/gnrWv5OulyfNvA
t0fQktj8NMyn3I6cctd6v7MBb0trn8AqGD801rg0IMe3VVlNbsa841tW4HGtzWnN
rLK3n/PUSSY/Mhf1smlY4LpMuz8F/iZBAl6bVAdV5WynEZFjGHx3h4DyhoR6rU9C
3IuLhlzxcJ8fQaY4Uiu8yzD25Qf/ee8DDY/8LrLwN8Qis0SyDlT3q+PEOXHT0ybq
oSxVvrSHnkB9FRyjNNMkJoMXq9pobs8XTD2V2eLdbLVBEHOxAokmeaZE6NxDpZTn
qKfIpcbW2bfp6UKAuNFvBACOIDHX1SHQk1qwl4GBJcI5gDlOTB5C9s9mSq47CXtU
b3a5YTpXEhqz3wGQ3GU9gzKkTYdWoHtxbt/i1tVs1qZaQgwN319cTLAypcf9W0Yn
+xXtJFppbQ4tVpWsWguBVxQX7eilHpAV5hx+f3XWYxiglidNkiWy4pZC0kgqEC1E
6AykzcQ0ZoATrxBazqMQwybAstvE9KoEXujMxIU0Ql5xKDFWATtKNHNmps1DNO7y
Vh+Y0Hg3IJoOgTM1Bf/IEmISmftzU+fltxwAFK173Wcx6pwU/xE3QHxxYLOjD6Ju
3CRaCixPmEoELbUf8AeH5EihFrqK7hrhDs0sfAjyZMjO8YloSSvbtRHlFX0dyquE
rHMQcJZ06lyzGIWhBs1+B66MsRdO6FlrjOhC3eap+G7eEm+vhQONzsyf7njF1Aco
8ZWWYjpYqnyVz0losLLvp4PTDfEVHBZp1MDqhnO1nXnXHe7y3H9jmL2+QAiMW5pZ
d/tC6N75ofdXooewXL8dTGoPejY5ZqF0a4/tsDpXEK6MJ4fgiY9i2feoHS0RA7BL
HQTnO50sYbK0KaIr96o6hPmp5Rjny1bXhnevX5Htj+VyR0V2eSrb8JMIYIQe4OBB
1LneaSG99AmILlt5emldPvIqJbLIJaVFA8ihLlzRn8V94oFg7IlXqr4yrmFL/mq/
/5FsPzu+hYtyQhB3294/uYpzz2Mn8+S8GXsDym7rIPbqahgQBzBUbFE75/hDOggo
hbT7Si351xv4hcOdx4JmEQbZs6FQRnTgYFVVkHo6w/XxSm4sjN9cwkXrYQAAR15Z
qWvxUVVgNHm1M/gDqaK/pPTMMlG7X4JsZnHDurX2g5s4WoTPz/4ElwOZo9D9beJH
/NUxIqXLuFiFyoS/RpCPwtOACwfC2onEdUOjn6n4bd3rL63EojlNn8J1yCg0nsS3
L1b3rUMKwKfyRjM9XYyRn6kPJ9qEeMDm6VLfcApc2SoN/H6fdeS7VP2MjZD74Jrk
TFfUOvhMj5iLzsMrwilOQhXEt4xMzDUWooc0QDOOdMCHn0Hn5ouH75g0dSa6PImV
CJc2a8Z4U3/pCHY1khJF3vKbogXPW11lt/XhfiuRRCyioNUxCzBJQ3m8ss2+JaZW
EPCj/L1uSW7e83gXU08dyzscO5I5hTDlbpbCkwYMVKFVN+JLU0TuHx4NshbTi1ZQ
D4WXTlcq0cn9Mk52F9sarmSW86V4ojds2SObygA++D2CF62bRbpLHwfXFgP9eeX6
JiV+O+cFniib8qXq6N+OvrmGI0raPhl+NPq/stLLruamcUzxYvEL+oHzRdUz6S6G
Bu8yQ/PEI7Xf9PeXniWtNjt1eDKCEWqgqWE7v4qrOn8A8hxF55Z8kiAvmMOOCXrY
eNctjHLUwktl/ge+ULn1Gacu/G6loiF00Dvq5ZBNTPEsps14LVqfAmrPraEiIxf8
baK8P4i0DielfABbKHj9VAG/N1myf0wtvTgLBwBG9QoXOx6LBNpze0wQTrR4XJM2
OkcmfM67tpnh1wSEdLKFCFm+JZquxjTr9pcR4qkPC5m6aeVjYj3H3NtirmycsJFd
GSofPgZIeqQdquRDP/pDQYawRK8nc1U5Zd479OkwZkKv381cZss4gpkiI5k6bF9e
uoj8eZA9JrmnlcGYwHq7pZyWzP57/ccqpojBCIJBiAhdUAwyFgkHNbvu1p3EuZmQ
4cd6a1TvZOgR76DYr+jiq/QzA+sm6woAyR8dAD96h1SD17hgg5IKvj5guZeYNwI0
YUViGr6Re/eBMUp3u9L+rmMnLP1rnVUpBalm58549hIMwEFf7aY0n6GxRdgMkAXZ
LDUkpAObJWjPH1Xz2WDMdpriQ/jRz99p5qiqp9vaD0r1cJVJrqgKYjiOqEjShFXg
FDJcRYAF6BeS6YfgbYohRQxLK5OuVtj1h5VNF4sSrHt3ieQwDvF3qtIZqpsJEdzH
tdgf9p/5ZB8Itshy2feO1GZnGGDN+rNNL6kn2/KC7yXqF4+0p+6Sx1c5jutRztWE
Uxz1NSWwdgj5Ydcc3qKxI8WLDxUjCCZKRrG3jeW4tmOCMr6WAWO0jop11vV9FIga
TEMz0bMbqVSqqypClgPkAIIBnvfBuOXRHv9XP5+kx+iZhRXnQc7dJHRTheZf6SwS
wPkDO9IntFiEi6StWT1vDUhv5vcGMHLoGVIC8D6jrjmsf5FmihYilMH6A7WBbzCs
4npViHpfOUmJEBAVgAdHQRA2u0O+NqKRMIIKyH2SrkmmOnVolQw7m2U/3gkH1Wj0
bEzM16cwGu4anqzPdxGX2fqG/UcY3XXRJxBFHGGNvf9D6kaWWkAKfs85+pE/bP2y
GXNoXRktlhf+JATRforc/h3TbrHPh6xR0mQMmS4ZVsGRyNnatbF+RWmLWm7trgRJ
BdSVy2a2WOVxMprA7FmvEKCTDoUsVhWVVSYbq4tKJR5JTItQFJVPCmeViBUBaDvm
VesiAf5Fi87mB7NUacgfCnuXLXg0BnUV2V9ioH/DK6y6aVCQHKnc3rP9/y7/ioDK
pe6872pkjw6ILNStd0QG5BTSrAZXb9u9Ha617SzyEXK9HaazRZU7cZHk9EbDPhtv
uX6HnJdvFyYUVycZN5SPYZKf5aq3lWGmf+ZJ5Pb+hJRaytFUFtBgsZO09hySThsi
itsj7ccCZ6PduhRdFGy6z4FcFWO1yXyeCoNGcTOPs7XkNHNuZoEC/oYL67Sqor2v
9LK4xbxCSC5TxzqneBrSG2laLYAXdE+yhCHfoIMDBHzAeM24s8KI7sFAnPMRUhgX
FkYhuXEQQTg1cGtoj7j+prjr9m+eomsM9I9DN50ndUiDi7wm7E6zvJ8ygWimYJg8
bh1xukSLN9xVI49+7hidq3Ua3WhVn9rwmr1li0l4+TGBimmPNWFs1anIYL/B5zS2
Fl3KYziCSG/IYqI0LsWEQA/s2giZmP6btuW+vrugWKGTDI8Nru3Y/0h9siuNUgsA
5L5j4wLhWvJFPefWHTJSxVqPfbntozpvpOjjKnDsNDWvCrnnKCk0z0AwD+GMiqec
3UbsvIKg1pX7uuwjV6Zt2JL79muDJ6+JrRn2QCfED7d3CAHzAJNGK7DWp283gCRo
5u9boK2i7anNf9ikvj6qC+7E3bWkRILCjwisCkbUG8lER+dyOOVkGV32+Xjbs3uM
MqF7TkkpWCZgHKEiM1Pk0qz4WopRJ52ajt048YnG1XQb2VgnEJ8BBt3mrxBaKeaw
IbA/s0jXVbAxPCCAdxF5FjHt2zPrdfe3url72fTZzy9e1vGXHvKrAJHle5Kq+ynQ
5TkEs8/054ilJDXvwvg8wHS3+CS+c4IcHi0U2WYtuaVHI+rTn9oCFK/k+w6x9OzA
0s7tolmdXuUCtr/53KnST44v7AGZdqujw8vDCi9RIk54YX2S6iq/eEJCyg1ojWpu
NANHh4LF7zjNSV1jlKnkQt4idVSF0TdjCNFRp6peIOUCDsCZvVyqfCHCWvdD5hYO
YbF1K1l0lLfWx02ltA8/69apTynnCg0xnW2l4aKg3TjmtModEGg5+qL3weF5QULy
0z0ia36DJW1ZRpnRWGYdxETiEvvcCbhBQEwpSK0rKtjkoggAe8kqtWGxdlavZvAX
jlIH7scngJ4RpZApbOBkcKWHr1NgapLbkLqGjBEfaVN21XX0Y6ePH0G/JzTYJIBE
KJj2eGz3ODoD+/b+m6gQxdaikdVsmM0jhpybIxHxvmY4PnQIesWD3e7rYUcHza1f
G83LGdv2k4BrMgVuC2xG50cm1n2OQmGM4H4lk/m36MeKon6dRAuXKWUg/JDSEuS9
vFOl+UMjJipGJO63KVxSTsP2lUC2a/etWFYKPWVoms5ueoAZLcWt+ukUP1kUKn9m
9NaEGZlpZBYvZI63K7TCIk2Of22qXKnDjodoxMos4E9P4zCtringO2pccGIQLlEK
fwkr83/Z8qiXHp790aqQgXHRehLczjslC9hmk8GPkCE77RNLkp04vEqz6GNzr1Dj
dPaPPDvUnsDeMVdQ6y7owMZmR7z2xPj6zNlLmaLlyYxiN3fOw7nEaxldbKCPjExw
gh3BL4el2N1P1XaM9mGN9swBGPwPcxaBZGWc5V+ay5N7/s3VGE5dA7jP/UycsPl/
Ft63JpI8gSbosWg1AOMOuIJy1XvDb0lEcCbZ3SY8sLhxQ0wFqMYlHFX/am1HxsZ4
fsuIPFMHHxrCxBYItZSWLQoxQUYn8BSOw0Rpg3nQa65xoniCjOh/lsiqfynm/EwL
SHAmerhQ5FS+KrpR7VPn1WAcruEpVtkQ8t7Lx6rL2RDkWn5G078Zw/gVcUTA+BXY
/CoijqymZpJATpJmLMxrTRBY0743mZnqOVv8TcNYisi1OdsFnSiKD6mVMiQf/8JL
GSDH1ikghzcw0zpX/LAvMl9FVtg18+0PY+y0Zv9Ug2TV7uV+VC+6dwXj4MZPOsV6
EvXiPGg2+rNI8L9FWTq0cpqwG/7SBga9YTM+CboVHRLcdiddg2S9wgGx4fFEmdp2
oegWUzTQgf/J8uDw/yU9lblE20DtJNg1fnbJvVkk6v3Friv5ChDSzhxS1Ojpac5m
RqypSVM2yERbea+rWCs2OvxVm1QGOHI6Yfkpj+E3c6EeW/65RY8wjaEbP89kvhv5
2gUTIju5yAGh96kGhN9Yhh+HnyLk+Oc01dDFtASsoKWhfp04gzFhJEy7kUSvbYIQ
qY3JGlClxg9tsaYIvbV+YbFn/xqZylEme0F/QjT6O5IdXUq6kFtDfrQburLavWIv
rnK/8W7Xe4dKR8S787Jnh5zR8HlX6J35z/4vk+50ItcrcSQOFgPER/RFIrGLmiPL
SVyzHgF1HkLVvpuKduHNkEUTCJmCR/+G+UG20E6qFaX0loQeCpuKd/wduLZv+6MR
zGoT5ienJ1sVhVRhawH3vvv+A//D7iw/wTBBR3Dthw7Hz53pMifSqjtNQZpCcwBC
l4cOINA0B4SjBYu+SSBGLjhb8c+/RsG78yJ8NMLwB6zMe1LMYImWCyVtRVPKfuOv
pUZQZ3oa32P2HMtMBktzW8AJiRxHbOkd6IjeCoGEWU3+t2gmnk8Hxx83EtvNNESB
ksEjpszinWCfwlm5TFotGlKglvQtL+FDQNwDNRaNX6I7HnVndBVbELTAO0nrrLkS
r6mgdfEMEw/XOI8U84I73tFnhkNdNysayEtKO1rWXG679MPqdbxvnI3x1vfnQiU0
AY+LMNpM2I4fKGSn18cYFOCU24elNfhaCZwQT4LnZ987vMjGRFE25Ra8OAZedDru
A2A/sQQcW+fbFfpD0KGgjPlfnigdXqxUD6ER8E5vqpkP4Rp+EFkk4ZH7UM4D0GSq
o97A6VtCc8pSeUd/G7IBqyYPfuuQvsucRr32MMy5H/3KutCiwmwKDZ5bm0HQ37ov
mu6FoadAxcFG/pueNOzQK74g2B5kAwo4yXUORVARAkg1CP96wZeYMUW9xarevBsj
Q9Iaiwv4G/ke5u4IzALE5mXblSczIHD4XHr73FhBiv2d6oniMkRpOARPOqE9wR91
SlKvtYak9CGRr6nD2+k0Dl81vrokfiNOI0P9d6GV9/SiFQROhsgDxl0TSOtgLwIy
Lp9VcRBeSpTUqoYwtCsLQnwbdxfR1rggbf0cTEDlBJUkdaVcqp1fzDQcNN+CHPv6
AhRt+2YkfH7sEihFLiVudXNZJsroL3QhxtapBGCiAFFAnzLMvEYDCJePfHJVONZc
Dc4Z+FrikRgjvTIBFLlSz95ZBjPEol/AGizHRJofsY3cIMswq2oZH1nFLSt2F/gn
6RlsEdvetRJGdDFOX+tx8uwyOGwGg1UvtJM/J3IEWgyK0Nk6tZ9tLDMCk1TfQpaD
oBE2nUwfBFm4u9z4nNRNczHIldt4/aTXLa2ULXKXwa4OgMmKmDkm7AzbWicVBNvZ
MC8U7mkjDUepmP6QoMROVz7Z/H4By6GA46qggc225+nK0bVQGYzDduxZXhjBaLZ0
jDJCvJIiF5fm7i/YtF6MwEeXycdy2KOztOvOKjR20FgTq6WtkD1mgwEJNPkbMU06
g+fGc+ZZd3eO4aGs/4royqwFbpchl8q09deupZJxznZYJFwsE5h32Ky1AEOHEgRK
3M1jA65gWc00MsGCu2jvzXBskM63kUpU/J2NraebVMgT6d0UP/p6kRwItb5iNcdl
X2JSTDXMCCRZJhwxilqia87tScizouss0aDdqQFQBxUcoRdBvl8gRP3G5SpKb7fE
N3g/7HGh0y3Jslhjc4YoSr175/pPiRCpiwr+ieFFFeqF6z4S1hNCPlZMidRgmtus
R3B83041Ncq2RMb1O8PstZ7CkKkuQa3ejcDkcRyeB/8Bt2I6p5LETnBiWGiEQxSk
grr5dvVRP5qCmzxzIqItySPVDzXPcgyv6y5KxCO3yvWtAxsVANvjQUz6ekowGGKk
27D1QNpeuPJsYzAvKAFOqjFnXj86rMUYgPWuQIBKeOiqfvX7zxIe05FF9tXw2lC5
3NbozWOiFtqyTZa9m4dE2jCMusjRImlDdGD9EEqSXACEPnp6VbQQRyUKtqKeI/yC
9uanqSoCRW7VUMxuVbIw6n8ipaa7iU8f1HGSKTq0a3cHEfvBzMHwaN5Wrutf2pPK
cYl8c/1VVrjLqOrh7ybMsOh2iHt8s7i9Awpk7gSZXY8QAGuf0IbNu3vGZNIpaQQM
D6yOyE5xMY3TSD3fMsEwhqxBU8GFuQKPwmc9C17zGmB9YxDjQGcV9WTNeJhMD+5R
KX8TKhE50OEiaaJ8YE3Eao3Vb2wz8WKwkL5jGwlQXT8v2iHNO5IaSt7n0XVpJJyo
3vi7pmCqqkvcLMiGtPYlTQJxZgK+f9zuWoFxYovF3GFf8MNHyGLEIdBwkuv/xqmo
WO6GB07PCeDQf+Q0IZovDgveuPSHXx3AP0jcR8/ZLobvzqTmHwj/5Xs4qa5EkVwm
XRY2/ggnMwVuDk3MBkVFqYnGYU5fPF3lB/teS0SEGclth7HFTKU4bsDF85TBQAZm
wllTjnMphdTe2b0n17CUHBMyMurwRnSSenUMfizG+fsByL8B0IQb6uyejiHjsZq+
vNq8XS17egvG++tVg3vhtt5sX4/r21VHj1MUJ3u+bwSRjQ5Gk6T6raviN+vqDtD7
o7vNV0gs9vJ/RfXyCf4hGUhE2UnJZeQepBrhbboVnljZbWMk73WnTjvp49MtVdAv
K0RlCrUlMQElwsgzpGIeMh7lPNltSpx5eziY7TO/10gkjEufFqloI3+sepS58Awi
6L1CnrGJoT3nJvZb3DWmH9rUzzpSnhR7JADi7AoXhelXmzyqoeWkmb3fiwqeag9k
sKmPp7hL4WGdub+bVR6m8cwgey3Kx23x9mlwEcsQC01NfjuMvQVEzxHm6sEGYrAq
fQXRHicOuTSM+Ubbxp9GY8U4YxKgaXbSfAh4mHjY3LazoguLqo65D+UgJntkN2bi
EtE2C0KiPKtpJMkDciY202xnC3qCAT1l4fxFiGNaNLg+Ccr1KnsRA1Ry3d4eWMi7
UZ1byHUV6T8cM1vJ6nIMImA/RJnrsIEHVf2t3E+b6KXzcdAFZDgwbDNLokUMA6rA
09O/fMRAA0StUtKxI6cn1o0E7y10QCTx89T+/YALGGLsB1djo+RZxsEP1u8dW5C5
CYl/jjYn+wBDQ4wOQ5SwrdN6Mw6om5ptZBGyXfNvKJ4POYTS0NL5xYIsRpjKs+rD
PUvF4MpvZznEwi8evpRBnAw/TvR+G6DtCnB255K5LO7mQEVRzMjW3j+jheOqZtP/
nijDQ6ssqYCIlSp7WG5jhBkW4NJVsUTQXB5Jki3EoDU4b/Xd54HysF6V51Z04Ibw
fGz2F1clOkXRqK+EJS1ko/OCLpabD0sr6fbwib3R16yMx69deVx1wxiDi06lkFut
hevVH+rBbXKT2BUDorp2A784E90T4EZEXILcnWfzjz5EMkf1QKuu5tTpY7hetDOY
lRJ/sc+bwhH/68b789Z4N0EZ4lcjAsv+v08/0Ji7yTmY7ixyW2GMxk3GJjv2AZrK
Zi3nB401Q5ZVHjzdrHDWQbOgTpFn1BGo8PqT1zTh81CyiZqQhR9yQkC12nXvkvwG
Ed7Ih47ZWSya5ueg6+D0m5R+t96q7yFuU//eVZCiHuK8gDytYSCWnaHnmx2TSM52
WdWbPhBt70rjPkEN8Ip8+Xwk+YJfUqn8C8U4MDrKvJy+LNZUOjSg0vgkARG2O8hg
hzXg6tL2yVgB/ozU1Jft6axh3/GgrwRY1TYVzYbQR0KKS58sR49qyDCc9RX2wqpc
ptx+k9RM8XhXBafRwOqgkV5nmFQzm95W54MisrDiqfK6p6kAGKqUW+v6KSwwkLBH
Gou6uThkxooz9sL3RPlGAZ6j7vGo7ANZkqymGaAnm2RpR3TlCJ1QWmp3DG9CG+pl
cJOpPp/b+ZNep0Jpgky//GkXJR/pfDSkwJs7fZu8dvjp4n5/OlN2CTAuqVZXIvyr
t1yoZH/gzbG0+/wU2zMSQP1rIDMmmNsHPc2qaKSUcFHX974M0WMEFk9clMrxwW12
yeVT7wL/p6DzOf6Fn81BDIqaco5aIBv0ItICQ2VTqCIJ1QSzj35EupIvJYbiS5GZ
fKGW6VGEJ2n9Sfje2n0nwiXQFn6ysn+rjPV1SxarBiu5WnUrQIHMh7nQFZ9NNGC9
f/x9Vc81iboEiuB32CJgOOP8V7BpXxZLmxtDCDo/vlM2qNAASvgwR553tpIEpepG
zA/XWNMxl2+hfkCy6KOsup7l5M9TGj0bc4S7UM0AOlYpeGtZfnbMvzsrcyPsO4sz
IsOYJ5tlF5bCw+4vQQqZvjoVdN/FSmfTOlyKGPVFkMONKrApLJWfNt0fcBU6gm8M
R618XjJoQJfAKFSQB2cJGrIhBweZ/5KDaiuDLTvQQGQ265+TRDD/ndBKErLqQYjy
Z60YpGP7Y1qzAiG8o2fzl9BU8s0gIr3d/C5G2WhsISO1UpKfvJw2K4aeCbnFw2Xx
9E9F0fb1rwjeGTCWJEs5fuOQaoCgYJpwU7Gs61rPevfIYl9tlt6O1fTIf4Mfltvy
3b8on7jxt1Wif2TLIli03b229C9iRte6ZATtrO4grmCaswf1IlZ4WldJyTbBNvBp
tk3uoHa/xpDdW7F8kqG5IlREITOcBgS7EPPSZsF7Ye5d/WoeLXTUXPZDAjNfDvrB
WeN/cJSOy79oE/RBsUPkcMvMQFubVt3Uo86qUnrd/pWuHTfq2NBR1cpZcAbeWS/C
LV+EdI0096jN1Z1Hewoopymtbd3rq52g5r7UEPj0RVOw38IGpYiJBpS4ORIJ84R3
cPAkrBe1JfcwbnLtxxYhhqPjEw0hZAedIB6pbg3HZq3tHEBk+nY6FUvhGeqeFCi1
j7TPlnrs3BikkGumcKEyOQ+eOCtsw5EPcp3yWCN+Fp26dfc4SsAipyf4MT/ufUOC
/Upk4wm0BRulpkAWhhmmyoDTSU56Visrf8JGlvkdhFRMpH4v1n88cuF5Rv7IlYL1
qizW/XVbf+/cn1/JozrLczLWjKVdsYFPnlcGZIHkHpB6ju7YlG69t4D+YDd9/xo7
QYl2Q1agQVr24538aNLjioKSoiczsLoPUp1Y9akOU6fBgodUh8pfJKU65If9kmGo
Zi8Y2D9yESPs6tu3+r2IFWzF+wnhAIh2O8UZA1awYj6oS2xzuvgtX3/nai9AsMO5
nMifKWA337LRCVwyKN0mByWJmHzvOaQdQBn2awA61n2aPzwQcECcZW9R+n5wO8Ov
uvdNLxgaWmitcbhAFhNs1r84WFYe6GbddLYrElCu+2hHb/aG0R/sOLfSBLlrbkzB
SkiqceTh7Bc5x/TCo1k1rgreUEOSKw/Rkj1FXf1cBg9NHvSv2DYdM4cf6ZCGdZI9
zpcMvT356DRYenfdPiDu/7LPbfDxONIL0H9DkNio69fpWbPudatLYXQtwtBG3ewj
F9oMKVqr6CPc/bcaGCWYxk7628TUHsispmnuVHvUzvf6sRF3WUMxh/icx0a/x/86
lqZyb3uy/RtjiBA+twuKiut/PIyM4HPKOZ6zzjFlGp/PJsfsrVnQnBKPVrAF6s5+
L/lhoQkAmL+5YdMejkqa5pV/jkxfW5+W7eEsufyu/iLYfHh/kZkDyDf6OaOXndl0
nf0rs2mdUlGNo998dTr1kBRRvdbb7inlca6u5ELfHR+EjavgrrWfb8FJV5dJJs8x
VzwupuA4xFGB8ZjaULy7UzyoYEQkpl8p2aU3HQQzYtJ8OsOmOM+6SUfWOpMSzVw/
f2pP0d79Z6k2S4Ifcz8h0KxKN7rxo9Wl02SNAnM2t3nPEXUHO6jsCn+WrXz5+RTi
9rfD1S6ug+NNj5X4Lp0oPF4s+Ij1LLJgYM8Y7L41pWHpOjA4JR1h4oICGdDWqRu2
b7I5EB7iplcB8ZxMacrpP+8bfBewMYoEcTlIJONNKF7snqvcAbcIrAUYt7RY9Riy
lWZbacB8aHesBiGKmx8no6zj8RgtQ5BpChmrm7lG46Pa892vNe+uFAhxmhOgb8G9
Dn6o8QyaejJEWTVYcESWt7nANCsgR3+BAIQq9R5VbxsE3Y9QzjtPNJDr8ylXjMaO
oLUaSTDq8e0vCX4Np9sF3jTd3A8YTy40tMEgDwAZlc93KepcvNvQ+vBJ6XvPiZqo
d16c7R1TqXHJd6TSARuzgYIBKGEgorEj2pzBbNV6YbRGNldTkldPNhpGGTJIW0Sk
p+A7j6VkUKVJiG4E1Sa8N5rq9ex/FUWEPuAOWDIU3+yrRBOOr6JVGJkt73KuSBBv
i90qOFurwaNvDwQqO3bgLqC2h0WjmQXDw7zOBSWk5KCyRWmX8B/ShANb5l1VOQFe
7uTd9Nzlwh6ENIrOMhPbjaiOriLokDP1qWLYWWSCKpupC5Jg4Qe7APjc+MdmjR7Z
HGU7MyV9vjy/Q6E6/Isg+qqFTy+cUwGYpA0GvXPQ//h78xqn9uV/V4IlnUHcjBIC
QPu585MQGgjzOGRXVQ7XE2qIavGDXO3ybGlectDawIi/JrNaThmUpDKEMJqyN4zy
LKlnY0bXVACj6JVMyx5PMdZ6XFfsT7rTDVxQMQ/BKQ4hfvV8G0LFcDf2//yV6mzq
rUV24AyLvrDl/d0EUOr1yYkGHvTBsWBiVoMBN28Vvr+buWjqBgPIFkB3vqA82zVU
PqL0o+AaONwthne+T9exeexWRDXF9HGeIIUu5xWs4d7GeK8I3ySPnvvOMMhCqRou
esCon55dkTcW5J+U6pO1Bf8NZ8UdI4WxLnbcLzeiCKJVXvRalSc84qfcsnlE0xzX
g07GMJCGriK55PjutmoSmYmqMh4UCflNWo4+dRZsKuajfreC4SdCpYSmuKM4qco/
Z5qI8D2LQG2jDbTqarW5C+K0sllUU99ABQP7eLC69ptbtjx3aYTGIcu9COyVXm3z
9lZDSlpA2/qkgWlvdislpqm88E9J8rrF2XiZ2NfZPT5ZZLs9M0qEueLfkrPjhVs5
SjFfDMT0irDPqoSonVseWVzEicsHwDS6R3UTPH5Chhz748C3xRmGg/s9RFDPYYk2
MWeqTkYXaqJ6e6vWoPnTK8ECGw1mLqVpJ2a8NZ+97EvOVYMd0lX9Jo98HxUHIXQX
Y9Z2BJ3UtQT61m1fXx4pC+da3L07F/muRtpxiJIhCAdnJeKLPWqr6pSNdEUYZdlw
p4rhhScW/IA6lKfiEnuerTPnb4uYqHQLfjei4p0BZxuY8vrLUmKBX+Wf+1XRsVRc
fp4/7kq3+bwJTnlQlycwcenSl+wuV2CvThU8AjmrAWf4hpV3bhFTAciLgWP9OKgw
6Sx8PtXcKbRBsbi19YdJtK2igTzPoOIuvGxg6xCSDWkxujYgtAfWtJUkuYIF+LQ5
z3taJHkF4QWnxUgwXC2rlPzbkUm+ZMUC3crf1Sre/c5hqFnGroB+OsParYCRczAa
B3/l18+UlEJB20fgzRgkMXuWy2jeq7wmQz7sG+tqhxgIcQF28ZYUBxgtu+K+tDBk
DJzx9WpEysNYWMN+QSzZ9tgkZrBX+DFRXgxU5GAFFlOTzJ2wzF3TDbGdUECxFn15
nCfiNgTX/kopMx+LFrUXYUR31RgyPDfrYSixEV2Varswwn6pmJyN36N/HYkBcUYI
xi5Zm/OXIp9VZAHiqoRsNzDGi1kEi9S2HQQ5zf7cqTdBKrDC+yj4PNarA7AEC3XK
FFdnLvIcizN4AcHmHfX+xZoMyN4/EZKRuQOWmjgc+hUEBsaCAMOuFCqvb4AoYdjJ
icqchFs8KxMCqLYR/8LedJ5ZIdcEwTZU7nqoQ1CYKybtc5k+UqebwrkAYfAf/oVj
3OGp8b7qtNIKUE4gVQm3AUIHTonCsXQp1aku1cUqP4OKWw8CKL8s4thhiSebUGtG
Qwhwu9RgVGUtnFIRc3cLd6OhMmVecCyko3X+LGhOINoUE4dO0UtzmbXB+EhuX11N
tPkXkz95Q5KSmxEWkSoKvNplmEomc6oKgb7i5pD4kkPgzZagCzRbtZTXM+Anmcni
pOHYMUNlSOZyI94L+RhrCQDuFe6OH3tklh3Xum7zsOcJrlkHk5NUGoDkNa3gUAeE
kNFkiaLUM2paKeJE/6W5+/pNiUB1fj7gRuSDVfAI4lieluFLWY+yzX2ez3k8Fx5z
F6PWiwJulqMQt8HqVoeWH7zNTsRrFESPLnCoHTtlBAIS1zEXAxkNKFoy8IYi2sbO
cxs0L8fQedT0FIxPMEIzZtRsgDRX9NPFSyCDaBR2+xHX2OzTxrr3YsGv392Fbz/b
gcbZvI/nI9/pCbl2lw+EyrNJhlCwCAvdSLuATlhieYgP9twX7Cl/j/kJ3/xKN8Fw
YyGUSLnK8BECEZAhbgSotGUTXOqjb+3Mdvf1v7GK6Qeby3Ep/0mlHmMWp2iL71Hd
WGDBtt/xoN2jm/FdHbHe+M7JycHIsOSNb6XZnv9sIiwvYnqQtVnFCgITlbRzP761
jAcC31EU2i3MbNLe84vPdj8hnNTY3KcC0MZwRvNejlH1NwZ72vKn+lOops2+Mo6Q
vgBFs1r7550PI2MykgUIjR3IqBVzNZbrLUvEopOIgUgDHcqSuvCC+1ZgqDhnY3OQ
1s8jbWvf4TiSS+Fu1n3Sps/U+Mu0gVxJfNTHKl3yIshGZJW8BvwaC3ARycCo5H9S
RUGbbRrtK0oTSc23o32w8FW65InCcsxnriX6t+CAfXLzHjcWSDMEH5HgToOpIIA9
gtU/kqV654lVz9FjSZgvJpHeoLroV5tGF0lnTEsI6LqUsAdIhll1FB9R00NgaPDg
vr+k5mv4QD6iKdmgcDGmFmL2zz2RHBEmWCKARsXy8L+hDeSseCAjOOXERdpTfFPI
vsY/8oEzZ6BLYa1eeA3+bXPQdSe7ZUGJ1vxrYKljo1POmsTnfGHOt1jkZ/TcuETY
EpirIlT5v6OZeBuAG80JDyHhuNSLHwsOJiAyfc+V1iUBbUZ6hgeCrf4Y/QZTh/Ro
JJxdooljnKQ67COiO75DvW8laYX/b/PkFlW8eNAKoKM+N4tZNQlK0BxmAWF91YLe
vv8pN8/RsfzfVVN9KmMtydDjF0i2aOsIYNfh/YrinE63PX80EuQumKlrnLm5HzxH
sSDDaI3iKm7lum4k9Hkr5WzAME4Y44/jgSVcHiOuGBUCmxNH5ehPvaqSq8iWkSwA
4VihOIt7qJMKaoEXDtNI27U9+2AN2DqXS6jshsG5IZjqp9Aa6K0p7SMXAf2WO+/T
+7Py3f4DFxCs0eO9KJvGzfds8VHv8zVbLiAXXHbRAztyB6l59uXsnRTTVU9j+MKZ
AF+FiZxgk3RmupNxmuDdk2UVj2U8RQG+XwBVwTcTjuZRjEzrukSMBbFCuSyuBT7h
B4RgVIhgYdWI/Rdw6W0eOpnHkCd/MPLnYWm23mIgFZuPiTSblT2f7DXjPymQDbCE
SOKnC4WSQ7d0e2/c/i4+gwZM3qIlwUVkriKiLUI9dk7+HAMw3Tu2K+HsPCDHIFez
eBqM7shYno41GjCpojUsSlsYag+AYWB73xZ8V8E3rZ0gomDB9SUggl7Sx3qYfixq
ocerd30Tc4ToZlPC1bsyIDc0qatUY7pCTW7F1cvohWlFMB0oxuFMhn/7UbaklREx
/tein8ouv16lqM0UyMU4Fg8QM/zhM1JBMPOYDtYUlcerjzQI9Qfz5DxwERt1zzT9
sU4Ckgm85/2r1lmzg8QxGb21XFbwpZ59FiQKNdez6vDT52VSa/06DLkazCA5edAq
g+PBYwDphDcJu5cU/K0kcvSMSSt7QCVXN26DmzFSaZb/8ng1b8Pt4XVzaxVlZHy6
whKTvv1shrgXEvsPuFX758k0XgEowZL9GA5N6wVeILMFJzXaV/MTaO4qy7KUTzMJ
6J17TnRbirirjxMnb1xIgQqru+I8d/xZPsSNGaVdklc6TjFhVx9MjHALROr1hOcm
8paVni8PpIrjmx9MdE1wVpF47sGzMGtySWzW2k+zhwLSxUJdafv58/+2W/4wleLY
mGHj9G48aAbHt8C/eI7f2A7KcT8IPKDEyxD+bMrBhuLtXwyWUquyScewLesvu+7u
OcCgf/12U9YjrKTKynu/odyycPaCYagbbsK8G+V/xa5Yz65NAXa1hZYD2T8TzWnd
Pe5ZlSMKhQO8pLNyJD50EVYMFYFeGxDatpU939Vqv+B1Ixb5TIoGT3A3+iWanyB5
6k2p1Eul1C8xEKWkwMNmPIOtLU8BBpzu9RrAnCBpBo8mZw7V3MWLQyF5WlmEGhXF
7JaZP+5KZ/rxjBsXNxJrVMhEFjD134T1D7oKzGMzrMZdnLd2zfPE+omG2flpBkLk
q1C5YVHXnHhumCRWNiNB5Cz672oeO38sCWrURotOffGDHd3mDOj2zUDR5hpfEkjM
DLHoY4YBOtzZvelPcMDMAJj3cYilmnUXoDkRmGciUx36nAOboeDsUgBm7V1rCVbG
+AqwBykg8IUO083lrcBVUxopK29k5hte7pBap4A3pTVJvLPFAlYuLkyptJ2fbos+
UNwoEPE/iG6mguUHPbXatHQ97C1d6GpnoHtF69/ofP1iFOP06C9fjbQrlkbXjYJk
mheOQ52LO9XkadPsRU1MAaVrgqI8i47Lyr7mqQGeB/izdFZJvK+uhc5vzQdftSvG
Fmj7TxzrIfB4HVMRImc14QlyGOujxBRDS3/hl5/sIinD4uFlnjtb0fvDMTeo69nj
ucuU4OR3yvCTufSMWIHE4ZAYut9Gzdry7iNawCPVZJ61y2RZEky44b1am0UEY/WS
NWxB1xfGNNDG+K8YD3alZK87YWRIHJFpjXE1FBb1u8cjNeS57Fln1VRVMHmBCWhg
/J/uRSPoJBP/aEaqXRSwOd+i4dLv9lse0D3tjtPVLV9MV2LWb9kFp4HntzhXBHnb
lIHR3V7lwLK43IZlrUtnkEITq05UfLOVKOMAQE8hLW0/7V412Ie4b1GYvhBzbPEy
GbLmWNqZcgrOHlRjl2pYGO+fYuiybEYVDQNOppxoIWtn+DrhVT2FLCbldwbZv6uj
EFXHCaWg7h0MCl8epbE0+r2eIMFPTzklf7hur9HxfgSxSNyi49cU2nXqMaFuaP6J
l078abcxiZN4R9GkV7cOUh+0wFlDFqzFG8fKUu1o5KuMxA/LAJRAuTaTvoyFC3E/
1dWX0Yubl7GMiZkobMzZ2GN968ddLFE7NPu4YO0s0sAJo4nvapApCET28DPaWR9t
P//b38O7yzeN59HgnkqOCkoRSdbfV2XRtwPbsWJARffktDzd/R4/beO05wb8fIdB
UYlDFRdC1yeqmmi0a8w+m+elxCqm/atv+kHznwlzhU6+as+5tdrL9r1Iz3Xrtlx6
eajnu0550XBxoPPHSL3Q2ZbXetCZSLpjtDwcY0tjLjRIugaJlquPBBE8iwCE+IqZ
q3NaY8ytgj1j4Y8xTbVrpf02hOk62M9R8SOVUejqoKYOLh/+UeR2rovLpzA0MWOw
5PVw++8eXrlwN9YBqW1ExZxTmdqLJbCVSD5Int//wu/vAbdFuoeAOMOLLX/9mM8x
/vRhMILIL4cn5eKPCkfXKhBjJkhVNseY5oc9f1QzxeKDVPRRj9mIJGUqtf5fD8yi
fZ7KEFxDORFgTJbXUHTLLxoOCGwHsl+dGXqyeErL4AHM9q6rCmE3ZWF3+JSC/40U
/xRqQUpn8Tbaqw3HIgbZwBC7uR40LQ03u0UBEPRozmNYS2qsOut6ToxdWecx31f8
7qpRZxXjjNvZG8r/I1Ro2EaYinPk28IggUCbcAKlcSfcoCGUyepQkovrY1rrand2
v/E9aRhZHXyFGdy7mwnHXWcj/G0q9A85dPCZcs9VQ4hAnndq7YuWS1laBZzFEWhq
gXYAgNmOqHNVT0fC89orjQPYg23lkMG1kVHFiWfK+QUrLGCBlKM88WaeAcQTTqN7
Ck0EJFU1gyoOBGOgmFQ9wSbUqwadk3qGdyaLG6Y12fBDtzLTBEmzOiBv3PUgdSET
/HbSd0RNho8K0urC2uZ3H29rJAsaKG6cB99Kq2oQfZcparwGNDiQJdCJo5N9/mg8
0pTz5M7cGS42AudGgsHc8rZVZzhistIPXOAstKVmZN9ItrO3M+4R1qW7QKR9gaPG
OpFpbLE8NhbqaKJBiR/WeLrI6ECrP7hGGyEoE7NqOV7ewon0BjrOsfX9FEbRno/3
/2IxZss6pwFF9RJtV4IY2LU9yu3LvWCUGo2BrsgrU2wkcbwdsMRw3bCKc/nCP/cl
H/WddULmtulaeTmJnn1NFzadF9id1ZrPQQGppGFH1k90p2cxf2FV+oJTkjnXdHWC
dcB5kIJCDZEZhXcGSkNwu5Hgfvqrat6j8LSfgrPVMQytcTPslb0BFLLr5ivrKqna
TaVZJjxalReuf1Dhra15oxTnptCAVWdrEClitkSF39CwWl8WSGNkx71/RGkGUjQ7
wI716M9SiyLu9kEVyKBeCDTeEd9iBPl6J2vMoTs7Om8ooIKL8gfcoOoFRbMT+yHh
Zx+7LyDXzQpotJTTAem4durdR/wC4la7LiJ+kGewLW6oN/Q1O6QxAEFO4Q+ZlS6l
fjfyjoNIzEf+mxvrPsuuDQMNzF33ouutheQySUipJCG6rJkkLaHghAHKxwzJkwvH
lZ5E6lavdvyogjsvS5TCO5RAMYqGUJQxbJX6rRBWRbrzM/zev6UIWkzwhUStliLs
UiwUn+mz3k+NUQnkpaKR+6L0SzQruqObNrGHqsoFWKa9V850gJucGVjfKEAEuHfL
RvzkupXE5LQ/G8KUiEa0UD6UJXOyuBsL7Or88jIT0TxLSLcczINhJEbKQJwHtnQY
TBhXQxpWeIRaK2FM71o9j6FTJSTLF7c0QAVDBKuGgROaklHrQ49LaXdp1RtqV/GV
PeCoJkr+5lR2owXYf5QRGsB87FPNPdxcnx+iLEMyxkB1B2sDyFrN8egxd3Spv0zF
Zc7gu3k+o/odxotGDAPD7AwAoMt1CdQBi7DrJ1QHGZinzJSO27w6YqUoGbAZsVDT
y/uJCdImJsiPvw2zheKVCS967ob57ludiE8CXpfF9ouy/ASBsVaoiK9/GFrVubZW
4cRW1kaoPVLRwRFAK11WK71vArGJ/ICRjmk3vysbaVRBVw9aWeRvvTnhcC0naWwZ
666jpErcf7nvMOPMl5T18oVAo26okcxm3JxxsiwZw2einVlXlGqdDzlqhBNUkYHn
iG0El/fGTL5VMn3f4+JY5Ib5vRkj83slvJPijXQMGIpdCVqWB1vbuGwzvfLWl9IS
b6SkpbgtWyJyeavCj9AZDag5NKRS3ktYrM7C9v2BwunXzB6ziAjcVe/+cIBnfNvv
F1ykhCSo6gaNxbTqNm4sMyae479Xjmmzl+X3/DypM3Q/ZAi1jpYckhmdsiWdpcGe
sPpMDFMoC8AzQ9UyzOzApvMeIGEie02QAgHiqvYfqQPN6+pxgT2HFYIwbqLVgvB5
dBccjVyTA7jyqiNo+WFp6pE2oGgcUPqox3pd5s4sRae74oSR6yqH7TIk4KCU454Y
Xpzo3CkoDDyCU5WX6gxOGD4KdnwW9xTt9Ole9CmcNH+C9nNSIdBwdnX5l6L1/b6n
pSR4owNZR2YnEVNsz2j7iu47bV+G9cxw7DjYyVV1HqJ2PaEZOAiZUduad1EXxJ2b
JspwGWxwSZ5PZIejmWXq/1NnBIgoMLCdlgNrylCfsptfhgvULXAdvM4zP3i/0SdK
/FLRCIVeafjQlvNuqNcd6GTL1grLnqx6kxnp23nxlvPoYh0vpvDh9bM1KTKvRJ/F
9n48w7yzX7ojCB7+oqh1W7kV1/eTOf/pXUgUsIxeeWjlp7FgXnBR3qZIDn3huHKB
GQoiCNILgbA2qqiKdHVEBiB3STwKoX/oTYZeoMoWbr4ybVWGbyFwlpMtNbs/fuUn
lvLtY5GAEQW4YW43eNocxdLpHOmOGtkYa7gwHFhY5eD3xWU7LVn3BreTy+KQYP1/
nKKzjDlpPBQhDEAFg1mIAr/AseBnYjALtlgHRpbo649Q6Vss1Ci+cq1SyQFlYeH9
yKZLTb42scP23MAW61hCvSDbFRSPJL/rrKbm7qaZShpedjXv63wi44omu4QMWkU1
fPJpvADPAnPDH6scIc9quGafnIbG8PmuxREWnL9e6JVrSNSvHqvrvaxPiNGqMf8G
lBhVyiMy/Kl2/72eciPYxib/+e0Wo20oOnju5fabPeW7m8H02EixSdurJdyMVKB5
t1ulAbfEenYoCROBlF/ak+4OOgy7m9paWZA4mr/YaFWFie0gfkDGVXsX/DPBjilj
BrFxNsVXKDpyhmXNLr35gFXUVGkm56FyjxZCdidRuynf2sT5F5J6hOmXdtdujs98
T7P6JSUFPhrvOQTsxOVEsAYK7dTQRLSuedwcFBrfBX60sfeYEGARZCi9C9vomgJZ
B+ChCCvS9txZf3mwoh/ns4mVHSXAR55d9XN/mmynuBKYtz3Pqo2BcsVubDuwSupY
mlw3n7yr2F1vpEq36EK/r3Ua2pfchrbDDuKaFClG4CaIW5U7u4BfnLTjFCpGkjbB
ek13H56b6QTFoQlZo+u/ib5VlyQUyURw1GiIy13DOfjhS9es9Thu63Ne7O52+VAh
d+SsWBG2suco9JwBzWQAY1/wrneHst1V060HWI+YBx4oswXVtGW+Lfc1d+oiv2IB
mnmHM6jtDTl9leESpQEGIcDgjQt07SLH0KcJknHXdhRonwDFVRlfUHv5hSuNHiju
pXsfrpXRM9xwTc8CT43RecFo+B3zuAGorl1zs+6cMFZIuN0oYc8bFPlzkU6r1Mm6
La8fHyZSvSUzZpmAATMwTRNuiXq8UCZwAJAEbiUwMTGSBg9JOdzV8M3g9bkwV1m+
LBLJ5xPH1iFkRTZ6GEFu4XqQ0V1DcxoAume/7pbMh2lwgVi+qobB0GiQu70Ii0oj
IhJjkmvUSVukwthjDxTfS8bTCc688BkmsOl+6ejE+D0dl60w+X5tdiD+zGHWbw5L
yRYrbojCnuAaJRfZgKJN/g4ovuWeRex46Fzg+o7dPzp/7CWQCVPOSQZqbYg24zMx
KAf1nVo3UT43+uOelO8sYPv1t9Sn7vgp8R0T7qT92mmvv00jfw+WuHqzt31VITSf
x850l2cAZWJO+M90CLiz54itoJVtXCpZLmEH8vFWDx/dJePHScZDIQiz2DwohgxM
gKhg+YR0Cs2IyLsOm5BDgeZnB++xVDPfvmJsxdKamBzK5fw8sPIqQJpnml4EVGUt
kd3t0sGk8cknNMqdq/LV5MLqYH5yJFvygddu6DpdIA3zAkHiCDznmSTvnOnobyJm
jmpZY1hh1Zer5SpWx4cvmDKkp8gVoWP486Wy9vOAGGd+tz0usuQ3n8Ln5Uxvev4i
VBwfGPT22AaqgklgvQd8nlXgUwBMxnIJI1VSMEWxrCfHqwsg5PjzvS0whjf3HjYZ
0xfuZZXvtG7WT0QI2ozrpjgCvq1M8J4ZNurr4JnaPtLdtCBcVzId8HZ89kWzrh+U
ofFR3MWshzCbbiDk+lk6bAOiQVIwR6tLnNU3NyjFJoYcn8wksC+wWkvSRv5JPc7Q
ReuBcBBo5Bp97h4eJdYp6vAQOHzMdXzDUQ9I4vOiYE+ZnQr5DhTqXZN1tdmRNNm2
q52yKOk3sqmy1Vsv9FVp7zJbyCie//BAaSHxWN1Ss52O2J4zQE5l/EGKIl4tIl61
Rsc/ciAqFvrcaAY1Du64ZF5pZ7o+L7WxsZ1IkAt2ht09jsoNagJ1BeQNdCWQ3BEw
ZkdzhgVuRfOJ6DzpkAsgKRlCBDu/z/W+5j/azJpxZ4vBTUN3QxyhMfqJuxUHgcON
mRPtepLqsvwdVfQaoNeu6m4qFOdUUmJxDb6g+hB/syDj5KBUW4CSvMphGRFakBbj
2TyD7e8jA741HVjK03sK7f//53sTAq5eXla6oexJfb1SegW2fDzc/XWLZ9+fwcVr
d8TiYaf4rr6VbtJ+gZbKJJ/AYWt+UniobO5DFOViRdVLM49/1w1e06k9AyW2u02m
vullZB3DXT+7rScLYyaM2DorAhqkpiutYXVD6OHMbTiOTmK9TWyoLbkjjKRtOGzm
duH6bemCOt/KRlBTrIV628v5WlRqk6I2HKJxHbbZEWtwHNgAa38sZWSxr0RnkMyJ
gMY3k5nRYj0Pqptiu4+8lbRrFTOQz1PY5dIWYWZqM/EdIO2ngLbFozBDlxZ+rwdS
KR1i9hKdQPXwuBXgpeu9B4+CDmLhv0tW9i7IqIASso2lqssX4VR6Ngaodt+G1w/w
ftG5iLKzxkqIwSlKOnHVcEhBMY9uvWZtWNsg2xjDMG8ytNgN+88jA/CRCzw/6158
NVou61O9Gc/pZqAoURBXvZ61DXqlBqtZhLjo63LNwhOWGl+kG31ePAC2uRxEsdnS
l8k4Vu2xEqQMxfe5eeDcfqK1drOtmiDziChTfG5DkwjfpJj6AmeaIPqq/PcEsRi+
dyNfP/4Owla+X6XUQQcVpNmwQhIuBmnxwctdO/88+rOsI0M6ulqY/JRnqpNMspVT
Gh1ZapXxlsUhz2vVkZXfN/GSS/ghxWsLuQJCYSSKuL7dbORzIbGTqrcgdtDEekqs
CYRD7nSkLqd7Olg4lcKocHaKemHIyRdKnW9imKNNbnh0dtJEtLMoSY0WN/4t66xC
0/+o1ImvTBSzXEFaMroQ8SE+lXo49Bsjx7Occ88yK1kjAmqtipAnuc8dSvboIH+e
m9B6ozouxwXFoFFdjEsgnqEvHR5tGhsUgdFa6ib8uvqjCpdxHYnNA1mly/cb9JA/
Bl/sCDeSWERlxsUxH73bH9JfG6TCPLqCdUaVfq+ZU3NjY6tMpj+mVIMRRpyZKOX4
u7Lxa4Ml9EPOXaRrHrCuTgYFFCup4CNfZyLbXhsglPRKYbg+tiMWSJVNRdRUng2H
eIW727V9XGb1xgxgXnUWgVQxDgiZ9GOWauENcq0TYDuJdNwbgCT1DBYhiSG3kd2S
oNhPJJayomxEhBqgrWb/acrafMCN3eVEy7tDxoz5izBjq/ALVqhS1pBRI95BrNBy
+toI334fWqHiyZXMLc0eWkB1cHGwqDGb3eOBrL/7Ev7z0q5w6vOr7P3m3bnJfIGC
MHOH+NKoA1Yb4OQW9Qy36DunOtd9xeI+OQoU5rEbsNowOI9Sf5K7KStSYeXJYIQ5
cEnqc48Twnw3hVirAWf+96ZBTXtaZaer+l/iLWHSkcrbnW6qL0zk6YbuMpVDOBsl
WFmpN9U9u8MZVLBNv9Myr+2A1P8Bh2kAgrdc7resqzEDhBPvsOaMGtQwDSflhYFf
tBejkb7UZ86KqzsU3nk9etjF1+9tB53R0ZaSzriR+TybqnVNQoWMqYyv0LuqL3Bl
3TQbsRocISTG78v6qLZFrcrTfg0f+HG1i+yzf/VeMhXN3qkMvFKJE1KSOro0gmkU
K/A8nYE4xks5ga1ocQW/1TkKcPf62GUVjRjRBq8YzgU34eLfZUaBYVuO3+LOeQV9
cPeCI0HAML0ZgVL1crYajl4sXx7lFSfsqfHGzRLgQfz79cfDSKgpvptsISEDohx1
Of6+KKL7qbqf5/kDysKFJMMz4K66CDUy9trHqTVu4a3bg/YLS3GIhd0xaZtzhdqA
JP5XD1zgohnZ3bEUPe+t7+ID7YfJaO1/qywaE4fepgl3Uk9mh5S1S+f/rCW37WRu
cRaRWudGR0BkwO57B8Hq/qP8u+i7EVJuU6J37LtxAzl0wrQQtP1rRR9Z/nIC5Jts
vaRMOUmgQuQ/1bJ6rsUbc9gaSBKr6L5dJGk6XW9p65teV39kvZqqstO5qpzQF/N7
f4L2+C/vVWLKfQdVl/DBELG/L+pqILiOKGO9mwCd6EceqdM+6peSWelgSooc4c1/
vsS0yMOYguxHDdMzUeLQibH0pMVylOcWJm78U7JGomnlhG9CwEHby9J1lw0AWIIh
+D1Jj5TkdNjcu4TSq7JxbBJlPex7Zk/dm5TfMIvzZtt5QfmXWzGGF/PsoJVcLkS/
jstwNXoTgSAyioCngin8YAG67Eo8seXSHoF708LC9EK/lZj/jCNWNIZJa5iUgma8
UdxMNCyCu23OAmExvTNfJu1pAAPxi9lYGYKUoD4u1O+XOu83C4fp6S+GFjz4V0Ms
iusmS47bFyPozhldDTNHSSV63knGLE+oGgTartJUdTDUEF2Kp4oMoxkXEd8KLJxx
qYWVvgGkknTkTg5aa04v84ljCgch2JH5sLUkGBTb/ESM9kNG8ZcZv5IyhLN2QpVn
RpTderXhjjnrelazWlNYJkvEhNMV8A5KRY8XkSOYSFukB9DBFSOe6gVmEvGyassX
YqMfszI99XVLQB3c8qJO+By7SqwbZwcVPCYHvo/cfnt0yMm5mSRxFvD0r7INeXyJ
GgisAByYvzVqSYo05bco0Yx4R8Xt1xzmi0DMmcOCd0Oa9kMSwUlsRv7cjO3VHths
3ekkqCpEhPcCAgJG+9z1rtnuOVXAxegWp5VDbaWkKAP5W+ReqcwenpWUKjbfa+4S
wK9JEOYv94uRpRLttjzjmhCSC2gUmdSSP7fLfamahBu2UQifQvHkvWcwSUOG5vLP
xlbhgDWRctg1wfq+BjFdF3WIp32Oli1fYqK/bg/+T4+/SZTqdm3uFSYpAWpAnMxc
8ggQAmnXqVC5mq4jUSDE3KZiIksJ6MauoC3iPrfwfj5dTrxqMH0hzCetaitDM0nb
b+1xBWz6Ml/R/q4shRiWgk/OWkchK0xdPcuuH5FaLIPitZEfytILrt8R64/h2YKP
vgS4FoK0NvdagrKoE9DQw9qxI3pXWbnB9+ASImQVrWBeAY/az8Oy6X/+g612P7jZ
OOOGsrm/NunKW4sF8nkfZoqiP/fxbLCzMAeUMGNYT3+MetoTTiLReWoPgaVLvFOE
VzBaqmuivNvq3kWxS903ZBfbc72ZS+wmmScKhbPhI9u6fZI/SI4Mk+DiSB8zG2vz
i7rV1NQ2E8PZtAfmLMRbDTaD+mPiKc//+UcvPp+5bpARnIZMWZAMPejVZK0pSLqJ
GEf5GuUzaYYAvFnfkA7NR6PjQfIa3ZQZpuzZ/6tQSiflsScQhbZSu6uPu9oN3T+E
swXxblqvNXYyY4LDOMyXfdNKW9gjFpwHHwOvg/ubuc03CKvftkB1mg9CgCz1+/xX
U28zvxRN97ZCpreCiC/8LcVI+kXHLOuhtqrYcplL1Dgw7rmF3S4Teb44XecCky/B
SgrqRjObEZ9vcmLvWO7sbvyilhWssEdG9YFJ3565T/0hZlTP8O4m5NIiQCcknEBz
iI5lHFetYrpYyjthOxGJP7oUcMItnYDQ7pot/KM6D2NeaMN1RTQXSuKB+GZU2/X8
yOMwNkeTnQ91/87RAg1ucjzt2JED8yZ+JphzoINMf72FYw3CnlZboJsN9ihCe1Yk
MVrrMSFDTN0Z9iMwwUJb5QSNg17vRo7GHQe5AuaqLMHyQxrFfCGhVCPosdWEtFvC
Oba97NosnU3yEK+LphhHlbS33voZWaOFAIMFDnuuCFj9Yb7FoHsVIADEz7fOeooc
tKnrAxu0VkfkyGkr4v1INT4JHN5kwJy0ExE/gd8ZhyCDIB+akpbUD/j4mm3QlCYB
qUn4vBGPgi8o/cUAeeVO0CZKqy26VwCKNyNHlwJGn12lUR+w+NBdAtUVOJpGEZkX
Nhl4gvhosOGGOAyZ8fmpTIeJDV5NFdC92faiYNupQkIHYkeODg6Dw/qto4tYG/eP
gJXLENTUSAGntHNUdQFEBBmTAr+UYAF1TX1/svQRZGxZdnYf24oMLvcuo4UVgXJ4
mqtmL13QoY+QcPWflz1t7nPMbVm2BuWeLxXWc7FN++2kvGVpCoJ7wMkMSCN6nT3E
wb+9CqDBhuwHdrpbszfbjwXN4hWH4U3rx/v+vuxFPbOV6Y9OMWC+c7Mn+B4w5oFJ
RMGhvoqd5QzIBlw4Wdt+/t7P53EU2IY5+Ft4/mNK8OZouEUZA5T0CHejLPXMBHLI
SKS1wEr/LHURFn5wY3ENFWCMXzPxOEopFL1b3V6zCeVIm8z8ArQy0iNAYUSRQW5W
ZqJz/U+YnRyNtS9UifumtgNakQ4QdTS2OOH+Yrg2MB/ed8on2CLgbYHfQQjNVJA7
r7Z895DYogRA/xn5RTpcyUaIXe+JF1CS1xBrKCpsXw5ppxNMwCIAYOzTwaDwCAhh
90J3jRS3P0nIEXYtmFkS2tLqAHGhbTSuAbIOALeuzvHoozsIBpxzL9C/GEqyQ/Qh
jLTuznA9QwbO05P+H4yBB1xO2WVAnxKMgDDmbwOATKx/urTBnBD4zwdlcyVIeV5V
qMjjnyRIrOdwzmnTASPGOomNIKR/13sWNjAOPqtp10L2hbiUShtH7xGbq0vxyqKL
u2AswVNwySZFbn3qxeb6mJUgg8aa2WF+pXxwEE7nMbj8Co+8SbvVWMoGE87N8WOc
XjhvYIDUhmFJI752Bs1F9cx3Hqom77sBwXe0tAQNkzhctCMe234SPRRNbQE47usM
ZqIi+qY0b7F4CkEjv/Guv2EOwDcOkveVH9PVZChTCKQrnGjOwDUvYGuI+y+YWB6z
xgUs6rAALohMkpYo2LLtXwPl0/5V7bHp86KpZ2PqEkaygVojK25GKLBWUd/WGKSs
rfMwgVKmBqtKiKSkWCqmpxYGg29utRj6WzS+E9APSePKtlT3MEBJwzCT3ZpPT7B4
mVABxlngUIyS1jKMwhFh+HD4y6jzmqVvIF7KgJ5CT+SCDO+69bxUx6i87rvC0pBx
SsvEwBVhyLFeuhdgrX4gFHCe5NlYPmylhLKQW20c3ey2zmXFAQsO5HggTzncyR1+
+YVXiAUN/ovutRfSjQJObmpvo2WQk3solmM6Ee4HcotatE458p/Bm7aPP5j3vBkT
XrgzC4BlvC3c1kzy2x0JY6YvPEHy3z8Za0iOxWteQKrVTsQJtbcY2+P3y8g9vr9k
FjcWsupHQsKbqovuOaYyVUeGZ3tVVg0fNAMp6akgwLYR3TGFBHBuXFfZAlCD2fOt
2KyHbbh9xgSACuMzQKCzypCvNrSXlpmeXmrH6j3YwoddnSJ8YsLPwsZuu9/kIOdP
8xwppA+GpM3+zdciGhZ+lk0ZuwYexxCzF0zZcCocZ3cbPDpvxt4N6p4BaZpjOXMh
tR/oxboTdyAoGOEnPfykeC4FfmCuPi5KUxPsgZoClbH06stbtjDhzpnohF8rBD6O
S9IGb3Dk5v+433dFoyHv1QyQr18sUHPpbaaMde1yagOKPl6HAWtbiHBOa+SF7WOq
7u4rT9ZXJ/tj9VFrVquO/ZEl2uu+8NOohX9AFs3yzz39Eb6Wgo+NWw/XS7Kdh+RB
IGTufWR+6awA1fwA1u+BPEoAn+bgnDjE/CsQXitbP558pRlU4g3XLGbYXoQ54ERL
tegJ1FKVKhabAKfEhunVQcmzSp26EILm7FJFPQfXz7RNV5M2Y6sLz+oetN9jk72g
M1xBZj9+BcvNrJS2wHLYdwLH4i5cO5YlHWGSxj0js1S4nUTPBfYvKB1FrEjBNw84
t7Pcn5JmlUuMSppIRiK5zerf2JGlMrslTShasrlLOLjHpym4MmxBKikrJMUw7Q4P
rhSBVyaveTtoDyYjCCflj8ab3foyXU7nS8lhEp2k1qIdRM5Clc12hEvnNhV/3cht
gKk1ky+EBLXORVwMGE2fqHpurKuyth+N+BUkRQNSxes9sPUI6rAkbwNLNAQndyT0
Y3u4e34nCzv84ch1ky+milBfkWIu8TJWd82VjpaTqZL2qrfc0QKMehluEET/8BVd
1bhelsKm1JUxrlHC1jUQWhUHavcFCUZQNGftjRJhOY49SmDe2YkmxYrBzv9PArnq
H/xfaWnzvCozRnX91HtmEHZOu5Crogv/T+iii+kQ+dTJV8LC/QNs4Y2HA66x1kxP
Z1IRE9olXLLldHX/xFh7bd4VBpjqaRaeWYuFI0tFv/6lwRV+roZIb8D/TP7YkKuw
GQKeSo92jeyHR0oI6a70DAkog4HMkgy86Fme7rmzhrhO6mx6vMjT923/kPaO+Wfu
OrlghVYItbcmChZd3dLhj+4U8Kkp+0wJcCwG7fJ+1xsx/2VQOKKttF/YtKThGuXR
6ARVZXBsUSw5FaKf2iT+i0kwN7iGM8SBGYQrcGbSp0FFgN5RHNH1BhMYzFN8GPZJ
gbzoQJ4DooJz/nAfHrGlV4+rNO91e48b72dK68VumqDw8SnPllZrKWkxdeF3Zlk2
yGTcVft1w5RnIy0gsQPnggy6eJ2U6vIMkSYVQwruzIZDchEP+7kMTiUesr44ZJ9C
Awftj8uqQY4xsgaMfmC29x/CFnKYrcaym2/P3u+R005OzY25bWmqoAYC+9ihteod
zvA9bwYNpreGd5KebTE/srbxkUKQfU60g6NRA+4MtvHTqdq0HRojJpx5KFwZlsf9
pdZyiuWYTfrVnc2cVC/y0cF+cl5l1xjXKYcXO+ar6gRayPj4C0m7C0NuFauJ/zZI
jhncv9YX/u28F+zvnfF1/0SL9WO5MEbHEN8v8PG8rsDdO8ViLvwbYZ/UVxe8Ntw4
ttUXqXxSoaiAMSbfuxeXhYLNowEjZ1BiRD21pzvKBgrzlfVJYfOktY3CCc+r8++M
TJHJMjSkPGyyyZE9wJkKDfcKdv/Nv1bgcrrMs0f1E/T0IFWPxhMuW7osRWA0qfy0
90PI1mO6KW0c1zS31dDjmdMyVOW+Hs87XdSGrK7CPYB5W4LgBxyK1CH4cC/2zlNR
5q2aPrRzVYPM5XeavyVFLzRgb6rwGbQCOgT5BJoayB0Fd1qAsPaij209DrcTsXkG
yvgMqHNvvAklZfRp9V5rMPN5Qi4XC1jIx7CqzHNL4xP7yF3MxpuncaP+v3zCHuNb
YbxFrrNLVLxH2CGjOCfDav0j1mnYMBTVoyTI7UKsDU3X3nhlLu8nzq+Pwy2YfJQv
NsSd3W41QNEHcLBTEgykfd0lVHDMpXV1gThL9k5AVLu7Je+cIqZIbDRYfItRrUoi
91QlrUv+D0afOeg2zhfibIz2We6rc6G8kUFlYbK9w3ZdB8CUgQlpHJRmSVvnnQLw
Pk1/i4WX3ztZjHzPt5IWqupQ9pYryFaZbCOA/n0HM8OjN56c1rTM5zIy3XnRm62M
8Ip+YbACpkd7OjahdRGtBPa7T9v3KM45X37CNuQ7d7VlR9lZr50dRW0+xFhGwEcN
wsXUTsiwSrBqouFD/l8pgMz13WeWjJTiZK7OLdNi5fxFF9IRVheF3dfdjF0Ju572
6t6ZHLrYaqQI0uwuMZMmU16KlCRR64kyEPKwroY8Q9Od+i8o08nl3uzIgxYdtg2b
XkmEIk2YU8TV/s3AXGtpg8t47SueF3XMQYmiL6EYTxv0BhVuUovXP6zDlxWyPZLK
PMWxbX8ERfoqthiSMmESnVFb9J8HCa2eixeryRZoJzP5lZFyBqvjoc1Sd1QvucDD
GKcwpmcyr50XLQrX9xrkbr17XZO85l8xZDYKtNIvhksniqmy/ry/FnH5p4buNr+M
DeGGcOcDtjOcgnFL4grDozcdgN5AJErbqw5byjogymIKyf9sOortHNI0xq9XhfQp
EHR/z3zEYQwaoglvPiCKmhssi61Ou9+MB/Fh2HX+rhzvue1uIuV1NvPuBWmpCYSN
ssdk2AIQRr/Teain0bZb9t2kbFBbZd9oemnVyk6Jw0yeUO5vzykg8IE9WMyyWT5J
RVnM4NnF+0Cr9071Pga89XJMJc+eCvmfzso9Lpl7Zag6QroOpF/QjLOw49W/6HzU
qnEmmEYpZZNFLsaGqyB7J4M+wUWoVlO+yW64xKuEAVTLeMAgDq+EnzRPb5EZBFpM
AVmA1qFNMkNtRcCXJgNpKbtV9JP54p86B/MyfESk3lqwGD8t91LRT1IwAnRLcWrn
ApdB+JH2CSHMWw5EIOumOtxWMQxai4lsTW4Y3J72UNZolWej/3gGpiq1/29P7+Hu
JBHdsDUJlPkVqhh0pK06YlLE5uQo+xto2fVQWjvDtw+AA7LM3P1mAyri6C3D6gHL
9aAPumfx9kxwgnZdKlcSfuA6EBk0RcCbzNGi7Rrg4s3ULyRComwI8qFFlyXznqeQ
oalTX/efPyOV39I0oZNRhkizcdgzTJRr/qJNDBshq16bvKXS9Svt+m48Bms96YGf
IkSLnjrbgMEXdU+0Ct/XU07I83pKYAc03zhe3+XSm7+a+GHuW19KryY3EThqhfH2
0i3ArYtyE/6m1uMgzoOH9DHZW6U71Am2pHFv7D23LmH9jkEF6mHbPkCykqnHmC4A
bqDAhPRCMJQN5guULWCkDPgoEo5YeYYFUf8id//WOMMXKmvvYYUAbww/DfwMzN9f
xy6PhP95cULKopu5BesmjskbFxpUIJt2+wiPxi7l8kOQ8bII5uFGHNwwK2ZAidjx
ZXQeNHu3ruC2WtlMZPCGoFbjazK2AFzYfNy4dlzlT9C/3tKH/BaR144KPgJyF1vJ
xDuwSBheVpyO1Q+SwgdJTt8i0wgNvATihrQM+BwgQ4GlcsUyDFykHGcCAGKqqveT
FwxVMGBMAdQ154pL1whNnjPwB9W4hvjPTDSRw2FnSqvdtz0qAegIc+EuVu3q1ioN
KnzxySSBgNHHTdt49yBf7KBl8UIFYm0OGu4pLGsSOxeVmymlO4EMuIIe6j+6c1TM
zkbr0HNJ+GOsLKyS8L0SwGTxXjb9Ca2lVsuWhAhM4UwqjjUE6OnpKYPKScM19be8
jfQdg5n6yEY65lw3e7MmU4mfgiMw1qXqXigm0s1WP01WXX8R7GwIyqIJXaAobJQS
g3Tprd0QzYiEnVeK8s48M1hPVGSO1xYTedJTjcJq2Rr7ONwrHSRXfbNvI/NW3a4Z
rrWc0CVVO7BBYhcpl5lAM4T54qcZVq5EbpY6vco77dwgwUsvw6AtsHj7kEujkDYI
aFhh65UL0AQDgw++yNCZnLB2czlG4C7dgsSUMeqBrF7vxek/PikBau9r0WeAi87O
m3ZLVDqQVitrpcWMN/rs5nwZGfNusRiTrtuCdEwa+jpaXHqS5CrUclojR9iJ8gf+
eHUY+YvZLRRlBmiBT9SUC0HXaDoh98NMGA1Ev/U9nu1F/7hxnDARJN49NC8Wu5Tb
f2Y81r9Zq04r6Lq7OgVEGKVgwKioiBUaBDV5ewVLa5a2xlOw6xE6FLrmtpHraWKL
+QSYAKtz/dH7JnXrAu6f1cOFz+AxtydSFip/kF4sdgcZlZ4tvNt+3fC9iD0auOhQ
lcwW2aLFTCZpMHlw7C+apAniloEi0XgjB8+Hpc0Epr1ibrWFIX7B2k+b9MkTYqNH
Zhrtox5Stg0US6wgZQi9SydZ48uQ87tsmaml762fSSgFb0YUHgnHgScquUR5+eGN
5UX0VZUhBYnBpymH280tZi/kjqzNSWqYV6TpcY9H4MAtcyaAwZUZczdbpMj4bNMF
5QXIfwQDtl6v15kKcBhaPjGROV8oSkEBxbPbkqGZCnIPEG1wVr6knD6Y9zE3krA1
xCEMWDy+BAeQI7ILRLvlDp45iRNrvftMRLEY2LDXLinCyY5L0EZfs5sgdyIseOZx
HWqdQttLc/y6WLN5xCyz2Rgb9ThOzbFNmBM+y4JjHDl88WKVNPDI3ZB7r2sYG5fb
g6WDCD/GRpgakXlOGStFZ/FiASkSbhd+ZNa+Qnd4CNATDcYfUdI4CF/5ZCnA9nb4
EDWazdI0Mbp6Rgtxdh+A4sL/ZQZ6n3gTDysQboyXeij+tvR0Je8Q1pcHwHpEd0a7
GY/bBZROl39fa7cx2qXdjTgh0F90DWltLQGRK+kX/FcVvPgtNw/JoIzfbt0gPCJz
TtS7V71yXyYRqMQnCGBpWsQ7XyxIz8zTar+WAxAJvMDUz3nQZvsCqmIGXwWisZhu
JcFUezpFJMz4Db+Df8jjooUi/fm6wmze4gInzlHfqblQXQgZ9hX/9WQ/T362WOef
KgV7BZSuvASnuSE4T7mpEjOOuTGLuB1qhwbmLYYI9RO1AKyOwC1/ImIW9V0yqGf+
PA7FLHuwqy1m0Bpf3B5YDDk5asqqB+pyYDmbqPashSK2u+fezUSF5Kcw03KqOANY
UlRFNG2QniVu8XPtY3pnPynCmGTwBv1+fVEAi2u09OuBfAn1HkTJITlEZ9Ftbea1
Bn2zppmjIT0P+NhXadQR17s2gaD+0vHkmH7xKX6T8uYaMPh0VkEl1hKGF7tZELVQ
YC39tMhbDIuwYifDAoHuAGHxjLfF/6rIlmFmv+714cUe11+ldkhPVFLemj3vV9a9
fHmKKjW/eFB/IGDtt2QYOLXup24TSKujYiuc192UJ8tvzGatyAg6Zcn+vLpovOEX
mRZycMmD67JztDXn7gTk/fZrTSQUwwDb1B01uLPCDbzT8OxUra0hXglJv7m0vprz
9ZD73VkTDKv411e1Ms538CdHy19dOjGxo7o81j7Vgj6voW1Lv9yWC+YEkxv6hJVc
oLDoZQcqsT9UjBj+tUwfwUsxPl7eHtnXvAoaNwT7wq1eln9DWc6kK5VYfp94sq+D
4Dn4B2hjhTgqOgxca48P5k1IQkErLjCpvt3sJyoGcG+cmWInRmWq0iROSVVq5c1e
OPGwe52Hl+fX9po0ydc2vL4ojFmgAZSSnqyI93xG6Uu7Nw/SOaYQVasqV8widhbQ
yAzxE3ykb3tjIA+HIFhHjqVdd4PvEt4bd4CxuvoLajSLiHCDZHsQdAAFG7oHFBFk
UxVajohdG41MJ2C/c4wS3L2CY2vhs7aG/m3YXKWgEl9flO8IskC1tsTPlUrLyzXo
RJcYunkSR8jVl+5aJan62G+cYZ8Wxe4ff+0GoTkSfxP9h67DJa8Mfu96MwvTUtJ+
U9DBB9Fmhvc+IH8OAe2CaMszp7kE3sumMTV5+ArrlwsqcEZDrbrOF0dBdNGTdyws
hem5gKf0Vj4Pq6k5DfjX9KaYpALsQVXadHEsSrM/U0VpwfE7edFq1Ecpe2IUm7g2
JMtuNULfL2VRBAexSTcWuo5geDFhwJKORVQy68PmzX3yIJZJgyz+llDplzFN/IKf
r7zISn8mkqXxINJbq2X+4P7PRTaJ7uTEmif1OWLJJU84nXSEqGNzgGo0WS0Ewhus
fBPwTFpMzRXCPivnBAhIw1ab1gtemSpzhsMI2s9fbluOVSJLpUY7jvC4JFZTUJTI
mNxQ5fIOXQjg2umt+d64S0yBA6NRnNq2Kdmh2iM2uEmAxVrVUqUx0EdJD5ADJs1u
FyNeY49d+w8M9Ohej9KPpFs1lXMcpYPaClL6Ls56zAYW0uwM7iXMzTe+mO7Dr6fA
fpUTGbisA6QT2RqQ7wayIMeJEK0fdOzAHlAOtlbpCtGR/at5vFVUf747M/mYj0SF
WnuM89INJfE4KrPdnehqAYf0lE2W6ahwUCId72ctQnkxMl8GYSAl1M0ctqrV7NoK
qol3bTzDwUwYS+u4B4Jd/oGMFRfnOZIBcQoOV41fH3o+K0r5h5pRCtDKl8buiyH2
spGkktMOIBTjj1wuhRRR6i+QL5jTUpqNXKvRQdjT+UNd4rfNV0uHkDHuWq5XPfe0
aXlx085ExpVohdrwiMDyD3VwAQrTl2j5hxcW0NTxsAPFwLqBsHeWhA3v03n8olmH
yQ/QsBoHYzurNJdhsE359iG7AKskMpxJw/uzF6xIYDc4ITyt+7c6NdSYy3oVvatf
VmH1kgtHgVuDmYlAVacCA6xMbRMp+Z8luPwq5pDDAH1yJenk/3fc01zfB4MoaOE8
amaOUUcPkIyhyYpkoyRXZkJ3CnhOdW7Lq4CRQnRZDNO4+VYh1NjtCucjUucvYIzz
yAF2JLEcSKFeNU0zqZzthKJ9YEvKdeP8JhbXBG+X26gVc2e8CK7p4bfYcmeVU3pK
Q6oISj1yDJsh6b8kHSwnowSc1PMCUXU5eIm5aaLSpgcw+xD8U3M7omefO3T1Bukm
3jNfpU8hHdaNdb+Ko1F8sjIj821jCJrV6TVUjPSrJibqbZ3wurTRGNnOTxmakV2O
26pXpj/ihCuuUGPasKgEEWNi8NYzrgab2MG/n+203MjQwCpiTjeKNP7YWGmrx9mB
78QaZbT1743v8mTXYZdRdPMpCn6ACmTYzqPec1oDzgvArDXt3SFo8YjfdFEqBKr0
FKCOO99DcxNx+eBDzUv83bILvPHxzjxD35dJe/nYFClMKAy2AXGl/ovw+fCMr5Xj
VD2wX7y9lYSUfIFO7Cx5rTV3/FYom9b+KssyJrekLi4yufrWhePe8W1DJxhRzb1m
fjz8CY1ikYkzvoRctqWj0rl/nz6Dxw50+RL51BrbgQUKUxm676sH9d4BNn8pR6nu
8T8V5vHbnjAwgwDxcQ/osvEtrzxol/RFiLOZyhgvtqaDHXN2ZP1waH4nMHBfBWre
QMY0eC0WKq+4gJryYsC+lIu/UjSiyb7sO4C7ElLx+PVwAdxwUduyj4hpW/N1el0S
BCCbM+pV2UKlMHefDzO2182czyaaO+FNTezaDhfAkb3XHdf6mLyvIONqXquK8To6
oEhAuF4QqiP32pxpXsA7g4Uxnj5vzm1DvzZGkOEaPSPSbFyXaHJM41TkOPqvl/pM
yfQeQE50OcUI0Lg93q+3h2t+T2R+jzn/YBD4sURmxOyDkbHTGdTF4BBKmXebuA4u
KMKwNIhLV6qZvGKOIW6e8NaXdmO3Xp2vt3gQtFZ5I3ZliUP4L6eVHmt3cftb05lV
fc+7X0xI8lRmJo2aGQtfZ0Wz5bVsgLtRrYrByturAArBPaMzmJJoPytt6XFoXIFs
G4pqHemiIjZkXMT/GGf/WzgySGZ/iZbCwoXPLnRUR/lgO3v/jV0bdWE+3JWxZPAg
4GTrLg/shCrOLuv4wUat6i3XeGkBvlkdR704XP+s6KuWnunXmsSsIskylz1YJ4lw
cZdYKDXs2/8o02CO1XR0sLqMmsMYd/PaY3qj8VqY4hIlgnFu4hAgXjowWSyKFPnB
4FLfCOU6WdYhkgW1K4jfg38PZgBiRWouPS8EsX1MsgSVEwiR+WADq5HPlqUu3lOu
J1HVPfaGMWEJl2naUWQ1I2WTpvMv6N5DMRvKUeAHzPIoUSxG6cPNV9F0FFmVX/lL
4E0HUEpxIkNDSew/ChDYw/dLnebh71zBQFrLjQa0AJQBFERz4loc37nsN/Ven6Wn
NZZbGIfNMUP9UcNh4cI4Xi8fBYCAKhCEPzw69VkhEOMhAYXkhfrYmsnwJNLhLCUL
hE6nYh37eKh++1CpRPVvQRY51osCqZUs7iDBrWQ4PLwAUrRBetehDNz4dFR1HBVO
lHJqJ36B/HVnog6m6sJqqTGK2SzEyjRWHsh4EGCMN4hTqFWLqw/nwsL4FfP1be/D
mu5A82YEyebtmO5rI1KmhzyIklNGw90ivhogNj/oqpYxVj6u/GT9+5EEpGlB4MCX
8Lye8g8BKySBIDJl838htjtNFnsCiBctB4AZT6sN5mqxLY9EQS7dTzSGLbhhrbwf
eOPXqiwsehO5anQmNiMwVipRvEpgd48HgKdr0FuVLE5q+7h/9sGjQKgzQfUuGhGN
F484OhJetsOQT9a33IW+l+nqqjm2EXPiCM3pFni8JAJm8PXPeA3iG5Z0W3ukE9Gl
9eH4PTB35JTek2Jb1jY7Nufap7pM30AHWMX3lOtOntFEZupQ4nosAXbqL+jXD8vD
PnnOJpN9Imr4zNlWMwzfwoXxhq/KK4iDkfDWsBsWAUB/Cm6nfuHIdACYEXTbWLFy
yod0NNEhaxlbb26ud1dw+rTGKEMqBZtkc8vWZX1u5nAt1879eVlJVpJMXHyIFWex
ZvVWrBhpxVRO4x/+dhhw9yJC5sVU274Aeg1NIdtk/yuP0TN4OF76ukziKrnO2wuz
cnNAhm9wpG//9y32xdQnKfWjKUzYba4orlt+YczQsIifsa1kJYN9HW8irq3KYXvt
s/eCB6GsB+hEE9OnnD00lwKwyg+YrN81/YX60UHhtYLwojKWwXr0ZoB46t+uk9/z
2ONV84Kh6zDsZIa441YnX3Tpl1siJylnKwChL20tXH0xRFK5oGjTcqzmLPYdpDQl
xcPmMm2u8BXuA8B2UGacpiokSKeXWkmSMr8UZ61vKw/5rRZStIE4dvkh62eUxIAe
ZM+rmvWd0LCzi/0gfrKSZcKxTr8GDTewTXE1hWPfY+WE3yuw6eppujoj46G9rwMp
v2KmW/JpzqONg/3/WN2J/9dsIBYCX9tP3uKL1m7llvWcGy+N7YWVKCm5Vyixfa7O
PtXYEkO2guuJZaSUHqRZd7843i9XviC5x1jLcudbt655aV9fo2CJAbSiwVUKnZ4k
wXEBpYhyO+oXwaTx6GVOCbrOUv4GCZr69WrR8kYNRLz0z57cZ3KP8fSri25lO2fF
59DGedxs+Qnu5JM1VE2w3C2NtELTgRNfMOXEljq8Gv/6LCyzQMJ2BDqbf1fiQWNH
rvg71GShK9sIUnfK9fS4GDRiUKidwjPqIA5SYxkbKq+VsIBUmANyPf1Yz0fwqUmu
hXCpnvUT1dp0DByluTCFXOaAjEgi+S+rZ3MUVa2LoIFztyfuH4Iw61jZbfOuqhPL
6AwP2xP2EPNkyf6dO3ilgyUW7Rx+b9et4ohchVjmB509gkvAR2sD2XaQ+Ks1uaC0
rVVTLR4IYBBWmslq4T8/L59uGckAxPymCLLz3wxN12o6P0kCe+6GUvTELbo595ee
odyv4JPsxX4WNb6kEQdQ5KF6hfQSCZ2syEAHs+h0oNoZpHol9vatEwRpRvXNuYLM
wVIYvaX16dBMAsTg+NjjubO12lPRJ+Cwq02qI5fj7e4O8ElzRbiCp+AblvD/DStn
YZ6M7GCkP2JEyUUipseVAMVgRQCuBu045+4zvQi6seQ6L9q5CGR+S5+Hsw/xa+qZ
MUpftIEpmE5OJvzz2q529wOpZ9n1vXVOoSy33IKQAh2Y+FFHL1EXDyCU/wE7AFmK
8MaZ8Y0ozk4WEY88QA07h/xunzI8DyafhRwpyNDkh4VP31igPYSvLtUn7J4DmDwc
GJwgy5XHEExDYte/ApMiUknRGmdlKNAxURwomv8wtPqu9ZjyWH7StQ3tn9BBNK97
RUPti3qV49OL8jVMeEcZG2kuwCqz3mPeY6/NmbYGF2vS3mxVDqJTT8+CQghL9Y6g
HHwEEsi70JE7POhCi0FW5levxM9AbSyfT7pte19rQnLfQfrtvdYQA51R6KmAfXYy
EuROsVj5UxBiT+f+qIDo3PYAScU2ZE9lLHg1y1yfmP0DT2XWYjTse7H53KMngAle
Z+NOfirlXy+4+AjWJW6wZEpDcO4IHYE9yxUKeBBDMS1Mp/YdpU1eW/e1ufnggfh0
FsigO/osiFbCJRZqR5buQxdZeTK/Pw1Jmbkpk5WU2qwyKmnRQjQzkppQUBRJugug
AkSmmvot/7ElCZAmEZ3JWs3PvxCsCh3TusEacMHmyEXDUJ21I0/muEgDdKeSKKqB
cHgaQsD/A29zhEGPT3zNBKpUEAxW+hyBMfGLywQXX9OC+JgyGLxJ+uEoyDKSLeCf
kwE/QRYvYktNb9V7/pE54IuVM4DlOEfJmGfYKda7H7WRiln3B797KxHM0YFp/KtS
WaDFwUWbypTX00c9VDwReNaS002EnzfkJpLk8L1yhqh9ivAxBTYMWCKGvQdCEyKn
y5hCC+APmv/acgWsM7FH6OKxyw8rvTNvFvTNx8eZG7KmqQxiWqJQK8sTISouDNVW
xQ7mll32bZODiFeTpHZqgrk9c1BZ/PuZDgDwRnhOM7KswiicdKKThYdzda6x9qXf
RhsD+PY/2BkzrJBprREFwgtoPXweYbj+80LQNTPZwzcEURlRHqyFxA8d2Cp9nvui
2VkAfl7hAilPl+3UPDWaEgkQZEfKst/0U/1D78wK+/LsPYVzGSwgMjHjdif8l0SC
m4SPpQM+r/Q7mmMlhb/oh5DRjqylG4GOci7PKto+658FxgRW/h4SUWvPeTWrOLWm
DM5f73VYcYZGcmRBcImfovCLrB51dZ3tco3R0+8cGAmmaoW2KL7WDauj4OABnmfG
dREaoaGBriaZ/SDwh/o+vE1EtouNYWzHC1kgQ4WbyEotab2EZ6r7TeiSxczeVyZc
yg745CC/5Q3jeicLtLBcfFAro5YFAkib225CC82SSNl6NWVtx49XzoOeETLzVdI4
N9vP8pwiTND4lA+2tn2wUSYV10/VwdDi3CRREn+eIhw26cGbGpMqR4GCgMzEfUYB
fraoFdI372OsBiuVtIewj6ru9Vq1/mLyWghxFw02F+drjpsRLODkfFFS7TXHJnUJ
Y92hmgpWiZRIFkcjD8wtZnWpSOnJ/TJM+8uf5wuulWISb/JpjWQr/MAVeLZ5trQl
k9o20OmxfzhGrGRf6xspmEp0ZWxinkMEjr0dD9UxD8Vmc1mTXgjGVlxEJw0W/Bjs
fssx+StfCCbnVQ5Vt2hqxNMSNpZ5J+1m0LnmiXcLFXqmf8nCTnCGXAuFuMhZFQNZ
ekfkAWEHGcblIxzIjqhG60jES5ZG9evpVWmikE/fsiP427DX2IFJ/1gFRqR0F/vd
MoPD1RAEMAhFkjdozKCuWIGUDhDc9CPpCw6SURXQs2WXhKFGcSNLCbgBOCyh5GrG
rO+/ZoUb/PssNvH/CS00ojXPZfbhBA8jHPHpzFMMdnC9BuZH6DN/T4Z4s+R88u33
FlxXK6VJjTlvlJqWrsyGi3LrL41qCUNbvxwTgtGLKQ4S/p3y4ZaIHOI870FX3sZK
5GJYtBXlydWtU50Wn69jwn7xlasoS9JYLKAV4PfOfnpsPxNfbRCiClcWiRES4GFJ
KvjCbza4NPr7CqM5+g0zTLIznKXSlyvsByCzKKP72NfcdsS/st8K8LG+6bR0NLzl
VdV9PjzS6RDm6Zr4lv+EH+xT/SDxBkd9jpoRYyEXp7hPnME181m/TOh+HG1U/XG4
pJ3Xq2kp6vjk/5pNSOUvTsdS1/oEr0cvwSlCr7xy8MUJAhxsDvjUB0X7q+F9KFJo
blstaJ86QASiU6EoQy8C3C9pLzQ4KR6omNrAkb/QQzLVEynasrcHSgbgDIVGPmuh
PXdYQTlfqrxVODq9puoshZhbNuo2cAaIDSh+I87UJw4nugodvEprEhKcKW8KMU4+
CDs5lXLTRalQGfvmfB6VInF8S48Es9+Dz5NLihRdIOzNO1ep5Byhf8Y0J7OOGpvR
OqqbzJ73LIkXuMpkk/qOJtaXzeEe6xYr6s43pRkuIvPdZVy6hXOZz0iD4EUUD0fU
8ZdEvo6eWTt5zs9XDa9XauuGTpnrX8XzNjDbfICyPWoFSi6Me66Wab/MXD1YUCpL
jzEJciEQHSuZS7lacETl8hxOi0dKR4x17nsn5hfYQJO55Kpr0CDvEmM7bOgvy70K
lHJAZADeDbD6oTDPQEwixNWL5Gtvd4bbYvFN9Jk6TRpHbWkgA3Y5MrT/qUNpvQbi
fjYdrmwk8Z/NZHvsP4Ko+YDqH+sktqNfbr+YSJ9YPCxqXwyZl3MzY39gg2TIOECs
qwQmXTPl1UvG5fw4sJFrugN9SmvBVRmjrXsmST22H/gitFcZGFbEOsfLIHJ2ytBt
r/iz6DHxAcGtF93epxXdLjIUf8ahkJRyx5EOpgcY7VrxEnYu+ZSxzRTrc/riCLH7
BmonHrt0d8b8fYY4SBNoW0fXSalITDKBGKUCZPJvkMuV/po0FoSuIUygEXTdwONw
2vZA3ZS4R3BCLPsD25UQtsMoZIPQ0tU3hZETqFZlpz/d58YTZCNjLTnJUSOemQMA
dyBbiU0P3SpWYhoRwM10ya8BSK3ymrv/Af1K0WlqzxyIhiOCg1I3amgwjRTX7ac6
pZszYD4jQqikR1uQRbn2YduvH/8noZnn/XKdM9NzFM+iwiJl0YVvnlJCFc/sSs92
VOjkRmgfeR2TPvCwovqRQz++9CsMYFVhL7xlKD0D91ew3iU+VeXmjTZ7fyy0Qyam
DSjLbjCh8X/LeEu/H897ONweeAlMNnGu71E6zLeYQNRQE1n3c2f8YzJJI+CMfY6V
O75S1nUhz3/4Md12Q0pG34k8hguASKjqjYKguAPI4um8QkMkTBYv4XHWSt5Bj9Ob
aEDNac5Fk0QCgcVdVourn7C0+PF3N7WaGfHPkpHKmMEKSSPQmJUYTO3a4Z6IBb+x
vGgRAoqsvwm8dE3DS+rF+728mAtZsc+OhpKS+7moLY6htQk3EwN3MxfM7/e0CWhv
3awBVEvSTPcEDxqWDNeGem+0Kyv+oNnTrwummqZJQdiRDRER1oUx6qOMR12Wukkz
KoyVPFa4lKOQx1qfigxniq3mgq8akIBX8U5b+k23Hc2W16SwznWQ5NhIeYNhchQ3
SaIPSREAIq2g92UMPwKwJO5kcYMvTxj/9lEc1YgHfj/3W5jUUg3J++jFwKFrFqt5
0U658IxRSSSQUEywJP+jSsxz/E8hvXteIaMPpWzeLTrJroYpU0c0jT9OtFkyMRf4
gWJ7zHTD0pnFzSjw+Tjnw0kZBnT4DEFyq+EnkWcfln8ov9wDol2F9fdNdluqfGih
uhVMC0cJTDm4aghySkz64zMH8vifMdZ7T/y8fePQFT7PnoXltuNqav/fYaNlrRDm
zz+hEX2LgZ71sBxgmYSecN8ZL1qVseF6Jb2d1UkKMYiXHxSGGGUXJ0KWHCwBwXnn
CqkmhzLEHVOvFhSnAmhIOYKnBnh2JhyENcd4g7MvlSaZQ/J2qi7RKEm/V7T/DVxd
YD9f3GIqkc59zSMzXX+kr8MHaixHoF0f5rltuZWoser8+s6hvObOSiaJyUUKs7ra
ouxFsPlFYTQsfa2p9ytf5xpoI6WOju8QvGqcZwiIljtPPBTmhrUkkJoG4pUZ90FK
JXb61eAZ/kc6/gkiQ1FeBe6ggciwkLhwHQIznmJV572b5R0KQaogXYlPfM6VhY4o
cAEc10K2iIo8Do70fkJBlet6AIhO7WzzzDmnmdtppsHNhFgboZCbwRMZh9ucUex6
YdALe0pbeu14mCNC3TVheCHv7CU1fjgNjtTorGjG4bKf6WcmbgPC4Ki9Ae9WD04d
WZb+N3uvrioSyABHs8egwFcenKstmhUChwvtd3wnfvpi/g0gdF05aQAZnCfYCgl3
8ky61tH3SfDTsXOpMJ/R9ITi+9MeNzliUxUTyrQ/R4yoY/BDjzWHHLC6TkXgrBgL
E7MXO4jNU3lawr+LtPZl0YgAJlwCbU42IXqGh2QZfptxc61exBd8M2X9y1ObJcD6
T3NU3jH6LUvH2tEx60FW8i3VJ98V4rlb1qZq72aSPzNL3zLZJbNn9UMxYpi4r9oC
/p/Z2zfkc+9BWyqwFBjtEdTbbs47+g0/m8zCUaKDbP2OOnMxiWrE2BCl7BK9xerZ
pi8Xn37XiG2mykx2nfL+F2Y+cqO38O8z97JoiQVFbaeLeQQ1dPnWJNnSgjLmfwDe
o6zvL+K8u4Vp/b/5givyoW+2IrRpZZ9/1F/XBoKn9M+nwVM7V7Hs/tebH6Crllua
zhHHbwwXiSkFvepApFd9nUCwes7UKDwPySnhihd4nx/wo4WtUQo85Qs6KhBYgy6X
NbmL+aZHvLcuMUxrqtczGNnG9v5ho4PoQY49fCAUjB7jnJfYbNk+IA8FOy7iFFON
vxv26PzUJeZF5dI6SbX/UR5/SUCJTrrxW/U2Z7VoxRKUAd4vazuDg3CBU/6J1K3Y
39DC2sAoTKy/syQ/gs8/IGYmTwd6+SO2auFvePmGiwnZTtAL6sqNLDhAguJM3tk7
a8jruXhTsDDMBnZ01ItbjEpQjMkegSewxbhLdNQdasq9rmszL5qy2HXrN1fVTQjP
tO6SV+xvZJZBrFw3KJ8AoSRcEznn0GT3928k5kNGXub5IPm8t56s2fiKp7SIK32Y
IiPzZhKBQSVgg423oJa/JNfIS20OxPkzad/3Jc95yEjjhCv/smiTdVMv9QfwUkIN
LBDgfEiHsowj/qAC3W9nVLTvwYGNZz45IR3jrx6Hd9+9b9JomXa62QTcMc2qGTvA
pk7aI3Dj9bCwUYKWlqSjCuuiewE0ZBgKivHGXyJ8xfhclmlIQRtgFno/9pJcjTWT
AJurqoFQw2Q223YOKvyg1K/zCp67v8pm8crpqZm/tZWx4XBsIBG+IaSRWrBeoO41
nERWozEmUPq1WfZaxTdgz0BkivElsAXgPp9efmvWVDvbiQN7YnWBSIZEGEhPwcyD
P1a63M9vbQHs1DCYmbGywrBnnoFFz//RHMdxjGGNEsSc2fpHsiBIhS9f+m+I3pe3
m2R3NS8O4kaSPMky2hJl2kjka8lWcrFV5xcdjm9Xt+0EhsS5jbfkln6/2pmTIu37
ZfhCmkDufvXXW+rL5NZAZoKe2D2qaeAOVIbIpVOPO3NdG1O/VJ16iPAMxv1Ec5vf
owvtlBA51K6hKOi2kA49LgDnnvUdlJzl1CDVOWq+yCCwtRsU4aMb2ORN+qlXanDN
hgPnw55j7ie9/Xc4vXu50hSPg7YMMUI8RGA+AaO4Tq2D4HSsHJPUOFO5AcIFHC6k
/nR73QQPhz95BxdKHbRGSbwiuBfiiEWPTKGBHLdrInATpbzvM9u8c3saJkmDjbSK
jtFylV5DRnvUkV5yzw70k4Ofu35Q3d/+5K1+GkcKo2ZDSRbclWZ3c6+WUOhiUpCL
jdEfhPPeW64XmllKA8b1ADpgkiXrj53+feai9q6AcjUrIwZhR+gjnwCKR3a9Np0z
Gvhc0ix+HGnBgO9jYNO1qZreYa+0YrR44jKr2cw/V5+0MmyUPDzax4oMVlTi0fys
HiSk/VAxpViQ+onihNbTH+CBmdMbcBEwL6iYDg4ZvIzCmmnnDdpG20jL7D7nRwDQ
8K5XjIFplbXIjSQzRvYxKI31i5oFlUNWvrVAo6Wf8AEv90qqUj0h/7vETIrnqupO
tv0blivGwXoTWbSPGJxjSyFEnsMiyTkPGGLmWP9gT7rs+msL29pFbGUGk/opl1hc
hGzpOZBJ1rGG8dd9EJCQd7o15Td0rXb+dVN5A29giDYr9vbPZFY52wVOf0Ph1/hE
eyS70znxvc1p/OnifSGiHBh3O40br/oKPgpZo1tIel45hue1kSfZ/Vs8JDSPYnqt
VAPpZLD/1wGVDO21/UEU5kMEIf3fFoUP1dA8exQQS9OnBTcLLb0fcLivJ6g7T6xe
UTKKoeBDCYoh2KwnMBZWgD3KkKhP4cngMOWY+S0Vrzvo4rQ7WKswEKuc0cbNrpxz
nSuNAo4sEr07jzSPwFuvpooU6iegBaRU2S2624HW9uptxTgUFEAbfsNru5SX3QwM
liokxfvnWPFBFlQEbrMYcrmlaeIqsFfb5FUs4fhcKZB67m5UIhqDdOQ340N6gsgy
t5MFI2vH78nMYGpNLSIa8w/e4k27W3Fd1+EHeTTR8+YDJoONYk35MMCYO4n5ZGPb
HsrIMv/yOVS11R2EV0beQFjLHDwz5OY3FeyHd8gbHZDZRHg/xcn08Md9+NuYr2kg
RpDpmHEpD97jj8M0QCk9n38cJCpxygKLvwI4xAQBXJnVsdP8XkrmLnEJQrHefujw
N7rVAXLLifottgcx8GerCUWqSu8pff4+YZ9QB/YwJbG+wb9VEqnuBcOT4PWrNcA8
YFX6WILV39QmTuQ6tn6O5HWUwawcoq9FnpvECLGaiMTPX+Ih/okOuTYYSpv8/3nw
reKvMTDfY6AciCNJCZOp5SFKNLd33bhz5JExxsc7sAxLx13pHYpWXSTy64Yr5nrc
I2noyuvun+AZrUmRgJpuToZmDToJFcYRrORs6zZoa/tDxXg7i87/bK4JjRM8337q
dA/EtsR89OBDGP9KQSMOuB1fvE2AGiBSP8/mR1smbZ0FOE9byueb4KDz2LLgeTBD
BFnCDiKBD7D8O9wVAIh/MNE0pR/t97M/zR/m+Hr5GC3JJIowSjRYV78VCvsrk+u7
HCfIN3NmNGB1FmWkrXgUIiMpxPpmDN53AEj7jdvslVsxyhxBO2SYYBInKQ+dVLwI
x8s95WsSbOXKfzbE7KowWf2mSFQJot1OpTsBZO3gx00LILJ6ml+aSEymfaQQHQNM
8X6fmz4Fq9ZFRwMcAr43jTXyRNRY4bGMBvUl8rQ66hyubpAUYhXR24emAHytxXVL
xgiXRw8n6FaxCnrnsNve2XNpWmfEpalGx9M0Qa5rcTAxEvio3wOXNkSALvBmYDXW
1q4K9qxpqgiXWLr3HryFdJ6ffk5Z+dcvJq2Mt2foMvvfNRqKkK7iLkH8QxmS4Fsl
ElwKVrBtgrA1AhgnXSDctmSPmx3+90Bsa8Urg6PVT3cG4yvCzZw4ZybfbvCf1ZAj
OcyBON6WXq5mTRmy96JRcsrOM9oPmjn4pkSzj9dqcRKrEQvX0bph7uKuGCPOuGk2
9vg8lZL2qDJUnobNhIy5KBy5NJEs0D72u8bTD4wFhGxraERSaxCW2MI8aCPUztgf
yzVlQIAiyIG6VrCgjTH/IQ14odGs9QBRdTIaHCs5xuwP+4k+AQb3kA1Bb+/ld8nM
l8WPwDn4SSRgbsvuY3jZZQ6ct4HL2Qp+3oEBSxLyabkGDqspN/R6D0EbGbI1mTLr
spI4rnI9HuGpKmjtrcWYM9GWb01WhOmaMEb7Hkwe/yrvqUABRKcVKHh6kWBFpKrz
haLKWGjwUaCTu2xcV9YG9wVkFkTgN+/RAZNC4PpfSWrkK626KoDMNbtxH9IZH8GG
APuyVGElPYQadNP0NHh4irlP13Vc8lSTeSqDqLj/vPESWJEo2xIjPF1eJ4316ynI
c3CrxH+LlTH1wEi5MY67/g598xJVNV15t8pgBiscpLX9wquBsNlOgkenOePT+KXf
Vo3OHub2g2hXSwawM6AD49JOUUtagA+ra+WiEaCZR4n//tPaYMX+P+7JH4t5ovWH
xhiCbGwJ8jtnPukF0Gis+OKqxuubFMRoTveajQKB244okx2ZaYzIakPS8xKudmgF
loR8IYg0DXZM780nRe1bBQQmg6CK7RAgpUD6CUIjnR25or5NhnFIPMvp0nsk+XAg
khiuPtXBNX606zHqkdwPkqn4s90qPy+KfQx0w5sbhICBMn/E6lbrtUYzmHZkVeFZ
s3YO29WVKuoP7tRV+OK6QR5NRy2TKGZR9/YgESdgzVvE2oSLTXPbhsgFe3Ze4tXt
r8qbpGlv9v17kJ65NKLfIHyNOou6SX0NJW89cAX0rJm7NsLawSh+Qunr4VHVPCXj
kkGUM6Kx+OKIaNU0RwjPJaCrjeIs3Lc9lAff7y/4pO0ol6MBsPGlsD4XSM20zIkR
HSsO8a+LBhplBLnECtU3wkl2EZNnlxRy1EHJqu+pX9bkuvDyaPJbnTj8N4MEA/p/
l435PTnqBd3Q3qB7bX+ZUBzhfwGyj9ZSbPI4K32qC2otfrDG7WL/ft9+UES8IFF1
odnXfavH9cL6qYEpcaWDM9nVCVyus+5tqsYU5KWoeAYHaeTFUWHDriaDGMTNfC2b
UgKjB/mVP2eEpf8zhCr+wjqoCAfS0hxyDJdFBjQ8CvSWG0Ml11UDVy0MxeUwj4FA
UZi4V6puaXHaCHa7dkrK8bFNJRxXxd5JRPsW/DJ26y7o+B3/hubmC7gH8CORLXkV
KvzokdL5c86MYEINIZYPG/lTlboz+reAuv5SRq3EdwaiJcntd78c64qukXATQYUO
Y/r69BrudLnJ+3QuMP8BxDGAPSXYm8o+3pp27ffS98aZCjtP2ARvdZ0m024P0Jha
FZHMlbjavZmZhcFJ3oGMlQVbPfGm85ElLWRFPnDqo93csFBO+wr61WQSmzobZmGi
im3J5U3K288iuv8cPd3+9vzmBdIMxIvpI2+KdvFP7p/jV30U63PB+iqSZSTNIBom
05oqUt/apwJ7FTKbUzNCtluinTxcPggbvsdW+SAFz3SUSasO9RTdeIMiNs4fOGzQ
i0quJD7Og2paZu5iTiGpZPnuUkaoNrHxDkBbE7p6kkKMDQ4s2tKuq3QhtSeA8PDd
QOLj9S4kItjgjtZelVePp2UjVw4JoRZ7NmtL4ljT5CKzHxkrf1pX1guIEwlr1Z9F
+hlDefEfdZr9iOcX8W4jkWD/sY3YZ7JdcwgYJP3M/iaF2iM/aoH6eJIjWfHRT3B8
Pmkq1g76AixM0i0cek15pS49ROi8EnRB4sghi/wJrIATyi9pB2YCF1KneYsJmHbr
H7q1WhcolsktAN47li81xHKvEw0SQnucm+oTAFiGxPMJ8kMZwyMNiMSJw90qxG8t
W2CVYNtEhvWvVXDNMd6eBpwLlYQzKLvsym3KsOYOTs8eeUBjYmB1Rue4t96PLgsM
Le8dosXkp7vn3JKfbTyNCN+iNaB7vMlIQczohaL10Sc/MIkr9GFWcK82xD+0r8e4
RDD7M2aAbYS5fa16eN02PFomKrNxQ6He6SjSCh7QdCwbkctyPBBcS9/nIuAE5bjR
zMkdYqtpmnd6J6G8Xf6hMhYT8tyyuRM3t3er/2m59wr8Als8YCzFAK7UozSBB8Ch
qC3xXIzAeoVMwyNt+kYi/C6iIlcqqUFQuvL6H/A3Y2FBC4RFXiId38OPUvi5F7bf
ewAw/TDfC23biRNQp7wLlg3rYiK6vt91nSoojj+MdO6ypsH8O1gTKl0RH80pAutp
B4yNzvUeQMN8TyOOYQOfi/wYU7CA/FpzZBAlcKff/Is7AHbFnrpkIPRFKGIxJ62v
26XSDtolen0mbyOyvB6AQK8ffWZ/aM5nzBRo/UHj5oiSaWJHRE3bNHc4bN6gRMEU
Tn4sWc4vDaITMv+/wq06Z2WVqlX79Pc/A99UYa8ppJglifiJhmvr6xD4YTRR4Sfr
kp44egTRUMfwuoNcI8vwLAbKvasPKWPodgu3+jDxc8mb8Kjvgdd1wUiSXAu06RuA
2hS22d2bYGsXKHibwAA1QH8RSclw51Pmf1kaVVRjDqSYHqI3YtxUDhReqNE4YkrS
vY0DC97qK0fioMCRta2KlrTomRsQoGID39Z7twabcyMEsT8r/SgxNAgrIsaZGOum
hL56eLDohso87z36AvgDLHlIrm0+xWfzvuQjRPHDEWTKb2yDJV+djSexWAIChW/o
LYmbLsT3iMoOjMtlaXPUYt9nbfIcKGm2ANyLhDPNDQ56pxVLUddVkRGeimiUhPv1
8Jp2ldIxlMp9NhfjHWRuQxl/2NSMXbc0yW57HT9pDWDDS4vBqOY6bCooBjvgxMHw
nw3OOh5SbzNJaMozze4odHCM62ORavJ4YeWHpeWB8dKcg5BGGgiu6z5bg1QayM4X
m4IhE68W5pFgNeKlOEfLNICd7l1/9q4LXo8cKZJ+voLFWblLmLCoP2+g2vHJ7c5O
uaHvDdcCCxZJBA/vyYKxSADpJqkBeYW5bhqeajBYuqovhdUlejGDuARLeV40DuVD
lMy4HOxNh+vwG4c+Ajalw4h7/v4ofdqqcpltLuwgSMV55NfVgfhHyvGIllK5yCse
T0fK0XyBxyg83HVcjaywWpqANSDdRcf4YTQkKwv2zGlIIJ4p7TzhJnLTXEAyaQzC
yY3L7YRWmwjD+q+z6/9kYdxvmgMnyAui3zIIyUaGnIxU8crpgBShqWum97IHFKzf
Lr0WXJBci9yck6eTJHacR43WfgcDa6O9s0zKVdGTjUtv09KDBRKWOqH2Mtzt963U
8QnE1iyA8yeybZkPePSkC6bkeUzNryw/3UhopdUQ/G5QM3LKp3fUHICjZHEc3Tk7
Osx4gOdOKNzeqiZKUBnxgVGGLytzrF4JrgZqTofDIMI9Sh2BbnzLvzMQeUIwwrHv
xAlY1a3NTugWnOgtFxZcxzsdYgefKuYXjnMPvFBqCE5xQUVt1CeYjKIbMi6tggbk
trY11RWAqb/CXy5Q3dxGAAkW+9p5weYY7itaC8j6JAbaNy5COPyysxcdtMRxe9in
/gsRGUTGeoVQsbbOrdM2eEGy2liZfKKVLUk/bJlSywi0NKwq2F+8kQYfposBmq8I
FKkYbPcXmnnfGsn/ytFFFd5JsW1+eh8rrEf0ve4N966cyRwyhMpKiSwHNb9IxgwJ
hid/KyGhdS5hyoszr6lT5zr8cz3ccGPPxGFZaMVBzCdVAVC80Kwi8mtUe38g+iiw
mbfsxSXaL0UxkEIdP2sqSjPPL5de9ef/cUEIrMfd1ib3qNH8f7U12S0ZgM+GAka/
c2BTf/fUtBTTZXjDAToatV46DqIcBhYd8qze0psL24gLSKm+2XV893Xd77e7Z+ce
mgMb2ubGwhIOAXU9tWKEdLcYPBjzI1bCPBxgy5XQLv3TZlI+qRUsIolfEhEeRTiv
MTh9RzCBPj+Az87gf3HQX0P+qsNSRTJhLHywClQ7UZBOFUI/6zUX6d57UbiDUydg
xe2vb1p+t1XpLOANB4A0c1h0GlzDV8IT2WgzD1BEDegi1SFIrgaqDI6VZtDpDdGA
KCFPfQ3pveQwVvf67I6dd56hoJvoZk6zha0ioR6idiJzyqEkUviEmJEswp3OYAKx
m0XilAPsULtZLIU3jmw7yFHLZsM0hC7xMXz56SOrwudBBTuMy9ylvbFUerOCrBRk
wPYNkkxiSE54cUYmL/hi4FS5Sz8EKkFBBkBvU+jNeT/o7sVGYEqthMAQlwOHr3Oo
9/eAskHhYE/llC+6d9dcJT5MPuqvdlOq56PhTiCitJ3I6Guf4K9Ei/4MTafWi3Qq
dMEKzb0C50vNsmI24KGP8VAw2G8+yQqunGy2OZksDFxaX12uklqblPK9oK8NIjvI
3hriNDkdZd9Clo0DCgW8fywSmP/0LoEPnWnBN2HFbYbzrsp62Wa/VnpKxojvswh+
j/LM2+fqheCcAIRDoO6IyXMSpYemdKFBFztONFlNTIA0nml7lNFuKOUKnU5y9OTT
9qrS1FtYZw0pNT/5RZqdpeVDcm/2MPPkg3qNchWJRNg3YH9ucBFAGd3j2byDh39c
n10sNHwKEAlcj5eeNtTT9pRQL7msQz9fgPFS5boGglXxIE5Xs7f8rf4eXOHnQXeZ
R+t9P70srr4VdvK47TGBkWLwUZAsU/jOxb28OeA2qWgMIarOmbvKjqPmtclj0eV5
uiPAZ7h+M5VBz/yXE5asIHjdlFNDE6MigIMjgPYvPQHA/E3aAuGrbTDoyXF83feR
ozL90sH7wjABHDeQy+W4+VQ3eG1ahtd6r9ru9nqoTv/jOgwjxNKQF2NVWk3+ALFo
qt6TDRbiiMSLQityqzmjYDwd2mK7hrJ8T90P2vSgHhUDpfpvqaWmq7ehGtSjcxN/
+O6ub/4yePR61unE4K+47f+zRwXOhTs9urJc5EDK/peVTVHYY10wDJXRRjd0PrDz
fjWOfMJUsDP2+LLypADXzwDQ4HguDAQGvNVwVyXeZfX9BpKE7ssojJtNhjkNXBR3
T/A3HCZ5RP31npQ1aKmcjw99BhPot0KG6+7MclES8exBSdzQmkbPAARyWE/ZdLp3
BtcKa9yXExXi2g/tMfZuMlxdJX1ZStBbMnovzf/mXKQRXajUuufJsK5FI4d1F1SU
E1XYg2MolpgXaOEaJtKl23ekR1GnkzrYj5czOcg+mepw8rwbzPFPvaLkhAnVZTIL
oq4QT9KBIO7OlOybjm4ePhX3Pddt7xLsJga6iQCc4UzzXio8ucp3zR+srY5m9Wi7
nQVu6uycMvQ4kJGTw6Cu91MNQlM6GllcdJB3g03LIEO7hQMfOe0VdkDDoBNRcgHf
7BDvV5Jnw4DAWYnmfhbU1y3rIxuRFIZ9r53A/n4B8Ij5UX+YQ14NctP/3lQmpQi0
OfwXkxRH6ztgeU0njCg/9R6S7jzqx733bxGlPB8cMKG9x1kxSe8xhMfi0m/C42vz
lzs0B0rP0U/LY6nnSpXYkZrCMPaAgbI1Ur41R6WAux5pGUyn112Z8+fHc80rLGTr
5YxQKaLWGAaLVG259IS2QcSxEt5w6cJESOSQTgKbHeeJ9jojGtMTA4fjMPALNzp5
k0wPmEELBjnmr7YibXBWtYBFPCC4BaZ5//9jEIf7yS0ov61at6N3nmAaDogHmdud
wPW7Bd0C5gyLtFDHIGz9imNTv3NqYX893+5tLP5cVNYuhJ2giud8YmsPNQwfza4t
s52vNd+DybDk4Y8N3U3wxpb6ynyarSYp7JXVMpvYKFZKjWEGTdt4Ua6aMqhpL0oI
T/k+J5thtyq2Y5WinUWcxgGL/gx9r7bEjnfCV4/kot1Cc7A11znRvOdxteJpsR0M
p81JMgMCOAwAHq42oLUzhgN8otSmB1wt3f/KLaxURX3RV6f4lyEkcXS9+N6Qt3FD
iKKQfJ69v9gMWvEHAwZOje2Lg9skK4kLiRTY9ZkFu2mrU0GwjDirHL8L+tCJyZfK
MSQCU+iPRkzFqAKfhuH1LvB7i6mErGjdZvuXDmSRypWNBkkwnSbj0cngs6dCJ+jI
p5bPS5Uxsw9fuyynXTKVdKP6Xt4xKnCCNLUGDbobDkdfHskgt/Oz7YpEZWprk699
yWQIgdS2RGz+IvBTj8EGg4oEAgUNMMnE+N63UhKO//dHldbtadEeC+cw20/x+BHR
WRljuTdYZ6OdxScD1fW5iVlByH236/yIKgdkVS9DIEKRwQz9GUO+a2E52FklPG2N
ZOtcgHoNJ3JWB6OaghpXMOfF1ceCphm8U7+5OMiN/yOpP23vNNPVTH/fuWvF+vte
NSCscx5CyiOJ4peAYaJu6gOkCXjNWjPtdo/f8964HvwXfZKNogyMbJO0KLki//D3
rDv755ChDaMv2XKNT6LL9negW7JnmwHOgQ9MomZrdyz1wDx0a6iX8P+g5KVoFOnr
l6KI9dNQ2rvP81EKnvey2df/jj5kwjnGdTVcOwolyxSjoNsz8th6MTrdSw81TDaY
YZFPp6Iv9RZg7xs9KDKmFVIWVp11uVoukKdpcA+OQawGJeSxgz6fCuSH1sTzaF3o
XoaUIpV2RCE+yTGoQXsRVUFi2GxbsbdFqnlzontgOs+ZoDoDujxoSxpXFQsvYTRm
q15OgwyroQ3EIn2gK+rVFDu8sgM0LwphcOxnjFKlxX4nKZKQE6MquTRZ41125T3x
70qU2p5H57U+fmX8i1zd+FjUXyE8r2piQP99FzRulHVhjG0xx5fU8HcjhQxlRwsJ
0GS9xZ6m4hn5z1BiFcDLOizMeM2QlJXfMtk3iiJ1Sth2TxiQIJ4rSrtEgkJq4qQ4
EyjsEVFdltUSssG8OIAX+5QTbBIdTCJ4sUeRpg9zZqrrEJxw6qSLobve3HBh7/ds
CMFQEbg9En1PND6NuKmSQW1y2Mmq8wTA5gIQD1rCScEIHX2JKPP7XV+z+gfaiYbD
JNwhYFQu4spAVuSCvzT1vZr7lB6/Kua1r4lorf0F34yA2pVGHA84iKHXjfcGdfE4
5GnnoAPfKmR7keVmmQJ33Tq1/PNBDe/XVcIh2UGfE3ArjBj80vQwRTX4ryOGkEbr
7CC6z3/DwcQEMmcrRe/HWB5eJWLPfcOjbJgB3jOBhvmE8P/cjtndJMDO5vnRUq5K
TQhe2TvjRlAUwU9411OyRPoZPnUzfI3mR9MXKyyiqLbe+gYRc0IV3IOLW2IpcdWA
SMUnOxvE6cxJuxHc2nRU0Ods9oND5kadRZW5qzgZVJoNDrYWkFBzwWCSw2LuNfzz
sJvECvUEe3BvT95NHgu2yfQ11zB4TnBH59S4I8QOR1drqOlY2vof9Ei4EZ/guoUH
p93iPV6ahyuEzV0tksuW5KzJdUEHF4S9e2+X7ppiiu7Ke+shTuWGSCbFLzFWEzHb
axfXXwAqQl82f7LP8KnchyAzu//igu3PRk/wR8A/m2Xp4v+xNm7LWXpMlBnFQC5g
VDtc7+uTWegwQR+4CAAs0PAhSJlSrzi9Wc3jTdb4qBOZ/sN0+wgF2AeiFqDHqvCT
wuDeqGRhiOmW7InS8w1I7o59hfizKNBEJc9Y8HL5BYURusWi6loQZfHtC3H6iQm7
+M030xRekPOOA4vjaO4U6NteYFTJw+rQevTVHSCfAYeUV4Qsq6PlbzImzYKdn0IE
ZvNHGWkUra5JavFdGem3JxRe+f+6HY30USJoJz1zfjGB26bkThfBbFDMeQbFEaTv
/7oUAkNfeacrQeG0617eWZ80c+l6tP8DvmBUEC5GmPoCmH0H5wKVGckaAbP0nL67
qi2BRdgD+/WbKh1Z6b5BmkSVmf2coiJtvHo0XsfIpUIIKlKpGOkMu5pGeGC7tf7M
KAm7XobC7dpIv5QkWEnE5TZN6190o+0iDGr4vMsTEGKlltF607WRo1gA79QISoxV
vR+HEHmZj+sCNrOTNRqOV1nZZbZVRPsq77LVviZFHIYC84puppZnUMIjkJTGJ60t
pEldgIv2CoHBhbS2lG/ZeA2HOP/GIPOL4x3AQqvCeCjsCphW9l1KUdJywd9pbnDU
j/jkWCDSrHWdjrdp4Fc7PB/y/HKd0SfeB1frr9RGtxY8SqcBAAeZ+J9PDGwlVTMI
FdMADjLJirX309PIAfrmXYbd/v+0RfcCjjs3RgBKpgrsr5ObBxzi+yElB1V3/lsF
ZcRkK2Fx0/fIF4PU5KNGEouSqR1vu7XyaApkGHGs60vDBNJIo78xmVES9Kf/G5Xl
MD0jJX2X5NvvzWiygTv+FKYrLaLtTSkCKKc9DpwaAZji7ldF5eNqnG5ZnpcSKezw
wfG1mycmsP7AbUK8fItdZlIIOlDFFxWzJ6ziIJJ6EquR7wAyCR6cqTe5bkcPBcpN
pLqqK2H+G3I/PZzeLtr4YUskZ9xW3wkPW1LL4QZMdNwpj5hIvesOy6wt2yxxq6W5
C7+6y2+CoFxC1Uu8ArVubDydTh33z6/GhRr5HC6eRu0pnhJS7pmgn/IcwEVQRkNR
qDoSjpFP+/zpNYyS3RKE2RvbzrtPNTS89ps5zQ5HS31pMJy/++9/EmdLaV1ulByd
W/YGVGVe2bjEhYP2gwrBiSVNPLA/mkThYPGzJTwBpE6K/IbI+k89ROIUpgJh3R9O
X2L+LRDEqyXaruqUtcUmOfXFTMwz6Bhe4sLVe8j5sYv8bPdlmQe0Pmn+3ILljZIG
fb2h6ivWIhu38345Hdye9XXSLpUi5+QldyaAQ5Pjin/3VEvlIVQQRtyKZ+o+EZCB
gv69JGn8sNlra0+MaTrH6p72fra7iIdQCGcbIGR5kcKY9D/jBV5xYWb+a5/edRB1
U2TUcENRP+NBGdCIGqtn4iJBouJi9295WzPSqoEi+gNX21wgVwoWRXf0nKdp67Hm
/4bxo3oAmIoPUDGqJbzBhWxACBJ8I21mOaI3r7Bqb8fmsHwjC2C/6u3MggGsa+XU
1bz6EgfhZjdGgbp8zi5gUPE+jLVN96eFAAsVyAdnAL1Dxuvmn3l6lmrHbVhR+YO7
I8UERoZdBQxmhl0L2iYR1XWiBggBHiyDmU3GE77y5GV4IeSoyHvInTWHRoRqyReO
vhaIrvDW09S+or0+/V5RtkCqK+nGobz2eoYrLu/1896MMXggxblzk7tOK8QtPuqf
fjTzeqxoN4y0vCHOtK8ZCG6rrfIyLWAtT2dgouGf0nQbydcn6Quv/zpuezGNoQwM
0K+XMd7l13337wvg3IAeXz5p3RaAmVqEiq7PEJUJskcbTBxXkncm3AAlp42aBGBU
aczli4CY7Dovor8dXlOu9ATlw4yFKjEnQcyK+zQb8vYvN4+QcyPPG/IVsL2RAOYu
8Ugt7lKnphPbDIpjJiFR8cLO+EpIBCaF8gXBc6Leb/dpQLeqscQEJdRB8lv+EXfa
f4BHxZrhaLMakuoevSIvQ8Mzp+I62joPLib8WogK0rsDdGzEAL0iiYV4govA0uCs
t8uHKE2am7tEXg3XWxr80eyfowFJiL29mcGsnqqkLMByNGhdvkFO4QFwISE1RWo8
rFXV5jgU3KxI/u1ihYa82HHtCyE+v2/8oOJHmmEpnI/TI0Ot8X5IvyG6G5nJvelD
wTNGe3mO3H8m1+DDEeJw8k3u5Hx0w2Pqarsk7QfoPVXNFwBDJ33JKa2QIXUw8QP5
wvR0VF15reMDyXhWcqJP8urZ/TE9H84cIxtAIFgfj0LZ8ZHOw+y5pI7nVGcnSDBL
ubVNYo0+EZ35Of6OVyf+T1GBI9QYOhzfEhVnmTU911Yzj69EuinxlTb76tlzRfta
0S8Dzdd7Lq3xTlD7ElW1dXr176qMlOZlEu0KqkpRi/T3FI+eihRzIZTNH/7EjGHv
vSmhZkliKGvZlswIQhSAQMZBwWJRW3AR0EuvbG5RWmzJpbWXlWNGVq+PVa2Rr531
tBHjuP0hYtjbLawxQOQ3XP6VwI+BqxJH/aXZw4EieIewmWma9huId8LigpyqFoBQ
NHolhUOnYhL/hXdy3I7zm3pMb1EPe6U6Kx7OYl1v/6qDHOMKXdLGTBQ323yXDGMN
3nSvPOB3RfPs+g9EjpbFB9szMko6Rl2s5psGjYSFOUX/g2cXmAR+J6gTaxA4v6ho
kjmkzNrz4ERWmYYBkPj+72weL+pxwdRCOjKIzxwtbmbwIUmrpiPm3EZ1cuA2hskR
VYOpc+p0esAFgyGxIiWS3MZGDDxd8UwyiN+LDfigS0mpIGFiM2hz0ovgRjFBPKOB
RpKi5s+sqHaVr9XTdkIeKfVa7L6YsEr0PASDtSKuuF+cHCNRlEAixwZxrvoB1vyt
5hpJ2wOaNiJFutd/dsNkHCA/ZVguM7zaW7A4+aIb9qhrRnkhEo0epfRt6B52uYsn
YX/xqC7vGJtx52IcqO0TFHWp2GPKq6g6RZb29XAvUunfzImsSk/f9v9zgPHWBT6J
hROKdNdwe6UdldNFxJFFtCHi0tG7ThD8KURn+HRvtx2SRDpjO5eM0AoylPQqa5Tg
6M/EN1aVUibHjVM19+T0AN3sJooLkxm9MiSu4rhh+zQYgrWqhgf63IDQ19iZTHpq
0FNOKjbiaCSmHftfKbxHTHdJKxI8OYwYWAWULSzx18PtdW+vxeLGq3zU3GS6ds8G
UqbeOhNeJZLgyWqFEjyRkKOsPscuMiv0S9Mp0ZKjN/ZoA82d9BQBukYJ0QmwdBgN
d4eiShsG+pRBX32DgDJsRdHcA/yaCXP2CAoH8XjxTYIL1rxPXEvqPO/YGH6qS8L+
FMrfIMQ0634RxmnRjvV6auQHg9C8WxHH6hLkmaoHDFR/MdVk1MnCPoFcGPEvYGui
WkDjy5b0muckxXuQ8UP3J+F3gRknB41pTzxdWc7H9ZajJJCdizfXJFQIx36+usV9
MWolbVs6efXiuGjsfKp5RDcUGQURsPZTZFZFtYwlimNa8XSTl+Kq/molYrzWwkjM
zQaee512Sk9A7UbcjhqLTQgV2Te0x2GPU7x2j9jQwC/MczdqIpGFpBYFUQZz4cME
10D0J+/z6vHzcrH5txRE7yk9JQ7CI+vdUetxYkiS7so7c53Xn8Kx/NfmJmQSlKmI
Z9WKhxgMTzUz0bDBu54PRMXE4NGLS37yla4ego2CYWC5RQFPmao0TMwV9rqGU7xJ
MaxdM3Qib9f2+q3bHSrVujndZAs/o+ZlHn3/I7OhG6WDpReQB4H9Rv2KJZFi6YxY
9wDeamorZnP0Em3pLztwiA3b9m9ef/SAZ+anrf3et6zZP94FJg0yJ3+IQtAEs4vW
OVCvqYq9tJfEMeMnZPA+ZlkN9mneYMXajyLLu8yorNnqNaDUxu4Ih80slnS+Hty+
wIoP4hMMe8yAAy23f7QYu16Z1XiD9T1rI/3r0qqMIq4wfyzAZezUsvYqdqLhxgBu
8BTflj+kbFeUlLEKtcsnQURyo9RrDeTYhEIbikKL4lzCYl6nCbzbVpO22+0xPyRN
V3pqgbqZ1DwbaPqajz93MR0JpSCDaHauSP4qHoi99amkCd58Y54CkedtP6ApRazS
bOp1o7NJtXGFthMNslAnM9PifFKB9WKcbX2z122F9YDO0V7YEKCFhiErVzvoxJed
lPfAghQvmWtTNXTDnX7GZfX3pKBi8QEWrm8T5oMOg5f9tMysmhie4sy02N6LO99H
7nEeL4+mgwD5bKfGvgxoNW0CIXcc+gYyVjydgODfmxFNeT6UGE/RnBakhQLaYXyz
6a3j2ietCklvM8xxSJqCvAlGoAzQ9ml1em3i88safR+TxBe6fkUwLWNgd1d7NhV6
vHyxvNSFDfh7W2p33m38LDRfNxHSnLrZpoS5jSYS6tKAKrHHXA1+kH/U6/UbMOZL
JiLAeYSKXt08XQLyk2ybyn9C3ehAh1ImZBnsZpE6JnKONWAoJAdlvU2hHVzsnvQB
/I+fbIL+3OL6rWM/HbisO7Qe6sLS9GuQ57KzpJXLU9rorucBMusoIG3L+IYOWqKk
CO2VY+vj/1AIKYbUxYcbO8E5jgnDRi11g8OJmuj/szYXrjVQ8kCTiXGZTuJ9ytoj
XjfZywCoG0cY8ayMQWnWaRvbMVypDsFNanO1X3/gyj7BLZajOmc2K1KLpK5Ilu7z
OCzR3VAxfk2hBLY8SoCHCPTEx42vXBGj0HPYnw5qwPyFABKx2KQOlvcsALxmgIpG
iv4k9Eq6ecd8QLwglwx04yB0N+cFbk/+pQ9ITrUmJsn9hoBevEpluU6CF5EvAyGG
KI3ngOIsBkArZvQot6pYPU+E9nc0yYXEwh0JL25A6OQuWVHnU+7HgUpTDXGj+Kox
TgxcoRnLwKerN6v8TnEiWn1T1mVob/WM9RCs18wafhsMsCTW6TM6r9qPmIv7M9Fl
glqdLE9547d7iHMDxEfjhdEeKf2tF9KsLi8dvMbsc+fCgYL1mgpMdiY5SDPQpPo+
fK3F0pAjBNC65iwuxtmyixLhBvyRxcxuQmBE93CwgJqZNk/4UCklDVyHah4NqCvj
kAzxhzA6SMoEYXLKM2mwvSi7nxxYAOG70oCQnWtTlA8Xv1UzdGXaPZga2kVjnRxF
rrBbJFOURVtigOuVP4wEAVyx561QKnCjJk63EgBSW8/RHefo1k17bt8IRNpFhkcb
+405MLVuTZ4t2+vXihS+bWZowQUs7wqlUFRVqgegOUR0eEdzNwW7e6ZDFXCqtWAz
s5uTOSkDh2iD6qXpNUlCmk5j1b22mQrdW5E70cUmc8qoAl+O/tS4DsPN7eZdpZx7
lggqh1g87TTHJ0lX76M2HQsZF2/vwxNVMNQgfZdHuOI4I0forwFfzGsN0y6Q0aT7
/yH6VmH/TE1eJX4sbxffkcqse8XiA0n87bGHHDksIUA0/CY6ysy/NgHVHw0iS+6X
jjgIzSppxooxFuBABE/a1l5hHQV2W8MLcP3UWCT97S+zMzmInwitL3vC8EbfjDEU
DDxTg4AJC+Q7ZtqQEdWFYaX3UVrFfPD4t8hlxK8AoOcP8ESfcwPioL2SoaYfjGZU
EoJ6Q1dADK0+Gx9cuPjs3UcKlC0C+vjHDDgkuNO/6KKgbCfuwoZkf/yezsAVR7rM
Yag08ktmU3VWtSurxTWIWIi60V6OLSaRhff6VEvmdsO63aX5ddXWuVI5W+VE5lzq
f6IbviKRghEF+acleRBs+K+JRsEcFX5X7X7OtuyMyi27oQHFIpj9wsjS7hrt5PTY
tWxsdEfJNO04A3r6X2Jz4Pfz8X1rxpIhg27Ig1XWstAUMiweobby0ljzLBy5dCoq
LCKRknjSVRlmoO1pwcALMUcxb54TB+2pefZ56tCNYMaxQkKfSO4aw/jVFWJcToLH
ZWeK8e9ffja8aUJ8SOsPTWB/mkTTemY1QJVEgzOFBYPEnV9a6oH0JguPh0liNZL5
OHTw5rqufsxbAdI/NeSdz7NX4cVe3VskjOYWmJnO+2HF76/cEvb50XplNtS2tSMv
nS9buNZ2SeCvafgFFiiHZSjljfeXLxUnwW8Ej4QBtCUHCYj7fw/1IyOn02d7MATe
gtIphHxKmxQor3P/y1QAW3EAKw5h59OzjpdLjI82uCvt7bpNI0nP85zYpaIu69Ts
r59o5OHokayp8UbmlZWHDRncxiNwM0vjEHdsGGeUfDxpHZ0JH8J3XYdFOQgup4Yl
IEEkk/jD+7NUhAzzTtOg8XB1zZxDumoNf//9FIQepN3b8vQl462adwAcQtAe/GCK
PcsfJmuFbVmYq5Qhz6OVSB/UDTdM5SwzxsyumZE1UmhuSW2ejnPWiNYI3RkBKGbr
KaiDok95yzeScx8wYsZM0J7UGJvnDOFmLyxG/4VOe/z1LP0IOMsYvQggaMzNs56b
2egJNKpYOyoh5iDBMn3eHCSXTjFO/1gA+lkJkg+ZUqIOBOaCqqj40GsUwk+yIB33
0lU/l0OQkNqClTUWVjk4/coFfKQWHJ7uEMPe2IFAL+0ifx0vo3+aCpDbQSFpLPTg
LeQn1vTs9oTcleofJdyrolp9IOt/czOjUPyeW+OfKbPMY3powWdqX/O/b1y1Xp2q
26y37x2eA3aRRAlM68uDXPkMrp6BHx5h9b0r8KvDNT/ba07HzApOZc5Vd4/KfSig
MMDDnmGEyP2tH30AR1pTpILICnl3EYSF2XUpyc13U0Y24VLg6EUR8VPJimMVpIOw
trdUvtJVeW8HBX2mD5RLVKUzCCKoJLTl4igsA0AS+dMIiATwCYfnJS7JZJYEMxc0
/FjeTLHTc+A9vA2NUWaA2eAKGhAIzBTM4xbR2LTFDxue0plt1JnHvnMwc0O3+KFh
8XPgqxMkLlI11KNsHkqHqf5k1N/txcvoKDIEZ6WwMH/5w4r11x/1BcngUXLvuTS3
Bm00+L15PsrNT+YJVYCxCq6VRx8ZOfzMzZD/rewQR6kzuz2jP/Z1gw3T6rhxJdcb
Ns/owyxvyo9jKt7UOKj4L9/VuWFF3B8zPadnXdaLAMl5rLTwGeh2IBOaogIcc43z
JOlQyiEVDMk19dqny3155Adcm4WIViW/pLtOGBTVVPpaEtiTVH7kTbvyO1jnUsC7
d5p2FqTWNL3HgJ9tguiQ0OnDHeSo3hZyknaTSpcueO5oLCPSTmLTynfEh/q324JP
Gr3sNGrla2fTQTuJkKmZ1U7IFDMVmiSSubZAUjo0YscGXwFQxUR2BodYtJlWHVnR
p6B7WgVwDvT4CKpA2j+2BJWOcR/1pts2lTs9uaHE8r+WuHnkrWMu1QsC7dQdD09e
nm11JHvKvSsYCKHeaFwHxFXd4bDaMLAYsMqxSV1mcfgkrhj+XLYytIHBdJlrXtsi
OSppWpjBzv7n9Vwpl1LwXQhMIDirqanQvxmcg0o7YJtvaltByRH8BEWQBJXENlAB
iQLX+p/VVmhFK/A/aF3AJwQvhp6Kmc2rfNYD0Z17xQR+73ATKcNo6cTfAF6cBB83
kBNAwnGhvMtoDK+dD/UcozFhXHrKRs1QQWQbq5v+ukPEFd/i5qXPmm2oE+HV8XzN
mRTSb2UeZl2aOzylhXpSG5HZPDdHSKUJybdkNF6m9m+QW4qwXNFgzGVQqQfYplJQ
KhFMY20jA/oPNHEuahocMgP65IF9z5krt+if/S13aD5m7OawysXvPnIdEKOVBvju
1iSVZhRFXSlI3zK1xkU8EsUoFMh1z7bSOLH4PIRirrmsiNAfs0A4/KoU562tJEVO
h294YdzDaEyAQ79vSrjtt/vJksItDOmHml29dF40HeZ1m7+MWUVdbKTSyuTvF8J+
FHo+rS4qOzrbv9eBDwsV8MfrUM1hcYleRIaenXFfk6r4wzmPE8OjpVt0MmYpcO4K
Srac71bY75bMuBYbr7wqwdS55BwB5FRhkZSCSXY1NILCH98AGkN8hd13Wsyf/d4G
ieOk1fI93mmnB1FyhVPRcnFwBeYumNyv475IIMEQx0U9eKAwPSIFmp85Oa0u99Ei
XbWaaX6tfxK/SXEhbZZTpVImrQ7+e3v3qu1tee5pJyXrZsusZ6CEOpA7vSGmIWrW
148j5p/3EOtp3O3T+31bGr7cKC29Z6GfmKAfcOitZZVTHbep7ni+wL11k0ib3LRW
YRPjESUsTtTjwvc3fBgH/SengGDxUWT/9oPHgirKwpSS5B5HypGTCdDkGOz1XziU
40W6umLOkxWGrP+kilncOI/C6/jR4GdmFulhnyrXr5evCmjXQV0fhG2Nj2Qk1qMY
07oXwSe8G7nIQeO5lRLJ6hW3/EiaHGnf/LwcBdYrtF10jLm9NXkr5gffzqYy1Pyl
bTmemfgsRXLHOPW+9y6dlvlKCspExQhYbYbJKtzZd37acEm03LQv5gu4hnJr28Nx
C0b9rzQe6Y3b0m4rBJ+JDJcnd60/32j6R8x9VUXGJvKH6RKjZNSdpY1iPDvhxWx+
T38+k0Lrt9tGtgLEQfZ2iUwe52om7rFRGgkVaQ27/u2NY6fjui/pUt9NhksoDxGQ
QVi8fs0fdjVmqOsYRIlOeGfgLLKseuylm0fpMfRm5rTNhB23nJxa4qBHeBEItD4S
BZRHG7KchUR8/ro63Q9S5BTnXxC5VFoEa3TcSLsD4PaMOMio0ln9UBZhgElMI6XQ
67edZr62+yP4HMMr5nbL3ZK85Xgq93LDoH/RF8IdNkMVD3rFubbD82GQimbRbm4w
4j5aMVXpamVZVjDcN/M27xnAwO/8yRP3C1Ch5p5hVnJJuZ1useAQ3KM7dwlbtp7q
oml1rGg8K2bPiOTUI386WtT7TY2H7fstDu6VyBM+6BYbNllH/396xgCmPBiQuOW6
VOA30P54GU2jZtvDn8kNGt28Zkv9hb3U/fLyq14+/gqKruCsFmkdoucWRyplTnSX
UYGPT+vXerfzwAu3OIYnvJnFp8AfvRoZEnBv9K7sTm7AWojRqZk+QuhZyQ0tiebz
NG0cWko2U94ftdcUP7q1s8EQC6x5nDXb1Jp4G5cHaozSOSMss4v4KW6F4TmOKTw7
XJFkTr1cERQX7eMk7BJmK5eidb8sf9f6Wn+gV0/HiKbIz87To2r46Cit11oaDvks
HADxBPD6lgGI7a5eCq85FWLCiet3XNXEXbJ6UjSzPNg9AbKjfjYnZLfTVV9y37AI
/zZDpTvWJkB/rgBtfdkW2Pzx74eBJl0ZMbsrbM4GkLHI2+V+Y7knreeltjfWSDlY
rvCkzyTIAtVWME9aeMcjIVW4Apnn1H7njQrR4EHJOMVYP033HGtXRDd1oaqUGsbS
b5A5KVJ+iV3apWYtMiVXDQtuWu8muHjnb7cahP+isnRoolh/Q2qpeMCoOVKFLSAA
9N42hfQ3vpTBrIT//p4PHhkvJo9bQXGiIsEM3tr/GOEhnzUABdoZMTLjExdhtyiq
phtHJuGxSzef3SQHeyqhqutICBwdcpirvPKsFGbzEFUl+JgR+rPXbItEDuPirjmJ
YjXImHr/KMffmMYlYEQRCoaJQ4fkGCTl8HudXwXkUs3HDQqV+2hBttn93QL65mLR
eO6ndx+Aoo4ZcSU9EYbcI9rsYhSp/0PIU81B/D92wuASeYGCFXteCxRtTTTKy3df
ShR/dkQ1+s/x8NtHzwfj1J2JcVcoQ+jOPhT+j6U6QDLs5DyvSp4wr9RoSTWpOP1u
mJQrZZ685bZcfoDJV3bjf0sN3O11f9VS1i1p/6YRFpIRujmJAYdCytK9qcs+VdXh
ARGunpAbLiwSMaR+qTDsYu7CsFFsRQBQXLFXu3l2jZBnCk+3Xng/w84thRAWU5Pz
R1kThwTCh2RJxbXsRfbTTJIXedcf+BNQbZ7m4rV39PdQAwcuxi4a1USBJap2YlDX
kfjmzOVVHN77UJp5MhD92GRoGAUfjv0BZN2l5AAS43qv+Y7HuZFFWoVpr//micBp
fyDF8ydzmH5u+hGNmqTSExHO6t4UkzGfg4linl7w46Spk6TVzEphZf6tCjBoL/NL
WRLkDEtaeK4zqHGRJCNDqlLXv5tXQcuFOxvLCYYGWZpLxsTOPrdgA2laWH1fTG17
r3agXBBLNgJ78J/dC/G7gAGC52QhYwcEJKWD8HWomlzt0XVzdumW5HwA38+aTi5r
On+b3RvDWZ609K1B3kvLHJQrVUgbI3NkvU4CTsJaFsCgg07Eqwp5ghwGLJAg2z7F
RJOkieBAOVm4u0WRNbpDPEYTuaICl/R7QM+3r1OGqlosJtMH+7f6o1MkgAN9HVxj
Mw+TqXEM0o9LPrKBiUH8laL0uwK6MOYso8tCL8HTSda6yzsvxu+dMraLenoQVvpW
tAnQ8ahUa0aLAYPNXqXSA9ekxYE0acQ9w05OBtPcMowICITHtJBVnJe7jr5ntvx6
qcQXBb9zSOI7keTELKzQPsGkU2OVWsQKUUl7gjCpZ7k+r15jUZwQRQ9syrmZg9a0
xmrvNhAyWjYIs9zP3JbAkDBwleAKbpdjEQlbfp7T3Hs2s4ZwjJTXfo5JWFIIy/W4
uCiIYnBEScEx85bYQ0tKvaXL7f+bdaMIL/rZeMZIfN8fFXAABgD3GPKOcVPqG675
SCeyjtV/8RuFngoMhCSA0/J8g2cfJSzP/MqK+T+mYq/dLUWxHJbejxenEca51icO
pHk3KQWD82RD/GkXIK7P98bl58Bxn5VEFj/ou1OPALoemitm23bP18rOPIwHVQ3U
/4bUkvGQQ8Mp/pJTQTR6VcPxiDw53J+1HzWgyCrQpE+z2z3zgYlElqnYvXlcFxlT
1UQMmkzlM+6Dsz1f8qHWs4qxr2uhptDYkjIhvwl3hztGt9TVP5MRCmOx0pHx3YET
GBQ1FHibNm9J5wCATss04E5LNkjWjZC7wgrJWuOALWDRBsbGpjuXzNAGG/+fZqsW
jHkngnFmIdfFivzaIbRcf3KNjqalTpbaojO60T46GptzDpPZqGVg/mNA5KNcYHIe
XyJa3LElAgTdSQFfo/emwz3/VSOOV1mscNc74fi8z6JuFtwN1hXcxsCEW088/1fm
gzY2eR0tmJ5dxsasae/uf8blgjbbNTeGcj+PNmKEbk/YXxC5T1MoorKeqZoCZ3+H
3LIrYwx0z2ZRO7uThooRXqI3uMgSrFQ1JlqYpTENgA2kR5i+Gonf9CnBBDUeBvVE
vlZjRdpMHILz63ktuledTH/qABlBlp9L3f+x1MVPGNvSl1psPx+YVjIRR8DokCLM
7aDr+CXU8uowYK10jt7iDHNlPcqb26/pt6jCgWeaARrC1516roiRESsCxv4+o37z
Mz3kdqYSHMNgRXi3qiZlVz8kxkh+whj2XokZIIrlLvnfUw80y/7YmXaRounAegIW
jlXeJ/KMbpyzIkuJN6CvlavXXif4QqRDvOt/YQVdtHUFG8eltPv2g8bZBbMC6Ey2
nuJQKsscGOE9f9zfEkOTaiwqs0/4TZmvW0BxKz9kjWd2MVGwjYHxUncC2vINMJpG
3R9cQS50j5CTK/4XwrJfn1IKnf/XyUDONtkhFSHLgg47K/H307/mn3rwx41AqiwE
1BQtnfzVBjD4WCLYS0O39G+BFdSiqwTkkSlGkuWsrRJlDbuMfJta40DdPOFihcWg
0d8GhnnzPzKPL0DRGpUzI6iSkc7C5zXUwgusk8l1nwiGXutvnUlS2/vAvOQQU3k7
AC+tLvfIqCDzhh+d3KatlGrbYMtvHgGqOfTQ+bTfM2DTY2PEYxcV5eMcXRy4gBf6
MSNHNL26lxBeZAHYDC49EVfUkSr+UjqUHvTJUSxL2r/SNSKvlmTHzNNER5piE1cr
l7n9HC6VsGfX5mCi3ZDkOQpzNEBfOg5JKFpybx/lyPWQ920i/Suo4T3mew/pJyBZ
BoPjsLi7/SJP7vy1sp4qomvX1g8Y4vTGXvRadZEP3OPdwC9G36fxirDriZvaSoLA
ECMDg9ux5KLqdDDNQQ5ZrZ9vBFEucRoMidK5kwzmoQ0/aV7WDAyRvX74AgcmdwRH
7t0C/rflafrA0SrJXEf9U43duDeFU58xGxkE39AuYxWeQbT6BgvGPlIJnUK1LJKN
BIRnHh7SzBNGqcEbj+7xdPvrxOEhFO4Z0Gx6/ume1PLy9UAJH1dMtBwpBUW7LeqE
vYP0VcyWtaR3SfR8gXWF4GwP1WehmKhchHHiW7AQdMMdxEzbM0gWzpTEBE+3QbXV
S8kyKj/TK0r5nJVHvKqr3R6YZusT2Pw0Dkwvt673bMq3MUAla2KK8HOUsCoLYUqb
ky+Q+SXkA76HI/fqkLEMVFAkCJngK0ZRPQWoSw7ztJf/SKJRn2ShMSyLccefwNUl
kvFFmX94xRksYoa3pF9dzOVLaDlhWyAEatjM5Srf8THkEgOhqUFC48aaDoD9bg2O
KUc4kbf4ItcUJyXV2YfPTclnAN6/01eh+SU1ta0Az2XF4u9bVWcTreYue55/wocK
seLf7pVrLW2/m2DBeHJTr2+GUcHrAJlU1q3pLxumdELDK3VZd4fbKEFR2bBxEJtQ
z12eT7thaHegVXJthMGlD4Mqkj3coJDeUa3j1deqzX0gW6VBp71+8VTpfoLEuNaN
QIFrNP1Pzb+u8/F7DxNCWR/MtDCBBWH+dXr4ro1qR7RJAyCfD0afNm8bBS1fjcr2
yIqsQBs3kZB/wCSQpD+ixd7j/1GdhFRWIl/a9CQsuHQUHX+G/9QoOS8spJZ9oMW1
pmr45xlmsaozOearf7d6U6FxhCtekVdaN3XtY7GAA+Tp01Hzuz9vucBPL/Dbolh2
EU1nsRU/qOrmb4no8SuV2DYARAA/Nn5uDCwU6WZTIgRf6+6/4pG3YGzMNn6KJeTm
9K0vdh0p1qmq6VnvTSb4akHpSV94AHAzvtGk35naJBoMfRBcl6o5kNMuGH1+Eock
zGT35p5wHowTFNtDwWFXlZ0u124ytnJOQ1d/cDfQMtsj6d2/PyaAOte3i3ay2mmv
fSP0fnL2phm4JnXmxK6sQbd/fcT4dGI8Q/a+MYzEjqY+ikeeEjHeXSJwwmGlX8UL
oMa9uGU/ez+bf0a3okhLVaNyqOv/wR0PpELCl9wO5KHWw9f+gS4/e4P7Ign3hPsw
OO4qSmRLKzeFTAxLu2yXXWfzT2mPEPsW62OXdfz95n/f0zET+f246IZnPARiBW6o
Yd2UIBLIVTHXFZECAq+aMfKly385q4z2WFz9YuRLNuLIyzzy5ZwEHNpSQohnn04P
lgHmjG6tItFUi354TXNQyIe9eCA/jarAbDn5nTkAgrQARigq9hhVWzMmvQO3Uk0h
peME1UeMCHko5LjFTfRg+GhjSWg2ocGkJEnalGhuv6K3ipn9/gN8pEofWu0DrVLi
j29ZKfwsaD1eIQxApvHKbnhEJwtNxslCFLcPuPOrWX0A9JLdl8bN1sVUJ6IlJ21I
mnDnvezDfJ2Ah7poo9mtFaDdl6cJdezknZg686BcQUB8xRlljFHTqw8iRJZoU0JH
nRb35TlNQCSHMf7IHJA4P1/7OTKX56IrSNHFl1fnGl8Juk7lZRiqYTDbRxSFOqNn
lzEcSB/8hrC/3UpCxaOe0o9lf9tTD0asMjYsLpfoq4KbP3bBRPYmGWK/LshpKHZL
Yw72Jnsd0htfWxREQSKY88vj71T33rsTF78Z6cuo4m+XkRxRHYnBuF45iR7okRZa
/AqySbFH2Sr9SPyfmhm3rkyIIMC9TeHuIXKHHtZ6Ybr5sCJ8tHNJZpYo+cEAweKD
ZsxOA1lVtOg+tYHx8QB3fWk3hl9BE1pLpJUNN+YpO8yT/1LJmopgF2Bqy8BKzHvI
ZmS8FPvNXnwOOmpi/fe5emGba3wWpwhyH9ycUe7jHYmdsqyETN1FQouWRDA3KNwT
l1eVappf0gfqU9cfOREWVAjFIssKEtpYCC7HWph9zHa355qFRIvIMN4xV9cBAZ8N
sJetRozi81N3apY0xi24K2gUbllBwe76I6kBJk5R+W9xIm+THDyepuhu79lXjSan
jajv6FSOJ2dRdye1yaAmenL1Bj/nmE5K9F3prQbTGNF8UbJXhFcqQ69vpqYH9XpC
gqZd+SqmiSkbj4z7rmRywA46hgD7yFINsqHzIBbkyZ7anBd55vTpB2zYN43FpYKK
AeDcnwR+cnavfj2AFJIgIObvFJrZnA83t00mK6aD2+2JPbX3lpvxwQpusIl+UFFj
+EdV7HiyMNUPD9B2KMgtAlDbGy/Wr3OOlTHiN7s2kHebSUVcDnI+Mb40B/0aId2z
DcgsodwExUy++S1cpUy1pPAo53x3MMVVrN4mrQY1/2M67Oo1YF95LKCUsxASg4ME
O1HUlzEBTUMLRiooKmL98uxgOXvty67Bq8VxpSRfVfh3cv/mEjRK9eXQEC/Gw1x1
XXARvAta1lMbWiVq/lvtcQoyqBjMcHO7/amEtj5u8wnVj3dpOkOA37Dg6gzRsNRR
y2a3dKAF4w90CAg4nh5GhenRIIf7FvE/ygb086nCDJZclnJLPtp29jNBOjstOzSa
WwbNyNSQmIVhyLzSweg4E5lKm1ZCqvGhrsenOBsNXzjqVOX7OITuxn6hqlgY+l1U
13Lq5tAJRQ/XSPXTeBpxnokj+KaCYrD5rWYh59lSe/kJV+sBjUxC9UnLbgZD9ee6
QhKBHudouxkHTX5jcw3vDMtmOAMtmX9aJkjHfLuq9HbsDadyY5PqSqQnb8qBFBsY
ju2mro1N2/5T0Us8NkpaS3ckxVw7Njyqgvr6pxm5gn6AYa9rnAdrYL1sIzgZo4s8
jt1dOnHBWeDxwOseoX4GEdx7iHP2nAIKD0tFG5SVIdsbGoqbu+tEa6wuloHuIZoH
ieXEohY9de2xC/fVlTLSUoC8u2X6b1ObUznQqqRG8OAwrvrDmcNrhWSw1rbe8HXC
c5116D/MsbxdaA0e2R6r7QBsSpB8jfOm+OheH+znpbYIp5CTbXvE0j7mMC203LgV
Rq5WXCeI2ITyLYjiXpFl6doF4JDboq74DBaBakKXUtUWNMYm9Ka+Bxgs9tBffUf9
kr4vtMONsQ34hkPTWRak92owW04qGzdX5z+i1KRRvNvwWWO7XLYJOiiRQggB3F2q
ZD1uManBWjNYOMbTC2egEmE6wuNyB8dcmOdpqv6qafJ76rLwQb8uCeQXQKWhN5vD
Px4gcksnpOim6vi9Sm4iN86uIV3SZ/s+kqkjRKNgdrQg4RhxuNCHPYt/ESX2dCSV
RVICfiZ4O6kQWAuZdc4GOjqY7Vl26i5ZmUK15zcZvE8ZrMjRgqzFULQJ7UO5OIbU
dZ7ipTb17ULQ1f2hlRET1MtyBmCQUu6JyAeDik6ZdIU4gJE9ZLHj3cilybAB9Dvo
78DfSV4QSb5K0K3WkO7aybMiX4R6HXgcfTY2N7GSatGKLZiAE9MiNr7K27rhXwe2
VRnuTYlci+/5GVubBXR76aXi+1SoiCr/02bd2TBkzyj7xFs7LBn+9c3d9atPy9dR
fVoL3w2nrh17NHl3PO5o+i6drIk0Kbo1tSjytqkjAKZtHLytUrdxEyWfe3etqxXK
nZ4DrjN8wKBO0wiOqYZnFjrgpotCHaUB1vxRHCNi/5yq4jhB7nDeyS62rWcPttTl
lKS24y2qv4GQ38gIF2QMgMv1MKUxbXapTxMoCFEyU7FDoQ0XJbNj6tk/Zv+iLc8f
fkcT2ta8DnRWB8ho5RNmq60I+1A0chdyEtD7PVp4YT4+4EqevT/1UrSu46sGq2IH
RCLHzbDgoeo4CUvhuxpgBehskArvxC8NPGHg9LzyuRKa2UulDVGLovFM1nD6bfcd
h/qfwY1SG95GyW7onjuWrv4fYhjlnuylz6pO5XQBoHucrc2jQP5qx0olqo/+6Cy2
DwVFXn58zCvkNDRr1WjECjmzK2TlrgFxU7Lqq1TjSnPnOyQukZbtMH1Ap352iUqU
ES/QuTgIRgHn4gUIWT27GtbkbvChmJ1GzdmzLkK5HzefzrmyEg56QMrC4ROgnGhU
q65GmS/JuAkJC9V9MR9MpgqB5VjxLfyeBolIs1Q1Fj2W/e8+6IBNV+IUgwFG5eyg
g8FEmY6C9xehf7S47FqLVydzxefIzJ5u9Hw5lAn7CAafrDo4/nw6XFTGF0of++It
hWtCmOLlVz3++/LsmHS68hRv19rqHA/5Z0LnFKw6+mJgwnScg8rQveXGhBIjEkb6
A/2m14yXb1iir10omYPjGXXCIOJPcypLDbEHBpCcGOpEobZBVIujPer/a9i48nxW
YqqwOKPGoTZULnReAZ+qr4orR+ss5/3dwEvadpBHqJM5ZbCKPHi5vxNJiOTEFVrd
xqWVoj/3CZiUwcyDnoWtAHtRk86GuF7wRU0Ewxj7qcd/U/bZRTCRezpAo9J0DaI0
YKFDUArJnI/C8KqSwjFxOvcgtGksmdzRQQ01I817Chh89jBYzq/tkXZRJdQWrtIA
1B2CV5C5PtudAYVHDg3iw73ZMQmBls38cUpDAagHfQt6I6HEu0+glNna5eoiw8c9
ElV3YjZBj3HKH8D3g1lYBSk1gkX+5f2gNblscvXOFbeyuYCP+5iJuMOHHPcKOIPd
6QsCooNrCUkEf5SqACV2/eDRa39kdSVao8Olw43nHuA4ZKuHzk4DCF9hae8vF4iu
ag2BdH7tKdFvEFZtThnNnDGSP/rfJySp4gF7zhyNu4hF4zSVue3dBRW0B0BguYd4
jSIS+g1Ggx84UlATpapLVbNpGaHUoCacmh74OWiZb6aGbYMqcsvAJseou3wuKLKo
APpP/BjazsYBSyoV8UzA3pH0hB+9+rT5JX1mJ3tZ+QGR8+rLlSthG2ypnUk6ypej
9QkumqmeCB7tCimzKH/utR47cY51Ul8JNpzAaRt5RcCr0wQpy01XMF+gkdGIsk8I
79yHUY0bdU96gTWywPCI7jPRH48MaAfizKn5mDTI1jccVt85byh5NLxwYcepzK9G
kR6BsTANqs8WFh5PYFzI1mdKnjcSmq6jvAkS6ZvSFygy31gI4Rigf9nZD0N1dHQI
aoyWwqEtkCz2q69tQfDqs65nWrSR7Einko5T3N4Df+s3UgKbEmspChuZD76thE0X
pptH1ESO9Jr+r7PjrUhGRr8zNty9OWRJZoHww3QpYapkOnE/L3ukexaTr0lsChRL
Ol3Q4omgomz1ol5RvvxI5UfSfL9TL9LnBhKQ6mkNl7xgQqgUMAk2+gnVDiv6KrKg
ZNQZ/jj7OsVOX7p4g1mQDtW+P73bxpPOTqqT5a/AminX/NiSQ6m3vmBAioGjCcb7
pYF+uJZqs+L+pFc/h8tQJur7y/H3Rw1LVgMwsfM9YJZHoN9wemWopRvgjYiJ1qww
xbhZKXWy/2N1tg4kzPCWk3hA7EHPd2K0qlYIHnUG98rEZfBaP91puBDIpHV34oas
pnuwFaZjEgFGYOKI0JpPKktnEak4SDoSGUclmyZvZuuK3ZLBxj4GXCbrcloCMKGn
U67YBchu03793Y5kCL3gX9brIXM3/2hsevyUfw1XF9LgaFaSB2s7uyE9B7iP0x7z
r0F2wZR8rrfhb7QCgHxTCjlE9dTBBhQsA48EZHuC0cgx5aIzmBc55Wd7b6ohA7fb
/xyp3cQglzVRDX1VA9ry7BJOYG3NNWyYRPo+OvI/lCQe/cy3bmZXUHReVzg2ahbU
X+8WK9cB1X4h9+viKqGgLPbbcg1pAtJr/YkIHmf9a1AzGc9Po3KVtrhxzbkCFuXu
kKEnEm84N2werir6iQIx4K0sdRQKP5EJCDOFRTY4Oy/SO2QxiI2wIoFd2wso1Zyk
uz1SjVqzcXwEYYE61MYcPQZmHingP6FQrS46Q3HuMdLSno9zKGQDaljHqoncHC13
I4DXW/jmPsmuAaB8lIiXGhwNnc7xE3YgWS2oIWt3hKsR5fsdlq0fA4Wuy3Php9N4
lvj1V0C5Ps1BTwED5opNaFR+w7Mwe7iGgaQZUmlnB73hMEHSVwOXLAwffl6rzWyA
ofLn8xpy7N4VDik0/MG7FRDNWOALCiyqYMuWV0cYMfwVsofTv4ixkkhsqh8F+hCd
DDRFM5hWAmXMYu/aziI9kZZnryLLxKJRtkCYJbFWp5Z5q46258bshFj1vQLYEkxz
6HYkUbgh9m8ug5UybqIrp3LnNFXr79gdiLuXdhshuqP1tc2NaozDIIu/wzrtp/qa
Pr+UJrH8x7RmiHcD4LWmVVIOS0A95ItE0BhxueD3Ou2oA2aXLE4Ufp7JBirT7YMJ
W5QhK0byOHPJENo6e5uqenpYa3BjFjt9TSF4EqkDHe+C9Wh3Vbcmfe+hYV7nBU6d
KW1Z4g41jwSnHU3E7kICFi10qHClNTuNXzZQpFkhL/jfghG7yiIGDYisqcevCitf
o3tMw47EUUS15LX8+hPAfw0zRLVW8A735oPNOy4k5ClHSII1htLzsyT6cwz4FcS2
AO5Bo3vV5YRK4u7o/EoaS8+TycxV2l9P4r4V+M8N7R1LdzRvTtioH2l57z4Tmgtt
DdywjTHqkxLeayRIcbtnlzYkzikXKb24PatIifIxt/r7LUYatbsf5G6Vl3mQec7e
7LOlSWZIh26DecMQzUOhbCwsLboFyU39d3+/FUAdqsNQioEc6E8TT6vBa2qRq54r
bNNKV2RQ9rFegLaWnScclRfvtE9lWu1GknjkiCv7j6o7uly+kDU4DjyAQ7Lz9k9W
2nsycXt5mgja0AkyJsZET1HwGQ61cA5Lk9a7iYQWNgDyGXiw6erQ9CTkjaCj0gS5
c/dRd8ECwV5PKnlkmUqbJMlw0Fl2OCGlfJZ9U8ZINdk+yYy5N47Q0IOCr3d6k9sC
zvFfBeJOZPmDw4V8dUmj+HENkvkkMpkx09WMPdYyvDY7n0aUeo3FpxhOOw7v4J92
87DiBBpikK0075ZN9V2xOQxlxHVeVrkbr9fml/Omg+0hwCYT98jQ5OSnOzqZXjE1
ul3owZ1rAVhrts2xLP5eknbPTeCtftYWL+Dq8trV339zQwAqrDzs7Dd0RGaKFUkD
mXMXT9495EfCoxRgbZgUalHGOk/bvISBkWYUxdi2BLo8RF2TgFeaWgJE4gp7nglt
CbUjDL7LOfZ3wKz0mFcTPlEAxSjCWf7h50V6bl784aA7VRl5sesnDYDChwrp05NG
yKRO08NbBz8hfyj0Hm9stDWQFfUjzDUcKdUu4lGNJ5iYx1csanyqVvNYxytMiH00
MkXNjfu3J6NzRri0gNZIz2Cjs9sqQ+QLMvX3IHmCWhpExJ2/YNzjuROwJD1+vup0
5U/kwUcqQuKsMewPRr9qNWE2Tm9gGj28MXH1lygF83dI2oSAQgCaogvnMKHf4IKj
SCPDuq6KYcv6hWhiJNEoD897PXUz4+ekvPYIFTBNngBqTh3PNgtRJ6ST4IcGtDgE
nn+TEHOcjZTtXBMOvt85NGRQ8gZmmhGiWF7vKzbobn7YAq3ue7CS+Ku2EhrYuwub
mnQthCYMfRARBxB/8isNuuagG+L/fsRvCfVQJ7rBrokywR7wvm6MKHdCCIN5xMTN
1WzUyK+JpWx1fHXJe0b4EOPodJ/0HI6dxiz84CZLbCzkxbdKMN/nQjJxlWoE1X/B
iNCg1ymzJYF3vctvmQJFZIrR5Bi7B2PZKFT12lP4EltsUYeee0V16yBeUBYl0rcB
xeDHo2Int1rmx7sKh452pfnMcgNBwy6pMHMIHEYTRm8sy5twzxpH3vnKNwjimH2h
qL4zdK6ftS5gFCt7+Kfm9kzQoRjbvGNQQ1L8g1H2WoTzlM8MYfKZMsoWLW4hu8VI
vuRjU4tTBzh7UtJ8LOb6LaHlXRsGKwhX+nnXgVxFCAFpQC9tx4sFt484EMu7XnnW
wWBgNr5io1FNly3dVqLKhpq7jJWX7L0I0wzbbCoLIXBNKq9Dlc1RxxAkcs/hmoLp
d/tetY7wwn2b/2k2f8h1Cx1jHmd7weWi/d9QfP0tzsnvHNvjYI0xmZk6fj3G8zGs
tQ1NjfPBTRWsrqIw925D/94qD1tnm0Ss9HjLdAga16vkSv9UvbeAqfx3i3gPG6pi
tjqJCWvjfzG3MFqvkNTrIgBasgEICUbdDpFHMthRfdnUBdyqh/gJcRATBxRmB+xi
5Wy/yGC9xYGYQ1PbQZw4r0Micszo3Pkp3x/PhsStzVAlUGDtYgRzB2SWF+EpK5DL
+GNlILShw+Dvr+1sTEv1waRNUcjB1/wJOjD1bb55n/Xex5e4yZsXwu9u/jOy4Oji
XdMILa3j/MLp9Zt8zzzeic83ijCQwE3E5ekVLnzb3NVF5ftjGoASvasC7BJCIsKo
NcNUeUX7n/ReQ/BO5B4TLZNxCbbX0X2UhpBiEwPJ6NxMjSGtOPOt8zFihiOd+gNu
2YsFQ5te9RqL61nXm4p09Vw28LBFrHlB6KPTnBvDwKE7ZSfPmSJ+gBv1b28jRV6g
puS6i6eIDUh6jwI10LXr7RJ18Eh3BNXmdUAPMMDyjyVVSY6bOfH1uA/oCrzgyTZp
Hus9lGtnePx+D6EYNGSVR8iTJ3tDec4T5GvNJgMpQGFZMNVKWBtzSnFWBXR8eTYs
najMlUgJggtKW6c+lHTosiVZNZU5DQM/QU6pzWINVvVpNRkxe3nsK3MY7HqxPkN2
ZpFsnKFjtm5VxP7vrgfys9JMpC8MBUoWFw0uqWlN2N4hWs4iFyaL43VcPGUdqSe8
F+A9qmMzTe+aiuQgk+kD8QtXGuDuO+TNZy6PGkZAL9CGrMJ6rLS4CJEfOTfb2W+o
klAz8UYdkEedjD4g+1zvTHakP3Hs8VcBH4qeB7jau0/H1Uyxq1FkP42QPCVfDzqh
S36Emj0w6VpeslslZ5LjiI1BDRjApOT6BtkcjSaSgUfB8ETHTh/2W0Ny9t5HtGkJ
RhKmZm5dfcbEuS+rP6xrSRbw79IUvprHFJrZlzt2Pbi9WtDCOptHO4HdXIfGhMZk
P/MV0HmIw2W8nVQkM38p/gCeq4UkYZxiWrMj+oLQGZdkhwncqNpTgmEa1dySNAj4
4VK7uBi7ziJrs3SiUL9atAU14rT1e7Hlgvxd3W+144hOdwrA9RUN7oHp970JTPAH
Y0ibg1m09fmnx7FD3Qd7iX9VPpUdw96ZeiRStAziAITTNTG37RpCH8Edg8woI1Ec
0Yx19efRe6BOL54LWs8mcWYZ0RMYUv9gxwlNP4waDITL4BQ++oARLeMDXwgB34UU
8K5U2v3YHLIwMjSP6Qf8oOKlFCY1VK9bFMFPGKSAIPvY437hXWEPRS0F3S+s8Vnt
+bgOl993yfdfHcA1SszZFVXoGSdkQVkaMILUGUIhMOGjTTbdVzldErtnveSeCahS
QUiiDtxWxd4L8MiQ51UaGX/xfVWs/3RR7FwVf4m1NZ3y4jOXpn0VieMlIXh5Ve/L
9wf29n3Z11ZI2/Hv04roAk89qWTAesT+bFLEAl+GDfrLAyOxUU72Jlw666pnybob
vtnEWQVfTF15ZxJ1QgKW7Gye5gl8GJhyofQ3PiXhOozfqS2Gmytln1UjI0Cd4heP
WeUzJMCLPSv+1rdzVHQ/oPUrCs67gEUBvi9ERhV5LCrFFLL5y1+3uoZOyK9EHcvD
NywwAY4rdUsZxO50+JOpsVq8ubc7xhm7h+XQhKCOVj8Tk/yjnVCuzcsNl42m7wsi
I5QaeGcvCmVGYXl921r2eq7AQtPvYSmjzT3czIQaarReLVkyV0/fA0WsKVNtE/Vk
CD8O6vr7O0lavDeQelhDmBQQGR3vXEqN26ppLnsXVn5yfGNZKGQz0uEzYLypRT3b
HJQhQ/HTjKX0T+/BxzoQCUfAYlhf2wzX+D4eKeLDv7mbUyv4VsZtuyVbLf29yv6C
hwh1Y//sKqXXhAKg4hfoAlqU24FgDU2qasxbq/pz51rWgXOtE0prinmVdjZQDR0+
ipklrhXu8qpEDkDH5O3xXZHg1N+IxjsGwOkTi4dUS5mIGfAhiH3OAJKZu5XaC0hh
Vn+HU6xyQa/UDrvcumvfpZB1+IDXnMvMxg12icWLmlzT/pCXig+BSmrMXrxpDYJZ
sDQZk0RYiqbiFfwpXFLeN8+P6pomd6QIulH3OxwSYzd91TAUz2w4+ldxDKIKOHca
uZ9zoFuZjI5bvaqukbzX6R9dJj7ZRSeYn+9epgRTRGfnLbDBBoYBwe9IlcyR46wd
UKkQksIVDm/3b/IEC8DeNM9rcKjRciC4Vu1/pFL2q/hyCn1/dyC731pQPVwmi5/r
owE+L6BK/hwKKjnJWMis2lbdtnLMLe/ilOFgKvcLxAnsbhbfAYB3y9V0bgBefG0Z
xsmOYNWk1J1DoDwQm0FXTTrY1lctfOOS0QbE3JjP5wZ3rpuKjoMUjdHk9JmudRRC
yHOC2PueqYBRQ6HZgJ1ADc35aerMG/aC0dLSN3v1eB7ORggHdfnSXsmtCD+7SQ6K
zjlmnGJREnO8O/DcwZ2m5+oRsP4txOxQocTY0zH7vCHgOW7tW/x2p1J/+uDbjv8M
OFkBLiBXoxIC8GeVNCcHtYFohvTq2NIsjV5hnhvaagbfRcTx7X4yqFgI2y0OG3kJ
USRS64iydpj8Vw2fWKXBId28zwk5ZPFF2oq2/nhYhOjoCsDevcwFOF1Kdb4HndH0
D24nCAjXituZQoxaNwqTOXh38COnqQFRNy0bpqKX9eNb2r4Q+e4yeU6/UUXJJmfx
fjO4KkfKp6IBI9lp3B44C4S6yfv0ymlX31kDxPXCNSxSD+D1UbKjc86Eauuy2rjW
5/TljOOf//P5gYaBAR5b8CgvkCko36hOQVpV82ZmubE3asemNTYx1iyGxUgCyLzp
aNPwZ4bvR8FPp/deE/FaPlqhutRG/TlVHIWXS8Pl8Ck+xcFfarZU9i1B0FwV2X7J
fGQ64DzrnNbR/I8u4N1dzAE6QlIcPO4eEM6cODJatzWYZfzzuRI54Lh2HMLQw40D
L0Kfd8dsrqxKxToq0bCFZG5SCvIdi+ihfZ7l4/5xZTZI/Z5nUxLr70PKZeDGL6Eo
8eIU/1Frd9cCGAO2T5ZLYB3S4VJncJlWqz0OQGv3i6DIILPslp+mHisFP3um+MTK
a5eSkur5RmaCvKOEcv4cKDoXPsYCBvB+BGvG0xBsvoEnJwQorgaVS6FTIWMAGbJm
oWYBw8b+fighrtdbwY7OJjMh8U8UFwGMh5wn9PEtktIbX7E5uXiNXzFkBx48cxbh
WZDaa2SHAdMDZWhBFCDE6a2IslKOfayNNv5O53KU7qzeZw/FyZTtecYouNX932ZY
n2XywPvf03COpSiAAOtoLKhYj4vxl12GkE3uhP68EuUm8H8otHlXCtiKKOhMUUXl
X4p3DlN9iciSayd1wj+YhFF7UCsXRgXdD0oGNvog2yK5Bs5hNraWsMQ4ZmI25Toi
KiRk5fneQi9I9EVMRhwVG42rj+x98H8u27+51oYrAnrCZm/zli2EpIc8xMtREE2v
FtFCJvMWzRdE7XcHC2YMveBp5KQ30CMfdIlELhg64R5A5ri/Ha/IaBFynL8QJIX7
HZFiVnItj6/Je6+S3o94p356fx0urRYEBBM1+YvcApr7SIboPownpbhUPtgef81d
QDsvPwHWqHsqV193flSq93kA5L7dIYnQgh5AaRzmOhQsAb0ctgWF7yCMTJ7EJvL5
L4Fzy9t+KuDIHtUNDrs8CwIeJSUvPihN/+LcXZkISnZhWQKAUFSlXrTwk0Bugaqy
AqJdFsUYK6dG9yupJy4XI7WZmQL06uo9q7iKAEKafJ34tOESyoX4NaAG3II8TDed
HVepb3ERsnsaijgSLEpxE8kmRSJMKfCpRGOlYZn2YgC9IfXUxDqJTHKQ4QfA6AQ2
/rkI/sAVt1HvuNUV3ZgJQ93afv+82EWVuojrxEoA9+zrHQuQwalYiiKdRGHRKEY+
ppFxXgwrVSU2yJAIOR6iR9ZnQoruJt9vakqL86voTZ9YOWR2KrwKgGchN/rrg9PR
m2p1QBC6SPRvtGKln7RQppZOihWkXzcT6byin0MjRLn7QIWNamjjs1trnFdfF7fY
i8mFWWh2rWcKecEcXCdAAuCDQ+Aij2PnSjj7QtMezJn8ToGsTNKelrtK4XFsXFDB
CHvpsrtNo/KSnUFgMNZK+UnzBTnDfq4Et3dpZElrV4u43SGpz6RDf9Wjh6NPedlj
+krVUjBa9HF3NV27aNlzvLMd1Zk5bjLRLyFLv+P9GmcoiXQZyjp+JMqmNZGdkFgY
hgWrZ8THB1CczhTtQA+VGMAf3Zuj0qEoJABwojBdsAIlzuNQBGAjTktbxUKHZ/2R
VS/6AbDhCp8e5vdtC4iRb8ejvuKlpOJGfVx3/3zBh+hgQ+0KQzB8k57WlIv1Xk/x
vmZ3n4T9ezzQ5GPqwuzUh8pkJosOFMzdlDPY4rX3KxhD2PXw7MyhWY0j9oaO3FfJ
lP6Mi/nxB3bnBeF+4z4BngluhakUESmCYxiYz1fNk7XA8Pw+730sVjraf0jKhxYi
aOn6VfR51n4BhLCYvfhQ8fi5V5ksmQYCluE83/b5s/uNcJfRgXFohtr4qkEwljUc
lvxwUDtqxoIb7omKzTQ0Po2vXCIi8rXeodQBCZLQljGZfITGq2fhAgQsvOETHUsH
6grdRTyMzeizAybZ961nzFLS+kjS9tL5p0WDs7M7EdNNR0NkxLoGAiXS1kmmSU3S
jN2e5nnASOMZcJYTlUPlAovv807DrtpufZ4HspaniOObNpHDdvEeRxCM89ZTvOkU
BOeeUaLvTL9FaxOr5ToFm5IM8rfUzzkXzN/FMYE50AKZxTdQZ2LtkUva3tM60lRu
1057bcEYXZDYCeGL5ZtFkm3SXlUDnLU3UOKiVxNVgH4Ut45aPhfHiN/FSWHkr8xZ
LYnt70SnmWKKi5JdbxSQVW4/XDksm6AvDGNjOAbfumuz0SjaX08p8Cws7IXZk9k+
udVANeXgtq5Gee3eLFtrfw5v09DS8IG08YuhsAO0vbci1KYwiR/OeW8QZ24zOJ+D
0PYPHc4CVl6UTTLE2xnTnrCjMHzxw9A0UqUxySkb/UlCro7pv3TSgIlUd+XtrAMt
naUt43Yhvy2uJBQfVijqgiNq7aHPxfO3mwbVrMX5lzp87ARKiCfkNWNh6aWbus1O
GqUq2IBD9lmA27fttCCvnv9ZOHqVbTF4pPSXwdXy7quKXyZ07JVSbQJtVpE0I3HT
1q16mKKmgocAV7ISmdBhT3o4Yby8rRVdhh8WabbRV8v8wKEVtjLRhz4QnCdgtTyY
0Qy7wtuGEJ5VlfT+c4QBQJKBqzIaVAuavpJjKSJ/vpSvq3EZ9MqhXiJCg/vvX0F9
i/IvDRJ+nYtcCXPxYGMdn6inIX3y/2L+OBpcwds9bTl5i22frvlwi+Z9HQB1WUNd
Vm7mzNjF3s/lLxfdG888Wm8PxZ5xrHcb237v5//bcr01lveU9GLIzIrkm20F4CXS
rj7nj3t2LECdJ27peJMP7Zdp8H5LPAkhG168xB4EjglK8yOQ7/Cfnxc1bI+oQ9Pv
/yvtWnrEfUJAbiYv8yJwyIjOYpO6Q5jM490GfyhI+pdpZSOkUiZ63cPDYmNdQJDG
LrGMw4m24Y/YF7EO6z8fRQsh12h9gYQvJSXxAFrqtaAuPhSzJXHpLcW//84zUmua
5l59Jr6gL8CriU3ct3Jj3hbIvU4MiP5MHZZpamqPHrDbw9KqscyRsNl44jE6JnkM
QH1Smg5iXZHtdJQTFAsqaNFFsPu9R8pBEetiv3+DEdE2Z3Eujf6iXjLMjPg3C0DM
XWu9ptJ7dTYm7xPQ9FO9zC+eraJbW4rydfyGPXcoMxSlAQAsxuqy2AzAp4gxRh09
0v5FKO7KDPgPOHbq5mqOoP5Hdj5VQCGHIHMd3tmULbzX/frhDpO6qle+0cJZjADZ
7fsCO2OUf1FqOd3VoBOnK9bwERwNqmVT7/22HkLTUiZcu1z+bCYGpfubr87DJYM8
VkCvFPRmL/J8+P4Y6SONI8wQb6odJ5jDDrXi5Y4eZc+1az/yxXrHHA1ZuM0GQY/r
DSUYBq2jFO+Haf7AlqiWSUWkQLrAGdo9CJXtH1e+ovY4CiwzkuH0ED4H9bSPMCgK
3p96UhJZVDay0uI5NrBOFElJl0akHHcWKLkp8WyW2JvCsuRpA1W3Lo8skR9X/NU4
9OHZDvBsPTAc81bB38L0XPdPzvskiYVbUcI/Rayj28sxanK1jEALULig+pWUiQ6H
8aM4DV0ghyN8yztPYTwVDV7tGStzBlZHW1e8AUmkHHXKi5SPNPW+i3A+scliPfvI
KjHIFYHVcPxkdLDLHAsDsBoReHDLParF2tLrCFv9JxlQXrQ41gWQBZC/9WCnXuXg
XV84IVMxameLVVUESRzKNgbQa0O3sh9OH19PcCop5OSG8by85Jxjb5m+514dArYW
96mwNK72qfnUqbDiwi9O7+7We45KSy9uqLS0AB+e5rdw5ZRZeCwUQYuCm0fDTJBQ
CAwm2Nj+6Td5+n/ZW8ySy4rSyt+3rHNC55aZgU5SMttSk22OL1ONLHjbmfz0EGrM
wxEUV96KVoW9XAsieJPncVhQnX4By6EGcbB9LbYf7nMQJ1fqEJmt3yBgl1BP665G
Oxof6Sbx+E+/RVROWBCAI1wD1FKVaBMQxUHKC9cNGa3ms+FG0OUUSnUduULq+ddI
KrKlpIklp6N/nk2w7ycfUnXJKppuYO7o8UWI/BLQXahHRjePmEXAyYx4k3v3hzV1
Speli1sE/Zlrpu9eH+R8XF97jXIMBq35gUow0nTPFXcIbdMxPndcLnOaLsR/rr26
50OM7DrcFxQHh0vSFAAUNKxGxsRKcyUmQoOdmz+O7mJ68B8rI31WzXlu+8fbyAFk
xAgyrAWU4NoFRUhM2Kfq6gv5CqHMkvSZXSnKxtOYTMU/chockKjS9hxq/JO5Bt5H
IC/WO+Skyg9HF7tbOVZhcCDgELR/XgUCWy0H2dXcT+vI4REdB3CSIHzqdK2swvd7
++O6MUqPQ7j/Cd94Fae5Qedcdrl3W0f40IW+xS8JSoaH62PiUxYJfq6ikVBNc9Po
ex12QBRRP+jShHgQ6i+7QVDZtoASmZxXpCNUT21JbQ46Y/hZ/ZL6wBQ2H2/Z69sO
w2ew8FqLOrWPzcDDYVSOhQSOhnWHqR278flD8enzslS3S9JWo0SaxgqcMLb5i8g2
NqmM1q8+mJ1mBWJWAIcixLGgXDLPqY3G85t6BCmeKlE/6SvVCllcW0e1fCVvGvYU
VuIH78pTTWpaRAnFjkxT1Fy8LE14T3U8KTI9U1BNCRL3OP73KV2Lb1sXmudTn2Pb
LLHfe20DDxf/jK/OS6a7EPNOjjptnsLwrA6ehgE2ZI2yx2p+d76Pjx8kNRVbUST0
YE1a9GoKiOUO78YRU92/+3oQp+zELadMxjTujZ8DEUE6qYy4pCoaG3SjNnAexzth
2ulAYdXMBImyf1BW7S9UwZy6Z0E/nLtxDYAEWdAqt15WU7emPNdczEOoXBfkyk4o
EkTZDJnoqPqZAzxtVRVGNXl81/zXDoSVeBrwOe0grvjZnNUlqBNgVKFGJ+rLwqIT
hxVUE3Kfk37veQRU6yvow2uq1lj7YyBUackFx5INCVO3VUrhr/Me4tIBeGbKcLr8
dMTzLnhAcn8QnbbC3tNcLCVAXTv+cIGVbbIxJhZU5uTnjjTMIqGLwMZ6YbzhZcXk
LChYmvC3BuZR4enbNFoboRY97IdswJs4Y8A5dGYo9Kxmkae3+5+0VCKeehT8oSgz
GZBXERc4s9T+LNVE5oZATW/djhcHpYjotCCdObkVnCCaWO3XpBfUrOHbV4eS77l/
hdinORopwTbnOzUQIxCHToRHFn6MsHqU4ylxu0mNIEfZJCgBMLRGgE7s9xY8k41i
dJU9NucsfROzzJ4KeU60cxipTBUByQGEAxX0HuvbwDR7QDhlxm8MrgtP61Ba5p+c
8zIBNmneHiVJCZnjCMDTG8J8IU6D7JQ/uJWRzIvBZ3u+HAvMLr6aY40gtZxArpUh
fRGRMidf12Y7nz9ZEstSQkINr9gwYWxVg0w+Ml4A1352wYKhnXlIe43tH93GiV4Z
INHHCLUQyobki2ES3XZwFXElNg0NQ3nFCH1WumEMkUVI284rtfqAItyUKfKZSE3g
UtoFaTLd/AlHzdcLUtOpsIjN4Sz54AN+PDyZm7R6IoIpMbtpxYvegpSNoJhY3/7F
I3+GR3sEeSmyKDoNVogS5eUqdygOn/yeMqcpiQx/4TNIuHVaoit5oDZ7XHR11FG9
1GAuaouvZeZRJ6tHIV/RZR/UWOHwMdsA2gcfPtvj1t+zQJxJ0XI+u4PoCWBVZmNA
1So5c6PyxCO7a5+dQC9mPqP3W68hQdRXDHdFejQ/5Qs0PuJlI0KBXQpeOBg67OaC
JXiStpPdOnckgfjOsoiQ80lf6g0eroi+t+o2Cq1LuGv47prWa4jWsxM9L4Bmf9u6
yHWly1KfsPQFQ0Ee2tXMgZ8pc9HHlbsIapA46kH/9LeQ0ZVTi42dyctUDuQBnQep
9WEcWi2DEETPvrJRSEtn6TAup02a6P8/6Sf/r3+BqsaMuBKLXPBVoOTaljmneHEP
XWg3qW3e42M7SyWKH0H5X9Qxs3d4t0T9Vevhsforbfh0A5vw5uN81ciBWeQ5e0YB
0n5a01tM470OMp6habbvI/w1LVaWqD2EOGRrWWlrmjd6GuA2jwvDS44GRg06GZsr
7NL8YKBfRcNIHeNEYc5iWDIA+/cTaXLyrsP7e2OSdUvzz/jrY7mVijVKw/5Iz1XM
B3yUhjI+cYnEn9dTCmdbBemGhTeKXIvU6uO83hhdvmYNTdYRNuT8kQqC1Z0jJB5y
57bbQCJAdtK4TZ+vcrp+zr04P3zx7bYZG1qTuhtNO+m76pFfWNa6tXPPNzv6yoEp
S38jCVsR87HGUlwwOnIIKJSuWseNSsEwiBqyrSTw15fVq+RMwyJ3UnFzF3GVTToy
CuzwP/Octi3ANfRV4Wov1+m70FX7k0qC53/1gbXVd9Cls6i8cp7+FWSBcbdW+Us4
nCkdARN0hFmw9hDKRN8lVi854D6vHJsrJplxRfalB83J6h3JQ9MW81vVO0Gg28WT
j1rscBhhosz9hSv1fOgsjVz3IFhqIC1P5ZFQxU4MAKE+ItF8k7iTtWa97JdmlloB
fYll3Kt0QUlfnOj8qKICTShPZmiIw6Lc2334O965ym++hNz3meZLgSguqbkL0msw
6BHEz1gkWPP273MJBXE+5SOMuv1+occ8Qcy6ksfWA0C7/GI5bxuoHn34z4XDb+Cd
lrOEQMeiKhcSb5COCOYSukir7eOjKJZ7DKwiR56ch7VB10HLCwpGWwpb9641XPk8
TPzGmeyvEQpb9v0pey4+gDAIBgZFgVDJ0Z0S5vugWvu8pxHNFqVLjqfylgSg3TCh
GG1Q6yAE9WwLn0JJOR4XAG/xYVJnL9BM9CH3iI3tWlwd2YL2UjNbIFx9dReCn8MU
sASuwfXbofBLQpfUA5iWUJIAztArWktsxq32hAHtS8FYngEsnJOoaOdpelV/+ABl
6crJyB4romJHSjkMJ5UY6VBeVE1iKyqY70eKS0pfKtqqxt+fp/j81y561Nt0ne9a
9TDFZga3VkLnneulNCNygnV5ChVkdfJqdSbPCAQgveF8ERzZ2WshYB/y9x2KEDcg
CUr4qGHRwEkJ1mDhsGPXI6etzBKHiedD8E2xb5JcR3oRJKACt72IM6JuRUjDTJNx
Vi5ERO0sCNMhjwzbv/nxLl5nQO0Z6ugF+r0qkPv3w0HopZo5bAPwruVyPi0ph7Cc
5KUJonP0VceW5hnNqYrxbvRd8+ebpxeESPmSQlGYvMbD/pufkVffmRYQevmhnnhg
Gm8BLmtC5OIoCvkKh03jn1DUDUfyEddlFRjWta0IKFcjlJ8JZSquxma7q0L9Fljj
GbNlWtNQE4D5xsnVXHRHLfSCty6whNWbUNeSqqlokfHdqSsqligIb/ZTEisSstRM
MOS3Pq1yT+d8yPS+YHz08Mfswi6cRnYYtuYSADnVq13c1CmSdcyNOYqE9hmV+kba
RbPUWHxkLS0z0xSQBBFlT3yWhMCHHlqhl4zTIP23YO/LJ1ZitQ7V3ePsQnO13A5j
ZigoByn+LELCjlOlQ3IKN/lCAE0q21YQB2gDl00dYlGhueC8av9768odzxoO0quq
AG+yVwUcqIK34lnghIn6YF3ObV/ymx3NZ/DpFk6NNry1rJE7KsIIhl/tNpF0XdV9
/eubHpuD6zETje//0oCXI554Kf0NbRza27NZbBc+gemiJ/7tE4BKEURRPVmd7BwG
OjisxDK5wBjZwazyrE42mwcsXu0hdLtpjwjI5A+MHA6WydsgTLRNWHU4efbxd9sR
caRfv3hSiMzdm+QurKQIJiHA0Z3LdIbSngGljdjS48bNUSY0hyZIbklt8WapsJUE
w+Ih6W54lY2UEg5K/HzJjUmq8JEwbF5vZI6OvyV4MrR9yjfhC65C4UufZUqjgSCw
3PJhIqva8hwzqIhNXXmdd9qom6cKspFUhVJAj1omTzTvgkllI6ywPMW+afYC9YAy
eqglPGdECX+xKYr8wogCEULv/HkTi5CYdZNwqDBTeZvlyMtXdz7fhQBh8pvdvL7G
dV33dZF4svaSCSrgLAWaQa5EEkbRzzqTzIqNytlgsYsOwd+HFGPTnuvm4svrUzt3
q4my33PipUwSJv27b6LOkpOy1ZWPFY9WcTHXYJtJgeDCD1AL4PoT9FQXLc4/g+ch
hNB3gp53Fe7zheMZdZ8aJtQaQnwjmHCArtSXMSQ6+/jLhvkhw0OM+XLcdl/xUXMy
dO9G74HCm4WpMsDctZccgDkGbCWQFD3Tmfk+h2j46Gjfp/z0pLKWz5R39SJbIV2j
/SX0xQaKOPYDz/NjnZ6YTx3gfGSbVKHlgpX9juznkwjIiZoYjl2p1fuELaPF1gKc
eDbyw5VtLRmZo3/x0KhGV+R8nE+CwJP3jbFsJ6zZwX2Iseo4HET0Zing2eMM0vZz
STUub0Qk7dsRpX24A7fePgYG41tggLVvTZxEw78JILTVUANjvtpFGgNuqyZpiZqf
HeTnp3vGg4wxvy1pKyZF3BDLZ/SBsXBS6ttGHDpkWGcHNtVPVcR2sZKKxQLxmzww
HbqyQFHSQx26eZ22m+/iio6NoI+mrVwH5Zun4vtJQftyldLLvELMjfSVn0Bfcs2W
QPMMHw8bYVs80oxI96wJt02zpWPVIvM0sAL7L6OgWnrv1bajV7fluPodGh7ctl5X
aZLsUua4yf5QEk8c8U+5twmo0k50fGGjzYVdB1dOkSNdA/c7zBLVVk5lngNY8q+G
3KhuuFrkw0iEfWA6z2/eqGQ94xQ11SDz9JsL+QoWrT2nIiAN547Io238axoIiBc9
4kUdHNRTmHwTBaZyeQCZr2pgBUSbEP1pDT7ioyf+xaC4X7uEfDrGHJH/gtbPb8wd
jwZ+0O8SHD/4tbgw14fToiMOW9QAkMBg2VROQfxvcCdmptdWYpiSxr8SqDbnRwe7
Wz9qv6ukSGZiwkq6qDJe2RFEXMSbFUSEsr+XiYLaTvewAhjujmNV4nt5Hd5zkjZq
R1RHcY1fUp2mTcI9mDHKI7uEiOspTvZFN3my7a7tzoEpTrCxLO7MQXSGhC/qIMFS
aZNdqtACxZUGG/WmyVgrot/9t4Xhd88oHU+Kob7C3PJ27VBN0u3LZYALDS0KMV/B
emTLlabZf1ubd0256wp4k5jHJN4t3RFfWuv5Bl9midxg+191XG2BmG5BPj1qVsb/
kNcqEjHbQGgzMeK6cs36EqfdX5/hW7/tSEkaIUi+KHwjM5dMbQjkdqgXEamHkMIY
fcS2NNM6Y9b6gi4tm8EWZAlo6cRgihZHbat90n93JJQ2Jm+XXyRZ1Lbn7CyGHqsd
I0EkseJMaXn9KXn/rbwdz/+0zveb3c0OUEY3bfgZ8hDxZ0iNBirhkdTf4P4AD+Mu
XTjhwTn4u2rquG0H3/EzsY3fTogKYSNiC1wGhluYUMzF1u2Z+jmu6yvNoMxk3KtG
y2I1bzZYFo9U7K3ETlUjqs5Ff+FJt7gxa2F5FDgJNUf+tMeuEIjf4/Uy8F/omejm
SDRUvbMuewm0G30/0y6iTk6NypUndlBT304knQMlwWBSo+QR4yH78z6c1BqS0yRc
4wmMoMvx2mbaxjdLWjYr0JyClkAMM7ujTGEewv/XqLWqxay2ZCdgGjrXmDE2QBLt
FxxNAYuTvCKFHeWSrw9V2gNYRwIaAP+NgbrW5qFzKM4cSf99nyGw8EI2/c8Z/7TF
SL10KPL4Yix1hsjKfivIYDUbVbHDc/VwPSOrEHYHhgJel402RYl8HHIzqOvNRYwM
AR8UvtOmXdOljDch5krO+CkTZD4b00Gf+y6kvzm8TtILylOcaMnArk/YDu/kd3pM
NkM/ytYe9qSLV00L5jJSqm+FeGaL42wBVAq++09dab+PlsITUAV9bLb/P7GPSxZT
3ddxTjEHE6NhchP5foRQAZEN51gvlPTSJUeyVdzzn7N/MzWmYrhHJO5GbxCqoNUo
OpTd8dc6VECKIf7HFoICQyW1cmnUyFQ9cx6pe8QwSejbaM8KMqm/0QdxEFnB1dq1
bPNGB9FPhW4liLCnKlxzPfxDeV95A8H3pHKBwLYkI/VxLuWoHR9xlsAsBsDMe6Qq
J+lysRX/lueLaXChV6VSHXV3ECHM8rJ3O1eK5lvc21b6t6eypVipKtnV2KI5ps0u
B8Em0AtZcGKs+Db5MVlB46Ky4A+kHw8Bd5J/5Ne7nJvrDE+h0s4XKO+lLJcSoSZr
tl/bpkSqMxAR73R1YSFnaPkQLvB/D4/VmRlhFMTeLqiWhF3tDMsZO4MKiP5/85Me
+jCzaaOpU5MmO/DKX7HUpJ4yFck/VpnA8tQN/nEiAbK2AncZX/PuiCSn64Tftouo
AsnnccT4/PgGFuyXy682ah6hXZrHaqiQXvzkvFAQV9I5Aywret39aKAkf92n19VP
px3VPCM4uNSnNEMlC6gnvxrX0pjSXdVsf878yu5vYqh0apz5bNDK0Q2RwBV3Ueq9
SKVX3apHTZ0WbZ5MXWoNmp1pTnoL6D8OFHR24BFY6/MCv4gPB9HGJDbduLt2m/oc
ELprWmmka9SRB/kmcGCmicilDkskm2X4fqotangu7uKH2FOoKn6OdrYFgkTkMvMf
h5HMZx0VSFKyJISjySF6FGVoG2IIEuA9oP4Mhza2g+wQFivN1tvWzC36mKtFcvUR
g+vyyLrFTYIsuJ096LA9Y792ZdZBYsXB3ZZf4tpfosrMw21UCAny/kfM4KqlruG9
XhjJ8lIffeiOpd1RF3E4A6hG0U0HewxaR9oBewMm1ucLRKwEsmvQo1VKePza0UEz
SdCn8H1p9fSykPZfFI/vr7gvTFy0kvx1bkw3dCa3IwRJwvGi4hXJ9TnXnP747cCW
IdynTSMjL/4R6W959XUFUOdjM5NNhhEFfuqVJ7Z7D0a0YxNaGtQRfGIXYEc0rEDb
xAdlntv8/GhKlophBnNlqaV81nWbs4PvSrRAp2V9VyBoJ77K6EtJK9+csWakmhg6
YmlA1f2lFOxY4AsujLQWc7aly7DGzJPibR4wgu1txRGT4D4dbUBr0iKpvpEJnTfg
q/or+QvaVLY7Az/yJU3T+PxrEueGj2mPRt/Mc2Ut0/3ChQR2UH9msdGmwqePh4jP
OvR2AUu9DaccDoh+jAkAHNRL314OGkw/pZKUhdHNrZmaq1gwAgpKAFBn8GuUnsFw
/IwpgVCY6XOYxVToDizFaTY+P+sCRzWxsJ8i0OPhxsrAfht4+osHHIiHeCUavHfE
Z39S9ujDKnyIVugGHHyhAaVevcwbMfmkD9OC2HbOun5uA2yAn9GVpLOfWMVv9OWn
+UgUA4CWWihqbmdgm003Am7P3KAxKy70F3yWfxPyIDF+lIfk3dMestVv+wfkRBL0
6gW2Z9lFXCwK+g69rExeEwh6JgXRKmbByT4AplEu+voE8j7GN3s5P47GbBqjVXo2
2a0npYG9FyciWFRW+iFXEgigqyUxQtQWpeE7dV2lcnjwfmIZV3H0RcozquwuaXxY
SU+69LT4eumyN3HpZaEyEmJYHkRgHOljK12e3STfmcqsQr2iI03BH63HpqMLnYTJ
lgtedF2K3048WH1XYyvylcXxCl93jPFcASSaW16V2PlLcLjzqOZaelenEgg+C/+D
jBkhYPt2P6Vv2z9WfEHmVSx7E4tLHnzg1RwlLoyHDtmj6BG3mi/hvc3gur9gESzW
S2Lb1GncO53YhkRANEob+GtGl9/5g3DnSissSGrW1CKSglA0FERRzLT+InSE6ta/
QVjyA5GqxRTkxTh28fyBZhyxu7PoDzMpj8oDsMvtOfdGoEe6lIcgkncDlrGo9Agu
BjKia7VmmCPlDrxdDr8Df/jdeQzBVLbgXHGde/wlH6NIYl6PT7jANzRtfd+pWSDy
U+3fjOHms8zCyLk8PImsuJZIWJ3ZKx36LheTLON2gi+MYOURJStvN2f/dHZGPz9T
RkuYv31oRFYvQxRrs+z3OHPMD2CmzlgHn5XcpjY1kLf/r4HksjCb7FvRAiyx5Kyf
aDCg4G5vxCssTuBFzLpBlvsNiW7D2YZmok7+vEWDHyDwXsmr3ojHui6XJS3S6UfU
2nW2YZQcXREzM29R6tXdEwUKFNRutTxdpi5BRcwLXe+dUNXdMS1eDB1nHt5/NBcy
AY9meRHTApA02U4+XzCJTvIMrq/MpBeK+Y+okkVEle4I5NiolGHNJQyJEy+280zh
X6eJ91DtJOyMMHDekZGe/FhiFM8ogVz677iohPB8uFnK6/IUi/Z8y3UiMuCxskRb
SY4QbORuqKU3z8ZR9rm68f3M1/VIR24PgNUg0g42JyHTMLWBSInN8xdSP5y+aJHw
uAzFjK8qlqJVpOPK+vluSoi9UVgXrvD03xYVXaoV9/wzNHdGnc/6VbmwjudiDLeZ
P6f3+SzCm5uA/4uQDF8hdaHGVRpSAKq9LZnoF4EeGl7Ko9dw878eULfM9Dq00x+q
Qj1kr/ZpvnnzPIESS5+whIi8zowGiyz5sne9X1o0XeC+2vk8zx+zF41wj6mln0h1
lriQfIA3r0/QNyAAesKFhp7CF+WZ+NugIIjJecuYyFmNFR+xf8jdI0AfZBCuCTKU
yHr2NHZKqMaHb/uKOvao4S/MBGsxJ5/mD5M2y5ms/TKlJteCtIAgTmekoe8RtmZv
9SzUGj2RHWtxuGLdsWxaoZm3q4pJOqF8tUp3coO8IcNl7cwGArvmfNjPIc0Ut/ej
DZxDk3Q7b3NWzWspAkQIqFjaBLXje5BHY+2VX2AfOABUkoGqcK2Gp0Kkj7XXKYqO
RqoyIyEOe4afeQRFx3sQfudVagzr5fXpT5bTAC52yNEehJoQEmqI0ej0oSMZ3H2d
XJbmNfxcaGWtfJZxFQQFaNOVhmd383TEjBTJGLIAcuUNqjYwBpAR1/YH7/Um1gP2
foayMKewk0L4xk8qI5Rgr07Oc9AIMu5il4LljFKr3l3ucqxTm+Olph3rj3hKL45e
bH5iXJJZlLza5oS5UDQLVJpBocDiTM1G1cLtM57wtumB2RUME4dsU1WAHvm6pmMg
fmfHdRj7bFz9W9mKQJUJ31bushc/m0L7tzyv3X3i9LeSW71uv/iGiuzvixhM2dtE
3qzgQCYejGg9apmHQNVEuZo+CGBjj+D5FBhFpGIMEJKdfVXrq6PF9WabQ5DzuctQ
XsaYNN9tbHy0I7mXKhpBurQ2fAupfxUpvtOyndMPfy+hkT0dnmfsOhlWV4n2We93
jGjkbRfOgPhpDP4Mi35Wh9FBggpWQW59+arvEL40I36pII9Vk3I80S7KuwPIscr2
qqL4YegiH5pr4qw48UpPfJPsqn3mp9sSppsFYsxrkPrnmuCCtmW9y6j4/LTpCWgr
VLDxv20R56I7g/dplARhS/EAb4GRvaK0IuXE6mScLN5DUNON09hP19xBgnwxn2i2
5ezX0ydRz/aialbJRrHe74w7kC3LkMsxWYKHdzlT9GNLln/TUnMb9BatBByq8XoK
rgYHlAiNRZXytinURFaE2NEGpO44aQ/wGtFTJHEXMJFzNzMNpR2chOKFOGFz1rCN
C3bumZpWvwFVUerfdSfXQ5WAKhbEU7ZwstaEVxVNO3cZfV+tSdXuBe4/UuqZ1qQj
hQ7X9TF8SVRomSFKh59BO4/KeJk5jzLVIAKNyDT6hl7Tv7IgEf8lhHHRU4TS6n0r
CmflQLzyMbC+NUuqncDDxG79/jWkoL9ugs2wcd6BaK9VnC4LpXCsg4zoHKtUhIqe
6y9CEmEXnIYhRwAykJc5F2v8rH5Ugb0sRNDxLVvwh168SVIZOtREL35TwH+Cmle9
M+Ej8FEMtwjX9L5xZZ1pf4hahGOeD/8Dd0V9GSArLQFiv0DcsUIavo7jOzI47VsM
ccGAw//FlVqlicjChNgcU7jH2PPkQnBnzbMfqFKWCuvGK0MF8P6k7IRVxJ1MT2dK
vCsPCVIJ45YXStPxlboS/eVUHas8o/MPgPPqjzRSZv+mEIlk66FwZg4yVLdytKga
/B2qgo3+aQOUSIre3GllHCj0jKPFHPPmWHKZ74Xy33kYZw+flYC7KFjOOAFZUSuR
uMRcGzZqFTtiqgcT1lQt4xT+Ac3EvCDBNKN5EnI53fpF3qKP5FtsqXaWxuwm0jNM
ZMcOX9zRhmeBcxLM5emhrkURCK5UW6Z+vBltYsl3qNdvckyOBhvyChrJfnDnCJYt
bkRCR6HLEmTUxQQ5zmER5diiLxdlq6dgCnAUkM0wJroX8gtViZPosQD4Al8qVzyw
YWpP/OCqOqrm+/gJCU6dssElpxJWea4g2VrEnZWrKSpCsbuvBTsqfM+BiS2BYeGU
rENIPwi58ezd/FYeJCI2K7Af58LJ8v1lfW604djF5TxKsqCNSBHgRCkN9bYvJXQX
CB+GF3QSOynMrz6fVnhlniZp3wN0kN7fO1bcQCOYjWaWts5nl/DO3Vcm3NyySRt1
CKnVg3x143CVXLhO10HfFWToAU+h9NFdC25ELYlIRW4cz6A1RLEm2jO7DqLOuRxc
0ezRFueoa2jhW7KvmDRl8ZbdXaEQsvtGyYIGI0jP7DnHGZQJF7SO9CoLpXCne0kd
jlHyApV52wYvXAfEWSV9zrLFcP2US5dLjaDHz9Z6TfG5sTS/mPjsXay3D4iOzmDf
SQRIMhfhV2elMRM84Cd2+Ps2Oyi3I2paQUPw5ds2upWtkpONW9B5QjGlAZ0aem+e
zuAcy8YFgdmvNx3laXglTh9uO3t2M81uZpOiy5A0U4B25DrHFVpRKzPi+eNv8xxT
3V3GslosgUbWdVfmajkTdPVHK0OfSFiSW/SZ7vHTrjzC7dr/SNMgbeaeBB6J+CNw
LHMooru1uEDc4Fnr4iRQAit/FA7uw4qH4GyyLjx9tUmFMhhH28EgQFyiu0Zk2bYL
Kprn466o6aqeHJ1IbMHvaf83d8O6J4ESdE/l5jBASmiE0NLaj7//HOeEZz6lT1Pj
kXZwPuzQCDojlkaD5/YyS7q6y8p2O5iigTgYG01owGgI53ty3NuwuQ8xgEPK4tMf
mTzicAnuTgQ4b6a1eNK9rQqjaj3S7wy0gwq68kdKS8mhte7FpDWWVSrHBXiLYDnG
cxlei2c3t2AF3yi0sFixFh1bJ1pf7bEkeHxmVgSDwQS1eIiz4urJxvLYrjD/mOn6
erQMwCVM4KOuMO+acJqnULJihvTso2smSnbelz3NJ4sgawClW/KbR+i75rwKp8Xp
CVkS7YRrMDKLuLixFXNkafjTL7wZ2fpUM4/cKuROVbNniUpWl0m7UNNlNLSQmvt+
hN4DWFSCuysT9arqS4KnYBq0J75je+CMBXatucFUfKUigoIebxTBYiQruKWNOUoZ
cQ9H6/I/A1HYghO6oNa+9aZ9NHfljwjuHJXOGTPq92Z0h7Sao17DmzdTIVVjlTIZ
8UQ6PkcnuarGoM9zGWHv4rZ9bBbgc63njIWxPNLVTtNiCezHONd8N2jwP+4YNgmJ
V6jPLQZCFDltT01HUhG0MaA9MhyjTBCmeVf2uoHd3cR5RB0ebiYKcsUT01gtyGDB
AcBvcLrVvVbQOWmDzYreHywMAgZSACm44XUNg5ZEhbJ0Jw4kRWUxhJSxe1ZrLpBx
PhxzmYEhHvOe7XacKj2y3ebdzHo/9aO6TmUXoSMcjfr2YDwmpUJzf8pz5VU0JHIo
D4/JoBQIiFGO+vUnyn6C6LSPdhgKKCDLZEEYGA+BLdOEBdOnj1fJrkFCPKAX7JXV
BLBcxzvYEnTV8NQlpcE+BMXcIYbVmjWJIB+wD7Ar3XR5abICHesFWPApwA3B/zLh
JL2Z7OZbnQePUK+XMnoTiA/Vnw9cNxrLV9sZIwVZ0uc6DIjpvRqW1jZ5RiRgXfuv
JqgaSSOmc6XC1azg2rUTnRnukI4mGwoeo9u5D7XOdSrAmZLYymuMEsOW+Tupqthy
Eo7cu5JO7M3AO51c1PLflvLyAsByIvisp/hnj6+3njIUTyD7TIZscyDJC//5taLY
rTjGTtHuMkZ0Y5B3I/LyjAdBWD5wuxsocj43PTNARWE/SKSwjcclbqPs6DUoWGjj
YIk7yeLBrUvbhO45nx513xcVBXQ18cUOSZf5zbb20F80Ofur0Qh6ei55y2nlT0tj
V4JqPkF8UaTUayLhmNhvsTh4MuBJkOzI5Ih8IYkxlKOxqA/RJq0Rq+8TmlaHRH2d
b8YCVUF361u9kijSo+2uTE6PIBtoKBy+MQywCBiLpgREhjnSbq1LwgX1IYtM/spT
pzKFloVbzdAoDwt3H8MHtWuTze0u2zjij8N3llsJX/0V1FVf7iHH0sIUpi+/W2Pc
bt9UBEgOSE6CVWJOUcHfYMjX9i2Xd2YlHlPHlCxC3FdOf10jPAqsFmm3pXbpdIuw
wapHjqUXAEYQO0xyzSsrq5H1aLnPrUswvUh0mdbGY+RjuNs1H6CgHykN0Ip0TrXh
ktYkr8z1ZyUVNkDxYFnrs5lzO012F2j7o7XKXvxVF3XKoTvcvif64NsRiR/EQutE
ILKmt62eJqAQIwonKxXvzZoSKTGJvAqgp4OuLqnZcSGaBbmD/ocaFekBOJ/fmxho
pDsprTVhmhPvsoWVFrhocF9zSHcLA5KIVGA9WZZSHD2AmAqRQQf6gn1K4SEk9ROZ
+A1nBjVJ4C3wxCRD5mfIIeHVJzv56oJGxWlyDRtwpy8THLNiCsDME1eBKUvmnpkz
qvS+dKsUD+vb/4iCVsJzOTxh1zHXKuM4a3IQ2JMvbtNomPrLJf4rUJtUK4wMEPGf
5JG/AL1IL6+KaUbltUqKQvqH8Cfi0vyoO7idel+5QFJLyoqrZYThajaS7ZbBMxa1
xe0aihSCq+kO7iC697UHTGfRfgQ7lbRdXcrUpw9/9arQMvyylWjtX2CGdN5cbJn9
n3KAinPhEY4kkDj7q++sKVGhy3/SglUMDSRy8e8DxlfsFz0XUN8uhFS72KXD2IMq
Q1oq1ri54DqJMqAfHT427Pp2hm0Y2C28f0VoOocJfuDKKcpvq+JTFL0MaujRO+0E
VWQby05krK+HDjH6xLDkIeh1y+LycZouB5sk2rqXgfSIfhhjCT0eSkaLrRAAu28e
byjjSeTWXmN4yjL2/Ujnsf3ZJ83o/BhQ0XlH0vm6yXsC9r4S4qBWeMk+/clxUIAT
lLdhbPukzszbwmzvuSAN1tp2EXyJJIsJdPlMspGFrvn4xcN6HPr7umi98xp3NW/R
JqxWUtpkOEaHBsUHHiJ+wiD4UMdkx3m6XmLzdfGh2h8jdhc5aH7EDk57ay3k7SOx
84BGm9IlK3qEAqE243IQDDKbnDNuuw1BdJOL2a0oHVEd6DxSEp9hj/yGJRKnDVey
w9IKQGVDM2wN6/H5XgTOWGGacr8F6r8eDv+wUp0QBo2JtpPYLJ/HMZIGJZCIQ/yh
xV/WcLH1qkxHgM7adx9UVqjJI28w9CIwRQsVXaJgh9ZzbNUcA+c88A1UkR3I1m4f
geI/cwp/b3wPsFsxOhrFCp0ekTRJmAfH3MgmtWhpZEM3PunYyM0SBibZA17sAV0E
VyZcQlupD05u9yhrrdPtG2e0X97Wu42A45hpPK1O3CAGEfqrCwPaty3r4TCyHGCH
Ny9SdgOVf3Eb6pImi5CjVy1r7naFirhbrmie6KQG4t+I2oW3oEmN+/Qt79cFYOmS
M69fUCwstqJMTV+Nc9FKe5AnQRql32KJKsAXsi90PHUJbb5h3CTARndyG0EVseYN
jRkm+PNtTs+C+zBWmxXNAaHwXnEFf6WMmQ33CdYPFd7WNGs+5q8VinVPpCOkeH8b
oVS0X5fdmJX71Fus404wWfA2RxmWYD4YBdLONxf5zWjVo4a1AJqsX5UrGxV9u/8i
JLsxqKxCoe65Hl2gWJUwXwWbqJQVWK2/gbHKz6qLG27QaHG8Eipn0zMRMVV2yChG
ZggLbi6QE6HLG8x6VUrzIMYaC5YP3CsyFb8kuLG6wQ/ZZdEl/xHbOOf8dYzcIR8V
GqW1zUZz/kLxe36Hj041InWhTiJP6Z+8h3B5SRSDjp21M5gOVvp36F/98Wjq5xf+
3tO+vX0H2FHBCwulFgkokKPHVLe1DO6vuKY8PEaJAhodcbcf6kX6mH6TaANCEiRU
hxuXneIEHBr6Tdv+A0/Ykb/rtgsG0D0WFuN745DtK2EsaZ3zOq1L5WH2vyRvTzje
kcdqMC0MY64JAEnBWquGPMna+rjeW5lsf/efThyw4h+rvtxH1hBj6e4wLGOKfAVx
Y4TOQPRJ/NVl9h5n1Vpw5wQwkDfcdQtf3JwuJfzlR/SGA04IDsVfvEd7rGNUBYSG
Y/ZdTVXpmP0VcUM89MGe/R18qo2O8/2Z+zuYMd6UIB0MbquFFIAE+j+gHvyGk/CH
2HlP09LhXWLVwzsY3mq9sStA2TpIL3UtK/YzbmLrpTqPh6/7JSQQ7MIZnaw4iWli
o1teiOA5beFW2F6woGhbXcGp0gcq+Be3ea7QCj24VMk7hcY7ajvZa5U2TLDFsma/
6WWL1FAjtanNRmpwzTpbFsDWdRL6UK9LKaQo1Sks0jUeO4EwOWH8zDF03KU/siOW
nwv4ZOneHaHRWMTpgAYOcd+BAm1wFVajH/sAXRO8oVPGYR6LvoUyMHBs1Zxl/iRj
LoKjLUKIWZ9qlGeB/bTAxB21mfpkBLM290Kji6yKzWvYK7y8zsLUAN6uBJnmr8xp
4FhXgyonG6q1H0tci1snQQuTFVtLHH3VWeKCTugXzSR8cxMX9JN6zPnCsb5W3QqR
Dl2eNcJCaUMLoV0sE8tWxKCMOwRnF6ZvHjYq2T27DX03HYmJWTWBNvUX59eMvi0u
jCvBdEzXyPqwrys3iE5UKwNYktBB9UfQOBiLeC7re9T3a1R6EdfvnLOSjcwvNZI1
HagI9Cy67djc1/GFrJ1lx15AL8n8GYzIPQ4z2mvYjXozK3X3BXLVQfVDcm2HTkz1
nG1sSMmUj07oYkBigS5WbGuMh7u/rI0Po6ioFcjEkQhiOe5cpjMpBukHdEJWonrw
gFan87dDvr9t+UUOaRR9cu9Bum6MBDlGI0uxI7/PnVK3IOvHpPAH2lmA01Rnsl2Q
4Hxns0z3CxjeY8qsYuHQlmqz8UFeGCa5P2koRpHQzxCmyoribnT56QY3HCRiW3cR
d/d2djicf/XE5aokliNPHOWzJK7yYhMpm0Gd0MMs7+1MEJvLzgy6dnt98/kldgrW
aw7JJ+IFADGGnNba9Kn2fduuVWy6oy6ObyGol7uRMjo9IaaVyfmTk15WbHP6ova6
g1HiXnzFWajGuws/INKs3mHPB87DyrQAW5XvqnV0lA3jC10Eh7dvWvjPq/HIp9O3
cIyJOt7VovyplrrcpVQY0PtEbUmHwYoPHnOn779o40ZlcnYzKoh5GD6uHY+Wq3vO
9LHNeE9MvFPgfSBp1Cyv8yfcrJkC+aFnk/Db+ZCt9IpA+Ei9MrVFnMtY4/+P6/cW
0KDTTHnfy5W4uFYFntn4E5zjwJ3z9CBdXXNQ60Gm8jMh5S8g4QgG3YuEZE9oMGAl
YoVZtxKNl0coCoGfIjquzGhvjKVSvvTV38nd4l3IGlSZK9ASgijoAJqZ9mDl2Pmk
+UU1nojSwrvb8Ym7jao0lAP1fB3K5gyePkZtquydHhCu/YfZDGdGELfPpSWUugD1
mfEGXJVSh4MecEJWjwn6sIgKVHsVSsfMl/VCgSE4owp5LPAkFSBDLmTTmP5DBoiT
LNkhZB2mD1ALLKCfrnObffeGPRHc1WkJou0jzzSMPInJe5s51k0ImKwlofvH3YgM
sgpv2L16OW3tCkQSsxn/RZ8a57V9SXagTtg7FRLpoaNWW1lDadoCcFS9x28p164v
xGEuoFlMoJlQaLCzMOdMFU1OHXBFRZ/Vg/PxgS8F5pyHXqjV67uj7qGdtT8Cjjc9
VDi0AXCWnnR85gkL39HuRMGFmdW8ojehjVKFD1jixfCfJZ2RwVOWp/fmQPrzh1Nn
Wy2edVOdm0JNCJlb8Fm0Dz8eYYvP5BLEd9bl7A2cnaar8v0ohjmRI14fsmjHc+hX
UtOuT5686i7GDJVutHpLTf1H4IMw8mOLbXImMkSiahlbaQ9u8o6qd43EETjzQ0+9
oUbMPWCldHayYpAHTz4Rv2v466rxA33ZMh7gKb0lxyHK7L5tpyxPwqoN5r/tcxEo
tmQuNQdQzDSW4+v6rXNqcCQjbev6NXXt9jBBePIRfbHpWVe2KgiZDQPnY3lnsdB/
XTGhawzhvUy+DFmHy457EUYUkgnApk+WWYpK9Ovx0KEfVPzb6gVAF1pu2NIY8VfY
72QT+Lg0KTnk20Fg0ZQcLOlSLjl6K6nIDz19rQ34OeywE9OV/rGmFk/obUY5kpOJ
AIaqdD6vA7NvG1xpQAPC3ZXVHTWzxM8hP6IL/+bdMsrlknGg7AokLe+uMvTX6WRR
+fvV9/hJGXLqn0+GXKedPjQKkPmVWuuMynW7HHxvaDggj1Zx8LNWdkKaK3pqKDI7
2Wv1gNdL3Z9+AMGXaXbh71MChTv8yxCv6bauPXtRWscqvKXjWr+6gEK9uOccKvvb
C17uLfRDCOC/yL6lZAW2thgNeEMgSX4Haar9MjDM/ngU6DprWOyAWpWY4rfuaV40
VRab1rb4Up/FEjPYUvUCZrRpp0+wRaeBfG6VQGHYtfWzqpBPAl6fLQtrwqZIGK/s
c6KdltjWd6oprxEgKCa5nqk5FLtbmivmut9EjaKTjDquuqNus1qHzpr0TwzB5edx
cD1I+2/xjcYvzMAyluc12cmIFWmuPskHzwh/xz0UApXtN/kANLHzUwbgv9ycSMbc
g+WeuD+kQOF/aA7Yj/P7HJwdr9F0db/HBB4iGfoqZvZdGIpmZ9OyNpLPj1ZuZ4f+
Tm+jbAcIVIMLCoYz8UdDuU/8m1cca3KzHhM1j/kMddkcBdPGVeN4RmFkPniAKf7g
5Eh005MOq98crST/F9j2ulNgj9ukPB0BYMQcFXgnwtJIc4qzczzkrUGKnW1k/SbG
BTQb2A6RttamyFG4rDx72zjMTZ8mW/8CI2kmBQWKu5kmtAo/ALY5xzvLD2tSRx/7
FiEVILZT8xidDJ1fCbkKILPnKRrKXyPe85jr0h3eRa5hjZkYrcdQeHxuLMAh6Yoh
/jvOMcSBw9bUzone6X+8qdWaER5ZZ10z4FTYZiUbY75Cx/Edr3E41fZg8yabDI07
KfBAu5fCJubtkFdGSRxpgqY50/p2YivdqUHhGEQSUH+BHngs7gN4ZZjm8cB05PQ2
Mfd2tIgbclf9gF8Z7UnyVzbZxKHNSYjz5QEV+R6bKAUh3pMZFvl75yl8GwdoH+vf
Zz8dbRrSUHzh8S7BzO4AfnSIX3HDmZR5UA5hHT/9HsrqKggQcSG/6pzmk76bUKto
4NMMnCIo5Y3te7a+H75x000sH15a82SOcSbT/xmcXLtiGdbztEXUwS7J8pyfUiCn
WzEOlV9NE3IU3gGxhDDXIvCSWS95qUMWqLVXsznF5YoNZAwSMvXxELYoToqEWr5H
zNFq64puBa/5OYmn/aAb8Y/Jyb51pbN4ibsY/ADiN3sfleZYdq79VCJll5PQjqpC
B+TOh2W33TXqlAlucKAX9jUGDh/dRS3otSsAzibS7Xw6FSWOsgS3an6Or6JN87Xg
19Pbx/VHVSo6NumTNnz7MfKOEvL4kPNMmhQx/ToZoaRex+/SktaXSXT/W619D2Ru
FmD65W112op1goD3jy/ZGkTw4d/LH9Wlvgf4gAhnc9Nmto/XWbDI5bM9KJ+MS/n9
b1vzTXn7SbcW6v/u10vmQg8h16Anjuvb2v7HZxC45KELNEn65w8SPnDMFvNnnr8X
qVxieoRYPg4iQXT+JFtqrbBPs+I7PguGKZQ5awjDr9LTCH8ADl+V+riQAVncrNYp
VKtOWJwgl42WCpsI3KPU2BAOHf2bqr8fKvEDLrmHwNCnS6yxhuH4YyKPZnTago21
Uysdp1Oo4rD+MlqhZ6qC4XJ9KgjiV1L8Hkhpy5QOAZtWGjo2Y2lHJQRV+zEzn1Ra
2Qu1Z9twYdG1G2ny+3da3nYAd/8zbodVG0JPQ5W53lozwjYZ0z5Pvx/lZuDqrGZ2
GItTJvY5cSh8RRWDpqEt7EWil935MIDOkryf5EfkrTxdBYP5xFuhLgSAtCB3o5ml
sSMElLUgGRfBKtgZeJ/zbDME/33zlwjx7lY/LPkAMR0hSvL1JMbahb3KiujWFZs2
W8xuHMPo1YIrM4GXS/GEDbD5dh6kGgvvzs1GHCCM4Wb3J5aXsQboZ1q0umHgPqLf
dPElfzXRXqKcnFY2b3YKPHVAwcwBreHYAm2F5GevnKWEA/0Q8F2HeU0rUmD+HZ99
R3HieqVteHjqczWq1Wwd9qPQf2vtH7yoHbgorbyDhbWcGdGejKzLdGVeisfzzk7G
lDNl9yabriROBlwCHdAvkC5NsEXpLKnLBbKBn35zPMY/6ZHHG6ExBt9QngtHLowr
LuaoC2CyJd2JqKHm6AnXDU/BC/+3DxT1tzmLcsx7vW3roZaperfzt779Z9GnQfpm
bGLwiG2QBxRuxU9txWvZqB67uDVmOakRX+tCGMHXHP04KlRBPqqJb43+LE8Fb7bB
NOOsQMNni+zu/NXfxPz/ozb0WrbQCJkmTTwusPPEIkTz1BVFwg0PkyZZ+mznvn2M
nabYZ/UNsKm97AixyfiGXZwBtPvHeBlMqScR1Hsh1xseWo5/NFTdpdlAnAZeXV5D
ODQ4Dl541hdzcqVwMhYsqWix7K3GFmC8RA48CDzXpozDQcFR8WpsezQiqUf9PS2Z
vG/fYRG2XPYlJv6uohzUQJPftNpEtdXbzmrraFWkX6DTVbgfl0VJ1VQxZBcG51Dg
9nQ+lHhS1ytPy9tDPTUKceY7pa2x6jeXEjuWmgZMyCX3GOpV6KcgZO9arChPZZn9
Fc5TFCyLrShCwajtMhaw+PQOd8mlAyaB/rbotEpLJD1C9YEDe4qVdHI0IFXF+W/h
9xMD88gXuMjbsgT7uMYTJJoNA/0oIUJb80oTei67IPp2vboXEwlBJT37VyxSFdmB
ORJloBYrcev2fSAs7G930nniM9KdMrh3VB+Hevgj22CUY8G9wHie3wAipLLbDWDX
GSWG+6TITcaQP+dfppgISGnlig1B/W1dUnFCzZfBdkBe8iEQxfLK2BwKp258kN2G
8Py7pqifFSxL2ddyFIFu39NAiNs8nDcjMphiU+z5YZ4ReXCQkGxgTnZ0ijCedZmE
BF1j6krhIC0db0R1tZ7TkmPMsXLaix2ACyhm87cOEWoDra5tsjlOIps2XteXIkAR
Gh+5/Slb4u4CAihRf0EnSnn4CBcYDUC/xUqlCuHuVD7FJiCAgB4xMdZivDrARkbH
TJg5s0VvYd8s9YzOwW6FZA6mtiEp5Sqji/AVL574mb7iRoIanMZoNumIWvc1+Zyz
F1naJ3S/XlgMAX+RB2AvTxZ6a/4HSJyH4sx4yNB7Iba7mH6cf0K1ezr3lcwXiux9
3Nh5i9LrNbIMBLooKYnkJgrBZu9Sux0YgE8wgmOLnccX8erAQ38CTgZHzLC9qtWT
b9LCis7kp+bd/F6RktT8xiwxeFRw0nIlHPYu7TN0E2/c0/AAeO8bjw0d3sy7xE6I
cjNKuT9FBUCcY3pl2Ok8fkmqpq4xhsduLrOHKslSdp0sffZF+fsViZqKJcRWmboj
5Cc6uzpG6BmEMRxwhXpT+LStedUGYN3iUXgLB5Crmxp62BkWpB30F4aAuT712sBb
VXbq/6TLUnQXINSuehQp0yrlXp0T+wyaFiaB+/aa6WnMvn7l2x+6WpmZhWo4lGr7
RbkGYeMDi7vJyac4lc/8+Ko452KngmTFVhAxJlhSfB4cXMhyxn6fpKcECGbJ8mad
A1BGMbOewufs/XZj65GQuM40K4M8XDdolwyb29tlyAFSCwZbW1mxoetvvHJGVYG7
fW5D1bTje5HfqueEwyeEw1qJoDvkBToGvxwAPEw8o9hwhA6bbY2XV720FNn8rFqJ
sB5tAf9Z775PBtt5MtWaiXI29dIfns8m1g8nG/36dqgWB1G50ODlx4JFVHWCq+YJ
JLLNvj1gjbcqM+Aw31xXmF5dSXcYNGJ7zUh2z7JYrDwzug5GWMekx+hA0F+EdHu4
2H5b+yJ5B0aGJBR60J1PqHQXuCu4wGlQXZp3mLZatJV7h9EnLuRBtCUc8pEy1VEX
txt6txVr2lXt9eaxBv0wRuo0Rxx21qJ9x1oqYKVpUW3Y/IQ4BnRG3TzzRP20PEv9
YdSTfz5955tyPC0ZU2SCcDyqK8HjCQ+bTMIzadYH/O9U+I19/ryHTU7ElfuFUntW
HeVgrfKYud4VOC3UCvz4HXagMEaqRw+Q0ypcwZfWPD32Mo1v3rzBJui0OxUfWnCT
qHc/sXnl6XHfmduKbYWxUuBEFl/x+vdwg8Nv2a5fIfjNLlYshB2gOcbcgFdCJa78
LSVmUgGvYDtVKH/YP+n7AjUZiXIZIVhjSWBkdXZMm9GrkqDO/gsAf5RbYl6v72J7
qxdeHhanTHtflXzsgqLb7gV0EcoTzcZ209ftUheKloDITuwFyU6pic52RiMu/j4j
KCS3VD+uECvBalbiBB64T6MMwm1OLCy+nighM3DWg9VmiH6X9fXEtrZuKJj3Ik3y
xVUGk2cd6+J2E7g4DQx8eAuRu5qOycYrAPEDNuB8moc+/yg+YVhjZMjR4UX6qyC0
NiGSwMfAVYBcx0yNuzpR4DAdM0SBQgWMWO9NRRkfOvGhFM4Z/oRW7DIIz5kL7E4V
JD/+Z6eWVTZp7K8eWD8fmYp/Jl8AhQJwRIhGuOloyt6Dcm64/6ZC7ItiVdth7SY9
oY5HO1AbIMPCok0gIVmf35p6LX6blWuq/9WPpK890QCJITiDP/Pz2p4S+4NngAOI
Sk0qtH22CTynGqrYVaZVOJidVFJltwPfsKt2ddibKfpEYWs9FJ0xjuxziVwdFt58
ISiFVdB3LldxKGQhZ/Ltjg4oG3hVj1H7FZti7pnqQJ5gi9z/g4/UqdjIG4GY3mL8
eQX98e73rjH+m0jssU9Rk8UUy/i+R8zRV9K/AfgfXoskXA0MLmnzF6qDWhjmKy9l
h5UG5gXUXbKHbJnoCPmiFGQyxmIHDW1xhF1Ydh1tZg9sDxQGqz65kJOj2K5BNTl1
Flsm9jtYtjdA664LCy8slPo86SMrCBGu0OujRJ28/UHrBpAEhryu4rYP2afL7Kqe
aBWi7jMmPlBdLXfTAFWMj7bQ64PCf9l2z93fVMIlw3ycXQ/lVCwmGOarsfpB7zvh
GaSAquxCNUwcI+FKW1MA7ilcAFNhQ5gN5nA80v+VH6D+0Fv8/lGN0/mowLpFnmve
yyAWG8HileBCOfckUfdT+wRY1cyt6QSSOVFzFq+tyvIB8sgCBKs+4qz+/oEWJlRQ
M8oXbSS52hrRILpXOjg7+KvVIM3NiHS/uzljJbqUNGg8UrTJWXFGHJ0GGzQQWHxZ
1cFxR3UBaLtnsdfv1Al4I700SQnQB5UgyYN/EJ4P07UsTKalIRZZOpoucz43bVYF
RkYcmopsUtvkS0VvxKw0uzDSUpPA5guZ/QBE1XutL44pJZIqHGvkaB2fX9YF7NWy
iqvJIfU+msHhciW/kAIMJWJ9abIH3PtTPqfJ8WKf7BK+y2zaUJnMp6LizAN0B9Wr
9JcLyBwbRB0FUOoLSSK7v67JbnZ3vWptaURsbKXtlNiap+uN5FkNB9EQ7Z/jlOB+
n9wAGp5rfRzDeI7P1sMUcBMm6B9ubszX6kpIFLBIa3dQntwEFbsC4LUuUGoiGKmv
75RKjjFo5M/kKd9PwgeTX+TP0Y4v2FVJwt/vHIZ5gJcML4IVKjs4/kbaFL2xxLIw
Zi0IjQDvTJebEenqvn+Az9jmtbTZ/mCv9Q5TsVMlBTa5bCLWr4QXP1rhnc+GuPO9
bekvq40Kn/Q1xvxJrvHytIIjR2iKKH+k0tBKjtN/VFhUMdQml+TCDBOXLeGGfFi+
3b1EqAcEDzFpiPfyADtkI0KUt0mVvJiM5gHL6QGOT9PyGPmHb4WO5wXzfc6T42hc
P3zmfwi5W3MgyQjm4TJ7CBjsKfVKl6Ky5kaPcmLd4NCdVimB+pjxz3SMZvcWObdw
NjQ9+mAX6csAdBiUEiz7oDDTW6y8Ut0MZt/N2P9kvUFZyf2ydLm+CXVZKlAAlFrq
0w420LFV51fpgn0rbagBlHvr35sFe1cJuLzx5PoaYakEYPMYpUHQe7KwIObO8MNl
9CHiFPtI2GYh5qN05rpKyx5wYkungzX2ycXJ6IFccZc3gkNnVizWJs2AoBYuz+ey
wxakW1zD9+6b7Oe2LL+K9Yxxhxk93vqDta9U/D4E1reLwEqyOT1I+hsBNKKsZhAq
Hcv2MOr1vL9kUtHkn0eZS8p7HoaIs8kDpHbYWxq3R5f8+S75BxbOOetLi5way07h
Q+EH8M8iIo3TUFMAeXWYyKMo8/VvZOwn3Yq86bC2ZtJpVAZECCPJfUfUzf/YvoLq
x9loMm3tUgOWOYNbfb5lhAljv+zxYL9WmM5uanCCeLPo6OaDHZZ8ykeCxj3S1Z7Y
XyKRPWWRJs09WWWvl68r9m5OMsmfFnr18UjQeuqHaN+dlAf8aNqnU8DXBXLMaaRE
2lP7B6Z5bStOLnuBln6AEFXsNpfP40X05VeXr/rrOfQwMMkOts/4SlonlHAnSlHv
sPvyQeJ/WgCt4yIpSVgBRSkPKSg1xKc4Svs0EqYkWg2T94eVKTLt/hE8Rfw4ZGWe
J7yHtUBX9EuEk7Rlx2pnTFxCDV5KyLMk4FlSGuPjnxmXde/5W7OXf8pSxkZmL7+Z
uZTPGnCGuFF4QACJJEHCikUDUYybc+QcQljvT+Wcf07+9qxneqQTH7JyAb79mg1C
YzOykD589aWF63ZbU9ue0md5w9ZMiFJ5ECoOP6eV4n0b1LlCDsFmzk0yzhHeLQ8l
pO7Ko+1XdR4WzgdOkin8+DDK0gaclELEQdA4hPnXjwN90pczYffw15gou524c2Ds
eHHBtQIuA29eBvQHTDxRd9wI1w8vHlTFlp+8ib2eyX+iaGAT2FB64d7ZjYseyqJ/
WrgcTjhZ7ITZP5LqcR7T88fGVkYBI0qUC00CqnOMRSECjiHulAzo48AWplvrFajF
5s9gEw87+sQ5/MqhbKr3SQLWZ0RuMCJnszv+2akHwfCSaTw428aPrI+jnyfsif8x
L9DzG0FCLQAmMkgIqxejF7wZFXSuFQzTGqePLv25NPVwoWuMIJ/7jxGkcRpqHZwK
sA5q1uCCR+VmIzjpRJMknD/I8BRVHD8xakkg9/9+Ju8jYBpqBXrV2MoNql0vXc8U
CzUxPvlh/u81zE4vRigfxNM1WAoxUE6SnH8jMPyqxZFhaOHxPV5FCdmSH6W6XVEb
5iz4VluKTT6lKD1qUTgxHx8DYrl3oweXB8pjwpJbSuZ7V4en6XyFimtegzWKJg49
IrDKfC+HqpwDtAoMvNrClRKwS3iIPiMsJH9HUoBdsQKDdjZW+ORCMOWr5ut4Rha2
Qo5bBILDP9DNg1j0kfBhT7xHXg0BVUWwrOiCThIjv17nECIgfGRS9ocWFDPOUJvn
gV3aL9KEXnIRzTGxws2al0S7MPf8GXKDY0ssp+RDPprQ/7civClr4HWYcooVm4Bw
mphGlPTFWfKI2EIDDjSY9X1HbcxFTZh41qgFYp4mVmyFRTBB19aFcEwbs1zCNbF7
mSSTSV97h5z+BCPh78sGQquNjKjb5vc/y6wcY/P8WC0KRvhht2s48CYEBTtEHrOY
e70ZedNB7FslfT3u4kD+yKrKXnclJ1uUJNM3z0Qw0nJqVpbY6k9ABCYhCtwbOCxL
zvkig4I7zA8p0tLst9j4LHHhvBuLOjeB1JuduybvACh63nR/qxvFO4rxRHvSymWa
lsN5eG3ez7/hYGsv1MnRv+IpDZ72kpZPa3TGJgW7pSCQNU5dt8kVD5jbTrplM9ZZ
S9ddjhFKUADedOzuXOVILDac2M7tS6LAGEiM649+N6JgPvVpTPOpsDjroFxcRC6W
9Xtv4dFHnyKbUEUATvCoUt8y7oUzmqtSRKZhnlg5luyoKCAi5A6LTJ4GxhlC2aYn
txfjy02CFQfKk45ECsWzm6925H8XChjeA9LkBO43na5qzuxz6fw4rqCa1zvHBuim
s3H7mQUqV42j6TC6vRh7hL9dq0niVVddDmzqRI5/9/Z6EaRyrRUQPap0ogRhwfsv
JJqH88BHfdB0a04m6D6rBF23Zv7rE7IeJbv9z4/x2x3gdjCNXnCGIjondDT08d0e
DXYTp2Gz273/QwqIb2laArtiybwZd7q34fHIrekg9bLxGsLYyvEtAhAQPpjb5tx7
7Wq4AksQC+vbO5LLnpDKyI/DiU0QYFZyInXhDWIEa3Y8Q8IMDxI8t2sPbU7bn9xc
lYuUI6jL/QVf494UYHsIm0vKH9IQHaoxzoMvQxCKkuBSAkouJZAF1WMgYk1GgoLm
0Sa0C8ShvC790vsaVtu+QpDqWoWpZyZOomuw1xr3P5yR18hkH3hQFKEhYXnPkLR8
mpJKB5UFyD7yIgAeMjIGN2gWtYFXof+7RpM47VtIQs0Noi9309ZTpfUXJnVKKpTS
7SrPry755L7Z03zFdYLvHeaUOtALYrsI1EVC+PfgPh7fVj2g8CUcog9eSymNYT8n
Zb5oJAvhmwGUurGi7PvaDxOsVnK4GoeFQWQGGRLuuvgeX/vnr40deKsD20tUUnTw
WCwVUSuHSHJY102i+0tdd0upzyhpP9xsVG5kbsNt4tquHSzXhhJAfsqZkOLMPMrl
HU7SUAnxQu18mK5Fjov+fTGrLD4PXgQnd5OUgQBUSXR1Z8/3YvQYV3QLyLeo8hIW
ujWozz/qnTEY5A8X5jZEge7dxkFSsoiBlH5Lux24d7sA04tGgEyDvy1JhswK9nXO
u8AAyIsDK0oUgoKC4eiAaB2UQZN8FYOFMgGynDLJhHWrlLYOCb2Z2t2rkAT+D9Wq
EtRwqXll6Fwl7D9WmV7j4n6ox1EBzLpCjZbAKeXoGYMh0jvjDsw7Jd5gZKHa4U5Q
VezIz7aVH50A/j/hvfqEMK+PdkfECySDCWN0Y1agdfLn24Tm28/blg6VeHgfIAOP
5Q8j+HF2bBUkHHp+Ae4hdHpsly+d1H2wEohsF9i/AIy51OyJM6fP69u0+7DEKR7h
/4OJsYWgXqhb2+k+MqV8SanzCi76d9R/LxtN59nS2RW5FXViDhw/B4aGdHGBXyPk
1qpbcQSP+1zdlzfRAFFj6PFLmjgcwBZSvM7hGugblvouEcXCmS+aogOS07bsWDrm
nxKFiqtNaJT4rReeoGxu0iB8BdMqWspuzzE5kAR9xlG2LL5WRLp+kCojh+dVfyjg
DEUFd7b0r27m6pzMZL0M8es0bldj1lfbil+s9/ihrKyaukya15997vcBO3w+NQxh
x0G5fHTchChDg1d/WZbCpo4jT318NtS2BGeX6fRChY0lhjE5sBCO4ArGytxYvsqB
Jj56dH1GLFhF+9qydmBfQTfrUwJ/I2pbMbBfqzI+tkVmhOgxGnwNKOEoGqAxI5AI
XuiXuqgM/RwTFZGfhJGO8wve54E3X5Jd6ra8T80OFNO76OecUaJi2htBLNWqxvK8
7tGMos1/2BDhLqzk7kWpp5oHzIIOMbpjBxgvGMWRESz8gqyiTI+cMApkac3falKQ
PefNEIPnWmS/TTxoPbaO7ML4T8n8nV4coRwPlP1xYdWecqWi7Jx4getUf367q5Lx
P9nYjxldIn5wnF21E2N7vl/nVB+yW23xa/pXO/ns2YP14OPtOMHOXwPG6I7yY4Gl
30iZlhzfmOCpNwd5jota9NvN7a018yrOzhy45MJGXpSmPz+ipi5UIH1T4bSO2omf
KR+QDtfjxiyb5A0U9o3BrESHY0iW6ruYC5WdtXcmLflCW6/HP9TF67Xg5iNfDvfs
v1rxzMgh1vn9X+1owUO6K1b0rnVIGcSjh60lwAWJ/ZK6dyNFNcSS9A9h0gPZVmDV
doNss2u9qa3uz2YQ6Ng3KPE3FYb9SJfN4sXAbHS8drESq9buxC2iOmBKXiNdrT/5
qtpxNoEcYb1cEb6iVbcp5IJTtHS1cj3MwdEZ6g/bB2igAVhRBGqkxM96f3jtMS59
fLdkvy2QKit5cq8nnpCRSPmhpwsZfSi0EkbGg8ES3OeYsGGe1eqHLuqqAYtsX5CP
lcFUqsKjZXhNUCaozMyXLGEP6HhZFQcrPRAiUMdfeM3LBQxMANcY4mtPVMOoiATn
lctPtJyL1FX/O6Ss6nDJjmZY7Oh1WMx2C6OWWn9YAhSaFE+b+3jFIb1iQbBBGNNZ
kxKr6yHxXr+/HvD0ERfMGEEgUWyUiXlLANEUr+uMMwkpzYNoVadapmumsIX+FgRI
CKe0h7/8WnKuVbSivEWC+d4KXoiTmywcESv2D2emRUo44FGofIDK4XeUwqal7EMK
cc47hBBKHpN+qfBXfPoCCZP64RUf3j0+6n02qzRaEzaaVgA95bn6h8d1KAaPo5TK
4nwCGPxpdFmV+OskfRDYejSwQXBtpXdcJ7zTxTsdlLMI4DYyn8+s0NUZrpwt/Gcy
qn5lxtVHFXgDkyUI1OvKqdXq0fltIF4/+te/7HkO4Q3niAivXjK9Z5HxQb6NXRzP
c7OyqV26XDQCv/G2lVf0uplPMwUVY8uaQe0PuKkKWcb9xEY3aRGQyVl8EBCRzTW1
pGqFZC+J+t7mGoHGdsH93zT8Bpq9A8C5l8w/nIRPKfXgQ1DhTkbs4j0q1wWLqjsV
0K1gkM7+nw7MnajAL+VLyRdsi7MvrXXDKJMg7MdLpB9tnFrp0dlbUL6ZSxLdszWm
HlzOEkheivo8TbfbfQDhFSvHPkEp0MTwicKYYpxWaDrsqjC5heSyHUkO9xnZtAHX
Z3Y7LVBcIc/51eqXJXa5oOJZeClJIhi06mipO7BnMN0gTHxp9f6DPY8zuBIF+TGl
SQ9vM+Hc7JENossXjrOSrlN7n/hTnXs99DK29eoXpthnoY1lXYD2W/sKQT08vTkf
UdqEKciJsCYvEax8V42yjEIx4094OAbbyQdbEiA2/U7dcLU32rr5UM/w4/qxaI5D
JNyEu7PzMH4rGQNTPtm9VzTV1EzTjW741ayqeYt1HFUsc6KI4A8kz3cg566H2dqY
SEvEsmeq88FmmTdburZ5FpPQnnAccz1u9nT2U6lCFXP84YvUot9HTiLw+OEv2ZXq
nL5zFGKhMon33YJ0yvKsJTB4umiUPgk7jVvgWQbz3eLMXeuRxL7IG6hJMoJtpy9P
4qaGhmSxxHZ2/16smoQbyfMgGXgnr+iup7/jW5B5aT7+spP6TNc5YsWxQ38p0Pwe
d5SQ3zZbFGP7grEU6SDNGkHfoW7crOhKtUs4e0sydSkccWcfjOKav+/ZnO4Jpws6
X632J3ap7zIk6ht5FIdxzEeEjCG/luL+weVAqHzEaXRkbSRd5xmy5Ljz4QPX5TiK
LS2RR7IRYS8kgP9vuIBXu2+uWXu4oMh1VY66hIjp+sBrr0pQEWyNQ9TUYOr6lz5t
12RXTKXmVFIqzmWlg62cjN1AtV+mfgUMvjszgn8ikB7Tv5JRy8xzWxaZ/t5fakW6
xEOkIkYwIPJxvw31TV2twp6K+AiiUG6S+0HRHYd5R89nihtD1Ho2D0WNTGjUmKNn
pdhdeNTwtPKg8Ub8Db7SJHI0RZLNPwYpAkTv64sUpjHMjFvkfbgB7oKG/0kMOus8
o9EoHvjzXX5LdFea0nrttGlbsfZw/TP65rjrkoFskF5A6AKVfEMloHhrwaFK/QKE
n9ODLyohkfLT8M/dli3tF5qCLD89ZQc6ao66Q3EmatgC46rM7lHp7JZqaOR11ui6
W1C9nKI0nEtKwuHMmbvHk744r20OcaFSwJ/605b+NNvphqBejB0htFPJPtFppEh/
JK7O1g/JJmtMPKH3gNtNCYS+dpw0pqQjazYhvfIpkK/GD1bQfCFFtylM+nXULQAM
MISxVknUaY61fhFPXnnt+SCFwNenBiD6AdsUKo3PX67rRuEwjjFA/Ta5mMa+xRKX
Yb9OZQppJGmSy9kPbF5qBjy4ZjKgnyEfiIGkUCaPN5vl4cJGTMJSqWYlo7SRM478
C+CIyr5nnps6bfcrCuubT8dEQzVL5WiAVfZITQcIhTCAB8UYl4AshDeKIcdgx3Vs
nLmAC//rgVythDDJOf5KCzY1AAPRIcEEPymXbrAF5X8zhXAHWk1K8BR9OzSj9Pzl
IyzGdr90BUen7m9Xs8IwEJ3Je7JpPVXfcFiMR6RzaqQOk4HvDP6FbYlKgCi+X6ZB
ARZ+EsyIiaPzO49PPclSRibMhi8Pzse7kSlGWL5YYqBkMR7jc0zBbwUCvslB+1pk
nMWFyHlnrlmPOJhJ1DZac9raHm3hVzg5OjmwhjjsVjTAFrG3KenU3/0jogvxzA8u
smJzRZO2stcRnm3duk/E4WCHApGOP9bz+7zH7Ug5k3CORncG/SAXF0teeNHvW/lH
YOmHEFTGV2nhknVPFfC7ErK8Eda5/tv0yfqGSLwbYhmHa+YlAeSFsRrZo+7Tzj6s
K349JjwdZinzVRaZHZlEJAJF3Mc2t2Q62s337UaUaLrGe2ZY9pdj+6GRzS8D7ewW
kz+n4dpIx1OEMnjcmPK7F+6Bg6nGwiDpcTyayVfQQp8fhi/KotBwvjLUk1Ok7q+o
mT9+16aeNpXcxREFHaELFxZcdUGF79ieo8DEMWTeiCXxbccR6fjIP37i1Gp1JkLc
Lvs+UxJ7u46Dldnn6ggd2MX1BuGH5+/12WL3ZDbxMFxEOF0pFsMQN3Q4j+SWRegQ
j08Ktfsy6lb7dO3bqt7mCFmsxPqO7NMudyOvgjCHzwdb6AJIEwBMdJ0+KEolkbUE
wHHW6D5XW/b0palCJXhELp0INVpyeIUV2KJn+hmZyvWIb9rsYvj7ptizdQ14vR/c
ClgtojZiX2tqHAg8AQUPjWTPY08wlOtzj0wMTway7OuRzcNt8fn1zWB0fV6fOgot
/ovOwa7fuGTT57VS61syxt8qjjCxSlvkNqxwfaopgFdBLHn+xD2G6CCdcpUzNtjf
3teoOxOD5xC5Z5d59UNZZu7+AZqo3ofFGTRcI0HJMt2byP2DuJsOQS5De0Z34SnC
kyDOjOBLys7yhZzhS4NqQAx+SZkF20XBzykuSX1MQzsKteoppSZ7l33IT0Z5ejSP
8qwFGLLP9ryrdI6pHydr8hEh3RQOHC+g/linoOwz9OGw55SJkuDmVEFgCpEBv3wD
D0y4giO9/Z/ezS3jPBgr7Zc3+meLu8YUjApz0oYdMYh4si2TR4WQKA0buMVOKgQH
fX9koQrCqy/+LK5lZHyefTDEjd3FamvGJYE3F5Ufht1jG5Cl6n5wLhAjSsuPRn+i
GcqvULjPyzkBkIqezRwY5r0LQBf5p9ZrFnTKxQrigDR7IDLNPUiEW9S355uua8KE
N671rACCGtPnhzoRRvHcmqyJn2pAXBkhDwf7urgeRkIgwVgQB1vqqitcx6/vB0ys
IDvtnRYFjHuWidYn+W30i6lyspR8WmSeo8JxCA/cycV4ikvPdqdvzlWj966FXj11
KZRaUdDbAfzpSslvDTjihkiZcpuatO/26/StQhvpKsoAdvolEKDzC7FJO1QtaWdK
fC+FOILXDhIShSpwbzGrepuTpezI8eJikBWTqDHPpwAM3rCAuEuBEa/R+SMiw1YF
xK1jG8OvuULvccs/L2JBUB9LMpsl3RHK0G/qFCJj1uO2bB257EvfhwIUwtbjMNqn
4iayY2V3UhnRlEULPwdSggyUw0O1jBUZju0IpCXvwqVOCzQK6hHdxdvMJRy3Doy8
CDq7QLQiuIXRkvfpOeehv7jwbfoa4B92H7cxPjYL1f5ZuzMIlJ+4plpVYtAoFdLV
KiiJJR7W5GsPa8PND0ftt/Jsqix6DsAzxzSUimvlUdEDILy5NLECLHVq8yjEgGEg
XkyVsUQC8fir3Ytj/xbC2Jy+lbILonU7HJwz0RkXr8/7xlQYuSQctc/LZip8Z78N
hBIzhchEAhkMftDnlauIxdQeh1gNvLgnTbswq2l9QzO0yeZEkNSmTYMl5EfRdLmf
hJj07J/TQE2lK/kqXs3anMFP6OqZq0P3Z4g44iP9sHVNbjo1Ub0uahRgijbU+vwR
3Zwpxp/BSksF2qL0KDpVmk6N2KurtEoM7zIB2e/Vts4AW8cPCGa7X8bWNn+knieX
fpFsRTI5HgcrxHHj8agJfAW0LkldrWbNRG43Yjvu2J0sideWmVT3J8IMmwj9QY7e
dnG42oDhCvzPUUKNVviierWUfAJgwqgyCH5jgsY5xUwa+ZJYazGEztMgoVvnpMGX
ugA1RAq78L06yJaQ3jwn+0PiMqNe04sb0FlWfcH/PDAMQ8j1iE25ngKPk9wjtaSJ
IvzCt6HylL46CvJz4DnbrprXeDvTgf9pjZPOVPyHxWz3P1JbRqmXSwIv9qIDmsMS
EODFOpia2/0L87xUmfHAfxTtrcMOoI5ieUWOLbJw29OWEUkiQJPj9MTfel+XSRIV
YAFT6H6KK+6sytc6D2dxjTtTIJ5lW0r29igf0FWRjHkbtA0XiylAWU4T0E7KtyLw
b0t8c4KD8db7Y5vTvc0NX+WIkvTtkBGk+ko2rq+7a9+nYUBaM6QgC3WGoPcREyVG
iGDQGhPkPx9r2OJ/faGl4luMS8aHqKY0+mLBXTyFHz3Drq7GhAFuYZZuHgucNKR1
EF+IFKwbAhReHNW3yUNPBWmOAsjHiN14vVSCi0nZp910BzoZckJCYpkXdzr/ipXz
57ZWUr/QMGIAcSTxazRuC4sYjGRQ/7KYl7fsWSpOUlsXsNqnCq1qLculuARckU2h
ubWTk2Vd+yDA9jXYj1hBAizT9C9UgVa9XWvYY8eDksfP9G1xP3sTS6qu0MJnyF4+
y1o6pWYOVn1B0UgLhHgaGj+WQZGkQOMb5aGtrw/S9yiLPesqdpWkx7Jh1VJLUI2z
Bzu3DWidvQItXHABOm2HwSiw/YuXRnivpJQkJlCrz4qmUHVIO/B5X92sYaTyZsEX
RxOig/Zq83VYdlIOm0cgSK2rzOa0IWuYOb+cNIOS/3KdfH82LgHmmWrklhj0Gd1A
/ac5kpYuoF6BIR0C0NGjCNPcAocbygX+L7s2TyjafYVuDlRjPLLtlKQH2PFjECNM
LV+Yw2m8nbxnLehmgzWR9mPvF+2MMD2QLCgsVZvwgNjEi9My5l0dOo6RtEFyeSz0
XY3UJmehcJmv6GLBTGCUVwFFJ75e/ZqJUxX36Ya1cOm/6C4xgvYhpCfSolBXhlmg
pljz3ELKX4CysuUhysnwTauDqX3JrHC6YhrexWlcOcLHosTN7dS0AusmCO2tTwIr
wflRbA8cesML1I48x2AYtmrSNDtUtRocAlFvwFy+PfmvGmRuXt5tVaH3v4J4qqnT
f9ZxnNp62DuSoxdK3ovW5U2lWDLsQJ8LhJvcHVIvbcJ9i6Yw6VriFfMidc3D/C0S
J3A/tK4ESpi9mgCIw2oDmrpranb1tFUlSDTJpUQGRX5Ztih/hTGoCWBXYmR1ZH7m
pxqa7vHh047L6dXr52hvpQBIS0nIuXlvnAizXzAxni6AeB7IHqUQxP5bAJGt4ya1
kTHAgr9KFqnwV5x9puAN16/J9euFLEmR4Sf4iCdgycnFcf97HBvghXlt+whps4mM
Fw8vCb/q45SLL9EcXCBYswpDfa8NsTEiKryLr9tdMnpg9R2izLSSfV+tjs49W+rO
0zxxfhEpjVZBZmMKHy3guHus20FORoxqPFGntTzvOzBH4qttQOBw1V4L9G+C/70Z
h5QzpYenF/zyG7CpD1aj+GdQ/S70COUDrM/grgvekMNzQGBFuYAw0kBov03x8F8e
/VWBRpOw2q0ROXLzdbdkIoS/8Iq6D5AExo//ZKldrjtF+y3B7SZtx+EafsdK9Dm+
4powivvdQE70V0Xz+NxrPzmb7ngeiKg5XI7MhKvybY2nNgh290NtLDzhaINoWWzA
VdGpihOu/mEy0FS9epJmLip9FD6KFPd1oTt/7r3SUxNUgfJJ4kj0+N81NbG11yPb
eBPhmotuQv88iRU9zf+9X+uT1srKd4XNdEfbgv/PEEnfh5izp3DIfj9FT553fgcr
YwjpoA4qoPGwZjr7hHXD6Q4H4iv/sETBWrX0sg4yT4zjOj7qWWjUoF8HCslPAHuz
txt0fbCBvpJMRFU51lelJZ3s7+XYbb3sXQ0c8At93KFz1UofXLRkv/OuuZYQDqpl
VQuYAmZqgpL2wobkBinxJOFBnheBHTg7SxTh1JDq0/LEJOLe0vScOYPQDgJ8mecq
ZNLIgAbc7nKqZNQZR3lYZel3UULgrVs5qKFLiBqLfRWcSOrHcpRhOhH9ZLSQaPTf
u98ejSXooHArB24Dsjd0So4CXVfQxVdj5+QFXewoLBW3ijmWHBlVSJ32o9MqOtua
Lu4f1XJq+Xpw73l19qyzjVV5vs2d7LN86FvmipxnkmAI6/depb2gAFTIKmXCKgdR
OlExJT1m4SI2Vv6Z2kSzNiLO6VFwgkL2NjnYADumo1Kl8DeR2D7D6V33LsOXvZKd
Gz7ZMrQj4W2PV9U1O8jGktFcwXtcjS7gEt2jHvOtp8oiToz2XdoiUSGT80kIhero
qlJRss1NEmYGciOskgMMKaVhtFc6W3LNf24tGPYZZ4G9IfEsUfv7tO/16bGi9duF
Mi6O28ojzyoukTU+2FLNCvPeEj9LB561wTzE4eucHU/7HGquTc0m5AyzNc99Ifna
T8K0ejMbdJo4I+vQd0dfbOfEqG1Wvj+1tVsTnVJA39bLoS/xeYxv5Yygfl/jtwLT
FMtGSwd55YoLkL7AdKuovDeceVs/qCkKgZpYOjlDFiUtnyfuJvp15LUrF5KkLAaA
qb6r6qeNJszSy/weWpmQ2d4kzFFREiokSnAdm6GuuperhQiNntjsI4sXSFAxKlFi
HwYJ6/LmphwOT5EK/asjgpa0rvi16DLEqA16yUOn6g6UivQzuG9hYfnMMcnB/fLm
oEE6gQNQJF4aU9SMI87F5Y9yLRRwacd/6Ji/FIPNTAS4mWE4BHrmrHql6JwVsv1e
V72ddLyZHQpjvI+OTVhxRDBEM9esNy7n6tbVz5jmpbq8Eokc1SaSVeRhZH/j1c0w
ozmLY2qJqNgSzoip9SslBwVHB0BxntynPHcB78lB3/+ylmIPrQ5zW0kI+YctY9gc
VID0os9WuKTjobGJ2ZJbrz6tSlMtdDhh7gwmDaYmdHRrqzckPHAwBpZU55M7+8Ez
Uxr6pOd/yRmKaVPMW3JZv3j+FPfCSNvi5BuvovvWiEAG4Wo3/ETIXIX7aF7nH8uY
bz5S432PwUpoM1bO8fn+u9Cj/uPdoVOZ4cJnPlUA6gvde+/lweKu5DigReiqGbO+
XMVHrrGZCFbrSyrEXuqSyEaxcenw4Wfe0J94eWyG80+bWfx9c/985klJ0uq9KTLq
0DHQy7c2DUAKlM0dYgIKzXL7sNA92DntWRst8M8uy0YTlvhOFHXcEN0bGe1kfdrF
85Rd/JKYpPaqW0w3Uc+fnbuvp059gx48Goq/T8w4rj6do7jcGm3GOwGVVtNlUDyH
OmUdKx3PJFzD5LNFMCCNd+fUDTK0URYp5W/n5+lsYKVlWlpe+ggYL70I65O+8+N3
KeWNfrMTlOeTwNmoMlBpMfQaNDtDks13lEvMTO+CDAx+mX9pa6shxidUcSJLYOTC
HtJ+1IL3wxV3OBcxeaBH0MJTalZ4qxEhZwEDpG77C+8cdme6ezG1gyjGI2QBNRYq
3NiZz9KEiJ1V2IIIUlm5WgpXBeTbSj/JiP/dKecDWD3BgP1JRAa45pyv8SYa1w5S
KExWa2A02PmOqf8i9gqIvGMOfQwN7W0mItfi7YO/CoF2XZLY00mFoh5vYGQXhjo6
1NcR53FWE07/psV4PVdBWrALZ/aQnS4ggwSyTakPSqVIw2MbnnG3j1NdqPUTyCU1
45hUc0jb4h4se623qE+M2qjVxY+kAPFK0oKMuC1rKPmjfOqo0JiNOCfSSfMJJT82
bqVDBomG9P/gwkz0xEZsmSuIjwRSXFsTSrZB/U8Bxs4lU3c6zqJEafvdY0Lw70z+
2lp8rbcLaVcJ4icjrR7zeG4+LGCFhRAEcauO0uCPcFtI53XgrHirFjICv2zAN401
odRzWGgCoFlS79f4HkKv4eIGiBhIGIqKGwb/i1TDzMYN/d1qSfH/wTCmLHNOwTJZ
Sa2o6d50eoO1Xj+fOlM7G/NHy6CkYuCha5wxRzDDeVwKxrvPE9iBMfpm8eBL3Trh
kqXDk33D+NfADKiEky1Rl1J9fjjwgNiNph/ZZXH53knKKrEzM03sYrvuPjOC8lbL
KJoy/3A4bnTcPpdSGAVLLqMZO4AfrKKNNy1wBEEEjOEDZ5LAcgX+hyeJjv0MgmNV
TTDk8Nqh+OZx7dXZH1yFjnpMe0Uk7cCMNnHNPkVhrx5eAoGPZgNI1L027EZw+pqI
qF6w8YUGPSQXXbsMriGmiztzyT1sB6tRJiTXsN2wU8HU+5SsJgYYGutL33XBBUt5
TzyYMf8uMgwMV8t8pBWznaiVW+G7V/2HtRSIBf2deGOPeT9h57K1NDt+0brdIYc9
aravLEwXVYcpFoibZVbz+ENYC6wKJ5IlhOb+X1c7YU8B9k4RJdxzypsqxpDK1Aki
gY3oEiA2URg2qP2gsgnaHLiy9hqzJ78BNrjGcTf+kRu0VxaDcdgMXL9c3XYYYU04
XNEyyHWqlnY2FLXo0lBW8yI44NK9KBf+6JAW/GJTTJqYVl3e5zGKdyrfyyiGAQg0
bSa/KBAwIIN+5022+9ZcCwtce+svtCY0p0TtIW3gBkKlpD8ajerZNXkdo8ipFbqH
d11QZrA0drA9lsDymxL87Exs1xzv4ByO+JpdEFQgNNWOz1l/PLwh4NbqfO0ExAg5
Rlfct/IidiGKKUy3hrZ+gvdN15Ro8jdtP2fpY7hHvdE9LfR1eAV4TQkCsoOXDqJp
j+fjrrOA37Pim3aCkMgG4KHLsgBDAMlyTWEJHlEsmUtME5QwsOOAR4A1cbBwUvMI
+3CI6eHlZXx/XX5I56z0eZMHZQ1VjOkYUkj90+DwIvK80VMFVLBljMQpQOntnY2Y
FmkJiAY1GBTuoYWgSPR1ET4CqciedgEXEPN8RlOzmi22euYBVTa5+Q6rSmMVWVgR
rCoVCZWcqRjlsn/hUQpqNvlLltRrYjyoaIqCY9Rfigb1rLukV+biNNMmRR55IU51
AKxS7QEaDBOwoy0nHa/zgvTpbE1ULVa7LboJxK/hgmfSYiGKq+MYY7cCLOVYPstJ
oReOB2K5PbiWfv45r46+l1qrQFAiHw7biBsxs0Ospo40u2iqQRAdDA0HbTBzJCJo
1DvmjwJI2BqH1MOD/kdyA0lEHjhuP7cBqnfxF82zyJ/XhYYguVs+fzZ0VRGSJqeU
Y+Y2FDpCUN8QY8onVgMxRKd+tF3wSeB9/vg+6secJJMIO5gzzB7LOE6IF/u+PWn0
tj9+diRVQdLtiGTjHFsHG1CnAKthG3KCfYK3UZqUhruzUwg2w4J3Qc2RtQ9HpzbN
lt9mI6C2JnlxPKawdS9tjWuI2+oVTa1ocrg97RVZbqcvH4CZ8UjDAiBWu2QaCB6z
pkLDuMyr139BGSZztM0gmyimsATLlNfHc/saDwEjcX7LPRQjojie0KB4i7d5kXTG
o6f1iFw/u3T2HlsSVZI0j4/ehtWcX8IWA8gMim/dqoSZEvd1n41EOhQvphLCdn7X
LnZmVRe3alSNUSFkGI+xWhiK5juusGURck5dqDnVifMouidkdrRfk0uXTi31+++c
ewS8diUVTUg2yQrDKWedQr+yJQvE8I/Sr5WGkf+qUAB5PxTviCLJnsXa8ftWJ+nr
Rg4KmfnVuUi/3OsZK5xdDPuLA+cg7jCiwRaMjRHRtegts+yo+Oyr4OtY5Z3nrt1c
C//oiYmDJ+8hnmuGhle/ko6sIUm4ToCrmS4KMYKhz7aiSvi+2+Ayt6LpJNc2udxU
sqJxLuW5f4ZdIeO8T5dnb2ebUP6tF1zVFFlReTjWROyhlpZMcCmLBikhSYuWTWda
6IWSDJI1i1VpZPISBD9WWn4FDOiuW90ror9RfG6XElfqp2ogNZXQvx24B1FbHeWr
oZ90pSq9vqPlFsFn0qXl5jybH4XyD+xDDFQGej9nJ31RTYIaglJprC1RLwWUj9+4
6DncxMQzTuUfK1fHxqfdax28YnytFPpdyGw0q4G5NkH6V018leZRuroq2AZCdwf7
+RuYM6sty7TRO4kq0mv+iiTI0A2UN0uZilTo+X2RPoafkBaN6MXnWgGKR9BVWn0v
1Vj63uWAYWc2n4jZZSSQ5pnebrfUwASCRHxrH2XAQG7jxwnIAEQplfmnzDVxTAj8
WFPGdUEM/P92FUF7z1Z2O+ZagkIA+LzZr8/GEuG+AaFVR2o+6Mlo/MYgBrLCfos3
TLslLo9sise2QrlCeFtNMmXDpMkvTOxp20mylDOuYjoJScRw6Bls7OJh8+nuBj3P
JgDngbniddXxWwPbAlbVZSBBLliPQCDkMPTf33CuWH4CCFbmku58GC92eNFdhCIQ
Eb7FWky0UQ9E2ydn+4g/llWr3a6ZBEkhdwfAD79LJIDuCqqSzB6mBo8whVhq4e3W
9rPNqAezE13iJassETg/aWHYbSjg5fBMcrY/LhmGaEyyE8rzOH4e39fAIGYs6fw7
cF9AS5t2fgb8VGgTdrCDWNZMvo4Uhw1sB9qTlCg6ePEzKzHkaFeJL/f8bDHNWzoV
9O/dXH4uSOVQlgYAGh1rXz/yDFBsytcn4X82NEqLfh6polrRabDbIobJOoiRLCKA
ducLjj8hfzMq3d70uUxXB1JMARK+F09B/UoqNMO5K0TGEcffb2dDhpdMqU0/kL9m
JZI7Vt9WUZ1dipQRcYpV5ZNvzGdz7Vlluu3dYUv05Rz/2dMm4VIzLXKeUSKQ8zZY
/UP5CDf6PGnP4ZRycu4oghOvUG2Gwm9B+nXEbOGCoLMa2PqnvjFVk9cYlqm9Bcf9
yydXv1exVRapcEHzj3ZOGRk7Evaaj+cbc8P3B8Bm2OElnSkB1sXiK0guLXWFU708
gTFoK2FGYKvTTPnuphkw3OGzvkp8qTQT8QZ8wO3FZtXZc89DrQPwCe1JOqqU/U4D
AASiwfQHcDlFV2hTtjyOBdfhrRn8el2FKcsl6MOE7U6RlFh9ZrC2gNdxvN4+aY5+
V8ZUTakY1US6mmeNmgpZytpRilU0p37ip636eRdthdn9uFSbthD+0Kmh6y0QMBSW
qjC+DRAdG3GCMqHYV+EuAOqBVsOCsQVwl3ZoQQnpeZOz6aADIqcv/VCeu/Ig0mqo
WNsHLQBelGYw7BDfCByvdb4pmYg/usc8EsVG+xQSw2+nwJqqrUDkTsJNAcIQBjQu
sMCzsi3oQdouu9CJw/se3F50qKwbFMj6zxoPtl3AWESvlIQfYQ/U/z2YOhx32xjZ
07avRjTrNwH9s6C5dopDwQwJe7tU7yA11fv++6wmq5xWblaCvxpHtGile37nl6s7
3SADxRY0hM/WoieiwwPhgWL3+vt4CGPODo+lJ6loYqg4HqolF1uY2a7BN3vJgacL
UiZJsxw96IrngrNojJVzgsxDd8g5lfUGSADFOKjCS7BvSoMTQGm3/moLrgeelIdy
xX18tQhWTt3L1mr65h6GE+eAeRDtxSqaPN7XsMw5UX4D8wbbSFC+J3gtSVzPtSUw
kwTfKRJv3vuPAoV+jzZQ/4ui8V8/1UXCyWYAQWFTdiCjxeySJhfOIQ/6cEqxVChH
C0jkEP9zJroHoTJMm+PxaF//+Im/SWa80nQpbAkRch5/LyIflINtDTsSHABUiD88
KtoLOWVtQwqJA8Kx48bWZZE1uRg7hk3RkFiL+b1XJl+Gi5OkFd4dI97V6D6PTAHW
W39dw9LVJhiSKXIcstkAadOienSUhnGO+AyUeVO/AtQ2YgDDZTisAipu6IUcnhGd
4pk5ZtwblgRwZBATaHMimT5JlcFGZZNvJlUGy7KXDnq/6+tRnij5TAjnU3rM72Kq
OvnEnJTcljIrlB5smxve0VXs9mLqTAkwCeesspEoF7WALO5LWg8KfY8PLOtndQnK
L79j0QNqOsRf6U5miS8PWXc7mB8/PVoleJzrJGkX23MLd9raVX8kdveYNcCMn0v+
Rwb4prQVuIC6dOU+yHzhGZwqHAQC1BFd4JuOlY+oaOZIYdxJtpTAsH4EDT3uWo3S
+QHM/lZHbSzJi6phF6EXoQnlb2aHDH9+7ttQ+SkK+l+kIkBOnknr7JdUxNiEmTg8
nVOIdRfbsaddnzkCVLHgU2jK8Vv86jj4c3/LAFmnnJLuCZ/AwGk4iYyzJMqJbxEB
c653HqEiSr1w9s7QZLqqgbrW7HJRdgqSXkm/Ms4HqUhjevZUqkaH+ls5X0lTknND
zNZtLi7ySA8pMw6vOi1cr/OkVSFtKEcxG+bmJ4oEOTErz7RgjNIrhBlotPZ8vYzP
u8pWs5BKcAE5U6l3uKUrNEXuAT8eO7V8LQxzuUWvTWHA3Emopv9SEv/2NzrlpgLp
2py363YYnQx39+ks0lUNhCzYp+bkY8SBi39mVk7IG2ucJJo+7YnrIzN+GkjO5CDx
Ylou41fSfuddi4uTQkKT0Mv1NBQV3e+H8CIf38VR9xZ1w8PUKSd4GH1ZSCIIf4Me
nKAo1fTKm/bVv2tryu6RAhHuY3Vqk2Ds3FbOaT889sXpwo+G8TzP+4KGq8od00ir
1xJFTfo5AmblNiEv0h3FtvAxjatTHR6Co204HANJOI6eE2qtDy0I6SKAKReruxDT
KIsvIlaPwY7VJEAWyuLhoyW5xmjgzEkSGW9buiHhydYq0OOqi1c0ediRT5+7jNZJ
VxOZUtZQjMHAEzcAENQRqFRR6YqElKOStjC0UkqIIH5wPTSCIjlcNIRBqXPkT2L2
9Qemk0lv7dybunzgpefO6aXqPG+/sxqGRKFwgIjVduwsrLeXUEmQaz5YBlkzwP0t
XknZnJN3AJbsFTCmn3Ly935RWxpzQrlK3FhiqaSa/UKELAH/QGrelehJtKtGb+x7
h7jI5YmK8JxMgnWxVnM2Qmu4TaMzNLQrzuOg0StR+wX1w4nWKSeqCwb6mmR4rTrG
9p7YTSIqEFaeKy2qH05aUgTG2RaXkOOy8s7RAwU5jL478kWx/sm7mk/5/QqICyzH
gCmjg09IfRBzxXj0Y2FPT073XJaIPL9X+3sKBy5X8kstO/Z3VKCqAH7btNQjmNVE
XxZhIDznkrKU3xAMsl5s3cowKhRNgaPkHcNJ1dfYmQ1aO52dUUfWCPDuSvlGkvFP
r1Gvb1WSTGw7wr4XBmhU7C9VyQl4yjHRjfagwzBVrC2ve32PD8YIEW/uC85aAWx2
c0IvqK6gRwzjeBvcy62xVmAX2jhZc4aID34A/efXzOLJEpyX582aaJxT1+k5tXr1
jkC1BrInfJcsxWO8j/cY6kfg7T7EChpJlGgWOdGLt3Hmxppvb2IW1pg+LDtIWxAb
hU+NqogMYOio9sY2jb+xa154eZPOVvZXRaMGTN7hfXAGvDk3F3ybz48jac8tlVui
UnI9xrNo4R1vpL4LgeStnjS2aLWBKY1jcwa+lCxNCpeE8CSkmUWIY/YNS2n1iigB
ei32ro+gPQe/h+9mVZTAxXvkcZLLgZau/Ut4XofrZ4sf9Rsu0kpDp2MG5kPNPCRf
DmPdgk5NMneUdsniTGo9A003tmM+7Ilch3sSRz/vLAKKzQVdqbfxe+Yj76CvLlkv
VGJp+yOSMTpASk8IHZj/CrrMtBcmJBoM5PWTny3T3yuYC2aX2Jkp8FVeCOn4CWKp
NHaDwdsraSQGvvkTYkyxOvdWbnF6Ti6KZWw/KFB+KPq9Mp9eG9i4oljoSKoimaY7
HoIs6dQsZvklYohs1dWiFmFutPKT2b60bKbTnULc69IVLU9tkvmeUy2wvvXjZDTc
TZ9VVG2g79OuP8MYQD9sL6jHNl7xQk1Vgw27pqkE60xvAMw+HSLH+Ac0oS6xp0cC
bALZR+m5dkRZpGIm+TmhVlizyVpfFAD6821XNvZmnCanxuQIVgYhYo0NwOL7dxEA
8+ceCp+/1IiNoUUoCO1FDT07ecYTJSo53GOnFqgOmEmBzkgVSJDJPL49Qj0QURh7
NZGl+nTjxPCWsPb+lizqij9SErgM0NKoGQcYKX7wZt8uc1S51ZVZIDFAc6nqKEUm
ZFfQrHfpIiBHeu3/zSNpicWD+VGSkTvXFmcdhjHm1HE+6lKe7IS59ih+M6pp3qpU
1N4hmg8AWDwr9KmGdKkMpJIGL3bxoeiU6fu4lYRllnFDMkVN++n3mLM2CMAP1m7h
uq4NQlvQvqM7lWxk45l7DzBOXayoJRRVpIzYQuXVYJVbGtOCkCojceuuYuhNSp0C
Qnb5r9TuVyfh4amPM+0+8q2EpugAOO1XvE4cKAuRCuvk06Rz/LY472BPqzhdnhd1
rMBqoMWMnlD0XDOXQ6Py0HVQESLoHjgmMgB7dCOWSWjUBB0x9KgQtmlq9EDQ3Y2g
CGgGzV/l2rbm5cgG2oamuhdkGz9GnM/hlSHYnK3N2kYlQR0gXnweDvQ4JkaIdXCj
SARzF6xv0Oa9TNWx8sYW55+fNpDqsypIbHp+ODqi5Wh4lAI9FQkEjNDwI3nlZ923
LAiFnAyKt2Z17KlHiKNI55sjiYzfmeO19FX4gRRQc3onhTZWa95MCYUEcBDNmVJL
nAyWKf0aDx0UqrNJDMVq2uKI+g+bjdOumLDY8KQrSIQf7O9P2MINzHU/326lQ4j7
1JoJuqG3a5Ac+onJv10rAen1o5sQuw+Lgo48WKIBPuMBBaSXjD70khujZ0p2+bmT
d5W6C0j2S7dJDe8HEDpFoCSOGdIZaYzB7Mu94fTFdLg/XOXRwPETcTY9pUDlFPN3
b8om8r6fNgsqPGwYbKpAH55c/HXk4ldBgV89s2ZMwGWXSL90hgwRKDQzUF2ApIZr
LOX1O80PwBpS5Pfo2/KD3rHqBwFVZko6CGcyzccAi2V84fCy4hFw2GuriKQdBL77
ZmzqZR3Bw5nWlXKifC6X/9u5Q2l5m4Z2BZ2ByHHYDJ328hdv2+hq5gK/0lJUwoVu
Nt8YOKVz8d0vWQlgYYuX+/o7atwJ1jddHCXxfKQtRz3C1skUy36+BHluNSszH6wl
8MWyMmSx7yzNqG5C65hVmQ9O3jmOqO2MKBT9v2RFEcTIff053VosSd5d14RGmlf7
h03SlrFvbU8jYyMu5h0abFnLG3fe9dOIRcxx2UPx6LwVw6yD8Z+nssY5JEIwlcST
uphBCGecJaQ1B/b2hhv60kAHUMjMzoqzHTo22pDF4DwQzeCTwf6TFADLz6u/Zldl
U5ay9OsAfpoko9kqaQ0N7Tw8IBUfvSocdL1I/so8dnTS4bDbZz8KAXw8YHbLcwpr
x7KZSjbOrKJnr6ihf7wmGislMBP24nCC8FEDPiKX6KrZ3l5YGNjt0XvyHdlf3x0n
qkJA0Wc9cKJm3OZRQmKJyxz9C15d8Pfa9uiRd+mmLY8REIcD+I1DSFF7I4VH5ps9
qJJcFLFMKtGoR6hloxQT6mgeUNCmIQXrPe5FPbRxbNkQxiMnYzXsuyK5un1Ds7Qs
A6QzdTo42x1x4dR5MiBOFGyhJ0QbkAJ2qvUUIvOzcb6eGDmVtkd+ApXEszoUFTp+
s6fVWHyfFN1JVjxXDfFUon9tEucPqQV0kaPPpYR1TyZ0t0RUq7ERLOWEzjxq/Xy0
riuh3LcHMq2xF8n/TX7ib+IYa712UNNGWGaCCqDJdLdzsE9PWJqxe72bTShfnqJP
e/mBPZ8CHezFGLYxuQ8kwg4FZyrgBqC1wdSmwXGTKtJ2bV9Co2S8GqSSJxIosUSW
W7OBHshGO3KgddvU3n7Oe4Msj2XTvqzPW1P6ehj6j6YtoB9OfjWhiaRoBmY5pId8
0zIxdIzXuFWB2aObFW8EAAB+SAlqNJNy2UkQC0AA3sHkv18DmKInEpsTbi6V88Dz
CxV8rglxoEf0hs6HQFzSQD9Ru3J7xWNSE376FN4TWaRREzVUg8WVcXwTsXWPgVgB
S+eMuqH7Ni4jVJ+bOinLey+DOlRoYM8fLdmeQEBhjQFUnxBp/OD9MzdyBc+rOjwU
v1ecbiRsLatTYHBqKDFbtlbTFpMkSNZh0We87IUlpIIoHPRNJexKSuMnAyDeCGQJ
3WMwhmq1RM5CqfnaFGR8RV6RhuHzMJSQPu7pJMLU2/0me2Rr9dBYj5aNvIMyuBeX
Doxww0v2lBw2pHZrSK5OxU9OKP1kD97dJZSziBMhaeyoZMGEsy7Bci9wVJefluFe
Oth/z0oihkyBktoDSilzMSSU2PQSl4M584HYRScbCsulr2JrZulQ07JA/UDRQV32
nJaBXMbKaV2B2idmdGgPlTtKpvDW+aI8WmjsWtPz3LvYNE78zAlN8KBhSNM7dSqC
tCOH6xwMfADEcPIuDuIPkbSzVKOqhLLpl4SzESO23Ifi7+zqBLoIOEWGQObNE/Ry
94UNjTxcDKyeIPaDW96LPZpzwRimQBUrny1Oz94ASawTax+25X+V2bS3jgCgH9jP
Rlk7NHZJuZBu8osEHJHuPWLyi5JcWeSloqa2T8J4CPPHE+/QS6VwD26Ta8FgZ/0I
OSInwd96yA/Aqisnv7uRl0SE/HxlOdBhg+K7atCSCWNDItVjx1QYjxLu8lz6gBmy
V1RLs/WNXhp518VcneeVANSJLip559r3IseBUWCGG9L7NkACyDlYlZ0+tW8q5czU
1L2rYDhE+Rl4ad2WceRAtdwFsNqd2PrmS/4HlrCt9ljAlTitzC1TxXlXTLPMqhcM
ww2GdpNbVnNHahKEqIqky1/DisiwWFKN3npoRyFlVRXE0RMuoa5PL4IamMCFPgpf
nm+eqXiHuevgdpCNezdCx6O0DvuDROblAlFTKtv/kg6D9l++tbULsApcHJE0Hla7
ysF+sFjaRiIDZrm4zRGvaOxw/dv/VIS6vzr2oQoamkInNMNdfoKJcqikDLyXC0X5
DcqVCJU0Xn1FK56iAgqnrqRpygAYO/5Gqsk4B2qsntwB+JpECfe74iBXKGhWx+HL
etQrJhqj6klq7KfQ4tr2ip6Fz2pO5C2lOcMqJ/IAxQCEIJQVBQxH9awM53bP+WzO
Hv2NBaw4Dxhp66NvpUNInqIaERa1s6HazjZaxLN5WE3kJ30mm5Rduq/fPh+MuNcz
yuceZR3e5K5qYreajKYc0dLU2cY1Gob5udVmbStX5+bxNgTN19MIKuy/X6NDx/Kq
mT8IhXU8jc9zuNYYp/3AsbHsGD0i3DRSByo3WWsRxIwhhTlvlkXB6kSXFX9OYAlU
MR23/dC7cdCzEPBjCFNpMIji08y2G3oo3DIDc+ztURphG3ue0KwhKq9y6Yj/5xaI
ucZLXSG9/Z/1DoY3rq8IQNZ/kPF4Y5Sr8EGy812bxBb5zrMGEaxNjEgyrAdBgylC
o4H2iV5QFEKIJYoeilF16Ovx8YxgWhERKcqLIRM6lJrZm0V00kjSpdSwsL1tFgQn
xp3ut3qrdChL3EiUAwtTIUxuEZ3WUIOd3D7RpJFVm2kl7/br0aOuqxfmbVtvu8Ni
byNcVldwr/m+xK4UgF4ki8zpIunowDu9oZ9jfgazBsu/Kr6NUsrG1OqH31EaHZRE
vqy4B4Y/FF7yaLXoXPYJix7xr15J1kzDMxW9p00xXkYhsPShLN6FmMWY7YLebkWt
c+kX1RUle/19OswZ8ZUgPHEaLWGv8euDNtMGXNq68C9n8QoY+Bo9qQvWHk0OUXfG
dXzXFYp4lzGgH22pgP0AALQSTxWKPeNJJqFzOgn94AnbDoUcS8q1v9ElB5M7yOdR
0nwo+IB6LxPJonAzwiJ3k31FjLWuagKPiTan6sdDRKyMIZ1mmCm6xTWcX7KGai/x
BOgZl/dYHhz8OR5kmDQZ5DfEdVeyy2goTysZ6KuDZ5dD8e7Gj01KbJcQ6ew/o5R5
z5U/bdnRbNTlFsr8t9Zivecf0VAPy+9LADGzR0kYzw/11tbZelu47edhGE1wF+3R
RmV/HKfl0Hm3fDBqKPhBEgohdTSYwLdOvcosBNV93/LSiNTMeMBPoMpf849zD1O7
pquIle+9Ixgz1NeORnF3HecEa/bRyYle+6/20u4AKgsSSV9moRyRl8e/+ALZIsY9
Tk8Cw30REK+tthujyFKvBAYPtTgHV/fILtTmS/1AtOqLRtcoZhw9MtlVRV+9hXyo
uSuDuJUZQTYPwbJVp200suHSK0mnRy7cfG78GLbXKFowaBkX4kzwKjzCUDHfy0zt
3kxDR1zOjgf77RAz9fVowUubtblaLy86PymAEh357zBBJLd6rVb5kw9oqKfP5Qpx
XG9DxG/oVVq/XMlJ234BotVqqBSvM4BBzWysMz1saOzc6zxqcOMTo7LyniHARZoX
QEaRz9F6v6c2VwG9o9azNBA1hcrWMcTsKQYxN/NP36OJJ1XTvaKu75GzmFRTqI2J
9J5icaLHkCf+GW1+O8EQTG3qglO7o7Rw9wncwhot9n6qNp/nyWAG2SU7NqjVDGn/
IGj0kIKP3P95Fs0iD50PO8/AmnVOD9AAn37lcYnjQObSsiC4P6/N1ZugO5pq66RL
ZnYb7GTSnT4q4M5T8Y+R03GVjow7ZD2TXvQgFk3adQLvb5ALKoiNGlm03lDPQKi6
6fENUfJ1iQyhw9w79B9enfwWnR8f2mVYqgqBnUGRgKIdbYihtCVeUjIFNanwx4av
90F2q/N0JWohGtgdEnz0oO+F4L1HS16on+CR/noNUc1cKge0NHWAS/RRbk6XPZf7
pYlD1x6bHiIsa055UnRSgTJnRUqz6PaK0MN9pqvFXGKMNo/LFgSo+cSI0qGKAhB8
sslsf0G6nlHrjIZdEAKhvYMRgYEGh1YW8TYEfJAKbNbNItjtNWSxC1/Vo79WOaF9
JdBZX8NgcnoQIHeVnuCjKiyoRuySV5pg5rCGLqbDyRLLKftISqg6qX6dsJQb6xVe
karQ3mxEua+xTFw/XbOl+vUtc1X9+lnaRCSHtWg+UWEcNIXDJiXGXFZ+kxUDgRe6
Q8EVkXxUXgL+Kw0s6Y12lePN2UmHby5p2AQUJ4A+x/rnX7vl+iodbVu53LK1GmtG
vp8zSbwTMkMtSbJZU9P+6D7XbZvMrJ0WogPlhJ+b+dY9Fc+iVIJo+kwpVs1lfSfB
KuAGFUcgA4NxtzRyt8gP5d152WcHapdLR/C0YLaZvfM+HuCAtvEv/uoUV21+C0Ga
Hr8GiA8ebkwfEZ4nk9Rp+Hp1SF8KpBdhEq2jkMyeZCATmonxRBZoeB0axa+YyyBf
a6hnS/xFDmzuUMuY8Bw8H8cEucnpzLd+ZuWF+rwbRDRzFshCdTVWFamKJLAFzAzP
Ax0x0JDWb8oOS2rKSN6vQAZtxFox8k0Y5DzGJRC3ZEpROIIYRblL2i3sh2ILmwJX
tBo3JxmV+2yBTjU7Xaz+c6001gxDjfVIyqlqB93kVIEV791GbQr5WTQC01X2UcIx
4IGuahBYGFQxXbV+Hbf2KgdD1wjGZUejk4fi6z7xeh0lYWki+EaWFE+DoHNMB6VO
CZQKOKQU0T/qBNkCCKvwQtwkefD2MOMWRZtL+7hGZwyKbERYKRmUd0zVXZYwawxw
XjGs8IQj+2r2sEa7N4S79B/f6jzSKaSleVMU15hLt9QUWqeEV3MMU2xpWqEFFU1U
2FFSbbBo7iPnbFjUBekdmnye5jzoQQIxjQ9QLw7zF8Rz8GTH5D2ybnpZsX5lKLip
KcRBRVi8eYa6aBEke7nNwLSOax0WV9onmBGBB3s4R7HLCoei2nq5hXKRfMxfaXt2
tQzCNwCwVy9L9TEUtHThketoAuT5bEl3XGzKj5Vyb5emc5plA+hS/9hoz3+l97mV
F0dhDv7Jj4rpTWmhEj8jI+vzgM4o8mPWf/CbhrQhBRy6RzOxMbzUQ2/h0ift4Msz
ngMxotBSbUg1nS1tdJPAWry7jXFKFgwkDLyOWnDCdhfdrwZfAbo+dK3wmJ4ZTjIk
tOrA2gHgQGOdo4Gt+2+UW/ZTY1eK85IwDxFTd2tCzrtVrjHsiAZXGnc941M+A2oj
zFOSdEsLEyGhOuGSVKGpq97pVGQd7UrKF/VnAOr/sNC7Qt1RvGraW6ObsazqYJ6a
u1yC4I14FQyPm0GV2NeIXsTqcA47Z1enHj6u0yqaWhS6wumWM0DhCx6kmI8OP9Eo
M3W0Fu2HQZZz3ZruM0q7m9v2km2UB7KYrJGFqXbY0oDduZh4wwS52ZnCGeVS4yu6
keC4E8OF0GF7rsS+9yQXFopdyvhGPxUguSDMzPqJpyl0kU1eXUY9Rd3gioWXjhzU
z90qLYj80pMYJlmf9euRXJJllofmHNPIv3aYsmszPVMoW51Ks35rFozrx6KWeH9S
d1ZV8syEFaTkWJEol50INfOc6wu4HSIgri9F44u/f0dT1/9bpuLSsL9U86Fj8acn
tnDOhMHb/D2e9no3OklC5k1BRThruUDWJAn8kxhcvegv967XzvOg/BTlJeP4FVR5
q6+OrZxK+jcjb1A+vOEdwyejLDUvCOJFBtq/yaDxi0juvEpUPZL2hVoz/u4FZslO
qcVaVp5obJTyMUXE5dG/IA1SdHqdwk9X1WTsO6u9nzcCOuLHos/35ChTOqq5KgpQ
wxmztCJGiZlCRPHVUAf3ZBuzykGI3e8owZkFUMYDic3rnU34y39w2qiIoXIiKRo5
uBmTZJ2ECc9x4Pu8pAhPGqKanseqVou6p0w9SPYxOtrDfE0x5gW/EZUfTKCaYEv3
HYaAKl59O2kucBaepwfJU8I25sdJupe4AnujEI6d1AQAqkxPOPCYRRU2b7UYYjr+
GcFoQolPx4D1310PkjtrxSAp2BCumA75FqC++XjSW5/id20z6WrEuaqQu6+0Elha
LT2hEhp6BPUp0xzc4+tQXlciaksPQP6ZPnBmYgYUTTShGU89wIK+VC999IFxjREQ
75dK9IBjDIQ4Y4soDIHd0Dc4vQH0nK3u8FgA9txuvB4ODM8YFQByJ/AMFiEQhOdO
gKEQboFU30rbWLmw45P5PyLP5Knll+f4smEFqnII492spCJx//ujxOuG2ccvvKtn
GEEgPZpyXocsucYQVaR7K8cnMUJIHWIy4Kedx8pD3IFDrImcFX3PO7G4S+sF57sj
9oKR4B4i+6Hv+JsijKJWs0yrr+i1n0WOvcIrPeOnSvBEyYEtTCG5IaPzuVIy/hwZ
naDUiZ55E1SO+bsUBQgDTEPysadTzTk4lZ8dDwFtfCqBr0tOPLO0yW1j4PoQxdRB
4cdYXdCVF4zqNKWo9PFYEDGGymxqk35zDBJlXsVFr37q0HPCDBpslriVT8SkdWoj
Ko2Q1COGDaXD8UEcOdMRnBDRWhiTxnVcxuprXnLZUAyH/s1mZ2AVBv3GOGwT62Cz
Yb+1RDiDXN+zTmlAIBzZ+1u3O5mKGfPsoS6FWPFyaZRZNo11JzcssuQIj5xj53xc
Xpk5BGmATvA6tIgq2vJ/qqISRQ7OX4x5SmJHHqoLo72EQwtgU8sEZcnsO3qtneic
tTpmlMcpDspBPZDrMbPHbQcHb7S2LqxlYpYX0xAxBmMprsDXVfqZN3yWlF0+feK6
EbW9EguTyZgyOGXZIPbvTuRKC1ClV/G/ZwI6DiX6jSrWG6PzTE3yom2PqjWeDYqs
JKhVjEavxapactivXvPOHEM1hBLGCj4n3N2e6g/X4yqppqD9OxRXmyLlMD6NwfIR
x5iBq0lm93oo8/XmYY5DrgUnTXc3dQa33t5/lVuY0F3dAqLkIj0dsnggXpw6nUsy
jD1hXQl8WxMWdtu+WcUdYDjitYnZTWMm3SbTVvLLGp8H5naLHh2YcwFalXkwY4t3
oeOFpbcNNHc892CHcY6vL/Hykf2EvEt2imKgaj5Zk3qRD7wzMhekMGz9FB7Dwm7E
GWPGhKvGFVXlHQStxH8qISDvVeVAVhqU1YscGQMTsW6SjVOyQ5w3Ca3jCkT4HcWw
LV8xn+iFI7NVOkzPgbXu95yD61aMSpR9a86wED+3b9ymITyrl7H6CJPYv7Yf2PCh
I3d1fca/IZoU0CgrLJfd3Po08V39HesKhdKI2+TAfU6BHMouEtj1M9yQ6MIVrZsR
fRarv9ix6xP5NzZhg2lxw/mOv6D90UYWEwp0iREpEMpqHqfm8WPOBCFHkHK3pNNs
UauYmMoYZXbUVLToINhln88IpCw432tO5CdoO7Yrqvch+BwGX9KU93mHxtvmr+GF
3jX+G6CysCKHBd2YZNengJZV+P9EZy0xFUPzBFmmQIDMSBCFOSlmtj6bgw4GFPLx
RZCwT5kxlORJG3DtkLfghsd3G8pzKEpuqxqv3TS1ZB2eiTcXBiiJLqIKPyyGJ5SH
AExCMzHyn3N/4735gzrLU6vaZtb0zepmfrGL/O56f/CbNxquwT1qcu5Sfl6XkI67
kJMeXe7v0khJI4BJ+Gr3m0hmYObKFPgBTNhbOJ8wh4Yc6vzFbJUkhyZOCXTeQ8fZ
JZ0u9OhGwXFdA3PKHWoGJKC7tXVqw3VrsEx4m1apuepjYwdPriZMZunh/Lu427Bb
Vw88EwlmV8RG/ez7nbyXWo4SMdVDk61QaL7yo5IdLt0Teos/mei5ADGvQlqIBKn7
tpLqDTmWHbB8QTwBx6OxteA1RZXzK/K+WUu8s06q7mwOBcKCy5eprUy39O3FymZn
jc/vVPgKIUlZhiZqbPFCVluDXbuQNnPeG9Gb30mwfFRvqxEyDsgpTpUeDmVDtSzH
Q3dvFA7DwKDA3g+dC+Ypk+xyxJMVi756g307rbS12FRj/KQAlaaADxxUrSM/qBuU
VW7LD+1RhEqT2HWoulEP01K2j+8LkUEgmc+EJOp/3PUh36rU7eomIPX+fWp1paUN
+BoKRT2bkXzgamWVWuYCg42jtfqEVYU9KXkkFPRmYC6Pbz00KJd6zVeUxWRj5Twm
EmBBsrbxk2YznlUQBvhrarh4GrLC5aKPXLknFbw45bVAucznU2p5XKvgfb43/8td
KPxn0orQenRrkC2XMlx+oQzGb6RhoeRLHJ/Ik88yAHotLQJnn3BO8i0cSiTrGWVp
RKh7Q/Bjk1jBnGVNI3kipaKCGXnxvpy6C6Atvhinhsp56YpP804trGr7Xm5gf+99
+wShGRw+frTSDbece4bzHG8xRnlsHdyYjsOEQir8sWYOSrtARGr/kLpqQWHiUJL3
f99ayoOGtYc7lYOI2RfimU3BKJk208lr+CVir2bnwuKjqg0zJ/BuNDPuzWLJIOgy
oSBktYSBCwA1AuoYtq6uVFb+AlMFydzgfzmrxtXwgAmSoNbkPruX+s9Nymfbg2+0
Dmz5tSq5h7V+pOJhupFPCivssGwysxBZivAhKGc3aIf8FFypt1Lp9A+5cX40/aif
bmai9eEzFqicAL1+KTKFDLRqnPmWYtlb5q8L4XAxK4xj0Llto/Qaqsfxonl2ujBp
2VgIxaTo3pF4KbK76PFjVsuOXWYcOEpHuzNX8nnGgdQx67TT+ahESh2r0NW0D0eH
hebh+ftTdC4DbUMCvrmj8ye/5fj0xIluPDwcVTc+G/3UgfaS6M0VsAg0wpCjhRyg
TCR8u+np/Ex1FNyyNStsydjd4BVk5lncc8c7oKtBWiA+ZFP5jFIHsBTiS2jg4Z1j
N2PDcx4OCS43Q54RE+vAnzvLi+t3liEy6xmsImASr6PmaIp9ygjt3AkuIemPA8pb
C9thApCcx/SBJZ51HAqFXb33HBrujCfyz5Q4Sw14D9Ai3RuB/Py+Hj+Ulg8LAk2J
4XNq/Lucw/P1YYzhWEdPiFdY7VUnj7lLqtPZGJomg+jMAAgXfnVENecmqehRNHj5
z0fFeX/T/c1x1hMZ9A5ziWd22EmTztthVzkRBRO3oOgnOKvQXpmXl9kNAwo05pof
YJ954pBdcHMVrfc1A1xeDa22oIfOKPiKQETrVkq9+9CLim86tVjvdOYT9wjE0TlR
31+7v30PGHXpZG84PPyR8zxGDkBVKN31i6uUP3pw1xojFj071mEtpvH8IQJUmSm1
Mf7Y9qPI286cz5URf/RDz29QAMbpg1WKjzu+VtxhkRULuFMdF0NyYUJLUawWP+or
LJdiTINXakMBW3ejwAuP80srIx5csq+TvW0VSz4nKiQgk6FQwKjHNcn7NQYYIMDM
iraLg9C1HdPnZde2b11OXoMBX5sKPDK1/GSBmEIcToeO8SzSHa4kylVcY9vN3Qao
aSpSPYsR53PptB0X5UYicKkWBfsnQUCtnNRx5g+o0OSPiri0T8o2vWeln5Bc2SW4
urxbcT7P6UlYml/GLta5GUE89o85WanjwssRzH7Vr4o8BTRzXLNhGNsnJe8xKRxC
Pg4taTp0FhldKNm0KtbgG40vGRmRVl7zPaSJK8IH3H6VyPDy76cZsw7RmOYVNJoc
Eu9WJ5xO6EMbIb46A6i2Eba3BGgdEI0NiES/FtVXJg9qIz1j2XmHavRVNrmnM2xV
Qa8un98uv1Th0IukAPtCXEXgmjavAQ18faYuFeK5U0U/OQthma5NYG0krgzy/4OA
LSygTfl0/7p6Ox8QIjOdMiowMrnzjddrmleXyhHSenCuEzscMHsmfETvN/SAwbc7
S0lMVnMuATBxq2oCfKlhJY/RnMfMtD88X8MY2eXMApPhgK+L4sx0yS+JWb9lYTUa
VqNCMpmsN9Gb7PP6HKlnpnXQl5v+cXB8GLL58QxihQgfouB/NLkTJNNbstepIAWo
YHwHwOnkJ8z1Z5nbP181URi4yjKUYku/WgEK+lXtMtYQkbBE1Nutanr+dKDjR44U
5uZAohpGIlFnWeJkhwYnk5Z5rX2wnxjaUVYpKrjnDiMs9Rd2a4T1TUS0xTloQ10j
9Ng7+wkqPwITD2JeQWTEzFrtA9y6ZxxKypQexo/mlkd2+pm1azKfCQkexxm7+itw
MhG82AvC16nsLD3oyGyJ3oqPjQeInJIF2hfbs7pV5iT8wcV0QXp0CIygp046pc8r
PKqNxxDcjPSRN7EIVtHlr9zJA4WVjOKA2vdkyjz5ANBD9rwCCO90Io/eNRfNYSdp
Lno+lirFaiVRaj14KjfhLkMWDPbgYq7r/WVkFnmIutugtLykAu9G6X2I5c1hBv5W
iklqiaE7Mikryiw6thOuisKoxk5pTnsU1NyLHei5hqQ2Av0xZR/rqRw11FdIdZ/U
q4F4EH72hbcKFqFZZbUT7MY9NOKEQqDt+UwT7JV/yUP8ooU05A49dWZo3qSEWej2
8FGwnT5TZPOnj/MNy0C5Ab38RoXpGt8Y53GT4KtOBazCJufc//JKoRnl19mPByph
mLo9jaxI8Q49JbZWTO3yo2uHEapeFueDbPROEjMCV/GnUpBgdszLvAUYU5j3uYya
1y0dp1LNLxjs05cMm6i6pMKhWywz3pHqDFYpazDe3SmVCkaoUKztO7xNMKPu1Qnc
/yFqAKbM2BARHTVhEBDwSCy8ooAbVgpUx97ztK61oBWpx3AFB+VfArRegFfhjinE
N2hq6k4iyKAPWXik3SpRPlqTWUdA0V++39R3BDnFHq2m/bSNLZMtHbS0CVz0XWxB
GB9voSGUwcfHp1rGoHhmoj7VEof3rbFLu8rdZJEqCLjuz7tt7iiYyY8++x64eJbC
LPnWzmm+Rm9y9y75PzgBdSD+OglD0UhM78e0EobWMUZkDIb+Xkcfgo8Zj5QWFLbQ
rX8Wk7K4iYiKDpBUzGpAZRPFVhc9u1KHhwIgLWdoPXq9IsAHYDwZmTwC4VzPVSyR
Q4CO6Vf3b7dxCYxUDPw+ntvWvrCT7zdpTfjBM+kEW1XlStmE14EEmJZlG/EuzpKk
u/+94SwhWOqMY6ndINimUDajCnV63ILm+sFnNNJt9kO5NJInrYVt+1c1RYMhyjxp
mwi2TRHtMWFGdBpF3pKGXfejVFv8TDjpACW/0SSkV7C+hajJNvYboopkdDDDbat2
bpzeVXX9Ew32fC3XOXNre+496G+BqFGb6EVOqaBwNdWNAk09xU1eakszbJ5lZA3K
Kk/gaSJ4yI/0Z2yi8n6Qq/hM7JBn9H4xbxuq7qmcYzkne2YyDM3rfIW6YQbpB7ak
M4EzpfJyjuzfRxs6r6jw8FWymNG55SFnqfs6Qg3gsFoEbqo2XZL3fviBE8rBbSWa
5vRidbx9ouY8SY94rlZ1OuwkEfy2BepiqkrNJdCkoN7yt9tn5Hp3eE5rmOp/kE1S
6lX8BB1XoVsZ1XD4bdvzhcCSX8yoBMKy4oOl5lsKF9AtMysv5lH5xF27r3oI+mBc
O5IAqlP7RXvVtbAkPrPTE1v3K5KrkkFLF+QnucVq9oEcYj2yHgEXXih+wB6Hpz06
sCE6e5wTL4qA6EYI99sYyC9+BD54IUzA4m+K65cS9474JSdsYb2Z+ix7Zrrv/U8Y
wpbvtSnencyHZiictDFe9jYhGTk09WTqhtV47PkeQNw9s6wyOW15OLdAVXOvKchv
4wx1Arl7bw1GBueyHZ/SYFhtl4+PwPgABm5cL4UDfTX/eBtWCRpqbXRpLW5UsW6D
D+hfl88TKKGLqgRvhDJMOVwSruCZ7TUepZWadzeJMeMqScAZ+nlDmRK3VRL1Frah
yYS9UoVdrZls425We9m5Qn2XmayRykb+vJCzkZ4gl3D+UGVG2zMdTYO5JhgRKZUO
jPewdDmEyFx/WfLI4tBoq326y812D0UFdB16kWSNIlUIUQKFzxJw+CObjlh7/yUV
8JiOnWcqG0GODyvab0u9WLthKHm6AlaMDiCuc39VkKd/XQUFaX9FKm7MvmG1YYbL
p4QHr0U/qnhsHdxzrMwtstnLq18UgraiNSbTDJ8PPyzPpNnQmLXDfT1yUFFrO2hj
9TQHnLGgj6u1Kja11W3R2Goe3WkXxzMwRjzIgGYMoEK9JRluVdDGvFyD/1pJGcMt
L6adcGZOiVfOH12ASgB/mXUwCUOfBmH6cq37kGjKBSg677eNQj2n8lSd+wYiOOJy
0n/1z5TD+SyVuSiu9T2N9wW4rySpgl19hI5KVDdKc+H8eiC1nBVF5Cj7Ld9Nrcoc
z+3jzUmkeKJXkyFduQdy+dH+een536LbFJ8oEg/dSnWX+RAcva2CWxbDP8gVo2Z6
IvL7r57PdpRURP1By2kE4BhMFjaUGzVQio83BrY5V+4ehqBrwc7P4otg8n6EiWlF
rtxVLqs0jxqFmQGEp7EEm/AOploGTAkmhB5pjSq5jYaZwmi49dXEos3WpUU85NTb
4W4Ja0HM9IlGu8iBqWyfsfjbZeADcXb1zjnWxvkUSZq4cBFP0WpN4O0/m6U9NTIy
lp7e9mGiK6I98LSPfuFTMd1TaAo6JFNGgihuuN7HDZGIxw+BWJ7Os6cPfzLK2Tz/
lrk4g6MFyZdWYmRKeCER5SYpquKesGuN25PM0qyIjo9rgKMzINgOnrKn/jd8okNh
IVUrwQj9VQ7Eyk5uqvMQ5w86oZ1F6ZxhNESuPbuXb6RSRpYUxdl0iv0amA1KfJMs
fioXbl7C5w6uZwMmZeqheQHhdC1WQlmkASfbyGKLDIeIunQr3nuNP28LEqY1PfUx
goOC7fJqRvrR0zd5ZYUAYIgGZ9BUcY6CGMn4fK46tsnkY0o3IrLHxLaWObbQRZv1
CZTdu6A4ZVGU9XPi8KIT8o9egj6VQMS8OGuxFxZO4zbil9zKh91YfhPMv19HM1Vx
zXBpc+TasCoTobBg381DX4aw9e6Csp69GkrtoNNC0mwG7HU+Jjqlg+nMt7WxlH/S
Dm5CC6B99eLHp+B6g1sZESa0XwIhCHSkPJwewLDNlSxc+OKUyQnZUrB8YfuRLdWW
DRoh5a3D5zo5sCEDXirZnkCdlCIddivAnrOeQQuQFGsf6I7tTp5HEXxhukI0bxOz
wZliR7wsq7bsZ6T2ZiL96+sN/Ym8IAFGjCA2gSex0uz7wzqc/rshDyqM3JR2l33e
D/IjzDIURq0Ql0C9qI5ok9BwhmhcBQW10/taDa5V+4mh9Q0rZYwsLXQMOpLqnAlw
soasnEbTUdoJ5KK7RB76pN1qIlUCyhCAVsKuF7R8TuW8mhSzPKt/ybE31V/bW1jZ
EpKaKoxtrh/c92hTt3XJUuH6PEo7nM0HzbRYaiEWBQ5g5WDzJO84LJgkAeHLLisQ
SaWBy7U/h1jKVI+Z3tpsoVMhzE1DRnWFmHawf51jwbPqPvl2QKI1q0a87DOlUjZL
tSRIXRw6BHcw258bLnkOR05EztESgg94dgqPAxw2EYcL/hUCBAHe1V0h7xv5oq/+
bjLJP9HVQ/tiVMnyCM5nQJAkm2/K11A0lBURdmmC6rkJDhOdeFS2WMZZkIBr/sYx
0dPOPTeb6+Z1+/ClIIc6vKKc9wHON7XzF0fi/+NHHRnNK0wvnmBH7GxVlAsKj2WC
6uDwMkr2I8vyBQk/R7RU6zkgTHxKtEECyInacfWK0Nkk8hD73onQ1X/vvuGSDSzD
x/mSbDEgpyAdiXKfv7HDmzYvXPWbzakp3dm5sHdSXlqvYOy1LB+8byuVs0cnmUDA
M+Nb/Jst+Wc9pef4VOXrS4ypHDq3U6n47nODOnLWM0rp+dsx8NZTB3/a2P6QTPtq
30/sN2YgyMA2xFpwX3hynBZ/fE9h5ArGl8J+heggkcz8LGtcmTgqSd+slqSmdQow
WXvXgBWbrFAMk22dYzqmffSl2qhKhEBHjfsOJMhoy7dYUbH9ejQTYRfPnWwwKsmF
LURFXg/ExuNJ4++krAY9E2Afhs7L+ppSqkmw3O9jDj8GG6S1PmhO4tVHzQP84tPM
nR8mtqp8eyIZTyMtmruLAnccxawFGyiO/KFW2rQ7oYERMyH7x9oXiWoV0tAGThv7
ACG8+AMEkPPr07mCxrt5ovbxtF4KPn8XRurxiI70icGONJEM1aLf2the3KxU+5c0
XJrjCHfgk8/PtgifUjiCqlly6FLOMqIDy86dZTjQVuZyRb3/m6hDkknMbfeW6Pq2
eXe3AQPJo5ws5dv2Mn3p+KrPgnz6GhWzcq+tVsMjeZVMM/dIg76N73OGnSnywDjk
nDz9ZSNmNBKHoEfjq6wsGnS3zjPLhNFgjkKXJ8+mWHx7urnMSjfmzHbJPkzv+fKo
nyruG6KnbREHFidMlOwLiDkZxBZMF1utrnK55f5kA9eDfcQ/zFgDfkwedLOnVITK
psUpkzljJd0G411AhBa2gwpnQKoRliNY5FP+dXG+doOKKoioDeIRUrN+rWTnWti6
YDoFwf1JHLqf5eTsfgGwxPkB5Q4gLd3HKgwPwl/YTCPdu4e/vgxLweF10duiGkKS
Jv3geRQWVBPrshS1pwesGn6qSM2jTsyB4mz0ODtJSh8i5gGBm5Hf40pweGnw9hvV
kPsYdY5XCxl0Roq87wHHwOrVK/l2z1Qj+E1QtVCEMkFxJOCE4VuJpVfk2Iwu6NnC
KJlUDYfRCuoki80Ea19pxVIlL+O9NhIQDdGLgCvgdamQUJBAI1Ts2vKtU1FJNPFV
tDzKpp8zlJxLRnxW+1X4WoV4n7vxOntPWiJCa+SVT5wlhuaGspI9N/Q45vU4GcsP
pfGjtgxGyb1Thp3G7KW3QVyvi2GtMOYpDi+Q/8sPcOJ3oO+wThogxCPK5QQhohwE
cfy0UOv0Ucc8rGlN2UIsjHLsvpn5Kbo4HK+tziBj6lZ0S/qBUmhOzPZi1kC/6eqT
RDfsmE+8hrrgFSckROG9uUazTgej4P+kE491k38Zr/TWzDdeJloaUdKu+bzLtLq9
k6Ig7tq7O/Dd5OQK3hNF6xxh9/0m9a8bDDFEBAMULNirflYpXgde5Oqh5hFj2luq
ZENcYpO57h+hgPPGVDHb69nlaQ9/sBFE1h3xFy8ghaPlTGhkU629Oay4abhePQTd
L037QkWe3lVzgTKhtcyWH+wvyVX2R14LiqqkndE3ZimyIk3NF+jY3Hq5yQkL1VMA
LXG2zJ9PNxl08/fs3DQRdDSInr/Sz4bGuQluaVuXmmWqNmnM/F97pN4fs3Wzux0G
qg3ZA4doH7Rurk5OGei/3FPIRheXsUQrPpJ/wedDpLqXpW/aYHvvOVD+nm+pgmCK
8NqZwS61pqBGS0QNPLVGY5WBBxNNysp1wdP5XkThOG1UHefJnGrJT4ttq9w5RVrw
PuC4kHn41sl3cJRDJ2pD/3030xneki3WhNhdPsO3K4ZQQ2qyL0aUYp+QzzA9CLFp
AVKbYITvOVNPXUBoewUbvnU8sHtuby8F0SZb+8HUHeWM7EmCrcWx2bCv49IpfkC5
ZfucMb6q4tNhy9IaKXGb42Gc5I8s2twrciZ8gqiT4yYeis48FUsB04wu4R0Aj6pv
ks/kg2AEj/XLTsemNedzWSVbNv8wOUwSUnaCohz2tcriQcMKYsWnum8Xip1rita5
xKyNivcgCjcf9cbLpfscL8dGI21RExkX8xVcP1hUeRQP1PohlRnYlwFRmE3e1yA+
RS5Nk9s8wHc/HvfVDJgIEx75UBa/RNwI7fsBcJXIXAFVDueRlHSciQ7jcd5cYY3T
IzS/o4NmQRu0B40vyFTa7xfZ7rUPyl90BkBr6x71TlYwBa5vSyutKko6LSTJVDAp
OrkbMMgeHRJuwJy7bt3mDoCB6OzpxrLleDEE7Q0k51jazQJRZVbbJ4HdLZVsLOJe
LzLR9HrJpiI/W5719jrlQS869UiSLU2U3h4e7gVS5/bTp/Wr1e3Dr4VFwdC6UwPs
IDteTCDkloA60zsHeO8fmT7QvSk9Gkj+heDNUSMtP2MpjFIPNtyK/cNkJdxh1pZy
e1dX2KIevxXsvbw3txN/JKTs/IFNqac8Oreb5ES4vayFiFKRG+6naheTte/+eTLD
ikh9kiOPDT69Z+tVENNXk/WU+89ajudG2h3bSbKUTG1wzmBD9xa0Js1jVRPdxj8P
HdHJbQTJ7qvueTD8KoWrI/PVRnFwftFySfgVj3cpE8yZx48WS5i/O0C5QLi/cujK
XYFo/MgeBX0Z9EKOOMUNf013tr8rL9iAdGrYFUSUOPahNg7r1XI/YzrOsFrr+71s
HLEVDeDp8lVhVeIFkNxSMrckIZlxNlWHZbd4/0/XdZNBP7G4MEJ3pDye6IbvEuly
zny4niSX0ZWMrxbavvq8Ktu5A05Rf/1uu/tpTyO1NMC+IuHMTr7LfItlF6+juCAV
Sr1BQ/tf3rmqEukwgTWEcTlT5vKm9C6HN+oKKqDdTU/gHix7R1Y4fSYoRuWD6Gyb
k39E1Rl07ysc3dV1aMbcAMKyaWhgQi2FDEjf/1ClYXz+cluawBpvCEQHcvbouKxS
mK+Ax3hGlSr5N2/vXD3Cy2SEViXoKPkmbEpl4JtOSki51dO4715M9ggTfmhk/Ak1
6S/WeNTp9YwY0/y15BQEAVzaSv26v6TN04E2l9DshUndzwvr/Lb8e1JbPnz5k5U4
PEFa6I+IkQdGw4iqMjPLxMkoNI3MWjLRu0VNX5nxiHnopjHINofoRHzOSgbRDaKA
4LI9d2/PlXghDhclO5YeSvR3Nqldo0hsTwEgGhAw11JJHphHBHrLzBdn7TVV/uJi
AUtZnrCIp7ypdkH1+HWKP38AcYnO7XusmsXfSiUiSqmv+FIC3mV9T8+RHNBJa96C
UzzOVJBWBjVntMy+lXXj2WDigukdRqf8j2U9jeNt2i05ZlvqCWHIpotnhloJrLnb
g4Nf+lrZY7y1fuUTfKxDUc2bkKaFRXkpy6TmbeoOHwTizLyRLsiKNcBiapBHpx4v
Z1FKdxV95oUA+kEgzqAc1Jd6DbRl09i6DDKHxI+7sQLC/TfbxhTiBzsinKGsi4WO
BKg+LOADqm2/5DFx/gr91FMpKI16PuLVR+VOF4mlgejbS9BoN3zExqJ6QhDS5sg3
429kyiP/Y7d3BUdJ5LoxFdn3QwTqBSo6rzwBN+gaHwq0dvjIw+ZuXUp9+JpGBl/w
Mo+iCdFoHvSbDfhXiCYrdK9VyfQmqMQ7oQbtNkCm+OhvK5N7rY89LNl3cT3dkFtf
tVFYPs/10btDr4b2ITLF/SoZ0cXil1H8CXIbspsN6PtSM/oBV4wR4k1dhmrA7tnn
YMbFrtyvX9e6DDSGooZC7d6A7sBcD5VFG1KxoJtKfMqmuoTqN3Q84bBpRxAtaNv0
BXKUgKGY1RqqhnNi21IR0830+CKq4bbYutOZn+4sRRjJOpCm4TsPiJ7r8SNmljW6
J5LkAB/jzhO/OQs0QHs5dfx+c3rGmdpy58084wI5wxbm0pa5NXcGPYBO3GSw0FeU
eBXSxYWcv/5sHQzKMAt3DHCgqvC8b06VBULnVMmDfK9yOPBC5cXVMVFIUNb6YYc0
xVIadunXHpsIjjefmnOLi9JiTN9RVpEcjC6f7kY6akwX+ZGqSPs/duhU2LjomCF5
xr4quIgxpuvgExNHhaBVxzch05fSwCF2Q3q3ABwUix2tcACxIhM0VpHrld9iAJws
7ZMmfNxGOc9WXsvr2higjO8H7exSlUG6u+BuQh/TitRHIBAQk+mh7U7AEuaGaVIL
P3AQ0OzlxDZ7FHVHsG3iSLzts8urd8AyiMSdcY9fk/wiX0fKt2htaZOCYG9XWOiQ
eNlwKDimnC3SKIIUgR9W3y09k2hBH0WrcrJgKYUBifLirhL0HwgUQoaFpikHcU+f
SHb1LacUVEKmPxhyLm065R5+pxNYcO6mAizMxizUg3fJjr2fSvTH52QHgX/L2GGG
WkwdGDgmSdq8G938ZasX9W3w7gPnUinIib1/QcVjyO9yjoWRn9MNfV0ID+69VUqv
fJF0gEmDjv5pLqyG/kzzEvAdh+1VOfE5AD4TSg1gqT+Evgq7G8eKdzOpxI3i2Iix
tO1gjBoe6ioT/4cNtkvntPijqSc9tbb8pSwjCM5cel0Lu78PWkFsP36oZFeDtRaf
OYwGKYPAgI+Z2vx80kV61PFEr3COWaK6wc42gQe4y017piqEd57+jpJIw4qzjeTr
vTCOqfzJzCNfLitCRL0T6QdHXbtqyJhykm305Q2fL5ZxXnKy7ineY3Fk6ffqSmWe
8iAKKZLIFNNTssxMn0EnQjUp8YLhdiogR+ge9VbC+nc57xtHtL21r4iteRZXZWPl
t+1VWi6uuykG1Qz5+5UmL+K58DtI6hkPyGj3tzKSSK8/QjQolwp3UrCKkE7Tm2HJ
tAHM+NTqUaQCy/tNIXTo3XTJ9nlFIo8uXfDLf13K7uide5naJPnuJ+lytiJt4XSx
Qhj/3oHK4XW3s28WX0oO60j4TNFSpkyVM89Sx9/llQGUQIE3gnGy+tZgInYivBuI
K6TKgsN/IL7o3FqM7R/ZRlS7xBTU0xEbWyTAjLT8k7bKFTwjfrx7uYqf/ex7PMzB
gGwVCJXij65WEipLuJVs4LEvkwJjew4Gd6HU77kTIIMjLCGhybu/Cy1YGOQmlIsg
BBuzQh179P7/IXnv2MopWINwdx13ajcy/4qMb/Qz297ZdHZiESK6wZDr1/4/r9+8
iYlhIwpfqarSG4CoUsaVZD+L9mCJPpcIBCI7m9EAiZHkEQpjR9IUgKfXMpZgY72F
tTfpNckHPVgwFpb9YMkk8bUg6FhW3AbXtYcQ+PDTKNvjo1jOePBlx376/xlnIZiG
Ss06LJR8c8jggEwfPaJ06FXEpIENBKw/fS2B3h6UiKQLQMCxMCPOMxPTzrgWut4d
nfeW+zdZaNjdj/VhZga5yIEGMJynXfydOaDQn8m9hjZ00A2XOn7cVNPmK1aNaKw3
WZCEknkQ/odhNVNnLImszuGoNa6EomEfBGko0KcwdImJ66/cIbcdcMFZ5M928JQP
UGoLo62M1F1vxc9Rsagcj+FdG2AF1YGCzZcxKakKktU+UUyq3PTqNsVBDNpVEvPN
njOjWSbvSAAXAnVy959nDLRa2EEhIbhuyS64B75GG2W8WOlgCYTNp0zVEXr9tHnC
VZFzXiqNT2ZkD4oBv9yUaNVttutVlrP34JnIcuVQVSC2HzNNRL0dfSdkVDxC02l4
QEc1a263O2TrDf1hjgwTiBzph5F/COMAluA8ffLzNtWzwMYZJm+GKVVus+c4AQ8s
IXr3KI5lQPIrqNVnseJeDkvIHL6RwA7AEURipzJKb0x3qZSWq5461QtcGX1LTr0s
LOZIbFLvMa8PMwHUD34Uu/ctkbd4tlxwfh5ccEV4h8dstHVSFdS/aFkdaVVDJKWd
L/0XPhyCw7m3ATl1MR0FiATyA0O32IOI/YchGzYPvFBhcBUSVG6WD892xzoMCsF5
BMxgJHjwj5ZNXbtx5+ZH26AtGja+T3nf15LRU2rGyoexfs0A8FtvsF7xp9n+Rmhu
gz81ulCCbo6SD2JfHrwLtZVEWjYOhWeWxOEfxqGXGyDE1GPTitMyhowELT18ho3Z
i7jwUDnJX96XpufTu7/z+psZFVMv+u6RBg457FbJCVUhPqsbpXiUQ/PF0gF8WgxD
ocZpNurmWp+Y/TeLI2Tdzv9pAwvSDMSjPQ5bQR/rZRB+n23Yr5LaBb11ABYPZG/J
RFg6FkaiQmMcV6zvOY1Nl+MO/09RlMA5JR2G7XmiNEwidh6zmpPJnBnmpS5DzohG
2W8f4EZcxMpu63TDfCDuyTCI2DdacmQmmoBuHcffwshQhKeso4xZaaydes0k1grO
3Zvih2hPU3l4FsOdPh8queTJijWcu0xsZ3zZGHwSqACWxYDBcijdq6e7ywfjBX80
0DdCsOcmZzHHl8Y0QpH4ZokaBNI0wEfr2WygmhiRTu99ZBoXGMj/gwIf+If7NrJ6
b/t1b77IND9szW1usKsb3d6QToEW3IVVVSVM97bj9N4fWQo9LNDsBzwqIUscQ7D4
tPzsT9brtDfiMrjNHqBosDC72CQrpaKAiTsSdgF8jVtzgHU3PEx7J45wPMx0y1aG
0369inP8JDGeB7m4XiibIACrag1NWGW7jrefc8bSPQjc8LdRB9UslbhLCvnQLRD0
0yYfkpDqbs1WfbjVqoLAVwFRfDy8KdYZZSD8CFWsyoRLwM/0oxii4Af+RhZFKoXx
H1154D3EtFnx3/fa/8vc4OXh6NlfStVR0oLAjxB33Sp8f8B4/GdTTrTLibpBs8KM
+PZOu8XdGhuDXgC/iQ63/FTOXyqa0/JBpUm9YEcOv8JEcbFvTWEVcy67bVPFKQx4
L4U5DWKToLa8A8MXs78P2S34O8g0SK93KvFA1UQVf1IJHE5of7SVSj3nJb0pOgKo
PzBoZ3JFbBj9A3dbV6ypBXdRnK2Da2EK2Pun8ACXvKpDDrbGQ+WfuZQTEA1vNAeZ
NSze0/qgqRi8BqwGK94Xg9pKluuBNBDbEbF+5FXCmWCIeRf59HNhSZMf53T6eSJ9
DKc80eJxvCln/Ep0ZRGsHT/HWYj/KHfOBhQW+Kj/SH5grKnXbfcco1aceH6q/ymb
iC+F3aAt9fCwW94SAfj2wR9F7R7objBOLK/jbignCy1CF4ItLCET0f6IGUeHbMCl
wOup8uEIV2QM2Ckg+AQd8DrD2Ww/nI/9XH1cauiO+vy4LXJz97Zj+QXo9YNnomH/
RtUqeeLD+Uyh50v6P7r1ue50t75Wmia4VC/ZI0RKq05Lw96zjqdFH0pmCRcjQkhx
44fGgI9W6hoUqHgzUGEUjawldfbTtMltV93GvD8AOphIgc9iRCBXejHhFCJxxi0E
ZPnovdpb90O0V3PE3aBugw4BqsyVPyo7o9ru6efb0GuLtDDRkUbmu5UF+KXLZBpi
kjZPkZY00ckfHaRURwecJKze/qzIR1UbKxFQeSdQ4OJTIImF0jd42rI9rHgdYp5P
CmW0+I/A5GzNXEXIH0yeodoVS9HWqqgT7k0ffMIrLZsmKG/MFyLWMRVeKvA48Ay+
q4E2D9Qx/fq0bgcyOd/ZtC+u3Tfpqs+EnNUAkn+dpb0A1nl5bmETUtFgHfDH/9Th
wLvdDVukYMzLgkI8zblDwagotCwZjhyJ/tEXu5gWvUjCS9Ve6pmKRP2zom1ThHSx
kNmiBkowTN+N4Rsc2YkiA4AbM1O3BIYdNtu9IxK0MWY5ViB0Y20xwoVMkt04Sq9W
Omcdm8Qc0lXDneuBdub67ptgnU3jORkMsHPYW5GPTlpV2liFo6SUdot+SrkslqV0
ZWJ4juYSssiQcEi7KIP6kCYGCg+7Cr3bhW0X4aY5MgeZWPwam9nBsFEGTSFdcqXy
ysZe5iTMPRq3Y1CwMfvmebRvcUzG6hYyO0i5x8ogZxAMUAianTOD2y2qRRvHQomf
+Qhj5x6adOFYByoJPOG6m5qLTnrPoITjdHcwPHWVZGXET0tfF3IJK+YY5dD4+bxY
xX7a4IiggbcE4H0V+8MtnQUdE4sUV0Ct+RCYWxj2FNVT28/kHr2bY2fChmWUtvA2
SeAL7iXAzOxjv/heWZdak6gcs5BFh8HkoGXh3jH924qYkyUoRiB+ym7M2mHlTR0j
T4tayTWthBhGieN+++ISfhlg5qxm1een7JdvZgMFW8L9b4sL8jIyooW+JcagwL/i
K+V0ZPH4DK7wcYZvJqgtcrmOxHCzkmDnfhGdCWRvhLtHvUCUvtjxNj9PljvowzOq
JkGp6kPITSAR6AfoK+QBaCWIoMtyrLYiA52HG6MOxEodItftPCoXr/I8oVfL59ms
nFoexBYM5xIph42fqRto+Hui+W+EjSAhvQSThbKeVFyKqfWG4BO4z6fBGcctQDmz
pWK4m4yA9TtF3/jXS7FX889oLrQkX3Ji37C+xuo//aOewXg6BixGHpFMGgka9lz3
fobQ6qJruatpVvrlKslSbgyR3/0MuuarnGGH3Qqu1yBU1AzN9PQdsmYovzuYcyb5
lP+Ojmr3/aPZdiiZkX2Ki2Yd9kSnhMzS+Sf0ihaMYHhItzwl8UA6Vh5Tts2EQvTG
iJ32PmIUTHpz3yXbxs4JWDWvMscXeQw7b7kfdnHNdeiB8AtmlsC5+J2EiS6DwW++
iMB+6a1P3IhP1b2sZvBnpR18boDybnVY/+JoN/Pe7dY4/m6+SBK+e/QOjG0JVSgv
by9HHOb64S4yl88DUXlHFNpX6Nwzhfxknbc9z7sRYK3q+cxAZOwsRZ/THqDYC6WD
k3jdBzvGCafSn7hLDdmyJ9OarVarKnA9lgdBXGNmteEKzfuyu47jSp4sqg9Kw7le
HXLp5LmGVfMSRZV3JmJ0c4WTt6at7+KP1hzQVhICDekjdVChTSV0rxu1A8K1fq/4
MMLpCFfoj4kko+PzJks2iwgXaKOn1Q4WEHKWmNeLqEU8TaTzCbnABkoWpm/1UCdg
tJHQnICmniIbKdhd+4n6yVUUDxWbnowCZIe891CguNnvB3xn+CeX71sTeqUpRMbu
wPtjiU7h/u5kcLgPAjpkNvutAYNqsRlDhG5olt/hM4bkcTn3Qyy3y+SREolwUJzt
ZzibANM6KKdY6VqRg+AgihiMcYWsbtDyxUPZWgmWIAwf0cemnCXlY248Xgr6A9RI
Z7tiAu0mM0ZsVZspj8xcKuLYyZFVqSIXgFc3kHU2g3OMS9xT7mMOibW1OhyhMXOb
8zg91KeD0xofZln6+WsvHxSjeVzfiW01wDed1lCRHtcdl+awsvwrRin9+KcWOTLe
WQKAiQFMFKX/RN7jbbkRdkgGc9N1foeBMzGu2f3NE7LrgWEh9jhIAP8pFDQ0aNKX
ffI0RmcTAweZEA6bhTNCO6hpUtEKIrNY0RpxdTdAFibSOY3UG3p3iABHvjWLrJqe
QKAo07BZS7Yn+yhXjMAgCVoaXW4sgIysEmaujoqe7WSExs9QYv87AXqZBmaTk71h
ocD1EogL0dKFJF/teUZQa9/QkCQELSIfo64InnAb3lt8FubgFTjhg9uyDycoh0Jv
x3I+TxMLDOjhDcC5h4ZUHZg32Eq3+kBd6wHJUpSQyxl4VkJ8t7X15ujRX+kfudQv
Bz/8Mljaxzu41gDAiiMrhg9EU4/Cbu8OXbVGRnUnWP3GUW5cu2Su6xIegmqhQWAp
SqFrE7AqGygPHvokYUwzBHtVRdx5AytwtgS6DB9l7wehBtXEGPV1Acsvvjm1nk2A
80FZ45IQ2LQkhRO9q6lHsyaFp43L99aE/Ifeb9v5VYwUmKCCLK1efIoKFcN02+C/
exQdnFg/E363y2Yhh+DR8qDjQ0NB2d1nKNP3MrJEnAUKYRpUk8TYvoKJY+Y/o8ky
01+dqlk67oL+Zr40wTygzt5XTpYQDgFl+bCAb3NQVR55KM8gZvMrslknVrCWryV5
WH+xpIjWtylCT1xNSn++xqZHp+XPLzcFS8noxYMPFtN0i2CERsOdMTJYXtG7E9OP
FScmoQwkZTqN2X0sh5VULcDfGpt5w1nw6D3WAKv75EeiKDY9S3CbnW7R3UQ7uzRx
e3j156Bzt3Sl8xIG4rNJdx8FeDwM6trYwjnzcGlKcbbJ8A+DtbU9TnsvyQlNkqGF
iZlUWBeuk9guAyP17JVbpMXGd/wlc3QVXBmpgIp9Nrpl6LeXXUScH2U4WWzmzOm2
L9Q6JEkQcPsG7WS+f5Bq0DWmnBzkmmTe7/+smt9SaFNrHx5RDgr2XAmo+AjYVFoO
rytLDfLrDetk9I0SlFVIZWp/HUMRI1eFRfllNXyk5lHtyTOY2FeIOb4uFN9LWlj5
mSNZnCCwa9XubOpzXGin11ar8Exiv24aboUrqZLfg7nchUskBhoOfCZCPV6VqEAa
yWSBu0gt/8aslbD/xmUCDT1oPBBKdTv3fY9iNVgNmrnPCoHzCaZxtYmg8YR723ia
WFpy7EgKQfcF7hrj6bIQ0dNarun3QIkf/dkHgzzc+pmMrFBx5BXZG/+FzHz09DJp
Uny9oECHHWWL22gRjIrUSqe3uObOJytAWDohBsCBZ5gDQ5GWEPzw+Kqq4+RCYcgi
XRt+4aakihx9fgw+zcgm0h0nhCgfQ0MMTgCEke0aKfvBtr4L+0HFlPUtHnT6uDSy
lLHjVFh0thngELewhAzjwAiFSFKl3YjeFFIq1W9cPvOPYrv20SzFhGs3glXrIojg
PstfnE8EGwCTAgHRye5eGrMRYlhg7VG5QyI0vZJNfCBS5e/eQqzwg8ItYN6iCgr/
98prmRTJuJTFxzgX1mDiGIoN3Fv5UgWjdOUlolgY5TOXl1OFjBtWWnTgOt9egKjx
h1XrwlBDj4lioyBSIXyJz+kIzZaYPqTEaKkU5jYy00YA12hpduPH3mObmUn9LLiD
nnORc9z1bNNH/dszCIQInnlrOtoQQPyM6hqzHiIaDACwBZ0gQFbDMyQT9Bz4vQGY
J607/hDBV7AAEN1XDmg7BIZM7jimy1+9BCz5QkmrOLzTK5jVg+FvhyoulknO5Jcn
V57292YtInYpCctR8kCqa/X/MhPLS17Vhx9c16NXIcHk7NCw0kGopWYif+iVfrWk
nn4v3Mnv5fF6Rgt5nj1fVxbU0EYZ+S/WH2QuYTk7E8B0wfH0gLkz3AbFWV/qPkTH
EAYS1CxIAj8T3stIng9eBdIk9cjojmx/0LmjWBpX9QQEFBxYprcDXwBxWmNTDpx9
uRGs8UKLfP+jKeGgwG4Yujo0NiE75aBllABqY1hzPB+DXAQ33SSOP3lPvt5MwnvO
hwHNrl/6CSVA7zf3pTxxC3MxbOne0vCg9h8a/QPyUUJlBhGx8lmv0oVo+OGhQH4a
hUj9eC/L/vyst9+gIfjBjaYS6NrgkaoM1mYUt0YEwroqhS4SvWwwzzyZeXd1GcHG
R2UcmWeQL0wcBogogMtKXFbVcVdgd+9K6pHOFqzswTa9nmpI8tUHztvuLTKsV5ID
eqx0bOCKnb7FnQ69Fam0aG2mjln4+iJlW3SgelrIhgFkyUjfGOeRZOxEV7WFXXQz
3wU4/J8V3OEt4KMyeS9CesW8Zfl0VqKZNJc5j1ttc7N0AZLFRjb1K9V+Gqs4ci0W
DP1s2+NRV3/LNvz8DvGQFy+jVki0wGloXH3r3MX7F/3itZeHFrUSS2jI+0bVw+LK
ae+/c7Cv4H5ml/QDu0BqwkxvO/IUkB7TbUsLHHWbfpd87Qtc3pI1ylZ+dWmUqUYq
qNBscLTDVJ/MOZdBOnmUqfB91OikuBoFDHzocLgOf9F6hdyDD02Yk1hL72XVpqpQ
W+wQeUXCfl05u5hLEnT5q2ZI3eTf6tzWQGUyQaYWF4shWy6z8C9lVko/mgYVawv8
z12n5SNGOO4iOxjR3119DBflNJ7tWXjjhIYLD8k0EZsvtqboxotFEa0+LI+FYH3U
6l4hgUiGx9FEE3gwzm5ufrkGjVq5PpALFr44/LNAT5+IK9xlmHGkYP/AWnRkU0ZX
NqSrlN7ViLGDUNWJr3bkMuNRdGRZhD2WxiYT5bmw0XUmqOV9gumuyljXLzJCSzxK
p300vflACH6qbxVM15g3ggRhKxs8bPc5osSPGlDdTuer0v9NII3qJjOkbsCOT/It
E8lnYnQ5wFGBQynVVOYiI/aSYzAD9noj/Cu4chY1HNJ89v4lQEfhKXF18XcEBz7W
9lFB9VE9x36N6/bHuDQ2eBHFrJPOQJx5YQ6dB6BEb+nWUj5IHYEqBCNwz/frxOAg
7BxNigygFJbLfWA91kuZcceQuJH9h4CdG+8UBs7GwShW3Y0IQucJghyJNSwNkdV4
l67UksvERChBHX9tSA8Y9e1IjcDG0mJ0ZJpAmjEg6YBYxkEIekdI2qFecow8rPzk
CK4M9Vk4Zcnfow3QtKza+9q+lnFvRRgu+mhMEmy407d1elA3QXAHCHJHLAmwp6l4
GoJ+s7Jas1M1MEgBevSHZv5jVh1Nsjwhl1HkrwOU15fGjFew91juqC1SoMicMQmX
tgOf7NUbqaXjkO/KqxzaUkOG7fG74vVmudAIWn44fgMRCI0dldEAHorUNGDq10/x
6voo0/xSzCRPQby/q1SUlD4D59lXr5j5uZ1xsoBfrsTgwGYdKd1NqFVeK7hVIM3q
fy75vIwL0JwRPyKoKvB6moe1DvUBHBq0BhUTRPt7tQcmhc2uNZlgKwm/odA9cadn
1cfvZfOaJ1L6yuJ9Y6g3ydEALzoefUtZhImwczPLaw6AuAtsoOvkUMJY83kj388k
iV5fvolk9OTHbnmBSRsNbx5hK1MdScsB0YVFNvHRnz3ZOrxZDltuHfCiT7VUUk4/
D13kRK7Wd3JsHR4osr3FOjt6y8nbvvIlhLHBZwOC8T2BpNDdH+Tvsv96UQb/mRHP
4NNJSZLatvA7cOLdfkmdYBnLNyTc1x7rSszJF2DO1lHH7z7yrEKOEtnOLxrO8Sof
TQtpLdfet+UGDjsXAUTzbP0E9W+PlHjobYtHigsrXQTPa6k8uNCBXYdfIHAkFDEB
olJs4uu9i3iBXvDR0H8I8/TZu5U8UrVarMlNV5NuIOQwZHwectH4pkmrKhFxcRQM
6iV1sEdEyqbJlGWrumP2J26Sr8GuJAw/owoM04a8DI1qMkGBgWIlTVSomHvvlv1O
8LXXhNqXsmKta2KJNuAXW5AyQsVMjWjvpF/6e2qbT2WzsUK3+EirbEQx2l8uxoDE
vz6hCsjClsskVz9u+HNZKOsz6x7ywAlK7pGZrgrGTLATH27jXv9MaOYnx6KbU46B
xAvtkipG7vMq9kTMTT0od6784KHi4lNbRw5PdPVpjRMgt5gdA1pcb0Jz8J6jpifB
DfnOfSwxsPP7VbMDrR52+z7uqh0hgoQEfol3C2VU7wg/iiO5IxfgM2u4NUcErs0N
9EvftaRe+TV1id3WplxtCNHSGsJKnJzgwgYd5v4oXa3K2QMHP1Z+ID9FwDUfOdrZ
d6WgwtnU+EwoknmuVKYP/Px8NnS1lDNyM4SNc/xKl/hFMs978qqjCBoc0AvyyX7o
KPbgxqIvrBCp4iphXmKZ0JrH4XRxVF1Ny7cV16FOy0nu1Rw4tdDHZW3DkBDe51Jg
lJi1W8BspETKhl2AN5BSCwUtc7UJt8X4IilYUqX4+aGibNDJdkelPjjQrYTsDYsn
dp27RtQssNsBMi2nPqi4pWkagf/yfc1eRrqcARJBO9BedWaImoz6StfPrCM8u1DJ
ch8bzjTlQJOiHMjVlKjUm5m8WeEapYZfbB6ijx4CgVl5heOYvNl5doDcMkO64CD1
G819ufIjh54c3xFdzP3bfuhlQJeOE4eVps5fpB7eQ48VFnFRspi/qoeFPHZSfcAM
TVw/Kzkbqf0xJd4NY8caJF8JBV6W/YSSuCfctq6Pxt3wQvXMgcezazRydkLLo/RN
VJF//x8dCDkuvEdhfhR8qBXifLTejfa5AmWWY9XWxSPvE2kGo1YMktdf5xQeOhxW
lvJkx580Zdfh8ksmsKPhOn/Ma96PThCEkVt4uUTUjhcsuJyplVX7eFZXDN3HV+Qx
qmM4xbNpM1LAG8CABbm0kumJCxmnJsaKf9JyUVPwRDTipwijYf+z6pyY9B0lullb
GIqM7udsyGksf3zyBlbfJamI5RTmz0BuWXtFJVteqaWDkj7BTxuBnkhg5YcnEPT5
TnDYu290DJKKeBxjdD6kZOQD7cvpuywnsKkpi+sKQKvGawf0xFcfhv4mXL2C9JYD
OnI5DJtSA5Xpi2K8qxiexNWF8oSSx32IoOGMpxgqq0DUGvlfBKyW8/9LgfsXgpZR
KQPyK6EWd5p4hMLRom47iLvmL3u6QGnp0wKOwqPBypgRxyWw8soC04xqAWU4cuxF
Sn05Fz4lXTjnA3i+K633Qxy4J/S0N9wZIvhnlIglLO94uq+T6ojXnMnfH4+NCp3E
fH4lzqir/fFh50yjt4lorGtVR4wOPoOGcJPxBAOSwPR+mkadS9oKw3UUbbHfchLX
McUWziI1ZmYLTIEmKDMAV3huOp+5c+9auQpwt48S5Gna7sCbN0RWQlcqAXvLz8mG
c7Vn94jD5QHPFK6uVGXZ+YPKpHHKytQPj9+orR1Lie32UIDo12nAFfIQW+3qyk8S
jRDsCle0xDsScV4/PwIrCenRYJScu6YIS3LBa/3F+XgKy9aufDYcGemuJXPmGU43
jb5u5LZAAd1k1LH1FilyetQG6SvduI1CSamcZZ0UvGevLGnFn/LAAq/Vt5dY1fdy
mwpevZtilH81vnBfKyVZJsfYLeLqmHl/ncfPXUzG1c5M1fxCV+MxJEAEKvRha0Tc
RQ0gctrt1t385qOT1ixtNhlc183DFbHMIt+HutonNkRBiSlyRplXq2jYEQSlodLU
KYb67nxCwd08ESDITznNp6uGQqfHOk17qPrYcnKNGfbHYNVYxxizK5ClAXKgZmqW
v0Cdf6Bm084z22c9Nl1+FsCEfa0lfIDvKtNMeVR3bfU9U18BN9RgXbFA0R9SSetY
uGNY5H4e1Vvt49M8R+z+3h9Jtu5s8YxFUHRuNPhuwkx3bLYVs2Qtk2XcMUIQqwZ9
8SGVPOyO3SLaafeUZ/5A4yd/nDwqBzSDIxvb6/sTNB11bv6PBhr1RRurbrIEO3vd
z5HkgVQ0YM1r2McG1iki3LljK3uJb8ngi9MaSx+g3lCVildAPtEMiSFiJ8vHkf94
vrkZGvxUzfmLs/pXDvdI/BCKyDMGhwW5QQxUm2fU805am8QgCSMRprggw5N5tJpn
g9E7mRKN0yj84NNCZ1l037MV83jxO4QC4b5bSDqsSFwYL3x2cBpMh6bmvHLcoNHn
/tnWFCDNpNwuFczRRRI8cy/M4HHTvyuRS5C/sbkqPewkd06EeBbZcHarWoWfaJu/
uGPV9fAOX/3C9kmN9BFB0wkxIteO56yDNct6To4pgidyCu4OJT4uhui710SmlOQc
jZbHp6+6kh9S4SwxT8we/b0n57LWnxipE6GqK5eRxrU91e9t2iTItswbjbtzijB4
zDiVg+2ULl2nwh8LZVdqrNDe8n08NXYDHyJ9dA8TmAQYoiGeUn0M6xumqdn6Mofz
AuMeM5wfH1xzHFDu8RrWlHIjpxtHiqRec7kbJOuXMkrILshVbVnYCtuFHLMQjV8c
eLUg6dbSHZPHYwlutcZ85gr24ys0+gwZRBjg9AmP1hNXgIw+BS8afofQuchno1Ea
xZUlq4ASVHhYRMzzgI5oFkj5NRsOWEf90I0dC1wE8rYeMEQn2vt0kTfJutk7y5A3
uSY0LZY6QoyxxnQSChkoomMAw2/oT4hIu2Qwmi69HGMU4B4MQkmisNabXjDD74T4
PCedMCkxIvAkh5cCJiYMzpl15l6vYouPwh52ySg77xd1+1rs52aIwbb6V+Lj+LDQ
GupgMoYHiQx/cQ83UMMI5iU3CBbaXzp+q6Ag2AAJLai04FHGLa5E50HTSS9dxm6i
wL3MvejtnKfK3kIXz6BTZMWH6PwCoVu6zoxFcmUaoAkFdi4/CRjps/MjIoE6APNm
F/637kjUcWP/hvvUr0zlmVtGRYlbjoBRDGcCSXKkb1Drf2W52PFyiuY3uiJqukNF
mOH3QSD/o4ZKcZXzXAq9y2bYaM1x2sWCqPmWoIlC97agnpHoanvUM5wgss4hIVRD
3mlrZXAxhRAhMGkOWeYk/w5aNDf1tY/yK+cT26kupPqQtKwHL+QIrITMas7wRafG
oPX9iDekc3m281Hied7zONsMWaqcKj11pRR5XaGTwhr8MNhWXfvwNgTyNA+n8HA0
hqGo92Cy3te28TmDO7tTwZ2Rz++nqJZfmdCY5t6i/fwcJnuViz6E9gX11sl7/F9+
wPVqgvm/mpy2dV/nNegu4dcaqW/WeHgmCai7pD8NsjccIqunj4LCbhtz24pweKXJ
R8sqH+5yiDg2FvGLcnxDx1XDuNxmoPF0VGpZQC7YzeHV4GtWV1/lTfVJ8iW8eGgZ
wT2rTYBReiuYcw9XKVTKr+t/oVWiNe9CpIqL3Ikr++DBCreaS64iNbuvfq0zYRri
WeXmrlprdBsl0Rs/xZOGbWDeog2fJx5r2h0icqBYUQpvu/z+1181j4taoq6gwf/S
pmDwDuoEe5sJ1b61f7VypaSHysHulXUNgxgl0GPLUdVx+NjJrYaGKF9qerg8TFjy
ogPJmUQSKvJ2Ar5W2cAVJWUPzGoXabJohqbfch1mmo6Iux+IiSBkd8qbHtONG6Pu
SUIAEQ42r2eZRkoAxQ+bbxbmxWmF4zISiINz2Fq0+MLfJnji/wcgcSs1BGk857bx
Ky26wRTcNEwRdjZWF6KSRQxQb6fvOLCVId/Bl+e2Rniv2+14PuIIqHP59YpatytS
ONh3ov2k+4mUY/B1sXjPMAAroIgCQ+KOTff7JNock6vrSCeiE6ueQtCucOc6kPxe
zttQfpj5OMbKNJOxwDt8vSLizzO09NlDVm2QRHpDxBxUF0g3PbE311Exo2iwQbjN
PG+9o71uoyyp2qxlw60nxUMmSyARyntF8gJBz+yvpLlCyIlFbgKG8amyMcFECPeT
bldQYH42a2RYyZnTgpVoBvVzDOs+TWK0FGcORd8sjuIYVpYC+fApHWAXZm3sE0Nl
d51JbOIveTuDh7nowIU+gh0wm29TuSchRS4x5ME9NHItHq9STPvZnbq5T55CafuZ
+yv2Q1NTElvbRs4fVI7O/LeKZqNFtYCifonv8sr2PQF1cx2RJxd9ZJ4rOwUcdZO1
zypkiifbKSNAoVg0yZ+MZ3/UR4Nyk3wDUo6XZUr2GrCbgFfxlXdiWS5lx0kWvshB
MQudfp/i3dYY37yIY2rUG03GtS9+8oZwWftNGmYA6ABZb3SSbJt1z/LpYCSz5CxG
h7dpAE8YQVkq2SrDjIDmwGg0RfYzAk4GFMEFWcl1m0b9KZjpzMGpULDJIpgkEftc
/QAGA1W2W4G/gJuz6JyfgfY8k3Y9zcEFeKUKEkOrLzftlNPM5shbUFvd8tWLa/zI
XUj0pr+0Fgm5zvvweIlAZ+cZG1I40wbuavN4hOHjtxoA95vD+I2hxqm3rjDdI7gn
SWROu/7NegC9/zqMVFx97qoeSnY/CInC8bkWtypxGOAh7AoIeVNmT3iEQuWKWoSD
1mneyWZZ+x0gc/tw1OEAVGp4Q9j/crI3zAiSq19tanU5TYHjkCxix9K7eoZXSSWA
zd1IwTC9wWkiRXQNn646cpcpweEwCW1pixeNj+r4LAwbfsAnK9LSm9xW4BC1WOBC
2dNS64SPdTpl2KLY/eYwXGvMxdC02wpU6goNHK7lqxbhru9ZA89MOt4AL+/w5CVQ
LPCEdX6tvMBHtETbdBnn9t7HFcd9lxfGaK29bbgQI4hnnOXU4Rm+eCIxF5IqDLwf
dQGvlQp26jOzEqHpilQVf92zs/LaZsZ2oo81aMMvuhI1RLUNstvn3pbwgMHAmWZ6
gBH00vaFCIY2zeu1iGCnR2jLkabuRzvCRH0mk83GJ6cpqrgM4S1ANZHysSIBRfey
rXQZy72Uw9XQt8nL7X7SJ7KhfKTJTEzAVg5hN6gAUoibZgxpQVB7AuO7Hyj9+nsD
F+6+ab03IowC3MhAFO0oTxRgswx4L2NGdeXlPwgVqjPgP8cmMJwMHMu1XgVl86cO
GRMBuRhq1Pieph4XmzamO8paqkMekchGHCmKslxy/IxUlF785+va7S1JjT3h1mJG
a605wHg+zSWQwMqztNkhCiVkUAV14IiL/rTCr32Gs/57bGyUC6J9JI8728xucEKQ
liZJEnw/822zs2cvZMbbUVWHd8OXwVWaD+G6OmNW9c3ILtol+Ps5YyCBv98Wcpd8
uw1ZOK7gWOtyzqrHI/RHrMISlSo27VvVs9wLNQo1u+A9TycVtkKEgStUE417sXNZ
izhyOdGbNEIGI1vs6o/KwCcKURbnYNg9DZOv7hqdhjujtf9754k7U8yG04DWXV2q
VE15iq4D3osL4QKYcwTyEHJQGHQkBafcEfiskh/iXASTnxMZs9JWm7ONqiOEnjQu
14jeteWD+TzMbQMmmwykXpeNXpKyBuTtYKGmX82T0qjRjquUYvP+Lewu55Y9oqcL
Eiju4UE4XSY8zURRNU3aD3IJsNCi+h7fE2p/lppbGBXBC67ZIi60fiqdUXM59zSs
F9QzaJPSGhXlTKMyGVIPt7KD8v83mFdJmRvAsGJ0mxYk31Bos/+OnQn6YItJ2l+m
dP0nXEsB2fY8hFemKIoR0R83aYiJ0z+aVl2r5MnjDYayQo1LJJHDGEglqywKh/ez
jjS2K12ECIoaDsPQtNraS4jD5IEMMW3DR1adwAY7+fz8bEzHo2TcofDycrZnEH3R
X44MItLrhRYw9QUBOVFnyRVSV3mh1K9/iQjw1jYdCuJqzoE8WXEbNVfjmWsy0qqs
3Va/8ykASbJGp0XRsYrQDYwmQSXxyAyJESc91Lsm+gcGO9kGp2ELyfVjlC63qPYe
x5Pa7nVZjYfoBexeI8CGwOl8yVNPFWHVtaGmvvr3xiIx4wCwyqOWz/a2sqRwqAaX
lB2fdXceckzLRlg3sIMvb4aETs1Dp7S0bdutIr9juv3WagpcJT8n8FH23LUTKTEV
Qfpw92Vc4rlAAmVC45Pvbj0+Fc2qF7nwu/ZryBuiMa9kiGRqIVJvskDtvaiQbA3w
4Weya83hWSFdvxQAwlB2hmBgKJjPKER9tVixRZGD84ThBkBy5fXZD4ocf/9Z2EjL
6rmSi4Vfz75XQfEgVU4p0RhhO6u8yg1523/YyQPQ1kZRuyvbJtJSvV1J/ut+XBUC
WKkhnWYkP+EzQLrxm5humDw9VHQbeMCYNRCwl7URXVyfjcUXKwDYBMoFx3Sy0+XR
yQkPUyj1RVk2qPep95WDkA4jaG2sI6GGc4xqjrOVSQLWiFMlhi6qeT/mU+6Jf5+B
nrTGOphe95dJu0VoDBAJSFRW3JsN4U7XDb0E5VqzPgpLxZsYipKA8P30RxxVkDM3
j1WCvU0+hIBubRrpN7cl65ABTobNuvH3GtGptObgrI6Q+NW5+yHkmWqM9ZUEiFlB
Oii1SRKdjDWXawYX8iJfqocK/zeYhQhrl0LZwOXBy0XXym9pg9r/J7DutuNliod5
vhXyFQTn/A10EWzskqlhwFEdzbLjYKzAQGnD7OvdvpLyDkgJKDjh3N4ezUkUnyGK
hQiwZGS4brtjTrdxyJs2bIJCkDpd4+TP32vJKwZ5yP/c6yxJhgclnnTAHPD/8XO+
GSL6Ha8jr+cAsZw7NMpOPOy2vE5d0RsuD9Y95OKOfeQ0mWdRrh7T4A/Jp7yaPXWs
8TrIX1jZ+mEtys394JD/9LriM9Q0kJquAhZ7HPgMhTZQ4xbDxNhcIiVrLHVM/Lyh
PFNaeFc3IcWuXKQ6eeWfIB8ULKFhwgt52DwE7JeoLgsr2Pjhj7ELossYo1MYty9n
KbGIeFCoovCkucYeXJYWvV45lnDFNGHlUSraoU/jvVnZ9Hx/c7vYHRdc1vd+OVWN
zzoGrTzCVMJbeRvH3eLOaaWqW3jckUwX2yihoXUOtuyVrzsNBm0sHmwvZt3PAjHP
4sgXmglQtIiezyn3TkY6yAwLcG6n1VOqomPYmqzn2sZm7wFGnSvZ+u5ydH2srXrt
ANxdH/2vJyMPYMpmw+fqPd5JAC66TTb6bQmUWw8xKUheqHIQhT9oOutp0gXGkaej
WtOduSv3uNfDTbJIIlY2TcSI0JTfhkylDUfyAUP673hsqbuWZfjzBpRQu6KlLJYl
Tn5PoiC9O62kf/RWoMOlikQyiT+lOccPdQXH3sRVa/rusmMJFEDnFs3TFqespbZk
vnJ8LiaVgQsS4vkQ8Dr3zYlrJwwBXqXjQMmGtKKw/VamSbBi+XCBm8n1svUkMf3D
ZxouiVuOr6Z/EKotH2qm5GOqWj//54d0CFG1BeclHpDW+Ue9q88oG7soixfIXDue
dpUDNAj9Hve5rQdWUhNu0Bphlgba/LEmBJv6JYCmp2XLwVAcY0bSndYMYC4kSUij
KXo4PM0sjo4Uyx6o9+ekNXnON3RlR5z83CbzsHooM+7MGUDCU6Hc5wsKItGIwm1n
QkD4hr5UwUuSgn1531W0y0Qqx+YtGTAyHiz0O5y14aA08cIEMA6UKZ4yzj+74Jrz
0f6Kqe0+U2ozJk2PQYv6u097tFYsJw8cvgRwxWWvCvf09ojZ+Mi/uBDH6C+sHghR
B1Gp02HDs2XQBYauJyLgxRe9E9AqKtmPI5UNp4mptYsu1uiz6YBZVVT8LIfa+51g
WQF+ztSGdJEapoltgi0XNRYaoNgZBj3uZcvHb9kN11Z6sEVPnMQOn9VWmkW345+a
yR691jP94dVmDH1iWnJkdgDxVfvdke/4wwiCUAKqrnKll3kMd9TOSdO8sMYCSGe+
oyXGcxunQLKAZQUic5Ry5jL9+EhpqSB1UXftyUKO39it3QRYhEYCcgyXdAcSLX86
4tRDYBIjD3mE9moBr/F3N4L3e0VVLfgzvRZwfBQzYPiUi3y2ofhj8ZT7CUWr4D1Q
H8ISxEtee8By7I5OqPL8OrE/zdZ2jPnZqkoSwJbEenKMp11tvRkmvJrafIbe/rO4
n/F10zfgL8aFfdjQHYy1yDef/cceloMbd7q8c7KESiNs15CkBarkrAK/rC2mmd9+
5D2DRuJlcQEBPCOyb1u/klGHgc9sEeDq5VIdRxVVB3mhwjYZ6FDvxtThX5f8RIqA
7Gm34Fva01D8nU05pZBoHQYskewvbhHCU85CVDY+lGZ+TKBAfNXSkuv4StPqIrrt
X4BvqCuWZK3DQvMUxA9iXkNzxdhyd2r0ojvAooerRShL9NjHiSuWaIvNlL+tCnpr
B80FsbK7E8wc4X0oQ7Uwi0xpI/9UFgEMU9Hyr5iE9osl/3r43oVGs1KO7vYaww/H
hKfKm2NrwLeND9Sj3WrqJT065Lhh4+ST37dc8gvryLfpxnnLEWu5F+9AY4uU4U2T
XjGO/AIvLwEgrryC1DTfC/gYdbeh6mcFieBnM5a/6g4Iic1l667gONWdtIkSnNom
8rmJLIssdw3bowPI/PRfgwHhbyY/xYMKZQ9I4xG8d/bfVrZou/HjMXfu998ElIos
/H1hB2Udwytlb82ZVvExoBnRKpXnbnkToMsRlUEe47TjUvL6RsI5fq+iMArcz7Ld
CqxgbvqmjmZxjipUmieKRur4mAJjRE7WhBVczWBGXYpIHfnJjlTB5wQzhXUeU8B9
PruDFf8A0PkLjmRnubZnS7kW1R5RwEj6EjtWQ939M6xmdZP4cmIcm0+DiviANPQ1
cu3TaRYU3vxptfxbgdzTervH3eYJZ5kREGpeJhOJSH0JM6txBNPhCJp9dugdQu0J
a4t0zPDlevS/n+m4Syb2TfzfDLGjhphURSTXdlRjyPAF8lSHxITvxaNL2qKShtn1
Yk/4rZ5CQukaBjQqHuX3b53j+pOkNAGT/cbK6fIzF72pXsHqcx1GROkI0bC5Kreg
TfcPq1rABMtk0yGFdAshKYcaToN6H1lgEU9XcGA9FpYb8U0j36FrURI35aHb58vo
bRWRKYA7uVqTcGCu5peInjNfWYXTqgsaWFUCt7zigKVu2sLiCxbcEkpTfv7oTNpF
FILTKj9w9JnYxoPKyNK0qtgvRkGxz4UqPiLMYS/kHksWvs14Jjn9ZWBJv75KbFLU
p+pZvSdnXww+oWN+7onqfgtfZRJdQuOanNzT9OjZr0N0ScLymLjJcJ9fxt40ee2n
pazJYeQNDIa6UOJCO3BRAXal8cuoJixks5JSXA64snU3TUihHcazW015u0icL2LP
GF5jklKrVa6K5Em2Z3RtoKH+/CSAmNk2/1uFONXFIN2050UFChk78/OeYZ4QZ6Et
5ew3VvIWVtXuk6E96IIe1kTcN1lCio/rZubj4VQjQ2CmmriLW5BjZ6440XeGUKNb
kfP1zHSzGSqujIzpVDELn8+6uLhWy6EAatfkkdUpxrlwJDnChC9Irg4vN7L388Uk
/8MfarvggPSgET8P8Yid1FrZg5FL3eYjWZFBZ9Z/H30ps4WKmlfMX5ybreULDZQs
AQ92n3juL2P+1TkMgWAm2+Ut56nHb9c5w4as0bPWpNC2DiMcust5V1SI56q+m/OD
XwRkjH61pOZMTuaFg+SHwrSF4Y2Fmv9p6fl2Xi8zOmNkiF3P6OAYc03DBeinPO14
XPGp7tT6uNb/SmAqV/Frt6VO0wQqaa3+PsnWEFJiwDdtBxkiPBenKTcj/KC9E5be
Kg5qmz2WikPN3Wu2SgagcngmLjrfSPWpV8ahSD5EmO0rnDwmE4lbYVetVG7nxWGo
r0yKlu+2vaT/OwfIha0qSM3+d1PmOz+nLJhFQSsXStXJqCrIj2Pqs0wNPglLGcat
taP6GY+rO+KzNa/j6KXdR2tip/o5U6eXwEB7vNn2cgU7mxB7uz576tuvX8MOnI+h
BxwRl5pRNj35wCJYYVeDvaA4ijcSf0/mQ8mCdqKpo/rUeL/xyUu5d9ZCM6sqy3Qp
Ix6JcyaJcLUPNNs8xmZFXBUCb3+ZcSxRoM3Vakr4Fo4shLFKmYaWeODWaxEAf1Du
Sj7KEyIgFSvUc8sQcpjmI4mFnCz5C/CTGYDFQ677TH04aqaU8Y8Dxmg8GxZvMm8D
T76boU8HCt8h7kHkwxHfwz1SL5wbqrIJAPFQWpGRqLZCfW5az6mVyGAspP0ooFL+
PgS6cyPej/DdM1TnY29b5ka6IK0e9Z5kqtAoYbkxvytUVSORfTawhXFOJgPF4Ua2
JPxg2YpjciGbC/lg5hurlOhuazSw7jEvSFmXc5bxeBc9sSGO6RiBKyQOLodbe5Nl
Ck4kfU7AcPrc6b5kGyyz4WslFaLVyGX2yXbxQp0lDfcI0X9rZVUPDIwC6Fie0D6x
4BDhRo77lJNcB+2ScTAa6AYQzpwukEG7fnomzI8Mkpz2oMDcsjyGLG37bk+b4Dp6
90+jxtTrVavjFAD0GqOJRldbnMgZtlMSdGzHHJqbENoVQVakKcdt0u8zYTH4B0uT
ZBGZ8HrRo6k93bO13zyIYvEUyDwldnYsYYPj3rarAB1z6hXN4jhfiHovmUHb/wKn
MaXAyd4vEjUYs/kABk8U9fD+rWuOrfoa+8QSNRKWxGjMK0CixhDtaZNfxQGw86Ig
g5hy37vHlNw28FjrHAKrwzYxUQp1MAXGCXl2+CTkhLO0aHCypfAhdnOfZ9lVcesZ
gKLJHQY8n2cNHGlNshLDKEn460o0ywmfip6bXHEM3l/bJ9hxaIH2IuEEjf29yTPt
4flKzpek9dC0yQtKAuvGlk5lnHG/PRG6L1jrq/6BjIKUjOQFMy6T96sx9j8DgVKz
Njb7REjYTkbapArBSh/N++wVzFGdKC9hF/aCHdVaiA4UnS/mBBuhuEi0uVRCaCRE
JV6CevwLNKXFhDAjl9/K4FfThHKn6GUFRva5GgVvi54FMS9s95pKTMt1kblNVeC6
Mj44znppFVwnAT8nB2k9tC4DaSnDkMObMJstcdJ/Rd/k6yszTvE5vAK+1hi2ahJl
TS3sFsJM+jfN3gWtNHqoO8JN+AcLkeR5kQndVCC3tqCIlyRzrKe4opF6/CCBwsri
XjR8EqyW5+7sZFQNtBJ3ELwN5SpTYaPh5VbZCCd8aHOb7Hngl/VAK58UDTujlOs0
vW7ACtg0lLaFjIdGebJKAL8b9pzKzQxU8HBwTyFzTIjJl9y9rzam/ScEoAQ9n8/D
+cCudVOiiLhlvskUhRuKmUBmxKsBShj9OiTYf6tBG5DhRDLobYka311yYD0c0d7z
b6yYknS+x65rZ5por9Coxhc9rwCeYkgvf5eLsWX5grB5xIBuDzPKm8I0K+TRhRMU
lakFEd+tOEHhKDXlSELP+nT61OnX2NIP+I+bi1x0Eme0TiMMmU+0H165ogW1VT/E
p6C3/c+uVGznkkKmFvSZllmpbcsNvqPKHksQEBZfBXHl0225kYK2MEa75JuQaF9j
HbUPSIN8Vw3fNsv7fX+q6yQSlOm6diwpvlTfX+C2SpxvrtFExZdTlDxvtaNrUWmb
mQsiOKlXh9kJZVlWv8hk8HpKVekSINo7pN64NRw0UThq8VYaBkOEQV1kmGG8v+En
9dGXAyLPjeFVbPC7bLjaSbVdg+/VjoIZ3yUtuaoCx4X4K92eD0ww43By+Wt8PBYf
+yfh8hPdbjNrR6FyDIOjIzh32cI9EBrJIYbipickkmZzU+UIcNFhK+/ZY+w/PSJK
UP5nh5GJSAkEG6CADEl+TDDIHnpjOGWt0kp02exT015kpvImgGmA9o1PgwMcMUy0
DlPCEuPZ0NwZM6Opz9cQljK/BQuLxQfsG1YNQGuruGAlFiJfL0UCGVZqI7g7V69E
mhGUpWp5eRiSp7RxBpkdywVA3+BXOl48+plrKh3K+axcZUKeFSZ6h5V0+df6liED
QZV4nwUW+zMuHoh00kcJ1eTSovZd8RpGVkmTdnwGznF148WmS+0MzO/Y8uCw9Hod
jTwQ/1Tc88LzBI7dcIrlQLTliD1BhHW5EVNSGMYBMu3jfE79XtLgQPa5fHNQn5Rd
gxWG8aszajrBYAkmBAonM1WwYO9BAZRWk76blFZ59mGrwYdFWpv7Ib3Y2A+kc5pO
zfwUpHnx2rDuYc2aBKQetu+DsZaiAw9niC0ZLt+rsc1A2KQdaNJmwWcXWwkOtlvG
ayfdGQ+JrERmu6qG4zPlw61rDFwT79gEK8jpyP/OdDUVIgEk+YXsbm5Z0xqcyWxI
TshUepWfMWKM2Bk/S0v2Ktw2uxyXZhxluYn7WT9Yd/R+lc8OmXs2dgiI8uBWeWc5
uqEq64IxWl/GYtxBoAwuVk7IVx2+MfBuRtsatth94YgbFIt4SG9Crxx9r+EpUy2P
QnEsXQKBFND88kyOUENFhWCLZqBi51AwpnRfMv9NJAiAOEwDUTU0E5IWyBsex24R
wBZDN4ZHvzdsTBP5mKLqV7wSV02otud9htvb4oCvmdtYQp2LPefwGxG+zfBrljd5
J3FYH+04NMeZeVBoh2IgXw1WHb+GOPA/4WuucvnJA3GSFkOQdeIN8A8RrZCSkD5O
WEjjVta+fxLqazwq+Mt/CGXCFhQ/xdNm6DcPS7TInRS3mKG3Fh9Tsn9ZrdkmWuXH
KTjoQtVLfzwjD6FdnSAxoLVCo4bWnuKAZZWcpCgS30hU3+y09x+iuDXxkoq45LBT
osV3Y6c8Hl6KZuD5krpAHCXocyJ9q6tRqZGJaKdxX6lTN8CxPoxwUjPl8BSXxpOB
nPYrOjbQjRehhu17+/6XOkl2T7euFOZXXvhvcsyk1cJlwz9uvBXgbmBixw7PV/n4
KXafK2GxzBmBFiiC8RP+dtO9dXq7yUFL+vOc2X8BeukCL0hT6P1DVP+aWaGqdUos
Rl0hMV1IL7t2zMoT5QFoHnee6U3WuELz4WeCpkZ6o7A9Mea16lEuUEcJmoATxRhs
IMugR5xlnV/8tIEifA9bewa3TAHiROXpX+OKEZZvQ9SjmVE+58Z/1x0aWAe6eax3
0CQq+o1Q2uOWQw2GDosiH541RCcKxpPl+VcK4LoZDTMf3zEY9hFPlfrIUNoS3dex
taLg1yL1YyS/+S3o5FVmbpY67tjdU+EhKpJGmI6JMUB7Wbg2rtuuW33zCGMV2cT5
Oai7WOoA9rQ7Rk5j2PfF0pVqEUkv6V7KYEu42cJYw3lYjaVqLKZkVHzqGzY4kubb
+CVXCKbGDra+H02CIlvTX+5XHy+hjxAo4ofZPikz8s+mLDRK4rmz7AgHzCuemq0r
MOuz4MRyOZNDk2hsjUSO7FmUQOsC22iDb0BjH/6YHYnBwAkxPaqbLSIlvfHxpphn
5TwTFQSUzebYtX4L/DjAHHgWMwlvmtsTWA5NAEO5B9MVh8Y9UWM+Wph6djY7QTQG
+DGXj/wJuhW0YcV/OW5u3OfanYBscgIijTtKkLJW24ZOSHlVZRaAsk51Cdeueuyq
z8m2h8iWY6+WcqxJ1dI+YJFok7g63CpRjnu7Ug0d53S+07qSu0rhexb7+A+gmj1G
kWN/e9gmzk14NxN1crttT65rIvkYmAZ26WoBz8cJs9QDhZ4ocHrGGJ3YgaXRrIRx
4JFFyx3NPnIQo2eFOvbXPVP8tUxdnlnTZ1zi1OUWPzTjGUsr2NlI8RHrQmSKtiQm
AbzXchz+yYi0uaMSTXJSvAakWNBHPOfUq0UZn39H2t+RJkZnQ7Krg327BxWBz4uY
iyCN4OyqBI9IbxVX7/1qfc0QIhNSbng5XFrpULkzCxDOVskA0IX+5kLnMqsHiokO
fGtJZIQ6qjtG7dPDY9Deql2OrbI7mXRzqeUAIcY5DAwCFZRsEeDstFsIw6miiOmz
u2yUAA9HKeHCxlRAH1XrY0VMnHGaWE4+3TcV+OsC+MMtd2893ndqE/EYfV+kU+DV
d9GcdpN6z0tfyVFa2fMMrl20YVO4Mt3ubZLZjn1M0mIrje1eQevyOR+W3lPIxRb/
IY+rDDeyYcyDgxQ7fAIScN7BXYPHG3KwfA8SXcVb9NrmxWdZj6VqtzXgH+JH7AdK
wf5DroN1AZjcEq4kbfTBZ79CZFPBCyeOgjjUq2789ytLPXptsyTW4dAkeJs4DBcQ
0xE2irKyKss20SjNSr0w34KzyQWzrxxGJdiP23Tzj5z64rLF17omTwLj5N5TIS5G
jKIHCSLS5qJ5uYUzwTa9yYkntIMV1TD7Yna+i7tLF+XDFdvPzwL1qdbOd5tHVw+q
QEuC4rqSReEmJKQb+gAJySdvtKQ4Y4CdwrnUHwO/oQYpj/lG9YUxPBUD/jWVJQ8S
19fmcLtta2MSjO46O4ATCKGCm5MM9RZ+Q7oHvcVzyOQlVkIt0cDTXLX/h1Uln6jl
FiNUX8zH3MJ1QSK0Brq1ruay6/6JtvuxjzIL6xIe40/SAcBPWo2IkZ+09bpuphN1
npCMYMKpQevyOgh5QCVfbuV+wYGPLF6vUddPZKQ/h4xOzRne1q1aGQIQiLAZfzaG
JLsYyVAlW0XTlGu2ROB0hDfXOYVvy92Ce7YbL75/opfK/+oP4DQ5t19EucqCRo+f
Zs5Inxx8Mha29n0D5Mx9n+4qaBxftSlavL5SAODEg4KzTEpe/um4WbVeinUYN5ju
F20O80pB19SyphtxfMLsqFwuQCaBvBDMM0na0AeqwP5BmKyGSDouYHmS/OgjxvoZ
54f0QTOx1XS+/1xL0p87BRK/X0W3t4OLD1VMhAOXs0mcXn0a6gcpZWBPoB1FcGno
rggKLDjnfrdcd/MzyGJ61IIfyD8cO2ba1nfYHcoQI81o7jUKYYabh/qNa4xmD+pR
fDbkW4/ENnSGojrm/EsO/uaFtjbrrb/LPsskyz81ahrEZsNDQTh1ezxhcXIBCEqa
/KA+58/97mV47P3GBd2T9C5vFGIRZ6qcOMvRiTqh1J3O31ExrApiTlxTNUJGRTw2
DDcSSPShYARsFpWfBNDWqjxDDTOtAEtIk3gU1kfcgV6WAeC6VHoNAd7KN418TywJ
nWh0npK6tmYiauEqQQYWg0Kwyj82ntmeMSQTvjXcPwOfzVZBpzExrw6cOijc34bu
t/dTMcSigjHAvPUSO3tOC1InUGP2bnJ/wOgBtTfC3Sdx+RbHk0VL0o5aLiG6VlBH
Pwitze1YcKGTaJ6LCHekLHbYmA3iE5GzkpkEon9escg2SmCsOUEio4fpoRLnM5Jg
WR4O9t8oXu6LkEuHixyFYx5vsEDDgDUnuctJ2C1CDsDUGGFkoe217Li7MS0b2Gvm
CieCtkReuHYGlVqlgIKccmuXyXMizg20677eOI1Th5JshsCyROmYM1FAejLClNlR
lY8aWgX30qN1oIkKa+oAHDnVcWMHPpjYV0+hda8qUj8PljukPmYp0GJNJkOh/Vj9
LrB1Z+kNjbTCbCNivOBAdMKQfU3iKTgHFMdzPqsn7dMacUmPjQnAzFtDCk72deZu
XeKCRNFjv9fT1BFEBtLxd5d0rJ9HNE6DqLoXv1aWykVvlgVxBqSOstnuNhKAf0wg
gmTZKMHtx64eYX8Ntj5D6xKCh9y60+YNmzB32Nn71Cnf46Z0sBpixcEbIbBmRmK0
27WHuY4+4JzkrJlhyEcYAfXzdz9VVxoLjklS0RkkeVjtcCVxiHNeHEYObg+YRuTT
HTDyJVv7RpQP7h1S+IN4BRiIQ7vFy1ZrF+9p0A2lcESl0xpPUtOuHL12A0U/GhQS
DrBiOX0Z7rcEh/9xIzGK+htwYKlzyFvW8mfFXJr1OK8SW8M8d2bXX9ANRVaqLtiT
I1FmUy36myobZylzM9yZ19tTd/Nnit/PbcOj1mbhZedGk+rKcwAY578DnDTz0Jxa
kzAbYTOIRBFuAvIYXj25Jq0YoWoo81ROvxPoblFJodajGAAHEyGPR0GsLITqjCKe
UsZYrcFS/ckS560Yxt0Y8BD16hJNQWj8z5Gasgh3gUNqCAx8cLRhU6lEFsgQWgjc
oCeNDU1lEb8OtMN7mL2z8RKTMXPYX+59GQ0ehX0WuLv+DfzFv/r9FU6VfgaoffVa
9sOOmxtPVjRS4vtK/N7tpqzm9SCq3j85tLTLxod6ZKryDq9S7xNMPqaDa/shyG8Z
dWfuJSduR3OSWyvvi/1rPMqFAyo6aqtRBBl+4cQghuTnY6ItPRBe2zXaN1cWocU2
IO8iahbOk/4mxj8HS74fCluN9cyW1indL+kNHpDEJziS4WtVA3UXObojwM3rbR10
+no/YZoeIQkWcfHkjkYT7UH7fVZoZKJmqXIyx4sSZxFOMSmQz+wNLeib4XSLby5c
QyiBWRNMhg/vCgj8TReqO6aVCiYswCA2myB0bDwR85wcWn1FdObv1dU5q7aUFoVQ
e4/waq5hw4IPyRqpIqJ33GLX7bdZMadWJQxHE/5KweuOVHxVxNqruC5/bV28+Tz9
D2P65KIprEGv0e7gdbGNmXr5JVELSKdML3vyDMocYB2lB6jXz/iT7dbtQk4oyEWv
AFx4VdEcZcko4s+Ym9Irw+Cex7Nt+QOTcj/ho2ioNNVazti5Q1jV/CGCJBIz2PRG
uNgMR+lBSzLnM7EF/lmc0KXhyQmVplggQajjhVCeNS3avwlgal/GtA7jbHSoMhGW
xF4o2auYsLweVHC29C+TYVo7Q7+XVPFD2d2EFiVH3kgjvZk3rgAl5LKfN9H83Ehn
ybjRqfArGGXzcFUiIRQtRCindVoWgQY+7ZwJ0/Q3T9UzW7e0KM7R4XNsdixchBVD
ugXLyYOQLqsp7UYKvjRWnwE4vKhmAJKpM64DkF3UdbZXf0B9OCS131p/qzz8nAtX
daXjMa0+j8/xP2oTWHM2JvVeAoFA7RyFlBX/2w2+MTNtAfn948M8Aw7g8Mi0fhrK
ZFDDikR5FKGyUBEz42YMx5iBtKdH9nFpvlX38ZWBop3rGubYN9UuR4sAM+6ev/t8
YPcUmvdxjcuiSrH68DjNIxCu91c4E0Or0CddkCnVGzDVUMgeKh2bYgdZGQqOCvkf
NfSpwBIamIY9fsNYSHcQ6r8487bbVDPwPWk12J0iMqf0t8q0hzTmoVXk7R40RPcD
GFLtNGlGvhoEOCzTpFhluNHy/tmvU3JEtIbSd4N2Y28oYXyZQAl75UfK9/jKA+gC
jWEp8mKEesRLltqHiF1BG0sPCo2rf4flTwhR55NkWWV+vw+I/qNTCgKopLMmjnek
sH9j7DcI/M2XlU0Po98Q8SX1PtkQcR1CUpplPiAykoE70TFsaWHKpeeamw7BwTn+
LYxs4fWSBZfMXQNwPI8f1aE/T1mjGYmrvq793QYguujaxjEDceqZuWKI0cCytfdd
CjIHhAf6Gso6om1dFxRdhPPw8ReThVu/L21FvGc18khS3xtoyTBXg97WEwqtTQlX
LMsKTGgW8JrjvqjzOX4LjLHRtkInQGTMj19odPB9PLG2vwmSTW17VlTX4iEk8F3I
G3cqZ9ofQrhE5nGD/2dwQP6Mmyy9TTE8eR/5/ScnK6jDXUjT9x61sUGx5Ex4YW7D
n3KTi63Amzwe31bYj/H8Zm5JyIIgZ9irCEntIpK71wZzWPXP8yvrTb5Vj/bPnsho
6sg+1w9e7HBfGIm2emNEi019MNvvqeuJA4Cu9wlkQ50z/EztBrOcdMEppOrNjj4j
sneiGZWxr4e+j8nY+GTiqCQFmNAHrUsKBCSQUajJ2UtUMPzDvvaL2nSSuJZsfElM
mJEmWjVNOniF0gMa0qQfMx0nPwxmdvep+1T7QWJGlv3FPM06tWnbhb/dpAgOWI48
zqvJER1mtVbQuusq3iRjwiMU9tYmOOW9b1ZD/IXCa+OXVGV0D3IcUGS1DoqiNZ8i
BcOBMOg2Qknx89o9Wb7trvrQIVDTcFWhjWnnUGX9PeBMOhqJFbNuEUAuYdZuSzPL
+gC9M4/lRECfSqDag+erSW9f4lOpLv/DUVWMqyLo8ugr8nY2bPyzTs9/pZzm95nT
N5+Ozz9Y/qCMEhqjYatNu4xE4jQcIA5t4NJZJ4Ol0+PK+EPegUerQ2JxVNnXxzT1
FnRBzXosUVau0wa9iMWOz9Fhzao8loZGwmWMvfSy162hWdhrtzv+s4wDguGpkkBZ
wNlxrX+EpWIRsB4+79wWU3SbrjlYIX/zKEKAi6h2tjlBOZ1McDTBI+RAd0PTohGS
ixvkllFqVgnREn21Tuyo+Ea8QfNhFiZmC1Ze+Q0EMYoVwujYKPUOgxRWjuj1uQly
gcLK3m5sPf0dzbhVJjSQPI6UAPJu72RD8Xi8eaJzRbAiauDYTAB9O5rtd9D4bogh
mn+62XXSlj+8ZSrSIqvWKwB7UV0+Dm8qb3PtVNHTMFl6kGwQSvjlZVlIoXeIKL6M
+oLVF4QM6PcKwchwFg1tUwI3f4VBQvqc0R7Jl4CHh9SBTkhaVpslvXfMpdmpSDfL
ikTRRR1FhpVsnh7KCjg2/31omMxDFGNqL/YduBB8WIZDmm4zS5Fkn+LUn0buiioN
QqvyoDeLGi47dwmxslYwf3rIKxZTI1HR7hzbCQ2kfbRJKdffo2no4ITED/Q6mMDr
yg7Y8+tA8mjfwB4a4ESrIXryAPG72ZXmJvPafByuK4/ABRGGkjinQ2AjYX368Dxg
fvonFbJuX/h/JMYpABcHG+iEY6S0VmcuFR+KwclIsLMJe2M0X3vPLOBlPT5IjKY8
MnBc8aDHyQjoNW80iSRzAtrFmLZKnfsm36hApkf70GOcL8uF1co4SsN7EJiqstfn
nHCW9wX4RA25Zr43lcPDPNxIKOT64HPWsTuJcbRUqt5D9LaOVPiYKjP1hZ39Pzuu
BFmDjgfZgOlm/6rlvQm7ACOgTVK57j6vaU/RKHLJtqz0JLCbtSvNdDeVV8KGx3dA
kCo4n8SQ6qLWDvvkvxTNWdKsXFQapjgmJLYUROHlv7uoMkkEwixHw6ejhb+GcNcX
fOWLL95Or8W1HfmqSzycHd3LngayYHRguoVg56wevzxLFwX02cf7Xq9IkfzvtIBq
fPDPYKkzzVl/rgBOiwsAJfU1Ij878IyaMVBxLF5hO/wTX51BldTR68SCfBhe9aqm
HsHV1zFgQOzd3J+i+2GHQpCvcpCVvr6kO0cYbYgt/icKCF7438WpFqzcKoJrV7CR
GAbo2v+suzMQ3M61YSy2YOSeyVA2mBNRYjv/8uPwnv8jsWtxwuF5/34x1y3IExG7
Pifhz+zLnKvx88qD5Ua1gH/+pEa5twjDZsBAzfmxGkISV6dfV++VlrdKJlpCS7PF
ypyVcujjzcQbLD4v5mlM1JrcN7LrJRfAuk51XxaGlEutbdG3AkS46LDfjEUll/n/
ieVWvmOW/xtExH0QqZaLtRnmlD9+2TZmSVEsgeab2BYsxKVofLPMskbrZLlobjIE
knNJpPRzProBPj1eU1kqFRtiKaWAH+4yeUCn7o132rEitu0XLg1obAO2V4KZrDf3
lcWKk/oQpTJYFZPXPjmAhUlCkgksDHv/BAAMUUL27Vi8Rkju6ZF4+YDPtox/HwHM
hiLdbs4hmZ0l5/uWSy2Eicd/gY51jTokFOEnSfWaoDKhTb2RDbiMvW4J3KrNRCda
u/nr0EWYljBgi4y2kgdBV8dzzo1OnJCsVRVFPJfGK1DNFxrEnJI+IYRNgI8lfCGk
Fy+bOJqt9jR18qJVwmQ/pvTGma/sV/pTT75Jb3zrAcL4AQ1UKIutsbm+16BMkRtM
1wqt/al/KWY8ruODFs2Q9uKajlhWgc5/R5jaOmnkJswkGyl0Ivi+0MkdVYuZbkhR
DG2UoZImBJ2VY9nDTz2v7+OQvLcoA+f+fowHgfUw+LKTEQWOkDe3ZxDqgMDtI3a2
jNdPyoJARvdeJVljoI4tC0/jqY/1GRvdQYpjpRH1jon7ZwtmluBRVrOSAx7J7lMy
7M0AHZMp2QsohyLtyP0gb5pO2jvVrwEcLx6/2A6f4yRknPCLWPnjVndyqm9IBrsE
Z1Qsg2nufKqx1mei5RusvY3ioefbHbPSdram+czzGISh0YtUSrfXWglhw1w7YBOS
Qmb/TmERKI0VieqAb/agkt/4XdQmRieUBnQZuGrj5wa/wPjbCBm+S6QWWspJbSD1
hIJ+RxK6FWsR/WKS3xylKOTdWHMFqCmYPfXBFsM6nV+Qq5CMy3jOIMlkdjhQ90RN
zFuqAMrRN337gAOI7yD65f/al9DJf7AzIg+QLu6kGe8jeB4jYJKRfRAqoyvt9/hu
I6zRyFoySVMF79k5ec5RmU2cGJt+uqQRRzyjQS/ty6LDCaGzNbIqaTJZs1rvCdkd
yhzjLK1gP536Pb1HMIhXW52F4vzbCTRGgcOQJkIEXYFUuSg8+hSJXP7afCl/HbCS
BlHEMc1T95ZKBLXCqBGZom6WjM+rU8p9dNKP8gJ7SpdZfcxJu1NZ1kkjiIccavYm
F3zrToX8v+GwxuORb506Rnw8ntQc4XbmAY5GiM9t0i42iYi0Ob6kNw4Oa5YJyi4a
pM4DwmPwHvq1Al//wbqlbFevBDWWL5SXcLtZ1nTpSfzr3uUr9KElwItjptM+jqSH
Yb0NBH4yqYr3Xyk/eqIloBRD+UO8H59/KYZR51eK5FBqsY048/G8WQTFemSdlf03
jxY3Jef67jGSeBQ049LGeU03yNknnNG5lDu9oj1cp04IKtkdOC82WjnT6I3LUxxG
PsxATys0o1kpwon8Ss2E48923BpvFUMbHzm7ucdEVSQEm/+QbXedX0L2rJU8Usq8
qeRra83jT3/JpUnY6FgMzHanb/3lX7gc4IdsVOr+F5LK8NOjbEnQJ0U5eqKh/o9N
SRuesoKr/TGW0l25XIfCEnLVbB+nmDodhNe1SpZDKHLTPRt+PogGBL6EtohQc9c9
8QwiBEqGil7vLn/6/1iQp1x8Rl0F8G8/eBoHfYxcTc5wGQkHFIc0eWdmEoohpBiY
OVIaFoiq4t2BZ/LWTwfX8KsUYcKjLyh+7wNxQX4G6BXZwaaUpAPZn/5BvkqoldF1
GmIXwmjlkdIeUCTFg6QOuOIIw4ADWA+NKd00g1oTGyZce7D/2yeXbC3H3NvDMXS1
SedjUIVcuuJv2o5QmgaXrcqRz102Fzd79DiIWmwFYhQuPcovqRwlg3BOisYnK+Xz
EjSvFwjB0hpKXYj1FSQIY6ZImLxU8qHcz4QNWrPsT+jLOLS6hqlBDXBy3fRGKj/E
Igbfg3pGgdaEyLrTmkpX6TR9AhK2KRNONUTdxTPGA6NDDxXSaf8ZJaLV3R+B4qcX
xcLEHRKyy3TQRJ/29ETM6hz06ljetJ0i3f9aZ7+6XoItl9sKk9Lq7b/UFkMAQ7bL
1WpZwFYliO7sHDuBOFxQ9YgfUBRu1AMCbsPlXT3uPYIU5JvHJKuJV1tUDO9+txY7
F8YG6NQ+hGRKHOLC5TD01mfoGqJeLvPLIE8o28wDQgL9Nrn+Vvpm56LLKJbG1SOs
v33mp+2tqII2gfbABItvLuAFGmCT6SLUrx++xBf86fSGDy8WsmEVY2ZFL093jYVr
Qw58xiPMvsu1r849ZoUIPJ7BE16u/3qMevg7vPD8oLWRrOmJAlfYUT3wxhhfUGX7
NFakj1URzsqkIIOW/HwYqIAI7vs7TFAd2MdWZnAmuqYlU9yBfR/R6bQJ8fw8jFQo
3UKR0U7orDhYT7e/x3L15GNN7LZMXF7j3pOWXr6sbB1F5GU+TxL9uR1oGoEqw9yQ
PTCqH+1XlgfAknh/ocIulouZMNSLDrvv0Hv2l7au7BSTBooABvFs9xfUWoekN4zZ
IwequpckTCdv6CSKGRB1BGw2W5Nj4aSIn6GGa2v0djgJBP2voZOpnwnEAEBHu+84
2ZMwG47Zq27Ymu4X52FNwb/MfcfTGHdRgWLkdZCrx0yAPTJagJnBQfBIfbWzzHNx
yq33/65kgsKSR9C8mZ30kE/z5nWiLDyhCYwGNCG152hq50lAT+gGjJX/OmqaaLns
s6ofMJcflzf/Q/Zr/7IDArlkdFZuMjE/5Mu4qD26CZbq/lJefVxIlAZOQyq+i4eW
U/AcqDd/EX0PLrv4j1B0BOH/sp+qVCI24EEP/KusC05sPXtc9HLL2mg/f8x4nAQz
sMJgPdvp1B/Gx6mi0gDTDmXmiwwjEPpp3PhFR/kTFQSte1mXVsNpYZ13VEv2fEFy
EyHG5WmRLIKDMA4y8agfAVsprPeGc//GQOE8X9l6pRZESGXdxRnfm3m6y5nxG0AE
QZ0j3lI27T5HdNHKQgv1PUu/XY7LPzu6VD4eLNRtwKDaUHhHjDI2YdiIXt8vKJ+C
roJ0y2tsHWMs64iOFXldTfeG0XQmqz3omiXvbnw6Y2YvGB1kbUNwNELMtPg7/YDN
SIu2WBEcWP3xKYZQ1iNPLRDIsvTaboHZPvGwVGstQt5N8nSmZqj0n9UXXK7lbURd
FiKdjFHix3YZxUZemYkXsY8dnBC/0CWn3nxyCOTECbRmyVIjHBtYDvwlFtnPDXCc
zk2Tvd3nFn3kA8m24S9HeLyE5DPPy7TOCLXUnhr8MDU0JC80S+gMsCRXwZcIgGhj
9CHXmHangkShMGXj8g27Gk098JSHM0RdbrpvVR4symJfsKOVnHrK2eZgdfOfsx+n
pNuSQiBwHUpKCOOF/vCLmDsxqP6H53L5UQ5xjmS6ayo/28gT6qMWfdCpxrouD3zj
DK+J4Sb02MWt0IYcalX54OkHfzYygJxN9nO5ByOf8R41s46Y+7efxyVaJ+Qz6D/F
CVzLR4f5WC2fp3WHh3wuYqO2z2UjIjWxR3s1nJ7xkLIGAIbkedvBz2In9dVpHC8r
S2xsGaMy7eQS5G/GmdzbjgQiXuerv5f7Vdf1lvcLmd3wgl1Vfc4XHxZyv4tgeMwP
P1LXzPnQavk76brO3Uip7aXzpW1vDr4DwQB/3f3i/rVjokuSxdLppmf0iM9jeSv+
Ljg7Pu345MMDBdUov3M1iZxGN2aHSMRuvZTHZrwKILMDEiTLnCoXinBUIAReg8h7
qNsHwO/KQ/rtWQpPHHQmu5/l94ONRidxp+ZtDG+9S3qJe0Yew3oeMumsitthRS5k
htqkxHi7KDbA+nLOK15Yldn70jnXl+dHVMrhIhVOYkxpjEX8qEtrr/aj5e2NANVd
qye6D9WGvzN9qWXldptBGKOoOXr2/8iwm6x20W6BGt1x68tNLyqaxUcMH1D8/Wbq
vJ87nmgxM5ED2XFqzmawpzW5VcgWC14jFj2Qa5J8bPsPtQpl/uXPwLeLIbVzl9HW
G0OaMV/st0+qJhLCjvd+nQmMFGCjILYKZFznC8krxtqAczoxJY7MNg5m0BRIFaOA
r1+RbS4EZI3NPIsn+3mbY6+CbO01BUNZPiZeRBfUdQldLYBs3OLAvKPXNtI/ulYf
CeNaTyl/D6gQiYDmCngJ27ASV2p8PsoIIiFU4uAYQmHSW3V4JmqJ5IBAwitY7HgO
KHGp6EpQdGTootITjtETs6F4QSwANgD5LXkOkQ6FpAjluyegXXdq23Y4ltPqPqXd
TIsF6Jp7CCWGugHjSAxnW9uJzooUwtubJ76MvbFyWdtaySx+247dhecTxqzHyv1A
QHZCVtFPg7sBLBPbB8AqZuo1cp9YWSickY0kjFPgQ+5z7fek0nnJ9Pwizfr3RfQ9
lLGS4BDUbi+hm6+6u5GlrHeIkcNteBa/MvXGW/67vZsMXeiOJUz6K4ibjXdUsINT
43ckVgF0/JyGkEUX5OMzMvlZaJFOfbPLPwczOwm225hvSZ36OHJAt+tfnJo6jXEN
GXhxRm8BtFwVf59weljHiKE2irTqtrtSpeDYHry2maiRE41hitt3rl5OdsPpaPgg
YZGA86MhIUM9Flz3AybRlk+LOf87QI0qDNJTNy+V40xPblBwJjx8Cay2JeQ/KAzo
F4akbNIzmmGNeRgnmtuUDGPuVSkRBZldIJgnXJcclrdYdTAGw9mh7SKC18S3A5dl
O8Z4J0bZAhzPwT8ahBINZR7u2bdlV6w4bHn2QJX/2RH5VcdAoa1vBXyfeQ2DkV3i
k1J+UnwEJ8zwvExyQzQ0oGNMzTwFPJ6dEb+hpLFd+ni4vosi6TXiCO08yti+Oeah
HYMhsVYIZQ3qE5OfzsQlJJK/YJMr3uhPORLugTRDt5iUvW6oYWOjw8o2XVSEpUbN
8JF3W4HUKlelnD/bIQzG2o6T9RuSxfcGhQ42yDIK1AlVRM72Tf/ttNUu1VGQzEI/
xEvApbF6GyosBq8O0qPPDoUg+1apRPKAo4+1W4eQuNCzyVVWCCPRG3iqNukFRXZE
QheIL80szl3bIbMcQ3uS/fZKAAmVbILIApzCHT98vpn08NoLbMBHUUXZNLvwUvuO
4LKyK3ZRZf9bEquJ9f9uQsg+cHaS33IlZIGT/OOEHBRX0OQdqFBPbeiXB4oCpHuP
jiv1u1qlXWdpOcjdDbdAaqqYu5aJzlK1hptkwict0LMpoJx0dteuk3C+mODm62Zp
H875+3BcjWFGMlQVMMro7/VHDc0FaAOCb9gNrYMBe+3uAX154YDPIpw4xEtWxIjt
V1uzGlANgx19047KxqAxp5pJ6lpJ/0XoAvIqbUPjS26+8uDOohSSYCBMgCncJ77j
UMsNpK50FWoXf6sDOsC44nXvuBETNVW//srcl+6RnISuDbyn+f8BZQlqS8b65h5+
I6bR6rjqeKRr6o8KbQ4nIN8uVSuRj2QijWl2ML4TmQyXphDKU7EQlGcggiLbgzkK
x/YNcMRehfvu9sfdHoqkd6Kce+LGN4Ygd+v8b47wWyGKCngoUz2j22FBdyBeIsfC
W29SCse006wEEghBlyzJblvuJxjW1slnQX03Wx5jKrZKHeQB8ngzjtVehhS8I2+C
BV6rqAIOUWiy4bgNodoN+oq9kwMa8Yby519oFBMp5OfrdkuxMFxjdmJp6FT7yK9M
f+EczlQM11j7y5F+RzWwTlcW4wipX1AfwW6cneP6x73UfnMh/w64Br6R0hEFtazG
SpfVCExzB62t+wRxMA1H5B21HuZ9h5sd+BG8Bmh1WFQMousv1P8lTbr3eHvjk4rX
mk+lFH78YBUgGI7qN8AuBIKisY5rNsi35cr6kF3TdMKos83mYAvZlh3l7CU7FUX9
9QA4evZ+9ALMkGlCchAS4ModP723R5IyDD2PzCoPexNt9f3MORYtXMOBXKcV9WP2
dJ7/fYuKjpc9DUvItb+lvBhBk6dsbZDn7ayL7yc1b0MyY9qN4cC3D3DsCb/Ml6Gz
RrD/tx4o3frol4OqgIXo2GJc6xqyfugfjHbZ7p+9ayOoV493F7M5veL2OhmW+Rec
dwEmXKHEfbhQMwzKrwV5yF1/AH/mzTs86w6EV1YO+v28P1wvE7kBpKySqq2yw2rl
GTZnRO9NugYxoOFuXzKjdQ/964OW65FV6EGClSVYfppn462t0hNP9sl5zYdt23Bt
heLqbkiRvfUNXKyWM029HUde6aUDvXJI7IQOwjeXfw8orG1C/ZgQKg3dxm1puARL
x4D5PohctoTzOkaDnwLRxxSLeypJErUkC4Q6IZ8FnYuL8jlpelJXf9wf645iCIuM
1ugurD9nplRV6KrT/CVqudMtoHl9L+6IIHAHiu21ZP1YYla+kspqmBTWUA9IPFFp
0TdWPm1nu6Nc1myUDY+VO0A3ZacTBf+ICE8w1vm36iNXl+SnBwoi6jC6JL/BiOdu
RNShMl7OYYYUciFPA36OgWZKQI2qXBS1HHhQDNX2s8sdWAaAZOkFB4WGE6BxoRcA
4v4E1TCwDZHOuNe/denAdDwVTpIpvx1BhE6RgYgO8M6rRFs/+gTCgfM8xbPEpBnk
sqvTa9JYs3B6ti8LC28g1KMA+ssv8eDWKlyGPB9wBJMY+olFl+S6DyQ88hR2X6yN
e7D8ahWgZVWRP3PxaKcdof+k6EWxU6uIuvxkQu2a3zVaI0ll0XrnR34qWlmToNEV
jMEEBjGKBQoF5PwJJmLXa7/puTyP7dc7WIZUZIC6RbTE1zyRr1cuqQHgDR7PSBht
3bxLMJrCB7JZT+px46MJr4rhqR4W+jOsAHu9JJGdLgRHUvkeplYtSvoJhsp+xS9h
xuIVipY7G37XmbACw32pdjJJex6rCAvxYLPtjGqRXJzSmXUov0Rh+K4FOifq0bYD
Uqqwz4b/YpS6ON0Y+LhdYWnky/gKaD0Xs8thhiyjEQwj2J9wPX6tsWIxfmFT6QLF
sNfaM+R950ot5N+9JhV6Usn21Pdl7oiYlozuR5StmdzXmzomse5rxbkyHGVeCAMo
Cqf9Gdb1iTt/y8LV4rAl60+lW8gYK5EndjjKrq90wI2W2SxtGToyPQqCRq2NfcFV
S1jEHNMebo2rRNldkvPOwjA9ubVIdXO5Kqindj+umz2yHyDyxj0y2ASL3bxbEvKb
ZPEgoQHKm7OYd/P1vnj0X8N3bWF3ia4QtQDBOcpum0iXp55OgNmirYgo+slPM4Uh
hc/U0hpbSlkL7ldMwtiNeWOP7WipST6MT9xj5RxUgHNhqQtGmJ9et5rDjcO6H2ne
NiKvYcmSF2bPq2HgeY/X7G0XI8KobAh8IvzYPU/e25DfYUWnyZkI6096ezsmk2Id
VEidZ4XKVb00i/w3BGqFIV9GO7q1osbElHzgfz84cvvhcBXArsPCcs/wd7HF0Os6
fs/leHvvfmxfT89LyzXSwoX0ZrfXbagq/Vg3OgPCxBvrZVhYO3AFzrf7iz4c6EYW
Kg4JuVQi2Ulzw4vz18UgiG7uS4QHSqUspuuT98K0XMSTCL/cC/T0K2QwOr17y/46
nXBwATLY4zqRyBwFFuDkjgC8Iqu7KvWdr/vsMt71UFNIIBNnklSx26Q6bpgUB/PD
UTbqWAjWP6+aIwu/5Ah359rSxZre07OJ86TQonweG290F0tr8Kv3hVIhB6kcbbw2
KaQ03wvDbxlP01zhik22TQE6sEjIDNLTMID7kfsZdz3CwabjXgIN3Do3x/caDwZS
rxsl8erIe30TZUUWlR7Qm9R0t5QUnqE5XB8IYfe2gU+BN0JtgmKD25jmGeGC+BqS
fIuIl0fmiYGjBUroV4J22zKM+wsZkubDEZC1LxOPEJjPvhblqWToE2507IH9oQqk
r3P45visUD/LkKvQ+LJQ8el7XU6DktfCc6PuALwPNYFHKp8aJ1NcBl3XZv7eAqyt
cT0CYI3cAddrYFqrTaP9y4N/fRxNkvz7PccSbmPHjH2/ZgQzYtMlxWeelp97Fy0Z
qjZESbLsJplbN/+wKIIpNlFeP/F4aKA+C1d2dYaVheZr0ntG+siayKrf8vIKfAVo
Bhqm59YIuAoW1WQ0KtQem1SyzZR2d8+tVyX/6ulDRlw5JrjVHkBdihVI0Ia7bS0+
goUFbUvrCS/yfjqBm8Gq3jcMxyEwlP9fF37d3+i8Bn7e1KS6yhy8lAmqoPBYdypC
/e3qKdMJjXf0MNXOHekXvBEP36ciBH5/9J9OLVCLbxbct8bCFy/DB0UD3Xepfdb2
XfZcPCkdZt3uQkklhC6endxCSxo2IEPNUuqNW/eqKUrdyuAEgbL7hkThfQ4Bwth8
g1hc6IMMoWTUCo+BAN4luZZs29fusH4DAZmyMfZrKrTbHVcsehrrBklxIzXxfPVO
TzV2///Nxyk5WfSCZyK8YLVejtsDjfhmbKpBPKYsMIJHiLlNoV5kvYMb5Ddmu490
nLr+Y1PWcaPG/cs5DNfQ4i2/zQvIHKokgbE57nfvv59iHYQ3cMscrrpZ5JnMD3CH
C4OcdEqGEveE20YnVBJem8QPVa+EWJt8PBoItFmBFqphmsRo6//fIhZ24B2V5onH
CidH/Fyw2GGNIRpYw4IUrH+w89B+/cQlqXHVzJrXwnI570cZyoerGU87aanapTPz
N1tWmuC8M1baQOOfjDoqhVINQwBtRrBi+exBqFZdpONs2TMGbm0s22fMfaPW0KEU
Oh4FUpnUiM9bHTGd3BYQwUfVk7exOGz0sScQG89OVvLkU39RpctnXBuYnpLOM5q7
j8GkscEQ5tWOOr+Aq4bjcF5s/cQCsfPjvhW60QkPEtKhgrc2K9thLNi2/tLq55aU
d0q/j8v49NyVLVfgdLnPtdp33lIi5on2/jp2v0Ee7a8gDWaR4Yw9Ac3YPBMWn2xQ
yvzsm8f/Wu+xAElgFcUnrd92npTy16aysd74i1ZdG4Ad4jJAuKRDogBREyTyvAi1
f6Kd7AybZ9iFzRZgRCa34x7Zgvy+Xw6YjkQvudRt/0K5nndP0mQmOc+9OXnL6N10
flRhejS8eVQU/CA0bFmlaY+ZXV8mA2ZSMmFJFo1P5PlBxyAPE3q5wgQbe884fbeR
xP0AndzOyQmZi7B1n99vfGL//FSIgSdLBhuLzc0OFE5m6TGMGGXP//ACAi6U8nBe
PJOfc+AlsOP4qfyVXLy4GhRWeQ9UjPiS3Jt4rXOlyT0GRT2H7U8nmCytp+1Pd8Ap
/AwuhBuFiJssnsBxKVw0bD2xPld5LpwhtTky1ZwoU7/IIGqRjqy4RZwhPNvgYnDT
6YHvEZ+I2Ao36gNT56M+rDowAxF3ZJCWpnwXGQDXvsYRE6ke4Bt87bhg2xYxUWVz
ROGZBPn1uxdPmsnZ+efmvLcIdijdubRvb9jFdkOjECKYMTUFYGCNLhn2qLiPPgBu
LAwGvm+ekbIOHq/XvjykacOR331/1cvPlDuJ0QOavQLhnR5ZBicxBH1GGevmLU+Q
Oll/JWdWscEKhHrHmsr1+iOsFZKsxUKe/0VZ8MP8XcPvfk9HP6I4Fs9ewOqyA8BY
gGqWJBruUQRw05idUufLujLps9bwQgURj5iajHCvR4pp2QQsEtgecuJqyXErj2Yo
0piN24yF3FV/Cr9g5M6tTymq5dB1bt1f18fUV676TBepHvWUwoLdl74GVe4PTULt
nDLay7gquQyPDcnhUhaTjLHty6rPC7xhEz9Bb5uRe5H8qw9VDVD6ezAKSIDyA7DU
5o6pkKjzAr4OqtrOR634FfnpRb7A8PrZY4TnGiSvOnc05RdXrYz+c0RaQDJgzscR
G9vLTgE+iSADT0ueA8uedj9jC1k4dcXRv4LCoxv8IxdnY9O4xNfBvHtUv0rIANMa
kxMow5fd/+PsNlrsdyCPdeTpozx4tAKCBqgWB6XhQ8UiNCMovCUT/XpOYgOA+4tu
ECQTpSMwZPINuwg4wNLqnVhKB1PI/GESsj6W8KqzY8uCwfveRzM5mC3N9SjSzPcT
VXUL0VToL8zgzJLj8TbvoITgxinQTZMiL+jBFdM+XFaHYRviPV5JuDTwEXHTxqz+
qhFcrobHiae0AX39J0KKcggPcsUDzI7yTjJX6O5Mcww+rJxLTlYOie7Kd66TF6Kp
oM3O+JaQ4Y4AmPThH7iKgIVWYWqCOcB4sa+ohmNRi6gOsCDSbIB1QG436orejHLS
mA8jHKTC4P0SSF6tKwhnQuYonkYXef5wRdzfCG+6YIEJr1STDQS5ZTIRwbOnfTLe
sSuSrfdhefixb6XLV0QPlY6vkNJHrbeCJFZe+8Byy+wbH5a69u3HbT65T+2VjoTI
yw9EBlbIUwu/O+Jr3b/v1RYM3PVK5b6c+lV3JYg7uuXnZj6B86oGGhA64aUpnmcv
4eYa5WQ76Dn6U2x1q72GoyguTKAy/C8crwBfeXrEokD/uIE93pqREwP7k7ivczoH
KXhGSgThkGwchPF1tUmSsWI4p8kO0TjQqVGlnNktMKnGxQNuDYz4DBTLLlH8nI1E
vHolPdRKzTXedM3mD4PAArbvnhTJfmQsRoJeJwCE1J/e5jgjYysS2/eVGXihS1fC
0UOauPjU1tlKhlfqnmiIj4zMEPX6xyYRqDrE8P8YOb7btdnaBV4iQTlop5oNJQp6
rZFGjhwYwSDMxV1wWE9Wa2ekeZO4tPPsmRaIh9izgcKxZvo/SpPzZ46FLsRDb1jf
KO/gSVgImY6+d8cOqkqREjgxBcqqwfM4Pp8Fa10qCViGZ6NSM69uO0kIFVp/dqhp
8E9DKT+HVixRUR70Za4Lt384o1LXmbWXmfTDL/NEwbQ9LZSpetJy0+KFtnh0PzqW
nyNVZ3mClL05D0+UJS97GH0BVL2pKRkz+mn1leVbg4EOw5peXYTFviI2xhnwHo6i
yRCY78j+PmjNHfMsSX9Ik/qje5X0BV/o+u8K795ZZJJSgU0tfhYYe1WLXYpE5IsT
F/AMcRQLKFEUxYfxrGbXyf4m9iTYnLJTtt2DL7PGlbiZukLgjwHC3P2oew34eE/y
iwFl0KxK78bTubV621FXvsJEvw6VaJdFDQTS6m8cHzMo5ooTss6t7kp4GBUG5UrC
5DBzFQ6xkwuWJd3r7fJOrE9PJU4fdRQiqiQf7IVmQmcuAGMlSo7DnpVxPzv91SYz
hAivXdfExq4wnBdOOshNuplEJt/1LHkEuaZ4Pq6D1QUD54PlWMYo1k0GdU9dSo+D
C5YNVg62d74a0PykpFV8hlnNxRJv852Ml+nPxBmilZ+2hqVE6N7+vzNIQn8m/fvg
h9SwhP7X/ofrh8YZ/jCOM0TACbQkVB1SskjOvRCtvNqWyRwwsqCQYGih6wVDst1e
Ph1PxvorCsdBIQ/hHGUismRRLxpcD0nT/BDnLuhaH9LNc6RASyLrnc2yGVVxkNTw
iMwVE6MrxF0yML/OP8ZyIXphr5EtfteAeP8bv3GTWO1/gVOUpNeV+08VqIICinvS
+hIgoNN/nkpM4o9swRD+e83w4WOSx3wzZx/6hPxFZgNrrpNsemFqrv90Ap3wnRqI
JFct8pW17XDuevrL80n5OPU8hbgG9xUD77BaYtK146pDg6om3HKhwlv49zQCxAK7
UKSeQrqjRBTol2HYpAQh+9Q/p7fxK5Z/xtEZKAcRuPe4jsZ0dc9hGVge8lbgLEkp
3q305AmgBWIUcj1IXIwWMybHAR+r6I5lNQS/SQp/9LwyxaIvtbWvP6Iwu0cRfve2
812eRjcXNqwlULbNIqRb+ZfMEKPiE2DsE9rtw3AFeYTLxXnifZv77R9und+/3BuH
awTDgUsZ83dwtNuYfgPNnqw5Teg290cMZGaEWoB6r/XKfsa1Z8Rcv0GyRJxaWVoe
azA3Ves4zWEbKU66PaQ8vvCSeiHt63vhEBsVEoFLJNloC1/xmRNYiQj+PnSD3Z1+
YqQD5o5c9RdJo9ABweTaa7QR50xDi82u4KTWKJHfL/J58Dl+pw1471FnzU9BSJCB
zNKReDiXWhqClxbZsAl/VxerghpFr9MB969SiqsRoo+IT2CIMLtDIt9HHiIXX0+V
ylCnNvy/flcFM0tgC0p5579sgeCEeiOx6H2y6D9BJaH4PLrzRI1DBvKnhroqLpmS
Juhrbzz984DBh2drmre40I80u+ZBxcoaZ5eyXVr5SghnAd1O+5RShB35E0Eo1HTN
ZZ5opeqyA2paSQZC6LiH+i7gHhDTlI9bgUf3Fo8KRmMkEGps28G9BuVw9NAG/NEv
2d5FHP/PJvjC4Mr63gGtqkKUXmobMipLjHcZc0btovk3sFNIWaXPfz05JIcX5PdJ
zXCKPb3t3B+cWrY2K/YhCYKeXJ6iO0p+zaGzLoeL1lwAzooin30ZkYoegU/Hk+p8
sv567T058j1kq1SpahNaqLs4a0WxqCCJH34MCCKl2dr2aeoo3S42fbrxH9rn/awe
vnnCV0DpMh1Y2qM6oO3EpfVSKNTmWBOb2WNxQrvLMd7FHOSTy4hMy8tduuYO0woo
6p9QM9qewUQ9FdnYri5DlR0w0RPD2vp3E+CtarLwSCkr60PCcq/A2wJd90OEV942
ZIEKw936U67d1qpzdE83zeDH2EPP93jEa74SBnysbctRXSLCEaOyf3YTILzU0zhV
cvyvRvuTGm1ptIwSjYs2FHdP9kSNYvcFKSJckWDYd7RZaTZrt0Ltb5l3QlPahgRO
5PA7M2R2SBOQrG1ortCLZ7wzyiWfM5dnGJWjagNlveog3TfQsuIeWLrKWd8uoBSk
bbnLgimlJ7d3X98g1pJlrn+5Sie6idjrlijTbSh4QetyH1nXydcCRt1AMd9EhDq6
KNtBANsX0deLmnRAouXViYSnI/uKvSPG17yLXnHCZ2JfrIeG+reX9yy2uIukSLU2
E9PPVtkxuwW53uWEsi6Tqq5Pq5VBxwWMVYS1a0f2Ax/qPOznCpB0epuK24S6Npsx
9vJ0HLhxWpMA+WZfax/I3tYUxD4N1jb7bDIBpH1nkwXrvKrvpgWbL3SXV4JlzjqP
n0kw7ynHfr8DfVE/P8AAqFEjPfKP+uXAPyySeA+/XDNUWa66NN90TK7943HA72gg
e4DISCcjHchZjIsQ0MUxHfFYi331EYd3Q5/VHyw/cTcAxspE14Tw4krySqIKq2DX
geS/1Hm4VC4yh3ZsGvfQn7BYd4XTeuaKhmwJFZ+MngZWoljO0G4a1NPQ9GqIUEkr
ieaBO5dYNY1+XmRI0SUGLLaiudXLXkNRVnr8SbaJGTI/bYNDB2n1H6zThsF3Q/87
FqZPDegv6HS38QZIgyACXj2m5foTtwl9slaIb/e0etSX61JbphyEhhkizaQuz+oc
FiNGNKoXsClbVF38cVl/FyUlah2AD+9a3w9hGBcNusEpfqBUjmHBaN2etklNvTZ4
2GBMyKBTuuAOLTiOIxMFkoIQqaOmCgimuzp6eP+Bw35vb6p80lhPoDxtz0yDR9ur
v8xAWSbZZ48a+CM6DAd9N5OiIKq7+xBDNYagBVUfdp7fvg0zWX4BZNMwWQquNfRs
l7Sqt15dDsB8oXYIAK+l9SGJ0z9zBajdANc8aYhX1yr1d/htaJFfr5+Lz6UgVkJt
jYt7F2RlWFBAz8/XH3KWjlD/rTuhdLtlZu62qWWhu2nGmfxom1UPoxAt/wBpJFqe
FNwEk2ScGoaQ9IeMBgCInK4RJSl6WsUl3191AZqCorbuqZLtDwK+BOedwO97FSwD
u3dUt6h76fd3Qv33o4z/riP6Br6ZzCXT3Jm0SJw6ACTdwl9ccRmgLresTdfIMEeK
JMjhGR2jbVaw2LceQJxObt0Md3gFJaXBWymolc6QgMM8j8mRv7P/2F7mQ/pGyiom
Vzb/k4vl2FvzWazbWhKOIOCltE9YhgtkoWs2OpQ1U760E4aDauUg5iLNHCkmgqij
4L3W381WlKZHD0vqtPnh8xfi3dXhB6Aixh6jmTbSX9ot3y3NDlXYxBkdgtx5dTO/
Az/OoWDjNHpMZBae1TxeAqg3rHGMW3ZQ31Zic1U8ehkChe7zq6epIYoR8U2ZY4EE
aS3KXj3dkxEJk9+KsN0P5NFuXJVEAbLLWnQcTj/uNWFv9k8gQ9/CcEy540G16Llt
GiE67JQ44aYf9hJFMpHd5SXGSOOp10TO1wK2UJ7tDzOHMP9oenlbl8ZhMeaCfjdC
PQQXazUMY5WgK1p2SkB/QsB5IOJP/xe/oNmUqpfESc1/XicZukHu5joaACa3agV/
4ycSbOYY8lfyBc6ef53ZMcsoqxOKiBVGnusVIqi7qjFbgjTX1mnqz+l520TMgAe3
jm2gUfbHpCm1cjxuh7H2wFwdNH3Xk6/YwvYK48MN6LeF6o1SCYeF5OlMO+L5xcUs
F1dSNqM8qUOxTxbahvvRGEBDDzrmhRTueSLnpxk7nJzR6ss2OaaIWf5wYsefraQi
q2OgRkT8heN70/fgncAx6WBudSJ5qcLx8QqHzKc4BZYd5t14BClmpb2kwjoP4QcW
wCWRrIuwcR5zQA8rEH66eRbyRrZeABoDBz21QCbgJWjBaK3Dh4Zwi895a4YedCCz
KHQ9tCZhBJ97C+DDBaShAv1B6HI4tlVT0rH+6zyK6ejH25APW3BjjwcOsaHncIdO
6Pva0cn/V1p+9p0XNySBgfbzdDFhnjrvA0gWAPFKkOHCSeFbgsrAPX/GIvF9UmhV
MNsb1Fj3PlmxK7yZtvN/9bEG+emONbMKRqoTfVkMPxdfc7+FMogeBmEAOM6yE+Qa
N+NufFlRsSd1xN400mLbUgmaagpuPiGiwHkPaO4rMhnYrpU5lZZAYRMpEU2nSa9m
dT+VVjs4pynE9MUuxcRzp0TkndFQ11wiiaYayOFZsHtIR5YyWEJhWO/huNOF75NQ
130F0sKZjVX502+/16I0hJCJggGbfQAapl/rwhFyERqH5W6XEGAA3520aBk0uvPh
+0J4vc505bSJIzA++RU3SBkEinPW9QkcI0LuChH8gsIZ3mva6qmEkR1xERR/rVzu
tj2yOXo2eUtCXgzcD13rB6HwWDtnd1jHZ3IGtZUoQnmTcMwX+8IhT9QHAj3GdmHG
N3pzSvR6QVFkeHvOPpeQ5q3V3F0g+f5OvdrbtQ2Hl7LrvDNkXAQFNshgM74/Dbpg
EcyuR+v0XtWJ36Uwou+brNuDc7Vi7ZVFuAzvPtVcj8SOZxDCEOvDvZwsXTdyNyJh
St8FUEqjtBsJAiSfdXmVKVPEMqZ1hepyePxiEq1rdpWpQ8AsbfCIfDdQWqOsipHl
RL8i6UPmjSyb7inWTchbXOXMydw8h03AUII0+rpbHzb3f7eFTWvEOIimkAlADE9b
U8/SI0fhaWwxtuGD+2MXKhNijP4NhJxcqD8OmaFH1i1PiWcaxAvRndTtS7KvUGLR
ebXzncMBdRInXuqHiorIGsaJhX+alpbai2OopMOupWW6iDLE1PPfHbKtcUi1DyWJ
/9IdUK+vqG6fefa2yXW063v5nMocYLHrH76pZXXsPneB+RfEqrM0+0bXtdLdMbbH
g/FiM/g4Qg7vg3IdQnVk2gRIgEB17IE5gUW8f34P1J+t+ICE/iSuGRK6Zel4smFh
jyt7INFF0h8xbRzJErBQH9c8zNksQ52uMNhNw3MeDoCpF/tjDeznQoaTA2NknwN+
AFzqn0CGiHYKcuUuS9hfqdQeeScYitqdrdrcBv4i67HIi5pGT+H2iHXGoSUJtTxd
nkAfHim6npX1nvB4K25uwsoGOB74JALIYegkeU48WrCMYImoJhM7gMpyKhRkMHNq
3gx59gNXMT6gPP4zfxkuqCPovrJMdv9MN/My3l+R7p1lzfVsS8KdOU04+lbuCrJI
kYANKRm3IqfzpxAWodI9PTmSglAH9/prQWY/pfXX6PPr3HAWO+Kja6AJA4wYE8fR
z/LQxChMNYhIpxItyC8FRpIeGiBaiFkKMZ177qrDmnBAczSzOk1sbARS1Yc0NpD0
13JP2BoMUA+bxhZ4ibrbC3AkBHAfWLqNHCNnOJqDqBE8ogMvcANADjDzJf4yg6G7
pdP993JdOPY/BGi2WfXEEUkdv1jqD8mO+Bld3mRtKO8Q8yL5JgCSwxUFOq9gy9uw
wnsM1eYRms9e7SOCFd/vxOF0iNbkuBzIIVCOkvftdeYenMNylsYnApVtCklTXGGo
h6ck4lNgYyWZVbmoninSxqBqnpXs8xAFTnL6Qm/Exnoxv1/0S4FTD97Nnow9+7oq
5jqPo9pQB0Min7KUwWg8uAwUFcMUufqrs4lOfgUfkuFIHl/R3R02MgDyB791P8pC
KiNcxsCtlXXdHLUXwka8lQZEIr57nal1boZolgnSOBMWCWnbJtiZLZZG+2UM5JAw
M7cUfJlF7ICfFPckCRWUNrnEmj7FKhiKBgcWnDNjU+pcWhMZTUpEbhMnXiv3CuKW
qUi2tJlvbF9XuLyItAJQ8pGGoKyeTNc6z8gVTEIGvSSF3a7KIVAgwT2dcm4TbdFz
s5tZ019cy4tthfW+4WC4d5nzmxE8q3pLScOP8f+9yyLXarEIhFmKz4nu98S1kpO9
GMzDrJAhfdZ5Twn9PvlYwKvALeBPXoDb17l7ifaSBx0VIw9/K/LWWj5cxH3Erfp3
5yILnydMC37xyd6dTY97gWpRvVEOGlJVSrWqwc+tgKn1ito+cawyX66fMGePbhRe
BYCyU6hdpFeOq5C6mlZfHb/VFkiElsLCbAjN9W5gJjkiLOL2nnf3i2mxvXZWCNcv
YmPbwb2M7r0u02pLhkDkaiTHOW0GiQRqp3VCiD5J+zmEMiaqXloAWM1ImbvsoVVk
WDi/DLh4g9eXBBcrQ5uR7PoKQwahKf5ZWgndJXDFRkPybD/vzjtZLH0V7L2NtY/9
TdFhj28a/KcRFgq5bx+8rFaToz831Sg4OvCHeWyVingx9M0VIrXfwMGeYV/JlkXq
wk0HhaPMh+4W/lkfRmiij5gJN+6oetpulqNfIUhpCJg0ryFAP8PZ3wdKCoLwtg4A
XyPz4fiPHkYwAKWm5dXa2Z6vC9by3gAe05mtQzdMrBJKiK/pv9kypfo76cHWhIw3
umDP5UnPhGEJ2Im5SNwh8/CtkGEndCFWU+OSjzp/R+I1k/KfFSoYbLkpTa1LMnXR
aT5I4KtRb14IVTfmOt7SdbCfbQTJf0n8h00wTj5f6YeOCeKXLbL+IBsngqfLvAEI
q47NWFy8RyfEznwdxfGLjL0bzLrCCfZqAiHkpw9DMtO2Yg/at7Qi+WVBmIb7y0wp
E0hXPdBRP/zOJB9LGk2VuooYHPvY7ZLFbo2+egFS3Y8HO+mAsXRKsBrLkGOCk9Al
KlB8WvUVt/BAqT7SQt2OuVTW4GhiN3Y7EDKcNyOwCjnOgVgFMbTL9Sj2MciuMAvC
o44acDbYXL1sdEDbUFlYbkiS8AsnpHHeZkjaC17+/8ff6U9BC5nY6A4Tfr2M28cl
1G6cVU8auFANbKbEwYjf/ER7KUeSREEytVzFNJQgPNooV1uRPNpRlRZf7xDr+KMn
cIEapJ5AWW5cuyRC59RLa7sv+O682wjQRZdI6IDwMhd6w8q0M0e8sx/IL0s1FldJ
TlguErdIsguL/J432ba2S2Z9wpPoTSxdWwgYzmcJttY4txQ3Apy8AJqfvnaThbo3
0gpr+kLDU0LX86paWlwGek5EpE8PNob6Uq2BfxuF75+rSMf6MpDi5KMkDyyu56yB
m0DzPG24oaP8ER8QF1OWXpYvIE5B7Hgs+1x/puWWRLyEf3Io90uZ0PTLPmvBDbeE
FVvUu6u+TPJBJRKfwql9qrUkF1Q2DACWFR5qcriJJRrf8lrcdmysC2ZvQckxe3Zy
qDcALCr5yur3zYXLlaJ1VWg1WUZyQ1tiXvlY5f0NmLO7EUWx+HK53HMJp9V75gbN
Ra3LsuO3sL69RRaF0t0CfQZaj1Xz077GSM3hyXnsJoT1LRxAkIUP2TWp73cRnyX+
K67HzgRwCIOgOb0/pGNFst5rNvt9JPEYmUc1EpuTZ6otDO14Kh1qHz4gUNLtaE08
GBTCG2k2WmHlQTTbuK7pzSOMMY4xhgJgjEYYtT2ofadKZKyH1Tt6Mn5PA/Z3g2JK
U0AV176IuUg+Or9Vpj6DH2MaU4qAg316GVelBIUKpYIDYzCNRXukApppq0MI6yhw
Uuq5d7NmHNzfFS7QcGQkPDW9TMOZHzyfYJGa/WzaXhZOq+0H0o2J3ShpP7cPdgCN
5ZR7EljTPDu1AzX84xP9+QJ35tEOd9Qn4MSL41n06G4j24KVHDroC14qsewWtHmH
yxu4ASSuO7HH4Zzo9Yi+shEnGNJY5xYK7FcyAAfwh9oF3y+nyqT178e+Qfwge3J4
hxOCC1OeE5JtEHdPOi+8iJWOFJ+0BYKHx0CjaOaUTNHkQxr++OByHQvQzZnDBa5V
MjEULpHErSCu4ZLe+KmX+/SFNV6ITTMXKJE9xeFT2ZVhEppCZmysgNb3uHw3YQLA
Hf3dT1Ir1q32u88mHUVECm1PYuRHquZiYM0nw1C21/WbIYKboSANbSxxvAv/S5Qz
civ2lpmxMfPhRzC9H7yJ2F1/tUj69l+nHum46cb+ZSiNIuqMCIjErK1bqSittITi
fiB4D+6+XGGRXKDFFfZtVkUZatOURBDYUa1bDyqbWtAD9V7GGDmuthM/Bb8rPW47
xeOVPQaG6QKTUPzW7bIMzJF3fhAVxFhNurrShovOQK5xzEv0NQ8uwEOl/2DzIwkK
dVK+ZyKgh0izaVpvQahh6Ky29p6oFRDw4oAYJZn616ZOJ3D0wLck/l3LXONgGHX2
WbVudnNGe3K/gplkYeZgr8wAjp3x0JZxwg+g4dAASkaf0e/+DZEGDXZEXybvmT3s
J2VFRn6i3CxKtQCCAggKgVUaMLyIyKDK7IEt3coTAeUZnBZ03iiatDV1+/MiBGQU
zhvPIaLSJzp/W0YRXHfQVhZFtxZMzAe7s+Ug/pjOEs7DFPN50KDFEsMg1x+vb7A7
NtDY6m6QJarRjwUYnIX5FBhSqF/GEehEU7fQVGRhk+1cjb/ar8doei2mR2m9AtbC
oI+5GMmu6QFvZp3rYHRpPb8PPdwKWPNhK95qSRsHAjzQ0M8RpaUZxqbegmmHc88C
3XWmXarunRw+ajINbBezAlwEM2lGs5sWtjnLVnIJWdp6RkCiVe1cVKUjmISDy1up
wCArcqYZq+Gl42FoJJLDedUbtSsuKHL8uFtlzi0/WHXXbsjXAxLqL2su9/VbGr3G
+votSkQ0wcJQIywCdMCK0h4dJoM56pj8yrnEldMT3Ctg/xUwypPgokwGg8U1NuAa
SLJbIqr4an0jtAJDT5SZtCvdGa6CQCLdHhyIloiKJY5jqICstLomxI21Vl5V4OX9
mPBFdmFZxjGkqusFuyQ1MM921JpuZTxE6EYhIrHizhFCdgyD42OIWCiqsobLGxRl
uLaxPDeNdGrl967SLQwH4DfmXZNEBOUUDuC9HiSJgfThIR/Fw/EL2UKHszmUpAvl
vg/l6Y3/P044dFrbTrEB/82yDpTJCr8lXUB/qsDH1KZR3GysWk44hxFe240fFP06
yVoJWM1YQZFhI5s9sB02hPLKeahQCW2nVirCGo9t4Ozn/6lPzyMLNs8stZQYkmLW
Pn1gT/jFDmtj0a8oGrARryRj5YyeF2soQLOYiOveGgt4mOWJmvxNlreNybvXZnmj
i2sN2pqiNz3eUc7graAzFbCEiEpJFyA0xY0RVcmdJcGlqj+xYddofc5sZ787Hjwg
4/ZNYmauaoxJw5GH46Mfzjt4E7ancBV6wJSEQPoGAyF3q4dt/HnYKoPeSLqlgpIC
KnIRzr8RgnM6OLbKF++mzzY2hcdNGud8eg3G3gke3dnZWT0gnhdnG6m4vQar48oe
GSEbR7jT9qf2FWq1hMzCH/iyIyZQaVAEOscLHVVTKlBt7uhfQsOPtSMetjYN3LcE
DK7clud8tZ+vqya7C2yYv5dgmj7X9HZTNP43PjFGsRDCj7NiXtAjGYEVmFrHtB55
e8tZbzCo+WMouzAdmpHwnC8zNt2d4NwmqeLb4nb8wx1jdmABiPz80MsJw9HkDysQ
UIQOJ/ygi2ZEVrKLoMudnSDHYDmYHaSLGzn79m3dmNNDR7czKqVuODcI49Hb7UQ5
cN+OGqu1R5SoF7vijdgCB0qsh8ck8oGXg1Wxin/n4ofJteYIjvz7KqYaMTzGFdEM
1PPDN0NF4d8SYhl0xqaHwSZBL/PGEFwS/a521c8qlHh9jbZtp+eHpCUvNYar7XOL
30De9ohyS6ua7cBEBSSDqKJs9k/MvVsgG0OEWwLwHNOXUjiggg8CztQdWhVYdJoH
rEzM5LAeHqJERVQqFCPA7bZvF+G53qfzHsEgPH9MzbZ6krg4ZbJtReOY5qKSvGgg
Ye89FqoBBjQ0OazMR4do+v4SPHvSU8Y6Fke7TBeTw0MDZt2dIa3MS/schOpCaoVr
nDa07Pz6T4j0mYDiQyKjm6+bswo8l5H7OStC2Cvx2qs62l/w9X9ry+rFr8wHNKF6
dCjIDfWRG4wOs3mL0w9UUm7MLzClSG7p8NO/1sL+s0N8MtgzCEhNvz/eHwDOiXnF
a7B9Q26wfQOm2dbFwwb/uwZjtzbB3EQE624SWbskQsWKbTOPpYaXSt0nhMiyQWLc
PfBMrA82O783XCPKrfsdKvlJYghl7uBvrsw7YypverTk4gBSHtP0WMM4ifvkjisk
UQEsgc+SF0FbL2dNDqs8b7THpWFd9p30ct9tN2gM62lNEmjSvLxonw7KVSc/ev53
c1k4MzMqVKJwv2QvkgPUxZRImOJ3I/GKa2wuR8/FIWgHjaFX0N3+2HtDf8RGNL7n
QRhOf349MEGYeDvnPBjdmP27dyKZdWSk7qdcU5oouzXK1aoDccKcV7fk5HQvWqDx
I0UYf3AwGpLBRyltDtnU5z7H/JhlMWTaWVRfZsXUZhTDlKg/GfEKwhp74SrlAyn4
QZhcKP7hFTNFmBL6sY2Zk+vBVMj0Id+sIVuLwCA6SAZpnPFxVIOEpixW2gD+R1M+
VjJ0Av6zPud6MLhjQZ4uvsZKDmBX6M4kOhb1K5WgrTZQleB21MYf6bQyXRnsLHPb
pr36/0LM6SwD0fZhgvKLAGs+x9nkrNaivYqfoPxpldv75ykUW9q/Hupx1jlZ0N3d
0eMOICqFoH874kY8x1POKm3vIROqsefPAPqDbybF38Wdic2MqLwUpN25+APKshK9
Nety0iicVtvTfp7TjUCXbMnQ/o08S628AFKgV6gF3Me45HsnArRFrZH0omTA9/pp
xD03LfzC3MOr5UW6eZbvT4lEYLGE5w6nm9lGAQaDiwgdM2RjU7C34MYJVRuomGit
Q45/R2YLdHpzWid3JYgPDnwGRUttOQ2HUDhzbLswr76Ncmn0yWMLBLBCVSWDqinp
2oNVz0w/1BQGOlhtsbZHfWqltjj4Nc653RblMCkmWv/M6huB+9cpiTHWiNTjLvIC
JTQhrYuogO9CMN4kVd98bu0/0gdcWeAU5hZCcugdInSao9rRJ4V9FJDGOZCkx8XU
1w4643OLPjZF8zmCC+dHHbTNzGfihdpsH5Xc5otDS1xBHFUxfGCkGiXdFX2mSpGP
RJAQ8KwrqKXvblNReGxuSWBwdgQOYinllYjIb+vAc+mL0+8KYNVSI1yRF3hyAybj
f2S9QBt/P+xDn3tuDgO1nFx1gElWgEX51cPFMcWVVnkRLAKEvxr2hmRkd8Nac4Pg
8aOqAlmw8XeonalKwI7QJoYtFliMdJ0G9H/cVIJBfqurKNZwWc+J4ftADQz8TUtO
7RQkPHpgw+x2Gwa6klrLp9z05wzymq97APbPJv76AJtp2O3o/HWsFtUbpk9rB2Kb
fN28JTjg9wfQvk580dhy/dVKiqMhzF7yjikGZG2gV5XWIKeQSH2M/EcisdV8awct
reOVqLjxG8X5oKFZEOdg4RW7VpJtOuSEhlW7EUNRmHU18CI/YpYz2p0VpU0Y+6fJ
cWnfBecIbOR5n3/R9UdDJxDpMw1PLQfl8EwewHCUMPprvdL4l2QG/KZBb4c96VjJ
L0fGj8S5mZA6aJ5nttAiA1hSz1uUyBgzEWVTZ7gCGL+fEp9XeKZN0WwOSoQxi368
qVVDgynDKNV8TW5MX/QHJcGURig4dPoQeCaf3HEjm0hTgb7osAZcWaJypka8/o65
cUi61OdfmkseAzFSQoZcaunpcZsBAgz+OUaGnktpSn5hInWeUrVRoYC4+3LBnaDX
lG7qoUHbaQl6n6Dw/PnWVb2+W7+/Z3PA0BqlERIBCbxxnIaRBcCmZGj52e0AvO/R
+Ho9dYro+OC2oN4cQxb6CebJ3fycCMuFHXe2LLTtblssh+tJ5AbZdxYzds/YEg/B
hOMOFISaQYDhewlCWaNmr2ViCcH3vruNuc1tL3kSXonYkhmQJTgJsmr4rqssk7G5
2tWSPKuubUKAAInWyShVluoQhevts3lMdEBM1/8PeT7+kVphC6sYh2qX9hPpkQO/
rqSjoHm6IgB+ywFscVYvJfXSyeL7qV8nJm/10AwNW6EAr7IjESUZ24iNLEV+POtI
Pbmxjotgk5dlh0qrN1kwp9aYC7WV11Zhqxa6ugsvjQ6huz+7j3i/lrPSfavofkKf
GxqmPWy74VTScmUcFy/RuMWvZEPESlkulKEjsFedH6AfTHQd9PaT3dk9O7HMeV8l
/fgXDs17iGxY09Q5Gn67Ta/yJuHZvDGn14DGIaPbksWSMFBT7n1+auvhv0DFMeLb
3Cj0qiH4dynfo9ZONKDZNuLdP5tpKCw5eXV0diXZ3z7qjBckfx8hXyWgp+purOcx
MI/C68wWr1XUl8/dFj7EVMQRVEOozIW8+4z2LtQP2KK8ZwcMP+v+avDlJsF+7y6u
5QSTLwEikmMflZH7Sbknc5J+xl+puIzZ5n83SIsc/RmnGGIEjwRqULSGeNcTz3/W
+nzmF+REGESUO2IsXo+qkLjmXpLd6NtYn8lKFSyhvxDcDvryCQRvJ/ZYs3W+tzwB
+f87o1MR+9OSVGgZoXzj9L1gJk6BBNf0n3eP1tZnXX2XRA5IqMUyMGURJ8WKW77a
Yr2jLa7xG2+/HxD/4vNYJAsVbcohk/TLTU7NKx6lzVhK5SGM/BGjB89TC9NGAR7Z
LoCWI99II0i0x1gySnyw2/FFtKTREZJFAhbot0DGP2lKOlBR/u7C4bcsPgqIsvRP
xH9U+FvqyKShbYSlx85G2jrBRDgVwb9WXqauoUjvvhX92OdxjqByqX49JNqXnyRK
H8Qt8sczyp3gDcduAAILK5Par5gq8haflXQJABgJPzgWF1lksgIQTCqx+IcpkVT4
3VkfjLuZnpG7nTxFkteus3F2OpFFl2FntlRsHC/6wUQ6qXrr+PlFw+MtlV9N68Rs
1PLvgHTmQNNseUOKC1wWXr/Y5g0cNkihZ0BuNactzOTXtHQDtDulFtv/AYYP8Ae0
lYOtXRFAcYaJmPSePyr1XMcpwrliQFght1my7hpxE/3Z9iLLKTUsJl0tVkKQlXZD
HeT2lFXiqt1YGwB6gT+HILA0DWHeouec+KaqZHZigfXL0mmMkBiGsRNlFLI4J79N
0vjqUfpmsmPgGLwE4QXfhej4Id5MBWv1B5ERsWIBCAMCzjWl19pYhLPbZKCBWlIF
CdZknkLfNrhjMG8yRkwEWWjYnXMSYu2dZxPk8nUgxmcM0q3vA9OQ+Z4MGJoo0+z7
u1rFpzGOs/H9xJkWqonXBXoOnuaSyWJW7f4vLzhgKKsaYarPQ1DqmC8RpmY3xe8B
2Cq9d1W2vzZUltsuebOK1RJeg7JwTVUHR3HxvUvwoSmCFTy8/97FYv3QdPUh7Bc5
HSR2snjv/RLyHtNqfl4/vNgUf4it7figXZ0CZUUhXlQFowFTNZlhA6felVPEL3xV
10Ed2tR/trpBpqx6Pa1mY04MZEQlNqHDif2EsAJr6aZXG1V+9exh9Ul5+UkJX4yu
VBPD+3LMwfAjje0UpXWYExHEaFcrksqMD65JDF6xBl6OE1UO2C/CXJ0rBNlJ/vG1
jbdG0/UvPT+8gJtpEwtAck2kNtaniEuRTlCIcJuXl3XwNgtHf48sjUq+LeSdgNdD
CtQAUVxm1QLdWMgwIczv3NvzjwikHQKKCulUD9cR4ERg93v+MlwH6mt8akzeCwaC
V7cMDIKnBfYryV/1i5MF9lGlNC8vUofTtPwhUGT9FUU1SM7QwewQOpHDHLJyL1Vt
GhkiFG+tLoT8+WOM1+t3g6SFw7BI91Hf57YBA9I2gZl/Wf4kEtvz1r1Njra55o8P
0yRzqrgPJ2vHF9pCTKLZPBFspwAZGipJ9uYzkQDPH/r3QqS0WeVmn+MF5w7S9HL7
fMCQr1DFteiefbrRYE4Trf5tlNqmY+u813M2jn/QfEeef5zFulff0o2KzyNsBdMQ
Hnb1pA9IFsKe95M8boRNPy/nOyDs+V8NvjsDbtXnyKgd4Exdqez5sy6d0Zs6pPoW
r+QI2rvwAxD6axxIkFdjXadzpax/z6kds1uVnF8LXgIw/jJfWH7/p1zOq4W7DNhM
Pv+O4K9m5ol62w8VUTutdlNpwpJlDBGkoeduCCEyr6AIIfxa/sFakFYkKsTK1WGT
QXrCEfsQeDpPXxZya/VfQr6hn8MHjKNUD7C0PlhDSThbDxH3u5Po+tmKKDz39/8W
8Zdrn6vmvbgw9TWBnre7cmRVF15EiTeCMeAL6uX9Tk8Ecjx4SSZZ1mtiFRuCUki7
mExVFGdK68BFxsUaL9EfA2TfVQ2UkrMwvrv70LlnOJLBBPFTfCiuvtIk3xAxq3y8
BeJgEYzq8H+qh/4/ufdKOE5ZtnZPg7wi/f5nUBFlm9gAZ2w1Us/mBy9i136iuFIp
J0Tnr47GO+JrYmITf33ifs3Vq/5jpojwkb72qHqJ+PhZ+I7Xs/Xu565LRqOc7EO0
N1Ys7HA4GMaksiIWnXXzaqY6L4b7f9h5ghbThtamHYzV98mCjnk+963xiFFoAF+C
Wv8lVDNSc8B2+Z41xJ1KfjyYZgF6vN0fNbuwOHFu5fBpMPGSYnZ1UV1T/y+ESec8
QfMH0zw8Qp/97vaQbSfWGmoaiEVbXuO4f35zFgXbKaFBz0lYvDg0Meh6RjvsqHUJ
0GsAMJ+ItfbNufOBSiX0nfzyw/nrKSJx4xfIBKH6jthR4F7+7NLRe861NENDB/Rs
ghxt3H1+vADk/DNwCcJvwpHJnQWVMWFmYMB1Gsj8olsiKqK0CHhyY+Mtxe81S2Hu
cr5QHEuJLCmvZHZdkoA1I6FjIy/WjPl593OoobQqphljZoNM5Lg7ZydNWHK+2Wwv
3czLANnxhx8wFePq0U2sV1mNuvCsK1TPFZjGdpWYOXof8rZH7j+B6o4+Pk3Gbm/j
4aB+g95C5J6S2n/VU3Re3rBRcUn1f9g5cJEc3Y1OCrFvVhkV2JkJLRw3poGD0ZPl
1Mrtsxbqb78uT5vvVXYFPGVNkEbbXCj1BuI54IoGR+GRmJRkcIChktBtgcBMDL+C
6h/fJquiAKEfDY2u/M7uRxc5QnIvrUz6RzmbqBDP7O7MFdlAcHItHUrIVV96t6CH
6p3Gw5pTLdXbB2uC/HxAXUYK5PzNxFNa14sd1ah+mABmDek3DbBrSNY1AnFlZ7zS
/Dwj2uYs27TPrW6awk0yQIV0D9xwcwUi3hOQ1m12Ee65UFD1Mff5ns4JrZcIdbH9
ZuteXNDgW/n/7Sxn1bOX1AYpApa+jLNpl8gkW7JBV2Rcw3k0Rp6pWBjOV9kzQ2eq
B+DEUx4KaXrXtH16z7XK+5sk0n1nkeYkAwZP+DUWQFOxE3Vn7NJd+QL3/YTGEEJY
jQCWqhcV3Cwdhbmu0Y5yMKPcJa0cl9/Dl5X4sbkbn7RBiUNdD9EYDHEqJ2K3sx8B
mpgcx6gz73/LoavIrrPOA0cgHnGaNLsH4yBrLdVB1aOU4EBDTRiBeZ0rTUULmh3Z
wm3qAnlbHoqjPEZSebnVYQYXECfWHHXNc6mpUKPHIbQ/DoE0Qpdgr9PDnlWtDFW7
dPGHV6jt5MGWr3mNlAoGIpvwaCD2iwnRzA5buINh7Uz9XKu4+8/3O469R8A02FMq
XJ4gpFZNa6fD7/ntg78tEcU2+39/qX/928jt4D/Pb0EWodGJnpYgeR5xwWgIvRfs
KpD9T+uNi9Te9uMi6AmlqyGAv5lyksWFg0zOK/oMXApGBrtTrINuxp1cdc8Cxf/z
UGwNVj49UaRyBFieqz2vKc4JGkF+tqxT/V4D7LRYO8wT6sAXVHbuBao263iF6His
CzRrCcaTC1fxdxgHXo+O0y1uQyKPSlh53SJypB8u/6laBPLrOU7DNaP32Ho2umsO
+Ddb5TRJGFzuF0l5ngKJlE7mrhgvmyhGGSVEr6MOvMZQeggTIq5DkLnVwpW0mbKd
k4MhRnzNrZaV+3bFb2qGn76ZBoRXNR3O54dfdNQnRVg4Fib3IYZVMpATuVazGsJj
XntpmgmfCC7/yukQ3+kMZbRz1k01xQIlo+C957masVZkGY+8hHLIl8AA4/um5tNw
56WLErkOjXvtbxM8G2mj6Odo7ioj7AS76VNU0Tg3x8MQ4S8Qg63bMhSJWU98BNXK
hoOfgkbfn68o9tkXkH1q7eODtmNJa2kuvyjzwVN91SyGdDBnhmgSU06vFz69Pe0q
wAiACdb5UaHuDU6bifVUthJ9+2be/q+O1U2BBbmnwiKLQCo5xWxPQKZHsjq21/rT
ceJHbwbqGstBIWM+2VRwI0aHMU/baY8HxUwh2HmqabEj9ESIZKn+29ctb/lwb//J
Y7hFfJvhr+aGx0OQaj3WXl2eeov0sYkoYLxsjQ/7O++BRIH0u5cFHvZOW/kZavk8
9oBJn10T/ufzln6tjntVeVHJgS6aYB+OO3f6FpluhC4yHm7bGIzJhxvlUON67Cfl
m7LU8vKtChGkxelZ8ptMAzq8FmZXnEC4ucAZq1hM5xJw2u3m+o2YI7pnbQ4heBwi
clxG4vNkkXF+fkU/Mljjnyy2uLUBAHAfLCXNR24HxGSipz7s7r9CusoCSzO5/XAY
kk56MhQjdgIAZxEK7uliAZkAkp2FZ2EBZysv7bnnV+FYxTWgbhc9ymK31Qtt/Aty
WRc5Bm/kdPOCbwikDgCp1AD652e0YjtSa34f47jmqL9PTUdmBWOEHvf9K7EwbHWU
iIYKHUgPHxD1JTC6Y69k3yt1as/E6qhPnYJEwy5+x8hlApAb7nuW+qOxr6mkpX3O
PpLEfX/BvJQu17yJjKVJvLoLC2ndGqCUkxLvqDZ0HLHYX3C4eDE/6HvOcfDCchci
DiGqBja0/E5paNwuaVJ5ZQgq+Ezvtxv+R6bnPSmW37B0YYZX6VHoab1hkc5uEXoj
0Q9f3w9JMa3LF9hQVabhuDuaJNPRgmwPEu1mbVUiV7BwPuKn3AbxMX/hBoiYXe6K
Ve0EW/XqKiMisl5/vjZ4xrTMW6toUgbxh7zlKuk8dyDW0b3okyLtngoqccGH25Wv
s0rDk/l0MrWgEd0MZ08i/BccmS3UyvnxuvQltrMvt35AOt5xOBnOvsfC+d/FlvgL
i+oEMNzbx2P9iCdzU8TKJqv6f8NE/JCUP+weRd0UFvNRGCeRSYvz+2kyv6kUkGhw
4YjO9hA/yMNNHGXQK7VyeVJMXuN1d5rZlcK4NaXOG+3JwhrVuUNxGfvZWweCWdgz
hTXjRrhWXg4laidDxgkZ5atLI2zEl55Jh0ljfTGlqPdnZucUEW5q+Q45r3GS0Q4W
rsOYqrq3JkOD/yHROwTNl9SStYZ51rt37SdKLXtBgfBcFv7SyyY3wqGblrmhpy3F
6foA6bhdYivho6Qr7Rkpxs/0aD9GcXSEz4qTO63UflkYNOiv0sBhDiCQpkwVoyA9
E52tWF3zFcRExglElTfa5aTuWlz0mz0FwXy7oiHQ7aXJniSYXV0PykD6X7rhOsSB
ftm1M7768uJqQxU2Elyj79tHkqPssrgT0qUd8qWR59Vwi15k3yoY4WH8OVnphjnG
zzRHic8l2vnsbx05Hqj+L7pTUztTAcOjIMFgQH+3owj7lBt/SBNiHF68DfQ0axtJ
2axpoMYMFZioXmeS4Sj5uKGLI5J+4OCHAv/Q241ybv/YncZeNkPFUYkW5beY9xPf
Gec4GdRHxrGCM/Jly2uLrJ7DjMBBpatJp3KHM6f2c+652Axdcpcxh37/oQTsDu6R
b2OrBr3Q10fmxLSGmbh5aUdjFsk1byKC+w5OXdY/oIlSnQf+VLHaX4Hmp2l063lo
6pj0ZBOCx4F7fxlDovcIrZPjkmQFs+1WO8UySpFfTe4vGxiuixtZFbg83AxnxeSQ
X9G8w7SLQMRkGP9jkYe4AYOcaIGKDYmcMkt2cRVfhLAgxL3iE+jcW5ybFwd1vfk8
FGI76yTU29Q0/+8GxmXv1MAGaLukUZhPpYkDFfpDJ5J01ZcFJb485FKnwMPdY5rl
cAJLkvUuR0csTJmWUHqv9byWo9rZra2tgpEsqS0g7UMT+QU95p6qUQuz/EQf033g
xqwLznbpU02WUjujfwD7CblkftPLWF/VZEou5qcNcol6n9VVQjTQBxWwot3gql7X
Daf/LTF+yyAsGdh900boCmr9OODEiQlehIsufumx65WpRC2/UwbYvlW7Q3HwYh/A
rOX9TILfQwTdBx19HciiIeVgfJAuKW6L/kObg/JKvY3FzVtIjBBFMF4pWrCaCrPw
uhyH72r4GOXLI+qFdy9F0YTmz7t2B3Cl6XqHgeejHpi3AccN7xzT2XMZUD4ax7CY
hzT2pHKV8asU4DLXEGjitroSZPkX0Ve+uPGfEUeYTcukw6xijceuMcJcmBa4ib0D
fWgCkkEwzcYsZbCGR/+X0PrjWD4plkLnzACtvdoC36p9VL/P+826uZcHGk/Nn/cp
1VEbCC09pRfjgjpwl1e+RpsW7J595XMeR5dAsATPYsZseEnN1qLGGoDTWAr2p9gb
vlrOxaEU/15JPu4ZGE5qVv+a1ePjtFbnGEsRTJ/EpSKKvmAJk/Y+L2oLWCAYj7jf
8Bj0Oj/dm7ClYvBe/y7SoLhGHlbBWq0dKF413/NFOgcRY11HuermJLAAtFjrlA54
+60rAQyszS0+SvWC4m22Akag9vga5wel8lQ8nv5ec+nTWh45L/UQ+NzvDorR6ULG
IQTZHcgQDlfErlYAB+A6tgbrJ+zI+HtteECbqu24l545NrXsa2PpqdUKKRAhXBl6
Qv4kJ39A3evNDHoR3G/Kx4onTVfONInlo0vvEKstpa8p6UfmNjBqZLZy34QwQLjb
eu3LAh+oKtZjB/B8Uv+PuLrV5IF9/hEFxQlonpt8rxHZMEsHBLrdtDuSUtqmzHOs
+/+WN8NcoMBwhA99UWv4+SZix2n3bYebbyF081QxsLZkMi0WfW9JqdlAETfT6vJP
w0UT+bPH8f53BmKcaGJg6uLFhEBz/oBqM7+dslUlRJoIckDx1+c3iInMpPgmIPUP
l0ww8AQ6xKVPlh3VA7qIv3P2uhtQfTdsejT62k5jQSmXlUJYnxTI3AKBekNhMeRE
DsOL2/t7oV+ntUjB+oDNwh60MMvMD5BJGngXGEJIhbvanNkXGYcNv0vt4HeUNpj8
KAMPVliyM1GNeYXfjfzvtC+d3aW4vbf5BXEmQ29WGwnQ/OAxX4lD6rAiSReh4Jhp
NGPGVd5mTcoWC0wIohazEslF1zIxfnvsJb8bo6BtZnS7GGt3s9ayH3NmyUqZWc7b
+wrBe7GS0SOwn+g0CvomZvXZN32lY4whnsBzQGqdDROxiOWnDZ4waoUCFSUmUzfo
Ry7/M8hu2uIspGZ4j9P0DCaSsXfd1fCSQ9vxFXcyi4t4ORbQP1fXi22eiKIK06ve
xz+STxfSEckxoeqKGOjD2I4vgn+MklvHtbraKuRLx4o/pGIvXSGN9O2W4f7FJB4V
uhmJrD1jEhS2L+Fa6CukKegxVN1rx4jX/WAAro7cXNuy7cqzzKnSk/NXcXLGpHUD
xZ3FhaQ0eXxgfgJN7/HRmzjKmWaoI06vaF7gv/aPV2MAhPDhEzS3lWRt9oNFWCHs
mYUlaCwF3+kp/3f+7PlwaQPK4kfuJxhoqDyGAg3JCMBBRYvBeKG1vq6Zz6Oqa5/V
Ezaz2p8/h08tPyIg8Qh/KlzaQnkZMStbzvIN+Yhf+lBK6W9BXZXf/A+uVFQ4JVzL
XZMa8i9xzq0GDAyTh2+7dS2SsliH48Lm7owtUYYJ9prAiJg3tQ5H9IW4vb09hsrG
ylOqeaaRueZoRLB1p5fvg0BpfsIqHIesswHnnHeuPcNmuigeSREUWb4TCkqRGwvU
Hw6oOmc8TJmauikj60h0o4Mxd+WX7jo6Oche4aTPZgdG1KL5mcArqPEB7Hv6wplA
odDYCcwKJSwTHVI8L9IL7rqlMn8fEZ762IyVH4Zi7A7GXZGl9Oav6tr3h2Z+M8aL
i+HtBelcywA5wGcGdh5utHtalUmopApQZa4cHxGbv/ucuzFVjit9i6u3GZSWnBYT
uYtT6N2RUk+ZeQ0lRIcsnsdQHfvzBdWepOAx69E8mM7IcyFDv2GxFKoZoVaKGryg
t0i014pcZ3uMgbB1vlSxw40PB0j9Tstun+uFfbLWZDkVJUZM35/HY269FfNIwWOS
PLK7lCQmfGIxLgqkEfuhrsLO1ROhInZ7/s5lt00+w3wdI5NKB9U7p8emGRIU+A4T
x06EWN5pXNehim3vQzQO08kOISLB7urDO3gZhVWd2fE1h9VDT5SKT7u+F5hdkCgK
o9cLKO6Rygj390PQiQVzSfINe+R6nkVm/qNrszgyDuOyHcIRyqaIYf6UrUyTOluh
pJ8ahTVLU6pqrD+ffJPzbSN2Z8f57fK13mFJ9VKOIVqB18bhq+Et+DiUmWkrYX/g
fn0Iv74zab/NffD0yzsJYGBY1g+6voKzwp0t6QmJaYZ/p6KeBLHT/Tci89XK87DY
S4TPTV/l/l7LN7Vt7cdWoM1E3rzQaaIvynp4GWQfma9PkLDmbfwQTBegpVZw8qm5
PDUxuajW8nqnLB+lIs/vIFGr8Ce8xImyCN+HmkO3xEJik8V39FKdy4dYjY9LzcNi
sidbu5sLQys7toaalg2Kh2Oc6aY1XrBm6ldZizDovoYxlWj6N8QJUf4oKWDIWi8z
VRo1cua6URalMrrVmGsrcGKRop5oxlNpV1GXVTVUIjiXky8n5FxXV30ZU/ehHWGD
NJAIG7eaV5AfWWPAh+g7Gmh/En0dGYsUtaFIh7SE0SQyxvOrLzP+mIV6R7+T3VfE
8JewBbgoCri79cpFFlVFEz9ugUW3QYmGnE0JIe5MkQZE36eK0hsPyBXN6cf2AYPa
kkOFCN1N0VFy6IIR6bpsm4BtVjW+ry4r0YauJw1gegJ2ijEKIC3gPHmhIRWt4qNZ
7+p4Vl7q0nDumaVL777kXn5kvPBbO53ZT1R5UInfCO6oxDiVZxuulg/f/5ZOPD88
a2WVebEGHJ6X/wbpIq5GYk2yY66pBfEFJZ2j6mS9VhzzAQAbKZo6QeuAtT050UqN
0t/Q8jHXDmsDsI/hFnW/Kg8av+j3XKHMRZMBbahEqYRM3XPZ+dIyVWPyhJYMMZZb
RI0zpmkllPnYdXAh8IwKrB27SQCKuRux0eZFdANfURNrlmK7ecSL/qXn2y0gGv/T
XnSfGYUsGcDcDaZXKH7hfCQDsCQba3r73x4/U/1Md6zGK/8SJn7i+jf6WwncjFV4
QeQitrWo5yilHddn+XFZvlwAjdyoT6PGTAFtZgkz/ZIyb2dcTEUCdCkxlxUnG21Q
P+dljwALFoDh5wxE45RXNjEKiGtbeXzDNFSWLZRsuSGndaH8hv+hX+LHCM52XnrW
a1p20VNJqKLA72CjHSKVXDPQx1bQ8XGE09gf9F8faFfpVEbcDyfI5fr4RhA3AstA
KjccTylsqEd9bEs8YUZKpvknbWxipUkly5EpFYfbdJ2XyAhZ2xn2guu2k+0JjpRI
T+CxtdTU2tjPg1DW25DqwEoN8JPb0eYS6PQtbMOm+IDTsjAonJ2rQk9O55cJiLGs
ESIMsE6QoaqQLQ0f2IYIfd2y9PzdZR570DnBlTJsvbJOIig6Zt4eNvZHB/lFo27z
bsvs+hgot5PpAMVzaCX76wYtsOzwbK4UIgz8kSANR0eXflAZqujL9ol1Ucz4gMFw
g4uXpofQaQYZbeyC8mL7r9pp8Udz7m12iLuN56gkNwGuM6MItTYPtRA4jpvSrZUF
aOXp3wupsR0GDsnCoFIkZAHSZOOXS9p3x5f5lENMF7SUMaaKtG/Fpjo8jKTF8X/H
P8kmaFt+TdJgwANDrrDI4qJCx5Ukt9f/vGaWuwEt49qP+a4RVO03iqLNRRb/S2aK
26zp/VGCN2lehEaw/Uzpbgc7A88wZ+znX6PKThHHevLRNJBCEO89VOr4MYZhgb9V
o956xEvJgr5Z4nxX0oqF1PufMwz102Nz1WbOgF+nQAOZK6Lq2Xk62PzcDcgVNsbE
ShGTCcH1SLZCGVRzjoJjpBnoQgr7LLmHQelfXoabpsnSzUruxqw5y2cYi1zAGWdf
+0c51KpfFntHCiyZjz7jER8qQ3QtSOgrpVoo6kmyocjAa1ccaVC58YoCVknD3JdO
HHlkY80Mi9ilRrQj3+0J69k74Z+4+D05zvOKGBm1/2ErBXiWT9EwaaHc7vUkY/ZB
1NcqBJniJedWUr5RQCZ03o4YDWDWzOXZQoSAyoatBWrTnWvimnggWY3pi6NMmDEs
78xD8pvYcqa21ldABb8vBom0xJ/AP1Y2c3LwotxnVsRoZarKIyJD7vqHxB4BERHK
DglXstqMG4Xb6NC38M0aw5eu/tgrW+ujiwVKlMxxUTARZbDE/mXFlLWDLPn+Bx26
ueOj4qCUfsalnrtuVkWX91fnLdo8J59VG/J4VLcQ3eZut2Zl1qSm1nbGYxAjT0Y7
/0eEdbdTlEt5zQTw0t1/nwaPnFW8/sHTvBzWtLtrTKkbfYWNPWsTdr3uMW5WAwJH
84rHt4Z2FUPJAm3qRzE7L9x30EUtzhi+eK7Xn8xBuLf4IvFFxBJJ6G5S3MMYrbxw
NOu9k0W7rjt+rkLkSW9zg27b15Oa+A9dSUx8ob0yJFEY05P8XxTWJVEHupNfDU1X
TKL2zHdbLZOA/91AfMMFj3K3i31xy7yNvyftXufOyMhgJn1JG1c8fFwumps+ZnQS
mwbg1nFvrOPb4dXd7VYuUduRw1sQVZDbVbqi4xFKR+e6KF4O09X9l5WQo9NM7vuB
qeEmI3PtrI2X1y0fGAYRjheZ3c36z37pe3d0ahCLwNfp9qGfScf0kl3DgvKemgf8
Dv+LboHr1OaRZWCySDgyicHRDjx/r5i2x4X2/FVoGH0bE4VY8yeHF59Q33afgo8M
EumOTEJKKgBFBpjd0PgcP1IuSinnI96o4P54ef+JRVoFNUVc6aYCHIJoThNu6ATG
TB5Rwl23VXZFG80Aj4IPKVc0jaa7lSEQ6z2lscPlyGGBIBefTTJStz5RqcLdVyfg
wF4G7O6BXlN82EZTkjEjaR021pAv57snfONP2ixejmo5tSVsRga3b/ldJunMJYBV
YNL6aw6CMu2ob7CL/6VQpuHSifIe+rZ8VQl0yYFMNmtHSaBLfYoVAmQ7kYmnLzSd
pimjTRbezfplzuaSe9NMNQxkZu0tejGQSMErNx0AH4OoVA5Z4hAmswG6RtXzVNFh
m6u6iKW6kGdRY7YgqYdf4TsV/cbKCZoOMtdaHkB7VRkcMzL2UPkMvw7WWbZNvsY0
yTVRLFESzAo0h3WqOF4/Q5jE47j2PTuwlA+q1MYnXHXZfydp8HmUX8EaLCPS4S6a
GIvPd3LRg1pocA78dhfvThXxXn13gbu9RRNl3s9WRa6J+614HbOUDgGqSJsT9Gxf
by7oJ4EKMdQAKkqdDs1mqIZEkmSh42TJwB3UhEZVTtZ8dqWai9BJurLSDLIg7XNH
BCumi8rmDLkYB7mQCuCI8zcWuynfVlDHyZBmcsS9lnsFy0FvS3XcP+MUyxQYFdLQ
r5PTunCLz1erZfuLNhgMxYws9N/zLFOv9w8swsPYmmmemAjAzS9JMIenX5e9nbNr
SlftrorWk6QiOJWKLG+gh4oYxwNM/eZDOuMPUKNX3FInijyDlKVpr6ODGfSXI733
bfWXVFoR1tmcwc+Jih1x2OqE42mO3izPcdVN08lIigS+QsCdlgx73CVpq/TrHwxG
s7hkTw+/mqfc3oqq8z5Borigci9/Y6/4bMUNMJtYMvMjTrY4MfzxwzWnqwAfQARq
KoFvvlrRPif7GwzlxYkQK9IG75GJgiei2Xoxv9E5A7GbvqQPwhPZM+0EP04WZNYo
x6wDxDhQZAVLZwSzzzL4jPgIdMu3HMJVM52Qr7TL628pi8DsAdONEfl6iZadkVcU
zNzK34ysRUiahfztPgMpP4wOOLhPiGqXkpuLlBUFF4EUVXhh5hUcCi+wNSI9Y8kk
P2WJtotgy5FSXle1oSkqINmWnEIa8WJ2xnumGdYHoOKicq9PcpE13m2sMPTthF0A
q+JTaw/tkczqSZdN403WapOFtBJH108mt5TNS7WYZHZj62SrK0dpOy1Ng7jzJq2+
GPSzrRBc7Wvk6CRPhkyBA239Ez39dVu31D9GKWnSjRBmExuakOehpsdDwbrPuR/K
Y/EvDQXbem47UO+1spfo4rOHmEw7LW9vwLjdtlkoC93GcS2tv/Nd9heQ6lUu/DmY
maLW2Mg/N9HuGDJXoi+gtBjfVw06btgFlpY+YVvKA1IOGc/RnoH9dr+6KnSzYBFe
IcO/InrRSFpWha4mOJqhuNiU85GPsAH802wEQ+QMRZ82CYzfcgvqU2pUSAeAL84O
B6BoRB742kERCFhmD0CmYqduDsbHRXfiqYNr2nfNPhc/oKQfP8BaqOqFyLdl63VU
NhVJnLHXWzhS/hV+2UBgJH8zkqcE7vXxacRfOjBfb85euA1VZYSOVXXamR/C1SMD
/S9qYHwcljuYZsFwX+A8f+4lm2TeEwNa5HQKGNzP1p4zbsuM8fPYna2famYlLquJ
ltTL6KpVN+BSzxaCaLp3IeNlc6q+xky5LBVhqyhpPYpdc8O431hnZXudHTaQ6dCH
kPgECHWpkn+WUs7Qyh17PRPwrbdz/cUFLe+Y8G/hqUuH76BdQm8osOtIpAN+7SYF
EsgOwUTeytSPZDL4WBH+ofrCWlryqSY4whTQyDnspFePusBsDgoj6B/Yi1t2Bgih
kRVse6QYOWL12mFQiA9lrCJLsMFvfySFpyGwBM9oQnRbSmSpftBmGpXXfxPsJ9++
gABHorMU0w+8M3jYZSM2fLGV6bNtCVfTUbc93LpMbgXE+/BVE2f27Od3QS/Ubz2E
COE2ojURHvV7XlAfMpZiKFzVvBlWybz3oT7b+rw0fMU0C2OL2qrNUUgYavfOyVcw
3S2fB0IcIM8hgRpRu81e1/H3j0k/t4vZAjSh6rXXh5EH4d11Dg6UMAtEau2a7KxW
rv7eBGiPq9+CXK4d1wUxdYRtqM1KGxUBJQw38Ig04/pSEXXoA6yglKiPzBYYBJo9
rDTPxW6Cx4cTxwoOfkKy8p0Xu5rvwygIanlP1LhvOiuHhVl/BKhO7HPgvjZYShXb
a6vlUmiCvYw1a9+0DFhu6vpjghmLPJPQEYu96bNVbBlly5BqrO9mo+BSHsANzQGP
t3W9QnNSOm+RfiaZAEVti0qqQDH00tru3aEzRnezXoZHG78Nt32HH21/x6Cd4j+F
NpvkGBezgll7eo7d5lWD4NRcOifNMmVKAYpDv8euXDU2yWU1pUHVPL+F7tEkKM3w
Sc9tBuQu/Hrsp0MGpkO+Rddu8Dif1os9R2Xaly0PVIk5h4sivyTtR2H8yzn3w62U
TBP1XBUxucMKPDF3vFaoCdB/V/JCn2PGL33PJX/THVBRP+uw//5swuq71ay7q/EB
Y66aCaDkAd1HjVzu1UKUZJ4LPmthZ9lOtkeKSEu46/v8VI8hdrdAfxyok5ExMhKU
QZS/qsSp+leTQMWyPRhlU7uvkdqIGF0sFIo/tRX+vqDjrxPqXlwlIHzfnra2w7sE
4iJJ3DDL2dlA9qQgBu3nJnv2fIm7C3+mGNZrBn7tNgIiiPt4SMEXvt9T4HSJcujv
uIlPXoeno9lYwvfWc4ALmVJX7wcVnTqoIQenGyTofEc0OxkmoxCejrBcZ/qyvF+0
/Gyc+gYL9budlvt0F2Q6sM2CV/undlY30j//UhL/Q1KrIM2n3YYy/aadb58goGAc
xWA3woJva8VMm7xF3kKqlmI2oOBA8RAP/Wp9sn22VcuCbgeyBSY5t24TxXBs1Brk
LZogXwUuVhsWZ8zifeg4K1CcapOXRtsmpfr+lSPuZAOuZK47FEJ/qvyxhCML/SuE
cWtppEqk9InD0toP7O20/UXIdXgMjI+ln53Qgkj/5WVl6umSEM402H2s+8POFVBA
dx/Hs+oQ3AwEEyOGDP2kHDTd/Cb/LPVSMdqR7XEqbM0DxsQ5EoXHpBKhtY1BVnVk
xOq0HsX3ya0WzQHjY8QMVWj4ASymPmB148WU3CHZbZEPQCw2Rv8j4FviK/bt58B1
ezQsisT8wy0n6JwsLPC85OaH7Xo1N0GSQNlPhyvvA56HmqLrQte1/+DIM4OP4+vq
virClHmJMAlW+fbT9SgqYuE372mpgPPIxagfmW99Pp7fnkKRrB3EgJQ53+Tr9AQQ
9vcldYSZoC65PmbHqjjWCLALlXzORw91HAfjOd7Sp9sUS+tvU6iNtXtUTIzyviwD
OJJgQ6a0X3KG4D60NL0Z2AoHmx9+BseGdaZ8XG7YNreKarknHFn1h4ATfm/AtltL
2i5SdVOhiO1z1OcTEX4URiQbgOb/GQ0P3qZhx52sXfqyged6w/g+x9u79NqEz+B4
PxX/QpOBnf0UeTug0QnCtuU7PNby8rPlxenDUMDmuEvkhcn2lLS1qoYIY9/Hthvc
X485F8B5wpfyXrBukwAMWz5hYY7Lo6tL/sFU6GZwEkKqwk13pdMOFIf2EkfRme6a
jqZJhNSC3vi7ilwmAFwwI44BJCLcYbgv0mKKY94FLhwe7K7Ij1T670PAOj8dYoQl
MJrj7UWbfb/n6e0GfIDUgowcWJD6TiinebhiW27yaYQSGG00/CyO3Dvpy4XHH59h
X9i+2BnKbFaftxBExcIPY/d260jQfjChB4XavB7u2r01Z/4Xs1igyWaTOkmohvsM
7xzI0PIpYSAbFRhQea+lR02AnccgfL5CLHpbnGwPZfiIhjhPoGXFPs7MuK/Jg1IN
oAwNeKSsF+yFLNlccUt379C0MQmwGhdSTE58HOdt8OqFX1wOmJ1oLQry/S8eHr3a
KeVTsRt76nKk1htZq9LSiDuKgmA4qEOUnz35yID2kWgAZ3phrqPALVBX8a+zdwn7
ESGslncN1MNADAGSZbZ+TWjfZ2oQ9L8jok6ZQd30NE2YoiEFRYf9tU8LNJBxDMPq
DUjSs4IyGV055R+tgeSjts5yTcS6kdQi+7+9FSRF3eS4purN+zfsaTltBO01bOuE
c6A11e6EJ1+nDJcB1udu4528ErHAHMShv4ohjcvJ9AZj3ueb2fEfDr/8oi2qtQ4g
x8ErWJ+amDq9TeTc/HSM05TUvTguBLp3ecKWihwvCeL30HbQ8GUGGz6aTuBYHRyZ
2jhDNIddhvuUVGoN7aVWYOmoYZxVR2el6R8yimNLH4pCWCYC6XHvXJP/abeQmmtB
7nwN/cnNHR3EApjcbMD7CfyQkPl4vfFA3iqf2HFobdoFfq/EbLKx1LJjfE17wvfO
pWMj99L2942e/h1zA93M+v/WztNhQg66bYj+7WcjFSrE7G61rY6NNaq+xcluGJqA
5IVpeA8xGEvbyQLj+Z//M2MsXzQ8GcdU8sNV9yh+hJ24KnS5x+5VHbYO5VfU306R
iEmbTMe5pDseUUp4mVgYMhsGdwfr4ycP3kS6QwgIeIWLfR4aie8nJARu2CTP3eUB
7h4if+y8Wx1fxlTGpc5kBDYzurP9VdsRlpEC4M1AV2sorpnQ7QGFCd1GqZQ/K616
rrDvM3wPnaqaFClsRzCrzvs+FXwxVNPxhBA/UJB1mYuwQgAOcWni5JSa6kEjcB58
SGi60nAIiRyJypKXybola3qy+coMZXdpxZw+CEgw1X3yBPz9CttxqKr0t+32nDFh
5f7Ae5coWgU1Th6OZKRWc05l81PYJtOkW+xu+nFcfhGitbEk6BLeIGrDSu/9oM+S
ZT14GUiS6Ks7vMfOApHT53wlINp7O9C63scvcMaFxDyGlS8IbRGqFwNiEzg6cU4Q
jrWCEpTx23HaH6VF4U0B/RIaYxxMutxKOCYAnTMhj2vlpVFQFLAN2UcdOVSaCWSM
OrRbit9xjWjhl3a7iRbwqcYUvv1fXUNuiGGb4V40CuYpkvatd5M0naPx3aQq51U7
KSRd6qQeD89gX36XCQI3GgHpe9nrx52d6+vIMZKiIHbmpIiI+OyP9D8Iv0ctjqw3
rGYBhraWL2vVefX9DCxbV3lE8qNyjyek3HPpw+pxZCnTvIE8k3vY0t8VDt2rsH29
VH2SYjrzaOHGOdQqF6ZskcLttYiIDJ0ECnytQRwQmGtkg1JM4Vn+WwANR2oUdxFJ
qlMmbIQTGw92fxPJTtkXWt71IoIvOIKNdO70G8MaLZVPXYlhjeb+mG7zfvBbpLwY
AejnCWqK6bGvY2mwetyP6BpuVhmGJesqXGVAj8v9PLYC4EUyrGmBIYP9A1P4FCHL
o0s8eiOrZHDCu6nxeD6jaa7cVN2ckD4OhFKzZ55VL6MKzrdbzhZjBqJELJbmv6Kc
N9uOqMuPzMTK7JSbmeop+RYWjz3VIB/SiH4uTmd+MBVUpEENHmMUrhi1VdHs3a7B
p/DtCxXash0m5mupzv9HjFP5XL4by8mOHndJqifkuH7T9nRrtsj6i8K3O+hRGuDL
dDDq/ibeRZpiLLoC8mubwrOmLKI2G17tdo1TIo4JdAzi4Ug/HfBNpEtyoF08sAj1
8caErXl7p16PU/0LLpoU4Cb16oV78cl5IgFgDMetcNOK6UPzPewpoHPsdu6RnnUA
wIbgL1M8G/0F/ZsHIfZB5wOQCw+OfZks+PRwE6nFElOL7yUD0JgZct041htMe/OA
a6WH7kppxcHWVxdTh/pvuu4wNxh9A3OOs+pxcSAXnwfL/kxggtuo7kLbxdqnc3Pm
4s1d9sAC9j8WxMyTYbZcwukyGD8i/pOlo/HrcXU7IGbybaQE1IayuKP0pjNxI3Vx
9NVedLMpwNyzI2d60npefwVhWAduRgb3o0pnUU8waKkciKE2FbIXaQn+1H06cY1N
8xZxBb61K6jdlHJbPHG/w/1OxNa4+TXPkmtZucVOLRhFunLP+2IVzvIB+6AK4qfg
EEo4479uRU1T9PrcqiTQupQo3BCKvY2mu9RRXCsBE42XRWAzf+cV3jPigZ93m+ei
v/tEjgYM68HZiv4GOjjMseiRjSQEDM2rEFayPx97U8fw+8BHyp7fLm0Ml3edKsKU
lG1V/+pSGcZ7VsBgd41Mfc6g4o9MefaL3vn6RtYUdmh0JkCP+ak6ijw3bbadQCE+
IGegEbN+1ePfn/qJSyGkhvsZEBhdlcCr4iUsDOOdF+o4bpykfp9V+THrTwROBp5a
1/Hu+xXMDcJTwekYuctPxkgUibcvl6l/xQpXfTM+b9iOSiZoFpRwXZj+b1PY3Doi
PfkQc6vzwnm8c/NTw6zjbivInRqnc+BRWvc+GZLCLTKfHv+PqwrbVXBE/ojfijSc
tiZyXD7oBgicc1+dbi9b1X8oKjyocAwmUq+UKftY9c0Dg+4SmDQKU9207lQD6uRU
FvTthflSlBlWK+6gYpUJZKSj/B/29gsCImMmrxKde18auPHgEKALvHvK9PDZ3VEC
6u8AXuW0W3Rh3FFLfwBWqNjSbxjyD3o97ac+XKXGRhfW559qNRBQ1Evf057b7hsZ
OUia4wPKAnd367uzhhv1IpVuqWYfYnU/ZoO2dH4b2CqBx8C3HQ5vF9o1tYlxIXaz
DWZbNAW8NzlchjHBsA6MJH8el4pW8vfgf4CiOY1LBGnicIztaLKXhWkWTFkcKbLr
UII2NEvWwgfrw5nKYowca1fvHHvmImg6zmM4oUxuvMTHblrD41UhfmvrYEgXXHT8
1XpCA9l3hdD7edpy4cdWx0880EbBJTuqZYQXnAJ2n/iEjXvkVwI0MBiNQQgtLIYM
YqHHJAca6OoMIPZcnfQOtEyC0j+yWzRZBwyC/ZucLltyAsI1rIylP4Uv7SJKoKfb
e1fb5NAkdPry8WzaEDXiC85+aPSxqbdnTjD2/4sWlkTB7NJ8dQWOce5Z8zCDXIEP
7qYURC75nELIiscrv3ItFhkE1GXjeWGdX6gDQSZM9t990dt70pcFdNy0Uo7qLjln
6/6I/GhP9wHA2gNrdi9ebdFFZGDAgoDqZnWybZ2CESXNLrnoL2orRNqJuKB4gpVu
f+n53GEcHVwGh3Pa3xbiwN/4OcngDzr6ltlwYyDw0+p6gMsYNu3gS/pXCoks7CpD
1mC5hVoKSZ80hVysUxO4glYC0M4cSpusQP46oY4EFK0QulCuzTgWphz3jdVzUCGV
BuJjs8a8hMuVZSjCmI7AbPKL6CB/a9zXBgkmDQ9xuzVJGURvd4qv/WIm9Ld4wLCq
Ww2lmVxQ9lgTrx3FlyTYbkLyRniN1GyfyKiCo7JH7GJ94QXqtkWW9OdV833mvNdS
qZ711U/2BuqH4oTCxUPXRXVzcMcvPtmfUDE7E1iI++mPAVxX6nVFFeJXSG1u9GDl
fkK9Pd6idWb/khPO+hKDySsHU3hA7vOw3KOKDIUMqUxpeo0fo0gXKQlsWMRNMUEV
djQD8u4BfJKES67hsH1gKx0U+y8NYyH6wkjxV6vfLGjeLq1/vcQa18OPtnFp3wbb
wSyuLDSfyzTjKuBSEPQMuo+O9UXCZPYlWZamco+81UxkeZ+M0F0cWTNqxPPUk/NW
Ep7mLdwuUg5/1SB+D85xD6cSdIUO8NsOl2/0XiAJKiOLBBBRgxlWLn8yFttrOuyD
Xa1+rzdVzt9weh1o2uGRg3md31FR5Po1F4Qi+M90tCoJQUMz1OwtQ560IGYlMH8o
c1BHl0yDfzbyZPpIvhubUWq0gO8vZSeJ0UKwj2Efw/G4LPXu4Hda7vpK8TwAN/1+
bAY4fTsmCnPYeEj/8ewvhps6LnAd2BmCob6sc41vNMwu3B7E/0vaP8TLcCd2YrgJ
/Eo2N4W1hzx3ZDGQOuZVMhVo73Qskh4PgkUlP5qSOkrn/6UC86u6jz3hZP3V1sDL
5YPGCHyVz82akHTr3SNS3LT9v1EHeXEznjRgwmd0TzPMGsnJnzWsaEuxo/QGIREw
XpC5hqglC1mo+MOmQOb88H4XoPXMC4kA2CwcJzd8A5y/qxLZCZbRkhDm66p8mtir
Y3WATvFWxA3Tc6KN4hrelsM+ltNIpWKC415JmC2pqamQ5V9HEP77SS7L6a5g275a
dqNBfcP6WCPMjD2LGQtsrsnyvqUb/QVdBto8k1Jn5j/Cw5WLxdJiSQOf7qO/UEsI
DCL591xEbS68YHoHJkS7aIOE1I/5Ye9ZCnuH9wVxCwDzB09qPLnE91GnnnZIsNPX
7WYV61aP1+7tREhfkX3GuFgufmS4c7QhYqQT/7kNSKkvMMBXLVC7raTsWOhDgTj9
bZK6rpei2TrgXQ9NyxmcoynxhjwjBxG4BSpyUZgo1SM1UeQ8n4vfKHq/j24/lDcE
sYyQjuvI3FnjvpUP8Qt2g+n9/GFLJEYhHJUSNxES7NPM934LFyfJ6VgLsnO3ikKg
2UVj+sH652Yw622/y5fS1chXH4v9kuTzE45jMWoH5isLk1GAp7gRrVAFtB0eWx5H
FMViImGhvrZWmGyHWhoXxl4Ifeiep8RUgr29UI6oayc6b/dGZwxQWhOqgqKnhtsb
yJKRMUfbZYwMTanndnijvRXCX1EpIZRYPh7eKIp8q2kBeqX+54Mvm4GiLdnw+drP
MUyq95ZCCzTqWTZd85OCeYgr65czRmlo8S3e07e5XdNyv18SAauDRFlPwWqQJFR0
c7ED5P/OSrKN4PanNL1q33ZCPZgX3QYliyDJnBiAwzJ7NpjfOiOyn/FMILjWqd7a
gEXqjIIRaWdusiq0mSgVBAXNsqZKd+0ydfM78FT4vic+IjV0b8WY19nG444IQlAs
CLqNXcfjV9zpiwciyk4wcuWRDfH3VZlHB/2hhqwpNHNs1L7/C7bGhBp2BdEamZZ6
eMGSgCUNtQWFg02D9SjLb6LTzZKlllpm/hy+jtKi0d6Z1rWplnQmWXFGFEr/xfnX
6z6Hldy+yEDmuDzjWVC6yXFeLRIV/nRljatpU06tlnFrwCuP93yN5gwAt1XPwDZe
0D8D9O5aP7jfm7i+TVBr/VLSyN5yolDJ31CgJLOiR9QCkIq4iDtzWkfsjVR7g9rF
aNicu2ido4Ec1nkKuMt1zXH91EgK6bJSsxgln9Rr5uXvrdm4PbB3/iJ6u9jY2AwE
y/+chTCVwnB47qSx7kXimoB3Mg2H8iStfOKx8yupvjYm0go6llPXcdjWEL4zLDkh
w+ySuljWjZANCXXF+ikCyisY2xlpNUtK7q91IIeLJyTHPvBQZ1FyILiRnZVC6BTQ
xMMR97nu4yalpOASZU2uHzHX2xX/i/aasFiJoBJZU0V5dm2/GlWcLwLsSdSlk9fn
YxVqwytCHYVLrLUqJuECJcu8EzZZpQ7KPMbcpHIWTEAqGc3EEcYxRBxxXkuUq3M/
rLufNHZKHW6+MaLkcM5UkbKqxxcrfbU3EKneawThTwJgq7iVzM3huUK5RqlACcmf
9VWl3hGo6aVnmy501murhJKtJ73YQUPSzI48ER7jEdp5ONvRuU81UEkdmMD+NcSp
VtolgOYXEi0wPGiqoOixyVNvPWXsIFk3aEQkdWdvcUf36qcVZ5eK30DJNBMdneQ2
WC9mfrjTE2B9rxbUCey3LtocdDF/Rbd5sCytj1gHpvpt81pdb3+/W/8YuUmZ4hJV
pVq19XlIuFL5PjDl9Rlq9z0lEjD4xV7zlZ2T763E6xIeDgG9aiQ3NrsDDXMbYcTG
wke0RCa4fz1uR5LvXCGD51dl5AKaFDciHYE5VJQdMJSZaiogt/7ZwIsgBKU308O4
cYK18tEyZI1VL3B/hEAsPutepNJXS9IeMzL95tGOamLk9Syu3grXhvnsmkUr0Ji/
EBf8JmebBC+0/j9PztRYoN/xNkYAna91UFMCf93qCRciLSJ6sNEZvyNBG20PME3z
dCrOX6YHOzL8RW1Z1WnbL2my0gEIeZnI6SQrGU+1yhx0Lo4pRwxQzQHn8vY8xkwK
AsfUSLh58WWH59nhmC8c37a16pcBSUz9O8W8Ziq8IgLDCPVmZpWywDfY5QF4Se/M
iseLI6Lt81hyH7VzZGhPlt+/PXJ0rzS/OJ8xxPAG+vuDf2QVEd3D0CCi3b6QE5Zi
MtOEvlLzKMU5cSY9JVsS6NoAHN+syZfCNSUATSBRrgDYZOOorBmCSMWUHGCioWwY
xNrGbI3+R/+97SGEv2k64RV+XIZeDoik49Iop38Bj0XljylgfQSKuNKTAomlzm6u
9PNg5uRUWGUgNIdisneWFmmRa9fLJ3JoPyJLQR1TE18t45XAK2DcXlwOeQoeynoh
KZnZaG+eY1QBV+bYzRY/BGEaJeXJbXydAbszOg6J6TNBdsX8rKkbKSbt+s3/uXl2
VuQS+DgnArvnMdchV1XhfTOtNv1jLIFhu8xYrKyLo74lOVXra7etMvHAgz5RflCP
dVYE3MTXr+fIzzhBzCFCW66SqC5fM/UIdNnpRmtRupRe+GASOxF3quHMMSy4Xl5n
rx2QyUtIIQND1mFWS8ycXfYbTbCSq2RDOlD6TUelkeh+tj3ax+eeGE7c/tK1yJbn
cCTx4MkaV0N7DQxR01ju5LEgEiVIhG+nSN11de35Shpd7kuaFlMpWsYWeZWnsAz8
GSiRbMpwTyQlAH91SkqU+pJkz4OZyXfxUesnlndj4255+09tsr9MakbDTYxgc1M2
LFfenak7thrYSDS+iDcrkmQ9pSgDc1zQzoyk3glOBVrW6cwW65hogIcy4sgzVOVZ
+JqKl3cpZHqqGdld28tTkhAwvyHcuEANcwPCE6yWMrOvr2JbW7M54gzsFqbB/wUs
u+8GCn6+W/YW+qAkq/tpb/vWoNwhdjWrUAARKqd/aWcjGydiI8AytG7z8qHytR3p
L27o5jEjZjhUzaXdEGb2wqQblLreAsos6Dt4gNBj626Pb0CI8UbKelx8WWdDmycB
iBym1pfeui2tKYupvr4Mds5fqpOEAneNl3BjYayEhtsE5lKh5fNy80cfgC3sDE2A
OFrnEAI8k9Nv8kZpCiQW35xFymcVdLrOw1a1cMvBCz2AWJ9eZPVGfAk6SpBi6i66
/MrskPCenC68r5AmszdcbADpKnCQGArtiL5QYh5gyWBf+6aLpdHt84lkWztMh85j
KTaPwoVTnZzHhOIHgP8zu7P4xtyVj+bD31kgUmy8JZyIg+5EnTvAXQSvMllL+9q4
cNd77cCl9wHYySPDE/Z5VB8ypihV+CzfeNhcp/yC7Q9TTq8lCBdgVr240O7hel0k
FCLMkZAWAo3UA9PVsaMQDFzWVlgld1+iEAXroGVrtUoiVptKJfXQlJ/CDtjxOhvK
7ynCk5wjZBB5mHRVDVgvzQrrQRrqzl44vU/Y29ZpqRgg/AkoIW+I+YIrYlu71m6b
yRg3DNOMKmXi8ssjm0+msQ7+xe1869oDRq5bu1k0ibgb94Osqug/hUbGPoMDMT/r
7xP6V7aMG7OMOSrN3Fv0XCXXMbLJX4v66GT4HjqTxXQUK325WLWS4f4BpL/t6KvV
OGZc6RKIjkVwcw16Ap2PVXTGVk3+xza6rUbAKl2/JBvlzDVEbrqPUYQg+TENCMr5
aKO9BHtAZR4IXv6k33DU52onu787HJwfvcB1F2FLKtum94qDPMZ3HLFqfnhPREJ+
Cs2X5aJ26U/WgRq1icVetsa68lYXbD2x1BMnkg3OErJ+tr/se2gt3eh3PcZ9QZ2V
lzru2mCtbTEqo9pHpHzrI83PAd394ZmsgtrH7yS+s7iZ23sJZgKKc550icOduGpb
TxVQo+jqiWSEQbv1yxroHQS1gB7k93o587rGBN1m+yXyMoi38QXL9RMcriCjdK3J
+NaFJo7TtAXOh856SqWMUgEf/VLVZCkcX5Q9XA8nC+kiHt9fZE+C+bYaYZDmnTgJ
X1MzfgkiNQfC0CjvMVvaIeNcRktlyG0LmzHFs68BFcVf2I9L+a8DC6xgFan/1PtV
bg4K2b5vw5Pq5zLLW0euRHQaAIRp6fLkQElpScpWZ68yy3GRbQxsNBnIct4Cjwgl
Nq8ZYUvZiMy9iUfQOAKXoqF4O7K9cvUbHy9GLkw3TSJDx+QjkBZ9JYYmWMkPG90z
3Pvh8l+iHZ3WhOPb6pBo4QJul6BYqaquE1dvftxTUjg+pyoTCK0W2Vrk1lLOaEqN
erG9cjjerVviOh6GPC+E5+o+J2S/kT1ym1PMtmoji7RUsxl+RlMiqpo+SV9xIHgS
MaPm5dJcLk3i6AVZo6NcGCwa7YGwLSnS2plNaBch5FYsnd60Bx8c7nT3/DeauU/o
8cogsn/uKdn50y0n80+NxOgUyjF9LjyQYsY3QWEdqv+bIJLBEAi/746AGJG3QsWL
92Z2vl+LN26nCkURJjqi/zOz3oMcfRG+oYreQtp0osuL6BFdkiAfTGjorRjaapmT
AllJy2lWjgLmpnw/krRsn0hkhkg5VZ46EmkEBw8vGMfFo3BDO431SSW/D2skPUX1
/7DxwMcHhb43BcmxQY/eC3mgCIN2cy/hct63ecrosm4orndxsH/yDFn1ruJIvYvv
OnCd5AwCBUD97FLn4uiYdyPM/a0xJwbSa/ewV8Fgt1+QlziD60rrgGA3/Ekk7nC5
iNhfowFJY/raIaTilybKiK1MMb5ZLy7rA7QO00+4RT5Few9CcvL6SdtDpAY74Ntl
yaKcm3PM9K4madY8QdT6yjYOiH7RfnuP6kXzIeMDVCgbxuSnq2XvSj3lSu55PNCi
nXEdm4TbzKJA+EBwGMV/dGzAvYg6+JH4e/Ho7lEfO3j9MYHhFMjzSK5wOhuqjKdA
lLPJLuPMcZeuuhiazRDbHYu5CcegYi9cogHa+X2RK/2qdazcnL+9aKJf8x3QXFA/
wEotS1f4dsgtUEikJ2K3P0SFIevVcHcA09NKovclmFKoX2MQBIEgmw8zuwOLhyzO
0ShsGZZOPtksevuXgcCiwCM2Je3lKihrFq4oo4j33liFdt/D452eO4IWj4R9WwsO
LlMurNxCBUH+F9TVwKyc4RdvN+PTMuc6L27A8B3ztXA2dxdATILBxKG+EFmnUa5U
6g0XzWKi87K/U+lqWuxC9Y6e+VYZ7x1H7HnztyY7Ky8vWkRy2/bzAr7wQ1uFnzq/
IUtCU+ifJfvWuoDborFiIgq0ZZykPy4pky63tmX9JAXysNum4H9tk7plbwocW4aR
04mM5g0ir1EPBGHPU/G7m7LAiZt2UulmVIqY1u7LWIsc7szkWPvu4A2p0NPrbDj4
0r+nvzEfmaYAVPPtEOsSCkVNPiYMreLN6U/Z+D9D9i18ZTlrLwa/HZ71jqGHOqTv
k54gFewM0kFNk40ij3V+SlSe+MVGwfnjbu5sjGE4FDhI3eFfLMERYgD0vscxCmUz
7YmY1kcBg2Pi5tBSsSxeQ5tk5FjC3k0zaYFh0HK+pw9Dv75xfBVQeWPCbyaEVeto
5llvFqOxB0mJAXEPOaIHVtAVNAjB9RKODzIWEXTcnMXJAY0o47ArAAzJy0DavkBo
gpg77QdwTb5RM4mR0QC5tD1omPy/XJAI/DVq43jVvIofr9QngI5Z13uHXAlLZ8l5
nIiVeTYyTeUS7YRB9v3osSleYq/9dl1iDSPsnAWyKJ+vARPgGFIwnHgvI6oa3USQ
1e8PFXa4TVAkpb4JPfwC3dE7p5maF2WwAJTCnoV6Hz2jJwgWmPfc46DokFWH7K2O
T9kvcx7qUTYR+7qFBcDSyL2RGagz36TPnLaCOQA3KdZRzwTAq7WF/VKauVrL24Eu
0MqqBTYLRCq/+sBc0P216ugWY7n/ExN5w8xq1ZgfyQ4a5DnxjlxdiHURO8TVnpWU
jbbr2Qg34gx1uMMefimZQKQBgtia+XSmt5uaEijUrnGx7DARBtEpgUnCSmDQ5al4
AjUSiFd1vUB2CwKAumcoWMCq+Q+hH3coBUqD1PkR/tzQ7iw29wYNGY7rh3ARv5Js
O1ITZXdPZh3u7g31aGxd1124rUfbhTA6Fip9eeX3AhLCG2zUUz7nKiCrYmZXMPwu
OUuTW2QhCaEZYX5eN7HRnYoUUwkrQ1vkMeeeJ127jKIBYCUWlL8tWYOoTqj5smh1
/UzwLvLrp0DegNMxc4kyx5OmADjOl4li+kR5L8BP9BnH9sl2JORf0YRwJB296DQN
swk84eCb5aupg2M6gzvU2qMDZWiRo7UCqXEpKMe3UDORiFHzTqtgbg+ugCm+vteo
3DDMIyMe/GRSpvZwHs/50+ZrQ5YeQCXPffe/+pVt561GFZMTDme9h2ACmbI+ddIG
/r3UUiz13+36VNHG4muCLCdtTf9UZQtidUgtBr7BjyYHQVwxyKgjwLbvX2YydNLy
juR6YStRJ1B/LRsIa56E84BVaxvh8sw+3EB27DEdTJqBpOke7yO0YfsxgJQxczwV
gwKS2eRB/CiFgUNdm32HFf2OUlAFzJTFJhWF0M2Ko7vo5mpui4fd3x0IETISNwQh
oX5OUl4rDWO9KfDz6iuUJz7JpMsdcnombOmvymIGiUPGnRLl95HZ7eZnygdHDkC6
8/nXGSM7dtN21l1oxds3JzIJgqPJfseI3GBxniLe2Ru7cPoiDrggUL1ux8fJPDaR
yKKxiji4OmJ7FN6EBfJIkJKUsl+Os47hZ4OgQ0id3qIxWpTpZTcRCrTdP/sIcy+Z
LOF2sLAnEXvMLkMtdD3p1qIyXeq9F13a7tRvPsZHQMhUI8tz2JTikEAbBTJMB67i
DKYbyc9v1UJQl5GVRaWYoyUzvBUhbLwMFaIx5D80gtH3ShE/GxqUdyIE6fYV3a+/
VvDppIGDQmx9lMtaUtEQ7SgNzyJxf0p+jR1O02bA3Wj/REe1uNpFZ/IgdhlrFwnI
N+qkl9IOCliIyUxE4ejc04hrADthiu/tUf68SfF/lSqS3yZfUefemM4/HGJ3X5JS
L5oUcgvJLcqoJpAr7A1mP5dWhKHzo4Az11Sy2ZoGOxjsIWdspCnkvh4LGfQqjsnn
J9hl4ym1cQEHzmUDONqozZZK+W4Het1aCrrCShcejqlMIY96cA0Q5jonhldTOtkF
9Qj517ZdyQ+Binmc3qVxOz9i9dCnqDJD72FOPuanvrKshUpKpXGakv4MdWjqF7Gp
IuhWxO5biHFHUoz0M3D2cyX66EXPGL6jYwFYGvhgoseUyX8HxpF5uemCnTVTjbu4
sdVJ87i+ol74mXP0enI6bsA6Yr8N4EbQjjAdUv4BD1ZkOz4kobxCu6PbJUVt+fnx
H+3BP/I3GXc6Gs79GD9/YKwfL3yq2m0u2CXHeMrHus5qeRECm+1iZaeaFbC2QvUw
37nERvGR8Vp5yO76arBqLfBax1b08PHxw+oYGj8Jf3IL+h7kf8+NwcS4w9fgCco7
VIJB3iQNkI9x0q+Vrx3E8jKxDkSOj9q8Y9ggv0YsnItym09iScxVl4aZYsQ/H5Ie
X31DXvRF3U1Cz3EEHPVR4oobMLTo53oVPv+XW7xq5dboCtaaE9EGYB8OnyU1+ti/
3/g7JKxEi1s9TS5upeiINbcrozKlh4DI0JHIRn+EJRRA2GOA1BQdhhC6v1GVipVZ
mpHABGDEV+uHl/t5XUzwjWQ8RK96cq0bpihg8ApwAEX2K/205ZeS8s8N5YWvJGbN
hQY1zQIery9x1spt4JOxJ5ZVWTMndu9p9UJoP6p3Cc8M0QL7Q5PGXFk+eDTYNhIb
d+TwzuOdWSYcUsTW1jdeIp7lJqTGXuOe9ulFpPvkVg4yUb95KxCchZQxED3uQxR1
ndB9xx9wUn9NJgFSux4UGWV8yxeb5EnsojxFrBIj9ah62F6jREVKfsSeprjzSDwJ
kLMecDtC6/VvdEPnNDeSflPsJ3TpBo0fFg906pDn389xtdETWpwDSiM5Dj814u3v
qMqXhUQglBqZKEXaDQIn5/5nAt3bIIQjzv3d7sheT8mP2JVv7Jms+H9QSUAt8/Ax
r30gEQ7iFmI2LCbHVnpH5W4QVpwzuS3XiI5zSRWiOZVJOTx0Q/1+M15Haq9Uzafx
5l9iJMC5rkFcJWApasoQ0KkvFNXHhtyBUPVSWyyGCi3ijDFqkhCRoCAuGV1oQYp9
4iisEXvYHD/jqkP7V9xo9sUudHiUA27LKbJF711W9a25/A0BsFQ0A4Gk31xdPTqb
hE1fx+hgv9qPOR7ycOKcGsKR5dzGE3VCI0Bk8VE79LxQPNq0L7LMtvERu5wzikEo
D8xtpp0xi2WcJ5rVU6GMoZZe1axGa5OFWsnEHw/XfZiGi4cMFAYXPhRfVpG3XgHX
anJ/tp7H4xaBEMVW6rn6WJfahyYN5YHCKqrPmuAui4ooo450nWE20SUw8s1Pxfkh
LaNYVW0abtW333kpHbqWfA5lacOGDmLuJ3o+AiTX/qVih6HEmdEJSnBH6BYyIID4
BazewlB5uJw5vT15j9xJE7pG53lqXth+99VoDz42U8cKAyxzEC4XHjlvDSvREqxy
ti+08zYPw5Uxpp2q+xyjetKo6CjXBtxXzKoS4urPwyxDkdwrSEky9BdS1GuqCO9K
ragerqqpLFAKqEEx/xxTcmmmswUJDqhdxcqt0Rr7Y/CUiCqoyUInq3KGu6fiK3ny
U5xnCjBuZ9ZK2Vr3a30t9QHgxUgxk/XWofDsafzZ/B722EObq2Yr4/IL5WRNbxAt
IAfuiIwLtEDLYgs/fN26xNu0C/zsgygo9CBQ1axKEy+FJkXbCY2/eaiQy00IFREd
XZ0/XKR9yNkJGl+HzCGpFz15AlJpQuCVzFXrJIqEzO7HS5ThpElPcPgydEOBx1Ci
frLrOEJb2T2L8UG15okm4T1W7sRD8q7jgk2IAwVPF8gGNA8MLKqHxipox3G//L6X
IZ+0qzkDlYTR6wKlA0FjMjXJEZx7eiDtHor70MoIu3QpF9XORYIs0xFHHGZ9qtHo
7aNohvDfrUaOOeCCe5JWJSYqkfHP84B+lytvSIrerr5FFmYRmIKbs2AmrEtOY0rg
LnbjugcZ9hZY+XovXmLX2odVipqDelld0TQCRn3WRye7DQ8XvTpF4dBP92g571xE
Z6YwkXRRq9egLYJvuKLiISohqsDBMl2LXoYUHJ89AV6Fgjjq2RqLx2KeV4F5LwEM
Y0pLrCtyqcuwmxBL8jMqGgE2/s8+PPpkVbdLYN/+5YofK1DCYSvVfrm16H3xVC8Q
w52xLM6Pq2Ck3WuIIBMRwgEbcg3340iP+XY4wOjh3QGFSZXwtjTs0g5pSGSn0ZTg
cubs80RJCiwCZueRhWNn4+CMgvnLRTdE2Yp3LXRCv3V0QR9tLwZWM9taj+f3B4i/
asMlQiA8xjbX4o31Wc4N8rGv2RVszPaR4PxDZ1Y4emY5BOeyR9krksoxU1NjyC6f
Syfcm4/iYYjChxG4NJDLqOmpaTNPnzpvpvLJOY7P0Ge+fLIOK/vZhorJQ/Z3DrT7
ZIfG0lxIe9K+It7pQMKkN1PGgk0l1N38pPV5xiyZBuONjt1J+SFon8mTBsFGXICp
eAsmn9VZc9DPjeEv7g0Ier/h5iW5+rYOgALUzD6+qhhfvlNb31YZpXc7fX+ZOa+f
WbFQBZsnAZ/WZEWBRjnxtoMwd5+6jtdvWpZ7cgYucCAhk1SqhGSHKCRM63KBBSZz
wOuE+ujP4v7WaxKpf2XPzrdlFmMiYb7lVpuZjrRnJcOskjF+Umrl/XpYurmJzePy
M578qz3IK5njbX3ND+Ywm5ytOFwi6qy6KgXcHZzqMLrfQAxGceNrxQ+H3ojUNYYj
UC6M70TcMpl/LoUbSMsl9uZCwaWnTfK2XvBAdqPfAfi4yqSXkxwApCTQhn5Qa4Kg
COaHpKTgSjxJ0Vi+etKZ9GJ2pEQAlTeSxfB69PbP8XaU92hQ8Sg8exUQow3PrKY/
VFYGHWvD50VdWLGBPln1kSp+rq1jCRV/KjfBp/CDI3xmrCRY9eOJYJHJhE/Q6ghw
uD8D/kiebYRRC47td3ML9SU5ogwu3DmsgTgRcQ2+eM4dUPPTM3WVZxTcunEWyKQB
7Zjenb+Xhi01QUBzzV8qg1DFM1brxcDvXiajzMrzgRv5UVflJfE+SeLH+PFM/jwR
kHW16wZrv3IU4lMUiQR8zIydKqmTgzHsUzgFSiQUxmkNZWPt0B1lCdI5XmDayY37
yQdhVtBZXXK1RlYUNaFIzAfZhIdIyJ9AtqhF3WhTPOT9AzgI21WLm3wQ8jN7bmqh
YogmiT2NS7B3+u4ce5SnYeMwoH7Onigta5L1BHagBAY5DgRkXtOQAwzUEQsI2EiL
RxYa5kUJL1qVGIDg75H66ITzbciI3LuB/huqIiFEamQu83JBhHhy1mlJ0rorMr4Y
N20qzDSPxBVZVtizOPs0oij3pZy+HWp7xxuUJzWv3C7x+t44BmA3NUqXkwkuQHZ5
1540v07mIp6FpA64v2Og+DaOMuQo2rBAyjpUhXdkA/pjPNRAsAVqB7YgkpMVznOd
6Xoj7taNmAI+ETAz9v2dycGfnVWzGNIyxZt16JKM/5BSmUMPOMkzyCh1xfMDvCgj
x7xmOV39ndTqdLJxYE9Eihei418sSmM/cYNLmRo0bin9bhdwYTz8I/NhJ0qE8+hd
J7QLdrKgGdJhnmsn62YEHlvtUtutAS1peqTbHrnH7V5bx+iHKtgvebQ92JFnwU0q
+jhHkjQBjD5pRlhwcb+hFNNeZugqxoH+Lt9rHK4FTKxFwWV6PPHheiSg/uN8wyQK
WCsQR+00Um1cxJcPz8QFT4BdGRwSaJn1F9gS6Qngd2V9TJc6tD6AmK+HtsER9sxa
RGHpOp1UF2WxPDUeX7xpMa2e1yqnm0TNA1ugHym6TJNz5K3dVx2BwrLnzxg/1kII
3HALpTYCeCkfeVbf4hMT2bUjz7Vz+mRJQicUg0gwcObcRZmNeX7PPYAAlHfEJEnJ
qOUD1iXCaloFoRXUQCRkUoxzso1yQiKf2v+GP3jK0mfCawGrkI4t62yPTtjT8mH+
3NMypJ47laKIdYB7bhcXoG6XN52IDWD80lKPHjaVVE9PHhAXIKRHlSVIDJt6YNjV
dEzsuLfLftRj59q+41QP16Cu++RnRjGx2mNeIX+JT6/wvP8nDpibf3akj5XsZGee
qbpATzcSmMJGwTe3TizYNV9Mu3GpXxzfS6ESK0FBrBGg0+M2faT5XvKTvhvk3bQ3
VSGdkfR7D4+jPxKZ2vQYEkCx87y0ZSI3Ejq/PDL4pOu0tEy1Ti/VFkNMx1ze+P1c
sScLaxcXlWr3ijlkrMwAKahVmRDq02ovi+Yn4zR8Smm3Rsam2cISCvewkabkb2F/
j1IDfi4Iw/BGiMm3E/Qp/7VVIYCqIzZEtX7afLIK8aX+0DAy88AgEE401ZTbMVyF
cox68ZCE9FXhm05aovSBZf5sPqvUi1ZYlM0WJBczd/rjKnEYgS1DfyGdIIYrmdiy
ZOc2I5tv0fZf41U1UWTBYe3GQyHMk3jR4jPUvW+hpFI1nQUs+hLckLaKKeS9LEHI
arUFuUFfbFo7MWYgY/cmQEVhP3zHgPLSNucv65G8zP9eo1rvBUp7iKlGVrgnvPQ8
nia6TmKt0vuEePKQZfUtGCLK+1a8GEtGNgvbDn352lWYz9lKh3hp5hCNE3CmdOTy
/OcAe5mkJdXt/S2Ef0FCx/3x7CE3OBhbVhMTo8PSFDKfbY7iqqmtGmaNmOcyQH53
6yRy371LYzUZkMLIurJddJ/CGKg7Bl4Jj+wdyzumdG9Hsza0DNosflvE9/KdN0gQ
pOZGUKN33v5cpnTwmRPpDgAiKGdbpAn+b3fKku0FIWc16i2Vo0ktYRUR1w+Litut
qPVG3XLlaNfTvsAGIc0ej5TOwyCqcFsF3XOtQtr5Wl4y4/auT440AqER3piu0Uqh
ivee28GJwgm3/+7P6qDN76CrjbUbCqrgsegaQ29s5oCavNEM7x/Af5E6zkGitDvB
ZCIXuets/W60oEqQ10yDWRYJLzyAcMd9Hz7M8DrDe2MLwLBmM3mtZcPONGWYzSQD
hgIUvNeDYa7Fo8FWgJC+0aQTgzIFXAJkMePeJA03E/XuzFrWLPXv+SGwhkCTCAHd
aZTqo59V0AGC86W+BcbToyc2QKhG7+HgABo/ySdTw2aDGnyftljV/H7n9C2LD6T9
K+FSM/hRFOgujoLzeUMwiy4L19leLX7NWrWc/pSbG+XA6MTQQm2zWV/V9NFClbNQ
P43G+qbolyGDuJ2roK3DO7jkmH92Gl5EWexK1L66AO/yb443yvaYBZ55lI6o4KTT
YyVG+Bj328lbhF8nr0TfjjtgbQzWqHgXKOVsUOAi68SfKO0I0QY+2Fat1eup0wDa
aa4BIQzwaG5xRarDjSq6b1iyXpAZdq3lYd/Jb4SuMOk6fSGbWtspQwEg76MoqVvJ
JZNJSR/4wI2g+JD7RurUM3VVLkopk76rTJACj9Us4AdRgnCuk3hBQfe58kGM3nAL
wT7Dvw1x2RRHW5APbgVz8usXh7RQgGCjrdRl8bb7/xJrjUypZV797L8HrxKoSrGd
bwo09xx6ADePQtQ/499bv33uaCCJ5zIMk7QMdS3ruKHh19mH9LDhr7ko/e9sJ0wE
9ow7C2J0YmoTwBaC2b7LFPDqCaHMG4h6M5Z4ld9ccfQ93h6/t/UtYW+2ywDaZvoZ
ivLkKAEdqP0QUQXI258xgEwGqXUylUq3pFLPMzQ8srZI7IhvPvzumw/Kf7di5evc
+cXCIiO9u0VMtw6CLfqSGnFdNRd6qHJ3ozjRCi/10KwoUy/05fPpE9XIksbSDqET
XlDOKpkqD5BV7xEEetcHGAsLjH+ygiZG9xPS2xEI/MrUZZuejv0gUxARQOZ4uSnw
OgWZmO2cqt4IEESWaSbU/Kfyj+xj0IOUc2ignlQ92/74GRBitsPVix61AsXOtb3e
lhagpwJeGVoWUkIQ6+3eysGP3FkCTyDvLf0jQaYVD90F06P9xFzdU+/lTUmiuKHL
yFLur2cySmmAIvT7VITDxoRWQ2X3V3TxR+D/doRUeMkt39suUpbvpEDqxt84BlqN
Nv3bb8ioCpGmsTk3cBEE4xhHiwMaXhBRuQnwdEL//Aw2NRbnR6CoqNcrgQvHEVOv
vIUcdSRq/fnfsKFJ6KPtF6TqHbZmbmXVHIRstCOpYDz/UN5syKJn/cNFwu+UHiRm
sGgzyXKEHRM53q/obEPnZVUptNQt+3RGXJ1Vy5khUca8ZwJi6jYHyiqiKPevIoha
fHYwBJZLagP8uMYHbVtNAs5sytVvUjPjQEA7pNRpnLJ9nJedL1Q6XklCKRixlEHj
oBLKgByyCnYC2V0hKqTXyLwqBLPtwFPen/wYyV+RrwEkYJSjm6EQTAVI/NiQHQeO
Ji8sBYqLvQOudmSKlcB33/MmyVBTqQnXrBeUFE6iFtANaiRyHJamQnw04ie8p0Ct
NUlRXl7njrIM3TTVeqbgHdNDQlnv7SOUDDyEhhV0CxjQh4/hx6+2bZ5JUsISsoQV
wmQvwC1pGd+SU1KPb50G+0NEX41/v2bMdnfY/p2zanow5GESO8p6zfM9OI3d6Pr9
jq0va90IbMjAurNUzKhrGqZK+ZoCzi7wl7NUm8fAck6vG+/SRWx2vJHVcbq62B0k
Hpkllm+onCzvFhE+LPqJi0QIXjpNDhhPm5AsOmLLc5VXa3x6MQDkuMfK66PF1qJe
MviaC2FTGC+4WfeKxBAMe5ymq+GmF1iqb336MTL4WhZ1fXrd2ItbPQOYz29akB7u
UP53nwakIMpheKr9lwK8nITpvC3tXelK89uh+zh+GFJpRMqjUHNPoORF9jZAcnwg
vhMb21P9aUiHfjdXocMvj1oI8E8y0AfAUb1WLTT6HflySIG29PkCrVmMewVgJrZV
w9st7IWMK/S8VAKzJPtvTeMfBrEBwVqONh5yx1OehaTdPuyb919LhuVniZh1Oijf
vQdKPwMgRLu8pfRiLhhpzZCNO5MNsTCoifyJtmnA2v1l4F++miizPmEpJw9rtoj0
h9rNkPDIj4qAdTWkn8jTeV3HnHOEwicwx36ZUjbZjflxb5FHe1+p2L9qqzdALhZp
5+xY3dqt0dsyjWWU6vzqjUkp+KZNWB1v3lh0A6EgmBY5/JmWzUSsdcW3YJG5X3I7
PYZbISbdntCK1p5b7kbHJIeqlIlSt9MYhJ6IXP7/eq6IBm5yGmVZ2RM8TUc91JiW
NZOj0aJi6lUb8IDEO1WzE3SSnmVEFgVqdAQrLtDuekbrz21PgH8q1GTG9+/MPE2+
n3Kr3UxMEookGuILZOLVh20R3z+c01eZQHYuqsqpfmJe0pVbsZn/BY6dFSrGxGc2
oBSgZQZvcPsDVErK2xUyftrJbi71YDGqMQ9R22aT/pE4mhmRlWIuTXkfwxhkHW5x
m8fuonAJw3F607SQJoHxAs1UFX9vBqVlyXuusyqOXqwON0YkM3xBBlwGnsRL9MMV
6YNPov8l1zOEt2IhxkaxM0qTblrGElybcnh8UTTNEk+NEQcB2NmubttX3dVSEX4B
/wo4Bj0QRgJpanGHWYniuZ+LdnJ1Mj9KMqOfX8pWcxZQwsedJVoL30TIOkZfxXK9
f74hDnq30LdFg+lZMQvSkN5F2j49+QNKWZcx+GC5C7YEIgrmGUvyusBOO7OSkJFi
i0N0Tsal7R16b47x+psogQtsxRVnz2UkDJN5tNReF9NhTrKY1FLAwPxp0zBnXxsQ
Xkj8IhmOboZXTAqX/epSEolQE0gR7cZjldN40Vs9Uh5i6m1TB+y5i6+vJBzvxTGD
bRXIcK0o4hZvLrrx5esoIzipQyOMJm48jw6h6O0Wh0Y+iNW2wiNzySwVZgFJ5baS
07zA+LgBTVwWHjTLDTWnDBsq+YTLv4yZoUYkoXUfXfCMerRE6D81dcrLVCiHfu5U
CLH6oV0s2n7rciNByTtahOodEH0zwx7gC3CAD8tzs2Us9xs7dQrYp62hZYZPz6I3
yfTgrckJNGV4GXC9KMmYFWYuKIFHryxufqisL9TmmNW8bV2tAGKYWOVyio4pxye7
rnYv1sOET/BQ3BTYG1xIsJMCUDFp/rROrikGMAFyfziOka/YFiCYM7UQ54ziuKBf
YWrQ78Qczq5dM7MMSniS8ECfdVrkGVDAESRDtxlYSZwnmmyYjDIRfxtLn1KA0yLN
OcXt6gPCukmAkYfjgwmsmseQPW5r4T1/3UcuuyxduGgrQQ8RLnz0GzMRXFu/KTK+
gxw1ZV3v7ZGL8Rv6ICytSPGj1/GVMhartxgCZGeAsW/yxBadUev6WmugInL335y4
mQCEoKW7eIjkBXL3DSuyb1cV1nMmJt0LrT4tncDhf//DtGFLrHYreqjPhmBW6X10
vMvUCMz4ujC9kV6+Y6DByRFYuFgKSnZ7Ue0aeJKNsSuXhW/tz+EODMTPgHklyhpN
YjXQYbfK98tSkkFSmEpOfQp4QDx9q7EGPBIrzRrRMO9Wj9dc913ZjX2yUHfi5A+i
Eu8b1+msD86fJKKepszQpwYCRCkBLVAz22da/lxBRhgs8rcjYGfv/50ewhZ5WsTh
2BZFSVkSNb3DtAvVhErC6CUxInw4HyNIpGumPkf0prrCCtze1hGFe9rQLKRvyxXj
AKC04FdlFF5Rc5XsM6utrEhOej+qp2os206C75AWlvTzka/a1V9g5d0enU1uVEDe
DowGpw1qjZ9GVcvoK1M7czPDQMs0hRxVZ06NcR0/hBzgNK3O4snOwp0o66QFYYM5
FrXPGC+hxWmQVsnyt23I1XZu33OLIChVsbk5ZbFBRuK12FzufTqlMoG+w4xQKLex
mf4bU1JqdIqLmIC6WIwG8rz2r+MUoJZZHBAi5zBAUYsym2r75V5yczor4kTR9Nvv
hw/WWfOJYEZfEF3EW83cpYSWbSwdoLmnUr+O4P85tZ31YtIAIttmVhhZHrADb7yT
w/4AHJqKsYIUX9bbKhdlg7Z0q48EeKToMvZN8A21m2d1oP48hCi1ohVWwXZGBoGy
UCyFK0DtLLKOwsC6S9v+vpL1z98g80ODgOJGB+cpHBoNlyPSb7dSn5JRRQOPYas8
kSacvb0RG2rRGOH9ynbrKJd1s86FRJhPLy/kwMBIrYcUXUDcCXYsQ8sxGiVNbBcw
m3wMm4M2q9D1OgnFZA1m86pJp5d9fkJUHAKwey/ez5TbX5MeqmdoatL8SUZmrUS3
mL9w1uyJoYUDVf924s25rEyn8VGyEveYEGy58oExV0oj0IByUMj08rFQPE9nct0h
kjIMIAYWyF9ZwVx7KpwmAQC7dMGQMYOx98vA4zq3Fi4mwUomM1RDPevnkXQLJBTT
wqze+Wtf1oeyaXlc12G5FvN7Lijo1SyM2pE7vFlac8DVcBUl8+ch89Pouuy4rSAe
gHLiJd4KC8jW6obsDgkwG6UybL0612bIedja7N2tEfpRzVqcwKzGUcLXDJ9FHzdf
CRqUIyH5skeEYntsaoSlZ2xejhFu91D0rqyvy2JPXZ8lJu/Q/7EjfWWMfCEoNQ9f
zXVu9hZrcudCzSny2K3HccmchP2TP0Cw/k/vrkccQcLRkKrUrZTTkhmCybxc4xBm
hg7U3h7Bsf/25Jk+TdKuQKuNncRtY9OoeImWfJzrRLlouJoSmVcOWYf8/dkjyGGc
5cpNzTu0QCnR+OQUZUvF/67K25zMcC7krqGXT5Peof66+HMOKqAdXUhEQj7E1t4B
CIwo1HyVnmckpPUJG5SJuZMutgiGX7pYojhBPrYs6aoINa/g6JSnjEDN9BuvShWR
F3CpAEbjbizhroVMUII+q82/H2bwPua170wR3gs1lr/2VVoOJ+8DupHEMfXmp1WE
SmwQhra+zsSUIBCzB9xqa7DQFZ8iLaVaAJxBwyASrMNw/Ny7pz52TYDDDYWo62bN
2tQTbF48Pg0iZvbLFHGxJuuaW7cP2n2wK5RGzu4zcDmkNZ1xJHNhW/1VKf3NVjif
b66/Tyob5RCBh2274qmF514/m6HmFGAwFVPK2WfYdM6knlSE4oULN5yBQD9r6aMv
tdw+NFZ+k0Rtx4oyipTXELOWcenLpVJnSOzm+MWpfZV8qAGlwcbc5Ami7CPcJSJz
8uC/V1AwgroVK4JMmDEiN4zI8KtXVsQXUt5/A5q4Q1pSue9pO1bRJQ+vX6Qw5QWP
zOTUDmPBKJ61JN4OveDH2JXe8M5/lHUVlQ4n0ruWljqIRYbPo93fONQm/eU6EYyW
PsG3rXzPvaf5wsS/ALtfY4JamWjEKba03TRpZ2ejpVzOj0X284Y/U+v7g48RRtsB
kO3WGDZR3c/13hvQCAc2I6+v171UiAkJZOvNNUjboVifd2X5gRI1PtgtfGjamElk
4pMEzakemX2VKk9uhrTfaOt9Ny/aBi8vPLaFQAl7asPXooWdTNd1mDO+eO6dw2r5
tZb0aA/VhN6g0y4gjCROs+IQR67y3+KGqeANnE6BEJE/ZL1aJpSo7RDfUbMH9W86
E/RCeIJmkwCiilm1ME6w5vJcHNV9ivm1IK31SaoxVrdFnkL/sSyEOp3622K6YZ/I
GgICXgZ89OWLXJcxzSQC/tewfgtOrwEbw/DjRYAmStULyA4PlF0gjvaDtPX25VE9
lFskzJAPpB716vBsOd6RPdjKs1jnYenJwQ/issw/4C3G3FN+7HSxpXQjE535h88T
DlK4stn6ogp0TmL7l8uqHLvrQ+vH99593xJzM+52GLDALdg1DTN59pczxxz2WY4W
4inDHr8vzy9Pq7l83yV67CTvp40OHmkjhlNh7WiGCSR8t9FZKXmp4OP5yfG6MM/0
eyJuMvFB6TkvGqxUeJG5ZPljDEVqvbWPzk9kWqw8L8gvm8T4rsu83xp+hK6Dr92M
/xr8PFUc4rX7QgbR0HmzKFOF1groEw7st3o9SjI7bmVx7wirDY71zSIRR20tM8i2
saqgTxzXin5SufU+QmCh4rPDY/zw9XopaDhvMcRRShgaMerwCuBLlE7gmGej2Ilk
wFyS9fQUA2B1z7yQO4sN3U0+ryRAeElkpU952T9GIvjLEoTuRj7ehW1N5sk77Q96
VASti9I7iW9Cgix2EqELvVkYdxQSlFsVHweyuiIQTsM479+y+FFe6kYiQW1MCa0M
a2w04vDYvh5RzCwU5slYY8SHitwheGKw1s79Lt72FdQvIiyu0roFTarVyR2+rMU1
BICB5Xsu2OVKuma05fP0ElutWhSKydARdQotl1lzKFxXl6Ry4DZbfVK4PVeHfT8x
EMheOvxSB5hG9ZJ6Gr6zE8QOD3802xoAi/TusHosA91hAgYNa3DdttkzRheS3xY2
Qdl8s4MNsZZZtlpgmgzETtvdiuk0TbJCYPxl9CwJnbjS2ASlfDRIMhQ+RGv36yyo
T8bJLQUwkThW2HwjTPpRycDuuPEZ5OFqnYasaNTbgmH8ZkL9gjzSq2+/GToGSmXc
ogM9uJXo2jv6j7eOHLxl7kxNXWO4JFLaTQO9R4j1CExoqNiHOP1Z/SeJSUjrwEjZ
fAhB4vjcgIzpP2s5BGjg5+f9oREF9hScS21VIWU7y1EgpBOjX1IKeOCKghKuFvWg
NmSs2i7LshBE8Dbgn0uNAVN2Ga397b1ht6+eOuibUlX8PGnYkMpyMlQYOXo+wWoB
L4DhEXaEii8JSkdO26oaJUCNgu7lb65RdUo2p+slaWj+gx5qn/0LIlroPDmjcn89
U/JtKHhw6GlDXyfvgduL9ZzVXiTNGVh/RL4i7/JhrxsDfxAwxYd0f3eRseXOxyXn
XDJERD5hEKaM9OGD/KiXpAhrmtl5TjzLo57oL13z4rKRgz2M+mwS18J6GdCW+LR5
+esro1aH8gpmhnLIZc3sS32b8YgRv/BVzhKokKkPQMm+9RBAaXIAZva1Wkyhmqvc
Hte6rl2WOx6CtO1eeVy5VS07QFUPvtPTlllmz+qFLGJ1UjuYEny87yJKK/tRr5MY
qE04AQCdyNwFmSr99RzXLUzjNfNxFTDssuBFUxYz2Bhzd/HDUvtgwxROLWwn5jw0
xJ8nkk7pNdjZ4AYdD2mHL/YtonMQyQpZ6NFQx9bFH7mMkgJUYkZGJrdUZRDbWoCG
Dw0rFVdEEu3h6bg/T2sOoYpOhXYLcBapUV6hh1i2wSN1h4r9Py4W3Ae5wF8yyXe/
mLxVrJvZcVt83FF2OAglqLw0ARz5oQo76vu0SRXe+HcLJDLwX39C7UUVIbEzE70z
dfH3v/bw+Q3/xdFNR2sKT9dfBEXgfibsOzEw2QfkkG7Lmzg2BaoToJXfUR1AH3Sa
kPNi8qYVd+DD2t2wceWIpxIf1iyO8VM45FInWLuvZxBm2xfxu5/9vPT2yqQ+j+eN
DF3BkpWELilZgMYOcDnMiNbc1B+zI3e4Oe7jaoAoHD61JWL6OEwuSyk0UaFuvM9N
zZ+K3EVbAJ3dQV2xPejkUsFzrUBi+dC1yYej9ZWvb9SmYdw2me0GPxc09B3Y8ejB
Q1j2khZipQCJKp80vY594co/IsJG3NBSvlgRRVCOAopv5zcKLe49cbrjYwWPAY8q
p7TBf2uxC8uN9UpdQybN3Jh5s4stglHOWen6nauZqrsUsus355/UMVuntHO3Qnm+
XR84dTBO4QtIUvl5WYQ1dRPYZDUjVJj6CYzZeDZsxqu8vprMd3xJikYXH9RE9I6a
XHTXz62jqecJBN1gbVufjUUhy1jGhfIzl9B66IMFxudRr9nRrYRvsyrCexg6gjBF
U5Pa97b/VNXUL5qjFweTo0f16BZNFZn2C5HmSJiRC8od8GJkYldDG2J8FHLmOa12
Sp2b0YE2EeHeL7BRIFcUQGH6CXPVpWj435olnW24DlV5XahqfVL2DSboIiZNCNY7
dsIKTe5yyfpJZ94K91tp2oI++RQEXwM6VxuMdC4/9jUf3+3oLROpLi+P63o7NAPf
Ixx4ggb6KOdWozPjreoaoj4OqH21N0D3Ooe7BL2BbBRBbxrUr3e1VagCwtnYMzva
3PaAGV8ZoVrz6IpGWtnHpBJCqSMssUB4NwiopbaqCzxTIUvMahM3zYmgKWQi+6Tf
n0tOJURZfRSCYE2Ddj9DKUKHzbFrGFsDrp9tAEbGTvvYP4/cuneEVgR+qHFxNhq6
nvVwTh0+CRuzTaQDZLGZuTF428EQe/79n7ed2mdD8p411KWcasCmWruWtZDA1SXz
EkMJiHBnztXWauQSOTyaNdIbTogvTrKRSLzg6pOnxBL/hvoVa25vEcgCGVohCWdX
t0t2x4QTECiZ0hCvV7rnoQsvmRhsqBd05tbDXSetEn37cFo/eYC29dtoiaaGbmxn
GwBlrw9baPNwcubwGYzmsmSEChoh9LNRvRAne/jeZ0ymhg6p/nEcplsEQfJgRIBd
fyKM/V+JgsTG5D13Uk9VwFAMj2oy+UKL7J0CkXlCSHJOaBZxtETAVrlpBjp1D6xI
7XOAGolWxXa9Y7qdFgGaBlIDjIDuCiqh5WoxWvIAbwiAtM63rxwMpvmye5fmTUUJ
6VCKnoyxRqRlV0BaQGx4qmfs1NTUatmd2SFwqgJL/kmGRjbLvwcbySzPlzWyJDsC
gZaD1vrGReqnh4AB1THud/V4g+B8c4QdxPMiV0otPKlebsqoZuGPzNEcyfbC1cwj
DwipLk6To0MguZJzMTmRi5aptxYih83F1KtQR8pN0tl5IA6Qw1jNEL1+BeRFpnzz
3hGGsETSkikM7ZkaXXwzQ2Y4whWTbINaKvRs18WvNv7TQ5fF74s+9SmC8p1GJJFf
75EaVFfaVGAnrTJ3yu0qfVAax67JwZ1u9rX1zBLIR9D/fRvxldfSk0FRari7xPZP
2G1BSGhX1CooWgkB8L/9wEsosLyzolZus2OcUiIralO5D6cREXOzL97YGWQERSHD
JGjIvTFzR64T7OMiJTaAWF40rbWrQanBw8Uj+ZzSKiYVa/kFGXIAXpscu2hxmmv0
gRHEOIqOr3UMBgIPSVE8Nku55ILPfyUTc3zJ4AUzP8UJMX++19XP9y9TXRNYneOZ
x0AjJ7ObO/v5dFfdGU9NEVVjEaaDXiNF5jisX+E2r47dc4deQPabfnM+Y9mT69OO
APLx8qW1ZOel8j0x41b5RF8G6cWbUGk/c6+tGtvvRfxEphcB2kH7WeWg+yjzJPKP
KOH91VMrOTNKaB3712LsnAsZmRtCkAMqoY4zMEOFyXG6+vHRkEv69UIXERzhpZDT
PzlEsZUZxbIfDLdw+QRxxliawjRcktZ8+UGmcXPBdlHgOsgKK4F1zAzTEldO4MNa
rWmtGUSB9t5k/eyhhmI3PJQSQlkOM2p0Y/E7p896H6DhuhP8Bj1+M+T5yz9iB+ZS
q7RNFv4K+yV/U+dhq+Kx6wzAiiE6XQB6qRp/lMUPBVGKVn0gLPeY8UKwU2IIVYjs
kEcwPcft94i9RUauYwGRkEWDljeTRrEjQvubuutjO4fGwqfNWqX0Q0GFLY1t/LY/
ib72893bxtiBFhnQTfkaOJNkjYAO+Cc7A4fpDxr+zIzIUCyYttxfsMP6E6ND3Ofj
pwnlOHlSpnC8uq9maaYLduAIuUwJKI9PGMV3mb3+IwAPbJL+9NvMBJbnUaP0RjCR
GfHwJ+ykcKx1z/Ta5RjxJjeLzrV6tQ4gU6Y7IucJFfiafxWT5mFaqvPVseT7nBl0
3eUnZGDapRZuJK+CahmjpURHIIpmDfl/rfUsVBIKzo0q89+R/7G5shNj9gMXgRID
pwknJZJmxzISQEvTgs5RTCOP3d8DQwd4E/ZrSddCiuy2LXTgcSOxiET6GsOgAyaa
kmp+U8CLnU0dsgVaYaNS5rrzBu3sESB4vSkipJytWDRDyD7h/pNP0OCEndUs+rDJ
Vh5FAm7qE6zzAGgOukD+dYiU/OKc5ganf/Ir2JM99vtfeT+XTqB8TcS6rMWljZN0
XkK7OdqPpPgvRJC2jTOTCN3VVfSIOovodhwhz/gpnzvp9sWDfRp9xR+3UFBy82NB
kK9dy18/axCQTw5e38+06SKh6M+GPDeaiV7Sv6EYsGIFwGPaYh4NmIkRwP/IXq5F
tyVgsCUiJ2MAgJiTJGcsGlKMAaeJS9fNxoEisQxqmmvhuhNgukjpIybfs+BfGm1G
JJU/uQMCKO4lFfpmz/IEz7YhiDOAO+Ca1rBLtzNx0mN/iKAWyP3IckOz6gbJJVwe
iL1rlfrNL0LOrhWO5+NxvmspkAuFkv40O2Rm+IgsSyV7ZqqIMQFj/YsueFxyA0fO
2ka/JpGFjCs9AowUwqvGR1xBhTBdFTd0NQgCwvpN7gCuIAvvwZ9hYoBl1+RKVUGS
Fi5X46/m8UI+sWlfyEkHWayVlvQMiehxoH2iKzjQ0KTCjQipq1JI3SbsNRRz4izq
WYkblDe9rjApWg8LXAwrf4KeaKgVybEFP1LJwDsPcxdw9UJFkwgUC5Pvg9GvPOeo
W+H6Gt18clzrHLkhgQB77U9l5HTSfkCTD0VBj0gpPYiVUR4rd1q+xtklgdP+yF4l
CJVki23OWjKCZWLfL3gCFQbvFdeVs1Y4uBEX9hsdD9wgwjEHwbxxwmRUYt6de4Gn
tQ8s/eeBa1OXYfjhO4/9nlPuG85Wwj8dCfRaHRiIja1ZVSuLyjVVoiZnquosVKuM
ii+PQI7POWIbIjYHVqUsE4esEKk5I1hmbVKkoxkMJ4yzJ7e8Vq6A5eucjVsJZ3GB
Ap8W+pBUXq+OEV2qZbmnAXU6ZNe6Sw+65nXHn3Ss8SPWKVt3nfuS904MUa1iMbv2
Ll1Nf8oFt5zf6YzzGx1a300U9LIZtuFT9GAlQa2tkv5uxvR4FAh3C+Jb+QwakrPA
nL0Q39G/XhorMkhFlFxVqnyddYnUrbCPfRw0zmkaIQgG1itrIu+iCnWq5IKWvWK3
w7I4AeP6j/vZD+9DCwv/kqoPCvC+p/p+cUYt1oDl+qH8g0DDbXt+IN9Bff7ILEJ7
Yqd+oM+z+ndP8+K2LG6sLewFmUjCi5RyTPHYpl4663ruYh5hAAzy/Lcfyr0pkY4x
XVIsbJgRzhyKrYeeABoPtOw1GPbITCIlEXiZPdht3SRltYz+/vP6O51dDyswwu/F
2aLzaY5KJsJVtGN/vzlg68VawfOvSoMt5o3qDdaLpCay5xqY90sZ2wzsbbN8D35f
QnDo/iz5jTIn02dI2ODn7QUnelEJj3RZzNkhtSA6iiKvsoyoc60o9a07f2Hc9pQ3
wjW8D3J89tFp1z7uAHs6BYELBI+vu4qVXaq0WcXDlq09m6EzMrg+sFk02sbzLmQU
L9kgmNqQfdgD67o8laPRtdc6tg+oPDtY2kNR9yobPX75Bfkxlr1HdWgyjsW2yIIm
R8VuaAVEttXq+im8vqDSxRsj94g4M5qy2FoPHeMrJ6J9riyo1t6eYipYjDm2rwhU
CqCMrFMFeKczsJzofMeHmPhRxEmWffsu7Wdlb2KyBc0wlMg+D30PP5COyi20sthX
WPvrXyIthNmQkiDs0AhDPxlHVm/00wEp1Cn+DF1iQAGpAj8Aw4En2yHuX3AGfeLj
gC29/tjhhQIeRQnvpQaOZI22eX1InUDMn9Aw6b6vfQC4n2uhoh+lS98AW5JxfeW6
3pPOn4eYSGi53vZ+Algw9mcW4B4J1usoqkd7TMGJPm8slk1msYxVImjAyJvuZvmN
Y1twX7YpREerwXw77irFWW5f6fwqY6zZwguXTPrfGC7oE51lIo4JY/mH0F2nQ77q
C/sSJXc2bq5mrbBrc+mL9LR3xOFikkKlnucYEi6deKoA7XQ7uj89h2rFboeHIVOq
J/EgrWNJOuPDicfm+E2vL3/CbTd9WCuUQlV/S7NkpksiqO8OyxMw/msNGJsgammL
UJE/ig4kV37PRIVbHOoxAHmg1yMJKUjM6j0R035nthV0oTLOPWOzLY8wJi+prNmQ
+oAqV7qhg5PUVzK0U1i4VtoY2ZCWyjw97U8WywRX3+5v5Vvl9v8611SpDLSaSWex
wEe8YdMaSPRNDv8LugMQ59Y9X+l61Jm9fYSVRuGVfHJewcTF/xeV1H37uX/b8o7B
upolNgwhYpTj4FzVz7PaPObtXs7u4lIeXaLYmdC1gVjcKHh3X300qE3HSgFj8IvL
EECdvNfIuwudbRr18vAxKAXB2xO+UllRFAE9y59TXQ5HuepzpovrIPe6fZ1mkntR
TbkeERv6/SW5AkeozDsWmsgKdnzBUWVGKaMEQAlMLGgw+v419SjZloNfiEYcAuyq
5qajvFy3DUMuTSjyGLFCtL3Xz3KaDYBaMr5QVypDhuToVNMmz9rf/R+LCPPWcH0q
AfXns+JTlh4Aia46G6Q/N2Ac1WRXTnO1k0PSx6jCADY467+rlMJyiCDE5obYFbkm
BSO0Ylh5eoIH4W8JbsXo8593Ni7J+IcoEsSa9hwr6dUbfgO6R2wDmzYbqsuuDxxN
E0EZdVro25b1yMkbWBFN8rLIceG9whdcG9t/8HJTbtZ7FIlNqe1eSP/ylMLlYVRq
jVjCIeDgN8+YfFov0SyujeltLmuHmG5B2QxWllf2SaKjDT2DOndLViDn74H+d/7k
4Yq0ibNP7v7sEFbv6N1m1qw+5BsrSs5hxtmpqX5wtLQTlXcx8DPa6CnjHk7yb3Ny
D4t5yb7kAgu3MeqXcfmpY8drnMCsBiVlActFkDo5nKYcxSaFWmSoeHpTKA6ZIvPy
hJPsJ3kKuYSkiZKhhbcVrPk18wDQn8uWZYSUksTrmjFyO0cxo5Sn7yDjXhASDhji
w8SFzUCfe91Bpzj5UEc5FWZNOrws9u/ZCPxIJ0Nb0A35hM4hFehDOWfNV/L3UtJ3
mNimScMDX7OiSsC/eb7St273mkIJwIlqaWZt57rVCDCwRlerNklA6HpMhEzwUK5n
8FCBOjk0b4t4UUk5bm2LPCFfJ9NbNQm9jKSD22G3I0o3N3XH4ZtJieJmVh7ZjN3v
Xiq2TUU35WTXiseYOqCV4CERbpwbFz4CZm+sb759k0mioiECpj1PMGyG6jVAQNSf
zJ9sDuxnWyBbjJFbtzCKTTd/YBwtxQYeW64IlxU5zWp6Th3LjoDXLu0JkUW1K2Ax
/eoL2fcoV6Yjgv+EoWR/i3rSYhnEtujW+9gZIMyz0XWAtjrV/MUBZ4xLnj64vaeI
97WiDrSBabSDBTOqKMwd6GJmW9qp4rcTwlUS0jcRbMrt2lMiinwp51YhPmS/4G0L
3rqLb+AUo1OEewiptUztrKlBuhm7lIeRxuAbghazFzjEKHz9nSqLQWg3AsahVPAQ
o3MQs6YMIBfAKm+xTtA1qY+krWRH7VSeiExZ++jVYwVhVQlYiQgG+IuufUmQjGNS
7b4zVYeb4QTaduKi0xej9PoZqySRTo7I6j4ADOJsP6z7vtKWLpqsVV+ZCfS2F/F3
95bTTR1NLPr8O9DLgkn2Rzq31NRipNI9L3l5BNbto3UnYMzl0oOhklBo93qZibMj
2YmFF3VomvPb+5BA03+vzCko70ixuXsdj9ZJ1r3KHyFNlasNglS7sDWr90tn2UxG
AfY/oWwxce29jz9OybYx5Z+5jOJvX7N1q9cAEcHjy/4SPq+7198IE3Te4CVjZhNo
Fz2oNq52bFR4x08pMrYnsbq0VR2+JOgvvlTq1ZlCz/EPcAlqC7kdqJxWdM2+Ti6M
jO8dbob25OnLhgsbW8HhQ2bqNDinOIh/Sio9AcqPWVB4fPQhnjt8K8TmvnOd8L/D
xtJDv0KJoMsZ/JS6vvYwNpIARCWJFHfnYqEIU4By+HWcs+OANbjZQYuzMLPD80Ne
kkR5AKIlE5g3k9JwWQgcQPhdV8oGQ4lWypXg5ZHJYBsYmpbZZNhN62Q86xPR9lsT
2ubsoFH+QZHtfn6KMsxGxbpD17rjjGgzmDHxXcLEe/YvV4TAymfg831GHwayRq3D
3aHl+Uj2ZNIkEYlwR241wjEdm0b8F6n8NlGk3VLJwRM2aD9fLhZtXQmzGPTW9zXc
EyplwSQMfeKTnC+6r+/EzzVzbKEwSlPBs86svAbJxqsNavw8MQYr6fdirQHuBMxr
qEXpd3wxhXoeiJJw2CQinoiOqP7bKiW9yrkIjhjLK8lAGjmhLuv/Bbiz02cmbNNb
NwVVCeYX0p194Y92NvTWEgCUmsIEdAOIYyO0Dpdvo1Kj4Rqx2gYuJXTgx5zRMPDZ
8e8bWj4svxegVAInWj0fIjfRjgaQZBiS0JtS3ItcPNuV6/ZNfdXdKmo3YiMwsqoU
kSd6kzD2zGylyCN+7SntJ5zfb4fhAOT/E1ZRpmcaxdeSoIqZZn2bmGiqEb3HL3KD
r+GQjK4DieV+uTzpoKBsiBir2owAMF4fBnhiVzfSk5QGGv4VY1d2MaY5g7d5impZ
VW/TB1iOBBC9IXoSbzQzZ8jvPh33Ay5VZ3QdwJ5yqq0bDadThdyZvRD8DG9B/qRV
idsfkQTRMCHuZPSiOv/i6mmAZhUlCumK4yqLp2iqSBpKodDH+TJ4MW+fHc4RxdKG
3yqMT9S+/7kIFIuBd2ugmvtIiMRk6BlA8bhbPpKCo/Q4OJwKQSUNmSJA+IZybmJI
Ix0bZGx1owOQJB2+O5+EJAipCb6mN7+NLKHkbnmx/7/qIFS4j6oAQZLi2XSwBJkL
MZKbLQIxV6Gcx6Za4OL4HXwqBztbQIYQSZK86qE+dZS/eIHTUHwgZ9TgaVYXultm
YubGh2zaA5qlBuB+G9fFqDamEagNv11Y5phL5Q0/09kcGN2Uc0iQZC0TETQwBNW2
0Dv6QqxYEgR46K+dIH9YLxdukD1fXMSV4j0Mz5zFoDzzRCvwRDO6I1s7DFZl271K
YuWj9DONKrHRWcTbSUL7BFUAauOap/GHMreAlzKeybpklb2Ow6kgjAqCRgPYLwWr
WmeO7Ch7XQvH9lgzFI5DPF6M6hvIvqx2rULWlJ1QNWWoitWgacKcBrMgfrS7Qlt+
ZMnAarypT6F9zfpQAKAP6ismajgPnBpLYcV2ZtbO87p45YNF5XR5NBH+ZBJ0S4nW
dFjCXGNoVgVKFV4W4+6mxjJc12c5qZaLGho9T2WpZ3Hk5wnZQ7Snr3zaH4utOZVj
NefbLEON9opVaMrqMdI17fFFMHynjgVMZslo2OpfcI0CW1e2F6dLauFnNQX83KwE
+sX7MDoN9N2Dw5WidNKVkm4Kgqg1lGNhAyO3RcOD+/7aoRndGLPVkBjSjCiyCXCu
wiBAXGWes0DFA/520RKX1RJRas+/RtICqOhk1avhXcUTEJR748nJ1I+J1gS/6dH+
aGZUvVX+vqIqZlxInI8RHNapLRsMu2Gegy3MTfd1ARPm+lX2+8+WAY0OVa+7UowN
bAoeQ3qtKEekDPgAl75tFwQ0+M45pTumzAlZV3xF05+3teSekmh6a5D9eqichcKO
xHH8e8tvKyWoDC1FjJhPF6/rJXsGLQrwa6thCk2StlxQmxREM6cW+xOWJYF9AOLt
ZmLfCszsnGkAzDc3KQieRBt4I2HJ+UgnEtqt+FDt31zrgsXDK2AVyFtnJrCpil+b
JN2eQfeE7BUMMoL3uSgAjCRqVRB29fuqk9cN12A1OUS0ila0x9t5jE8PbaXkCgAL
IBl+SVGzZs26Pfm9cGSFvCmoOhCO5rXES8+Lnt2PZ7byqp56wINNRHU/n86rK/LK
eYVI/ubU9LeJJu6HieOjKqPXfmNH6lPUdbbtJBAwz42nCXiTXbqm8APmyLvd2i1t
U90ilvkPdYbuLAAJam4EvTjjaeefZwHI9PuHrMW6nZDpV2LYMWQvrFgN+cyJuMwJ
BBgVcYJbKpoPbp1krzgSeziHjrdoV93Aoqk/3SAUK0kYcZxlOmBzIwssHuDZmLKQ
CT+JIXOpT/kqHo5m3zSeUd7fvxZsPIZsakEeiQkMuSyWee0fxf6OR8fUacFdyH5x
wGacP1ZqC/+Czd0E6NSGD5qqODs9CRTGaF0pbXFvqFSJDu0w/qvDIDnbSdFfk9pj
TaqWIEP7licUz2yPflQ0gjKF2FQ1GsPMmArNQYo+s828W6dL7jZDguLkgBqWVRwe
W8Gbe0UFkHYbb80B8oOHz/iYrn6Z/PzA3JPFGVHtZlv30906eQZ0ryUk6rSdsXej
MoALCPPLAwtuodcm8s+IlbaJwgb24iaJilcmveOTQEIX7Q9ji7ITcWKAeWyhqZNJ
X2rx066TwQXfDXgHnxgvPBztGYg/tz2BWi3GNXCnQ4XgoNvvTVlGjcv+FfQfp1SO
GCoXtpWg4U5MLgFQ0oOQFUMAU/QlCjGDg4aFk3VH4+klGsN6+JYJTAyNUe0NSjHq
/2dnLhqc2qgPFArvm5l7z8kTakOyeiBXjqy/Qyzm+dAf2bad4J6oT+D38ZNyEbbL
zfwVY1nU4npOPKqGlvPP3WdRt0EkoiKr9FewAKxpbW2NIozC2FcPqAWKM204QA7r
G+Tfor41ckdna08a6RaqTBcY4zuV8WoSYgR+Ue5BT8S3ojJ3rM3cs9j4njdBmFpG
G88Xqkjq9Q/2CYk1rXo2my6jm71XcjyYukBGwKG9Y2QaD+m9teOZxK0w/StB2AFG
hdJT6A37urVLP8LSpQe2jwDkg0GIjQSc9FF5BAt+QWhSVlzcmbk7958Df6JKGpb8
tE7m3koi0Yg0+yBftHqLmzTtWB/B5YibFyRWeEs4BhbGvjZSj948SQEzzqh/IeS6
dw7nB9bQPv/xl0u5Ow62YsAZCAPq/rpbz9KCqhTZ8k1Cv5PM9JA3nHKtav4YrNVx
crBakzv+igiG1g5BqTCJGGqRM4WTcmJblTvWwqawtI4rT4rFkOdAxmTHCP1m1UvN
xFLG4vIL4VdxFtFEMQMRHz+Ugh+I9JbkTeG8Raf4CulkcDpkX0clCzzGdtOV2go+
puPGYmMF9VGZBKR71h6Vh/b3JD3sCaLrdQzlv8lL4kUDNfkEgM70/usRlE1HQ1a2
OElBqTYonnz5gi07f5m7Q7HLRStu5spF/ZDPlsdqWIy8FRjfAyZ4L0No0TcnBgEv
WGm0rQKu8Gs4LUHyo2JJGhFSdJQ+tb7F97cmG+A1fRdpGS//EZlqdOaMJgYofUZA
8hUEAkEFcHyXhSFsqepz/GoRb53MofyImbJVE0dbfZ+K6zTuhP8DyFR/XLbVLzQK
mzoZNvMoXAc0sm7BqfOBfXLmK8+MzrAJI6Vx7x82XOu6G4eD972DOniYIDrNaB86
3d79f+yA3GDu266KRdolXvGhwtlDJFzo7DHw2T74BGI0w3DPtBdg+RnyjL231V78
88AtSfbM/aEsQI1fBq+k1ENtaOwy3gcbdTEmOd8aUbaj7Evri9fe9Tfz33wPEWn3
BTgNdkecVesyJ4IQJac/5Cezu1nAvVcMtweAJWrLNIPD7VOJ4I6YRyyjybUpieiB
HXjYVjslDDvktLLa/ebN39bMS+ZQy8EJ5noT8wCp307bKc/YreO7giGMLkrx8UYy
+DCUdXfvdJuyUpe5ZgEOPfAdej8RJOiba0thVov8IK/YdcrPueqjgsjD3OVbe75f
bhCxxPOt3m4B8y0Y1+3kFwhf3kKEumRN1FbRDEgHdy9pl1nCOzeLwMH952ZuFpoi
N4p3LBl00FM/jvLeRzpdlHDGZroJRLIvgUXLdfhJwd3xElRovLvxP2Jhh/pqc/rz
dFUaVtz+oUQHtJiSx/55AeI6JlUqmPwLmOsXDp21ImCB/FloUxNlS+ME/IhpZP2s
rEDiFn830NpgCgO2qkVFHQsgS4CsijRVmHkt9YdryqpJrwx4OWn+An1eVOLb28Km
SmSJIqh+QjJU39IMkYhTxcVs7B1jBZYiI9/isVpWNdNYU88co6hKQTo2SLL1OUZH
04JhPFKF5hWJI8MpZsHl8bDOuTE/oeHyXOQWQR4r0x72+clqGx2N+yJO+D0Z+nCr
dQkwbpfNqE8TY8Bjhuv/5bdk9TGA1mVI1X/PNN20i6RHsMGGVZ1vFz53qy/yB6Kn
2mCfIrnY1hW4AYZBxyeKWWlvObiZX2FsndRsXIpQlzufrvVnEJlSnllyWZp7DGZH
XZwhOi4XF9wVMSBdcJJKwXhUtJwd17i9UhEtNNRE0tpRKjcEl/AyTiTDztOBglFy
eXeGppv/lasetzf3DQyKUh85p+gbSbLvdoLz+PL9OnvUcs2usBWoghMP1e/J1TpQ
PyIHiQZX0PB/CJh1iVVUWlIKV0KNIKtCbnaifKz+d4S6um6umwTWxDDFNedWPRWS
g1hMjJU7aNZwSviEgZbrlEwB7gr5CkCeb6vROKV2GGaOAIqsTuS8Kw8MkTbXt5iD
P/2trwzGoWQdjvbL6zLWn4vVoJaCw+DQPeMRMb7aDX52lVqPyD0xpYMQXQ+4K9tK
/bDmLGyx43xJXVV11ror9tRkMMW9LDN9/ss9v0E/v/NW5UWcf2LMSGcK2Q4R4zoQ
WIcAtizn1Gzs8h+y5WhIuciiSlkx85OrC92n5IxmPgVe4/FGILL6SGHGzqoqep5p
jqVSHRFmW/Eb9zA6VeHFjK+f+oyYWZC5yzQWJ1kHuefUSu0lpsBphLp8ulGA3xCy
fepnpxNGZb3q6OkheF9yCINeu4EtHxv9GZL4YjDEjpa9m/y3X1hoWxTuAW+Ev13k
ablZDqbaqYSKR5MD+AuL4a0ca4PIbjy27pNc7ZsXGGd6tw8ccdWLhlqvtNcT7FEG
9K9ZutdDReelNRYjl2ij1Lksq901ingIxTbjFx9/QJHmy0BwRpxFE3zlZlD3cjg1
lqXj8G5Q/EYh5wDY00wgXXK8RP/EJ/2sBZSmhkBhNwpfjHdiFIt2SAnobMRhp6wa
6IqRgdFjuZicCWaEvdoa3d3a8p/NJw/Vscx8BVgM0CXc0s5jYsJe9HB84jMfPjT9
EYqZ5Pp8eExiScpcup2lk9Dfp35NPgH2N1vbRltd+vHIB25CgRLIPVKTXJNzmI2I
iHmTei6yForW2v8Rz/QUkd1HxwFRzQcSZbTZ/jfR3XmGfOITcmO8XPLi1eZR1sa2
/Kr5hGtYysOsbGRKoWGpYS8B0tN1hNzoUvynEhPAmSSTNDsDBKfoMRbrx0QnGTGX
AtwrN1JJOTKyFa5IAIowQ90pGInzxMzgDZY8UMOuWzBxJrLPn8W4/gmb7zXxtbIy
G2U7e9dTvhuV73xqsJ+CQ+tkygHkrvjuV999GCyUqKQMdeOMyZVVFwQoqdkO00Oo
MNj8dkBETmI4tqH2tBdIMv2K5aRXl5IkTlraxDlnE/A4YcNHktNJxZ//WduGLw0R
exv6cPzRBRlSj1W4ZVHuVfJrrEMB6ZmA9z0GJCNOp3xy8R8wi3YFkU/4MA1llf+d
JIjR2S/Qed2foCKFyE1rAE/lau4ULF+RdGEblHrfpo0L9wkjW5eUlEVe5aSZMaHR
RAB4ihRm4Ffce3uGoE49sTl2GxKe1f81fAlfj2oKRrMrBsaKW6lj/A8prirkNx04
c+pyEY3OaKCSH65iIH2U/Yme0xvY54HUn2rf1/osFOPbsSG3l7rJg9Nxdz9WF+zx
9Au2LA0foPgdX6qq4eJ0KYmyc5bN8Q8lrKbJso1srwzR6IyHAlZibqpgfyJ1uWoU
Ghnjj0ZICC/N4kMQN7m80Gc0mgI4MV4bZi6YLDnD8L4ncGKfUR4/BOMd1AY73MQi
sASIuwzxkHsQbV17AtCeprBk/YF9L5GYmsCWy4GtAxesRp4o1yAOu/2cY8PSXFNP
+V5Oj96GAHH3ntDid9On6xZ9D6X7NKR4uZOG+A/JLFHGK5s71u1CYz61mYp9eGYA
god1xbMHgJkDGcPjmjab90kOPX39+cylIS9J4K4qA0LsSrBsqPWDIrcBbvrT93aa
jpxpRD96vBqA/hr0YfSDjv+DFIULZrfZ9LAx2j1oAgSFHALiMOjHU9qxT/pI7RDF
+1KYcybXs1maWSeKwmY9TzSCbhbR4/fkJqHT/4HFsllPwX9maGHt2w9Jj2Zxk5QI
waBJ3HM5VaGHZ3J0xtMa6nArge0Yum8rMpsW1m3pPTP5hjzybjqDg7rzDLf5AVzb
35IPTIiKK9TyfXKQhF9KKyxQTXRU4U6jfpoeiNX1hdR/zB7YuqLC6SMCkX9DFJsm
EnTiFAwYa+XStc+lFpmncQpXCplqF1wvtWD64yByyTbwxdpX9lwnypYL7bTdAnBN
lPGTYfxKNcEtaPpq8uGsuOQovSHxwHGsuL6fyd6hSgUli6yQvUMkOD02LggynNiM
OskB72Xqw0WPyKwm1EtYPB+zQnzvcfj7WBkRIu+M/Md1Gu41fE+krQUjUoVIaiKH
0UA/8PfU3cdvwkLX+VUpKnHWkiOPaU3CV5wQMTB7o57O4Fs26vnjrosWMmd3i7In
H1awxsu/H5/Vq5T+WfcyzSLpsVsAjEzKCRRXpnZm6Xhn2e9mxNvbM4FpUjdciKit
dV5nLDbZcK/lB+9rbZLAnFVEpWEQzYtwp6HNQLL3sqfvJmntvElPXZzErnQjri8j
ovdRxlKuJDI6rvJEOL8nQXPV9PgiXuEXqqdirZwv6JEr9F8AsbEkfr4GmmZhIUZh
7AeXp3StaQRQKD9vYswUKjNAUp9D50WIj+dlkFriwHShIydfh8TK+K3K2MqqTH4T
mXDIyWIg8+X4hKLb+4eDieZv/O8V+hnwuSpPPWfVvus2sIQXGmo9ZqkElVzYpFPK
6HdkFglkCqMkyFc2OCRDf2mtM9sQ0Hlkq3ns7S5GeVsG5eD+QXN0roj1x35gN2/q
MqazEoOzfG+Vk3BkHIIPT8mWg9wb8iyLm6Hzmvy4wd1u6UaSJKz/5MLccRmJigNB
sKQGBS3T/JGDvDCF/kBV6hQyvL+9cRd197cugj2Tux0DYgF01XWglmLPHEwZlli4
z4rJ2tIqJNRQuyiADQh8WeNZiH1nKIyPxqi9ZOFEgaRNt+Rb2NvTyQB6BsIRsPLV
7hFj/z20M+ezeDCN4KcVgKjaF91zK2X1UW92Sh98eChPNEW9EhgzHLOW7Hq8ZDSU
Azx4zY8dlvTPzKTdDsSVRoZCVHRgzGEG3nyNq5Ts71Qux53kgXOIx1eyJjFgNFxt
ezW/DW6h428XV0H5OODm7RuFe3T1KpVshDAHP0wIfAB5qjmAj26Tlk2MS1FCJqSC
6nW+YvfrfLto+CCH2ssVG+oV0QTjtBWB2J+LeqxHWXoRZ5J/V+3EocDZFHORV5cb
+5SdKyJeNKXkkP8WWixd9gSZBD3VHGVEh7QvWLcTrv/fy+cbyVG1kql4MLjRIPIN
WefoX+WA/gcH2VD6oJjfZarP8+wgEybBhZNRIx9hLDLOiyWS0q4nk6+H8IvOrSiq
mP+AeMNWmCdNVGmuQ47bCj8G7oqSp+rC4UW+5wPls+rX2mG8MkYNNGKFi25VuZF0
HOIMQEMZNlaRZcWuk0cwd3FTAW7k/xzB6JkgEsU0l0OLi+Zg3Q6p01Yre/SKUiPh
d767QMsENAg9/R76J4pPYuqlryYKgNockKskTSTfNsHZmgGQOVOoGEf+NOieXocZ
T0BijQSkfmISGLLZuMkPjgD9xemYzJgvyI16rzJP0+xPzWPJC8hVEOplh3uGNEKV
jeI3FE50RM5XrDKfHVH7VxCHzU83fYkMg+xkEEs9apSgrecQdED2t6skCXJnVzba
Zf5S6Q0fdWv2bIe+oMHd7dp3EsRcwFHc2X4cqLJrS72MwZvldzuop9syj65oeWt2
lj6kGLX8odZv2szm74FOMkciW7ocq9KBBiRRNu2Sbz8whzTHw/9x79L13HEQ7/S5
HHqam0ive2kLWWEpQs4CulgUgvFvwumVKv/LAf/RC1EOBUoU/bcvW2I9JFdTbJmi
xU4gIQTORwXSh9/Q4JpKncTH7jBCP0OGx9OH4Wo/zNiJmEn7ksHdXvluKi0N9YrT
vuB+cwCbdkfCrYNXjk5nwrHfg4K0mwckO5alxgbLVxYhC72OeDHVWiZ4m9nZCBVO
Grsz9CZlxUhGkr3ooZxA9XeG1Qe4DACz3iyutfxy2JrDi3mEboYVCqrTC8lO/rAw
l9CLmLulpRJ3lx+mCQ4E+oQz3OMvRjJnTnyAJ7YiatzNggmQVHI+npC20a6QVwDA
OsUkdfqo2OxL7AhMNswJC4IhdpPSANlQe21iLVj4KeFBWYPM2OM9gbm9AKfb1fti
F5LE/VodwfClkMy6+3PwwM1xJPHidqEI+9K1GiKHzUJbGb/8Rk5BX3AZAP6KyFvC
OAIEbNnL+Xip3ohjzP4Fode6a6oYjhRBLhZH1y1E3bRTWTYe4mlkXhU+/jYIRDA2
epNo9IWRpAvIHdmhzhVzdhmwlXxhgGolEPigp2gZJXLEArQkuffrSWTlnWjPQwoH
UKGnJWy25I/DHsT/tBWys+6MIPFXAoYqk8sJr3kfKz55c5FXjGF0YH3NAgoSuQ60
quhHuyS2KrsvfNTq9MOnmaQQaQwulxzOIA5o0ImoZICGg5Hkg1MZr7m39p1BjP/x
IEsx98YiN7LGZHnkdgzXXwSh5fEMrazZd8ZDNV2Ta5bIdoQE8lxFO9sZMvmUVAb1
Er9/Lyn8WrVk6yxirWTWNTiTsDy/NRieOTuQNWoYpHNXyXyuJLFDz6xYmCS16nNf
4or5UCZX9S2sff6t+8Y8gTC3j66LMKOEPRYFMmde+TvmlxGwqwFc3VBfmRkCOpgh
HnndCQTvg7zDXBXDgXXQoKpA1T1n0Sc2ANBnuwn1X1dgXBceXp7ipM7BxMJZn5ei
VxjmEugYEfAGbWlaSSH78L1XaB2BO0nau20K6sd8qOR/Gsnw2/zDfBxEX7/z1h6W
sn05PF6loPxFXuTKMqRCrN1J6DNP1QG1ehiWsTWQBbAw7IfmXOxN6LV0Oyv8xTvq
GAn8aqwwEiG0FLsUoWj4hFIXyl4/jlOE4lD/sPnDQOM1Uc4qEg+zIQx7DydmfB8d
Wc9JhUuACXHUPcYzdgp0RSD66fFo0cXwpb3l983Tft/mjAcINP634PabfixrDLG+
QMrKOs7j4Cirld1kyivy6oPViz4PKVsykzH0f551bDg5NtziKSYOkUfNQrBeryWs
UMeQ+XZtcBXQ1ERhDU+idmIMRTOAS4FYSjF7i/eKM4Og8kf+xRP5uUapXp/k7gjh
oVJZii8aq3O7FWuUzIJt7T03nUFsO3wr+CfH01NkCDGu4sc/H4h4L/dlGoJ6IfXk
3QP5FoBzM/rB/+sIxK3fRThr64QJaJ6jOjRTvDiM8EskR8g5bJ+Mdp2A7NpNyCtL
Xrwsntahg+zoPlZgS1CxMSuVi9/UvhUEhN6+Dj6DHQ+hH/x7exvzlF1ss6W4kkzm
zKsveyv72q/twXS/nQvBZ4h7YIaRZ+m+2y3cpd7gq7jqFDwy6sITE49Z+FgVkXQW
LQarpqgNw2y8QxxE8Ie4hhvKnd0zZuPmLTgb98suKNGNWvg0c04ZSFAYf7skGpQC
s3oO86q/fVLt1cDMddVUHYNV4K+gqBG4ZcuYqzgj/ZXQGLzrguR3bi0mXeHa/G6y
mI5Sv4z6qaPqcja6Uz0wmm0DBOORUE8gZy7Fesgju2oQhcDZrZmwFOA3K8QlrKlS
aFxyh+aaaIsSAJXqsfN/1LT8BYis2YmFHVmkv32IrI2HTXfAotg3Y71XslG9fMYh
8DLtOUJ/6usDzaawe9ByEjr5XJKJwW2RYmbeppW4njXKzcRyTQNfYXoczfwfKSB8
gHNXmv7cDtfE83eIYmn7FxRFymWyrSI2FzhNFJMXFiEVuwNCC0C3OgnXSi8pITKi
qiqhSypm4dt1astu1EnyI/VxdjGR5J+BKFF+M42fOhy1OiC3zw2M71HkHSlloYUR
u6mzM9+fhD8wciq/V9w9jvWm0UqU3oDO3PUrvvVakJP5jQStjD+XUKLYZ9E/pijj
PT8V6b0eW82wLcVedu5pK+C1V/Q1Msjm6CNKOmpSjqv6uD575xmgMpYfpCrk5F6J
zq1sA6OdgFZiJrCF8F/iOTNTFx8cGBe3Pya3Mej25A83ZsSDiZOyuVK67InbyXLj
yTnWgb8V/KDYHv8hj8w57bHrnOpU++QOop9qdHirgFOI7Ylhf4mdVjXA6S49xpqU
YIPhJWXwpAl3TzfixojBUW4KJPmh8fEMg5Kh7tlR7zM7cA1B/Mrqtlp7xv/CSXLS
mJgjG2fkvF2FBe7E6CrIclSnDUKxj+GI3EMegTbo8+dUFu7PRvH6UJ0lMZPQELW2
OywTYXzalYhmDNPVUKKN6GY/AirTIsKUECOkwe4/hYPTLG0xuXpw3eJwttmOnj2X
+/JHUtcumsiIysz65FtuzTiF0jR2PvkwRvCMC4ZnyweeB2OUl3CdvvEfDue4Si6V
17YGMMCx1OP/eq0RxIkDC4Vi8GAc9RnRzKF84p+fNoWNLK5MinKowaBqP9PWymOD
r45qeKLapt7NPrTnPb7+vm7/IY9fQxLzKQnQsTnlCzRyjsN8gD94DhJSxYDLAGSl
wEnaDqQjYBw7Qi52fDe2OzYsM3ysQr2twaKv8iCFD6N7kEQZzPpPVKT9oiiwHhXt
PYHtsNB09UnP/XbzX8PGnMOY3H4jAdIzHVyZiIvRHn9mIwdh4CZWXsF+1yuY6upv
lZ4o4V3VJw/wi8kXDUpOoS6FqUktoEe8hurYqIan2vcZOqohJ1DryppWThKabpp2
2sJtsuq2d6ydp8Lr5amaOyeadmmXbbc1USdHwUI8Z+3c6XiGzHpcEpwpjocyWbB4
cgx+4Qpl2a/NGVSEVG5EZInEE+D5xhfPslqoeY/Rc7Q4xN01cCLXUANhkclPQLrG
jCNtZnFQDsGg9A9gzv3L9RzF0b6wIkL8YRLARdbwqmogcrUcYApjQFqLmGhkKij5
z8eZYLDXgu7d7CI+/0ywRxt3Otg2i0NUFsqqqR3Wxkr16IbPvpkEJLwaK6r/grzA
824unW8H+INeMY3wF70vOpAuRRxsIC2cXa/MJzKFo2YEYp7mMl7lr/f3t/lAzT8J
v4G/+zy6agW35PI88QwlafVZdiFPFIpdi2HQZlbTbh2PxKztaYZt9VSaZcZ40Y0m
uipPrmS9P76P84ZWWUkqAajSs6Z9VKR5i3DneWEcOLx/+8B7/N1Atyd23va86Y0e
zheIvsu565D7YfrCONRX2cGiaPzxCTzKt1cTY/BzoZmN31ytS1NNwj2jiCNfoPM+
3skaBrU3Jo8PA9ORKWPhxYjtbiH8caJWSIjMBX4bALoE7H3tdpUACxunR8h2COvv
33vl2ZgY5q2M2sp4BzJsC4vuCdDhyH+4C5YKMfZjNVJRNcZCd4PXWEYhVGoQOWBT
lb9gootOpsPv5WADFEAC4NGkrlO2n/aVPBpvuF+oV0iC5nsDW1GTNo2GznfswD0I
pewxqSlLKgnT7KAqGnjPtDkKKD0S2DglguT42Xi9xXveJD9J0/5gs917x3Fx+ypC
gqR/W8Qh8AELUOiGaxh60gq1VMk/Y2FxWvyoQlFXollkI4dI+S6O2g3UIXGI7F3c
zBWBLQm2AjbcHssYKxiANh1s+cs4n/ufmtOlUqgz4xpteqczemIRh3HiOAMxZ0zX
JFU4hiGFqrx/112ltL19dsgDkGBxrOnE54bPXwvgNpcZfpSsCkx+B9E49zDzAYWv
ImfDSlLy0ukUwGKWneaGYfyKJSX/ZYfOBrF9saYKUbebGrfpfah9TjH20lWWJraW
k1bKyhD2lbXkvJ6vwsHRK0887407cX/VS+tOCEuQTOUPN4V/nq2odlrxPz63wO5R
d9EoiKrrsamxscKUSz47dp395ElMrjV0czHpZUGh7/F6ZI1l/G/dpM2gLdHrN5ve
abh2EQq0/uJQmLC2qCvkooufk9oTtSK3CigEz6ZtlmHQM78ztw3FdQRVpXyV60wn
fv2T7UHYgVIXT9mcSEL7BlCbGdlQmrneLKntrIQUQn6u7tH0nZdcCWbu7PHjm/XL
K2HDxhlsDWCMs4Fxbga09UA74VVV62QAzDfNa7vDk2Qk3bl3MdmB3trpJWa3F6nO
xc5E6RoClKXqNNLypBar5jxwwD/Gfs4iLD1v5Ky0cgkvE9mHHdMyvt2wxegqRzon
XBaUecpy8PI+RhaXrpxuHyanezR5DA8H7WtcpRxpJueEQqmhmU64zhTGRh1dnjyT
k6oefTgMHyw/M9hh8CX3wDCGkX5ZPyNf6hjV9uPKAirXMLOyV3jARXVoAWfSQyVK
1NW9P6nwI4v6TXnMuT8fjQpYWSJWKSRimGpJ3xL4/QaL+v69ldv84uK218/54cBC
HvD6M8nw6gpG0jqLiWvjDDlj25pM5usiX07v3ZABqB7euyLKH7VFXtLwm9EXhwe5
vUYqf09/QCW7p5cGlghFT1hnCRdC77agovtlU0D7wOwYp5iIUuMRVb7Id8OoiU8w
8ISzSJWwsfgkVvKAD7VEg2OJih6ttnyUu1rZe+E1Cuq4DvMRY7jdyPyOQaEdybGe
T1av+tjeNldS5empCUn2Sxuvoh5ShEd5ZGFYS6aQWsoh5RZoRGXhkX4zXQ15H59o
wt7YLa2NtZvSiX8G7Z7X+PRqCM8YgEL64vNyvElzlHtzlOJKtJK5JfCAlMbxoOpC
RmbUZCyf5OyPYvJYdWApmQcMCplQ1ArqJyGTCHhAohYYzsyw3lHTDsx4puhV+bu4
ZU17ojH6V6YHr2ZVPVPPt674G6bex6i9C7sNg2LTt2cA9f9u4TZoQqW7i05yD+7c
ijjwYfmpAWLHyt+ub4e8HNPnZpSV6E3y0faXyHbsOpuvz3DDlRxq9dtJ71H0lXKL
gcI9p9qRirpme8GQXn32djD4WbPaxNVI5ocMWZBsB39xC15jqOb3D4DCwlFv8mh2
dR4Tuqd5BoFsZmZkJlLGp9riuCPBJFBm9QTbmABfDM+yKUBmfezwRmmAHttAq82P
0RypxmAnKblyHknjlvmckKGbJ/6YxQElJoDZsZGFR6vBerTmXfmHrBRMMRSV63FW
Fui3Qz5CA+sCBr8UaH6Rd3gXRJAD/e0UuCkP/pNtFdC7ZbJlmbe8GPCAVRGnkH4O
fbdB/rYeTNX2s6em5+L8Js5eORqCsxVLJZk8U0OStaVGSdqxruAkqJR/DjU18Yaz
wlMCq44Cjw8lLKbY74fvpEVpNo1hNHv6NcP0KU41HfaX7iye/Zz62XyPvdm6djYE
nncloXQMIgFskOx13LFfuWMzij3E7IHKfrwU9hNxYE3HhceFMouHGIviDjrs4xKV
hmWmsFHk0doZ/8WGRbD/MwXuqs+OmMtIxDLwRRBByihBuHx5Y0j/jhCtWVmN+ig6
XE36b5dZ7C+JMYuSU53WAzRddrle+yoUffWlZ0DvyiNeV8PloEFGGct3M5nwu7zr
ae3IeuYjpsLgGS41qcnT8S15TmQM/EnVDwNTNvj5Em7nAzrst9yvlB7xoVW1d62o
zlvEtvaAMEyiRaE7ILbRuukOaVVSRf/Yr2v55H2Hf73foUP/5rV2cgLj3GuuQrVI
Pl0Ghf7KQnsEkRMI2n+axMO9FifB9JG9vqbAk7RvjI0Ryiq0PGpTYnmhIjfWQNPA
lWiCpwxYV8Hz0k4aYb3yn+/TO1UDjBaYROdFvYA0ZwtIC+ENO5zGeJwOuIifXD+8
KxGdtAjM4SaipsFmOVdcyQb1OAom3LCuQZmOMPjtKgFtXY+ZaiXR9O+y+nE9t0a0
3CQmQhBIH7LEN8dTqcc4e2Kjep4/6OKlmWCfibfb2U67QRNTlZvdN/1FlTpJ3Ns/
IvkX/4PGciZW2Glamm2e+0vWgmc5DiuvZXqkTjqBTM3fBdFBxvI71fE9GBrNXytA
bGwVTiun4RchIHgGXaoYRP+xAi94+8r6AV4RM7dnRJXFP5Nu9HcdehtuqyZNJOGD
hk+8OMePOAZqmZ7PXopYozcoX2ShTioq/tyy3I+n0G6PD6vkqW0ohcKL44WDX3MK
nS81jQ8vam5KtA6GM89Cp+RiSgPAeLslBfQpOaI610ncqU0bWhx3Z/vY0yOajvaJ
cVrcvWzlBf2+YrXlPFOIcpI4xeEBtgb2D2ga57XuErUuYmemJujspJP/0aVVxR2S
KL0PCkeuw9SNjLckpzy1XWJ+ok7BArfF/HNDr4WtjQduQ8ir6lHY78AYFuNh5XuW
0eOrpFuvkvqd74959gYehjppkwdGTnxb9zRh+7z1YXVBGeD+55RFpsYrYQum7pl1
nJ25iBblGTdklpjhSSrbPhDUS0FnuAQzyBxxBx6a26rcRV9daJUmyW6mvN5A3E80
eQ3Ci+i8NApXmOqAdSZVcbJsGcUB7BEFfsDFQfoADo+RCRjzqpe7zlACCQJpX9Ru
JJfVeS/gk098SRgKI3508Zv5VGwjlz7Rdm/OOyXLdUYsS7B+qNKywt2sKY8Obl/8
hPkk+jvEBfLHV6oxfxDXxm0tnb2KcH73V5qjYV41faYR+I10AaRUsUzS7j2S4qEc
imEbCbQODeRp6c3t0HyDBX8AC1rJ0SBCqfaROJ0OvaDuxRRJZKOCuYrwjRzGjS9/
lBAFWmw2dEgFnYx40Wkey7XlsRZ6jesqNdM/GSKIPn7dt4zrtAjBDhwZnsJl1WZB
mH6GI0lD9HGr3+a3yCFYcaTEOflDPkMP1dc1WuDqKAsUYAIxUF6uOjDpRjsNAV0H
2L/77z/hJCLOrIAy7jzmvmMZ6tVwM0EoU4hEI7WWTFm+/XiTb4tDWHh5gMBpogqs
fKi5kiF2WRChpZeeQfSs/0OOLTe5GnHzNKTnXInm4OgaoOEeXqM5M52hzG7L8/Le
mUTU10d50IA3iKfEePIQO54r9Fo4DfZ8xa/DgXu4+00HvzqXrsLB2jAbRjhKK5A+
DSD4BphVpzjJzTxwZyCcPU093oDoVrQwHXXLaW77SNAoxeFrHl4riU0dXX/eF0of
ownVirhzlJwBLX9tfXmiuvPOPVfjCripV2ttVGLmGHFCJA1FolEUuNPisrw1lNUH
vqubm1ulvirVhiw0zoZYs53IZ3gq2evgBwKQZsNHSZm79P9spDhgSjcaSuw2TgH6
A36PfUunAlmHim+67p+ixfNZdex5kXQ2kK0PJMzalIxLjPHqvrljONaQtWQ6m6hQ
MnvfcZi6D1oxjsXV2VhnhytpzwBR2SB3GWRZcdT7QQrpoTZpO6SnVTTqn3RqW3HL
JIwtpMl075NIbXWrRnc739VUKZyViOEMRp4KC64VwXIaQ14gs6HlnLAiNd63DgnR
t2nLQzZ3oUFdXk5vlREv6VNI6ckGsRCX9eP5igY2OED/EyAxPYUMUYDP++TWGWI4
b+HFsFoybWCwWSLw5SUAfFPRy2gBrBUfDHj19LGiwm66cjY9rQBONAtmyvQ3pyI+
xPmXt6+Ft22yfnW17T1nsmiFjhdsl83rw7yivufJTslsfzVYtZd7yJLWBD6Qypi8
fl2r8zm0UJFPevLfzreiTI84vHOIKwhcjEOp2ZgFlbtrI6M2u6XrI2Gvpc/0lvOZ
GMjX/lGHMQ5/0SLO+bQh0MykKrPoLGJdeZyJsYWySwrQEYjf2dGqqEtkoAVVefE+
AhI8YfWdFAO0BfmEePzb8vASAPsh5IxL1HujJjMazRNMoCLKeLtkyDVON3V8ZYek
8lA6w640V/iMfPJW60MBep+fv+aQvl6fb15BRCBNIHmHhNsRTAtfMkjZGUXmVwV5
SU+zqSoWoZkICJJk+1J9lkXqCVKRaaMIMcVfjnwkouiGQzaw192LmNaTzWrV8fRr
Smf28yuuU96aNYRfxdQLh1Et9zvdKkk0YWT3DBclcntolUHAUpt6uVmLFDQf2IeF
Uw/S6VmYBD+/ai4NF7awY7B1HTCqL+yvGatluMAAp9WRWiYnoqbGuxZaXpXaSPLG
FZOIsZeXBisYZ4GRIfnRVrqRZ26w706L2VwM2rkvLGZQznwrSbbaQ0FuD5/IqyjD
zHYvSVMvt1Aqxlp8+7F8poQi0y1XdrttL7dlAvwYOV18a0XVoEN9d4CtEGeOpW9g
5Jur7Jjhjvx5Ght801hqJP/9d+tJXpBhez6/ZJOGzlkMNGDa1kBK9ScNdnf7Vrv0
IGbKiowSKZYSRu2TEX9vM5rn8vGW7bQhoa3ddtforGcFusZq5BBTaNoptxcDGOGT
X20PacsxUUvuHM4lbK1FNys9KzCtrHicGn/erDb10U2kQbPuT4Fe7KHwIQgKipjQ
y1W5gpH4II7gbUmfseqW6ImeERLZBCirnKr2RqqvnYuk9hCYbOHq7AIDX9DoPztD
NHGR5o4bwXWSSV1PRo0AzOMlEAbZzY7RYmmo908ryEseWON3R4nVtOGNlmro+ETv
Db0XpmieqhiLlCy4xgswS1QzHZPUXKLWl+nRmMYiXF2mkyj2kHRMiy2R7yeAzkfP
cQvdMzwqylvehpPiC8lAscUrfArWE/q3Aq4+anZ4Gxk4cmv/RMQg2RxFV2ksz93Y
Eg6eH9l1SRwP3y4LYT+Pllzl5rFYNDMN/eiuTfgRziW52jlAg9TJmC9id1chzHa5
9H/LeakW5r+AjpYyYCXWMbaQSG430DJNazLncZiZDfGN2AyIwE7AuJvl4mIVOD6w
yyJeST99BWZyfWvry/tFMPhaCDAqoYaqJmr9S+C7/rEVYVQUCEFouPLLi6DI/97J
FQcmx3u9efDLDtWWBHg1CroewT4CSdePbMcjQd6E46IodansO24bpNXuPohHUFYW
f7BOS1RhcrRiY5XpMeqCN2Z6XfyWfSch+mpHg5PBMSMNXh8RE99E6fcmcl6g4wHg
m7xy7W3vzPFsxNlKZxxVOf+y0n6HPB4g/dIVSVoLNJy0tBn8wCOi6PoBayqzXqIW
8aSm9XgFJ6Zymn5wvoj0EsEiyiGZJ7rUx91M+cw8dXB6K/0yPf6rOxq9FSWlrpEt
0JRAvilZx9uUt3KvcRfK3wz1iWvnWbAicNxxDQoep0rtKo6TQ9ur7jhsiQrKW5A2
KjRS7sTaA/FmM8gRsJO9gxaaTMZBJ5nnz8Yir5czYm29tMGQPV+9pNTt3HYa8ICK
dnlsJB+0ns+/Rc31Ni9YgBPjPbs5W7adDps6jlUNto1qM2OCwC4G/UjNNczkyd1Q
lJw6rzcbXsHGBNt+967L3oHv3ocv8W5RpZueEORws29NmxszVVwpqJAbljHG9Qpk
0SRay2TBb7EUV2rVoBqMWrcaMXyImth55jaMNF0RORDLQiEOKOC1HcGx/yRyXZEd
wiXeeKhrAeP4qxXr8DFBPfyHT0VLQ7ztgBGnsC20gex5Q3gLapXg2aT7m9znJ8Nc
vMAr0uYgcQiVvcKgJXI+ihxKNY/V6FeGScwIwUOFpn5QeGsrwsLzjyTLTNn/ONlt
bv0HPzXOx7gsEVRcEhFRo/BnTzkewP2c6beczgmO+lwn6mUziFbvViBzJ/+MtYQa
w38U0GgL+jARIiQT6tNsaDHL+nbCkE4ekH0NQ9j93sFdBMg/JWDpICEC9FLhRZzH
YzCvU2j6jGsAlEl/ficb64mXBGHVwFCfNx+26QqlGE81r+Yo/tbB0WWY5TUa9EOH
Y0DLu0+LAz3mSmBelqa6HFHc0GgUXDYbhu0SqB/Vz0nP8KFqoFWhmg7vStQKYZYz
cENKQUx7wVTN3FMmOX2PC+wsxAsmrjxYUaHEE3lvd2Z7+kEnk/P3GmWb3BbcYAvf
ib56q7cVNNsfIWjh+EBsrQuFZ4olGgi68wQ07Cf4nI1EY3P8ZIfcXoDFevLdqGzL
4XjDs/NEegT2UbVkcwgvCWHq+WmZw2iDpPLzTCCLtG9wa4GvMDbFxycjjxnliiZ1
IB0caRoRW6cGSH4/5lmEXQIsRTlXe9fXcWLdLPE8t50TGl4mSbcFxMzqFm536UkU
bS3qeE4BYHrJwBdO7jdXcPHXAT7k24vCiSzyo2QCSHBtqqxMaCQPSRX5at8fwtpM
/VDIwYRrerOj8T/y2wQzur0e1FVYGkcUgNaya2zyJAc9qm2rk7qRTe2Ul5XwDFrh
sBPrCB8w+P2s3G/dJfYkqxww536ey5vSXuurSz6rcPG0SjnhrJ2eS7azz7hvUJmI
5tfZnPVZYcsX2a0yAXJRns20sfWXvtuvGrYnrA84nI0/gvFf76el3MzPV+GP6QGq
iP4VOh3hMp8ikLTqGkabywtPft4Nz8sKX30rzGD53NKshOntW9jQqaNoTwOiBIjz
IBD01WY0Eq03zU5flNkmZQucUGYzxELGa3+YkoGrniwiphiJPBy4MFh415DcSy+j
opBUNfSk5WJRCEG9Rtcoanf+ZpoS/TLXenfbyPePs142HyrIWq6IC06BkIEGRw7W
tzaz3GWHKuimRaC7MQn7ygEYUS12ZtgfaJyUrR76WG7WBOTaUXSnWp6n3UG/5PMt
VawQEStHgakeSsyfWwoYvlZTcsSxNW7mX71ekcuv2pLDs+Po0ENI/Yj5JsKzYN2f
XMIWdFZqhVRnZmO4M8adrSIivXFMCqbUzwLOLLWzDJRLqDYmfrImMqKiA0f0CdOW
QEiXkKkmu75YKLR/+pvAz+iqWxgCxAuYahNKR2OovRqTGb7kQIJbadAZi+worad3
r/Z2ENITAC1Lu4tgsFX2ITgLMXIAm3DHvE35TWVPA0alFYkAgVFp0gUOCl2m9QBq
oWLdyD7vFdBlR9LYfwY78oBCwedaMIVsfD2e5pbMPJWJC6VFJ1n/++FMRIX7WQAc
RLbWruKAVf6w2FZWobKgbg0HJC3sQeDXmnV9v1pCfY7bcU3EqeM+EOxMvcCWZ+hH
HnWT8UeX0j423T5MU9LB4Ao4az+ATAeuzC3AuQqDgxW1sZp5ssdzWhQpsnsOEyZe
i4/6d5UuQbPgMJM7AnM5hHpo0Hmi36n2Ml8TiH7pPSijOfycaL2lwes5OZnkstx3
dOZjcwp/twK9VURUOLrVlSON9EisUTOJ3dtX0C2RsbYFMceYdo5fweIWliArINiL
Cfe9CG95SgEwvfgg9wM45w8UOObsGcrToEaBhZlVXt6mRRQ5zx8dNo/0W53B7Soy
zRKyXlq71+7dOBSoLOH8PFpdW5LlwqgUcuj7jHhqMnlWot0LzlXabXz0WiiiRSff
Bo156FWO7ndFf6a6SixiKgQlJwOkeSE9AGssjNDiY46kRnVSihSmOdk4Ac7BAHHg
5Drk97ETpK6GAmjlUo/A7wssoHfl9pi5JUxMwn/3yR4DfFj0ULj8AKAtj5Gm++11
p0rp8Gzbz14xfCFiH5616M2/w9Ip7LIuJAeEJJ8xlrg9nIhqzeI9cF7IYXa0l7Y+
LTTba98MTV2JG/RTQApQurSs4euyKXPyZStn0EFKRuWVlcGwZCGbzdAiimZKl9j5
YJiFuidkZzSee+rdh5ADHChmXrj9JuYJvqCG9CJG03lNWQ+xUZiGxM50GhRX4vBE
c+zlzrWbgTWebbwdFfvkj1jEjYbtSdbHGgM+n9EjCwtou0/K6hD0IBzo+SLRT/9R
kF3oVB5Zh4j2NVXCMN4brrvs/wO0aJWbUAWYEtoVEtJ0GMpWTVgxW3uCKC1JTB4/
llvqjizlc8Z3iaT3RQBb1+gIIAC9gslUyLBUjKEhvHG5+R1vcOIQ4sFI/wPA6vd5
UIzP1vustaI5d3G0qmqGbj1TDZwdKPlJzU1PGJUUrLansoZq0gk2yXQ1dAm+ntZF
gdkTAyCpKsmuDkh7CZ+l1AOTldKz2sYMNHzcuHoT4wxG/mMmRdfRs8y87VWghCyy
Lx4KAtHk6j39ajlF3WXbsWvFbhCYT33Jq933dzSiFf2oyei7IS5BHUWKQUwF1Ujv
3Of/K5w9HXLWrQUXJkKOp/ADBt6OxoDW7BJ1KX8mLza4705DVxEt8o3haPnMXOnw
t+Dg0ZPwPB+ARHSdhCsSPecUZ0fofoNDR2KXtcmLYLiOm7w/BH6WSG0dpZtSoYQn
Z9CpaJAeO9cE7uhINwIdBusM66b3NscMpZ9w8sVuFwcOJuBwSA2ews0GIAfKParq
NQ4fWHpN6BwiBZw/vapVCB0wDjr+S6DhD862Jtw8POvwg2a8xQo0XteAiCltnHFu
OoMy3AstiYLe9VeU8SjNu/NIthWkyZvsAxxuotE9JsTDvSfoIW76w2RpU1gVDqi0
Y9D0Ty+rkNk+115AterQwuYZvFrFM84ONFzIFAFTHPS88hAL3qSRKbwo4A1gqEUg
uhm24KZ6slRnrzahJ85WyleQnocQawNF1/sxjFq9J9vAz4MbAUosfBeIXGW3FFhC
wjI+t7VL8e1x5TR/S64FWT0WYwlsPlFjmldIxPYqs8yvUU+wy4edc299lnY5fRep
QhKInExkE+zLweqCsFMvQEVIMBfGU2gjO6b4yTzeD/O9LH1MhGR2hbWcnSzNvEvA
o+qGNveRNvt4M8aywauwsL9FK4Qr6tTj76KgkNaRXMx0Mow5Uw6qBK61KAFPzEh8
P50Ooue5b2ANh8fqOhCGWv3bmk6pv+wJ1xWe1aKbgsPi+0/iDqO7WYmc00t24iIs
0qOPauN5XbS3y4YQG2YeBMTweZ5XEA1y2S9Rg1+HpMQvLXFfmNwC4iuz9RJpBnyN
xdABB1ol+78BgRUZF+F6/VBOMYz+Vq0j2W371GBXQX3KRErwKTvwW04pr2W5+rhr
EagQWinblvjdTgx8ZkUVuBpdBS+bT49V9w93Q0aM8zL7k6aeXsS079cXDTl0SLxd
4X7qEgnXoxeKWqo8SbMWwSR5HLFhnp1E5PtQBgAuAER/BQLgtN2ovt/w82AZ9CeK
47oXJtcORWehwFmPgCRcq3SPDjTtlTED+4qw3c8RcmAJsaIiA2x5BktxwLmiY9he
WobSWuRaNknd7Jbz59VulpEm/uJVXKsUpSxmETku30bcm9f1jSzUmKxxuowMPIuv
ApurIK/heRJmlrj+1rIHKq0kfi1fCo4ihGF7cx7RJleAlYILt+K1caMTEZ503DUm
XK9/PkHr/fb89CObCxJOnh42QWv/KHoNLmlGM5Uls1PuwmHFzIvk/vVk20Qyafx4
a+CvgMfU3VxQ8nyA9CHYWy1f80plfdbIJdeWrcDs7DadysOaeVhaAuFNU5LWUAv4
osR3/vxy62R2mDFZlYlkLJcHxE/bxCc0cxAJ/A6E8DFpFD6QB7ad6a9aw0QYdV7E
J1D/a475hpA6snt17soOItpZ7UhlWr1WuKPV3N6kGVy8YFRjMjci5yVBO3VN+H3s
eNRSJEswzYAqNsSIrWeqcrcQczdQ2L9uTunoVBd17fmVnA7Jm3w1Fuu3Agx4wjM5
4/CCkY6XuziBY+2lBDZvfQUzyrEA+qq1nJnDP33//t8UdYWo9WrPqx5Rp67TIsBk
DJ4yaR58nJ+scGFFcfiXtk5aEy6PPenLzdetBO8MGugJVDuCZGQoMbzD7zTz4CbA
yCDfEUyETi8AY/B6fPN86T1qRuZeijyKw5ME8ET+1H3R74fOWj5jAZC+P3Z4cg5p
Q/3/el3aWnGqI1dTd8xoIKfQgMiEJVFiIU36pFCaZ8HGVovwH3eYKICl+167R5rS
MnEzL3xFNX76zWadeC0Yx1K2oNWGlWMu8noDO5wMc+h6QR42CB3lHvDjrTPVBrpp
uJ6nahk28nZy6dSps1xVSUwAf0jgCPpehgeIrmpSIeNmyQ29p0LFaEL7l/SucBoX
kHfAe4REdtRcVPSBarQppLAuaPlFNw2TwnSZZCsvqqt67O/XZuvvMYG9F+DJBTBO
ggQMXiRfev/CPSMNaJY0QJL9Rs9evzjESUuHqsEPU0LHkB6Cr1NIXG2rLrkLrnna
Np9KKetzH4C2VDGQKA7C17r+ql7CdhsnzlTXK1Qv7veSBskKA277wLQw9cFghfbX
vEODqt+XnpdQNrrLr47/9OhxWWzEFxSRWpLIyT7JWE9s3QFOQpOhPw8pnSGZX/+j
fTdi+K2n1JdavEOXxyArW9/kXDE3Por1WVp2EnS8YMxEA/8y4qLvQkHUmYXT60d5
Bc0A3qzFcmhXuBLTrTLAxCgDmZ87UWaGO08O6705ugHjthE2gzv3Cl8n+BJFnR9S
wrJjNFwNu+wuuK+YLDO24vvyIt2FZdOwGb987nJ3dPQCsAEMTQqmCeoYLr4NcfH1
RmkMe7m6D1C+76kRQjx8u8HJYDuOOqrdF2Gv21y6i+1o8sSfl/Lgw4B7djsMrP1X
WomBgPoflCCsAaGQF6aqqjTwWBnWkusT1MZbbFrK/XvPZqOaa2kfXjfNgTYUynvc
pHjBh3QAU8ndYJohY8KxoI4maxLCV1fzXdHhr4oBabj5HfBEpyHim82yTuEdX3xv
vZSxAvMsIZsXgPz0jNScG6fMeru8ZNlUxFa8/on9AZLmdskRPGimaQnhnTpXxYTT
fqhyvSjfMrHsXfVvXViCVUdQWcISjgQeNVZjCmutBCLlargY3R4eJ097Vf4zdvJF
Cy+hFddX+j0jjtHLoEROtnfJlXB4eaEnV1nFTLuBsnjk3LHkTdRVdILloA6ZpIy1
G2keF0bgg26URepFZCbikw05NcuqsHqMV9YyKz38RLQt3ZJZkf88e03ookEzAs3B
CBhmYmyZqYATPdaWFF8HPRnoRdZ9ennDomi1iVpkjJFy8UC8TcCq0hXKoG50eebS
MEDKcxgNhfRWgdd9ZLXiL/3BO0Nhtay+x9horaXPgPTPOzG9xN8OMV7BtQFxIFi7
UCA4QwhnbMD7EAnkF1ZbT3MlG5cTOKUE1yWcV7IzPUwFSV8qwjW7toRbQumlBlLw
jZ6oW+NcKOYO4kXlO5bNjYovvctYkWINKGX9r4MuwzdoFi2R5JLVmQh0BbcfBGth
GC3CEzX+38KaILHpC+sOjgt3lcDsMtD6XgEhNLyafc3jJyamhR+QbcuQtpcs5GHD
q9TwJBjUw8as2o5youIuw89bpz5D5OuhSaIQpAywB/rpVnWPm2LoFW5Mb+zxd4br
RjJnmibqBbFauut9bJsuLW5dQnk2jn0A86vDr906Z0KN8xy1A+ZR6dEUm35sLwVL
z1gP5LBPI0yh4Su4rB3D6jnGsOnVGqEcAbDKgYvkBdgt8cc32yU01s/mwQ2bmKKh
CywThe5qeSPDHqvGoCINYNmuIim8trtsdHVEOWJo6bDsm0OVO3cpK8G5uA9+mCIU
QYtuAFtJmyF65k46eCSfH61WuFYw+MiXSR+Vpy1tjGH9RYAWVBPmpe9jiaN4z2qW
vF5VqtCcqVrdcWCAB3rZyB1Tpk9Ly+DMU0c2d1Fj37cZlHEQPTzen6FqkQMjWqYC
XyBrGqLOVxO+35ype/g4onR2XGv+U3OODwkdg/iRNcXvghsZ/yqlvnBqRAOcmr76
2ZYwdiThMO63ALlgoZnEdqE7NrNmRlpsq4o4SctCNXnSmzlNe93CpYbsi7Z33nb4
ozSaCyaP4WoZGDBMlduEFrpLWfE3DI8QfQaFwa36pBvY6uIv9ek/qCidtXtVR0rp
6iZMNbnUeYSp/RalwYTNxUsuAlQijsvRKFVS3lMmf6m8iXTF9t+CHQelWoSRSK8+
X+yCoG8UY9H6Q+0tDlb6+asNKkNu2Usqs7wJgPlgeiFmWKiXhm9wRBUUQPw/vjD8
MkK5HueU5bUNlG5FuWyUxGDKMAVOmncOcXReEH50HszUnSsaH69mcLs5a1hD03mc
9SJoCDbUBRjRN/PLUEJdp52Z7gT95/vsxDVypMRE6zqg+OC/v7WrcVhBTXDGtl35
J+ssr4d7tKMR9YmwlgmX6V0nOmSJbWBOdQ4T4/Ok24zdyf8ASj6LHagQSoxkqcvj
vaYULJ+G4ZfRi+VH4Vf2n/c0hSmu6bZpvRoG/l+T8QmRaGMklhhSu89dDQ181VnT
9WETH4Dc6eyp63DPEEFSwQrM6LMDeksDv1WT4rn+QJ5QuslrCFv2ipq/bynGTuU1
hR7WId6pVfAkckZoNwpSMtk/PnlHYkRA0zj89PqHqgXGdnso6lxdsKksJvl2g74g
FQzMhyqKnbsiP7LxLKmJruucFstIW7ztGM+BTyhrgUT6it/SbPvBVahkUEkNKWPJ
HEaXBAtJMtrWOmFyuX5jfCtqirjp7RBFXZTAbVFuJdwDMvU+GkzWNOvAHo1OwGfT
y7K1YrhZ1vdRULO7VaA0Lp+W4APJwYr2AXKxVZ9YWapv7H8+20+kq4EjZUua0nB1
GmC3DIk1gpbDNvKmyWLSHQ72bHwzUgtrEZyth8Du9VmWwBGOETQx6ePK26yaGh2h
AbbgSbi0NKyYVbbMC6artUVJKw0kKzpGqH/wz9PWM5twIc7jMgNbXx+WBlmt5Lfy
XE7awKAh64hQJVPlXRrX5EoemjN7/gt2HNbMcU/XWy7Ht5KdaYVf1Jzr27bl/g53
WtxalNi90md82kXsS+MPEuaSfFdO8nXH+n2kvz7bUFEqu37RXQbzuKYxh1YqZwLh
SzTsD7fH1+i+CK8OZx9eaRGFSNXU50dNNZ6KBTAka89hP/lSegv61/hfmdqtRDGk
XnRpwoZidETTGuuVOjmKkluT3Sp1jMench6mSYg8YQDyxVGkGxwtzRpVn5yz8LQd
vCYilWHQbRnheS0Tc048aHl6Aw2wu82puXjk6ZLJGE6oO7pvTX2Syribk2c+Q0kB
bdbiEUOmQQtWAK8rlM2zmJqP8A+lUskbVixuIZI7pyOPQro9J30o4CZ2H5GWO/Q+
Rdo+xNgcfLeWl84UOWL/+U6SB1tf+/Kf+ZpF96/2zZr/8x+iwOS8xBk7vb7hwO+9
dxO2XqR3ZGTk0C3k2WgwiWaR8YOu+djbsRcYCKL9KGhsxTAz+1G7UwjVpGq/6w0t
vYKq52E5n2uTl5xd/DpNZHD+nbIE99DL9/uhCgQtGc/RK4506jXfGbEqyvP/nQx6
mkOlPs45lGPh9mZ3VVwgKoIZpm2Q2ngQ5Rw3hmtMqNuBewv94vDPBaVF3VzcQh6h
TbSNUHuBaLSh77kRMm45R1eg0RDy8K6tL8PhANwnDIIEjcFms4DzUUC1nhtFakrz
zbgVb5CRcfkrrWRsG+v8nxOeV3p+KJuHgFSmHgWO/pLxz/4hrNlYatgtR5l7OFWl
xswqTzPS1pRvLcA3BM21Pc6S3zKdtnWwVDT6Tb59pr1nTUOcGpGOD5FJIyTwdYN4
chMKx60qUSh4FSsUGhScVE2wWojodGSy+koDjboY8gE1V6yg5an2t49FdGCOkLsW
Zxcnd1goOVKJEbvct5EoQL/qW2ZJwMzyLeQkBWtw32hSf+HN/aY8HMeDPDHb+nBm
vL5AtTXMYwPCCbb20EviOShyrGrbehD/oDmk0/t3kwW7dbphN6i3d/d9isFXG5X5
cS7HlxlDDYDlvYwOr7LIIKoorsg8ner42QewwWi8pvk4qoOpXC+iyTwmMeZq3g0Z
j0pr6vVGH7n35W8s6Smt+nzGrfak6U8XXwnZRykwg4ANcSaHwQp282LP+YzFVex/
uJr3NPwxkeDsEyQB0+pl/ybbqyDoOZ/MyBzGj9LdxZmLT03juhdW0irjliuIA7MG
EXGuW8u0fZIpVowCpV100Mqnw1Wzdlh249t770E+nICG8W/ZtKbgK/c1/Yq3WkKb
Z8tr5P04KIfhSS4MuyvfA2afkS6VejZk+rY4zv6Z7d/rMRvT1K4PQoQ7rUR7J4l0
zYeKyYbi9kiLI7yWax3IcoljpB+LeXMfY/7orhZGoNTp/fQoSRZKYHF8x1SSEc3d
2G7vkHiIdFX+RDVcnvxcmMUCY82i6HF6bRajhPlVn6d/eeVt4eklBcHxgabezDUD
4iWAe5vhwZ46HnGdLu5u+QkkbgoSKiE1xhuguwtiVz3KGpxPp6br8vnE5XYNCmDQ
1ZEIYMW1TRte0xhqBkYU5Pnoyym6SCjWFHES/BXLExNytF7K7dJuD2BRNb0QRGPX
fcnpEveTfxqWYsYdVQIGMO5idyOJRzRexmPVRr6HnuHTrac6zrNC448obJf6aV7R
ysluy7NAJoN3YRA4mqMkenZfFwAS8KxVTzR8vgvX4FHL1fivPBcg+bDAUpcDIu1n
TIDQXfDa0pZ1YopnHvLdbIF7G7AbHCNifp93XYtfRydoMzBZ5B8FTWRuDcBa91j8
6TIbYBpf6ea67qVgCUbsZmxi4Jgd7u7TZGTBpCrQ/rXjv3DrBzZ+/lYsK007idWc
Ywj1blazhQh5KJTnptGJlEP89MTcWF99A7Nz6HcCKoAD3RTeqW+rJE4YEcdL99hf
aV/EY8YtmzfmhECdNhLQk+lULn0qnIHairYLrjTcRijrhEKTbvINCNASXtGkxgZv
9Bo58abVtFgA+2uwdhMYiGh4bK7SmQpLCjkF1B7Phf9Zc+iGdcFDu1i2wMEplx8W
Vk3RgJZH4Am4Txh0RoKPbycvu3n9ConHU80mkLzkHlvWRcmk/KY8IZLqQkMqno3i
GVaWo6OwzwmDXDd5D8mJnFni4qXllG//NiENQIHEJg1XKn42+QwQk8NeZ8exx+JP
+ou+9HT84SYg5XeCAJyOkgUCsQeFCu4HQD88d+1uIEWMUasXc9/0gvXeHF2QIAGg
NcbQ+IGjoniHWLF4ONaD6XhgnejGmO39t4w4OMDZeZxwOxjrrYbLFE4klw+D2+iR
sULvmynZzooG3fmLQG1UbyHD9wfElGM0u+LadIeixdxucwY9Pz2mWwXm7nHQFrSe
KZhdCejP7Zqkmc/qHzvh8s9eTbGmJfcVfR4K3kEFB+YTBze3mIX6pzWop9WphrlE
3AexQ5c0cramCfEY3FD+wQpE35jRP5PMLneYesdH+dIJt3G7PrfEVejCgLFwcdm2
jH/9Tnt7n0Juk3+TnHE+wSOFTdGCMMXUHltj0k+ir+rrupXUt7aP9lePfbnLUJQq
ls6YThZcoc3sHqmJsLCE1cbLE8zom4rfCR4ptpDvq3tFfgaxwdeBZE87IKw5DUkS
ny3avfaQCUY2/0Eyu2FIewa8bGiwZM2ERMoUby04FsT97v5lH3O6unmAMGXOKvg1
WJhJ+Xa4wBpY7eP92sb/p+VVqfE24GcnycEOnaevbJidUwzHlVsBI27rQB3gKNd8
FPu1+PZuy9EEGmPdALtLWY1WYn274FbLqgHdv+fR85J71bC+Igy8Pzi7Htea/mvm
tphtB3MWL9I5YdTIB4Wede7xh8+iUhnkvi5siEocjywO0BtN7di9/fNpvADN5Pbv
xA8LibCUpPVA0l+nngRbxNn3gr9jRNlS4TNmQfA58sjdLMZF0nZHLWfLKRPq2e2w
fjKAt696mnBuDC5KK2LmK0fYiknJn5wPqxgx/ZZF9RSrfgMaWz5gpVyNzmhV5WkT
/vM+GASinEQ7YoYa1wrMnc7ylnCixi5fI7WmXauqTIrCAISABoN8Z+zZQcWaSKDV
u2/no18GCeblLFC1xPV4V3V+gxPTL78GVVJ0iXEg+DOe8CPaKLXpQWvJ1FCgMtF6
oreXL18GXoFSORRS+2tuigsZvxelBuZBaCiL/XobjsR4puvhyA5KlYPRP78tsRZo
/mo4Ii1g50tcTXDW1LEyA3Pxnv+5h6c7jPysEZh5F5REtU2hdywL7SFnG/U2E2vX
4cKGfSAE8JrU0TzGMmckUFEUj/oHrkxP7aYV2iYpfDiIw1W58vS4pxF2kGztM1Yo
8zTFjcc1IqtrVpmJ/X5wU4ZrstNQFDURhOvUKZlphyN0qrS1iD0iJoroNneFoN2M
4IV1MeMTTpgJSmBqOEl4esWd5mLbmJ91Jz6XcFK4ams9Fov87RgyeQlO4OyP7J3k
9adMxs4PP0pAnwasekGURWyFxjdut4CwxgBQDTfbQo/xB/qfjvScoxZLyahv9220
9gEYYSu4HaUfAVMc8C/1tbWRWuUkNs3bdUeRnAbqEimYc3+WKRkB7lDlgAYG1v4O
oMqT77oEZB9KFFwCRWoYdDtnOaBHXklNLjLer79mCrlVt4vBQAzlI3Y39X8HH8oy
kt31Ek/Q73zm2du6Fx7BD1Sd0Byspk1brgz9ZmO1Rn7Y6PBIx3AMs+5TMI0/BRW1
r3OAe7qm/oRa9uvqoyjGAIviSVKjIm9GVJuyLCqrnZkHf6+/SGWHqZ7FlDMi0Wp9
hTt/iqLKYYBiXAAKPBL44vfOkvT9X0COTuFJP8nqBOXvfzAAsD3ivXV1mXWM9QUk
JZob/XsMQ7NXF+F1iHTM0XeTWb43+tj0QWbHgY6fSr4VVpqdk+zmdNuIM81ze047
qbg62Qx3W2oGTrsBjCQh3pqkSosSULfAswQnLeJLSCuoFJ9Fcn0odYapGmynavkd
Z/eHVRaqraeqPQqwaaY09h110agfkVW5GB1pdQ2Ooa6J6e2Ua2J3oC0Q4icq+/f2
heyUMv+pAkTEYjTcuh2HQDc0AABdX3WBtzM5PUB24kTWtbRcIBPNhO65rd6yzVQA
MHIwWnMQb6RzfPix7Q/fZytVU76em8L1L4rftl2yyr58BntjL4ofOmYSlpY2+Ieg
zeZmnh/qgji4cqbgk2N0xSS3TNRz3s4a6PNQCPFHOuM6bmRBLZWuGUqHp957qDcv
Vsu0bBA3bh3IPWXL6vx5lczPv3J2bZvKgN5icac8E12TPb4bM16VLUtuS6Iju/ew
4md4waECO2lT+0+jc95geO0lt7+BbbhQMMbcu6eAGvG5KRVvS+ZXopAe0qVMinPW
Q3NeTLX8naCkMGkbYOyQeTewy80WKUd5OEKkuPQt3qcrtbELNoIFvZCD5Qs0dHub
rnHLiai8Jx0+EmumRWFFi7lEP/Q2731yuuLUvDND55DCH9gD8Jpwp5TGjfRV2cZ6
kkOEoDw3pupVSqaspFvEoLbPzmRCxrVTD7zeWRpNP//F8Bd9k7/HuYh5feg1xERn
P+geIlneOS1Rdo5fNdGbcD+EqoDBhpojUNw1WIGdsLzH6IKqTM3+NaIKkBa+dwE/
JP7XMjrmQgrkUNVLnhTZ5Tj8ouoEH+fQz/tdCOoUTOCkmm12SLAr/XAgiZqCb/Cr
ymwP6O/Ka4YXwBEUKUC8p7KCxw9JxCquk3JiMhl0ss8iopTgyAVU32snXNVcD5VL
ly4hmLIQQtFFI28E/uOO8Lkuqavjlg88LUtOug3f7o4KOhgIQDGvGB2nUX2Z/Q5D
z54HTM8t3KvYwvO1wWKY2aWzJaqek6dMCyS9+kRjfR2ohI5rA2FzjLovQE7IoNiO
DQbDmBJbRHP7TaJCf0kAU9WytEpW48qpQ32KsJhM5Vpci0H6F8DoxrrhLK1Y3MIW
8NZjpUsRBDLKbsCcoLfEEJiaitQqhBn67morICrJzp7YH4k2/I4/arRnYoAMF+FM
GFGBpe6e38Qr7RbWtA14F5l35AlpB+x1KMQJhET/KdJ/lYRpAAgMngRG2fjDlEh2
R08M0HE1zvpOJ9zKQBujpgdRx81V16pBaIc2eNov0zeIFUbwQSdZ/QwTIct1zGeL
cEL/2ZxGFhXYagac/JM6hvyXESh4dPDj6lpzWN6KuZtTBoiha0S2HRGFdJz2mfU1
SOuRiBXZ1rmVg7qUjF6qkk2fQ/vvwhD5wNyQj+rfbri35vEmEz5J1iGmZ5E0tCUD
YiJz1COBCR7zwW0w16ZfdTWxiCV7GfwQGIfKvgqItS+KDfLJ10Z5u4egq/YAuuti
fJH2THygWgJXRg21uQo4+yzhzPjIepmJjXkEIfFUJ7wRDJbKnbaSxvWEUp4fZdq0
60+ZNghZHoH+ZfOIVLr/bCgPq5GhBBX8AElfZX06+Ca5UrOm1BK2BjZv1N1NsB4j
vb4GGgtUTmrxiBWvSelaFnXVpyy9yOoRL0uXHvANgKTK7kgBsYsd8xNK9X7Q6ALG
BtCLMQVKfsEyNFCTUwFSEwjPKMLWEW+lOVTmWmyHUm6eHgpBAEN5j7PXMtjJj5D7
/3qWr/lTyvTKyvr+6iqnligtQJcUG55jXPgbPlQvvI4FpXEcufhxGSpciv2uN8J7
3aNqnTDsMcCrqOnQyR7GwpeJngmld8q9NuWiLVUi37l11CQe5VqIz7+8PnMs9rB2
c/QDEO8DqY7pR2McvxLgDcYUeEJ3fxpAIlh4cbiAzBbahFlRM0iY3WydHXicWNJl
dDgO5NJHIYiirjjiqFBgXFUVtsgiTnJT+UdU2yiDnrRLLrMZ/iA7kLOxTnhhuU7J
a+CCuQxdKnOo+9iS+40dgWgfxkXpZXLDtsxThpRWZ/N+S6OBKYp2Li0kS5EygQkP
Q0Tj6DfXJERVdV/31RAXvXerIV+t6pZyc4NedOL8WkRS5BkZ+/vXbRfb01Z3/nfB
4Z7mrsan3syIHsQqBTf8r91mSLF/ODjWisWX9vbMoX9roH7i0kNEuYLHwhtjx/Vj
eJNXCr2XCTEJ5dXKqToytzuHvc1JutGLgakRlmxPTnC2ypjeMim0rHx3n6NCvOsT
7qcX3v7Z1yuIZa1L3VtZ0BYdZQ+1a39ce2Q3zB+HCyEi4rZajXfNMOg5zHkFKAOV
xdBk9NhTQmmC4yy8Q5UxGXDFTKfMtgak6uFXLY/kyIZDatXQ8eDA2mG3DgBDFVCr
eN0GG3tETXbfcONDkW6ud8FmTpi7eOUeoG+HAN5re6MOIv4kyrzwJ4pDzE1NKnx2
ouvnFqsPhv6Ml8CAoOxDaQpzoz142Kyx3Lm9jhCjTNBwoi5sw026VmSvz2NMPtjS
TLomfh3zV+9VZTAZD4K/FXaMaPvjWnS9g7vMqpsbhEVYrwimkCaAwIXK3XNjBy5E
gQTLDM4N98F7HJNbNzRmiXCBY2K1Oc5IO83ZkyQc4oJunXT9kvF6exDHB45aPa+N
r5M6O3L400PDoFLqRfNSJuL0XeenuaOKv/vzwF1m5uEh51shRXor55Ivos+CE5yT
4lvw2FJEt8qS9XGF+7Z9WdqI2UYmjMbcWtFAhFDWxFZVJj7sQrn619rFrH/csOwm
LzvnFyTB7b79mPzCUUOzThWaJfx5Q3SWJS6MsTRGvHNL51MLcFI4/qurBeHDtrZR
fbBk9wn6SiXNPeRuDMEDOD2r4VV/504j+84uaA6cJyuaaqTLi90gcvEFUrsK5DrL
+YGxPT0oaS7K+Vhb2kM4Z9jZkdGS4O9DcAwqO08s4uahwgYgq3jOAkOL9Egw6/mh
juxHY7vKV3d2oyuhZ94wnr3P042lmX/fMI2f+OPOu74/qg//YPLYC4V/xCuXFdDe
nA4GyGscGg3UXaMWg6yKbtRNbTGorYxZ4dYu8s55gRwy9sPuelJW4vd/2cuOWJyq
DXYDzW2nh2hMY/KWygTpSvEvjjcetonl6HFX6yIiRIGF7uvRhYh82WSlXv6ip1Lt
jouipwj+i+ddSFa39YifXr5umqG2VwGrHilyjr+ILlTVhvtzBZ4EC+UB+uXBRK8T
+SJvRu91ZFzCwpa+T9J8yKEzYwjGTnYri+JH6ahK1OE2WtcNZ0Jf7iwbUw+1sAlh
maL2t5VhVlU9zxPbHPi27U8RcQKG1ljvW5ffgdbd4V7jhLF9U6GTDHywVVbN/UXk
aq3/YuBvTl5C1j6oGcjeUESvSjKFoLO4sewy+UAHErAaGgye7Jil7LTE1R0GDEfg
qek/okG6vjiBVTkMHIrlbEtYx1EG3lr4h8+/edqKfwSJKyWxG7D26uDBNuIL5GYm
P0p2yKJ1APns/qQMV017T59wSXStHLboDNn+S9i94Y2rDI37tQmARn6Wgick6Hpt
QPIWvkjE5gw7D+qhO+doIySQkqSAqPyQb41JblLQezL74DoJyw7p5J8Pyk9Ojbzn
XJNRJPYVEdtDAUtYASIQD0X3iWknmDmYxUn095wLuHqOQxkgplE4ve1MMvhg8DJX
SVD4wwjvt6QGfHjlpJpabaWujYXSHvcZboIhGgUgjWZ7PLApyDvLRxIampa5Vzam
7duEXQ+PyC8+wDiwRyqXTe52mHD0DfDAcvhwsGBtQs9r36E/GFaPl1EFWgEF3dTs
0DNXmg3WlzLQ/05QHcbvWVGv0xhJzT1ePoQbQdVNywnh6ruMRnbQIFiHI1Wdj0mI
tiVPMkOUbtmDwudjjd0sGOhORi9SXt5qmcb7PuqODk+n2BZbc3UvSYNvS6y8t/uR
xiD+MoEgw/2/MLCXlszMXX3uBZy5dwMUZ/SBGleUgSCnaYpvmLAKo1FK9pIvOa/b
r6Nvm7Z62N2xuDgozg839auHcsynyD7YvtbRnIDUZ7zqrphATgRdhM+LAk6BGQKq
09vAYECZTY+KZJEiHLzHfhCjwBhX3Yv8C1LgC6H+f9CzwhNxw4Gcwye611dHA7AJ
r+droU/lCLmV7t3GlDei5HMBLxEqNumnNR9IbR61ZcRyIsqLo4YN1FYPZjzseX5x
aVKVQjMJMOsZ81Y8395pKQS48erOZLv0xprOGUhXyyFxfzE/qHQjWwduQcciJtln
Nf3PPJE6vEPknKG/2nxamhb4+S8ed7z5OVm8GcK0pw9PJ8DVFrMEQ5Sf4A0C7Of4
T4TNAmrZKVGlTNAaxLgo68s8jPY4qJBnaEa2D3hBU1MVKrkg5nuaJ/i2v+M6w/Rl
Xodz3M7eT/T99mzs6+z8Yok74tdaaW5Aa832S5JymlOw7ulz01V5UX3ZUXXKpPTI
BRvODZFeq3YUl+p2F4nJhd605xt7WHisu0JV+jN9Z9GaoFLKCAARZYBOctb3OY/q
y4PFb+oYI5MREhWYGeoFwOCighW4+b6EDH690Cxj0lkr4d1ytNAPjCrVwtcm8zxy
2Y2aVQP/JdlN1LzABMHQoWv6Wx28GxSiOtFnRIKtEcUKeVKl0d6UfpQXieJs7qSI
Xed/M/ypsyUCw0MYqCOuIyMsKIXbsV60JQ2FdyFANF3EARctl7aQvlViPUFcHgZi
EnKR8g17JMGPDc84i6qthEIxgQ7gVTM/bTFRYmD3q8CdyvE+inoiaG5NK9ruftOD
buB2K7a8wcpa2gadLsQ/5V2TvkVXj+KebcZT4xG7iH9jyUb9VFNzChpAIMFRLNYg
y6CGrVIMVJ7La8fua8/CTP8Q4XYL+GJa2yrFgoPFTXo5l7pTpRUP0be/8giY1Wd4
Ybxe2IyRbjWoZlN/UgjjjkCfpL+DiwMGxz/PD2AZIYiMkRnynXCVzAml2JMboA3h
K3lDYu9iSHnHy/UI7+nbgrDFTS+fy6MMQtlPwwPEyV6d+PQ7AtCjbK0sn1lyjMgS
ToV4UTFMSvWflSJT6JEwoCBQQfeARplvIQW5nIhoHWwflUj4/g9Zn8btB1HJOgTV
A+C8SQvKJIVBx39LK0NIF+zBkur0YhmXZA+0vYwq33z8m+mWLKangbekZk02BLst
oHavdz7LejusgqxUrLQa0o6LU3b3acaPtfTHxyVJHdiPtEVEvBgG9ysWIoCOobP6
UVtHyTXWrXvIi+xtOQfrFJSwDmQ5dFqJQJ/oZ0/mM4CDYnQPSxm+U5EP2xUwvQQW
PtBPXgxnyOKdCeaDrNDOgwhMBNVAb6PBQFIqcXGqUT1bEsX6Ut4Kruu/AzBsM8VJ
p+H4V1pVDnxcL1fX7c9pE8YJRne5aI9Yx3MPA+59HL1KKlTbqZ39O9FAv3TTV9q/
oAINm7r7W48hzVCYQdozHaUNKMv+hBmhxmSi82sS+8SMsZWTdiGKASb7HBf9MPfz
zKm2cv6p8zH49QS/CcTNNS6y/OOOM0B1ouf1DtxYl13w65FpT4WAizdA4lC+8X1V
PQRReAemm/tmcldMWJNiV1Z2NpY6NUDLftvGH87PgkLtMmc+D9b0QoJAmoub84EI
F1GARPpRPnoWV93opNVWgjE3N+sfkFCpavzLVrwNatDkNqTX4jjv0Hq4KEjI6j3K
rWaEpThX9kxf8qu4475qjNHrgu9XwhnXiDHfkoMcf7+yUuuPROszDxe+gsXO2ub1
IByJTgapDJGJxHIhfGgrsu9Us4sziDMtujnWTD7sQcDjpcLRA3RRocANOkWBGHLs
i1GMasCwvqWVELSLG/XxGT9DtCB9KYHj4QsoQ3RFkDieqV+AbYs4WwtE4FyKkRdL
r6b7WxcLaXL6kBBZhpn9wqZK3rHM2GE5YlNmsiRuhZ+zx/yAw4b4iQQ9hkh/WPdy
08ns7wIafQN0OPknqxj6AyNRn/wsdSZXDLXWAARCb3AZ+ycBtQwrDiy3Pqwb4cpu
VdJTtmHMdQkcViC4kxOJ5dIMZNEqS2fjasL9yETtWZKFndlE5AZ04QIO2SCLW4+S
H6zeCH5Cvr8WEXTvT6gietvka1lB18r5vd1BVBl0di16/vrE17kU4lSU7ASv+I7Q
QfGlSqcIVGJtQ2uPPXkNTdpiwJmazAZ5w7e0/7mjCUjwCZUZUkhKrcvrQGe3W+ZR
kTQwEkPOd8ThTOXUDKVGrCNcOuJoKHlqPqyFf9v4DKALLY4z/QpUt8k1uiYKuf6Q
alI63WjjD77deazJ4YeWqtcvnxBjSw+PhV7zEHydKEd/1gbCvHPGQo39nxWcIxTM
4wsSay0ZzQPdEVVvJXQPOKCC0ST55JwA+Bw3GS37Xlrw3n0JTTzEx5lCLQy1oQqY
6tWvlJ/Fp9MZzQOdVJVrxYpryOEr1ZtOToMbrULpJabl8yO8yCkgZv2kjUAOmafT
YPa8bytgJfIW5wOyGcHz+AGgVh/ie0yW3r52Thn52Iju0flIRwOyb95vO+4EXcl7
zsF6OZl05EmIsSYSxh7JBTzJANnKJ6JFTFq3IusYuCYD7sesIJ86p1882vaRNroT
SjR/WPVFWlg2Zj3C9o7zeE9fEthdX5XVaW+tpKJAfbLXHiUIPG0SMu0WJLkiwDzd
r2acJm/MPvIVx9i597cg9Y7lgDqQ9S8RstrSlC6T5ZMqx1t9Zb/nNor4NrGIbJHl
0qVueSmu75PdSTYBTbvSQcaBBzZ+minaUAxIx8ajGFD2A2f2haC+p9hT+Upwvdor
oGsFwZGEWYBRBdMuDNpBpjDMcbtZfzrgWqljwVNNpD3B8utf6OKnw4iJ6qfX/AY7
5zyaiigBYQVhv1PNWoqY1ha+gYaVXfEpl/iKlXRaIrOCJ4EEY4w0h1oZat1o4ch+
X9AMqeEzciEUUB1qIuAu6U69gxhCouex57pq/S7EpvggT3m5qrwLBrykcxKxpKgj
rR9Rh26rSZ2s3kpjaZ2SFK0Nk9kn6Gpk9rvdUeUGjuR7bn9uWOoMiFzq+NV3hhO5
F1JCQlHp+nQaUlnC69exPohyETvSp4PfRfqbY6G603AxaeGxkagZkSI2Jg6l7C32
Zb3ia9ftjABjaRHkpgXazi6OiihHMOTvTG5v4r4FW81RU5MIzwbKSVEWLFGSjxp8
uUaCW89RXxmLhMcm991TX7G+76JV59D28/C1S+dMbrCo1usmozHQaJaBoQ78Zu4A
gbsHvuiwBOBj5ucElrSVigT7TfUXKB64x2z26ajdqYj0Sk7G/TLJZGQ31b2v/ixO
dPw0dRxnuQhqj0UPc8bMfbFrHiCLvL2quGagV/qYssa1o2HudRy7c3dxr2zXOhiL
ktY6ErG0eABEJ475px2SuYNJJZnSx+EeRBycO37rCzCg6zOr1kihSS+F5sLRd3tO
h1CtsnXGlsWaDwl/+GKwnoAIwUPfcrqvr9A0L2vojY0sWqQTujEtBLETRm2dNSsO
VLy7Pgb4kEE3sSxjpPNlwWfTyaI384Ycip606auynbH+uOF0spfxvKxyo6MhPQWB
D2qF50X/gR2GoEYs8f6WVw/k4AF7vp7mQ0BXrD7KEwG8Z64HuOcmUf9o5OSslkfe
YWvtH0rQDc6OBbkPNXfQ1ZZqyQyAxRc8KoQC7rbIseZbDIsRxGuFoZ+JD+1R0AVk
70QZCAVx2WzsHxgR6fWmg/wkKMk8oYXgGf2zn2A6zD38/R5J2zz02zxy5gRcBLaU
nVvzmr1gzgh3ICYjTLq+8oZ9AxCH4WlDiaPmcOjTggrw0gJChtUNeWNAKUYbCfk+
EMbWeyHt+2YgV2RzQ5X79MFvb8DV8375xystqMOvJMvLPz3o4rXL9C9YeLNKoyBo
M/QFtIQZ6x5dA+372TmNTtsYOYPQEyT/E4ee3hE1lf3H9jKktk8vrACcauznLKw0
sYHYPElMys7F0lB2UfZe/JDNrVU6AU+jqECS7YY4rm9CxycMKFD+rp3oADKjyqQb
6YZW/V7zvfnMTEyUJoVRU0LRWrptvxSibCGJpMNjWM8E6Blws87QmI/YxlvCgud5
IVQKlMWDXRwvwF9Q5UBjvvSte2T3+DDleORdC9flRxdIPXT5WBKo8bxz5zmXulmJ
nUnsbHW3umrTkcAYVWUyU+QzAgBEE8g8eQDiUkBDyPl3mx0s0Hn27znUXberVFBR
+7T/1MQUvV6lhVwnRuH2PrPUnQ+ltVdYUft/on1Ur4z2hsygRQPLnEzOAMvp6CdA
kgAqmvZyLFcKtXQRfUX7tIRQRsjr5durq64uMHIi3sSxQtiGFEsmux/wDu4OAH8x
gvARmDnzJPZMuB47iTj99yNDp4tOOeXSXFwNgN0yYjnHVim2Uf8tePgQDOABte/B
+T01695VJ9w8bldUwFxVrPp6SjSwhHeGjzd/qh0fYV8YIsvYRdNG8Ej+ld/z7ZGh
OmKvPB/J+McEIIhyM8obyc+KiE3+zpEVyzX9XKHzHr4VxqOFgrsfeqKrEk/2g9YU
UWGKZkRMgQfnZumOo9xSCjdRaUTTv4yO7vE0K8ItXEfihN1b0Eos3Qm0W821azX+
1We7EgFa3uuLNFNnsKELLRCprvqyIvVxxSfuZ6ptx+72BAS4UhfOVcZqWVl/sdSS
aMpmEKEoAa3Dx7deR2PzGmRLCl8y+bxovgU85vkmPP2EuUanM/xH2ycKs1PIFPMT
ttEhS6E45cD1TFhMB+VdDHYuMI2EtEm33hZH+lvzIeKOk+FGkE4ovGbXz9OKdIEB
UdoXyGdHtoyQ2Yc2t6+2MXHF3nIqXAl016FLbeGvUpZSp26biB1cT17IOsFOKnIh
sdb5kqHJ+tgAt6Zm+A3B0R71fUaZtVslR4BwEH7MsHD9l4WnvmwcCkxGSvK8va34
i/7j39muVkoVPffoKBva+QTAQxk6LEIE6ZUaIG0XoLoL+3FQI04OfX1umm0/6+vx
z3u9Q2Y3giYugTvz23dGAttnEhMS7HZB0uUpCEMA121zUhoU9gdfgGNqy619c+S/
pjMBk15WYJBAs1MrWtlL+ba3bIYrI3Kbj+ZnI1l9nBV2U86/3NmazrhKOTDUE0k6
dpCNPjUSvuEWzXKSQQk1FAmpoe/vCo0ufWwESNaPN8qloujh6AiAJtuwq1z6TZpI
/Yc87XcGGumSRvp1BLvjCh6guVR59NEqdPPHAYiymmI+VmwnOevl8DiKDaq8kWMT
6Of9hSfD4Suo+faZZhV8/KKI/OOOdVDvsZEJOj+VcLiEyMSS5t0TdQBOoyjmreAN
gFQ1tS+8FyI2HK0IUABIMBSadRlxzUBpeQrs1gsaA6TKDelBHPVhui0MEsSHvv/D
zIzei/m5E2+SE5T5q4xjucM4UNRZlE8y+vjGUrjvOZV+r5O/RGYz9+5YhN33bgDH
QLLQdyNbZHaOEq3TTgMdh2AbNAP/Bk+/EdGmb0pqeK//OGEc2+P3TWxG90pb8A+7
pBYlblWSc8adtNCovOkFXmmD89wrz69HdF4jBVoWorK15YQuFZBruTL1QM86+mb6
N9461gyjJcO4GUqQ1UaGeO9cSZG6bgV6afqzvym4rzaxPxrpfZNlj4Ir9VAaf6Sl
8F0Ru79yHtjIkDkeGiGZD/khhwqG/RRATlcZZwmLJE3H1O2v1RAGuHDYjwtrcE6w
GsHBK3X7cArTwkbyJJIHQ/G02/L27XwKv50CIefB4mJRJa1VGcGBBHm0qijvBZVI
xIgioWx6Wp2M2ZgrrEIWDyj8X5Vv8qb1GQnjS6ce5eWmR/IPzj7lKEehLlFGs5VP
0y57SQ88CJs+7lHSlrwU4YzeiENa9XgstxLttKPg77c8Xi2iN7Ei2AaZrpjyVcwa
CiwQwMcBrnZpfdJ3XNr0uIxPtP7iEXP/EprdLckVeVQ0KaMxvLzCkmqSCaUbp2Tr
Ir+l9J2xFYwd8RUJdaRodzlcO4BPScoi2EiDahBBvvWKjsmgXtTweX+mZSlcpkpa
XFyW/gKvpumoHtI/mf0laXjDMHpYLJLbMPUZsRaqIMORKebnVKmF/h54UetHj7Vq
RxqTFrCxJmqiJ4KIX4Jvma5kva/yccgNdw0SdqPfIl1bZjN/z6cYefP2UBjRP+Dw
tVyYM/MDmDeKC9PmzuTu0K5nG9GLUJ2fxQDnouZ8T40JDE1NXXYaTz52Oc66CD4A
+Gpyv6twBZ0hgl1+ljbxSyuwUApgrii6SYuatBaXIIxmISYKYYteL+fwvuvKXT1e
n+MF6xmYGsZM6w8i+RRmHZ3hx1HRMQkTHNZVKCt9pkHGDNW64TvgX0sY8c/Hx/g4
Gt2nMDTLrsZ+tnTiE+qmmR5KqwoHL4eto2Jr24AQE02byzV+N+99Gpubbf2sBFBx
i9uK2feVjoefVnGvF7vck1S5wQVhln2kf3kp5DMHOvsQF+FWA0qn0LWrXVHmLzv1
MaEtnVzoL4A3hjx1LHyhkZAm51NHLywqej5j6wBPLJqZSNl214ua8K8bwdLKRHAY
A/KI1E1zBIn/6O3VGbjfI8AY6gpiEwfTGtEnLQA/DFFcj7VGn+yh1+atLo9B4qRl
E2VvEoFb9jQlqvcConqbnAXC6hcYDolVXaP48TGeZ4eTvg+FUUFseuXtptGMytOR
TPOhJALcTULFOw8fki+L59LONmk83onQLo4xU6uJEMSuJF0roNp90MKfV7zCZhvq
vD0+Ept+9thKA6pWZbSFsdcfXjG4KdjULnPCdQmqWyMpigfhoOW8rNjZMNT1RVUH
vF3NOINq7P6iCt1AfPSrctf6roOhyEnPxn7fL3qUNEZ+EVVzSCGgwFPWkIDcv4VH
EeGIlJSwUfDFtMVbgFLN8fUGd0anBgTzJOpjoHJCzYAT6VQKVCphoXdYVueoDLIv
8QsBkXxhr0F0Zshk82jcwVJ3RWAKaP4sNBHCuIIFnbvaN2rRbpEOywE44NosBokd
88soKnKDni8nww1ft6lCe1PmVnSbqhBXGyge13fmWVXY9/ShsivDhP+nTRw7YG5c
KeWQtW3V1QrJDaOBsTt1ScuO48svxXLph1EGE8DTMJ+3sPkWH3LiBnUdmwqm2OFW
HqIDvjOXns3oSov+KncRrGiJrKYmAv+pB8sSKw99flghSZP4U4Je0w09/7JeWGoQ
tYICSzeQwIiLN4Rqh4dVk5sxaifKOlUBc79s+oRY3ab92gpPOdKtvnEfzX/Xz7Mm
v6t6IbO2n9vMazRV1+0OcGVMMTm3XDja+v/+HucWzHhghU+iQcDzKGbSWC86JuM5
YitXjxpqUNqLASpOLpVmFYHxLbneq1RWsbs4JRl2Cpn4Rbup0sz1Io2TuZN6TynC
i1Cj5FkfZVsI6OK4uaSxTQeR0B22++O7Zmrwn4S9KO7XzfXI1sLX8AfFSR677r3p
LTMzsKKCVXdEvKHNRqKapxxP8mf+CgUn+/Q5nzAYMkmhXJd6Zm52D0jw+Mzo2OBr
L+pmfUBNEAuGCZ+Godju87ZQYRyDSTwqdc71GhzV0g7I1n7hTtqp84SLCWHX+YWE
s/881TF5nhCENeKmwPxbWlHvfQ/F+4RkzHvDaljiJ4JjZdOMEoJMyFFLTJBRGZEg
xG6LONgSHgD670OnH6L6GwtBAks1xVGQyY4tfJEhHmTyeFDFr0xARGIYkK4jQxjq
SpMkpASk0usOHcQUIzeDLJ/1FMsLaAyDzeDxdOt9pIYJC3EObOnfKGKbrWNXjZeP
Gn/wWt35N/5fojxpsele2xFbecUzm2Kpx7QiWxqkhrOhG0fxAXmH7d+tsUqr4t21
DxTVfWSsl5W/JGoZCNc+b8LvK3v9vs0/H0VjLCh6EQxmOQSc+sok+GMgyPERNI4b
ZIuundMMA1w2lPH1QZAGfxUp8XlkG3961QbaDKYUSyg8lB6O5mXT1+gIMTKUT3En
Jnsw3REPqLISNeD5eHwa6CihG5a3Bggg5al5W6gppEiPvx3bdLPdKY2qMhBRxkOW
CL8IhJb9fQvyRuR/kHJegQkroNfXWlBKjh+ozvokAIK8l96+iPoUquRfavAxgnqI
MvmIyjqRgr8io3h3B0uOt0uD29gPr6K6mWkKV5UZFnRvxkWoYtqu4aiQt559trlc
qkQ8QSk/Hu7SpsnJRAi5LWZQMHyKVF2hjgLoyr/vCB1WfPzn89BJQ6KhCd8jnqTh
FAcpnGXclCnlc+vq4eRjQTp3vCYhjHKqRDm3BZ/YYolvMckujLwNbR8VsERl/asv
p/DjB+NRfGwABy5LAGeDQDtojX9ZZdf89q7nw5GV1SfISDk+KcmwOZYCdfdOUGRF
uW40vUoiIbwf4igBUQ/Pc5780XCMkyP/RzA6pc+1UBdz0zS3dlTHBvM/TUfkIy5B
LnCCDvhYdU3OA/5H9enNdptfJY6zw6Vb+Gn3MCmPDpy4okjrgMELI2/ys3pjYyl9
o2CR5Rai2H15vqQMqmOoByhDQ5kKkYq5HDHCBoUQVmWRHZN8OMOVE899OqEqXgrJ
NAst7aKsr4xLrSO4+HWl0RjYRdn7xY9VnvcKI5nlGMnh3msQoWs8gSGmM3QU0JJ1
WDMuOM1qNheStonpFWz152BB/HmUlW8seXWurhME7vlIAdhglpNT7q2S7O2D3TtS
19Tgl5p6enk0xWzn/AwXW31NE/tpyhlDH4EJEdxDVc17YgJtEq2AGUL7TZD8whkT
wqsOgXIQ+8Trozf8NCkZpnrcU6HvMUg74CRxhDYPaxxOPVF9TLReIEBtnDkQfJDO
0KRLZKMElgQ9XEtal4JCSRibr0irFMwnkg5GqRPdoRAJEgVSMAuIW4LMXYGPtjYg
1oftRNzDaMws1KNHNR6vzAOvx3rKIQXscaAfrEK5e1gw0JZqonBP9lfa4N3+7wkI
aV22MSg9efdvew4HO9eRXrcY5iFbVY8FNL5rdz/8fZ/btLsHsVJ8AnkR/gwWaLhU
UpE/WMtySnBduYwbvRW+81rhbNcEDkbzflZia2uE5rpH+ODMgPauCOfSyKPD0rBO
2qdeRj0pFxxGX1TGJmOEFwbCH6KG0twhk+slbzGbF4jwrrpnNlwMBZWYneCiqMYp
YyGLtEwqLJ3lY5LSYANg8oJt2eYHt2MwFGvoREMT6ESA+rut/e68N83hUf3asY3b
fwl6kHbGiaAg9fUVeFDk7IT/jsn3ErMoVB73AqUHT15HJ/L3AQ18VdXrGV3/49op
OMeuq9YUNIltitnN/dUUbr4CvYg29M0q0a+67JOHcuG4tXq/ypwDgUR6rvI3JfzV
Z71FnEejdRaqomC4B9i1S9u8a+Iaxu/0qVSYetTigGgeuh8/1uF5fPWOfewU9D+e
zqPcoxZKB265xxR+AhyzoqtqMRsShqVbc6M1pCpxqvcTpbCNEo/dRcHBiLXZiocB
4MQeQW96AfOvlxDezmafW6wOQMk6fIInsK/0XBO281YDLX3mdD3T6Umw6Oj9vuOA
hN3hyOhjZkkd6Mylq7Mo2VzhbtE6TtN6SUZqk8z2fced6ZQ/k6/eblzh9AIXKj/J
nmWDAioD+CznFdEA0HdUh5oHo/5IOb8M32U/sKWoJ1hU0CRtbCPImvSx8LDZzDaJ
2sPqzRJFRyE9BbUY6UFVT94UV4o1DomKefaNXezK712ULB4IHOmkZtGsZH4TeGlb
k2ShPYElulG4kai3758YTLBSg3Hc3kTT8mOxfTmCcPiJqsHBcsNcItNfAinx6n7e
8xAKbSnQoNBsmrLb5xkmZgllgPCz7eXoUYICRT6cwT6CWhZyyY5d9nud6YsoWC1E
QvuMLOb1gtiJyi9j1e1eOWjn54k2TumPR7urElsyYKxyKbG/mTXajs665UWBBPAy
rz9G17BN3EnXVy0Lisnm35s8G8qREHk/1oeX9J+gRHs0kLSWCOzZWIeuglJ8bdmL
Y1iwlHbELRTNx8wuxs4UDzZOOKioox0MaVVfjje+vE7rV1Qr+6N/7x0Vh2bCJ2o9
/ZG3sX9+evRT+hpXFRgcQmsGRuQRiTXAl5zQ1Sa2X44NH7si7dqp3oaV0zmmlEZp
zqonauRm0VBXHfKXzMQjd/we+YT/BEoOSivHba3kTbfia41qAlQX3+MnXbfnM8OS
yQ+KzCz+D506JlydNtH28h/fXzCHItAqXqZ/EIC2CdHoSK4S4AJn7yJvy6kfSYUa
ySTZUW78lR8Xke7HGS5n6tYbBOAehnFW04/PP60nJ2zcfC9Y3365ciH7BSshgzYO
vmFWA4FNvq2+k7p2SgybpWZeLIMWretxvmAUcb0yHLJZFKKEpGa4e2lbkBeOgYhD
Y1IIfiib1gLk62zrtjv2w66EGfouB+EE+aScAuZQOg/Nyq0/VLbGE4fJa3u+9AF7
tvw0irNJ1FnOSaAJIi5Q+H8ONgWCAxuO29VyIypXUgv2wfL6WU+/wcAG/rP33cPM
Mez4UcQdki56z5gPOYGUD5FqKoaCr/hXzswcQgsgmnlcAlcbHQK2UwtKNrd+bAEM
L7Lj24n+rMT3bzuRailZjVmOsJKUUPlvh7pwQpE+XqR5dc4UwMzdsEoNq1ogmQlY
iDr++ez3NtnL3HGOpdzb+KIa0HujQQ6pwvFlWtCTmpAwSSmaqsWuTF7o/99q3w6V
52rspMVvOBvLM94N+wn7btHmPlhWUzE2o72hnEe9xPu98+ZLPTA0g34wEVbithUd
j0Fg5ZyQgJb5qMT3oVox1zgglPDSAppYCqAWO+0YD+Pj9oXzLnteoHDd1LbPsXCk
qEZgHJuim7F2wh3eSMuyeWns+OZ0BklkVhE8gVeB5i5WfobYDI5371Rz9LmF0KoU
KHq02HVP/LAQcFm2VV0dLcnzMyObWCOx2d7ufPVtEdVWPBvKLNbVmnaZJPqDnPv5
8Jcd7BlDG+rH80zv2Q2Y0rvEl1qHiFfgZBRC3duPYphlvT3STNj2PLL5rOPmJ+cd
bs4zI/fbcyG6LPQ5OwBvGZ0CRtKKTQygx0nxOgXrzDpTmK7q5oSXdgtEOR41Oj4K
BRpG0uzTV7lfso+SXJ+NGC6WcXhfN0/nKuFs1976ZBbb5gpvb3FLa9Fs9SKVl3X+
GL4ECeKrDcquArhgAQ4X0FHAAkhnjeUpv0zgEqjLCN2Qu3Ad1OBX+bVhaGXGjl5/
Eys2jxcvXLRQHsEoCSF09HcTENfL46Wp+qrlx1I7iVVzwhP535i2TCns0qA7uaX/
kWX/oDr4p9EHhoMZx0VQK9Ajqo2+yckbBhZAj8KE7YfXO9GN8W8LJAZj4DmlTqVc
MtTsn4q4wbTfuuw+ERMmZXydgz7rBmPy4u+gYuD7RJptykeLFxeyRGo09aoH9NB4
CUiapBQAxW00BbTa2terImlEqaJpug1rjqOvl6GgAq7J2rJsVAOq5TbvH7jJkwUN
rc/J19vUfi1I7qqUzkiOMXBIHLt4lfC1MBZh1JevILUab+/XmJ8XeJCgFLpNiuFR
mjfoAnWUDsov8P69nV09VQZmIjM3hry0f/LMusXyOMqAGC9HELFWDAVuC848J6um
eMUqxtyqhLGHO30IfRWWmYhQIrGZBPGgzb+iGtSiSmXCqs5bI2YEiprjd/12PSAU
jP5X2yEB0Qat8JS/iqtDvKgx+vn+4kuc0fTzB9nzp5hVDzZgZwgF/aY5KWofsbCs
uMsyPNXtIHphWcNDDYpWgdSyRMp7TLiq/RMQgu0NpDvEPcS86E5JidovbQtwKee/
/jX3JD3a+KH7TZGnEvxvbrAfEicLO9bDvVhv0ejCF0yr5ZoKQdfkCJQTV0NOw5Lo
lXH4Jq7r+baTBaYJmd0KP/0worYdnQR1XftgBHZOJYjoWthF4uOzKwRcyFO+snFu
6QB0S6VP67Yo5YkDtpv4FChqL+1JxcssOcK1j5BGieTK+QYx+PTar7zkakfoZ/Mn
K5PGw/4NwZZwqu53MpHaqdeA+0IJUt0uXa6K638x0bVq/HiXhOPt8uvwaPRYvbKF
GKOUHyY5A4R767t7eRdwmPSAHf6jfJxEr4nXlaGALbpH99MM9KQ7a0VNjer33P8h
4V0kGwrH9d5TDwZd2XZB8Qz+6ZXgulzRCXTFjhFvwG5WnPcVdx6P68X6d+emNd2z
2s3V58xOT4EdfeIZXfyNzs9YFUZgsD35BIVrDk8+n1bUOX9+C3IOeXMNQ6mEeMn9
L7wxZgfF6kzvxMo5D+xc2+PNY8UJ7vU7dgFN1KG6s8PdTLswDGSzPTTVbHBVE6Nw
NnZoEEVkvPzFg1FHhkmItM1tywBJ4F2XxQlbZkH894glE6iswR1ZesFScxOEJoc+
3LZtuz149jMSPXlc2RHXnl6GOmZ64r4tW6/b2TJEA31+OAJyhQU4TImbmkip4m7I
WrPXeoF9dCMvADwjQGblIVWajP7GmFxu5+UXDhfwmTUkCdMKdkCq17pWYMqbV5Y5
AYO+oIWnuZzudC7lbOisfE2wFnAKvEe36cN6w2Kd08GxSD1+t1XJZXb23kLyHFyX
vqSOAxAyColpbT5DQqHafzlFpSiWLkBtZmVgtBE+9a9H1jh4IVjtojLvEZPq9kED
OW2gx8UGWP1x7eYz+qCioVC47wrut/ABkxuuDQ+QFUWvlTeTi4kA2EPp0Y67G9Gi
1JIUThnA4cjK90hiQcNXSlOs0CU/EK1jFAsHCi6JFRn4mQRJQJhj18Nu7S+nS/fW
Z0xocdCyA+bUTXRn4pFLBsZtBEvuhv+gbTiFCMaUyyx06pinNf1QdfhWgqRH7GDG
knKfPYhj2zB4dnaRQ+c96oMySeZR6JkXjqC1PG8orp0SxKmtzdvNDhHQMBDU+khp
GyNml7uAYkSgibz/sEY+VsNkBZZJljP/U6/jCaOe/TudCXLw5aajIsR2NzlSYJ3+
M0odkQyk0ddCrCMRMjpt0cCrsp7oJR1hcsVUaklroDy6xGjRwv8xDhuSy7LHPqF5
ZgQleU9RcXoH10+14m+uoPEEkx/8fgoCOFbZwUCZ3L/Spcy/B9/+vbp/fsIk7xwi
mthVbUo4N2kwkesuijL6IWg+DrR/TdbVYG2VqmaG0auI3GWjA2ubGmEmoZTFNb8N
NrKqpydhUUyHCz7e8iskFpxO8oTxZxLRR31G+iCBd1gynftmBbP1TqfpGQtUFNzw
cN9/oUfYhOnvp/s8nTniyq1mSOl47A3z8c7l5VVWdMZNVkF/exrAvW5gDAV638m6
ZESF0pbWvRSXOY4wx5tVtm1NAUOwOrbsMam/mSFi7pmLTlAKKcttqHhGtQfYf2Sy
+AnCa8HOw9q1fecPCezrS7SqeEIXPXja4AT6B4q5xGzrFy3FygGWB8hWEMaiJjbx
nB2t0J02ks4iKBZjx63Zn/mWyumzpMgjwWkLL5PL8CsDY1kcF/f3ZEaLwPTua6//
BXRXy1jluaAzRWlE9X77297RvC7dLem6gN196P+xFnCMjmswRqElgAw3PmdwDy9R
TNrNHrUqkNfloGboNCqg0qXn2FoAICbHaSZc2DJIHw+UREJIkzjMoy2OX3jqxllh
RylVrJ99eKrWZ+YURtxXH4RdseagzYoztNhqgycQ+DhUpnbU+HxQsRommJA8vymt
t3pg6eq99O21PoWosn02EaLD3jKrIHSDHkDl01AOPOA4tspS1sg9GowDRXI1VRfB
yZtGVo2dcby8HRfUY707AebVp0qBuwnBqF1nEOe8a4aDoYDqanhdl/BaZbIwWiTr
lWooCovO+iFW9Va/oeOD5T5m/xE742sumiaDZXSrgim2VH5QiBGeFsMTobPMVsFn
ndzo50Ea98LsamSiQQ+XULEJ/PH0HhqoQiaI/26XkU/FCbzegVI+IbpyD7qhZYk9
8LPC5OMcIktlJHcFhmySyI+tps29Pyq5acYnAedgz59gVlGGBYgbYAhZAmwurqKN
Qu8AUTGJJd4CVLPJr/Y1g/85XKwqJWdm0xML1ckitXb8lYH4Vna87Ve+dXJXc3f+
k22+vmuHKUJj4r85TzMbJezSXwNMzVGhJDd4/V7+dXwqRp72ZJRAmwBZn6AdOWGg
LM0JMDFsmXdFRiB3ItNuGiUihyft630ULxRcE6gk9eOcgXvNWKiFZnZKNLuer95M
FCc51uv2mzgVdj1SJTr4JUtSkREnKro9RbY5ZVhuGC/yglp86rGdzcavnMuVAhNQ
1UXs2zRalkUURVgR5ciFxirM+h1J3a2QG7gm3eLzJ/sq+XkAFvVEKRrtwiHy8hfQ
vxKsRROI93Iwsa96CAqu3Bm+djwamsw3CWnDETk9rywN3NwSBq1S+KOm5/33BdTW
nH/WlUdtBztREqaKzZdFhJylipwKbDnSe+nr+54amD66FE8l8oGbcg9JTQtEQBaC
qi2DpyNfXI4RnzqmBtYxOlYKQ69e+EmCqhE4yDVs5OEbbYQpxnuh7A839ZHfe6nW
zya/7/q3z9h3FgblIoVvOsAmTbEZOlJIDutJa4qub9yOgM2EsCPcYwE+lccY3ng7
sLMpUBAZV5Jr/KeC2CAkDX+v4fW+IZQM8RnKgyV3H5RGdwANDar/pTnSX9hgyJJB
A6O9ZkU4KTm73ENih2M3ND0FoaFvjhTSb7GEwE3Mk3p2KoYxAazFBzWhC/31rFfY
Pj5D2kLoleoVL6YQbE7rXlqpx/b00mAwwmbmzUM9IF0KwYteVVGyOhxueKk+ZczF
3ZBlo2aRfZeVVFbqXvlA7vnp4pOZ/1r7LlZC+MwiTeeL6BaMWruUccmzBNfUOVjl
cWS/XJs/WR/nE3Ois3m0091b5bxcHnO0obXtostn+QGjPMPZg5guOndnoRpqKEK5
4VVwXZKd4lIHqqT8tRpHy1gre7ubnjgLyVkaWYkv9jYhBU9zpahZX0HkCZeYlsYU
w6wABEIG15BLJXMPjOSJXIrmFvZwmPKFAHerLHYa/SSNuEHUzjmiEVrFrVhiREvu
DrBjflFlpP6OQuY4doB7EkYeskOZYlsi2x1K4NPDbOLupRlmF6IDjaUB3aOeP4uz
cHWd8QPx3Oir32BF+Xq/rFvc0h+tOPZwBVJhrZdKJ1mNc7N2PNAQ+fBjiEDYYb/E
hsta3xJ1BK1B4rOK/JAVIvxln5s8A8vexaeacM6yHDvF8qnnI8FTjpmia653JWd0
DDFglZu76R8bL7ZHIpwZeKaVboUUs0/6oD1UcKku8H/UoG4p0IylmxGaXpCLg4sW
O/hwdD+n5Thprtl/Jx/PN8rGsxgr0OtuJyQVYbHQmPRB4k6/VYfCK3u6iF6sWrmd
Os1cEhwQBVcsTNBgdhA1H2Kol0+YK3TxHVHTTbymjJqsjvvhAHzJzVaZeeVH3PwA
vANIH2o7Max0utDPS2xc97NdY36zjzyy4Hh4IE+1SuvJYxrB2KldBXwpmRNhRCq5
3M4UTcJpXRhVUzs25veY1ZE4cwCcYzFECOV4v1Q8vmkC4BMpM4LI2rZuxk8GSY8T
NBb8qrsfuLylzXVDE56WocPQ0cMxDrKPmdKUI91KbQ5tbWFOMin0u1YmulzzKOJf
mqW+W0chIZPJfTdCNSkmIC346QbcnNv4MZr1SsS2OemssBsjDi7Gtc+j0RseHz/X
Dn/xzI0074uXw+/BLMdvxKjtESaFeZOeGiO3RJMMvvpLYDN9jxhkWmhY5kypR5nK
7kxxTHk1B0KLPKQoVrk8SvsDyWj7HojIlkGqvc8rTCfG+PrgTQlK/i7k0JwqFrOY
tO8HcissVFfLybh17rlYPUmMxHq4/OKza7NeXg0cPDnhxQUfrMAwerrWleFisQhH
BxohCZkZeZPg2RZmiAjvzDkFCmM11pkZY/2/LDc8nGiBUuuWc0EljqZA7NI0iy40
2qOg3ljB8mWbcCHOq8HaD3GSd2qOIW+y63BAp3HAjMDM9F2g31t08BynFU8X1jXD
zivwTs9nly82FV+scXBnitL8wDpwhPP5Pu88PGreZDyR1JD677nvn+JC1BJaZCW4
Q7cMqpnudAqredscSgV9lqNTm+iPLK79yrZ939Z9tnwm98178TJabr1lS1IZIb9+
0Pu/vi0tfxi+OpQqVEfexA7eScchOSzYZUvUKKht2ho5DS1bOaHPYW2PdzkzeeNr
q7E/fyIBjO522vmC8qhwRS83VayrUEcSvOxnMy5hdHduTXsrE0NK6tfGcjumIOOB
55B0pT5Wfn1lYzjTcVshWwq2/yMyEUmSkri2h8NzEj9CZmRT0zeAtK6to9oj96Mq
8xKvkLHD1AZO9YhTP71BsBC5wU3ZqEoi8nOVKNw2xq4C80Y+aB2VmvRkkI3Shqnj
/woPfdl1NJmz4rULkBNiphX0Ebas3yfSnj0UlnptJKtKD+CO/xf/ZwHymoCLhnME
kHKiiupR+P5B1atnxKlg2KrZFUQ/5qHEWdIqW1Bq+4qKW23z1W17In1Tx74O7RF/
O3IKcr9aRbWiih/0ixD88f86A4ybx5x0EWItLplbPV0X1aM0NX5XzFws/1ZkAPKN
2RjUxeSMLnF3xrKrFPztprXPM6pDQDYmgZNc1+KEmltGVQSgzgnwZdvKFSfaj7+Y
GJTZxycpH+g27yTL9D2M5kzQw75FzgXvzpaB0ZjTGHUmPuc9Ajlxc1zxkbmIM+w1
KDbiUvVSluVX4kEvGxHBSDF2DB1sn1BtR39ad0MhmKAYttRz125xVXFi2su7UAKi
JNCMB2qk/+sARKrTyT4XVt3ZzG3H63YK/YGSfsswepKK6sG4NML4Vfb8SwoQzTES
rruUpLcZmwfJkHKIRhl8iLE90NWvvnKTvD4uWXEVPtK9OpsF6y/tHpmcjtwkV2th
HZNeN5Pr8A7d9+lYqmwy9BYvzBtaYxLPJSzKnLXAWIspDQBOkG0Bwm6NCBPt6+IW
eeWEU5a6AHZneJTOmhl2jdW7eVhuwXWlCLXC5HPculypH3pd5UqSZrOU1mZ7Mj6o
9hUTZ3euHHxUqrIpJZbP9h0Jp4Rd41HgXUFg9aZJQno+3/m/KjC+Mgejc6ew49t1
lJdisBwOpnP441cF2VXW39v1SgK26NnoomNDXQUwNAQ4cOq6g048jjQipfYZNFnn
f1eHnhwgjK84yotyWWjGKIVd5MYiZF61wbdyppvHRRJn5g4ekRaZILXpg9JXD2UA
lSkWJpQ25SNWJgZZFm44t19ha4zuVN4JD6ce+fBD17VcBVp+HRPGtq92F86jI8nz
1ISSI++CP02EN6k4AngFM5HG+IabuPR7ST07/zfuv6KNLsXRew8m3AGzuqbLIQ1x
TnC8VQQp8EY6ljlmIFTBBBYo8irl2SFnV7LAf3mwbpFrT7dHqDMtfP9M8gM+ceFD
LLfDviAkggPCmoAusPLiAJgITY8PZ+spmhuGXEoAg8WMTV1hxNi8lxnlmwJblIJh
KsIK9puDqKBegzCeFQXkZh5NPPqZJclrzuaJeQ01bfsdid6YnQ7d54Na0S0t9HNU
ND928fxWep1FM9Jkt61MBtnPdvWmFZYPsjQH4FHR1ocUNACHKA3bgnr7SbQqH2L8
MJphn0oqEMmzxvrgRbrDadHQcu1Frh5cEtsKY5pE4ryIv1te+AUpn4OWMdyZwrJH
eZE2KOiaNc65EWMcU+aSIMvHxj46DCYfBBLHY5l5aiaWxKmaRZ0HXQjHjVhQMTxh
aNNQ8Rxo4ym9H+7VpGVqzlTwQegTd/SqxhO3zgWyKRfxjVavqeH8zZ2x96btNIDF
zbBBBD+YCiZKZAO+bR/dd7Pip7zPN2G+WS84lfvTbHKL4lhISH4DR2TN562fFG0l
IGZ11JpCZpsKXWyxcbhwCVGsg20iGulDkAvhvuFY8sIPfHb80JFziq9nIOjHyvFA
VPAwyNJ4PoZoTrEFcIoknIEu02oAWIRJy67UI2hOaNH5kLwbRw5APYHgFfmeK3rX
FLFxmbY4auJlfh9rGj7RPzpI0PP6Wig7oJkPkFmxb2fLWmcEzZODZ91249wa/13L
6pLAdVRUa4C9kFSPxjYn0GkGUYFnaKS9VIYaASEZOkYa9S3H3KPywvsTUyf5Ebox
tZZ8+2hxYJtCGovqR2UGd1DarV2bU3VNO4edpOgziVbXlXyOEcqMdOSor4yGgTZH
2mc+WgZwVPakKUFx9N5TiaVwpovDdkeOkSq9LZf4lqMUbUgcjtLaDmEHMyRFUiOA
MZEVgXDwk+viFTwOpx7G3y0EtsQLpXOV1m3DcN+sZaV70wIdzpmABzkWpu6w97O7
l+VDNyPYKRSoI3fByLqQPnFgakzynG/phldh7Jlp1jZCw9+zJFM6TBcrFN65R8G9
gcdnyFmqOuFBnjMpnMXqQKML6nKKCDw911fE35yysyiEQU+FWLae8l9rZZgfnp2i
h6NQO8u7ckYsOzYPHC1wpLBPJuH22RerNOoU1xG6EIBUtFrlMuBJr1uAcJp7XaXw
N3W6stwVTw4sAOpSzkW0yn/5WclTzJO/km/wl4/yRVPTVjNNeTKGPauvfaeOZGbs
PeY6lYbzHU1REtnaQ1e3f4q0hcwN472HkUMC0iIyofgbeCIfUIQ3ATc49U/iCJ1v
c9zUIRrSuxnBQIE6IA15ekcjw/a6s5UNMS+RKimo4x66BwvYKyZxHi0BqY+fRY7F
Ymljv8oIsCTWTOTOAfb96j3Av3rRjoqwR1L5KPGO+1EhijjSru3nwkZNlnp5P9aL
J4Hnj04p6lQWx3+Q7v3n9+x7fxfq2Dfc1HL6VJo9Sl1BF9IjzWwq9kdn5UTCPiCA
OMixWQ8c8h6vHJf18IJYEPdJmil7PYN1H+4ZNqihaHK7LTF/jlwHln+SQ+ZwpSo0
KTSgkD34wgd490area94VUFlkAj1BygRwE+V4aaVjsCN2P9ZtyjmcLYDSO3R7DBv
y+Zdo6OCJiBNOpSHr2hXIIs1heb/lLYTl0pGVI+y1LXJb+Iwc6B10glc/wMV1OWG
gQ8PbZSs2IBCxzlF03PDPzNIk8BzhDS7xbsOxeRu9kck3glSEZ5VdsjgX60a9Zva
Q7YMybrZktFWF43Kk7wr0KtgOlmhyJD5jVAxx9at5BauZ7h5Q+l6iiT97MANCspu
pYBXlhCnhzC1KBbE+C5YOEigIZYd2N0Yqktwc6N2mCMdrdGSx6vstYDxSiS0RDaA
OUvlmyPnGvzGTkfsopw4WsO8R5MMADnWggTf1j8ZobMWf4tQzWxK3+tH7DqFTwic
lvY/mjArY8oMLpd3a9kzxy4ofTDRoJJRw7f15REIEArX2akilE1hvmWYmGx4NutS
cOTaDPDTDY1xQT05661jl1pdNUnGuktBu5t+CGoPk9kIXJrion7RySDg47W57C+q
hDJiB5+NBP5QDpha0s1PYw5ftIS1aH9RxJZq6lIXsVMktNxM1QFk+yDNnLshxH1X
1Dq/NxehEg6OugWzoLpaNjmNKfWVrFbSAyupoKaGzVHG9c2vSzZ0ry+ES3b/jrEV
oG3eRyzXldKCB57Y63QGwnOCxzXnDDK+K2+Q6JJjoO+FvER+pTxmrPnFvWFSJ6ia
mx2PinKuvd94hsb7AYWhobOJeOztaMAukaB3oehm8EDB1UHOpUUqUPWpJbBhuSFM
gImPnDV5XQPJy3KKQDrYi9wwg1KguczTsOpE/ONEdaXPh0dGYqhbQoc4qtyFBEPh
yiD0LPqKUm0VilcYmfGEDBZdGrBOidzRiuQfCGMU7M9yAeoVziTp0HuG1LFMv3o6
QO7siU218Cur+LjMiIdvF9j99gcoTGmlWLas/rSK0hSg8v7MCyH/9tzb04/dLgiI
efl7cdG5xLtZH6gWvu5oZ+zC8DZdY/K1WZZSjsO3iPyfqPTnsZxnqyn4NTceI8zx
AHi6joEei5z9hkFCqkGJgUXjG70DU4FdyowkyQHEYJKe5QEC1pRaqxvmudBWg3l1
jQ4z5o5Cbf6mojI9NcVJmK4S+VMuBEcxNWTeMcWbKxhWbKa+WKeM/M4tgG0FLpyH
y6R7o4ojlKl4oEbYA7shwrxJXGfSj1MzhUtIRYHhG0w4VHpUImHR2pVsmnV6V/mY
F4xqJIYXpqRFFK0vv5n7WXf97CodyPsG2JBv6BFKaIQtsbGdwwK1XVG422Ax7lDm
5/CdThKD3/mIVnz00BTDk3xf/7tCeXy58Y8xC+aRnIRy+czXoCw/u/V7akizs0EF
dyj2yUA6ziKTC/y4F9ufpmUUBPhyCyZuFFW2/P/xIxD6lGmhY2a2q2GbO0V/3sLJ
wIp45rApAJfR7BFfldYB9K5m5HsivRg8PBNHKKL5YEKqs9uRauZwm1QSeEMrhnH6
uKKxBhWm/Ul5UPItRsfu94koQiSf4x+2iv2+QEy/DBqEk2AhNnPh4p6LsO0G6uVs
PEz+hmNKhBkMovIQMrghCcqgcB6D1vnWxlTHDdBEXuWfyVucaz2ykUG/+a0ym+U0
zdaSszL6NrWRSsJsM5+3K32EuI7I2h37Q3T4n7u4Z5k6QRLAhhjb4rdGckenNomh
/vymbCLT0HhSeT03HlZ82dQZ73eFoVNFqqP6xhfXK1JSa06GtMrmKjPWrnY45OEA
GN3lGRNL4k2DWlwV8y+DDhE6ttPG5zq2Atkwl4zo5fZPHrIL2z97rYtNSDCAyvWn
mEedBxyKC7DRMYIUPQuKOrv6qqbypBP47gUA1aSiyUgoAr9vrDKACnPZEuTGxqG3
K/LvH9nSBewHkDsEF73gVCWXrpZcezGhLkN22xzwjD6LPY+IYIZtDoezkXWzbY1k
xKFNgQhEPoEHTbUdM2zOg81ADJg7wZLzCnKD2o4dvkHrDweBk4TEGFcVgRoOntoa
MelZG7Qym00C724FXYLge1mF9MRYNwzcImaU1mtdZTdWzUZwGx50yp1sXHgr1Kfm
6zjLDMWncP2UqrScsWJ0DtjnZ6+anGXtwCupA98+TMN3/RmGLuLzST0vuJtRQkuI
eq49xFR4nCzw4cxxgNyNu7Qku150GBEde7bTkdKLAgRsQ8Y1UTUvHjhYT14aBSgz
UO7yT6EWxIhcJxMbHr6CrLDNYZs9fiYJNPV45AG5PF2Vk1qukpGSr2dfFXDLF5+k
reSOvPFeJDWAeDaOPbSRObP/bH+SC90U4U3xRaFfwc7rQxkMvm5fO6OTh9R0aZza
qPlth032x06GGG8rb5JdPHqhcwHIIdBscZN+Jl4x4VRCtc2nrMynb4SUXTl2YhPN
wn0agbQCNKZJcvNM+zZ7pc0moTd89PyoSVGX18wSPP2p1POQQ/A95ZUQOY6vg+Yr
hvesbrHHgJjM598h8u7SdLY1TUa3D30WTnCS/dyjNrFBjEomQ9VvKbA+ZoFQ5LSf
fBr/C/bCY9i1FOcW+GkOZHb4VaCwkyonl2U0lC/6eTOzxIUp2pdWD2BJGghyVvgc
R7c2anQxvAh2zhmcdHpi+kUtD+Tq310CUbJVwRMbVOFVkglDo78ZHDCvAWaMJGFY
H13FGnK5ZNsX7Gp4hSu+uaEnJPeLFBw2qNVK023dUijSZYC8h7lhgk9g0TiQJieA
3jdMos83iXTV1p8cQT9/LrEJjpx5zxkddR8f+zsKIg8mPfb6XX0JuM6fum3orNnE
YEo1S3w3jD6ycQ3ppYNxmVvSPHNmMudUZbxd6nQzC+ZX/tmIzOV5VyBKmZsZhwLF
gIrJ8rdPzknQm9hpMlUZmjGDkA9OU/yk3eJIqEL8YG3l9FbcaLv7q+2hVe76YxeT
sLswmLJ4Xvbp8Xo7OIDdXitglqCw3QYiL7VJeXU1Dda4+ixnq6JKxNDYmcdTjcB1
fkvutDc5DdGkxJqQziuf1FuRQibA9lwakxdN8nwpyhaGatq3WrEMan76vMk/+awC
1TOvDG8Eh3ZgVsSphn4ZooPa2WQBc/RWvWqxwtRfHFeo2x1EKd4fIkaDDocS5s+S
hD+IwCOVxDI1DF0u9qvaN6absRVdy0XvzHXeRbmwIVuG+s1UDq4ZsrzZa0sSeh6t
MIcaUfileGJwxfMZnSh5GCEEeJ1sCwXaQ9eSo92t3IlUxOWYf5sryL1AxmW+0Gwi
sVdvta5cHIhvXnACnB7w0MtpLogkJ8C0Tl0n5RJf1+VAcs4WlQHSVxpyeVNvijcI
3eQKSFjUgVYGk0O75dDDrKyBro03aP7wVGYauU0LNWSQ76BS6CRdGJlDotz4RDUq
YI5Gaz5ITINBwgCFgoSK/xWVfKNZC5uIZgFfTpto+mM5EVGNN/116FCFeQs+9uZq
jWbfcrVcPHnAVjnuoTffFrnESWKXPsxm5ERuuDS+SrqAQbs4QVdR5CknKlw6ZD6B
SW1JnE2Ae+dxtEhMFGVyTlnFotNtnjuvGm0lcgqpzdkg+Q/RZMx1q+ngxyinT/ab
yzM3wBmiA0a8dZOR4I0NMb0r93tPKlNtSCIn0DjF5fmrf83dnKx/xmal/sDa2wmN
pYoGtPMUhXVIwdUsxWO5Ipq06CaSdgcJ8mOqXIaRdOgwNt8Xa/XZQE+/zbPMnVC3
HS5tyO2wDKCC4MkbLLZeyMSHTD4jiw4WtOMS4whZp0/SGQkCCAnOH0lFP3n2G+Mi
MO10UjpZa7O3FzpFD+DJwms1Z+P7rykTIoYU0lsbGIhUARZqbHuFqMje4QgdNucd
VdCZASC1kLEfsYbEeVSPvg85RsWY2sMLBfppX08B7/b5ZL2R9IBmObsaZR9rhiaw
auZ0eTHz3P5cbV9MvTL01TPgHjETHq9FB/a5J7YCA7LH7qED1vpdSad0OZ3rNeAk
jbcs36zXywVu2H7aVqnWYjSYbAywYIoysqSZNKWYvzM0FkggPRICFNs0cQPyw0Vo
EkluN3hInw/43HE5jMWSdCIcibzR+5CP3v1we0wf8uWwFVdlkXBsAvgP7fre0FR6
T02cNm3o6yod/s7KtUirfuskPzDusonC6QSOvfvQNNWyVVKVjZlSvjpP4Q03ukPZ
zTFoF0/YUSqJ0+Wa0U6giPTEWNsUHOhWcly9LICLjfegHlDHHSaUkBZTzT1gs32C
dhzio33uxVSM3dffGdigTNGi7OOtvHFfOVjCf6kWPMZn+drEMuG5qFtCULSWo/ld
bGBbs+OElHpuzhXXnmXaToUKfNv+VHKOyjcTwEpz7i/LaS+wrDdmXs0nJ1apICCL
AZeABWiLvzwJpnqUxfYLlr1OxWHDBtbLrJ7rc0zniM376Sow7hFV9NXRdNoOeEIv
5jRTWApEoZggEO1FStsM0pBBafmoFMOdBGFUwdjnj4q8Jb1beFL/3wGDTYZPcTnt
gV4TDM7znBT1lTRtLx+KZjiQRcEoe+23kinV8sc7N7bi8Igz0Qtp6pMaTu0gcqGt
XU4mS6zT8r08PH555Duju2H7W9BywlYFzJhz8MVRVur6nLWcUhjHYElYCYmsDnz9
c6v68LuwBnCkwIAPTv6uYqF9SrfCFCpBZ6SpwqOtI71HpPHa89xinFh/lAMgTZR3
f1smHAjrrG8TqWKbdtmJMY7NDucduU9Zlz2qiCESUX9NOaV2E3qqmSOVVd111UhL
BUHA5ZK+5HD7pjH7cg0fbMnyJ7OTxfBLl+L+3EjZYgMYlEl4Kxkxpc37COWMYf82
Qy6U7+tHf+GeTj43dqxy+MNDy+HDSHH6z7iNhEwJylZhoOvv0Zmq3VgiokHXbxK9
FuoqNtpvKX3hK88/dvCXZXwaFNRzJLVTX37AN/UuSsgpeaqthk435yRUfDA6b+mj
Iz4PcXwB0kpYGx9cO+uH/garXpuho1ET1H179WQm3E8Ri+tfnWCIXC/9WG9rWe0d
qaD9/W5XXNcdrVfeuI6bPZfvyddH4SL2mQBsnQaCm0C/Nt36wi/+tx7G1MOahClM
SqpRqQ7E9DOsYzScN6uYhiUdr7m3OZyIpAQ4NyW0SiYffZuzzKFwWiTx452pHlSb
uUiVCq0tlD+WlzSbJn7M+ODxcKH6+XxkXImeKVfA/nlQO5udIZ6Tcq/SkDkyJzxu
0D5a2LtJH9D0FheHz3vcgllJhiEvovwiy8knDw3MkFm2IpT/6wFwJUnJzw5X02dT
darbeCCPgv0XFVkBCQIoxdLD+aUkNdl6G/peHxA9gLqZKYowFajZgPuxpRs8MxzS
aETBMYVeuR5B+WuHKMqlBHqA1/J8UD58cJsori5fzwfLK36xm3Reeoow9vrOW/AO
St2coUB6z73+n/5DZruCNKp/TAM0CZ6YWS7s1HLafJ9xtUKebLt5OBfo1GvnXJ5b
M6VEQlpM6BtszVEVEdkVZ9TgyRpe76yMk9/oT1Yo/NRg4dWnP+cHoku689EeWn+B
ggJRG0+xEq6N2/LFTqHi+foXUzNnSOwB3Dko0Bei5Ny5SSZwXPb6h7KcycLzlwte
qDPwVnZnsir6DdHsBJTiAHtiDDiuByC7d3/aCBfxXZTr8r2uWpwlWG4IhyAGDFU6
cRjo2j+VUsM7S3u05IUdL638S7+c6sqWodFBojgjbGeHkNpm+ik0JqYCUACNFdRq
A+K6inqNQgzlTOT/TOYqGwqb0/PkcXeXPRgqQuwBksz80kaQZUE2B0ty5cd/r4go
piGK3l2o1q5k3ewIrEq1oFyY6Y03Xo16g5ISvxS0NPIaWCZ2rDOxN1HloogpWCh7
OWceo/WhUtlhr1Pa5FUitnCLhaPOYXd49dUIvd7pQiB47MtAttBbc8V9S7g98dfs
NNx9FiYa6MdOpIsiLL2zNYs1xYIxqrvM3PSOe9AvWWWrGCX562CgZ9Sd3Js6u9k1
B3muosoM+SO0/BN5BW1F4mU/g1kLy6B7u4FnKHjtwTmZ9x4MYmalo5EGxvH54Xqp
HeekgMJDKgtQ47nCxo2RVosB82ELiLYnOKc6vuzb9GUthP06EAQx+fd8bkEGJX7Q
orrFNUKufymwW2iYdnTzqFvtbO5Rp4IdClsh3DAbhUwA4HUnAa8/ehsciJ6BBKCA
xZmQEKWNe+0byWHG564WWQBBi6PJlP+eq8NWaZGrJccS+3c2eeFdbjavjqBseMeL
2bzgISAEP01fn0mv8rz0qnEaiknYvalsEYSniXJ28lC30uQDP+DKomJ9Wq4WenRi
fZ0SkjODv+w9tQU54zjZUODgdivL2nV0T+Mhp9Fd6JcVChzzp2Z9gXxviYc/kWX/
URDC2B+jaD0KE6x61/PITBE4BhzVd8rJfiZyb+jW+lfQ86SAstuZsh7bp7FE+lgX
q5H+ktm3IjJhi9d0KdyzxgMkKuXnNZ8jgMHSjJidXYTFBS4z+DVKJJRRpA2/VIlp
DCga8SlqAeCyQM8NeRM/eKDJtarZwu5xtWbVhTbi67S+l3yz4r2Pb37VFr/RsnR8
nBGvSJc/kkuvuzsIZBrpfOL7Sq7r8Vg8rX8E/9B0cILcxEK11a0Cv6JkY+3FR3LR
0rBvCVf6NPq+ndGeOJysytiTO47OZyw3ImQnY7MiEMDQrw9jcQdbaLSyiPbj2017
aHVi8iBwEQnOn1Au4wWTXRioEWNKUV3piw3GBzBOv7eMUwmohufMrx12wghqZKpt
UWS79wxSA78fX74K5crBJRqMkgBMCFagMaT9azkwbgyqGywQgYxdnU6vna4icx9L
jXMQw4wtzyUW1gYCToQgrnb9CJl5fC3xlCsfTDoIaCkKhz4m/wGniY+UgP+/l2TZ
6UVN8SZfeV/R2/EnFIhkDoOKIWHowmzHcQHCV4SAFT70CYJBi4UqtAqQqSKxqRRn
i6miMp5j29l/sbBJ65TDvL8cKLtUJLV2KYaHVXeIyLytN9aLOSsFOTdlx9q53yRP
x8UFwjxhLnLJ1ejgkmJntu8KRlDKKpodWf7XZiuOFEHJx6t5n46QdoAjgoD8MQGq
t8eY9Gu9/0fKeXcbuep7lA7slEiqya59Ck47VBftmKK+p9DiXHcqjSY2YBKZMUxf
vEIs/ECKlMM2BbQ5UuxJqzbRAi6hOLezzKliTi9D9eyWVzqzjtxB11aVFcJ+6OnO
3ZQa/+2KTO6HSPkmWHGs4nLQ0MH67yQBAnQE8JQEY/QrwFg64flT8rZ//28IPkbz
bqyDZoHQY3DVjCdZZ3vlG/FWgvtMDPSmJa2ROiKRmuOqSn0K+mi2L5rZm/IVp9SK
xJpSl2P1PzR3WXfVqXkkPTR/kamx8OH7uX0RJwxDvMydwZyzVTJq0ymM3frUE7qK
e8qURq68SjXuktzeELLWxP/E3A2wjETg+GvXUwPK6Q6NZ6Rgx3SXDbVJ6TgIXamm
35aJKRWUbw6zc6D/uJupBd3PtSOIAaVFNUvhieo9zBfH25pIdH8oakem7WXeiUu2
oegkUSRRHf9eXwXAb5BNZsyRwp5+a5n0iTnDeCnNF2nrkuEjNSbGeCY5kN19wlnd
jO0kqnqv0Hop98cda0SpWAhCrOBVC5ct0sxm/8mTcQwqSfeYjcDEDGZhCOFWYl1d
pJu7p6i8BkeLmdXFii1AmiqkWzx7GvrEsDmvcvVKYFArKYTuiDLsM9aA0d2jolUR
aA9G1sqVkNYQCpPd8/MCvGANpEQIz5pjAoYEZVbavPTndVJ/CJdL5fhuWQSIi5y5
nydRJ0ICh/Qa7/Yx7Z1ONTjkis+L2YAp4J2ZP+QIzm0JZ9ODioclkRlMUbamPDOd
Cm/5V2oVvKK0Jn0WvDVKbH9T3SXWX3+DUgcXemV6u3wQgLET5ne7VwaDrP4RgS85
RZdw2Ulq1QU7Pabpa3rwBJhxhERMN9obfFCMN3gNP4EtAEWidlkqpcnnhVD5XvZ3
TbnJUdglZjm27Xkl9M/EP02kBeUrH5fpz0zPNSuiYhy0e64lNzyJ43sU8Pl0HLN5
NQ6mFGoxgKp2YLqv7y+/mygcmQn3n12gbBfZ60jJHKnGWqVHK7A3CPIgzQD7N0bW
Fi4HEDfbeOIKw7tqzvrcgrTZEzywkHPYYfJH39nKULMgsoXGXm14xz4/c0xPV4Zp
h2W17u0aR7j7QU3G19IoMRqk+GKWFmXYSzd8xZlvzlSyzhY8dwDpwgqSq6bOKZ4n
2rdSpMlfZErplkuF1TBHejR9KG7s9d2csiPokqd+jASItj1e11en+TEb18gzzLzK
1ZK77geh/T20Pkavkt6cmI7nbceZOA9m+zvXCS2wnuGf/bTe6bdfhWrMcAxxzXnC
RLGOl8KG5QC7qCyo+r8jk6zLLjkN54GugVOLYOV4+yqDvOXmMWzIY51j0AZFAtXI
FMSUfHscvweLEUL4DT3OW+6qfCegcmoPbJXCm80Iav9rEzXoCBRv6tgUYsLxD3+S
edNYFQwx0TtaNZUJzR0jfwwN7pbJ3c6XssIfEvQuyYiPmvE/kOOgkeka6BzeKhCT
F7R4RSm1B3FmYUF9y96O7Nc7Ai1gI3Yiz2nQyoILxXBH18jVoRph3shTkOTsEWQr
VhCm+vCLP9gs9sFJWEz6y5cCzUUnDelJFf6fSvPF50OTBQyZPu07pXpmVdZ/uVLD
I/6EJANsmH7Ku+Br58Kt5xIS/V7Iek+myttMvby3ullSEqQbbANsMOSFFwOkneLp
Ck90686wLfg9Z8t4jEKTtNKdi/ggrdcWH1DaSG+d7EWgtmeExxpjIvCBh40eUpOl
Ck74nbWu8Ay/gDCJblIH8e9Ez+j6VQNmFke7yQWqmOfr/BjWylptv17R63hwXtBb
4onbuk6P5OJfld4EDWnknMpwV/Hr3ALk5mBSNvLvqqj19egdS89Vs9+JpiAFErFV
TwGpFXOLxX18/qlm9vpbiKL4kJ+PyZGTM62EqsoGmc9ycLTaURyF6XX/Q9gYbT/x
pfa/MNZQkeSucGjxgXaiQNZ+64Fbi51dO02oV6jVd/omxTwyQeit0ZMxzpoA7E37
tqcsIEAHx5p6IIUB6k6jobeK83mg85iLxwtm6h45EJdbyFWk0EWT3z0AHqeJlhO3
XzrkpP0rWGWitwgJgwEejhxc74fFumh3+rk9gAb4So8MdEqidVaV1AsNCJQ1s88i
x003Ygcb47YB9sYcWfxShn+8b4fpAJHzS9Gqy2fN8WeTaQHKaJ7a8WVtzmDUj9vr
2S/2MuJQIsc8UM2QboNoFHs2ml74iDTjQyUUhJtctpOkzuNMVpc+xqp9UPd0iqOy
u/OvcaYeXRBo1mBenEvWL7Mpdb/FRoJ5GyiuqUQs7ck0S3OFT0iXwDWxhs2m5lfy
Ge/GxplMl11hwPeP93okAvxRprwMyCw6MfJDmV/XnSlKYM9qgQzQ7L7yIUZyhD1D
kTtlAyr7SEGb1IkRyyv/jh5pTjECpWRgwGlmvG/SFXh8ny+JpNIIMDj+h11VJ6kP
vfjoAJVM0e8zzb35hsbHhWcBG6pUh2MJcYw7YT7nPSlcJOJA33XcVrxECp96rwfm
6mYV4//VjtwMofZIVeHHoFPOPfrLY1iS1h1/l5jVVD6bymmlf5q5NsbTbqEBSc+P
i+GaJzZGuDTNd6GKiFpsM3k15VqZnJKgKsKtDWN73cf9vdJ6pIm1soSHwjOZsWwO
iqcgqa/PE4hrWLhPdvjxFfHdsoyhshIDlimAAZ6/+cM1FGBC1dnO7ivL7CjsLc1k
xtgzIpioRNAheHNkIAcp21SY0kY34pUEkpeL8BhBeVVAVpjMhHUcFBMw5FZOdG6/
stL+64QqBRPpFvIbFsMNTtFk3pLY0gye5Mlg5g1oNTHh8mUU/mVSoBFWVM9QkMEV
XMJWc57C9beJPAgaaxn+JthWgxTgyeqt2YgihhjlLjoKPbjX3u3NNqtPfaEqkC1E
NdiVHPCsSkpP5ZVqsXtACZy1nCMDZ/G/2qwEZXNxgpTVAFEMOuFvw7/tD0Hry89A
H03Y5xIXyhkkXGlwQ/basqo3QBEgk+yvz36xzNgrfygktnAniVM4IWLt552h5Ezb
FuUZbKlnV09mDk/jka2pveJjeRfP+CFEndiSb9iiqKZ3DS4yIAY47ykAQyaQb6av
B+cVGDHWnUKb1LKJPICDMIlYO1CW33XCtFLWKtDB21hq9mbXv5kTOufl2K3Gu/tD
qwvwgATWbUYVAfHjanBNM1Qr/KVZqA3HCISGG9DPjV+6SvPylYKRD2ifaOGGqw3A
HlxEV8qvw2W9Dm6fwsnl4jQqWHM/W2ekGECNcOuPb1cX9OpjNJyxy25k//fd1s2F
1hPgLoodF5yuY38ly2VeA40Ow1V+qNgf09JZNTlz0wC0tPmDOIR+eNFXukI3fEPy
Kzedjq1PPq1FztX8rNj4BAEkNXZ8ELfvWiZEjT43saL/mIhKZ+ACGhPomny5geca
baLe87xVYlY3XqxKXP1gRfOCcXOuNOwxbHiFg63yTphK29NUzzNOss8taJxQhy48
KUrMUaim5ai4UN/iVGB+FZazZfDmFJMKy0aQJBnmjRSrFU6GZT1i6ttPWMHr/7Wc
i0R9kGZ5JNb0vxrCwMPO4StC2QD5xxM9doAfrO0tDXZfzfAijzE2khm5iNtnTy2a
1D9/R0X++2L5iXuJlg6MIA6ulRfZiIGiZSThWBqpCnt0YaJJgzATpZLVZt10tmmI
ViUVkf4K/xON5/lgFXZMK6FidFoYP6eThmkMkWqoTt5nl/Fs3ZeTCnBkXmPCZ0iU
mOX7h+aajdO43cj2fcmwlGTtLhLT2MO+XaF+Af5B6oVF92o6ABoZ6IeGygmjAi8b
IvLmEAi0ERWDeDlH8DGdb+p7X3eyBr/tqXUIr20kI9L0ta9aVeHGhp7yI6KwUz9f
uaBBV9ckcH7yW9/hDbtXj71CpW3OpuuXbwYNUjKmuO9SLUWD5KSY2IpvmnbWlnoG
AA1qfK+dyhYOIZ7srpam6Xzxaze+ovfAjmLV330wRt80b8SjH9QFtBhhGdiNYtFG
oAEK8/nIapvdYBQb18w4mJBgXJH89xjoqp/haykTjDMMUgsh5GQndymYXL2HyleO
3nrBhAdXaEfFIa0QyNOgwKz50P6b7zqmf8swsrq5xfK/f3Pc/7EjmEhXK+A/+e6j
ryf8ZnVlG0/KhCHTLShK1dyTUxB50Jb2ImiRB6vj1WTdZ6OEt/8Q3900J6lRfi1v
gUp0RJ1Jwam0vVr9y6NioaAQt4PNXgbg5oBmx7Mx5bKIvxWoSw37lgcJLka6ZPjS
R1InSy040EAxt4o1hgbm0Qv+NXOyaJ6EvnQDCA8hokKdPo/RwZ1CkRmF9cI8SnTe
Hq8Aas+Fyl5skXRX76lW5yqq6k/GbPs+EABw/l0bi2uiBGrijqfGjTtxtU6qA/tq
RvSZcZ1jnNy3y/ns+8jYtjQ7DRaSlxgjo6EUmL8m0GIFjjEpioUBOD0ja76Ac+gY
zyhnhY+gQq6r/4TBta0WjgJZaq1MWTsKPP4o39Pq9Ug+/Ha1d2XhoLlasPmuBe19
aUyP1JXov4s6wFIwvqFZXLb6VOerLaUrfF3pBRx0b1RnEd8VRJzA0LD1SKzIbwDG
SQrF4Fk5xwHvoHz/5Q1a+31cgZLAIyqgpjyOE/G6HJYvFoLxus6PHCpD7yVsGj20
huNNjzDo7gR1jQiBWjKdgR1oflqptb01HxwYZpry30A3KbD2YYDMw0PkTvG0ZZPv
Cl4VVIfS6QU7F0eiuVHxN4t+xnbreP4WcRQuORABBhClJWU3tfhCBT2pK4l5hWoG
cISXU/ILmOMBKj74WMjeBbXomkN/gRwGmecTeSA2GzkS5FA0vhwlAObpsYOv3xfW
HWk+1EzzOhg93iV2bekwBAZECs/Z8cNvJ4zOsICnfwaEQJPWx9IxNfY0IEa6q735
s+V6627TC8glf4Jt0LgNUy6+yc5j1dmvBMYZsH8fwKORFG7ElMZhsFVuPLXGZJWC
gK1+S0dI6IO7HWujC0N9jfQWNbiknr1b6ejxZWX94ecu08yQTzREWfGFmmT1hGn+
63aZt/Yd/D9H59ymCrnRt6LCEGCZLPA7qiu+jnHKCjFk6SdPGPKMgW9mYlNC78E8
r6TLQxB3KTYMDbqoaKTpRhYsastQBJrMK+JRv1C0VjomdWAqJt4Db3xJHIxVkHzo
NAgfv1mMTckPAQa/+D9LyXicIb4eZAsPR2d3sYUzJccF0yApbsLZRq5ztnNaHWGg
E4Q/+afKPGTqJ8HBOAOAb+IxbrMPi61OaCRDLt4fazXkl6IDdFLMmtwM0Yls4CFq
FvAsm18HHNlsrWd/3Gcy9CBpfB9vofl9Mhv57jv0Hokb1k68sHUq210m40tLJeSe
5EfG5JmoeCwEX6xX8Ab6LFE6bRfSHa7BSAGuR6ued2ZXLHeuWNpI6+BAUfIuIlqk
WWaXriBwdgDhKD6mBGySf/LL03WTQB0VoVm8wYEAlGbUZ86MIZKZMRDJEs0au7yG
PnRHGLbEYNKJoAB9DP5hCoAaD8fxefx/6Gh+zY1XjDR7xey9upCXdukYMjAqcSp5
dgAb1YjVWmRIxjW/Vyc5bnUJIpc3y3KDRfrS34r7TpVt+r9RDMghwq9uVVviATO5
oOyZgY1NykUt3M42+5CYBHE75MNUgpqfutJ/1GXLfKPPE+CaOc7Zni1Kwt6Bbsj3
b3x0OO6H9KjOlQj7EKrBrDc5weH7ciDCqFsgYYNuLcdAYtAgC0/5KKih9I9Sih6D
3m/QehyVl6W/12Ka+vdGtAhi4DsQLCyTRciE59rC5hDggFj0nSxcvgz//zxKq00x
2dkB2URs9j3ifKh9IrdG64YP5gm5EYmfJrE3xW6R2IDM8aZs1PEJCpPiEnLlvdGZ
kjr7r4khpEJeL55vQgQQxidOHj5xI3KsUK5m8p9u3nTgpqlAC2O/bCReh7NU4H8V
GLoa6oTnp1dcJs5FJAyBRZpT3AJwCH5beUhbHehWQXL6o8a3nWLpU9zNJLSaG6Hp
QSs/gyJy0NUgEzbFr38SGIFjhlRn1tRngqkeRB6YNMSuaW/VK8eCj+JKpYlRBuF6
fKlUZYZy5PmRDygD+pLxJZjXb4LU1bHTDSAbVSN3xdziFNTXEUenFGzl49eFJu5X
MHW0Y7hTFzHTyfIOtnRDkhBWJDIyyKDVrKk7MJqnOANRHL8B9zzCyQmoKnu7npiB
OOPmlD1bkYS1o+dmz3IF1IC3yYnI2YtEMDmlVgkblCOW1VNicQEqciDGptSZ0cK+
iLSOX35230SxNfZ6I+zAkFcK2SMuHtxfOu+NrkE2BfDV9Dkxg748vFaN+acxZ+nn
cKiyIF08m8bDt+gkFQbmJ8r2d78MUbcMbc4hIc9krb3LMp3gXALWLXkT5V4oxlAs
6zJOXtqM8jT3v5ELGf3OVofcoNWuZ96mMfQKwxTHMT9gKLvOU3Od0csFUmQ0j9NA
ScDLkMUeG3JMGFFTEsUuAr9JO7e2X4w3q+1eHPialurShv7IYleLkPNEYRuBCASZ
sCq9bNpSTJ8ax2w1BYFRpFL2PDwcjOAjTM0wCyO+dHhTA0OLzLo7V0mFyt4uCtx3
VO1SLlONOxyANRGlpqU1hZBMTK4UkDEw5vc24S/g1AteAd41wi68vyUh5adCMv6n
Ks5zZ8q06iS34PJSa+mnq7QlRl4BPmOYtLvoZ3qZeI7ptE/I2ZMwF27Jay+1RWgA
rdaDxcd5QeyW7QN06jXov6+6WggTJyCDVrTxd6HOj3o1FkWYWMtZyYqlSJrqIh3f
fB5p2FOXM12TNm4lpWU4wLIxjr81lADwa8z0dvKsBbLfc8YxodijvRgwLX0OFPKa
r2dJldTh5H4SR9AJCE2N4QSNklAARkGFjSmYkcoXMCVw2g37d+9F3VOEloLhBA50
i2+XTrKY6UMyMyblpkqJntvNXzgy1nJ7wYVawyBKsR9LqrHkKt8hK3iAuCgo7oc7
4UCkRohyV7VsP9GMIO+KZqG/QoW/R+EZO7P/qzhi1xRORUjW0uWMFv9eCYQBi/nt
D+vNBpVFYhEqbLiHMxzitjrNk35hDS1x3cajKHpBuiDt22M2VuZRnyGU7Ff2ei9i
W7vPQ4V6LChCIo0UVHhNSvonANmisvBvxL24MDLxRkPScQ9rPnWd1a/in49KcKmt
zQhMjesv5sJM5VGce26+StgplHr7x9oODyz0QM1DmidK5XroL9oUyghu0RagcU4k
H3nOg3oLMtcmH6wlUZIZEh21SIvJU/ORtON1snfIoOeB9OGGr9Ec7Pybux9Ni2AU
+6bvoMbhIHOocQULwt2RqgBBEVcgBhbncKjoB2uiJArfbW0o+ZTvx5rubSkPbDCB
mrVPUysN7kwtlnfS5k7GlfL6Uu/3Uh0O+WtKNtwh7wtnE8rN4lsfSBQWcIp7JQjL
CjnWVXwG0aai3qLY5ejauN0USJKSaPq2pLRZC3ygAPK2RbPJito6jEAn25F7/5At
svvc+voUEQi/va4CnFePUMgXbk/sKI9ObKwNvlaVqgzS9wdvpUjIJw3sW0601WOm
HGSLmiatashecu4QqO+KLz+zv2MpYH2URQvPFhNMQ9j00LAr2wqmE0PMBqTYA79b
kLl0lichNroGFvFjTUF7cJTkPqyWZRVbPGvQaYjpFr9T89tfNMKjJkQC1yPM7DNh
bwydvF4wKcX97nQ3S4SaRMdgLJFjpfF8appqaIhMY9WGBRsb5vHea8Xljtcfn0KD
gn2s7qV/c8BSOZHe8T6ATyNJKiYgB9Kgb0916RLxO5GYm+5hNgAi3dKx6tg0Tv7s
kA5qDx0ExtUXeA0bgJHdshDyFCAWFXTvfN50M9+AUf6I7+vXo7MHKY5spg1/k+jA
++/Mvt1XSdxiTWOL1y+zB7N1ID18e85NvygxAy5jAi7VXsp6W8Yaegv7BNUQflai
fBBfHP9vNlJ/Q9IGy6qGbs/t22ZKgQ3CaTdJiBZO7LudNAUZ54BMV6/YtZjsKQMQ
XeMSBQAw9A2bdkdKNp7x7ySv9SV31N+t6p2UrbuK+2sFtbjJ1OrT2QwnlQhEFUIX
0gf0oJsyMdGfZsUg90ORmtXOoi6aPR6CFQrhXDKnPGCPqIjfpy8l0FQuxd7HxIp1
30JWHJUNwHWkyMRtEMt6mDipuw4JZaL1sFW2G0cZ2SVmyckJJb7XgYJvEZ3kzb7N
dBLjd/ioRRvoOeBF+elzhz7NOqkHZhj1f2OmArn9Ewbya8ymhwUTk3/3MaVPl+fA
2DTuxY29tRi9nIFAHrWboFkg5zTJS/RAcwxRkY4g92GgrUQHl+QIDrttdctRC8aX
p1ghQeisJ9eR4lyeGk5PttvaQvrA1Gt44wSjlqc0GXfeTeY2YRW0d5ixFOCaA6Y4
FhCSmpXWERpmUfEzN1Q1EvOtJPLfKD8N6ZEqICjf/d9e14GhFb28qaVRBOWC5Whi
1jo8U+bkT6wwUczheodtJf4rFTdSKxpevSZYQD8EiDVU6GQin7KXmq6KAIoTrmHZ
2vPi+FozEfol12GdZ5I2qdERamPoJsaPq5IXZHGS/3CUnvhaDChk574/NetHlDRN
45YqqZagSlXhqwxQz/RYXjMstvhkRQjzEaItOzxyTtwDuO+QEjiquJZcXEC6bnaL
tKmDQnU39l4EKXRuxnwHn+ZP2A1G36cKlkHd8/DDGZKIWHodkq+0SPwhUScSXKe8
K1hBqnV7WswBvEcTwT1sbnbwdbx2jQeUCI0uL49MgX836UOZbSVxAFCXyjDPS0Kn
AlyKL3KMMhAQ5g4+6vbcqDfYwJJtBIxBuJqzbng7WdIFuuME/i3XyDD9qhizU6Wk
Y+Beo9Y8Lx7xB5Y7O8r9n+429NMbv/U6PnEbUN+cC0rBPyyS7kq6E2+cFRxIfk8Q
p7MNr/A0l/osdWlgE8fJz7HpBBCtWRPkvvi3dP2a7Xv065jYALQQrhSJuGcgevck
koqYsAYEsJ2dW2LlI1Pq4D6/acAD5pU5XUdfwQ16O6FLpfgWOAyy+Q+WtY8E8ts/
jV3orneOLvMcAfYzS0y7xPXdjMy1s+7msTNXAYQF8/wz7ImhFPW33quuCQDAErgf
njbqnaQb2HYS/CEWqhko7qVEATmDAHy4N7cOooeQeGRY7zqd0HdTNPFYPQRa5pvF
Pa4EOn8WEiTRj5JoSnQwwvyTfoELaz3hXg6cHHpIplwevEB341W57AgBpFiK+nKS
tB2FgNbtXRyK1SJ9I/QV0PXOIyARTbAix1Usj3pbbHGFgDVNzIPyUrFEvAn1fL4L
uYk4xMlNXQr6UeMEp18wpB/X78zXKuKtBg81qrCIwuPNWrNIjeVxW/xtc4dkNaF0
swjtNtRcXJHe+5Jrzybos58bcuCEvr3yVZZENrWJh57SI4Hn0k0DlLHU8jmAzl9c
ShZpyoatUNBYgLZXIvHlv28bfu/bVVCo3xtDwFlOTvDVN6svWa6o5S5XyDizOBFj
XeBcnbqZsKRzeetX4fcQWm2b6XGPZMHdO9Eiqqz4sK0VMofvBlXekmwd3jYWU7zM
eCJu0sqxwaHRTxzifIfHtZm6HmKDlXe1cTyWqB2w4QDPAofhjiVHPWKd1fO/y9FU
d6OpLTdIO/czqOF1qCc8L4jT/D/NXIsYT3NlHr/eJuUEFKmrej1bym4VPtof40ug
96oUIZB+4noKAYM1i2uKmtDvDC0RKoeebivSVohGQa47RndLAziFDp22d+UgGFQt
mgzjhPKT5UX3ve3lhUaNLgRA+3Vx4e+bo4Jic77w7hEYk7CfpwZNkN3ZSrkTXH4g
YuF5i+qOCbjqHAZ1SefxdnDCKByl56rynW2syLw2TWHeiGeqWYZ+RAbpo3X91fcr
/K2ibe0JhTz7IKuneljd3C/NlKPQKpjdKUOi/ukQKel697YSx9G166a/e8hR/VHQ
glcxplYtMP2wzEZkm6xWVLl8auChOoF5wOZYgUi+Wgu7fR2dC1f2CQ8lUnSkOUzH
VcYoTufYDnYrlt92E+q9nnAyYmr1ZCIZlXO0ZFRQR5eeNuYgtv4/J7v3VVwK1wNP
202StSQGbsSx2m3DgUrT05yv0tcff2qogL55knkfHh153xmgq/s6dDGWYIcoAgzr
jBrwx9ykJEPDeqD6m49fAwZoc+npUPLbIrK/m1bjStv1CEn9AnpNQ1alut+gsaXj
AC9N1l//NLXDXIL2DV3QVQ0ZVHjfComFI72nbxSISCfbKtnUx6wP8Ik8V1wMtdP4
flYZ7wtmdxuVHCvhr513gAK2eJkG4fYnjvsrNIKDJwAeAjGSbjLEDsggSM9vAbZe
tSgnCRQ7XIGK7D5yg/0IGc6JXVm3bG3/t0E0e/YubG/bJlmiTW0SdNjkc6nGNTQZ
1LnHu2KtMI0WkV5xsj1s+VmxdEKZ3MP4BUtADLO5EtbdOKk8XvuMhedSyEX46jHR
zm6ywg6xgntV2y6TAjOzIBJ/3NYieIuU5waTxSgH6C50O6nFbyXk8cCTWzop04Px
w1ixo+htLe6w9rdfzzqYCFH8TXRyqZJN4KeTbUW1ycSvlkQzkxPr8wHvJg7E6ZSo
GFgJxTQDJcpyiDc+JgT8tngG09IH+WLEf0hy1dMimjo2vjO8p1l3+eJqBJRkI6vW
cS2o0lhnWjRqgsI4AJqYuOZaFx8SuBhoWghNH4MUG9XzrGbxW82z8bi/ICvLvLMg
ZnhQF7iAA3+SnVeebS3nSWsGf4FsfExG5VBbJpKj5T+GG3CJ3Mifl0iHCAalH/lg
B3UTrYxa0pPs4x5aWYQNBH3SBZot/dXgQnADaaoMV2eZ6eRTHixHQWe/x0It6QHh
+G2g5b8UD42JWDFTBavKtPeDoE0Lk7T1TY4ygwq1RDvXbPDGGXh1o2/BUUgbrMIa
1jhF29QOG/C/Th4eAsUH/xAT88PRlxkQo1jzwFnvepjo22pRlgtKIiTw8c98BfiG
TTwITJaNfXMOpjW9Hqm8z4Na/WtLcm0pr3FVX5+8rVLTz8kZc1pWvKVyHgCYhNgB
9NhcMJ8Hu27c68NQwocKAzfCErzHiWQXxdDh6LGusljj7jqeR/+d6PADJcDhKsQU
ksfwN4MBJh2vd+fHKkWgwRV8Dud6q+FiP1u4i+ssrEiE0RNYJ1dodCltNB7ncPxt
66BglUgg3CvkFykzTaHqbUKoJ1E0MywYf61Q+uMRbD++U5Xn9pSnHd6qhj+nu6Re
LwdeB240mVZftncjjq91LSuD82MBShwEr3mKFwAY5k4/VwRKV+N94AnBug06obiK
W+duJcc07mRrhByQPRe9Cp8iurHt8Wbb4Cq3kBITRO5QuqMqVdh1vLT3orN3FMLZ
4OAVueiGx8da9T8QMXeNWWUUmlXPcss4wMmkNyA8O0ck5MwifqYwNwuLkh+CTMyG
T4nf19dIPFp7p34KdGfzoHM0BTlr0e3lB39TlZ4k+NLqCCdHRf58Szbg+Nz0XSo7
nHPGVkZEBpzvMBrnqhqUhcXdHk84wQdl1x/QTcMrI1C/3MCXYrbUVH2fLnKFPqg0
BOB+qFXeIEC+wC73dfJ9kaPwYk8FCVSz30DRMusYjw6nCUAy8wuNw9IK8boEAjKn
cunPNiK/8XDQgbY/sddN6bw1KBqtsKy3K1OzTdnIF0SdsJns8EkzfJoX9Z++GBB6
/5chPwVoLnpvSeBTkMA4dLxF8xCfu4h9SBhxDcg7iIrcX6JzkgLn/9dPvWn8V2Ha
mCleCDeS5vjyumccbFEd8YFkW6w/k5CsUDB+G+IclqBs5XODenUm7mEGNjp4675b
FvhUASbQ68s7sUyVFUWOzTd2lUGhC5fv8h+msKm8SFOGUfyJHAcTMYnCT2m+cG8V
K2a20Z2VXYq3CyHiVrt23Wu1XnBw1Fspc+X0kASKpQQm6Rmgq3U8Ca/u1ys03mA8
rwbbmynFDMIEDPvjKHB1dOeQIpUO82mEuxfLoETfjC6dNaNOrZwP0WeMr4xCMcEZ
CQHArr41NJ27ccUCiSGzZKb6D0wx52aymhT/tVlhU4TebHhxDSh6Gsft012cCM4C
jza+Us6iXxNBNl46DM5eOu9r8Cniq4T9rvRLjOysTFLAOekHN3DnxKj/kNivbZcS
E/dUzO+byZq/3UQe0dMKCnePc85Oq2rN2i66oojTxGv2i2mOW2ZWj2PgCbDS6Hjo
AdUtVFnlD2OjDt97WxFb+vHS7R7k8Jz+uyLHob6cNUHgAqxns5/BMI+G/h/fu3oY
VU5CThvXAFkjVvi8M7Fi/mLJHPzZPicLU+XZU5A0nA0U7WdfXxU/I6FXzZWDD/Kl
e/Z+fNRB1A2AItp5u2BEato3loYBFfa4GQE+ir7vDJaWY87XlQYQ21x0iEDax0u/
SS8H4xUvAZlfUzT1Cn02kAbwDzqCNysys3GjAutzsD2Vhn4lKrJJYwxMH9IoamDb
o2hPvqIuk5UerTrL/o089Okhs+skpQeKNo2M+EaId+qq22DosnIPNGQfRKLrjBoV
YyhrwKzsmKUwhSynkZ3/lnmw9lDqG9O72SRo6g7u9N3AjATg0s5ZKxO4JHy5fsH6
fcoxDNZAIs1qM7OUI1lWBFgoxeuo4rQFzCxV+6y5/Ef00snWjZ0+aRCJLtSXbrbZ
B8GUq02sga9WTLxZVkLzv7PrLGxKceTFP/ef6HTqjoZjJsZqe6PhgOFFlS6EWHSN
JdHyCF7Sflg1PSLc2Heh2So6PAASGt72WpZFBjH2pE2kM2qbCmX7obLw/tYhLOeL
qv8ucJZVmmhjs+l4xGn4/Dj5zuG52iRz6n+xI0X7pii3EdkAKY8xDv8WTeswBFnF
7NX/xUVKwcGMl6aFFYxmY23By38l3lwzluQQxBkPvU7Tuz9yl7geSjHv247m/Yzj
g0Sgn4Xn1DJMsuK3SUPw7I5bTui9hXQFohkJFhGh4P4ggtSFYzd6FYgfMQO6XfHZ
khAuSWiiSt6IcA6cy93Z8x6iMKAG0Us4uWRDB0NsqW1F96AP6JmzVhYnGEqh+KAd
OqJaMrQN+zDumJ4JOV5DDlQMfWFXx3BhuQJdWYn4l2k7Oc1dLVUzFMOtKTk5xy0D
0CDV2i+qt0ehZRikkqEYbKTdcrJgweIvY0bOm3KgKVXAd+rwQ2PEjmhuh3FyCdmB
mWWv0r/LB62ltFfX07kL9uo08L8aXXHf0XjzzL7I9uZ4l6FpFIEBnEdKHTilfE6V
oR0A4NnFb5AWryDBgkDG1NV0Xc700j9F1OWusOXCzWeajLqKe+mwxRNGeigys2ew
Jy8j1JlDarpmPu8d0lxCP13ovkQH8n/gDj1MIX5I2s/oVPd06hxVoWM4CuxiK6+y
4dIExmjxk8zNdtqmrxFhPk0C8yhta7HKxfa0FAWywPnGIF5gxHSRJQMN3sTr6USj
WlvGY+Nd3Tfov4QANWj6Wry6Eyka/pFPEn8RQjRHesPPYO8lYIWmxxGmHxm5ljrb
CHcoffpmmTXwBVVMJgWAmdzczxLr4y8uQ7RWslumMcftpH/Y6MaWTDi+HC4FxMrx
qWGmWQtxtS3q1pcjD4cWLUVYLvWdDraYHVyiZTegvWh/i1JUpZiQAx+vMEkPVNyS
S8J2LOIOxymPBr9JYFLi9ZIoKD1JhcF5zrPoVCdGpx6x9bOF/Si7PIwLyg6e1qAd
YLhrfk3qEE14bwoSt0sBnknMpVvVhICiUHLWSSPUYgB1BYQCpe+oZHJa6r1ItZiQ
dri13ojDFrF8ckYrU7aOcxwal1gxEhlxzQ9zMc2Ah2Yyhl6XV8erCqGF2pHzaeAQ
tOfItVuBaf59sUbKrl01xR/UXvBfOjvAPSmVd8Y3DfcGUkAoDWYq3cwn0hNAjtSD
HVK3T04JXOC79BxoNT9CUENuv0FOv+WWw56TcXlOqhQZmGDppd2sUghEQxRaF9sr
UOMJl9j5O/3ajLDXHDJFd+ttlgAMPdJ43VH59VwVwF+17ax3No0jHdCe2CJGb+wt
ccycjisp6s8KLLktwOXqBI//w/PgEz19twQhHvFwWisaHer9D/WNl4CXCjFZ7aUI
hXMjvxhD4TLDd77wtW9a3AzMYOrJqv2+gVstjTg1mmiG2WPYAZBgeuHRu0SeqziK
9F7QJWaFfIUnkTJB1qKT7PMlXFA75vEYsOGJsajUDCM9t9b2nTwIQxHnyCUCCyQk
dRwrRtEYIWVeLJVKx1T311y+wzDMm+2N4wZQqtE1WoLZnEFvyzWn8IxBUR+HkY+w
gn2pL/rwMku6u70/C8pnnHf4cw4qFAsqDJ1ugKfjp+pt66yn2lFLu6RAfqop29TC
FdERE7DiOF6aiOr8ElOjmYy4m2eoQ6O6mMhb7uwna/HawBIP7tJSaydm+iDgHVev
kni3fEsWf8o3yrVsvwea2K6i4jqOHKJLj8TuQ1ljjNk4pMewVdEnaGN54CtKX6TP
8XPKa/LQz1jdZUQS8SQPdBjH2l1mvymR/fdsafR3YCE1NUR0o8/I+hi9WOU+G9YH
86XmJWMdWOSODDC4GizCr2Vg6QDarQ5pN8JDz4EMcZWYsva7UGCxsRVQ9jZJw8Ya
npeZVHcjbuShJZ8ZdgpwWdJrWiJCL2zrSs24tA8DHycXaROGK5tsEzX1oJfjjDDt
GhEqIW/UNFsGevZ6k3YQq67UwqMVCNjQwdnaBJczho9+FBOE0Z6u+Ejqgl9LiiZe
UD8a1pYJSavKG1hEOWl7TYCNw3X/kP5JSjLon/e2jONvXcJIfTb1CW4kdy8sOOnm
qsu3AxMHIacJAxovgegNdwLLNH61VbX9yxUk714iQaUIrv3NIsq0s/kHgp8TfCdu
gJ+ppPEWZwodefL+cTU0Ek6KOwfSpDo8eNGNDSkqNRX2Bnbq55KYReisrUWu5RSc
i+u++W3jtGYj2a6xiLngoxMwPVsVqCHZgj7/v2XxQNb3LRfU+yni62y4eQZq23oO
bQOhUHiRoB+KuGLQ00AGxsV4+Uxhv7USyKbaZ8lzPCU7KlJ+p5WN9myObYuvtpHE
otO4hAeWAxgJ9zXQBQ90z5ZJXo1n32GM/vR74u5gywd5h4v+vpnxNdYwU8d/hQjh
8MrGSEBkSZSLoVtkU2pMyOVr9rYHkmNYxhepqpbpDmAhllEj65plBjafElw3EeTT
5czwzMcJlWZDYznwgVuBcDMdsYsCoUGvIXFGtutQTWX2j4yYvWpB2flnrQ4Oh63O
T6wWXRZtX1T2n9iE2n6jX5+FpAban/uJ3BTAMl8TFzwSnfhEAjUwPeTjMaWjt5vM
WVC/6nwxOhdGUq8bx2f/tzEUb7BU8imUj8gtvCumBW0XjY6rxqVyS7s76AUL+bW3
Ks6MNuusA7vCgVo4vzF8zACRKtKiQmftAhjGLpW257nM8CmMnCHLP4QGKMcSwozZ
Zx3TLusa5KcPJlFX8BwPb/aTJgoRP8r5uvG2pvvoUKh6xrEUmSkah+oqMjl+DbvC
hrue/tUEdoXlWo/FItN3PPs4XdNaxCIol3mGHuas46XRjhOWVau+9ddb29jceONc
op+/nYmN9tn97Q0AHN47e33gJtRl6LAySA9AfOf7VEZF3SYNFifGUZUeKLs/6j8h
sxTYrWxGmqr33iwMZHfbWoW5d7k+leJbrVq2ezEHUysPgy/o3xdijfpwNTBdKQ+9
VqFJ0BCRBTxUzjERdr6J3y72HtbhhGQfdCIiGHXxDDAgQMd+Cm63DDUhOjK62HkA
TFpa/gQ1143kihyul96QTLbKOErubGiP5xScZpupWAiZbiYNFcqvDWK6NXJtE6rG
heNB4PTXZL9nPmE9r4CjhUj9ygHOu/H6ykFz8TuKXlyU6r09df82JLwQRyp8h098
c5zasPfXCKg3dKPqwcNdg3MMr/4W/m+BqfkC4FLuxXZx88umRQOa2YJkkRkhkoFU
ah2VR0U19n5q/784GSs+VraiNxGwOWRjtR3heASTUqJv6lyW8Oznz8neGRU8uoVt
DgW3hMXT2dGCpEPhR90hlV9/VtaDbDSPRiCSU9qvDt2FIf1bLLYLn9l4nPIQipkd
FBEKa08dzL8rKLwAgT2yHdY4v1vKP98mLN+swoT8NMFLz8X4fIovd/vVF1HLw69M
NmHQapKDm6QTRtbDpTw81K4L2nB+PHtWv18fsQm6F1zd/yrcs1gs7+hS4qaWI7Vn
xgGXCo9UPC+lcG223kj1mZz/o3xKxFfUYAJ/VpfB06E8uk9JxdPIUryRC49Jo4rF
vR4dmkCAa2SbREYqU1k+gKvLnaKXPqL+n/0QTGWUk6iC6CgBHdRoro8AuAj+OLY2
f0ETjZWPa9F9XmzeSSlScZf5D294Z37FPVJDBU91HTag20B7BCNUkQzjiqrPZYRJ
ZlmGodD0R/KnjCAEkdIRry5XqUwFF4kbSt0j/7tNtj5DdTeaYaYcIMZ9W5hexCDG
LCl4vRn2aXcYnezzzg55Hm1xEC3KMjQcHOSuNB4BWnze+cOB3kNc5XdgAisfEREb
A+VnUKkco0O7Z1AbDsEqjgo+a+4K+eIUeiqeMbX766Ib9b5+14PB/YW90UT6Uuu6
V3ao3X7nkYmRhBT1/F69wgrTOsGnTbmr6WQCWb1tvsbPTlqR5M/rVbgU2/PyVOr3
nqsVPvM4DqUYl1VzkKeLA9pD8QDLFdLNhqBlMXHkmKBB8AimC/Wht9PHUR0feXEf
ROn+efwVNpPoeqne2b4j+b3yCRIcHWoE7cDFghvpiq2qDyjM1SXmixXAvSceD0Yq
nKA7aJrPTRPRDzRjhn5zlLJ9iF7I7UckdZ0yDEaAfaRLsHNpN01nisFJ7Ow1Hgug
bHSdLXpB6YrIMf9oEH/It2X2nLuQAfblatgcL1NumZYEi9aySTpDe4sNnJy1gNo2
T50pqz3uY93gCBHIk+tdxET31CYqazSlqcSg2txu3VX/k/p+zaC2c89KHpc+1mbe
t/DQycy27VmznGh+TlLNYlVJqKZiHGqGYLiIqVQ7mPav/5tn5dJxYPWRIL0bnUVb
Soo0nq6OLz+6vvQfEBqpr58E16ibxU094rTMG/qQhUi7122D5FIv1lwZp8paXeV5
XvUVUpNkWD6hmTqrdcyjWBK00JkZKJkxgRBYJZY/PX1bBasHhp3ntSZtJRCKKimq
of6Fq5Iz7ZYUkj5l4BHTZ4yeBG9/xerV08UU9t43bYKbT6LJxtRER3XY8cn/qvjs
0dJ3nPf12KJ88NdOy99PLbQN3K80UBbyBj82F+HUMKPrY8R5wbhRYEknCK5riCj4
ioBuIWOg08rcJZj1yIvMHh6SvKA/4R8eCIYMXgh0nWrDUAk+WdCLoCHz5o03jwNR
ORqLDtT1Gxb7Ld0dO++RDmrRGqHnmeHhBJvKP0cAnZC53xHb/xjXRl+Ft3VqoLb9
0x27RNndZ5WwwnpV6xXiaOtIY/A8o/TB00ut8/3fhVMS6hOFJDF9i9rSrqaiWmjN
MOqVPyT2E+7loo2tCXPZX6R/K0Y9dN/UcQUMltEcPDQyXEmSaC7f1HSoBQSae6P8
lRnao/5K2+DoNY1rjYS7wF5g9APOx8QjU0cQJhlVoj7lbKGsA0tk6L5eIJ+EyQhJ
reo9WwcG6TUq9KUKlNoeh/j7JVlnqRZLgP2z2I2VDiMi0VpqgMqblRDw0BoNqCjW
iHwF1nnTnqwiErnCK20cMcLrxtqEcFwYd3sRIR4rLHeGjhDA/bauyTSwUJ5pVEqf
xX2txR8K9nD5NxKXyGBV4gk1BMCYe7lZdo2NLB+TY6rb+yI412dMt0qZOZkDiYBu
SNpikPGoqbx/9gItjVJTvc8kqEPNXLeoTH4uvY4cyp5mE+n0h/U1QYv0IcsBBLcO
SiLkjknpTfGu8DD/Jq1U/FadoPquQ01R2a9cRrpmSODXkWzdCz/cuKkkpDdJ/E92
3c0SwYfr9IQl1wt/R/NsZTbjlGhVN17j1xI5qvQi5WFPdExPhNnAUwpAXAwG7YTX
cm7mqh9nO7dh2gw53R7gGavVJXPzQon8kLMLVqYjUHbFFkqSt9+trOqUXwSsK/cz
ULNQouJFNcgObGM9+TmE0dCVbEV6jPSEjofB4ZrMNH8uE1jZmJCDbGyfoSCQjQPM
okMfGbjlFZoyFKh1Tup8I5tdPsM0FCRrr46+aEuECu05fY+I4dRqFk0107fGZuNa
6bdjrSgwsvXNkqIRr/QgSkCUXuhriCRr9qNM12/gbsdTbQPsHkRqGV0s8e/sRGRS
XOyyvzHnaDEm7KuNOVg8NfvIZpBx9mfgxupMiAd+PWcJXF9nuOx72H3bzhL3FocF
UstvnSvnDiCRC2vdDcPk1tGBWaLkX1pSb/Ypiy1yh8IS2ekxzdYD3ZFnPqvtFIFB
jz5dOZw2/1HSW0rojT/Ucdt7zzbfkpG9UnTfgEhQFyS5+uuxCHHX4F0+8V6MUabw
56hGX+g/TXDK8rz1LkAmh/vlP0k1zUt8+KHI2nH9ZEt4X9hR44hzCIjSZl8gY/C9
NbR3sVuFRwGyaco/KaLU0jB+QIcZRNuweHFM74YDvcmAVZ+WBpEqNIh4b9j6U1/H
nxIhBuNv7r6dyI3oC/vmjN+RIUCX4/V1ZozEfXiUBZimmMfbjy7HvjoyZ6SyVQAQ
Bd6RtTxfi1nIThpF2yII4qGZBxGfPLTWPcQ06rPCgk3Dy8llO+McJIk6BtbDzvNP
EDEPJZ3IrRH/zjcPDqEhpnI6RbdyGw0VZWRvGHvnVs8dMvQ9FuW1fCieiO4fVgMV
YcA/26pEes6sswSZiw3GfGJr6QnlLBY8ym5v0wy7pNArUEK8z8LAJslAEjxAJvC8
UEjaWdbPh7Yvva8DIqMlKO0i8A6L1NwM0aP522k8E4lq79/mzp024i1cRHmvhqh8
dkh5vKTOzug8NCNksgy6A+2SqPH8V3mgFn5EWJrjEc7M3ntIIoQ5qRRyUJjPCfB1
Bc/UxCytA8gDDPAM9mIgKHdUBJhuBrvG2ZVrYGvXnrQaUDj0YwFOnCQaP+b672c6
sDamdR0oQXSmo54TZdtWgadJ1r74eyW/7luRneSQmpfGhVMus6mQVsnmI5viUybF
LZUITTo3bmhsZtBTFqqkxf9pZCf/5WW1mjJ2rC/ozS3DvrcdffvjXyaRKye1cy8X
l04ZyW4rk9Cb2Cdojox8vDO9CiDIwzMPYhRetU5y5kAZkx9bFl+WY2HEyy2dBo7l
JwgLwZB9UYJceT+4NYB55SI2vYUCl+GQwJgn2tkB8zzugNzTWAiQ61rfQJL8NGet
EJl9+KcnUcuqAZXZmxYDj+w92s+0lYuc5WugjsVifHzMUCIXGPHIGCaovDnO3Z1X
/S2Knbbx/zgcbHLRs7K344ME53WR8vkbjTRdWwEJTzebT0sKYMEe6Hd71over/iW
VrrXKeBx64M/Kpkg9XK9qU7obDo8LprP596SmZCo9ui8fyMhL31vCQ/Yj8r9N26l
qNO8wif8yJXlyXnUk4ucz0EjQDkFBMqlckS8q9kUfri13mj2CeSdgGwxFzdaiFdD
OFTf7cz06ZX76vdetcDGDUj2yKKTTtz7R+C+gFyFDVvckoLo22sh1FfJ5ypz+XQV
Ljc8l6jm9n1qZ2Bsr3ETKgrl4oiGsUmrc4vPnB+e3hSrGnS1GJeNY0KNHmD7QHE+
5Sc5hat/nxIhfWZCVqDBRmBornuNrAbLe3puR4MizQhYeniZY4T/ZeGJCbZq7wD5
AMTUIPsL+Uv62aKDXSmoDPCuoxzODDU5Q5kUMmZ+UmnTSYM5FUG8zkNq42lxV44S
3BYdthr/GQ8OLnzJTttvYy0CXXfuk0FDxfM4vqVm+x61Sc199Vm04BoFnYaycU9Q
je2WOL2i3yx29/Ro3VML3K5U7BI7JxhkmhFQxdszRL3wq9y49bHHbaNEobM/e+19
b0NDuvQedxpu+FF/2yb/rqLzGeDk/GWIleL8884wjXcwBIi2evYWLk4dxohpeWo5
mkWpSzzwWGAa58Yy+0ADJRiYULxCp1mgR+FOY4F8o1a1SmmOMNdIie8rZsu7tmfG
4CDO6kBAUgScCSfBmbS5GmOKMhm7OoWz4FYL3Gv2dt4mWqbOAQsTYHAfHoWqMVL6
S7Xel82yBu8asNNs83OnbFlRsln8MSxYPkuHYuacfBHhXnZzKdQ6SC6PGKuURXhX
OMXjU5d7ZKQhUxrDZkskqHaGnk6xAgIMPLHtmpQ1LhNBfyZJlocfJX1gIfBgKPLm
/3aqxqA6bniRUTUhnD1IzISEjYEixfTZgeqf/BVKv/HLxDciqIB4w03dii9LKg4k
gGz72blnUkM85Gi6zoWGqwSZbJJaIGo9NMvVkNFxhJpk6VeEeYibArnYlWk3hHoy
Lpn7ujnJw8K2BMe/MvRoTBE81VwGZ+WZqVYTEp1jZNQXovRTMOaiyl5D8DNTXVFr
+eu9lYFflBYnVuH/MVpyh8kHnrGlJ9mftuHnLIl3+GRZ2eSTxRHiquIWyH64QVXt
w0JpsJ6R6NmQV4YsGIMK9lptSJIe4Hnpwvo0vGfrsPCycgF8EBxORblkXo+wDmyL
iP91L9fTZ8FbvQfbdDV5ZnXjnhegn/tWKnQ8riTr/y93c/RY7gdGDsQXkHfSc6f1
8VGTRSvDGCuUWS/ZYQX+rJ+0pn8Hhh34xpOrKrnmbhCnba0JnxPUc+S6f/Yum9yC
KqTcQOz9QNF8JnoDbHxqa7wjt4Nlv9rmrKSYJDgPaGyvXSpIdjbKLjiKdw+pV2ZM
7ZnnKSvwgKYWNyxER2WlbXLwWl/RDb/1/kbm50t17GXr6cZPmmkA4hsz28/nrNsX
yS4G3oQHnZkr4xkYqHi6c89wXteAjcOv/+c2eYF5QbRFShViqiLo8hpyDR0Iokei
M0tei9fEa4o8l2/fhYqXMHXPOR8zhJ/dLGxyyHJKb7W1/CsAPrglboVyKzHPNL/a
VSXRt4Pq1jx45T63rtK7DcrYZ/XRzUfKqwf8PJn65XUY9rrdcawYed+smxCxUKgx
znVkCOMPT1GhPzrdMpWX/2zsOmwlqrQcYX1Tj4qwmqoGlLceVnlkB6a+br6ezP49
Xt1NmL7QDPA7gfIoeaziNH5wmJo6vGE+lg3DYoZrLZZYviRsD9SPdBpYgygXvE69
/YxSMyWdsK6i1aAOTO1OOnFecaYPs8LKvK71Rsm3ytxjUh+CXKpOuQX6G/fcuOjS
ZVQmytwYy4QYB4vpD/IztialUzhqCShwON/d1McI9NWCij0wrt8ixhPEGSsk79zo
5VYAt18B0udTOWOzuFA/UJ50Lb1oKyna3gwE/OOes3tFvSdG8vk2Pfp57qosTHe+
UiFjeow5KOazKGk/oO4ejF7qZI4VDm1pPrF9uQvlLwOxsNnIwoTfDi1/QqWTmj7u
GJWbLfmaKmMFFDZDRo/b5/YHaQl3IFnskE7cX1qlDZLvwH3NyCUlvXR9Ldrn61oJ
6bvqdqbE4t6hNMqPLk/aak6Huped9YNhOxXu+BdaZukgFwSz6v1sVwvou4fpvNnj
qKwfDiktWkLhVqHx61KsaPvKi5U4sQOpsFNpyFPcpXGUWg7YcG1C3eCU6/SqKGSi
aEVZkISVh4AsqP0jaxvMDOSoerysDL1o62cE1yBQvFgxj/QY5PHBYRRY7twgtIB+
C9Ij/NXhKmiJfoxfjcaEvi1CDQvmvbOycSwOhSN2+Srn124DdTm/B+TnCEJVD2Kr
Ax2AucgX17NxY030Z1C/JR0JXCKxvD43/X8wroSJWzwl+vZ3zGGVgdXg9YF95k4K
2/JAsYvwiW5HtW1dQSY6EChY952RgH4Pe3nhahUCk0MoSt9oYqvdVgIm959Lsb1Q
9+8MFIRYDnPOXzYKRqIO5l4+Iq+3Hs7AMfO5JbsMNM0EH5vrmzfKYQBn2F9vEz6d
mWMo5BHOIJgSGkPB+GAhGHS3ntXMRACB3SrBrcdHk6EEbyXXv9f/pbjdHUlhUJ5m
hD1A5XmZKFla6gGrqmsqAXAd4F+hsLIwbPNy6TbkNdQUqSD5ZkWcyll7hzGiK4BR
IOXftFWIdH8o5ePPFsxa2R8Dx1ddiweSMubQQX0THUWE70cKaLysJUnEVjke/cWI
R8L7Fsc00Gy1qFIu4K377tiRt/00h3AiClgP+s/Mn0OWY+Gu9sbLjGudNWADvRy7
Y9UDmGN3HUzxFf2rZ/QL65gDR2RoeqFZ4Ggp4xJq4616hXnBVLenuF423Z0qU52Z
6i7MmKd7UaC5uDbSPosyLaoh46we5rk9MTzSrNzgRJJGBxUFxYF4lW2QayHWrM5Q
iwcaZItfZ3NP/PkWNYYtE7iBa4yKklUtIHlbCKyvRzY+VZKxrezFJWV80UN+kG5z
JOoq5dG878b/YWDZ7hT4CbPK5XrQr9+1/qzK4hwE3OiCW3uOMwLmIA7g2ilDEmnC
9w5EIl2TjjtFO02lPKdb5782QPC6sYce2RgvUgdCMZb3BEedVn/3211D59NR773c
TKB9ua7Latv3JOHPHYbQVYtlC4c2O0EQGzpgpNzE0gvknHVCzI2gZgeLU2npTsiA
qM/bdlyjm3qrsbW5W5UAU3+iUiYZPA+fIp6lG5vJMhTcrEhZuafUlLDbsh7yY05F
uaEHyev8i7gtMRolAZGiz6agkBtZ1wps1f5dS46OWenUAwVoEPzxclP7vdFdrLL8
YIi7xkzx1rw+Po9u/VKNtBjoSnqQ3akR+vnyDZ6wmrjUBUlFfrbDey5M78ZH2TKA
kMtwaURyaBSRi9wziEMidl6gqn89iAG8wWaP1tnNarTObA4XY7me/xI+OwbsUQq6
Bs8TnSMdoXfNWrN1o+oxwSgl55XxgWiifiV7Q7d2CuxEB1kpvMuRleFmXDe4Nfdi
gCb+nZfOn/uORLlWvok+bcs/Jv5IasrD6lsA1XHC6DsYbsdGdmQy86RTA+b+aTqU
vO+q3258gO9khj7Re51cblWkx+Sj2TgNPUe27biex3/r4hiiGYscDPVTRdqU5e2a
7xbs3TCRWTMNq4fQiSnVpFmaXL68ejXqF4UdGF+Zi6y7DU5Cp24HDNhwdCU9N19W
okTuYdl+/3mYg5QyTYy7tnNHBo5Y3AoUtQBZ3LSC3q8kGSMroUaHtm+k6ZZzv8rP
EuIrBEDNnrVxPIYDUQWhtpj5JxfEuRS4H4gO48crwZi8LuPh6pSD5ZcqK+9S7gkN
G69nLb+PsPHE4dGGHtIWmnR1SWNJPwXH8nBpfgl8Hhhu214GDFObcdCIQnJ5nl28
4OFj36UNMzIOK2vlY8DirEi+QPxUh4WbBybQqGtMjHcRArAUtn3K5AKUd03/7AFs
pnOo4kNr2SgCDzntzNOUSIVjsiknZ2QinSHJVnc0SxY5GSNA6uMpksnmlXZaQK+c
QHNsZVL02aD4l4k6Y5mk/cqZm+PwFdz/3Zb5mDhwKFHn10Bc7MWWG/BiMmDE6Ehx
kifNHiMSF55Fd3Mg3jFxLb3dY4nUggaUTjF2jp0f9SyIV579rtxmJaTh6seI51/a
4WwsNuIf3X917zYwGkBXb9CQhOwioOcEJdb7kDIwKvYO0s908p6ylULUxUDeVNsS
68k7yyFxWOW5d/OWGzZvPn0M2HZp4GeAvWpLwWNlsoyCoFp5Ouj/TVy+9YANlVbf
cheRjOK5aEVGv211b8hwNk4EkEiDHnJloRXnZW8gotdth+w3lmNesoaxn8XHUwfz
X9VCWwX3bmTaNpe8mCU8cWK+W5unathiQ6R4qxKc9J2bsNzEWeRB36BRi3U9LD4a
ETgi8/rmrCbG/MLbsA81Wo7fP4hYB5IbMXpeoY6o7SQwgg1pJw/NaolHeZlixObd
U0XIt3VqQfoF7iNx+iQV8mrcoUdKBz3Wk2P84OOl4s45HYXbX/YimpwSWlEWMUzd
H+sPQPkt/XkS3U4FZq7pojvFMX5kwUyqsPSv3Ln7YHgMbUxDeNXg3dNu6GQwFlFi
oCxiyuHS4dad1Qh0BTU7pd1celEG3NHdAwZdMrmEvvDxL2dGq7oXDT1vissn5yVA
xbCXisO58F4QGZs0SUgVdmA5nirovlYq9bBJKHqIbD1xFI7wJc0JazFyKbiUkCGn
iXnmy/vKJ+trrmocTzha+N5AXMrTbC1LkasS0K4ZbIllUFhwftpk1WXvekHvaik5
pj1QBgds4WSBT6p535f/Ft5Z9G/h5RITQHAgMi2IcljCh4RwtPe5NhiM5f9z42BG
6+eKP5Smb9wh+fsnCqACU2b+s/lte5BGDVoV9lRNnHF4KctmOU2a+H9+kcYHBjQS
9ZpEtUnjVEKxITOV8oOIp6/Uc6jZnddfGddaLLiZQDXdj5WRlrPWeyBuWrW+PD3m
llkUkFlzH8pWPm3unsH6owc9MJDJQEfldjZU0oJl76XVcNMopDHVWU4IV6fxSmTT
eAx+YN2V1JUpsLcQ5yXysjQ3/v0V6HuYQBQ7cNbZ+PI5SSsV98CQBMTxKYrUp0Uj
TGJmHlV6do5Mq2I3uqvIqk8wvpqvQ11cRuh5ofl8chkgh8DdvAO0pKo0H+RKrH0/
hWqJ6W2B/tpSzT5qDAVl4Bz5Zs2rdBRU/7jz+mMAIktwPhMcnvTDNSsueNSAfzhY
X37JOVFot122UZDklHQ5IOdqGmMLrWt6PI6N94AReePwLOesb234yrdnlX17dKo8
yPaakeqqYfvYxidTGyl+0mBzqdNAobvbdqGVsCwJwiG8XaMUad8Ij1KwpP098Ggm
RHjdFjoGcT46u9ID2M7AzFhRT16rOqnjmhnoOtlChNUPScayNq9DKWRs2dUHr6hu
/g2JBLMptIaMWqHtvtAv2kIdX1p4ysFkPgVY2/M+ipP8ycpi2+qlQvXEBkx0WjVh
l6E5W+viwDuaK8+z+QuxnTdtMHCJgJQna4+D0Rn9cam09cq/XyVyYp9LfnaZxNFn
hHfjnxItQVmwC1uYwxt1mctWRGDTBrNFWTVM+5NfxtD8AoYCzzu//RA8VPQbA9dc
jJjnnScrd1ZoOeJgEsSU1/IKKQ1Fgtb8JPPZvFHHmzCfNDToKz8OF3bf05g5SvmA
7pq9gr6+Yx4Mh1SEstwmPeMkCLgqMNFdBmpehJawQ2gCye9skPB/okC/4qY83VVr
2VIyWkyyKA2Rnz2GVSveIUen3ciCgEXDhNJzZ6dmswUwnM+UsNiVAPHQCuWONMtk
d4EcLm5zlAAbTh6v5+eSBABVg3pIg2yIp9O6OFZ6cjdAktoOmydKJrK0Rt0s50e+
6YWXsA+fVcQlNIbJOFxq18+ZEy6/g/uJUjY2Ac3M2hLJfKnLCUHtaVQYUue0X7Dw
eaIsMuDtX8et8/Pk83BbYbvniq+zsawdK1xJAlYPVE4U4Dg3jprn5pd7e0YCewPs
rY0qdnxb2aXzZJqmQcDrWdlJ2qnG++UT5yB9yk6e/z07swZuMXQJTTtuMOorZR5t
LwaxP7+wz1HumVDii7SKNX+j/YC7zBLc6Vra+FFWfGv4paH9sujPMmMRYYRIzAU6
SnKIdpPQvlLAkTdhY6ksytj8/PZJe5ZQKR0/q5Lx1yGYDgBH3sxI/+YK1MfLiyec
Tu2J0JEf10jslNZ4bCoSAopp4LKmoi+ddXJPbfzzb+V5dezNcZnlZ4XrVqH3XpDL
Yk4mE2QEKtoYpApIBKpyl869FIZdEB89oV4xKNeTb3XpELWDXSB8q7NJbkRl2Xdg
rhH8M4EOwJyhldjcdbyadWqpTx4XZnl3kk6Q4HabrTprRBv+giIeGe3ffzv6LK37
61Wk+KfASb9W9mVKIQbmVSmeV3Jg9gRZRJt2rzcbGqcPuKGcCPSBS02UErBMYPG8
sRm4SDjpX+TbCgIQSverBMUTbd12TkGTdSUbamks9tb2BSonYasFIfJ3AGtAWFLl
hrSCi0O8t0vsO75yvsjhumN2rVUjXVmOQrZC9yz7OiAUBIWX3oAIoNeYDk+XOVYQ
OiC2GotJ1Y/0Zx8biHZuyXmOnNvZomogHAZuQqtNW0zA+5GjlP3APbhTb8K1YP1u
MQfCEExIJN5X3z6RbM9QwSykr3xalcBar8vZMjEHfSlnWMsu5feFYV32dp8Dg/WJ
W6yBELtVxF28maW5WHXEEsWTrAI1iGN1oku6MykFibxowmys1xVxnSiQRjoKvXW0
JKlBPnNKUrnD0L2OHFr7BnOvKmUMnqr2m8hxdYGKV63Lxl3LBe6LqO51OKDaPmhq
7/3GvBjqW35FD87TOF5+W5wUQcuXh67IHaDyV3XjdBsVM4CbNsEqK5jwrRVPg6lb
u8NgvIHRFllYQz45UbVfVLPOYwhndh0n8zMt/hoBScSlYDqqAx8y5AjqSW6WgFnO
i30USasW5tlaQP3duZUQZjiDOZOKdCO/F6fXbnON2fRw+76FoRGcScd/U7t1F9MV
jKwbcZf1FuDnZF7fUN8GWLvbzGJFxGqBgK3xh/CzRaxp5uFDoxq3Tfj+A/t2paH0
b+VN+dtx0kDRF1RwGmLBIE69rGxS5VTQgavzU4MK7MYfhXuv4b2l+AiRXJPTlW/u
a4aZnZD4KbtBdcJIXj7rwE4AiNLUo5uJYygGkxyAsYJSrNTzIZkjkUpNRdTM9M28
FgqBL6jXAneOpeHoFTfbMm6kHGovjxcczepyliYzG6s6t9ZVIXkKQFM/wOQT2cDx
cxXsycps/G2aMuqe+Kf2NDH4RA7HWsBsEMKSpPHBuCu0ApSrZezuvbXcdeLgEyPD
5R+EbDmvCw6920zMxz7q6daydjFSE0sgzVOIf1C3A2/Fsd8bivj1kF7Pn+DWCOVe
sF+kjAQ+va5wCTvFKFjvFBGBTWiVYrJkB5+nZAsL3mS242cW9O5WgMHqwAmfQA6Y
BiFdwonH1Y9V0PXdzbGav8Yn12+zbmdnCDKO7g5rPuGfscIPleajIr6BLNkBlyw1
n0SGz93gvUfEMFuPw/JV7/aNFhkFsvOHbUSZQ6RhnYpDYxrT5u3XExmxntK2Xkh0
Skl5pGQWzGObzD2eER2VcRCjLV3ye+c0nrFnA3p5P7q1JF8jTgX5I8LBrpw4YjO/
vgCJj037bblooL46FQU5ImldNtSPLg9oBFHZI7UtqLl/a12hrIq1PfL+G0iUNuEP
b2UqeGcH+cZ/LaZHVgZOfQQgatllPPWR+uIZohXaBhXceN8gelQNRl+4IOiKqkxb
VfZSQWGbBnC9fkSyKglghjmfC0JtBMuLLg5eDAUtfoFs+8v1kCOcyyCOQ5OHgH3Z
wvf1RaZHAinnrafCLtrTRFEu988mmDZztfZAL4q2LjMWGCoaqLHwbCkovAY6mHI7
+/KM2aW4uzOU8V7kRbrvgSlyOc2ayyKS2R4ShDNRAQdSxoPs61xy7ro9Y/w7cenf
kFoOLL6wTtXEIMuTKUyV658dSpoHcTx9QGuXN3XxwWJZ4xmaLcajmTmiX6XmpyjS
Rpv4NQA0lL8gSv+Hh8TcP5j65oNSeKrVjYQIEHxfYi/ccFtWrUIdPHUP1XPSPKXc
tdhvHCcxsYgmflsShnghxcBhKQC454xTCvTdAPpu5fwfzTzUw1V3tY6sDN41tPom
G6yMXTWsXu9wE4rITE6we2JAgb7ZLhM4lEjpmpI6SdrgoH5Bwwo2D8oGpzdgEii/
5inKDWTXHWnJV0IVhp579Ju/gLcHbI70Ci4L4QfBpnPt32k1S/q09GZwTtrYko8n
RYLRljYhpiAc5LKAdftwaTOz8VjK0EwRq1QtE+xaGZ3Y8qXf3+nB+J+fS/jDyC0f
aH57JV9mxUA3sopevFC7Q+CO8akM9VqWmGkNAxw9grRHRmvbjBUJdLHTu4Nro8Gy
NN0ip6CHN/nIt0u3u4MfUsvFevgHDy6uE2lfUgDGe4NCB62f+WA5mFFfYxW8z2r8
o4r4JSOghdn2t3DuNSBHf7IDEnibcWjfBElPPJzsbZGFdVJgs1W+1U1G/9+fKNQt
OkioWuEte7L5tZLx/6oBGikrBiuSbDj+az0O9MkfdJxM+Dy7b7QIhrcu6Kx7bJdw
8w0DEKGdDZB1ObW508mQWqNzjhh6GK/Al7Ah0IULTdD5p9rirVZO7Txmsz9V1wkY
VBgQ05PQnOTenBpkbaQlMBGNj929B1g+L3MqWQb6/OsXHMpw1Msu9mg0Ok4yNXpv
8+Blrq2sag8v0NOyUqANyDAoPcs+VpXGax9/em2/wSBx9c/vtVWdentsfMR83iIC
YszGjaEpNF8CGYEnbAFk2J762JHuQKByqk4gJ5R9QzFUTCKY8elE+6LNlnJ15ldq
u964VqNJEw4irdmqB3KePLUk+fj+ZhN2EHWv5rvlGYsSfIXEHZ0s4y8jsjR2Po4O
KOrX/zAhqlg3BYVUkqyaAK0kI6GAhO92qaUpP5YnLaDV80k276jWtvvhtD6wKXI3
+jhg+5b6LfjTSXhusgZ50C7zJt/HIY2bCBOoTmdYR1jd1n9C0LdKnP2/iylwH2Bl
0XmciUwZ1YsqKO+gBcCEPrP9QChh2QXw110vixHPKBXVvWZpYREEjXu7lmlfPyUs
9r7VdnFtx2yYuki/tfCZzYm1i0nEAAKmbtRWpuMSoy3gN/rafMyfz5us0RByeAGq
caTz/fGwPd+rhHUggaffaJBh95OxMUDhWwe2vpKs0AXXOA9bhOwJf2oiVE4X9Vtx
RZhgdDIiVTU4K4rPy802bv86EzUOi4nky6lH1IpQCOYSbAoTiXiDlNNVwAHdoltJ
XCEru2Fps/ZWS6C14cB69UaZ1L0Nrww0Ks4dZHvMSBxUNqEhrw1kWxkXzilFx2In
se7IttBjSLR5Tm9LruU/EgxeK7m+tg3pvOXkuveK9i+QlqC6oM8ErPVOjIZDsVAO
89/Zwn7QFjgjpb/OvEN7FoIzMAOq+KrsliXf4ZKVtzT1hm8Fs0DM67Lh/NMOPvDj
GgWQ9ds8wr2qwrwnlCft5w6VbEWFVJP3z1Lclhb2Y8DH4zMs+QjuCkVRi+n4aJU3
ysj/S+xlHBBE/LbL9N008EgfeBw8pWaI3bHnpCIfNg7uunKnLfHULyzaqP4jQ4wB
3586pukZTCjIjN6C0Gk30xHoMUDw7fdqISb+kZRh4S1Ixu1IDqxOs3q5eNqMKJYE
4USUNjfDu2qx3bXdjpYJ3WPqZKqhUQrI7QFhuCKa1lf17Y0PZ2Cx+UqKtRWFl8Wd
jczuF6TeyG96qpOIX/cSvPdkd0SVirv8Eq4j8KEi9Xw4CsMIEVYhG7WVJNejY8N3
pWqCxPOFBMuBtEUDBVVJ4RjYQpwL6W9ZVyD/7Jd9YAiNQ11/1esS3ZtxqAEpOAlx
rgcugnurXls61BNmV3JRzPLx0Qm4oQ+QvVjh3VLtpqpVUR52hj34hhpiZ19zu/th
gaiH3C+Iv76t2PkcpNfVsLv4tJ/VrByAcvDpN4PMwfnnnflW9hel/7dYuBwBPLZQ
wkMdIBg2sRArOVJXZmT8pmd4MNhRWhCfU030H+sbw26BqUc1Lvz/jOeXqOY8Ey4i
sTnDmMGlJLGgsoK1m2E/JkVDHWR1palGTVR7DPCH3F1XW5FtpSY/BhcGhQHrng1J
kzIzUCb4GKOg2rmAW8tKdLAvc5rD4zWS3O7pFuP+3GXgPLpXnAo8JLVN3BEpLHVC
YR3KEVJWSxlpM8DYnXnWWpAyMNxQvhlZhMRMuIxQTVvMYMFVMHFZnMlRWm8jX3gh
47Gx4pl//Ffzp3ST5GwjCsN9e7pFUDf2ygCr2oXV8P5MTMu2H96F6jijrlr9KgkN
IkPG2HosP+pB+H2OrRtUEsapEdpKkpzZ84QC2WbY52IlgW4NMQDd5fCMtUwpqvyY
6AYrS3dGRz6o8kVkm+ixf3UsCJ2tChYOc/LYMIqZ5a9r4LnXmjkNGvCVKAAb7TFa
E61Ufo6nNqWUZhy6LAYEhwpJXoNrQlC5DoiaA/7MRrJPEDIscUZHGxXGDxGkbDEA
pcbhlpqWhzv8RMnZEsIqRH8TcgxV50qdDo1wt/VX6QypP2OMbcmzds8iO4F3KHiH
KJ38f7ftSvHX5TDc8FeSfuNA5XMlo4bUKjclRfsNFBor9lYzdrY5NPY4/0Tucg0n
hW8VPqTQefvE6ZLtQvvZ4A4pjdt7VnvvMNbiUxQIMYef7EqRAb65GsENL6P50bbF
9WwSajbLXYq2XG3X3D0KLLgBYrM5/T80Jfbc99KpZaP3VDalbUboWxYxCcH47kLg
xSJJaKs0jQECY5TjygNKQpqqcjI6Gv0+BQA39RntvbUkW+++mZVdQ+UmKKpG0Gt9
Oabcn2pE2sp6TEwM5Tx+VkSP+qdlpx9hyVxDdGC3sFZodIT1DIWX/4TvYPU9nRtc
ndgD377peeg9T0em1xQv+Y03PHMdfqLZOxaAyAO+3O1DdnomzaUl+o0ZSI3w/223
Uk+odV9U2ZbVvEAkDZioHR/I1tpoVDVfjxBAplJCd8+HM9B3hVQRnWcma0mVkmPV
NftbJjBnZDz05v+xVh8Ytex1d5cwxToT/gEBC8leCmpi9R2rnSa0lACT1/CgcXzG
C11r4dPsI0m2kEYBOGTK/61H5YuN+UFyMKjl9TbLHXhNPmnChlScr15z4ej4xCGa
etuUYpwgjXOVpwD9m9TcQ4I971s36GZTeZMA1SxNvtEsz24A1MNMrrJVvO/IRDw7
J6t3Czc+4J2XXWqE5+/Y125TkgcSE0900SZJOqW+KiDaUm0QLyhBDk5E5iYEMrsu
06763VXz4OOUZjdL75e/5dmSD3sGRCn78AfpZPX5DH1g9RUjQBb5Ge6xgvBlM6/K
csRSlOb6BKjPrUtfdqtmiTTgTAu9HNOkH5PIWKHN7rNo9GoICRi8XEoTRrSSWSlr
ZyEbvHXe1ao1smw+clxrT0omj3MtI5M2nE4ROY0yBxIZoL49yw0+Tpq9kD5fLhoG
OGeq0eAUvo0nNugNPhZ8v6DY4NJ21YREz+SSBvMLgqNfTHeTvgOg/dUtuITs3zgD
55ETHxuwFGvsg4UERck40/NOEdQ1VESlcJ7eWmz7vt+sSf3s/gMz4vUJEcVof877
TpUOBqDoMSXvAgxV3BmGUD+f8vwhb8JpErAY/CT3ACbmBQyv4gFtpgngsgne3ZZG
H9zyMoWC3qqlBzP4gVI7VBHVU/ODp1MBh8pnh9IOxdMJsUyFSuOmkw7UblRHKnbh
lm4QSDg2fH97SUZRtzcuisMIZ3kQO/mJ0/Bk+jA2SQXVQQpjZfv+P/KX3yNv/Trs
81fwpu2gVJb6lIVf7LmNDlCyBj6UpOgbFopk5/NRuVu1Kcu9pFoLVP2MzXpqa6Ea
7on6BXmtg/htoQgSK0MJjWpSu1IcgyxFEBLbWu/iEA98ujVbOjABNZIjOZJrC7Ba
Fhpz4yJ/FfYbYW2Qac8v/erjqe9qODsUKxtZ/kCkvgVN8rTrs5GXO/swKOs99Rr8
jMQnq2X8grSFzkoPUxPFEv0FoTWfZvdSgQGTrV3YBRkkuX4pPFnfb2ApyUQhppTF
GRAD3mgXJD8s9MSIHeZPlohuLSQZdDkmzRDfPSFolXWgViIwk22bXFTLRoJORf44
S2+X62HRyrBBlVCH2hGLaaBmYiMoElLYAY2AwIBOgHeLZZ2C7SDyCK5+1yVm0bpt
/clZMd72X2n1X5Nn7fVe1Eg86cKLO//1VYTdJPNmDa7flhJRRmzTkW4eaCCzGbK6
DPKest6QclCBMIXFO2uBgABpMuES82sUU0C2lOBg3xBhWd8ExF2SKr//jMkB3Hx6
levNw1TKR6qL0ZIBMnoP5Fzu9CM9sZvDCjS0mI6M3ogSRIDDMLZXpcDw8xjHQokc
NeqZm+8SBuYq6RnlvmrQLmqK4N9QVlF0D0nTlTPAYQJ0ktjgjYWIAcsoy9OAeZU1
fegZdWlaGoPBPdATMgh93hndJrS3ipmXyWMex8QLznE9NArLkVVc/UhpFSLyj2ya
2306OqIW8uswvtqBjnUdvHhJ4ctM865YkGyMEDmAE8ru3UiNP7joKTm0F31vLUwP
NLDkViR3pyQKuvZ0F+MSvBkzIjxwEqJEs4miy/xbLVl8hTg94+H4pf0F3OUHCUrL
BK79j+85dlnEYWS18UR+2JxpT37d0mftKRXGdZkJRIDCWecLDMbJPiuRoV1J31Rs
6nuTEnZ4Z/RXDhng43KjNGuuCgy0b/5xw93u8EQMXertOP6fbQd5btunejsWg1/J
Y2TQ6jrbGn/PgjKejwBahTAdWKY6RUHXobvCF3LCZkBUlobscGpaJw8OTk5Wmbqh
A+ViunwlH8UAefpkNksH0PXt5i40ZxRISsmbs4SHMAzKwDiO5zZenkhiFWVqxUAf
ueGH3B/7bjk3VrerYvpv+olsCDXrjyi3DtBWw3xKubRp/3bE9nje74Gjwsely1Ca
Nu3Xv/x4D4HoAqIswxmI+KV7yy2ayWUKR6QX0U4sCgOLNGcxl59U1j6HuqckIi13
5jppggVfw/CQmDxQK4qUdBRMFCGZ38EGZ0dAl1E+5F3lwdNYUqsoSvR/v9FMB0Qy
l0Czxj3D0xqQrZTadCLMptXZg4inPv5GFFRdkgCy7p1LKXv9VjgiIZPrqBU2HCxt
BkVmEtPnfea8yNjAKSNz9NI0szGok0eAtZ8+CVt31WYVlvGC8HHZCbSQuA1QsG7r
RQ4x+dqY+nZhMhJgYRCHG1RME0sqE5cMsIqTJf6mBq+jWGNiF7NVF2O1iuh5hXc8
+M86s9wGjGd+Wv10ut75XFkq277yysJ2lztzBRLPBHw/n5CZ4QhWnQkckRWc9L13
+kwAw/KLKdHitBYoh3eLcFq9YGs7K2Ivqk6TZrPF1ANs3HXHgZWHnQEwzCvJ/Uri
GWTsL9vti7LVGstsXwF01p++GsBS2O6WM2XVc124brO8pCY3r87EW0EQduyaIqc9
A3FWT8aobfY2OFvJccVtrNbnT2ngohRGO7gikMkH09lVu/dvYmqbzL60NI5fEA5V
ECbR+V7HXbdD/Gxa2xmBIttUIrwSOwo8mBfr8uwQQ7LTiI874tTeXw0//x/gRXId
y9cMkpqhKKX53LGarpSLuOMo5NhId+js+Vrsq+kURapH3Zp2gvePxx3H8vmuEff4
/dDmyZcvGWsXACaQlx5yuDSKuHJbCT5mydSLqdutfY3W6RrvJxoRaF2VLZJvOmf+
oREU7eg3oR3Oh1AOHvnpJEF8uALsLmWNg/uGZNrlzeUMy1+j1uxp9eGcSDt/S0S9
hfE9p8/gnGvUdMJkIxid+DlCIHSTq9sT5WP207STwBNpiI2CFR3jlbTlmsp6W/IJ
gKk7MAw3xBC6Q1PugxKr1NBMfQDl23cESXB+jHusIvQHVFs7mIFyFstasJOesVfI
a27q6f0CqBM4aOV44uIpSgEqpUqYMrSJIlKLUNkEjx4gS0md2dyRLkYhfagAP61L
i4i5H5qD8nc31mPxRrkWKavG8Bh8O1JZJT562Y6/WaryQFH9rN4E31kn9g/s1WVJ
8xfMkN4sbYW+8DUHWqjYkQCXvPaOG6u2XnIVar0B/dp3kjbSGz3W8ip/7eziZymK
u6p7wdp7Fc40Twmvm8p36ly67uFOaJN6ND+vrnweINGEkozuk//Sp3cCqmt0iEfj
m19Gm9yD1FswpOKKKP74mG48Jdv36vcBRa13BHfsekfSpjFH9kDmlGELY+NOX0Bw
eY+RXe8nVQJHmqcxKVUj1z7CSkHfFTtjYMfC24K7gBhr0yOSycPA/iN8OFC6iDY+
ddZesF9xrcl6ZnYRZtOF84ZKrppQ4QYFBFRG6k8h7VW+B+QdUx9/uH/3v01TZzSE
40bVxpm7zfxKk9FR4viIipbqnysqIRrb65b92WWUHQQbuhCZfUr46CJpiN1aFJdR
CSauOYJoPQvJP4a/vkpbGjngVDYTV34nkox58Oz9LeZUZtbz1uFJLej66r62tz1Z
GgaOzuyig733LLMBsW4135NJkWyCEsESGQYTPIHypr7aRdSEMuZhPvksFeIYbCWo
Ys+kGhrWdz5Ndagw1kMAAH+HKGXnikvCokxS5f2ZI17Kt+Mkgkg/nSq/Lna5Qn9x
Ub7z2vgzkRjf2cG2wUAr2UDiaik4uq3fDFD54PnVMhnxJTUag0U/ZZKYy28bL+ho
GiuIhW7jowEJOoccqRLIbpH2HpP0iEdSTkA8K2q3I4ZqWhrHSnesPudgUey3yhEX
o4qduQLrcHHAb7Cjt5IQfVEOyvO5unkqEqPBEmRMrQI1Pzu/FiRNvX7KPIjwseLs
vOKoXNAREZNnDiUVZmdhfeus5+s76P01KXYx3R02YCV1dO+XzIQP0DxZkKgX9X2P
Vzzf5jo+A15TijEUsm8CBZCYKzkFVF2C08+cTScRDZSHQxP/RTMKWOn143/Ngrw+
o0N887cP3JF4tNEerrlYLWMx5NUS34aoObFw7dKlixeBq3u99cxJyuCIrS/KIpeG
5d+mEcCI99VwZqRTjAhDIjKaa2BP4d1kQCMGBmCJcLaxcN6YZlLRW1t0/v9P66Fo
Y60Q5XzKNxDuwObF90FAP1hMe4ucVcUZHOSpUltBJ+F9zk8E/yfA3ptGLYJx1ZGE
aLURiCv8J1iyaad64KY01Rtcmzvb5polA+CEkmVJ0uw3xucHufSGu9hH0bTi/m77
vvgx/rpIMHkV2g+dXA9/7iny5+pp5gQl3UNcLqFLNddliB6fmNn59MTlvWrXEAzD
zrVC90GBJ8KJOKJ10iSeJozhybwiLUshLIdL+SFw0o5LWYfTGpS70S8hiNXP813f
r1u9gPWDS/LhTkswCZ7/i7XeQQ+4gqPM7as4G5d8xLstnkVf7N/lqUzd+qecCjgv
mInk3/AyOGJAPag30wKs99L0glrm+EM8ZdZrqKwBAGbJRom6N+VCYjyCYY8nCX8u
1rFk8vobbEyg3KHRx9X8K+APjXvE4mfFYW2aZ3J6Xo9oFy0t8YtJOsSnHey3l2dV
qlsFQFJTnQ2EF2IYxYn9OaMPgof3xzFATjn8oNWUbq4iNDn1xTDcAZOSmxcGZsCn
FAXoVtIYDw9plchfccg91g02/Vy9pEnds/3mrJMdAaLaZsoyK29M0TOrKi4AHfnN
HT3GaHNvC97/auMXFLNyXfEQ+0j9KEPJ5hzsVmg02CRgFzw66pa96+AgkFsteyEa
bKc8El0S9ntiV1XA7Z5Hp2E9E5i6O0MJix89+ETOyGNbSeoxqKAhOO/KMC7e2Wii
S0p1XAmsQgFfKDdre7uP/CZHQRT5zp8cS3ieBGu3hV4d+QGjhNNL/3qUMqsFN78w
bMUQWHnLQZnvZ+ncXS53KmyQMv/2wuVi8OD9nxyCf1VfGwtzxXTfi3G+6aKJ6ijY
3s+zSuUW8X/L5gsjZrYLy/Mz4ZZpCU868KFq04i3asLGRPPjsH2JViDcdJZTug8l
rcfsxQA/L/TNO68p9dUDxJ215jVkyHt6XFHUv2q/O/fTdf2to2UthntoxCKzGjiT
WOBAQYrf+Zz6HwV93XaNzjhOqSnQOOz8n+SD6oK0jdWqaYDRNtnHKqt30tkKsu+Y
uawGf5RtmQuSDtUZimztkCb4bTtivfjdFw4pIa1oitfNPF8reuuJotyJvHwxS6Tv
YoL2FBXUhNqmvw+SK8yFHycKeS8ojFuCNkB9ydCpwtd+yAD2ydlZwQxoXMxQ+cH8
0PYJ9TUeymEALTEy2EQqt0ySKu1d1nR7UsE1WzA8wikKGFLbuY0uBaIKKP7/Agsj
35RK/NmBt+MVKAunVBhBj5T20n/E/0LTeUAVI/nmvM6/ZLkVquZXLSsX9rsp2su4
LD1RMXl10C0mEY8dJ1F2ekSQkYEfpCj5Ujv3aMjnri02cfNZxbRKGi8o6IQ064nU
wuzM2pXuahOvEVm4RABItCKI3W4okaj3tGkpG2QzWhTOpfuPjMVW12EodhBTCrdp
qJOpYR8XJZnO1kqyBL0BhHv0Uf/0iTouvD43jaO/kRIE6kj+AONA4xcnp3stseSQ
dU2ZsDm10XqrQlmrm9cTOHywwyOx6rw3AED1jGlOZVUkQ/DFWWx0DzZbgwe5/fDp
z+66TTHRvPlMDE2Bg2dl0y6W45eEqcg0ionlFKZ7AZye+ugqA1IDSrpkikG7jtYM
Pn64A1Sb/ZbVlPYzg1eZP4xKxq242UjOupM7RnkrsXlsRolif8BMTJh3pSXi/5GT
+6ok4mGd3ey9pzKoLnMg9vwG/RO0LSqFRgQtglLRy0VmRW2OX3TF/yxcfAGCs/uq
2CQsfq8LTFTbLE7/RLyKa1IEwh7900M60Dw2ZHK63ofVBIV/1UUZMAWQPQQA8lzr
vmUC3KyZaw+LU5XobdluYAAKjPzpG4i7l7mdMFgeIz3UYtE0k6L4tQun3aaoCEH5
NuRs9wOl8INsDeOAAgu/WWvleCeVvPoppWRdSijj1fvaUDPi7vXyahhRbK5tYTkc
bx+BXQ+7Vd4XP/jhJWw4M9/MeSE/Conte1EQ01pHlW7m7XKy6uiJYPCaQAuYy2z4
A1gdkl8mvUyLzBbvjRhdz2VEG3SmJC7H616QGmm8v1DaMfDVCelRpeWxUCDfqK9n
gcxnA0u2XBEheRBy4ZHTQjO6SpDSLqk7rE5YYZieiqMNCfiOCpsTSig9zGhLyBi/
3spPOCM6jWuq5Wxuj0hGfuQmETebZmu1+2YpfBQJPAKnu4/FzyYxGPW1PB8wsa1d
cO9gh6ran7DgTokSMSpMhFtQc1zUAc/umPugIo3dz/7STzfIczNGHm/UZEa3w0K/
KXvVWvn+HbQouGUQ+0cnmni4yxF/0hgSDTBaxLnwWMSfHCVHCl22oIJagNeqyXRM
5nz7Ngv6HqefccV5uYOvN8+TjS4jtYyp8pbts6ifDygAuAwclwdAicPlrsPFO3/J
zudqd2BTPt9EsqZGF4pyy2Qw7VumLkbQ/fh4UPiOitYIj2co+XAZncmQ5gmHysW+
i+UFYRjeH2z6dM9BUQBQ4Q9ZatPDc8HRmaY7HT5e+rQIasPTRB8TFNHGmCFTM/HN
SGpzm+1Vql+49uFLwrpM4t7QQuTjAyz7141cBoKGfkGPYzfz4/K6D2cJXJZR/KOl
gELGJZ/iJ1pnXrTVxHTfTRx3TIhdKPNVD7vvLspVw/oa0q72XwdDiB9MjIHLR+Yr
ruEKa3wDvjjPK2GEkBebiElRL+/MFXm4H9q0EDS5DJJsasXlIllDGM0SC0+DRXXT
n0MWpR/cqSugNnQWGNp5gmwt5/7sGYxSPtgluYNGAHA6wPCrOPCMigj+WoUl7YCK
zHDsje1xqFUX5NVVvcGEJVn/YzEOSHmTjfwDQMJc3WqqCv2Vs5GdtQRj6ZbNzTuN
Z/R6cO/VXb11XcBeG/+n8hq5Z02m0OQ/QD6Z7oGCS/JEWfw9A6XLUMNHRvR/at2j
dRV2Mkpn1Wkg9IesL0zQo6YAyzy5ASkqFJvrYArq4etKC1JQEyXIvEv2vnuCBt4e
4YuGJizyouo51qu4yyq5NJzBwz8+WIO5JgUd/iu1bsBHGFR3NdzybjP7BH7xVYEt
E3Cey2uD9azY+TnHnRC23QF50hR5aBGAiBGdLKGNZdVga36MVS3jl0TCg+Bjskr6
1+NQAtg9VYHcZxiup02yqWO0gM9RF9RdCdzPBkf9rm0hWhURV9vm2fjPZJlAtV1u
TSE33SM3IogtNszScWTnCGUjD8E22fFynNgz4k5lBQnIFggCJZwmo0IMfeEmc0Yl
+lhWxRNWM6g0Or9a8whac+k2W3lBryXOhXS5DGPGFQKUx9h0lhk0+o5BK7cvXc13
9hi3+tEbOa8z7mLowxvE1f1syzMkla4vipo5qVSNriZVASdbNysuUPPLQFbgnBT1
hF00av6sZZobEyvifopxR2IcW5sC+lR+i6KotDC3FpTZg+PHP/KkBSfLjLte6mli
pUqJPc4kK3drjCGO80f81kS5mqnaIlBXfm7QQCoRf/Gb1xKIfw4FdCR4h02m6Y9S
tj+cbHPy93n8r4/L31o+DlPaynxfmycj+T1mK1aloRrWKxGVn6RRLjTg7+sBccsv
ThgGxwUka7YWQyw5Si4xj0JrRTlkkE4LRB57ZATChZG1qaIBrJoWMVnMN3nMrWJj
Y1fpaxWtKWq0UzLlJKh52UWW1Ye8bgWR52M+jXk4i6yQrouu1wcZ94odLS6mF1tj
UfP69iZtQnz8NnFmuaHZCLkdDDz1seFJL9Dr3O57nYcDo/ntOHhpQgu3Rks0vHhU
QR/uvPKEjSwmL8MCjbzRrt5WrJVDsg42O47TGEF6TVh14iSy97UgqYLb8bNpH7W/
Dp2Xj1h4hlhNm34xsHJcKutLrp/kBzqWS+cXqWiWtE+CtVylQhYTItNXF0vpSy9x
hGNduqyhh9WbkFE0D5igOKomXVysLuKQGSYD1Hj1YZI71x53GLXWixgbnHuI3YWo
9zp5JVc3n8E0Dw63YLVLSQ+FLYN3yL5ljgy16v0S+E2Rz1sUlEkD7jR4ykkE6DKU
vKJdognmKss5Mjf3rR2dqGoEsbrFOnwblyxHh7nBl1Ahmr9g2b9sGvqz26GPdnao
gzpls1vQv7eF9STIjsmR4opMAv00Z+g/02uA6vOqs9UyCCNqQ025ilO/8LM7h+my
v+SG15tIUUAjwaaOvBCItxurxYPeMn6URyYNBQOF48zWdF5KBHEV/KjBkvB8LJbh
m+HlXGZK4TNIaUGvICSOomVDarWaRwKxJv/i88G1SxB+7WDV1fX1Azka2pM7QYA5
9Jhg77xOeJ9vUq/9Z6us1BVIhi9W69/VJAzdea7LSxMyOry+NC8AWeniqA/2RaUS
5QtNwIH+qGg25wOJMMe9x05N68SlLawrcxQuJ5t35sp26Ac6jjmnHHapdTR1snu5
QXrPMiMzopjITQ4DVRSDvNv/e07ZKAsDmzr1FjCz+2T25APDoxCdytBi8it+kpOP
DtM0iJ7IAkbMlFQRuZ+Nxzw3xiJ1vov0aK8ik20UpALWynWQ5/YpkaMDuoL3VCEV
Bkd4dvgRyoQ9JQpopTpNOXeUIFDv4+JQuO3K8GByw8Y1cKJJyDGYhMZbxr20QkNs
vjH80PD5O5tb3Bo60oUlnArh6A4UxoX7euVfyOGoekatGaS6KAqBcvmHTezSRFEr
BCy2/5D+0SpmMjy/XaVh22AHkd9JjeWPSHcXeGy2L2BwTwlR+IKVc84uacyAKJy4
RdUm9yM+7q0HQ6H/jGHrA9vmk8oCVpZQDCuclra0z1FNUMzftP8Nj4q3q8DA4tJp
GYGfQyENspfkEIlhDtyfm1TqLwBTA6LxLUCkzMWS13dF05ZUjD3gEO77Oq28a1L0
VNqOD5ECllqlv5wG2Cjhba2bRA/MroHOGicB8xeuamlxguD5koK2iwPur6fAr4lz
at+IkG8gpCAh0xDHWAq40BIg7UbyhMuWCLN7ABg6T/VffGRTznTcBrk/hOefDOU3
BzdgMhjsUv1YPAf4+RTS+RHDNyDhp3Bq99mhEWGvtjz9cHfS2cNWWDXkV1UXS18O
AZHzW4Ke69xGaW+M0ri1XplnupRpvmIuYoTxQ1WKVD3M44yH1j5GiczdhXg6lsTP
4vWLlajMsF8KsMvaNVGpPFaRmMHJahy7/zSI57lMhFhTL8AEzMXUQ39Pbjf8cKI3
9LIYCpnnxGJpl+1pRU0sdmS/z11hF1FVXwgkxXwtmhQr2jvw8hMB4TtNDB5sxI7F
hy+2KzFxAULveP9tIDAyWPj7duqvd0UiWlCx/MzwZW151Jltf83GmI38hXKmHOJJ
EzELSjP/qrS/ql6Nctt1K3qQTtHsfufT4upcBSQlURjzyOWSrYkUaLqCsOFFW7Zx
CmJ6WCKuoI7b5Rol7fi9DAdohQdgy3EgqN5WyVZXVZYh3v1ezUtCK62f3AMxfhU3
TNHrW/YXuYkQ/i74uhQuvMUc9gzyd0HFuktFkBbEQ42NG+u5PS826X4/hMrOzX7n
vE5VtGuqSdz5njM/gWP9O4v/w0uSxoH9oQJXzOmX0vRgKb8jnAB+W1AjPJCbS/zt
J9JU4hh29XgoYCf5nI+bmX+36IbYIT/u7OpRNT37lBNoVbeTsn1cHdhXWmEU/GYp
EQaimu96Xp/LwKVbWv0EKx93t/XGMTkMNu73xBPu6iLyLctYXcCYhNKvJNjbx/AT
XPST6ISuGgp74ytWAk0VO45QRJwFTXgjAlEP03FW/okX5v1THX9d+0FfB33vwbM1
S6XBRUVvR9GGjnllCSekL5RgT2yMwTNN06pm8+YUHbLdwgwK+2zM01jdXezlnLU9
WdXB3ie9PzVX3ljisKY4RNDX61ZqT7ZXx/KNH/t7sE16QjhW73lxKnOE+f8n3YUV
M8akBhgt340odoml6W6udxFCgRdkivRSnHqCa1leF88sxLgnS1b8qM2XwMPEhDCC
iJZyMauMzVHfPoTc8MLwIdo4u7blBuyrfa7MZmhcWeaAsyIdxbOOfdmQCx6Lyuzt
X4l3IareF0OM03bZaRtS0iQWX/DH/VGs/aszoFxitzqc5LPeYVfJtKNNmcXb8rpw
al7jKsm3nCl/uamdk5GQ0pCk6RMnNcDLk008FOjF19ALbGHEjsG3YoXDLZkyO7mI
uz28Fy5eS6umPcxT0TB41dsoVhKgKZLiKRMVbFsHAzEF55NPq/EsrGXmxjiNKpzG
hyPdnnuO7wXhDxq4cYJC1eB7L2xFmeMMJCVJmoNP+8aRxBCu+5A+modkYsKbEbIS
frezTVQt2AHqmju0AzSapKqAqYX8MO8su0dT9rc/4TIvyYPhUgQmuj0NU1DdLBiu
Ms6CuGTVLa2HoqcSH+Be+Q4H+mWAFPv1Zg9/uiTUAtiZ2O5QXxjZ6vH/PW0t77Ua
M2egZYBGAWZB75LOKMKvgP3nM+XU1B+kdCZI6ffFQZCHuoUAjhn5mXHQXpioxVKN
wdkqyhBCNaOiGxwt1FJi6LnaPS868FDZy0urPFKTWdhVvOb2LHMJEZAwGUwTvIqC
ZxZBHKNRUdOMoquLBk0yTbjxWgv1BgYflcaN/ASszeD6970jy4KKltc+azNKa9jT
Qp/oHM/7GujMBUSOGcFKxprx3uXH9pdPAhnmCLPV5za6tcgkPclPe7uVaEd1qV1A
a1YzcuCt5AtpiKJjlC/ekCSycfGygqHQCZV9MOtOvojD+aUXAtnvEiUYgtU0Utk0
yXZVrBj7tw/mCJSHbp1cxPJXhsxBnBubzdLuft5S4nkD5S6tkDx3MXDJ0rLu6vjc
wxVjfH1WYpFM63LY9U3jFkniEzQ5pWm3lPlzHZCunro1fakMpJi6HnQ2PxKbO7pV
hCJSa8ZJD3hmjUZ15qbfVB0ldkBg0+DtHrBVC8L51lgtI65cIaWCsKLOFTXfefz2
D085NwFAcBnZsi6SSePU2rMlv/FCcp1XM/88QPani+ooILjL8LJhXv+ZGnnr9JGJ
h+890JWoydaYNyoUKflQYM8REDC2AcQK8wyVpUlhU7QVsRsY+aGtNADPz6maQHty
JmH6TI7m/mP++/Wla7yoppsnywIk4ycJXKfDEiS9NaSEg1NIn0bnWtHMEBeQixTF
ekvQfC9x1mNUg/pF6lBqCyJv0o49tcnbluwYMXh+AzDGNC5/pHcMYW3V7AvKAnO3
tRcB6syf5Szn1EVBHwwmwGkF/gIqptVbM1snLI23tTKIK9CCHsNDfHx+Bwg4E8uB
wmLHUMd4LesPePGhLJo2w8QgRfWMdHW3J0g0/vq4gSq489PJvmRebsy5nKrtIZwu
lhBUaWrPwXllV6vG7UagQ1T69yKXficfFJk92A/c7HVKgAOWXYho5sDL7HIbp7o2
fSNahJjeg3O6vXZ0a6iE7KriAlAP+uM4MNy4s/JFfc4D8D5EemlXXCa3HPRr+XT8
qSKTNkm8OtjMjYscnDkVCHderTjLSx2KHIzhzjhnbZGn2OWZwC5i8JBIJEmd6Iim
mhZSJReLhJaE0hrHzOP3OKErlRa+28PHmtLKeYul8MVO4hafcPI6bXgEfC7W6wEY
E3hCke6BaIfjYV3jzU+UD7qGNbgafUGw2b3i5Kq+y/mYOpiZbm/NbTEIhIc4gKqF
sUXbPxenFbFJFyBYOnWzuZgUWiLf4vl1VD1npAXFG40vrIu9Jb+WMMukV05DkM4Y
QZn5sAPXzYRwRIWuTMZLHn+jmmWa3cLhkkB4q/dm0iO9GOdzmGOWObq16xy4a7UU
00FLtVbE/D0uIF6cpMb2oT1TwKhnrEPeSUpNA8UloBB8pQEVfH1q0L+CF1WbIc1E
CTeZmJJ0VqEjkBpB+t/VYFzb61LLk3K2x7JfHFDEGMwUOIHipwF3BOhpAG4r32Vg
mo4mdgtelJn9lLw5a1lzU+NOsxF2ts+PAWYHgdJw2qFSiDlR9wwSK/tgjFzetfyO
A2qPL+xRsAM4eUzkAZc3E2nw1o+YEQqR0sfdHHGPqQ1+b01wKGSJEp7abhkydjIY
psHq03dREZZ4Sel/DaIoflFiyB+tFGxDMigkHmXTpSPy6FHuSdNDAQLKA8CW8+qv
Kmo95WtE/K5wBL6G/yxBTA5CzXP1WlnCygD/KR6K1kWmi1prbr8ONgdB44mlyOmA
83tzKSrerY8QDSVxMYxS5IXyLSHtf1Af8CRvCornEbgc8+QYe5Tvu4ShUAy1JHqd
aF0WDkE+Isysg4NP8K9ph5tg50qaZfWRWcs4S79by/HbFf4RaMsr9nSY7cnBrcDM
9430bcOI7JmLlq3f4Jj1oAnfEP/E6BItDlVXQauN229yuIUnkegdJhD6bYL6dQji
jtIawBYii32sjYCMb308xcEGUr5hlGHhcywCgaj1vNP7vrOxIj+0b/ovLW17d5lc
Kl4GmoqsEvG8T1uF6YU9xRIXIIwrgFirSqFWYlJRZzgziDa2rG6OPfRAFAm1SXqP
/Z2TkXj6cXN8/QWYxmxtKqpi2uh7nhqLgFGlHJeoSFk2CqRmENHVT4y31PZj4SS0
/4LtSmlw5ydnPkRNByCofNbP15Wdjz7/a1rccndiBzFlyA9hMzy+BttTjO9/DhyA
9AAHMCyxM4JVdRZ3xvYzZB3FxkIwCoSTqwOEDUGUNofXJ0djqaf4CqTPzJRe0p72
fe5jiPr9Mw07oP1x3DSZ9FKG6E3K2mAtMNrzln5F27E5LniyWEoqh+NXpGJV7YKo
OKivKIV2ZaSwwnfHxoopZo/YvCJQwBJn931nV8Pn6eNMuqqOai1fssAmtGimismY
lIHS0rS8UljAJ4nPFprwlFpXDlTBLlBDiY5t95wxUzxtMj35+Hr+kKBef6Aodgnx
3yk1e8VMSXP32enmbYjR/57tsLRKDQPhL2JHZTiTMsmR0v+iiVtaleQKVPtlcx7p
JoWOq/mQOGjHjN+cgZFJ29rKJdwzZfVZG/xChRLh+0v+t9gOKqy9gC29KaQHvIxf
RnQDClipi9e2+UQJbHllOzeYWLGbGg9opNjYh8Wpn/Kl+r67d1IcnjsNiCDLXyjB
tINZ98APG3N/j5PugB0ky3mElLLLc/Ii5HBoa7Beu2jsgrCVmzkDjFGTu0cffV/E
T6OHe42kGptWZVOIMuXr/26KknSeAjDgUbDKGbDBvvQ+lToNhz6JsSXFxmCjmnVz
Z2FXxIbN7k8sZneoelTXjrZ5bXejkDjBF3I/FCbkKojsINNMl5Ys4d/0Ssm0C03k
HEJxZEWk5ddRcfRxQAt98CNJwZs15HNM34qecvWWfFunXRrQdF4oepGkMEjUCKrN
N3slxwC19uR/QEegO5BR+rocc9kmsdAY/5S3zbs/CC7/KHSeU0ovPmAwRn/YMu80
R23/hJuETwHaWFAMh169GSjDGRKm9gqZOxnZ+EU9q0722wBKzdZucDT5acVzWIET
hwhbz4FeR9Stk5dcmgx2neFgwPpQGkmr5PIpaQuTpPMdQtktSx6RnW/VPB1OCq9b
WQ5utXw0bWbs+sOTimgcksQL9JbPfd4NVSHOm75k5cRy/LCVGQ1d+25nfVVjbZ5E
qmy8YTaM9eAT+aMoW4Oc2/7GryCguYw9BZoOane4TQLrh5K0Mukm/eQWf+0vC7ar
fQF7fu1wPKAK0PInQdumfVuIQN2g2zJ6uTJQuCpkf6Jm60baYC+iWqL/tL94SZ3f
PWOMwB5mcXRU08hpMLGLH1ypkjfj1C1uVsgbUW3bh1a2Q5a3ve0jUjUzJggpUwW7
B+Jvf019+1KdJMRFSyT2XVbRZz8w7mAwPZm6n2mwgMS3DKKxwf+EEPWGNu4oNohf
miN5gQQRgR/gjKdhjGd5ept5Ywrdvi8rXl3nyZ2asAvOBW3tkRzUcxwvpUlfvthI
c2ScLbJ3YYTh4KEV2qTNQ7clNyQkTRtmDUiacSB6HERlc+iHb7AtyGbuAIxsbhYF
06L9DMxsdiEv1+lya0qwqFYNmPFwjWc2THKo3dG89ipAIOp7i8r9s5pB2ucZLI4J
UL51tgVWnfYTTomlSZ1A1zne1XryrMgRspulspJQ944wgTFPkf5cS0elBMgv1+hx
V7SEgkqlGvbUD8Np764IeAlUm4F26MZ+R3rVlJkir41RNxqH5V5wsfvsCPdC/gC3
+7aghIvFdTXLv/wuqYTa5CriuHPz80YtfnRh0uDSGrFnVTUFWk0y5Kz0Ec5RdIer
LPjrN8vqLY/pRNBb9SlOopV8RDc5RyTPY5hyfArKB0ZIE+iq2Q01z+DVJmpHZ5VX
LQiC0HOO9Zx2F69uWvpv6kMFDX6nldZVYtNq/551+7O4I65Wh5vTp1HazOUoB3k7
m/tQ2DM3/5zhKH41raVWuz/23KQm1aJM5tXsp1CpE56yJe3oEDUEH//S6kuVXxlH
H0DnDwuR5kB2czYWUlCQ6qoQyMeXTwjJjjQXCTL++3Q05LEsIbGLEM7RHJmGm1l3
N3C4j8AJsV+kwlEdDvU95eraitPPmQDqwdIKW775j3OXIBSx/JiR7mzgzOdhh8Ww
HrZHYW4oJjX5KUafwuhzXZLBEmjWG4wVD/d7r1rswQ2gXDc6IJcyR2K3QawrR68w
FRCFTgW5bjD8zf4eI9Q+t1/w+qk1B9YJCSHgImHfPKGNqWeNZ+7UNKaU3WWdonjM
7KfirIKHKRMq4k6//LpPLmy0OKcKgQr1jAdQZWzn8DzQHyWiJ0YE5Y8dYzVUmVtr
wT5ck8n+C7nk6mrFdnW11L31YXUosWp+eiRUWiY8vQDZox7H1Imw2bMqgJ+/WPft
MnM7N6+HdIFmd5pAtUWgw6pGCtbDm5QVcdjxp42hmWrKJpHRWUh2vl9O9jX26jR0
XGwZ9hNa4Q8yksEM8REMEnSg9GdPQLS54gG/VI5rMc9+DPKqVi/FauA/Kubv2UHi
ezPhK4Xm6ssidZILCHLYO0qBf32oPpeLSukqy1678uZ1LuE6rp4lqYsPeM1+Gbs0
2+j/H/IwYwov871n8Nh4mv/nNU2qz9jVl3dO99QDySuIvb0pD9Ul2ZVZGvwLbbbs
NpatHcSRDW+h9BIDM3R4fbQBlR6P0msk+qMhDEQUDLcS200w0H2gzEzrt1rWvPcI
iC1FA0mGswK1dj0Pi6sxs/tHrC2HkIIV7WVBbXqQG7amj2E6gPBPXfrQO2mimKje
3qjdw+U5sEggvjh9lKs+TrRRQHoi++FFi8aTACvNh5YBSmDa+UdXuWftVYsv+O7d
RBT7i40HOZANeRNeERXuPw/rLaIX6SuCsaCYEQ9bTEQpM2XOhRkmVboMdK2LkRcv
2oMp/5PwsYumHWgWWS81vpGGzndsKANktvHiUp1lN2W1WTB7DmUDI1XY+P6oKNQM
ZT7B96iXfJexKsBNB10YJuVlg24IN//PF5ZMLFxIPhqr0DZ/WB6c9t3eJu6+Y1UK
vhARXJaxTmXRp4nbBBcctdGzV/RF7409l5LH3wYQLwpJOst54rpp5GrvIjIab48q
45Ch9bczLvONsMdRqKLWing1p2NJyWuec5BfboxgnJQBSVIn6W3GE77UnhAOfyN1
8SjzhPsgbNAxhUshd+l/sZL7P2DguXIqMjTTSOBdHqgvrpC+n5ExIOFyWV/F0hxC
wjokNN9EqdRtaVoY3EyzPIGw1r/CrDPl1gU2GsDLN/Zk7YkrUBGUj1Svd+rsPSha
N743vg7y2/nBJR3/kK+yFrLu2rz6YK+W45eV2lnNIZRqd65CJDmXvJ0gUN9yykKk
sTpkTrAAAWAUNlpS4Qnkrv5qQDgWo9TTv6WrB8m8Y7HHQCOKrvLy7pwLjovb4VzW
+LXvixbeyWkKUhiiRC0RQrea0Jom4+Pslmr1/0vsqdogMoAU3gmoI3oOdl2V9cAu
6a46j3WBrFT520JSUj4lNpUB9hJ8ElwkVQF18CDcxOqkBaDcsHFckLxWHCkx39DK
zUC0qkjFCld/y3WBHyc39Nqa9B3YQRm7LrzZ36ZgHRjxW/d6BUplJVu8pbZKEF4x
o9jhBcqYEgDliWgcxdLszAG/FbX9ctlLJ2Yh5pePQNdZ2H87JBfFBueBU4vcrWpw
mONtF1xKEHGQ3Hf6ZA0UfeXrwDUB9ungizHWR2ZE8x84jvYxIdKUKAJvM9LskKID
dNgqYMVrskYG8y7LE6FRW050qOF2+vt2yVxpRIX5iLMmTa0Qcwi+4SRta/fLenZR
moAeWwwxQnPx7D/w1IIXAGnYffXPYkyqFmUHPm0mFFh6rhkWAFkM8LfSqrAhAq5O
I3tePjCp7+5vTpr7NzeNKkTstPaAGPa8V2FwOACB9jMWLbkdTCX+LaX7u1+LiLz2
8pbHfQc77mSNbLs8zDpJ99YW3v2wfATN/y4w2CnSbJL6PUZDCgua7LWizQKOfyNS
tbhCXHCaJC/pR2L3RuZPbG58ViSUaTp/fZqayMH4HHs9mLwNrLWcp5A/R5UXPWPi
P8odlC+iDLvR6HL408erarOnuB6rDcWlGQ33nV4krGrN45Uz3glzQlb06C5TWhJQ
BhK+GYbWdWuw9HNDWFeWOPTaXLKjB1ZCm2IJSppHE2ld0sYYVIOLprZ5w4QU1Xeh
ffT0cwv8qthFChKAY6M6avgHNi09TYitSE07Aootpf6TEnPcNhK6aY0eJ6XMOKwK
GNdlhbkGuS02s0rLcsccYoexdgFNj1lKpnPq3HehsxMFE6g8xQD1qY1pS7SStT53
ugNMfR9JcCHPaYTYP1ZGHc/2Hya/IfqVYXLVo8ttOfnHdMt4CMNXL6wn1TxFVCBs
0rQ8o1FYNqaZ/VgiGUlULzoDxvliqHL2uIEzaPowlXzmhvAR/+9qjxAQHU3SCEhs
nVfk/Tbd539a+8q9BL+IWKKNP7oXjeT30CHxcaglnaVuXskpCYucLLUhXfIVBzok
w9wN74VRZFqVqgGnYSYMFujXGi4HNIjMwhO7kvwS3pC0ag5UgOaDhahGvrCBAF2M
VGcDxjV+y7MWz70zRZUKjdrhlLBDcainfijrHaCJsC4dGc1cMqDFzUFKruK022Ce
tcoV3voB866QbXReYZ1KD+yapSV/ya4dZcNVGDzGIZYeX2/cwdHmoSUY+9G3jZr7
Jg2oX6BxczPw5rj5dEoQo4RlpQ8hHa0ebgESbM/ml2xIjDQdjAHPcwST57apspms
jBj4JhyrB1XwrWlJ/mnrD0Zpp7+gIjTyAU1NK+MRnvg9h/7exvKfJsj8iEMYXM31
s0J31TUXvzRuOm/muAY8TziSRlusJt7jDWYn0BOBuA6Q49GdZkZtLs+BFdixLYWp
GE1YjZ9pIykTVCFvYwekJWYw/Qa/qxhmVZcg7O6ifKwMhiQtSUTpJO9Hz6xGAfe0
yvI/4KJS7DzDh/YlFQQCL8XpDabHlKQIbQOSkspQEC/CYJy0YMJUiMKcbqhOd3+C
A8DXRaDebBYhTbpnQjNg4kU4aU/hQliGo0ZtrM9q81JPNJ4LoT3/xrkd+YYpFkFd
cbqEQoU1vZNY0+G5DK1SAHCOeYo7IuOSkj+te4/cHpnhmETv3cUe88z0y/eL+nXj
9IXfIc6E4xv9KjMU6gIYYnGbmyeRpx617Wnwteazn1MMePgc18IeJ2KMSt3v8q/0
NN1KeAWvSkic2uoCwZ86UZHGlngUKhm1o5uanZdz70mdaFvDdT+zuWYU4ZIBIBc5
DLQqyrtEZeOW6i59JTmfPn30gDzf2CP+vbJ2nSPTk4sB+aQpl1tbjQ3xZZnpJipa
2d5G/kh05+WNkQnkdXAbk1YmLwA7k7HR+2fWKtTqcQtdfZ7Dhi+QQL5sIGd+6Hg0
g/ASF2aYkMA7XRhtUwfkiyHrZk+/YiKOXVzw2Fj+3U1CFDecyZR0s6XYs0Et1VAT
f+tMVimHpRSwo2rdEyamDKaFsiA2rS/FK2KkhfkeNslurSCrZX/U2RqGt8DCMm3X
2tjcXoXS8hb8PTJ2SbE03ZZUZuDUbKVwculkSZluNwmij5vNj5QDIHQWwcT3uMYt
htKtdBGvoUCqW1VSulr2s0Pxs4ULISj6jnVQwdVOLl1hSzR80Ev/ufYJrI6nmIK6
NvXsTPRMonyvI9CySGSZ9sRXpNHANty/TtRJww6KL54JbEuOXQ0Dzl9EGSUwomlv
/y6/ngjiWfqWdULDLT27XDIyz4YGj6Cq5fEyIbgzBP5VluTQtUSDVBiLf1pixVgn
pRPrOuSP2vyZv+fapPWL8UW0IYcSQ6cXvIo0wmibyuhe0pNqNbcb0E0hmt0oqy73
ZHcndwjq57blJKFHO2kmpp+cx78F5/X/0ApkMZGkfULGBy/jBAMfh/aHvCE/UfIo
bAd6ZOvRwR2SBRkG0NEdVqCO5ObvfdnUbU2hjFtmEaoXrZvKVzVF5KV4v61h8+qh
nzuuoAq9yeN6RY4hD2mL9qU6/D9SIQSV6SyYgFYjAQo0YJvzoEuorMcG9ufEpK0h
gsPCXVBGMlCmp1AIWm5ZMSdwm55daLWUsUj0gF0G4HJAMQnOYc90aZD3dHW7rf3Y
TcdGCjigW/O+gdFk3DlVl2DpqTAfScgPcPHQB3mC0yLPXjrVXLKafHPIJwT3Lyru
eyLWQot1gp2MKM/SzfMAy7Nqpj1uGhJoqFxva6M/o49agwUaWBLfEGCF0YUGf4t4
e2gQbePvd0l3IJGjsCGq0qOeLN6sjn1ypoII7eNAivy+v0hD++4kEYcMl4MVmDG3
NMCwwxfAYUIi/6zYgq/SAHJX5IO8oQQoQjN4kjAG05OHonA5rf5vI54Woc5OdIVM
xnfBcX2Xxxm22Hp9s0WFRLSE9zwDLlb/VcOG7X3bBsS7XozGnS2d26e3WNPkz4HX
0rV1jRK+9UwG02uqKf+NkKtG9v7jm+GFfGEtsVyUUWfem5zAMqZk2LywC5w7sJ0w
3ggPAAIO1MjXf4qerAMUH8jJD+F+axmCqime6uUawcWBovXha3e28WLFFdI70s3I
izEMbsP1Bru2V881jQpCUV/Rv3hMLZ3aDKIbSb/UGnucCPx3VT0O6AWejm1imPAa
peuxhe8OLo2NiKWN70EEbhitk3cKf+wAKbZ+ufuAMiu5R6QeO55dBXCjsMK//eyo
LIvIogn07mbXWLqKWBKU01iAuQlJczo5DhJz2Wek7V/8DbwV7Ey5+xnJvID5wjMu
ZY2WXpiemgZ7DfC0Ritk7OnMdQi2uwgAGUcIN0avC9KY3egN4YYgIbj0kMwMrEUz
dmNfbybURU9QNdVUm1+6c7aU5lqf+Vw2PsONA6gQZmIYujY1wxomVSMOSvR5ETnp
JmLgJsDhjSGZoQZI1QhQ0PrGV9O7DYaKekfQeyJOJm5TkVwDDIzHjEPvpM7c+Uk9
d22ktnCtwtTWoQ4ClB4KJFe2A4OPCGWNzxa6/VYmQ01M6eNJURdGwTR7rDVCZUgD
3ww5xie9U722PgsZmfoOXutr6aS31l2WEMG0j42VKKt1W1VKmyYAReYHjjZmYsEL
Db/ABHHPQ0MaoTCt2EKkxvOSuELGHK0JPuzCINs4Es66icEYbf1wssmp4B3AkJ4z
T1z7MdCOLrpb27T364fiHJ42HIDpXyROwtDNwjC31Pi1JxWTaL13hjjqaRAamkN6
BRbcexVve/MfoMBVhU1gF99S1bM6xJoIwLhK+QNHUKYpCVeDVwMjJwEGWa4IOe3Q
LbMuDK7wpEgqmraPOba+qRU9ID2tEWtys71drwrLBXa3k7ZpriTS/OTAry2WtF0p
5op8W0BAy/Q+QRycaPWTGkSYHJP8wUHPunalmCKltfVnL4xyclsjfJrWXw8IAM3x
YwSt+GfG61h1bDpzBJV/vCB9SFyaMH5/WNeF9aFbzb1JPwPnNOmiEzC/fmdUP43E
iidKzzj47+sFLv4E1mK9m8VseLPbCrAWZCOVSQIusfcttqtxwozOa+XjIEDcANXc
t7BSxULiUMkCyDoEmSn/Q3yO4hezBvSRICNzUnegUeWub95SjwNqEG4+dmFIxQJi
ndYg5JkTehFVx4KaXZhl83boexONnHgPTHUph5ACr8Iip0Ng6kY9W8wDt/H6SStK
eVOnHLE8CKd1vFe8cKmu5lxaGSw6zm1arH1CNyz2sdl24HB1I5uO4fqsPnLB+S4m
w2LpD0JqqtVfICn+UsNtVFCGumII2Kb2oGIQ6ynlDU9mol2KMruLvh5OIpLh2cYP
9E3OU7L2vbMtjqM9YK3orXSxCzv9mbRQiEDotP7WUMEy86rFiHzsgUMW6wHYjzmn
fxheLu2+cH4je0eV1hJs8mEWKDxnFX/eymlUu19ntTtva5i/UNZhE4uk+OpSzPSa
wNtuMbJJL2qWuytWo9jwh+EKH809Iyt9L5hXHpxe+24UeVYfv8Z0zxLNpgABMeMl
K2M3Jw9tjhiNyoLRDVpGXR4HswLz5fAvgYnO7+W4XU+4py+O8rSEyoy3UVm2DEzJ
C722G0NKNc0XjSLWHEOQeE0S5Q+fwufaxH/lB2MtCkPhD0z61sW9oK8WSuy46/Z+
KTdMwQYSugqWbRO8886yjHaGK8OBlD0xEPbcgmirJWYX7xxyer/N/932DANaUXtX
T4c0ri1HRK2b03gvnwjmQ3d8d0FIDNVHIBp/iurghjHv35kIOwNqusZ1cpz710OR
1rrLUEHhqIqp9cqnXlrMs9gkhcRXZ32zS/PdrHec4S9jsBisQKUTnDVFOMrgbbtM
PgauWHSVNIhWSPHpCwdhFSvud0BRr/xml1e+J9gKxRFaXV5YfE+N3SXvG6e3rc4a
rSNIpjAqWymyB4y+oyNv9u/9qdNJAAAni03Ov9omQF5VLm19OmbsaCA+WKB7rd1J
BYR768rpePFkH9kck65Ksq2O9imtEVATH3y+YjMHODM0Wi8mFsbIjReWZ1Lk2DNm
sii9BuY1TK3C4cmlrMP6xOXrOfeTOZaOTX35+BMmJPFG6X1TnllJbgAk+dFt4SkY
bq7SOVBmafWJ7JA1srqweplEoUyoF6LbwzWIewPAtyr9gqTsIlm8CALXzT4OPrAc
hr+6So/nXO7WWopJ5SitjL9khiUkriH1jZPrQ2g/aCxnZy6BB8LbFmjouMiihqJ6
HvPhEynb2g8OZEmAPDk+HAnYh/pim12bBl8yYh3QbwyAJicmHLdqevNkAdNMhLph
QbY9DrX6nV7uILJnveZnjZvwyJg4qyisXx7Hc0o1O/XLUiEe6PPvcULKKbfnpBeI
445gHC+tN1WrO+V8i4Owdew9/mvqu0GQktYbGcz2oe6y6JkVow+qyIF4YXwVph+O
e7WMqEfv2RkDWOecV6fHJm/L10VulOSqP+HjZXzpnJCg+W/K9rPRkStqLckBIt6J
q5Gizx3aKUBbi2gH2cqTkvmTdZXQbkxgwrZCR1dwvanVVUsRuaimISZzVD3/tENL
lRGBlmNG5nN7ptfzh5EwhBU4x1cgUPxoZjlVLOk8G7sBOlzVRWCRI9+rI3AH+tEL
majDuJvtPQHSusrbL1On/tV4gBrCBaYadIxx02c3BKK669gJLnh8SDtFzQjnTJm7
CNoBe/NPqfnDsBBYhgL/ZRB7ucBm1UcFcVvapUTpEhQlPoMGOqirjw93lb3a6uSH
P1e2QHQtU5ZooSOgiyCAKtL4xIVZSlFXR8+ip00iJUwXWCKDW27iSTBqGKh249l0
2AKVQCs7sDzj/G2Kpljzjsu1b+vE2uTQ39shqHGpPwYLfE+vPfTimYvi39pVwH0/
VEdOd50u4ytUTLipwQhqw63JNQKUMen0dPzViWrKVYEVQE1FWCttmMSQ8GEY3VcE
HU4FvymSV3njlXAceznOIhtslt+j+xpPZP602sqSkvaMxlVCU4RwzbVidh5dqVAa
4FBXQ6wlWINoq5okoSbqEzTWDwj3/LOke6uD/r+ymnoZ2OTVce5iV8EArUlw73Vl
drummL4uRmV5hhQSRN5/a6LKECkoTYTReDJPgIrm+hBPFNDOfQl5TEMjE6lfRzt0
lt4BS1kfoaB97LBg3OFHhEenmurX3j9j8zQ5eRBwfr4OkjruocvhVsMqNify8AdW
IiMbd/XO/Ao8NoEoSbPeKMhn3nGAdcwThIn7PM2qMlRZ2A4J19aVvKjiePPwADd8
aWj1BkQJSbIO9QObldrZo1fmN6BiUMHiL/WZq6xeFW04xubKVwA9H9mSLspv45SG
/YGkzFdsvmK4QVVeqOBk6Rjo3TkD32Q3xiB7UN3vJdhpWelsPiGXmHPlkGrDa9JY
v7BgcPJA6+peTbenIyTM/XozM0Rg9gJZaDJoea1RHmhZQ876N9RZNj6SQZiTaaf9
3wy7C5/rNpHFSefuD3DOjBXxuvbMNXCY8ObbvAZSCnqNugJDyKq7ZRzA5G7ijKvs
S6XOZBhipMPcmYOLXe4HVYSAyvBWZ2gWAK6MjhcHTEhW0Efexux57xRRgi9n3gmk
NUKpz9w1JEqNOaB5Oi2Zi3l95I/dTtZQOzO08qcowJ8Wj1lip/Vzx/ApPVI6BjJ5
KZ/sxEXqpKXxMlFa5KuwA/Em6HjfIt/t8Be5/bJTO/cBo1QVu/JXehmNWuDNJyY1
BcFPCkrQuInhiqCgCsLG7qUlpdlMpeBmZkHxGjcovo9A/BCHtlIf3Ve/e6x41Lof
IqsjB9/R2z3lFi3BmBXEe1HdmJyfqPsb22lmkhGStgpcu6dBHvM5oiJSjgVqiM8y
0kxo8VfdFLdgCp8D5BTmfIHOsGP0qzzIFnQyJSI2yqL9nNzCogX7HLoaXwvnYZ42
5acBsDIYr+rVQOCB4DAyv/cskHk2noNbMXg9MgV5aD/mF6U+7oCKDCz5DVpd+YgG
KRlb2iv2zGW99hxO5PwBHkeW/p6W/TSKHB2orrKBIpBtdTkXzy6TTwZ6wmm47svW
25jiYrTEFm9wPNOmZ4PjKlnF9/NBjClJPMi6KbSvsgJZf05uj0zret+QZzir47rA
LXFmqBOzkSpGoEIkWS0TztCh1Xv44QTyHhsS56eQ4CYjiYm5pgqlMe/B2JIH8MyH
CzhzTGPfKNQGr6Iq5tW/0As5769ftxdAk6uRVati6sB/doP68xlleaCyIXrb5st0
fMmEG0QoZ2KZbsJP4RlzpleP20Ptpw1qoZp1LKDknoV7DcEgxJqrZzEcHgs0Rzbk
NA+9hcR0U5XZq/2i8vxtcPznXfLv+y0t0JhdF7cGwmUU8xVGZwfVkQYjh5BKbfLe
p2pgpADx+2CLM05JH/s9d/jeCzZLO/mmov9xKbS7IDFyBAGQuEEQ0ZEyt2OKP+yI
Mn68Jl34+n++wwiGQRRFXPSNb8yq1OxvZSxGF+w2pyS7pyYzUluXHwviILWVEM83
GrNQtepDtpiusiCue3y0Q7FsLf1SLEGGeHx+lKL8q0eB/mcvpMwiqOjgDjQB7Nir
ydlONOH0niV1uZzjHlKNRbuLQ0g7Y7qWadaih2SzGWfH54/4D/TTpos5d5fS0yLe
M6SM586kQSF+Qq98Wam4/gyp736mn0qOI0we4DvqbnDjSr+LO0DVzkFsUpznfn3R
urMdT+wcG1yh04dCWVEtPKCX7vxSIirAwIk64Boo1c0HwWQ+ewORll9RbTmjIIiJ
OSm4R8EWEVooxLyZyA+6KRfthZHk20b6tX0DBZd1Bj93IyqmHLlD5X5/KlRhYKAg
ZVyJ9DFDkdSH5CvH3NIQALOxXfSDhMZ8X0a64Slg2nqQN36a0RQnb9neAlg+srTs
q/b6pClGr8L5m2+ky80Nc9abITtfw0toSyivotQTklBexr1U6M99hnwtDcKYAXYz
QKq4KRCA0/mV2GAYo5+VbB3gSu+gYZEZ7MwCIKQ8n+XjRM74eXWoseiezzBliRLz
/mHBQP08CxD5PE2weoehdgdDHVaha5sKQ5rPedPvtw7jMEzHlJo7NK62hdCh7rIn
mDSYA5+u6JiSxi9rQ5aYN9U9dENr0xhqG92IGz635UoHIiV9lKnNs9UNJM3CYBcM
oRAgHEaL09q8w9SN058OZVB9Z+ut1bKCbY7luk9gAhS7MXalFNItLdNrMFN0Jxz4
PYTn0sre8BA9JLYm4MoHFUaBRD8aezzhDoblUb9Js+gqc+3pQo+aaUt89/LyTqso
dUf8zidqYZEzarFFxGL6TNfx78s7JvHi/GsyV7MBCKRxaJnWvk7eQqNk6o47K4Rt
iuSeOoPZSgYKGcoEXmh6e1NNteH74sdVhgK02NljIKM71Vy4j8Vl5hRNDhIVmb70
hBkChhjqEttgVzhHSnJxr6L0hX8CasdLkgXXDHFWKJ18fnbKk919ZPo8CZFSLZon
G6eC7HOZEnCW5WooGUhS6vxoSLfeWhi6UyBQwu+mzot1NUnWhhguA89wfr/oJqaF
HJdlTVCSavYiMkud8I8tpJ7WtzU5GHH+07wzjfUkawgcjA42s/1ct0KYUa7r7ZlF
sJOCDwTftEP73Bc5qCxD3cyOkvVQa65Kx517CsUT3hQ/gTH1JOHE+ugyUij2bHMh
pQbWaLTMn4AmUc4YMv52kNDWF4qR9DvInpg5C2x037AF2pay0gdh71Pharv8nUoh
jq5vQbreO3qIOSbYOP+IDqB4aq+1OfcSD8amH4zjQxtltG74bReqx/e7rrgVo/3n
emf6rl1BK9TngqA8VkiobE0XWcmOZ3wCOuey+jWKdSqlJQiKbaGtELONRdoESm/Z
7gdag+Qh9htLPCvkeUeRlbrRPt9Fn0seI4ly5jaCs3YsydmQ7KF8GClAPyPlGIlg
mCtMfdZq9RuvGiImUN9SvNovCBmBkVi06GpOY0DMeNamLh5Y7shd1zSzCufkXZ6i
3Ne45cwd5fOajoDuRqa9sUUBmx35kdgHwIbIV6ijfjuym4s7VisSCYgTK6QlqgS8
X1ImMWA2XOkPkgM9F48xhC+98f+IOfiTKVV1Z+t7sqdZKZH4KwylHvmuJliT+b7C
dLpn3L3iftwAYADHtzhAWDTQ6C2PhBJdxARpAU+0VUz2Wa8UIjyDENXkKd8ZoleA
racLxSzlE1vfRA/eRZqPYyaIUn3kSyYerd/6z90cSc/SonrV0o2NLHB3lQfSqcQ6
UqGk1nqRMieMe0tUNGpShX2ahTLJhY4YZ/8EyP4zFxYSOTBj+dsos7mR66wTCMuM
8XWtAC8ITiOQGmZhGchA6ZIjwgIJyaGUP7B56aSEVY7WVY5JqZanijAqEOYqllE/
y/IOThUW6ls7iip8Ylya7y9McgAqHYiYQvJGLACkAh+8uQBTbl93+Whd326AC4M/
Ud+82Gn84kKs5o3h8U2Oq6Px0YfJrUI2sHT+96WK6Rv/8zqzq1Xmf/aiC+P5AC0C
t0z40nzBXgeKrLqDzNoOf7tpG5KAoIbgB6Z0xfMmB0wTZo4cx+HuBTtBqzITeEzl
ABqep4qlr6ACQ4XdNP3tY2fexec1bBqbcntprXHDz7D7Rgq0aCadlT/hEZDeU/lT
JzEn+6C+mlCu1P27lqCQe/3K0SZR4NxARAdgM7Penv138LHGepJ5iocKYrNQpHBS
T4uT8Z3hseSZBTN94dZrYM+mdiKaH1YRt71pPmCla+yr36THo+72c00eOsbc4ofN
r78CN5p2uhp6b3I+uowO1oN2wjhvowseMddbIxG9Dz33OjeGoevnlwC8ihPFvUGJ
UYbTUYNig5GfBFbL342cK0uc2SihF9fNLH0izdXP5p+FELat3yM9jYAAXTH3PwF6
sZaJ/CngharXIWo5p19sOIQBYv9qb25OZcmSLeODQe1jk/5VERfuXZTneuvFSTZ4
KakeePbHqAT6+YdMK328k/JoR8An/aoKyS9h/OSg6UYXkMq6QlGtSLG8hIgXBW/n
0UUnDFu7RYPVT9xgAEcelxz5tMSDMJoeCTgoEyeSlnhYi0yYkScVZVFFBsTerkQJ
jcl+koHw2vnDfi9bp2ZD0NIn7etJY7146044XIMlpKLf/nQ+WXJsO9w7GY6GiycV
m0CzAiswYAPRP+4/jv6K8hh6ODCRrZr2RkuBV5r0Sg49ESY1VCNM0Aj4I8GpZAdx
c4qTyRYusydRWhP2jD2sF1FmVFWxAn5NfAS707ADsF9YqLVQvzizNXJ7uq6DtJ/1
B3iuFIiVUW4rfVp3LXOzRypWHYlBf3IusFVTHnDY1FDXx7Fxx1KpyA0ECdWf9+Yj
xmkhjN1BqVfsT10a7YYk9hMEoAEN4vaoTZLBMorJxr5RqAAfFzZQgcZtQKrGUn8a
ogOOETV9pJLA/sZBCyJeG6FvWaKXwjunsSnCuyw3F/TdOk6/WgFASq+zhKElwIsB
2sVDh9DmpLynx9aHHBjNGN3sUEJKq1d5gVJD1+GFlNYmLt+EdWf+HhKRH+/E1ZNC
LK79xqRai2Po3f/cmWQ6BLdJo/TDvZ1LXmjZ/uH/I/iGSVKIN5XUDW0nOttKZ2wZ
cdm3jJKgWXv+PRAvJCK2hAHqzJ4TPnsBeePvnK/7wlMmgW2oHBI5Yk+E43AExil7
d3rmjcxMDxUeY4Lc/pLUuiF4yos1HB8aIumQNbfDTgF+RpmPJSWMgMraynCTUeD/
HvjmJahWqfX8R+RlP99yL/VeFfLIUmj1m33pIzBXFgQMpFbsJinA9MLM/QegEsh5
KjBfw2XQEKxxmDZMtpKi77j6vpkaP89GFBRTLFbKsHxkHeiV5s8qFvZLBig0++o/
fJEdPWTsKfBkwTLy04RjgDYGn3em6+aMH+Gf1exnnmnGhWwQJaIUYImHN8MgZNiL
+pGA8Xw451mBsbKt1Tyb5VwL8onc90DDqDhBEx4xXFhRmt1Mia9gGmd6QO5ysHZj
FMBZvMMDew1dekSuvvNqZQ6lijV1IRaV8KkcyoQdk81gM4p+q97TzcsFJt+URJO+
YB+Z20ouuczTKD1QwFsgg1+hOwWy+O3Ih+tzY4+RtYAO6TX+VWxiKEX0x8+8sgCB
ME39K+lYePNxk2cHt6+mUtGLmeK0CNQDY+J6fUFSY38BZVtmfWnHqW8S58EVSg4H
7LTi2sYiaAPrw2HrDYfT9noLYCHhGhMy6Dru3qtHsxsaL5vGc+AQsAAMERxpSWKi
4dhdH5AcM4298MWgsapgdc2mjohEQnXRzEYiGqTpyKsvUNmmzEVp1y9a5BM8MhUn
QW2MvVC28l/Ext99Iz2hsQLqPf2MbCifNirm2msHFXL8JR2PuiLKFjPVDR29+DPY
Z262HmvUMgf80cJ9r72XL+6lK5sh5UymPe5sp1KKDJKzPVEnQpgZo04txaF3ropb
gx75mmsASZmvLy5aCc+QbTHu+cNuaxYTzmJTIDBldlBOgvWEaBvvNf2JuWPw5PQf
LtCAU3qO2pI6BoLVvyXzTsjCuZl4J2as2MFMxQWcV+fGgfP8EJYhJ+P3F7ur8H6J
u8jdjTEW0tNNntYQlShhOQhLEMS+N0TX/eE304LrO7ukYiSTwvuIjjr0bKgtnVeN
yOJ45EdKvSdwoz+Oa+m5VjJ6OB8xUsZPvi0U3YuwfKih3KhHUQsXki1jnTpH0KYR
JzhS+LMdY2x0KfUdTMEz78KxkT2oC2q8ILRIqPyMxA647DDQXhCw5+TFS3iCMyle
M/bHIN4rVSLE5ZZOWwXCIyP7joqpO+WL/2sTgjpTIDVlrthk5dujKFzeEzh/GroU
qHQij/0erCa2HdeCnqZw5MbfTDaYZqyS9GGXuTIOeQ5EnujidkaegQ8EvgZ/XykV
T3SqF9o6pJ+p+0kyIoGPC3Wxu2y8Mjo1R5yrBwTzVTKhnNWyeUCGVMiGDBorkcVe
FpADkSdxOM5HXpOBU3qOivHSBAjskOOeCSVk60SDostxoU5zfCgc0xmSSOdLvuFo
ZMSizAg/U3Y48KEMunu4dKUoXWjWqntUJtp/Ipkj0FT8Q6lookCqGp2P7RkQ2ni6
p6sHkUr+7BphPhty/B74zZZQIot6/vpYj6ZSh2W2bmMGarj8boBR/8buV4M0GNPf
mH1RkFaTbz9u7ZJxstRZP+/YhgZsxVz8qvjSk0LbKlYiKAKuJtvpYAAxzQ0C75xL
MtXzCfyqVvBD8H2gXI17u9t3nZW+LN0bykRK3StXjNZjfyGMoSDn3K3srNwZG6nC
aE588wggWDIp/iF5MP2+vBxnC3mhmHD8EPo8dsWwzd8kbWDYIRBbxMcWtmryJ3Sj
q1GYwtJ8+KUzRUFdr/zDkYLok5jaSlCCnKGnGbUnCwHTB/3CRq71GPvxfuWAHaO4
vFHIIgEF06sbXZdyxVS/X0auZHL5Tp9Untsym8d0K1wLfA8ImeVymE4MB8xYM++K
BvqxNh4NRayiJXFabpQRElqcZinullQobf4gvsp5VTgh0upf/PclkF+4VnGPWVy+
MbtbFGroMJ3J6gqiuxUTFlG3tiboxhbyhvhnVMYgKB5C73LCo9KC3QODyR10NBjI
i2pDI1pYpf9q5Xslog7L3RrfoKemhDab8py1vl6MuAnFB2SgoJZIq/T3FPHSqUlm
L8rx+1Z3bkvZcN46bnO77Cgoi+dGycBs3qafZBOeeRyFAln0IxmetJMpJGsrmwdo
SeGP0UDTlJy8uYjbRpdmzi533EbjPdoArU/11KqfERsJkymxoKv5j8Nl+Vo3lEAY
Z/LHqjpTPOB79tbHqy4aeemYs/Iziqz0I6q9qjSf8OZg6BH+fnIX9k0qNHZ8t9Sv
RKfRZLLWXOcbCRDeUILD27vLM7ZzPM/F6LorabPgxy0rn2/1x7xSoP296CV1gTgm
15HaUdPK4u2A6ZBZJZTmrVAqw9ZxoMcVeBOTv9rvO5jc8HpBg5eMeU/eYzxJJPcP
pkqwbUGel3HH6koP0r4mIHCqyqh4HKv/mVWA9eRxfEUn2yzAyXPAWyF2bHg+/sOv
rflGAJUdy/N7GYZhfyDTcKbMhGHY2gQqxMlvzrbjT/3otsoee2KYTYBv9P7PzpuV
79toOq31HNd2Trx6sD5Qb1eI3J+yyP3GdJqiBkDkdnEWG5O4cBWu0QasybZEoze9
r9/Ae8aaRFHNCvJeM0OYmRVYhKTWGylpNz5ClTW8ittTSHldCekUJjFFA6fFp86V
XGl7O4NDu/e7Cl1two1d8h9Qa3VIAXhW4wfufTVf5ed5BnOXishW7RAyMqfJjoyS
9xFi8DP1NljcwHCXld0jey0BXlvjZ4JN32FWxsCgOFA6D5L03vgJkePBaTIBUcpm
NPvstQ63pHtsFt9YJWBO3xNuxtKqeJxbtrZUfwNliQleIdIoirBzMAZ6q5vYw+nj
zZIxKANicgPWWb3vosi/e6nRtZcVeraEa6fw+J48p+ABk4FCQmgJCCBvC8+gM1GV
zpFZRdLop44mqO7Qlh2Nx5BY4k5vFy0NtkUMcjUjgWq+/k3yyTe72GaDFnrU5+/+
ZejrRTkqiAIzJHrZn2CDriplXBtyZizNp0vg96Fb8rovO7wy0H88cJdGDiIbga5I
XzgR9Hh+iBq6BQjDj6ngVKeYnqSqLavZ8tHTZdU/X1zflpAY+H4XzWdwhHQxcO2Z
rAlwNRQwz7NvIcIaGw8TpS86QZRIT+zoFTuqXJlPrbNXWHiiSG9c/YnSjrbudgHD
zLimcZ4BFXfutYXrUvAQfg+7Z2diq2sh4IuyuA7MbGR2lyIP32CiHoF+ZWk0eRRE
61G9AblbwtjVTjHZxOUVJjBwM6nv2Wn6bEXvDt2r7HHn90hIlI2vE/dEPiIgEDy7
FjLc5j+LocE7GK/BcRkxzhcc24BoclU3K1DBptVc+iYSVUs7iml3SofEQJLgDEq4
E4Dzb1SJyWU5WGIBDY/bUfbzuxZymWTH2kU+ogK0/HfL4ZckXkuJ5zFsoH3txtzh
lXLmZbiKv8qk/TrkO6n4ppR/f8sY7Sy/8rnsmWQdlryJ+dLyGGgC61UN36DHQNou
vNMUUxXY2rfDHGD7VzCE+xUVby9O5OxQ02KI30MR8tiN/9w9TaA0DXLaC4JsLiwv
IAagkLyUq1tfVOmYP/7LEtd5sp1jB1CmWQYXN/GKuiXEwZEDuo1gQEZdVYxvmju9
hAzJ5BuVx3IV9THIWgBopwQBW/O1DoTaz3Kf2Gl7mstv89Kt5rob47/vXVOkBLkP
ctaCHH/D5xKsi+ZDU4fvEChBB4vZdJvfn4dojNZpv5HIl0y2MH9RArXq9jUmGk+A
v9JpD4ScGCkI+DqjEdbbKwCV6uZgMENsqFi3TEFqEAr5GRfABavpUq4I4e3BFqur
2pxA7kkHUQwZjj4iJVJOzD2GUnKn5NLPZA0uy+ljZF3ex9CJnP4kFYDPClkn23w+
qB1a2k3JnaoSvmedL4/Lur+Vl6kEYb2DvTb/IctRcL9gKJzI4TI1jvGqgthMnh6w
5QhEDacdlaaGyoYTPW+i1XRfVwsIuj/TXtW47O5YcvjSRSdAHRUeC88DGkVVuyvD
XZcoI55ocvpf9j8PhmC7Z72TM5OQhhMBSUUhbzrHj4vNwKlZciYsJNIsjygg6bXA
RyTmj9aOlLRP9PWc1C6GBsBvQW9WFH0h5LjJ013U9tmU8PzafHIwLYUb/SqC5aFX
UhO+cndFuTyCh42vBZxu8j/Umlwv62ag4XrfqJQnl9RJhcZBj+eRf61x+Ld0DVky
RGG2RQfASnsPmBs6PlCC3k8kCROEab6h4eN7W7YY1U7EU5YATJni1PIex5cQf4/9
3RJhHmjpXZsS7Qov0C70tJpsme71sEl34a+e6rvm9vWmCOH53lGnjIFjM3YnKfhb
UBjePHACQy8CoUyTf9CdN3r8S92kJvQKKlQohwITeBxdMvgWTHUqyM9HrLsZFfQw
4joum/nNEdNM2cHMI8PUl6xu+uXWBThmJCFl4yeq9JtLvvJikr0iG6f4MBjqhxZq
3rq463PiIz6fVYkEu2laYzEiilswMNCc9JZmwNzLAEoNsbYBmm574rGx+phSHTkl
5QYAOz4HT7Tfhg/t3f1AlwvAQTg7IxyHErt7I+hPzudhAP9fwgQiJph4TGi+cfEe
j5g2owLizavO9wMD1sOkOoXIQJ+lBIFL37np7zfFqR70cp3ruomGl7z6b3f6QG6X
tm7RD42Zh1y2oRO7M6dcvBKYevzOQvrO0USvRyE1aVyj5nU+mgqKQ4WW/qs53GNK
D7mFjMWcOxxaffJfU/WPezJ6uGxaP8C4HCs9HAomKsgMi+xqU0TDyeakiGdXfsH7
0RbPDWdN+jXEpmgdgsq6WZkeMBo+TbdBRHSVUZYwVoKCmvhCdC1GH/OT11BtpOL5
cdEqGMfAxOYfIxjP41QKb3/XpKbCnP3jelI0n9HtQ72VvCxPWPkylAlrGjw/abpX
/n0o2lvYSSns+a1xU38vjOGGQCw1LSZykucDN2NeSG9jHox2ut3iq7kz5d+BVwjq
RgUfhjwPR8sHyYdRx5c2zhHPJjFntxvmQtpIPkd6ydZVHvYcZ4BUWEVICiEeM2yV
uRgf1zl+B+uIXnUuBofhvdHCa4G3emBRsiLi4gsu/mfo6KRVAffP2bzvZW+y2f4U
gZcXhb/T8nHvzMwTDahcwECblzW5pQSbuFFsvmxcg1Vu+SOzcSwh53Ej4YyihHLa
S8m5e9WZu+MXzUsTIRZOhgxp0l4XWZ5284DEvJmOZ4Ke0PWkZfX37Wc/JyQedHGf
GscBjg1by2nBcZv3R7jQYi2fZYe4IcWOoov7zswCYk8BuP6WotPPJtCFZchqhe1W
7zgRNny8SBf/GXMI55pjzXuM4IzjAvcWyINFStjVvU8rVcTLXPctSxGqP/JDah8Y
o2g7ZQJkxCqAfQhp2f1RpRDe0iX+dxYiinrBqwM4yW1S+G53tRQq2NlS9Utqs9K+
iI9Zw9gsvq7TQdOXe3VWJKPCyrJoGH0ENRBOhs5S95hRPZkRvMzfqGDbLme1/jE1
s6GRg59hBNtFSN09A//AEzA6cvi9LENGUJ5y6WPCPC0JeTtUFPIK3zT+3sZh/ab+
kcoslpBuZ3aALmioygn8tFlBAdEXwSHeNysvs6J0gixXXiuSHXBeUxfcbxtvp254
RBMTgxep8DPTQIyEAkTnkVpUjJbNqzDIm8Cl0IMgd7Mbv1bW0oKoCLuMKO4h3/GS
Y6Lt4IEVUhJETCFR9GN7UeSBQXezwtuqCy9qO9BFUqaKzGAXvennpjNMAxXi+Wyv
m00uzoRb3JCOYTxHfqzyFPfJorWvZZlzIuZ7H47x3UGch7Q2SYS+JnP3yRiyzW1q
oQMNpnqRl9N7nXsb/SPOFKjmsHhhHHAqGUIcWEUBxPvL1tJHliFVwqiE8s0PbPFG
JaB3hBkJNeBJaU3wCpJ3Tvf1DIj+quN/oBw5lVD2PR6hwGNwRYSmKD77WM99ncU+
DKuJCZGqS4vMPMYDs68obOPlovfWjd1lqjawyGsNNn9sKmMgXJ0nixVnlvM9griz
OZ83tO/j+3XV0jool3Oe8jKlCMAxxhjWIBAXTzdLFwpQGjysPM+xWrh79oaTLVFR
ddXqqUakoKJQRPlGbsyngnfalc2DWR9ztEqMnTIqa1w8Nux1ScB2XfhehiF3jgbM
ymIOaAGyYbciCKv6PmUAt6raGMIWzk3rXbd6YgRCQIznBgthN+nJQBrhuI7e6vjX
P/jgIftIpHa0k071WFJ+k+hdyaxfdjWE/Lhl3i2Z4hJxHtrdPqxwSV2Fyw3ZNRJW
KLQeOYi1UclEDsWuMLDbYt50ZrbEcqXppK4Ay08tQowlqJNwyEvHDEeTWe5vTTGf
qNFEvlNCGa7IunN+NrXGOTohvOnxQXIBUnlhG+qgO6dxJzwPnWLqinO8MrJ1MHmE
kIvcoBj19c8xS0kOFr1LFRRpVEjSSNwiiyhwjBlCbVgbmQXdWcV62Ciha2H/VhlW
gujcgUF9uKHAToXkU0bc5RHgwn2dP99KORVd2brEoTkuXqqWMPRJlcmAKISuBUcy
vgTMDhlEpNpqmPSzyT6eF5USwyggZdAnD9c9kgIPd2KldS5lGG3gHJk/QcR4blqr
ReKbYzTW/jw09/3AQ8tObEehUZpAI4WDMI3egTKVUGu3KQ+usYoaxinWoh0Ok2qM
hhgWLeXfee6Sj1GEoslhzGf2YZtYL8Npk3vFV0ypk7BoudMkXfUkuC4J4Jq9tX8j
QDLmyQRxKQgl5iLkUh771hlI0Mp/1jv6a8SJjXd44bDJQrUxdN6xDOiwWrHgzcpP
L7spwkmBnybBFSaydWBqoRH3loaMJgkwnp7dPO1KYsn2A+pSx8recBwbplg1JTUL
FaCZ97M7XmayQ45+p0j3fM9ttORSeFLqr2A6UsyW+DVjhNskSYV1savVY24nMzIR
q/3KxRT9wioB8fSsNY+JFUxN9NOLet4SugMi7+PPvDy8Dz7H56KldtCQcQRb/ok4
IIXLFViYFOKHBd4Wt0OF1U2rOV2g/avkgFYESuJOCIcjTzZ7hU1F21rOgCNct/mK
8ld37QChKGW1aLooBNQMd9J5JZ3aO/ujDrYE4UvfVlQ4e6tvVaIj9z/6ulOUXcdR
dtBEfdx07ZjAGIrTUb6Nzt9y82Ot0Uonw0orSRb2C30uBJGDrzVYrUe+BglwEcmt
Bf1KFLe7H5octdlNqXEpANe6IDwlivELaTM6ALhYfHpxG7ZhttOquwUm37Gb0uXK
XLMWKvn+sweD6gU1rHHT9CcmrgJr1lGie0XIge3m4MwefjbyJ1G2y09qiymYTMEx
Gkfaugsv30suwUSatg9rbxuHOKsCXR45fjyih0odUjmzCB+SCLRgGAp5Is0BcA91
sKOSP8mWyyspyK1865xzoRasrBQg2ibj8E0fbP0i5l888kM/NtCfqkbccQCC06+1
Xorl1K3M78KVCjC+nKVyQQxxbqs+ENepzZON181uRljeoMifNnkSGcMENRIZC9pI
prDLmjX+hbIx/7CGEltWTO8JDvKXY5SeH3+mxhpDeYSvF53rdcLVCaDu/M1gRuX1
BBJNEsaqXwHzy0OPxxtpZASKx/d8QRniBhI19x8/FVj9wOiutNVhdN0pWnMU9mtt
bk+ARs5qWLB02inoqAU86LqRQU4L61DWAp4ormTsfzRBvqjxSW2ncDNmYUCz0zfw
zvkJKi9Ddi2C6hLlzEj8V32nRLHLpWxgmMw7MqA9jagOFkfWUUCih/lDThTEuBny
dldbeRdpTXN1Z3jQmdYWeE7czlhvSo0O3LTJ1sCFsEMEQtkx2fYoTi2POgA9p78O
J0QCwVl2TcmIwEbhMSGhPlCSy0CuwUlN4JNUTn+jVBM2vhxlD9d0BXo9PQRS0Wet
4n4QypEVSkhGCcOflCQep73RPF/foE2CzFTI3VGKqBFrI4NeH+18zNFHfOL16ZAS
dwXVZJwf1yzFumRiyNyCgxPmV1iRJJ+DdHJxYPi9lbJLJtiAfrzdMcRvJuK4PuHE
/woOkXvXKb2mivDxK8UI9TXcJCv8FchLrq8Z4h4+F4LzuictmYar94/68cV9rJn5
+SLHOIipZ+I2l5f/QKEaYCUm2FFU3vYKBoVtJVP8J5OuX1RDIa+M3lFHFGEufs0t
HR98nu8Wr+5U9H/248WRVQjF7U/BzIKFPXHut9TAtV/aUoYuVe1Rbs8bssHgxgOS
DgLWqTdvSh08qPXZpyatZH9drSGmVue9IczO6dON1WICB0WgOQsPpYa2wekF7srZ
EnYcKlkkAiwZ7ezho1UJHZc4M/+HDf9I/+r/Drh0N9e7PJJqq5B5onfbBK9UmbC8
RQPFva9WKuUQaMU6Udu8lVU51Cop4gDK2MzsU3wzLh8rTAbhLgrOXi9PGN1fIW0E
NyIZFZInXJMPWMsv1bKAZw+Oc0b8fH7iVkURahcgbst5sJIK5XfZo0q4hFZcUJRP
52gKHP9Nd8M5GPzDOwKZP1g+o97jDvtQrlA3lax0apjHh9nVHT8MpbA2+oZVWo4+
sowifMvU9+5Ieyjv2cRwYSRFW9T9cRA651ImKmgMM6s10yGuQTEi/w8UiP3S3KwB
3BtkfZGKvSrm0t+qqE+APBoSNKefFnS78e0CTMxvcqKkn3e+LIAVAPc/9ilwgS++
vLpCaG6Xm4nPiLDyDgl5QQ73ei/geTIrsWMnnQf0GHMBjwg6lcfTt2PUsS9OQFmJ
YHWj4uRicXBOmwTSygV7p/TDHtt4SJvCaaHhU3vqzmkiaapkK3F43fEU+T/D1iR+
lZlsZrnqJOO7S15FVHw7+i5Sqxyj8zyHzXntOVkP4JHAaB7hUQkSz7GeVrDA+TMY
RqyCT0iB3Lw+PJ31waoYJa3O5Hlfs2PaR4rrtOnI2osPux6qRcbXlTOYyDdLofhs
6uzk7PQEuCxfllJT6aOPxZ78zJ3Q1RLypPXw+8r19rAfvZ5TBRtkGlHSsesJEcnT
ORST764hAc5XOG6KG+6iLb4Wwf7mz3a9tCDvoATD6vNHSOF8BbOq1mRZRdVAa9KE
dqcLEyyRwYTsZHEmuKpmV6tPgONpPy+c4iXr7HUNdkFkXLZxnpIxdRkeqvjsa+3h
L+i5WzgaFT8XKkeaM7aVtR/RRsFjGp8Ockr1lAH/+UL9dZNs4JLKnUcIkON2SSqQ
fTHHFPZQ691c4Hd8wY47jWLQOD1gkrjSqTuVWlccjxBy1M7wega9KUG5Dkzr7D4X
a5I1p65YsjawvBmEg78Pak3Dg7aPFXkCbVzfAKznStb3qeSyGNgj93ZwA1zMJYNU
AtqspZX1pSuCizyn6tfAtaOmP6F9f5Ap4TpGVQb2GLLjo01IQ3LF+n0iObMOEa/i
uphLdXqyDXYIfsZ0Ir78gjWT3hIeT7xU1bbcqJGBJPB/SwLZCl6/cd+/cWuQKv8g
pFPec/Pz56nYAFG81WAJU26jzZfC31FDJEvKPjTt2MDkmJm0Eqv8VlWBbWRx+02m
ijinJ6UeWRiRI7/RQhpaGr5gyVfa23j2zEd3GEb7IFtHzzmrK4BcyQNaACy4RYR5
/lF2fiha+ktRbQzSEjRodkKZ+aKnB1DNbdIIh0rR8kDi9lSgiNxuntq/riKHWDVL
kiac9wYfinnv9ZqpukjsW/QywqtcD/KzrmcdZoCyAsEUFiyoOihDYcKGO7L9r5TJ
zI0+ray4cBx4l56ljsdEBaeSOdA9aRsWzzJnUnvT1DJ1VV6j7SqWDjXq50PBdGVE
zViUYAdEQMQopxC/txpcGhDZTajYW9dDfx4C4i5sIUWKLy9nVb9le+hqaVK2npHr
PA83PLycHtoR1JyIlZHw5xbPdDi8zBoneXOZqECy3UBaJfAc8xWCvcqgM3dSK9TL
EiyYUvoWwvpmUH5rfq0jJc1Aco0K9BiPfHzzf33C/8ayv0+ZQ63j2spgqnio38YW
T6EZoHQYwgyhrXHE4kDoC9bBiBuo2rgkX6BVHOQHWXG/UtaBXRPPH/YPNPFhCckN
z+mTW/GebSLlP75S/UFxYg27Odmjut8KMEnxvrl0txU+4tqsp6cpliUpDC0AKvu2
VxInQtjz3JeHdX3NPztv+CSixJyhJQAd5oNDuvbeI0gibX/akEjqe4fWEdkFUvYe
6L4Sk3eD/etxaTJ/PjIqn6Dq996/TtaqQqQmWK2V86rxpobgELmGPIBMFMNt/KA2
htPUnSRGSfj7+DBgbhXo3iL5J07ifHvJDleVUc99XohtE3qqPsDbv3UTJbjZBx1B
72bL88js9YqmdMJV+F/xpwZTLiwBcJCgG5wFPQsiQmFoTnKumHLBo6iDy7yJnj7H
+bMoFOR4jYVzywsDTfMf106Z/oyDAUSH400hMH22DaRg6fWk1keXRjChQ2E+gi9H
jwUQSTFflqiE44/w/LjdPHf+s9NdHMDIp69WO6rcmliMkTAVRLp0hzZrO+Zp/kGp
8wi2RUeyD4ga/6W5Rx4LfIm7iYT0R7Fki4C3dyQuRqgOrONJPWO76cZPnM0uYDZy
IlcoMUL40YykNRW8BpOVSdnWaazqJ75KC0abjoMuhfYO3pw217WPjjSAc1hgvZAw
fBV+y70DwuJpqDAo8Vj3ENWwCXQ4qizJuoSNU1bB6vX61J3zlf1KkA6fvCOUwyA4
oeW+QQgEKBssQUBzY7m3MbanCOWVjYPD8XI0wftlsTmUDddM6D/tSEwAG94FvOvR
THETq8bkulQiCv/hyIAQZfFVvN+tsL4x3BjN/rQ00P04c4S3im5rVpR6PlRV9Awn
1GyJBWD7l99tVQvKGRJyv8xQr4xzTMtX3RrWnYx8l2Yf1G/M+3r5k9FannGhCPcp
JAk1DBwlkiGqgZm9P3WdrmKTzh2++XJNGmT3oQEMiU0TKarxZcwVKJUdLTD59CuN
mXnNUPkT5BbriPEw71NpOGsD8RV3VfUbr/6wTBV2HdwPxDvqvIzYUHWvIyxJYofb
snVQRgmWtJgxPEp89/oUSaLol5EYyBptdMKDabgcQk6nMkVcj94l5Nw6XZf/IpoV
tK39oCPCyngsFpwxVy0snZzIgseLpdY7CDq/NVM7JlZ33AwNyhCEp37h9Lk4pM+Y
tOt4Tfd/t30umkxyZl5rZvOigWJCHFQppcdrqFFcUwpcT/HEu8IF2SVB9Tu2y2a6
mxjsdehtnPHRsAgBWJSWRwHqYBYTaZQNkhF4Cj3SrAc2FQ4RXAYZ4kglhEUoEAgf
mckh1x3dH7WTUce5cmG6DNg0RJqMPn2GX3FahL2tVpYih+vORi0Kd/6bQkCoIoyA
1an6ho8+VFU8bg2le/LM4izFNo9AUjfwoS0oWQK2V0e4Z4OXLSnIj4QCpSy7dg7A
RY6GYx0+b949poti6GMPwV/Lp/hwsJT0AyfJ2ZM3jMgdgHAZkHxYDK45T6xsnMx5
5HqgzVUIsHcoHfVKEpSE4/uJBIBDJXfY1Ce6J/iLTbthXxOsGzF8nWIrde4gooac
X7beEDNkaNMCo4z/Eh/LOOrnc/jC6nNqeQsF7zTQh5eJ3zDO2Vy2vYucwHrvVxSQ
YG4ZEvVdX01xQeIAU2MSY/9U16C8dpFZfFGgxMLnkdjjCri+/lDcMQfZnNcamtXj
eASLbWMZoK1lt8YGL1SzpP20UJZs2QzHdX4N+n/uWP6M/5uSj+Puy7eqrDWLRff+
oD6SWlKAZX0wgdRQxcuoABjWHXmNqUPufE9FWP3FKP1Y/IIj+TUJVisIHMFsyR/1
/8U2J/YuaOUXYu4S1+czgzWTlhTs0/0dWUNiav1ecQwv3H1qdiWSG5dYNfwmcW7U
glbsVJoAQv0XD5RaMYZ50WUMR7h/0zk3+hoAlAPg+EWKNGJ9DTIlJCCJ6ExBBTwp
wEpPw1+V4Qb+Kli+HiHE2GnaKUkyZrf50QiECGGlgrYn+/1BSAVUwVWuGVqXzxuH
3/VW8sY9Kgs3eXSCemk9atPvi0uBHU4nFrIZgpFguGbKavZsqjsgXe0UB2uPFKj/
+N+qqtmCvXYFE00cjnZrdOs4nQi/9JL6fSxITmejMQpARfvneeNpSoocWNieP4QS
KW1F3i8OihCZoTMXg7OBZpDQNfZm1HDhsdIC1kteuGLbaeiTF9rjDSvptrHbfA69
RB1D/E7K4uIp0PGaRFfTdfMJt0HX7E9sDxt+KpJta+tvH1cgahotZKYNZSUhXolw
JyyDA98wgcQawt5al2WWcp9x8kBiImaj6lfTfp5I7JZROv9nL6XUPDIjLGm+erIV
kEOZA7FgbG/1hJo7O/zQiHF9MWkt8dTdnqrii80E9piJJvtlwUD/d70IBBLtrVd/
c0GUsvADRRzQ23FOrp5D2/ebArW5lVyrG2CZiQp674T/UVRdNjwn8SbAy+061CAX
HjWCn4Qjq0MVelgzznk8FgYvD/pO0csCGreVZXKtweE4f4iVe1rr2MOKjn31IrzE
iW+X0DXSVsbx1efHk5+q9DgOqUF8/oC3cjvHR85zgwtQ7nleYmchbXZg5cVqRbP6
9E6PbwgZ1tAOek4BYY5DsE904tleJkFaQTOvAl+DzMFqA+Rl+zqzeeLFM1582yYn
tkeZfKfqNdRJQniwfBG52gUCyfEesKzEdEOCFILzaCggkQ4tP6TWGTtT01by7XTn
NcMiJeyTZsQUywq13sWt5nXNxf1eLUzILyXYwasi2z9qOGA+ox9ys6LvIbgzYZzl
xdpY6Rziys/YQGKVFYr9kiKQr+A/snF6GASJt26rf7TMc0sOihny6eFsyGuFvvFk
oSL3UbM21XnPJ4PM3VLmzkpQ6wdNf6ejWRD4Q/PDEUlbXN6jSkBIOHayE+FqyUIL
xxqtoF3+SuW75j9iDA52gYoTr7UvWrTrjfX1t0TfX8HMX68QqXiCTqi3f6jiICZb
I/OucTSdxy/JCDP2FLlLfRhLiynIyUpQd7lHl3R820MsHO98UOqMropsvVfBjvDu
rJ/GdhHORSpL58+Ql1fnd7HWGxt7VrKGNqxGmLZCJdZrq0T/t4gav9bn5cGUuZ5R
jhx7ErCf8kFcpzf4c7PiQnIe8xwyRRZnuvZjC+SaxByHwHkKjBXP87a6+qOrDq3h
rt73PsU3xUOWfT1+NHxc/AOrnLUL3PrIkfGzfhDhgmnmrwSrDnjhhHBcM53HO8wb
xhxvLjEbuGmnIOTIxKnpr9VxRvqyDF/OAC9doiBp54DdlJPowcE4VYB4FTlXZVvm
/VNybDaBigViGfAARd61rXL/eqzD3N59D+be6KXOEgO4bMRaV0RNntV3qZl7UCoS
pzfQqgznAhFr9jNhChelSPAKDs4qxgzv7A1MjnFgyLVmiagKUC+QJ6XDZqB2Cfkp
9rZyCPSvFaWq9q+uSCQm+1kZP09xoVVKgQ8lp4mopQ/pFnGh9kO/XmAmq1WcY3eD
hU2m+ppO0OjMb7JFqon9B5rZUlnUJ1YDX27FXrFgfMdUOxGxJhpN3Gz52cchV8OU
Qawt68T6Ldb2SVpg+RXj3MyDSAz+9PybP7ichbaRqGSaTA5jJ72OpSX0BD5PoObf
gJUF3aSc7rnfeyTO4vuFh6euuZWo/4uWe14e0r7UFIv+65R9NSI8XftVUMhO1K67
4YlF74r3LHdQ3rifLtfsebkZ0d7SKKbr5RTsjDLogQNmGw346uP2HDlNJwzdPPqf
vd19LRfO28ZCye1nyvpmi0NDv8IxJZTf3DHsIietrEfuGHwq8Ggl90uXXaeamgG/
eoU1qyHSOw/SnP2F3WTLJVBW/hJc4uOtQt8XXnN+PfGoVvmI2JDee34waMdxKH+d
RC6gxFtiCJcN61bF1bDILTEP1luTRMSBRV4YPqgMFoOwQ8p70BxE+eQMYuhpyhkN
GF9wki6P7fjHj1zoV2WQlGFFU75n2f7U0tAlmFraPpjCCMrq2swOh2MA74CDQg2B
acxewfDiAf8SQTrBbiHyhzNb2KMIYGdTrDcWNs2IuPSgX94DRiPXXpQuV3166bRR
hAasz4QGqj0YBK7/Gbu/5pI1F1E00ubzdvWjE0Fi+N0DQ3FTmsFo2boIMnnDuWHB
IuZ3mvCuMtOu5QagFb9TnCxXdN5O2ZSeAcV/Hsb2YfcGZSlDA7sJA+oED1Cgknmi
A7I/NPQ4+Hr1kgivu9ISS9AbOph9bw2VKHxU3NKZ/Ftz8Tw1HYADN19+BEd2yJSQ
0qcCU4YW7znmhu1Ow3YLpDVRAfJRcIx2v8n4G0e3hZnYTjUSW6LhRx9l/hjbtlgJ
AVTu71M862R31kThVWfJrHfpcy1crzSlTVOg2+5Kz38v3cfwq0KeIj/rPSOecgoc
y2BJEpVWY5c2bBd0zWXHFj0KXKz0XIhZ0RL9FeX+7L5swu537iM3EzpxsHKSL8pT
1bY1kEgIZ4VckUW4E9mZWoD5JyzGR1n8F6PRVik8fC1Qwss3XPDQK2H+E2WZivFs
X1pjKZJberhk/MrBR5MsktOp27tQIwlGzISfKShId0OsMiOZf72vq+WWk/yrtXVI
Sn+/y7Agzpk6/xnjc9oVYRPZloudV91xtlevn1+doVO5WUgFg8Z0K1ZzKMAbsutZ
h5k0oqqsFvEsJ7v40XsAEPNS5G06HJ+Yr0TYQjqoAH+p1EMFqmVK2tMHMS2FgskT
o2U2mHCUhiCuBoIdYIes0PuXMDbdJdTIb9afkgYA3kAocJwcc9cGSBVQv/ilCI8R
vVDrtaJWJ6UvyCNUayNeAlCPpo/CPA7zAR/JExzognoR+/AIlmbCstJcYyi8yJfp
YjAj2tAY8uxBs3CrNUQLSz+jDPnTKabcvgtOsIrvdc9yHl4oCdM1mHUSDs4ikiID
WEfHZvZwqhh4By9alkv4WDJHogK3Yp7TZeOBDqkA6NaRaPRx7ODCf+sCX8CUQ5OQ
N2fP023S0RIkaT/BkOA085THOxXQpaIrohK/ecrN+2n8x0SD5n5AyT9JgGjciHSj
K6UepeK1iC3YdUkYLdWPEi3sSp45udKWV61xrptoqHOjTBiPx6sA//rSdPwgPTHJ
YB7lBiDWEBaP50dJEU0hWWqcYGyUwPogbOGEO4UXCqXS8OtxxQHAXilPnDWoO1Y/
QbRnoh9w9GCU9uiIEJegt4Fe3chiaqHgqb3K9zj+hobSrOwTjKQG9ye4YevmN2m8
VD0m57V/jEMKiU1UFXYbacAMJTvhk2R1eulrBpJ5PZlGVGVPArDe3YHvwp0h+0Ch
QnCbRNlrYYfDZV+39YBvqKXxslzXj39YJ1aMvxLeoLN2gz8Zv1cKlQAIogVUNmxn
8t5ioV4ap689IU5ErPrBNKCtu58roBCDM/85mViIuOglLED3ovY1SgZks40OxK1q
ms4cIwZacaYjExK4Kq4Kl8ktKY5sTh5ZRIzk1gHfBvdXrNQxPNs/tGJFm/GP5jcL
jVyM1BE99FUJfLSBiyE4ntpuKUQyNwysaBc/bpXESsjhhhC1tE/rTlfMI2Y+WX8T
zf3hZd3d4YXKL2RHqOkkCk3ChFdBiLCbOvhLFpF4uwYGWxdFKI7HvIGmZI3yxEZb
7kMcKaom9eU5tyBk9HNtK3GHSL1lYWjdWHvpyRKt76a2Rwtkz/DjjYUlGzVg+VJP
kcPXLiRf9bphtgcX1hq56YkdPL81jrPG3HUhqcf2EYFbLt3UWk2lSH+TzCrckhHt
yKRrdiT4i8GR9uGoQYtoCVhqz+1XTRxg0V1UjTZ7DA/aREev80l6Pvz+FBRvAdCC
jGQaKvniWiLUn5FLJaQ9tkGbofMXknCl317wlQZkhpdAFShCopYheX8Wlwaue/DG
6OHFScOucpdGKecEgXHalnU1z9w288oOfpUWh3N6e+NMskScuhx2rP7j1A7rEQtc
YMmHwh32Vo8xlfj+ntSGYZ2WkEnBAH/dXjdXm3Gu6axNo/Fkqqw9k+UV5PjLNPB3
+lNFRbNOJoFbV3e5ijA4kkfuUrWq6XlrkqpRGw56zf2z+HQ9u97hdVNk/s7ovIK2
zpR3/cYSOqJ0kOreDRETvVtXLJrMC1Pgtar5soPQT4M6teSMj6M6SAe1zxbNDx3B
l6CT7DmAWjexFMr9NEhjMtmavZ6FvB7l7T4+JhqC0CnRyehPoAMmg9eP3+IPsX29
9x7u6iI9+SqkkfZCoCM523TA7PyEVw4XvkIZlNkXHyAZTP5rAEckh0+Gq+pUHzox
nFdZ0+hvkwmS4t78YyO1LX4a4i0nc0lks36r1rd1+qTON3SLRhIv6YdmEZdNijNo
PBFlqv0QriA7R13NAGjJDYwxHwT6Qzdk/2KLt0OIbvn2LvJbyzBxvGJlVori1Lxt
dEZpdqbMYq9xbPK2NEEXng0b1pvhznTLDozYsD9IthuxKKoo1m+ik6eTNLo0NWW8
bVpbQnM+YN/BAB/ORb7Z2LWe42qT8ptQi+ane+QNcsFPSGjSI0wIKZNm7kxeHpZk
LgtVs8dP5FU86MZqgj59g0z+2P4Ss5a+TQnMHrhmBXG5ovvgUTswy/x7tq4a/Y2m
EnekM5JHBMG2m19Sd+8PH6VV7zmkDKFz5aHb/4vE2ax8vx981wXDOEMMBjqt7pT4
icJE7gV7WcKvDF/Tgn8T3fIlj4M5PDkibH31zprS11X5eL/CxuOCTLucdJh95rSf
PUvhHDqqxo0hh/YZ0L/bCS7lIx8RNw8bgde5Dp8ziutxhLiT45hVEmOa7D/RGS+C
hJEis3fxJFRhh67njmaoIy92IEwPkyrs4QwMCyOF8/kG4ECUWTxPWHuQ73vzPKL9
eI1oIxyggm1wnXXJ3W8IpNPKZeqsmwcg44erzbIMmpwhvYup3hd6LUR+yYJ4esM5
JDmZld6tbU7VVdzSjEQZ1EusPWxLTOttYpxvHueJv/GeC5U9+cA4ISJGflRRxvgV
CiFiq225tyxqaq5eo8YHEi4QVbl+C5M/9M6lR0W7qd9G6B9nc2clrp7fwkxaDn9U
lGkna9njJobvMKy0LieXVwGudWVLVky6TEz/90DVw3HMN6a9VEA3ARAfQUEi4+VU
UPGOc9JaHWGm1oBQnVP34t5O1/dmwDmFC3TDIN8kJX52GhvrMqlDngf4WblOZ3nk
yo2SpPGFL3HazizYkrl8frLzf2OuYUA3tEFvRjl1H+IJwP/RR+fOvPCTuok4y9Zi
lA7WaiVFV2RD/PM9njCD1iEiFrvmtQvpWilmBXE9f6xViOLHDCAvlwDq/jCqKdZb
Xx6N8WIFErgKXWsRBn1LS1vUWtygZyZoDH/mOd7uK4rg1bA97kbTL8lwSDhaK6ZK
/UmwiJcskvyElrjoGTH16tEAJU8ihOksoQtth//J5mAWcsBYL5EgnbhjoOhkMzqx
zaLvO9okTYS8U/IF43Du21H8tQ2iV5ITnlQEuz5alKB7APcBfjD6otWP1ZsAwiFW
3QyqlHXc/sN9qnSAmNQg1eamZDs7zDQobHKpbmPjvi/dja6dnrZ6uL1NEWZqqsNR
h/mjKWrSjE9/QwaYNppPEL+z+GPOzcM5KmkE9fY+YsMh4cI703w1F8NH5h1Ulu1V
QakLN0ckRSbZL9uTFO4J4qIc8IXZnl/9Y34vEzHfOm/BCRgC3E1ScQxiyOPxrWK6
cfXyTUWRRtWKNaQGAPZ+W8fLErfdLtf/psWpzg5HkaeoY8JyqsCUO+veY6ommSbL
H2H9IEYRmsjJaY2yUbeYleoueJMVk8fJJhD41L8iXD/mhHEaOHTmMuhv/47p9Mp9
IPSBi7jHdfEj8wmRGqH183QyVK8qqtJHNMj0/P47f+gVmHp6wMwVdp8oFmLAxcvU
qrbhvGQfko8AOQC8DiRBla0GptZ8t4OjQsC38wwfN1P39fIkpBwFIgIhyJxUnde4
aaNHdxqdYRACUlhR4tOYoNocKRgl7fLyqQy3qkVriIuAZVFcq5eEiD9u8qV54I7N
geFY18BmfsMtnsEJVyH+AdL6fjcry/mJy/y7yhv76yz8S4A55KKzAH4ieUkwtfqR
mlEDn8CgPMfDU0XqrC7QBiRJrInWiHgeeIIKLnXj/i/iTSBEz9WesIIlWjEvCABn
GWFzPYsajk/kNyq0CPK25W6/AuZaOoZEdERZqgitr8EOfIK750rZJYPyl9IYVFu5
3k/CJMWGGR75/eOoJy09H/MI6BChuSZJVkH8fw7a0YPW6O8fj3vVIgR8ohtZ+UEl
1f/jRbi/StcPlYHzQXoSKRZSKug4Ot3/RluyJ1b3YjSyu3k1xtBdnRghfmoXCZf5
MsObxQjOjPGjw7lwSsnL6iXtxG9ULrZ+acMnRNF46MQVrUkcG2dODmewyS23EG3p
LOP3nU1SxJQHEf70Ao2Rzqt5x/x+iCtvxr6088gQYR36fAcdQe87irC05Va9U8NP
3KbKIK8FrTLt4ev0V8phT01NVVWerURzSqUkoGnAanRlyCtT7TB6XSCQo1Zd4Vo1
29UH4BUgGia2O2K2KChEGu02Xx/uHl7dQyMae9XVC+jJxptugBWoN5tGu9bsoRB6
JJqZbP3rarZ3Hueuwdbdm99h+3UMIzwOfsAyDM/Cemc4pIuQ8erNg3oXJxlctd3V
TW2/hmCLZLjPHzPHT4ros+W8bzH4RF1FcFJ/GswuNrZgtnmiFstjvcL8uZPueG/q
OpeF2PAOYGgrELEadpWiYgncRbahbh2TlvTy9sJtVNaY7LCNa9A/Hq6u6Lv6E5Ib
y6YgugYPqsDwVk4uj+Jn/8xsac7Q3xlIdKwlMr2yTsfKIB/BNK8vBlCe2M5DX+rY
1pDbQhagxw7GjfDeyq5fJiLAv0gk0BvyJH6ogSgfiPrdFZ6Ux/FF+U/XX42Itlib
8gUT1OFBmdF3xTGvIOrH5AyGuqnPBzGFPlv9ibYeNQaS9T6VLg8zVJM6AAAHiJ5A
Hc3prsmQHMk7BdfiToMH5R9Gqqd7EJvnQY7euDFDRRXcg5mYHI7YOA+Uh5IEyz6q
+C26XyQP1kp+0Xr1sBjkSb5HDQX2lna0tBIAVGN5xgVArj74OOno5FCcFRpmiw8t
ZW2ruzFN3jBvZtQOFvUJR7T+aUXPPiNS0yQrPUzisxHFvmo+DGzDCWDFtx39FOox
mxtjWIibDFFfm2iDR1o+MIno0wBWCOPyK9d79tCpUAmaFNI7PrN5t8fvWaqa9MWV
ILXx353iH2nJ3aSikwEJxCsRZUmGdlwcfyUs8sGivHByHLqV2AHcIF24ZKRliyu+
TFrYthR2cS9c3xqOFrLgfoM1oJ3De3PXdcUWwvdS9mf/6rQcQbPc2fJenLpwFsZL
rb+1SukpyU9WdgDPMx5CLHS0Zf6pMHUWR6Oh9C57KDprD8RoddWLz3WVi4q984gW
9d821Gg1bQzlulmCZ7Q/XJMvMfAJ3RKoSSn8whW77LragExBKkzarPDOzxMNGxc3
myC8Bcx2NXIxxojAM+RYeI2UhMmuOIHcfopb11Xt5gZDT3KzhpBK9lH4IyMRiSU/
KA/qYQQEFeXa1zrCci+JS3PTlG54Ga2Noi9iv+8zK5bZLm3hyRI8C0zWtzuBIjUF
O5JytL3efznIdJR1wmnLU9krByCqf9UiM0lJCH+QfKPynGYTNLUxAuoc937bwf8F
aj6FOsxsxAZBdaJ+2e499TuBp70zYzlmqEA8pPldo1EDextCi33tjYPUazX1AJpH
QgMSXGg97ta6pSF3R0k8KMN7Aqr5I+zc579roz+v90O75jgciVXL78YINlkRxZ+f
KPS91LUVtNDRM79kg16znKEiODn2dVTgcwOPko2MqQ3Se6Lbmb77fxFBowcYYDqd
n4ASLkw7F1dm+8EoVOQiiA2XR3IMccBe4Ef243hjTMubE2wq50/0eme8MgoJdY7x
/k9HwrCVgxeVBWjxfisUCHv4aBdPFihP3nnk3dsZD8Zh5OKWxozKFBk6NzFtud90
AQJ9H3hey5ToMEfwvrmZ7T1fYUCcuYYfJegFdfrkW11WSevL204Hj1fV3CXlmV8p
8mRbTHafGBX/0KnOHjwk46M3mF0DDtbxYTrYkHlTjsMXO/R+GqBdHB2i4xIdrJAs
hCnB3yvfLoETnnWVhdDRxybRzwOxJSd4DyalBqlqBXlUz1PvnLuJ8SAsZ3D+6ZDn
cWPBUyyLyeJdBpgR2lbN2gfUCjfIAq+Q3Yfob7yJWqaW1HJvDmA1Jb49n1YockqD
elo+SbmVqgca0LgADrqSKCMxk/mR8QKd1dbmXKuBnV8b4SEmNne6SkFydNtxI8KI
wgyYE2B6DIg+03jWlYWrTUJ+tWf9/mm98tu0EPFlotOKV0BEBDGVJkLpgShtEYUO
hkjwFs3xuSVpw98CulDckx7eLXR38Jw6iu1T1PNV9MHQGQDTgtscMW6slFRQ6Ifs
3KW3Pgbzk9fTtxtiTf7ZkD6dl6N/+IHBYUt5HkVrxuW9LflEZs7Iw3kzav3wpNBX
Z2JKxuOlH3TBEs4N/+iNtnFZ525HH88Z/DZ1fd/mAiTK++p0fckypyJBeqkax3dq
MH4LStZXZp9xuvr+yXfSJqL+Av6NgVJwPg/yjoxr53YyqIXLGjmTIZx4jrXruexV
b44hIvpmKYqwTZUQJhIpH4QfO3E08MD3GpHTGU540vhaHz+0hS9cnanHqkTH/3Qn
fBrbkcwcVPUrwhpmKcR36EW2O1ZalSHAngfm8LhNTu29zTlvsmxVO9YfNvnyaV65
7kZmrLaGUW25VBR/T8AgAcwzJ9FeYy0FqY7yar9D3d5wX0hzHx5+CsaGESLOSypD
KV/cv8oqt+ZsPPf2onW4vvA35l098qSbKeazxLBbH5T4xYAmxESW7NT8DiAvumLN
ICxb9TFTKxc+YAWoWfw+rWUvvxkK7mRrPDH+icnUnisTrPsF68aDztkrlw7Pt2l0
CAMl7KV0FkVv42+gkZcdCvz/vK5wNdFJ39L3A87KpFGBET/bN2uDjajBOAbdCG8L
0z7vCu7dxfYGcjL8w5Z7jEGbTF543fGv/Kg28txhq4AKFR4Z8fN7dcQqrOhReztt
u5LqB2yP6laHKrBxAJYWsJew1W0xUaZEtHGwu7VVHvhH6/r+AT61FKZ65Op1s7zH
V6dAm0hzYoRM5QCJZZWcjGKL07TYWeR/qJtgeoR41n10o/ZaeHSK8U7itWieet0f
Z4BH4huirFJw5BLGbtSofma5ChoiL/riGBsmn6+ii0YZY6yd9asgoJhqOtvRdIve
O6nX4jmTUnOmCNFPGE8v7n8L27Ecm1Ml4yCx3hOYNM43eU4HckNBfCYCQ0nUSWgO
zScpxzThIEVeALx2fKrGb9H1wqbASJggkP3oHjFFSs62oGTatGvwlYFPuifQcwjs
Q090orWC8JeUSst8IQOfinFZtElMlaT+eX1mIAR2Nd+xoMFXI9fz575UM1djd08d
hdu2PjielDEFLq57C+nboORaHVgEjov3AGG0BlQuMPMPXL+mCFzu1CpapvlQZ5C9
+yEkmwpG/gXHfV6yd+p+pEmJf8B6nGHBxe0vvsjFoq522YR6sLw30wAKCilLnGCm
SrbUTl77AmLJsHLOG0GrR3w8G6vGlifLhqbLYROGmzkU5wo6KSsj2T/gzaH8BKA0
nOD98Z54CnnwSap9WXXPSX9BA62tfkiLOPoNDzRfynvBjeluypSDdu25bppltk+e
O7TtqTSTLc7qZR3MP1FMdLAqBZWIMjxSGbAwl3hUx2fZlzFaTCEbYxBmiZzo0HYl
2jYrSmtZtdj2X1QuaKeSgh6fhOqm8Pe1kYY7i3p5EIXaOL828JxTM6KDvV/lCf1Z
izcMRfOeQE/Q523BUERj2qIyWdzutasU1GII2ometUm2pNpNWtgfFkke4u2pz67e
a/csaaatELbidh2YboVvN1iks7G9RsqVZM4EDaKEv40ibcDUVUvKbNQADvJbgwqk
tPdKYu7iH6QvvJTOGLLr4f20gA7xwpDiOtz9wRNsteYwmcRxhllSgs4bo20nMhyd
NChs/3OidAyRh0ZQ1HaXmVpQj4dVBYrCwir7Od/+C8wKvW7oi+Y2jWf9zk5H0ptf
VECXLa2Y9RLQ0bEISKl7SuKZMmfUdJ5htVijUJeAbvfJU5CeNggv4F/LiyypNQTx
+V5fP4L1WzF8OlpJo0YQ0ijnd/jDK6zhNmfXhcbrew4ge3p0a6vvsAhIZGQBDVgp
0Ol1WrVElbTl0HQ3YAT+NvgoFFTh91G1BIoHbY17Ajnoks/HG7Ab47T6z6kObnbo
EmmILTDTs0io766z6bu8QlEQkq/DE6XhUAsZxlpS4ZVyY0Uo3NPdCKlc0drMwbNv
4s37pDee8p25+9QChU+15AgLAARsV2kfITy9ikhjiH+MWb95c1fWGEgABPJtYUR3
mIaKZX0b0cSm1NTB7VQydRPkBDWO+0Wjg81kOev8dftiwXdZXizeewqlurPOx96C
X5unmkq4scPG2Q6jrPUK9vE7csAEwKMyvWq3mFCBDwUdUfcIgICbJK6qyhtOUOrF
NgiX7QXvsul4KkOnMLMGQWny6kKFaPwhb2w6FCAtQvijuoven6fhmYSKEnNUPIiz
j8qGcSMT43Ap9xmx7k7bQmjuIxHVWiGInKOZIeuRKcw4rpIV+/c49YGVMPuKCjvb
0fp1nBrU75BLc5DwD8bDju+hblY7oUDZ79Z6tGFnVowErgAn9ujr2wooJu2a8VC6
J5xnlmrJyTCRQX8SVuQ7uMDc5F8H961aGzTJR055NxHQR7Nhvq3UFtEydvu83snW
k/HKy0IA8DLYvdRg0H0DuBV8EWGPQKC8wE1AF8q0LooYbeRlzo6u7/SNL1MhQLEw
pY1LJ6h0+OWUOqpeuYiTZzZTRGXBtXMjB1BYCXnTtc6AJXJXxJmgOtKI1ltkasUN
EgjKOmoN9MjOaJu9BiP1G1nfcyniD+nI/zyJZZpeRnkYcizSE/fDB+8WR2AvwWVU
MC7gUc2Pep5dcXDmRxasPLkigzH/uDSWFoW2g0/K6gTTBu2WmPnS3mUun0qOA8Cr
HDiQbCOWL1WoO6JFU4VJwr6L0xk7wMTE0biSDl3OXhj2DGMZMjhberv1A94YLyXf
9VQQmI/BxPvBemY6w4NmgbP8dKeTFuWvDLPOeVAYwrg4SyJho7rF9S0ssDvFhvXr
8gvtkqghLQDxdVNCikts1CrEqXmi8NQ9hhIGb9KuV1cHeWc6NDdkJVX1Te/pQW9M
XnHnwH7UZu9e34VCfjhpU/docoTyP5IdgLzcoO2G2n81pqszJ4u3+Z1X1W73bCW0
0cqeikbRkOx4QTdMrvpVJxvfxlwQEq3O44iobRg+eMeSJ7/Sq0LYxvjPvVAcmasl
EzFZTaUdTPnfbORPOqe5wAseH/Vcq9ZyUxxb/UeGxIY8P1WnxukQSAJvQ6dCAnf9
q18RmvmNY8qBo85AEToHGIsxnTQkjbcBuglEKaoxqNDDW9KFBq9jAIFYTTvMRfEk
yg2vRf/6B4WDiUspCS06zmsj8ZBDowj/cwL9GPB6kWpvC0cLsxD/T0V7D7QPvt9/
HOjthnf+mDkkeqBhi8gbqy/+PsWrVzT1iQjaf2T+lC2cnKo7wEgI7JCxxYhj9X8g
2ra2s52NdVKWOxc/mGIT4EEIEVENzr8NVTQIVTWXUK8imPb9csGSjiPh1XKlxDDJ
5opQgJi3k3IHTAHuotx2pW5jFkfsa1qhC3JY5c8bESQfIe3E2svE6R84tj3Wq7F5
Z35L/WudR5edinsK9+NBS+e2p0YuKYGBwelMJfYVH8Q42hnhYEBxLZII3S7MAfwe
71ekVJTmoKAiGLg7nyViiKbSbVx7DKoVm89seN452G6XLGjQY8j3BOSds8Ipg/po
AawoIU7I3bpEr2DqEzS4vJdK/i5Jow8eiUeOShersBi8CusvxGVYxGyqmfxgOQc+
m9t4GAzDEUMtinipTNROBwHehf8z7h1JoBoJE1EGqag6s2o2qdnQAoG2lr3DAkcb
qNaHKep94mewGf0pT2sVDPPELaxFtzBaE7nMqVQbGL5VUyGj12skgXG8FaP/IU94
+FHaQJgp4NHApgzfAUKfptGjEC7fJUMtWHM4ayv3HyXakhQHd9WFc0s1SN0eUpPu
RvG+l3hkg6ab4+39BJvkfBXlOhRYM/2CNX0GVbqNGW0NLg6TUC0ohDD/jn8Mbk6V
kBVIODqgfU/JMx4aqMcDnTgBLYuy2n5krJkr18H7K6c0//dgmG6TyXZaQh92TG6H
0a6fUdYwneUdeG+v5ZqRfvi2fR6aAXt4e1NXFuyPHQnT6VE/cmxbXSORzMxRv1Qd
Fo/DKS+DY6QqnHpMfRCiRmvLIUMdjm2EqqQrxwXdpSfyXmUm5Y8djt5lDkWpMSvy
++gsEYllIJMwiRpojLQe3tGOangPweN8zzx+g9dLlX+pqG3DcqItDRdTf1+6Nsx2
4qM+y/72wEWZPUuitsHVtNkElHjAd25G6dmp0bfZbmx9Lp4wCeOlPHigS3Zln0wD
vgu0HaYH3OvFsF/R12+aBrsXsqs/D7BK8my3MyCqE33wAm5ToUTuhRAth4SB7MJn
rPQNN8rKUMaZD+MaTuiDBqKzrvCPq60p3ySYt9a6Z0yGxgoyqiuwCdR2GULqxflc
pqEei0DmXwoXEj4bkndw8xDbG98zRc/rWL599pX1hLEAxS9/MRyJanCj3vUoTlCV
KJI0mhw5ILu2Y6tOWJJhTHa37kIVdOPZ4EsgHVOr/cttJ9KTsAVUL/y4Ztwtf+11
kgz8DLrcHIxaTApCydm7BPBL/P9F8w1vMXWp+DyjDXza02pRrrnAmJ8fXetWRFyC
BZkvI+hC29wm1JhyuUnKLXB6N8+Iso92RjVIDCuw1AmggaURLG7R+oUFklm1LQvv
aa4uZILVvQ79izGM/q3xFxwqC+1FCUtE/H+kCEYYug946L06UPBK19RH4TpJPQ0k
r9sog8oC/fvee3ai60GNOhiIT35DsxqbZXfrB/Mg4K4uuWmglo1PFqTsVauS4fOw
tK9ejfM6z0AYS+sw34A5FflQsGWquo6pupacQ3GzBgzkUMmu1npIG3OgtJoOZGZy
nuWK/82c/3u0v04v8dmhmOwoMmLiiMqIT+/Kj6s4BhOk6lackKimEN8b1LT5z1jX
B176saFujfCOyMGjhochCrs6FyazE5nSBhP6cHdVm6acaZ79pqUUiT5ldZjyenm3
dJZfyY0EZHBun5N3tLsr4BozkyohYVGOerFnOgyZh29851+4aD4CAthQfcWzoCt5
BaB8cMur71m3uqF2iQmziF7z7OsaV7DA0jogKoWUL+zc0qR8zd+JwgDiGkJz/D5p
U9qy+rHUrtuvtVHs/j7ifUvX8/o3lltB2OB4MoiAAyB0Orwb1q1uNlonk5+jws0W
iM+6IcuSOxNFY7lDqIdGg4dfpKIE0TEzBUZvLW5lKZNpybxokUlI16EW4TRVBcPL
y0iasEeQ+uzV/ORBSi3j/F8fNKFaOmP089nh4eMJTIoNIgXLyqfK6LsCs5eCFaFn
FE7Y9yRuO91+ilzZ9sME6p5jl9D9sotcpXEZN2FqHa6LkeztJfLXmEvUJQlKB316
5F3x12wT4CU4HpehUtnDn4lM186rkfT781lz35ZGKd+lEKtpP448E/Fpbq0hY3kk
SAxdMzQrMV4CuWZMVpociMkZYnPRYI7S99jUAF8rzzs46Go3BY+KIgZ9OY9122iT
WOoOGgqlGJl5Rbc6GrLqPjd+wii+tEGnIVIb/1AHvjhmURhQVwctL3FggR03xIcB
vnfl9ZK/SGhpcGgCEnEpRhlYBYbzhJE+u2/LYWzGLeZ5d2oTYbOFBqUppwM6XESz
4VJqVWHY+cQv41kWnpvfz/VGcbBFeHZU0YTugY3MT2Arr50NE59K0zDVp5n586Z2
iQ61CT71te/XF7peY3a+GIbpw6VCUMG/lgCtBVXJ9P5VqkoMDibMgZFqJyRIP1da
PE+bq0nbdIR58VFqXiUT8Ssw8LSBN7P2dkXCcvLtg079CRlL+K44PMrVDbPoC9NW
2CYcDJVVNnRas95wJkjjwpWUau81DVYWCk78VTjunti6/778CrPKSrYujnMOb0oj
rL9jGPEFbAhpIND76hoHTYKIcrYYTqBuQweHB8RKYr2W37yMSaJ7Id/Vby4Y1wpZ
l1mN+pplC0fU4rGnlyKNfNblabyUTpGbtjOJk4OJba496vI5acwLQp7L1ma1essZ
PobfArifZ5zYOOCCCafaKBaSLWCbxre3njmu799gb1t3ImAok4LykL/sklCoVhOP
NxsbV4V73cWbYfNe3MVNPmMBeOk4yvZzeuIXaguBAPiwdjSIAK56BtNLTaFTZTe/
/mBJo5M5vcmcP4i3L518xy1/Z0+DmbjZ1DMjB3O6lpz36FV5GINSHXJKpXBcfs9D
ujNwllKVUN/jJJKc7LVOogIFZ/GLTapAaUyYR/XodwDVVwvogI3IOtohC5fZDOyn
llZpkCVaSlBWJPjYgcOL1B7EYdoJRl7IiqRFcwlXXY8E2behfhD0ypuWbuE4EtuS
HnZrn7GwJfpZpaLIdj4r7rn5zUGtYNcsnmiseKRhBppwwhwTo0ihRHExH9dWiprZ
mxLHfvORqHyQzCiDETS5xUD/Vbmgg2douU9qYbYXs67YIy4YI7O8v3B28tj8ajsS
iGCurpXXF3nh6bWpGumj1mOuFMZSheMjRgh3CFJvEk4P+Fa9un397VLD1exkAXYt
Jis5QGDaOut9Kc6BvuIx9czW6Ge566wkmFsdkwjt60KEhKPcTprAtgGMZbG5TmUh
mkmVqtHE2rrF4f6DefbbNFsh29RjZunU5BPOEKhO/qqjtN4UQGrXpM7fhffu21hy
lGwfCGh1Sd0LBBCXKGelnhJNZRGticjPDQZMO6K8PKHTOBzH8T6rgiAOqUGq3x80
2aTRYpyQ20rspOhj3DOVpjYHyizKiklQ/M4cg38vCNgkodUdsAxEfJyxAPdogpxm
/W8LZUO2/AIBToVzJ6pB/yaaMbAcMzPTK7lQne33gZRzuBqDyy0K8SwP+bNBvkaD
4vIYL3ZcTR4+EpVmxpYmD2dNK5g7J5fQaX1MBfnulIyS7kzmwrPD068Kdv9LrL5X
Isp95W3f01aOhFmr+MZGXl47SEzSJTtZjs9wsoJmK/46IqfzcLSbbpKyGpeMWsTA
yRiu+i3MAAVY0va8+GjTZ7+rqRTQ3N3AJad0IySVYhSKClXaz56h+2r3PiEeL5eC
zQ/M3sQ1lhBBK0vYR+wHxV6HmqccJWAyg8eekhH7P3u6P2fpxBuBUXrgtuFzhbQW
CZmtKaih1eelkGHVnhU8U03DOnO9zHaPn/TufN2/u03TYgTC0u4o9aI0quFfg8s8
NcQieavLLlew2RR6bqdaEyymc1+TeJBXFiLQsfKYiJ5uUGcg/Y+vmFrcrYYOFgDW
/XQEW/BrDmlsct7RVULJuLC+TC8hR5s5A5hrjql/BM5ZjnEebz7RsSskT8awJu1B
XXT5h0sbAvTk7W2IX5XSsPXbQITg1rwSwI6uWRME4MG/QQCV+PkdykrZl9KaAg9Z
3V5+4L5QCPdN6QwzIQ5i2HtlYcl7DaFnIsFgbur10GpH1TKxDcrTQRe+iOymPsci
XFSAYl4/o6cTL0o3dC4ZHAJ3e2eywiVPadFdp9Cl2FQLgSUlg2no/zvZ60cu5aBX
F3malCqSAlSciOlcaRA4nZ6rvQXsw7qOzb8beaZorReXnY26kdzMrFPG92Gd+lwX
tg/dMEnTas9SNdBc7UMJ/EOQf0T0ebCVDsjLRBJDXuzqX2kI8PPt5I5GGw5iTg25
x2UJftpJwAZRc9nZSdQfI8rt0E4sq0vZMAY9x1RRFaetvwEOYL3bEoz7L3wGq4L+
GZKvvspmVfnpbG51wQIqXvd8ZKKnz1cNR0zA5kOU203OrkrsGbBqFi4eEjnvqBJI
CIxrQUwGx1Gf4zo0x6tYk7U+ejDOgWqkJ1ZvK6Ge6Esm4iWGnBF1CeeSoddw5PFR
QK1/lkFm923O27W4kBi+HwnazUzJEA92O7nxmTnhhg1jYbfYr/So3nL8LHqvARbb
KyJmXCiyWBzcalCBBfTkI8t9m0IztShdqJlGwogEb8dzSZ3o7eC9YYF08cFUJRCN
ebsL8wtu9m/vPQ/sR0avqEc+CvPndTLbej6pK0D2zgbjzqeGNcf/pLGYO0V/7vBk
M2zCBLFf07vouL9A0rrROlgkrAOKNlD68obZz3GzJZz4rOKuEhcCyRN4SaK8Ss/A
Ag2iRjJRdoju3bWXjyiWRK5haakhvrlws85tct4r+WRcq2fNCeSLgPrls9JfPt+y
x9aBjJhoFsGbuuQj6OtEt8tzvTAgo0JGE7O4hB2FJhWb0qGA9CkrKlAjjrjkRZZo
R7OC2mkc4fZ/LJIjcdCl8yZrerLN12kldPsDU7a9GtoBXtH3vVPKldZbOYCnuA8p
VSRptVz2uIfWl47SlgY9PHZfWjWEqzIWLRTLadZipz80XzoTl1UgaHXuGaPAr6IJ
eltK/Vx6aw5dwzhWuK9kS0w2eE1oTWXpW+es+P0G7agX6eqR6Xcl4DMjdq4Yyh/s
HllJfUpENp5J5oaeajFqd0LUHBtSX7CP3ulxeR5mOsgdvXNhGb081SIlcSvCa7Kf
IkzI1JQdnFTmGS0xunyu1CDq29f1ib5nFJFv2TOHeumAIejywlejGPiXHTk8pkkF
gyyHp1wCgaIvWtJsC4gV9ZaCOG8Lia8MWK3HqoYoDugoX2UdBTLGiuw0zaTgLWDm
3g3h53yKtO2xF00JJql2ouwFQUyhm6JT/Ujq96mKePo32B4f60Bk1vsiS9HTgBQZ
LUB97oW4g7U03PxCweCkPX6ZG0dYZJb8Vt9SMcijMJ8QfDelGWeD+F64FaGWD+Q5
Ow1coEvAYZb8r6M1jOXS0e3QcLfMxvD3IBOexlutqrgDJg58dGZS1rme4Nadr0ZA
ZbR1RO3JyieJI2Vnl5DBnc4IcKfhp2NCL+Gbe225FwZoTjyL8J6F0KZ3N3yGZEng
uvTKm95AqtyFvqLXqX8xAVpuwf9ApBlMxGQZBSuMT2ts/1cehgFKhJPFpF7fXa+g
BFqtIOlzPdLEdO8stOnUTvq6meKfoFlsDj3MYDa5ydYY1145VLGKcTURThnC+dwi
dSE13so1Q2ckpbZIoZsrg2aU9ZskffGaqIh3d/GF+0WgTGEXN+mBp7tCQJjl47hq
6Nf5/dh0pd1MBGfytLfIULsHtKV/8piwVgh4S2qNnd9R7gLn5FBr/7n8UrD1QXXN
Oyu2G/iUXIobVR24rqqlX9+2WMyLFkna/v4JLcfM/ht3qmIKTeBZbmGoxMQFWzOP
FP30VaYGTHzJvsphjy8b4cDl7Z9Y15V/Ue33vXCnp2njCKTrg3GspSict8wZu+UG
Wdg9UIDzr40i3jWpnIXyQ8IXMbNKoR4fDD4Jrtfbzyh/CfhlnycSn7+fVKFTWp7B
RQNnE+TEjYHAdmDf5+/1EiBjJ+FlFvrqLI2KZqWlwwAidx0i7yriDNaRBfCbiL+A
bmIn3odlhTp1CO80K9HTpw8fsdRB9XYjmhF14ybdLSBEkHGKmYEhIEz9ceUTzPdg
C6Jw9lMVenC5LR7lj2UZw/Kma7QLMeo3MZmWQv5gcL794apfghRbc+JeDw1T3id5
moxVruoLx8idyuUY4ioCzlJc/7UxmtsqxyWLSQFRj0WgMCVcVPFS3wt1w+fYUPoW
boePU/U0vA08MUI6z3k7S00AQ9zL2Z62qC6XlNB68EiUS8m/RuwHHn1CZRtTwr2S
tkplbgEstyLm2Wfk/Z3/XJw19gInXoIUw8aWdGaQW6Z0Cb3yO6T0TaZK9KunNOzl
pw9yd9PajbeA6v9bNsm6UvE0m+sSub1ZBiUVPHSzAinXrxMYj0PozlLCJC4dByXt
Du0JROcykZPkqamuts3i3OqZwGe2yiASFsEPpij55ckloWG98feeYDWHdWBbnGc2
JR37axum2CD2zXMsuNYEGBfNRrLWgnRwLyD/EVNu+eov3ntgi7//sDwuRnySB+J1
IJDjD45frpxuby5gARfGaAAUZplbX5F0EHIQrHwChEvMZsgd/dUVIjKSG9J/FS/H
xWcU3h3ASvnHyHOvRiiDQyyymzv7DXgGmGAXow5E5EkpDjZ2HCBbahd8WyV5grS2
ImTycANLnSqfYTwnrw2eTj0YBMR6Pp706ulZUyTMQMmh3dJXExxQhq+3rcNqOL9O
VxRofMD12JN3duEEjwqaX1XTGr/FoTyA356W+suA5JnFmHitOMJ7bCIWn/vgCV0C
g+bLfNk/cNt173mxfN3A39C2Zz3LqW4uYLoRccKJrhV8ibKL2A6ryE2OF1CoTFi9
SpPjPKrWXj27UEj63Njy7hP6j+VUoHieyHOYMNoekSRYCytqpDPWNHooJ8yFJDrA
Mtr/hAF6+OV9lTz2kbqQ2B88Rnb2Um0Q9iX7s2M92mxheNZ6rbxCFdDD6mz7L1Xu
qduZXx0LoFwNhVwu+gRLVhhj1R7OIfQC7rhn4/6UtdMGvvYpcm24Cs5K+jO8LaWo
bCOmdlUQpIM85KzWevNk9tBwBZTCDHYHzu/GxpuoZTs/M2Z/xyFYjzjJGHuwdS7V
korMLHlZetNAjYIeKcsocmMoQv9OIGtzOoKFab2yjA9Xwk9SYSgWjOJ2Wo3G6x4h
Y00t3ZUFkoEGafiAfABgLIeT95Q0pWbm1JklUcwdvWrqJbugZzxQ6mwsAsfzxTj9
EE77ptfk79bHM4FigJTqWZ1BIKi1vC78XS2KKdgf8KZ1Yk36GP2leL8eIh2aNLUW
N4l/yFZcds79jj6mjx6HPEIZK9udWUrdBTzU1Sm/mrlPoHoqyLFucgu1V4WofFz3
ZT9Q5/GuxkdsIxhE+9WQvUlLSdi7SWkQwFNrRD0ab0caZz0CxN2b00ViNMUuwlFG
zk3yaXXlPzCsM8dZE5/fe6UyRlum4tDKV6EnvroFj3otcH0NsrDbwHvmV+iLqgbM
CcctjCgNi+d3JD6uxlD+cz7HbWwqfJsFhNvwpV71RtO76H0B817BdG0QAgKgZcZi
ye3vZgZk4ihtJ8bl1mIYiln/9hwe7WWLQD1OXJvyUisxyT24GyHa0e6NspkWpSUw
buB0DOpAgLr9TBMDyTNscQwS8RT/xNtvWrTfV/4bawDW4jqe1h0Em7nZg14CVTHp
ab5GGxWEJ1Lr6uPyVP5ilSUEv/oVg4H6/pTMujzL7x/cQ1wjbZk2bZTUoOUpP4pd
ZT+tKgCI8JdC6LhOecJgIHDNzd9AjlEH+Rnafpj+JILe4oOZsrF6dYbc+ich5+/I
BtaRGWBw5dAsNZMlXTcB4RTI7EsZ4uLp1P+MS+D2IKn3cx7RiALfE9b6clvO2sW3
GQ65WAKHPH0aXsDk+DsIAd34YWjSV3Eef4J/SUj7PPnt4fePNFJlPDF4hx3sRsgf
k6s0JBpAm9N/fcaL1oCPwgLaFYwFZw3yCYBPT52//dR2+q4y4SiY6KnoGQ5jpDUA
VqjxuM2eb6jQMtLb83E1vnR+SgjMm89jo11lKE6MGub0E0KuSFas0N8/RQMAJWuN
BS2KvUvhAtQ0TueCi7HGXT7EVffcleHqaxzVaqx/0Uu7wGp+NsBcVCCkHxXtQ00O
1pYmcX8TlQi4tNzuR9BPNEmHJKtYZYwKg9i40hLsmryRTk65yKxm4oLpf9Qed7vt
q3W/2rK9SHCJ24l7aXP+p1CUzwkplDxY9Cm7mYRDEm4z7gLKShHtBsMhl1AZj/FN
VXas9UAaA3Dw0uB2K8YbmM/mT0PXDbzwLkPuQiWk58+lLGF8A/pXfwRZH9oe0Klb
xtaqLp8/MjlAUW2aQKamzDkVNACeKzEYdTutebbNyw/ie1HHEa/eZl6GD9RgIUSA
KAOwRKTEwropWB2DPK3dWoSCSweWCk+UM2HzK2QqjwqrcAo7ugFDXACiQoAWeCmP
tWCXIufW3jDEUldmMioW4g/aQWr7v+qCMs6rUYrlqFatoCkmc/H5jvwVJBUnBoTK
fUu2HUvx/l00rcn/tLoUgbgctxvDkuzTxfuEsQv3FP0x/wVp7mFYmJ9cwaVguDwE
gAsaRsHxM0HUPlX9U2jUPikOeJpuPZ81H+90NNxQnbs3VdQZEJ4vuuobObAaZVow
Dm0dCmBz7AplaOIGNr/CzUhdasoix4PWvJKcW03/VTewpOKog0hAr6V9mcXYogm1
4kMwSgPlTXbrPMH+eUzmrjeMu06xAf9OStOET12Tbk98ugs4jV4hVnaQLhDwmlCr
xsNcdM7LWGcvz5B1mVkq3tuh06kfpDQwNwncGCsAokQsAV8Roe9WZwEkZIVlUcA6
zA7KUEHIkXIG4IBfQkHxm5xoTNJfHJBzhDOv7IyqSlhBll6TFNMWxvJ0Aghm3RXf
PevZCuh6xvNwGK+1xh6+6dms8NETO4PSy1Fl6ZQwSG5RS26AyRz1qF6P7MF49g36
ixuMF6xN5VIoD7606YDBC2tC7XU5dsi+bXHM7QmOqnBcecnw8p0e7zF8jq4SLeo8
aZ9CvfjfZSAF+nb/yGnlhp5KvOVFpjKKUo1AUwN6P0UJkQ81ZewcdxK3tXJ1YVM0
EUauU21JpxSsUn+o9oPE6pzifSSchwp9DK1oi9O30OQ6QN6AB7hLsKQ7dsfjUC4i
TJyo4PjsvKwqQpsok+7i+vQgAFKD99K6ySe9p6K0KchGAUV2sa1HMtApxF8Nm2k4
k47GpwXcmQGtCSV+b/1eExE4of1y/aRBfhcy3z2y8gqN85wVXPr8lNY+etLgxQBm
KnsjNm9aWIBBdOCOlK3SIb0u6ZPrPy2NzY98siTtfYk+Hk32hC1lmMx1LGIyxYFu
HaotAg1hSwti+Z+sUnNOcpPLSOJ2XLWuZLtBClNPG4qUwufNKz4lunjvPqN60D43
eR4aFOzxOa5bypuHCnPNfPb8PWOKF299cFLDURQ2i4GDl0R7PruHYZF5J8Ts8vnI
KahMq833E1+ZzXuv2ZviJJf3P2inWdYHFK8KQHxSxozX71JibJmNINlmaTeuvqMQ
IOtRu/rOaF1AqllozZRG8z2c9mWQ5HgzDF9f1cRO2XMb5jUb2/a9bie8Ed9PfdQe
/RdNcCVJe1yh54NCV7L1kEAIq4+MUt+ficoSO+cw8x23U03kixG0wBtlrEbqgQFA
omBjdHj+HHqWexIQgngF36QDv1DY+aRoIRPrrrpFBRLvE/sg3f/l28HhKpy7eUyO
5wVXwE6777/hpWx9wXOaAs61+M9o/BJUtR8+hgjBr7sz7qY9h/XuUitdZSv6Gs4C
suIVDOFuzlg+ejOe6WEbP11384xOSyICb5otdM3ODuBRhPr2pHMWWgO8xYuELAIR
SGHP+Yy6ENB2AuSe+b80xCucfUhc9sBzS7S8R0EC61xYHyBweQjkjHsE+WepOUD6
AlaGgZXQmV0PSAXTlkq4OLbVMkrJUfkuz5uBzmSGEnvYRK+iej1cENU75mCw8sUP
moHnj5+BNWBakElnga2zQSo9jjygV0kqwiyIwZ9WHpCEZo6K0Dtl0FzHee5U3khZ
ttRe9AyVwCOYgJULm9gbDCPtDlbm3HgfQGjQMfVMIdAqROdsGyRqcEdr3i9JuBlM
4JMwMzEDkIiPrxOTcHkZfGa6CunTMnpvUoeGsv/c29M8/K6wZg6Q3ufv89MFCYAr
0P6tbU2ibeONblw7TqVvES/VpeqHHxq0QYAUZLY/yLJsOtawJrgkYVPQ120co7VI
8A25nUBM4gGfBk9clDepqBWW83X8XzmeNxAtrQWBCcz3mueDQnpF8qDOhasSDD34
hpFUBgMWKfUwgvR22b+Nhj7x56DaJyB6Lsqj238mgR0SyZJ97RlnZABIcB823O5y
/3gAO7z0Ucg6MLx8VRDS0q0eCzHN/ZGQPfo7GktBBiROTJYYz3cUM169cgpnzwJ7
BmZj1xUzbwhtj3Mvq9LSFNbAG7a9HZQH2fSTAFICwKLERDslk4uNEmQ2JukQS0Qh
TOx2UZcX1SJiT582ryLqxf+OHlJwIGbYiyAxRFs0Ejp5XTaPYytn2QYYu9w+T/2c
ko1xsvdNk13OFmXgw0+Ni4hGfWAlArUKUoRyoeh3JYLF/v2yOhXKNIHaZhN2lCCv
XPJ5RXQ1/hNotEJKQ1B1/nd74IyTCEEZkCNlqpBOZUrKcvP0U9beIR+oOHMKVwKG
qeoZKw64ojBBusb8LxT5oqWxyOyVvy9/M8yVH1YvzJ+KTL1hmzBSJxUEAOvYXjMo
dQxeaBvR0AQ/ReJpxn5hfonB3Ofw605rQfPS7Kn3pywMZrblYcEH500yUnc1AoTY
tUnpGyy4Q+Cno2P+RUxS5ttU0egR/dGbKawISh8ReVF92nrCTgjhOUrTUNirW3su
F2+N7d16IDHcu9/ge0kg/mzmQZxBvM9wOTKbnWapcjnIJ3O5VG/py8dkhkg1MNG9
hBM2Nt6x+xkLwH4356xmnFgZdEo4NRfHJtwjUQlPHtXP7UpKav/HhV0TC5fQhG9i
+QnbDnar5CJEhRCqAjaMkU0csElWwNxUfgG3Q0oTdNUpmAlWm68IheekI0dd8Oso
79W864M1WflmrDOyaLhSEy2erFGBUMpb5LJiduXptFXyK32agZzqQX2mUAZZSDfu
jL6c39Ub2E8EjtSZn/CqbY2xclHaANlpSPMJEAbkd79UkPjTJCukbu0vuKC/Jw3q
h1lzudGXsW/NPMwg0M3ZCYEvaQck6fTVR0VsWThuvy+WxXMHFZwnD6gqwdFpnF6i
waYf4+mYaVFLB4CqTo7HNUXTWWCxnf0pMuhvdnrarsVYVGPBSQ93E3pCKw+3J6Vb
kVoCR4rr9S81TFmpeSqVN8hm3amwJQy2zO21ZWotlj8hPcjMhVgHoeLEZldC0xd8
sK/jQQ/NrzSnXqIC4E4rXAoHZKEIauYSqb/wGHS6IPGG5G2PAnshmJ8RGara0Gi1
FaLvvY4qFK6scINBubfOpEtELVxt2MdTkXC83PcMh0jYVQ331hwbqvgGL/JT54oM
778mY3lh4TRoQIgqOB/zRUh3yJhPT7X/rzzZK6QK5QBe2OEifsT6ZHUMaRrKIssZ
cZGnnOn1vt5QnKt6hnt/9VFBX+3Py7DGbcwDCOvl2XTehzSbWliBxqWuJ+B5+ipK
C+7+mx4qvjno51SBOHf12AMrr3owL+I2cqCi3lZTuK2Iv/aQQDtRIizj4+PgTs7N
bvfEnySbZWoIGdCYYQFXyGQKOy3kuiu0br3tLMj032+Mc1469kHyvJsETcOwBN3u
D6lPFe7UQaTmM+ppyB5yBf1CTlfjnZWUafFkHK8lgZ28xl+AO/fCad0j4R24bV28
8cD+bdl6hOk/PeeRFOXh6qBHbjdWIDcmpIxh5AvEZ6sCjpcE/vQprgrDqoUkGDvO
nbfEt5/oRx440ERm2MOzCHQFpD7XrDrm17+3XvTwsIGYfQ3g9H+UYhsTb+0H6Agp
uT5N0tYktrIoBaE5M+JFWC6GuVajrgHu+0ccm0tMxu7Gu+8qfIajrrYmOiF/Mz35
Ry8UF/2T+Bgc/itmyBwr/B4HJAEqvvAmORajn+bB9iGv3QwmT3nbxkqesDYen35d
Chq/5xaD7RqyUuh14fVQQIU02b11qmYaRmcPb6VoSjmynpqZNb8Yk95MfzwjJVts
DMgYDvUEL+M7lL0flOp50fhjD9rSiKEuXeaTo0dU/CK88Hu/EJx3HUSSVIPp162p
oavRxJTgr7HQJzktKMfm/rKp+l5/BNEnnX7bh43+aAWUUjHbdHb2tyKyVLGnqUOV
T7ZK8gZFgMNIi33sGsuc5YYuDlJOtDdoYvWEwRP7M8frtOOFEsLY/aegP6zBbufb
i/qPgiA7EcIQSiczoYkgGkVdsa3wNaZQuVVkfjDplRnOjAm8SRpujbtiNukndHJN
+StSFLT9nWoGaAYZ8hHMwzHDIbcVQhesTJfV0lWUtIywZJ9vFcXnYouM6XzLzfPC
7djeBb/m9QX+DaLyxPCUN3hfSq1bwq1ZhNjmhGrL//Rk5fCcSXyXIANCy1GHBT56
vNzpQHAG/CEIflNtVPE+COOf2wA6O2kfEAtSmNS5mCpLjttKaV8MV2WZWRIB/l84
0wkaNJhCvV2ZKuFnvf0qCBhwNs1E6UHMmuY6iiZ555uIp3yVNKdbTD5IIeZt+G9o
5nrrq2fNL3bebRJDI1HF+6sKSqdXDVrqZDe1y4vNPpe75WvqAPPhBqrun0FqKz5q
zqMabSDlCmQfc+6rtDeke9x6eOYhQyy9wBWNd0+YeUpBMzyKbmecHw45oyrus/Ya
AMeddkIZXeB4jYFONmbrWnN/GeokVVzu652Yh/2De1w1seQO02eSw/bWndZVyfyz
nc9AVcNfBPcgjEm0Fxldyi3Bz1aXyI99DAeUGSgRZBamk7esr3Hgy1rEDYaC6bjy
ngxKZjUrlRBHxrmK/Qz4f9JT0HfMa6Q4Oom6ooJ/sGpe3f7yekzz2OX8t/PDCc31
3QaHMepiL2kTOgpC/ppome2geDOKuEW85SRsTrnl8BrGEpZ3kze4EowlkLVPO6aM
TBEiGVcNEE7Os/8PbmtNQgx/kQLbZ8Ljo44wPKVpDxiz6ulqUHzSi0IZcCQiNhSy
vzrU0kZUCf1MQMYl+dmUIiV2z/DSIn31zd7nnje143dz5KyXz5P6Vc3qx+KX+ed7
dU3GbQ+nqoR3tH+h4NM4LBMNTPn0jOu4/AKzinWq3e/5o8I1n7PB9T8SZTHL3VbC
f/hln5lOEHtlE71aYs655WJgno5yc4OJK6z5a5UbKOn91LyyYA3QKY6citUIRtNY
qNN9WKJR+bMfTwAtyYalCSgZi1kfuEV7RirzCzkuLYaXygLoQGpCfsoy3tw7z8kP
uy8MSd19Le3jMJ4G3W3Y0fdJf/mmwmoqR6YCZmfhCBWDw8l+5XRAgFjNA3Xou0O/
wFuHdVMmSRMNw2N4kXmGuW6nnfEGqvaYjbRlTtWgsX3U9+ljxiSJbsZi3kMxdLWm
Xp8dyZqpLV5ahCq8QQkmLAOYkudcs2l4DJ4DcbiBiZBd7fuxsLskxju4nhYRxPgH
4yMvdxqN88gYcIEKg0StssCZiFA7EElDt0QnRQ5YBAxYbcJMNEkQemw2CK1wPBr4
kCWDSOGawnLs/8FljtPvGK2mhO09N16rtlRGsFaqvSF1b9MyQrm2zqLCjLNDaL4s
7/a0ZwwqIIk7sDaD6d9XAWJTqXT9T9IBLbOnMa5W0n03xPj4tlA7xGP1M/gqlDgy
g8vuiwA/S10cEURQG9DFydD+f/XLUEmiXeGEhs67LIIU90iDWG9Njjh3TBtutpZQ
Aej2SteocnyIJaqXrp02JPGf97eojXL0pjHR41Odd0r8RkhScSomqpH9RJLfPpXW
D0XhXF/vH7MwOUoK8KHy1GJlK0tGlh+418jNr+Z3IQMQb6DAYVzIh1S6U3c2xlNZ
iDykhVA8ACkodZWqfVbLHdcW7kjky/2prXXSReGhuEXlQJSxJovyZeAkz3nhX9Z8
oMPT8iAL9C432qJ6bdWHO6/IwmCFlRO6z7irIvTK6MTW2H7pef7XiznrVOC9t0EH
EFLHmeVx7EX5Ng5ZNwvmI1oXMGv2e/y6gboTJ3Px63k446ZwarjCV9gYBA9ufN+l
KHz+/dLPnBxi18KQfut9UDhPF2nIfLrUxA7MkabvfOmGjTMhKZcnnbd9nmPD3dTB
M2r675gyshrz7+Ki+oR53bQQcwNVGFYvQ7SKcHtDUzs9WW95NYUxNFqcZPG+06Pu
Y9dBfYKvA5licmwQyLuadbIhg751GWHWG+xz3JDXFg0Evi5Uqxu4EgI8Q4IED3iR
pdq2rts2+ShXaWbW//qY7LCdA+OmXNAeY7PQeJs/1cqFAz5jrS1fkh1pLo1YGD6w
hguQm5Hr0+9cllMUzsMMJ1J7+J6G9TGUA3IHDgzYD1dObvR04PePri9DJSqWhhxQ
ViGEHpuvBaRH3RMW/7HFQIFaUfYoQdKFW06pB1Z6uurWuA59SYA3LlxXs15TjU5k
Ylt1ID4ri6ajMaUGJHNq6PVNWo1VK2CfGWq/oRc9dYP0iNNYxwOVyami2OqoIiXk
4y+YBuK36t4jlOIONiVP+yyI4NHcjAdeSgMTkliqpxCnymWySLjZKOv4sR1kKPPC
RiBGskDPL3dIWPL1n9PZBda3k73ln69RQOWwQLLrZojc/KuqWWKDlQnXLqhechXM
7GZPGyD0diO4BKSoWDZ0NY9SpeDzrRA8r2VTDG5Rreus0teXR+oCGbaFw7ju/IgA
j3FYxhKTSUNYde/35fsqH1ZzuKxNH0mCJ3VQReMNXGYbJk1gVjCFzHblQNBDuirV
soZaEYeWTCfJtiLrR5vVqnUS3TB9qevP1p27IKVQcVT/ZeCtR/lcTcLavetiVjq8
OC2nOCA2tdid/QsTqppTQxoQoKvK2Qh2AcHUzfVSEgHMFp/2yc9HhtDn4s1EkQBm
Wx0ekBe/8ox2wNIC6xmWa8bI7MXP55jB4Nq5LXuCO/c+TfuaF3N4ojD4egdutLXm
5vj4g7Qf3q5/WEhFaVPbykx32YSS5eoLKYNbUEDubXBwCRS1PQQV5yjWrYnqJDTr
e4wxZ8E+xymroOdH2WDowLepZgnvYZF4i3vFYck+D+ydJnU6aH3/qOmu/mr3GPeB
HlMIALqn03gECAyOiFvB15awqWo2mWdKvfr8m3yNmJJ/x2rmuwKYFagop7BNwqd5
IMVS7EaBGVDeq6lub9pRPiLEMDJXTxydctkqnXiodh3MfCQNd76l6rWuMj1p9zPd
FZmACDBl2GkhhVeHJzu93aZTA389Ys05xPZ87jRJnMiSz8XlWAV87HQRVKef0Ks4
LpmOD70oqYU7smwOnvgSV78DHRHNHI6ueRn91FAFkHioMDM57VJ2H6ToyCvt7mBy
ixL/6yJW7jO/GH2dWp0iaYQPpuq3M8DtMLi7W8GipV7kudVHHrqZQ+Hh/1ruQ1s0
iWvnQva2I3kqfGDjfSSkg+gPou3DcLAn4VX1NDm5JbIKbAoSMrgpZfByTSIO4nS7
+IUwnAHXl6DEFS5+ePGPY81kQaP77m02O60oFqq1GsDHXJ2gqh4hHX6DKhwrsIzl
yCDGulI8JSPdDRgu4iqlkVsWzdGwAktkxRts0oKqRvE4N6zV99QhvHYtHUsVmoSv
Zq3w3Lhk4vEduksplXNtz+jbvUtAxvWZw6OFLmMkkqFdoUYHOfoI5utjVVnE9z1m
MneL6cv3GCz8YweRkKJtggDCdVoOmO6DeqxaT3gCUiqywekgetNGu9nSLIDNZVS9
PXUQz6WVN2ylVdtDVfB9w1D+1EYmX+PiT2RadhpK7AAiV9wNq+RFf+yaDG0QWJhr
4gejNJ2OhhOcODfuP6Z/16L9NHeurMc40LvKebi41aAFZKXy4UzfDn5L0OXnsljE
hM1XA/1gZ9f1oWq2CnzpE5LHiErI5x5PeQ62OJFAjKnPR754kou+AaMZZNIu9Jg6
oeljFCIhCme2PYbD/mXeyBeZPblBucjEAXIFuqfYsmVWfQPl4vcjG8kDqc5onC3+
dRN0NebnY1dAvQF0/EV/8mSR+f/IMfbBhjxmipwL4OTuMifa1tAW2sWIgTA1xN+v
9yEA68XCR6/kZf/7Pz6qFS8NNcU1RtnBGBi0lStPkGRMNJIQHMcBw1H6or0KRZcV
2hT0gdAyEg/uJLWfTpxFF1x/2hcEoathM30B1hQk+y99k6JyxBimnKQknNYqKyeE
z3wuVivRT1XU5yaxyJIrZ219OIXxFsr76KwubKGxrbt5PzA1FTMug0TuiS7Kwdap
a456FGs8VkWUnSXYETwsxWg5VL1JNxyNaarc3+Ij6Wq98bvaNGRi0LDIN95qHBAE
t/WRt0in/Hl6Z7ejKXf+5kiufeBCedNNoXP51Su3JXqpwZwgvcZ4d3G6AUt7fBt3
fi6H+4/C52FKeQv/UwNHjCqSNXnj35US9pbFmuQZPfv7dyOWjxaGLMJ3NGwQv2vQ
hrdlDkeZu9bCwufPyZgoKVY8XDVpOSz2jeSPLNdFwvA9/hjgyC1AKr1cjLk0wp7q
sSx3RN/hT1ArYpW/u1lIS8zLacsWSrHBcjCPNcTrnotUn/1zDqEuVldPZWbIozff
lShfLlGO1GFPEeRUvZlsfPDdsFqfPng7qGTERcJ59kZojDkOEzT1Fv3XtNVYkVGS
p6jY7WkjSoTI1/q5LRCoQunPGCp6n3pXKrAlMV20cqn3xRt9b1stZwy9ETceRdqf
2Uyy9tUOGAJk0OHfiFrtIcUG2jfNMslnKz4wMWOi0SVBs4dzzUvd9x56EMRvTTA+
3B0rhohvFPa5vFSIHzUrxjAb+rTChDxQU/sgaT6d7cUcapHWkU+pAcpCwUYpOcgQ
9vwDlLM6JNtRCIoPUxZjz4oWXugbiBItenZsaogqoKmD4+EoBOtrS+Cm9AURwtQd
YLralF7voe/9XS+xwWoj830qDg3n11PJ850w4LyGB01+1KNwHOvjcX8uj7XH1PAy
QMhRHm7T9IcOo/nUlMFKtYMwTvnblbnPvr8ToszhjfQ54q7im9iQxrENbwHerK6Q
lmFDv6awu3k7Odw1jQsWOUz022M04EC2yHLTfF9uTiw/VF3FrbtpXfxe5L1lf8po
H27Mg6p4IWnSXf+686OWDxNApPGuyc2UDWj65jf8wCXMJp24UUHMIgK7kll0TXPq
aEiiLRoxKdfF9Y9lqRWRzpPDXvOJeQL0asgYEG6X1xOsvgcXMrKBQO5ZuewN9qeg
fMA3UGJHgYT3va7gfjq29AjjgkVT4kSmbEQxWp5g1xyLref/0T65TypAtO8jYep9
cBGI4gmhBGgBwf/glP/OBDVdu3C8ibh+BXLq0pMOIpYCd+bZnmeHjtSeCQZRHBsj
aeotvpqRQK4rfkBoNp0Ha7a2PORu66f0p6fRU6mzLXLiawMeAvT1jE22d6f7L17c
D85cJBO/JOyTsmL09B1b2Dhg3uAJy0zOrMxhtTPq2c/usF4czrVRF/ov1GfJlRJN
J5df/ECPlxha6Q0NFqUBUs1xF5UO9wKXycWyIbvt0xqEN8QpQYnsFp5QJ7b87SJm
KLF9MzbHG0WNh0UtJgOYT6aKacGiugSWaxrmJpBrs0BQrpCZJ5BmK1nZc98Q+2dg
DdC/QxE2qxiEM6v5YlmYZh2icJm8V8hHI3pnH3V0f9kkFjE7qY81lrCs68tRv2Ld
arERPFKGoUpGd1n8h1virzAXNDDtAC8FZUWmMyFHcM4f/xP+thwSEqbwzdPXIbWa
8h3SFbJ6jCoHaXXJWCNrn0DzpG17kVmh6yoUmyhn3GPGD3expI2e+2CisQEV2Yxe
iv7684Tt5YeRrumTRxUpcUd8xUmJotA2js2yslNWcYhrk+1CxqZmJ6PqP3G75ZGd
e4yRzhT75iOd+jF4f5T2GPJSCGPf+7msLGtI75sTyXm5zeSQoutkotIkAej7o5IA
jJeS6L94/mJ+P5jVDiAgauz+nLjh9mS2Z1qWC04zUB+C5niotOIf0sE/d7/2kgQ8
fQ/AykHarSmtQ51MGvu8wMJ3eMZyItTjP6iRCGvwvSlUQkJxlNmWB9NZ6/zHWMgH
M2CmqFx9HtBFnlrdT494EcIAcsk0+wLfyyKncwu327U1eAK7K9r6ySxJeUheuX79
Pn5rPsWACG5FkHCRj2y0zFjG0TVJBwNg/Agj7Ont+auYGSz96uQsjF4Jcz3tI8Or
lkKO9sCgpBeQ3uKRV5UqV03ECPuggpmCsps8cmK9PfJGt9/4RhkAF5+vXcVZZ0Fu
xfhZKLRAYw1UH8R3usSZLKVCXTGIlak6rC4LK5dEDDEtHLuzkLKe6fM4uZbPrC66
GMP/gAVJ9dmA5gZBkKAJogkCQWZtKVfpVKhXRpu+FWr3wiO65lpGmh14WeBM7jJn
b8azR+WYgbeCfbJ9Rm3CFO08uYaO09YGoO8BDwh2wZ/rc7b0RHhlTuq+EEFndZ50
QSvOV5qNHnvZaJ1E16FkwA+o4xZ+99ycsMGrbNcQL0hyk7jCAAk1Aq6E29b7Lrq8
S7JDs+Aov64hPyzhFTgKBMRfUrAmDYxz2vqt4EPOZ067rnw5teT/k48ewuyjAu6r
NotpP2GDB+jo6kLSzD0K53HHl2t06NKtcdQi7uF5kLNE3i3UhXRiH4W7WDxXiHC3
PQ00dp+xBIG7zxCndFH4TztvVm37ozJ5x01HdSFI85cIFBlqnDmcT+lc8Ya6bIaw
eBWWSci+/k7HmijSA29hZIIr6detQ/MgHwIn4tM+z+cm0pEMNAbRdw0VX4kfeJSK
91S3xcaKVrxah3RAlUzjAiw+vXxYOl1dTRH2dzWyL4DsZfh7tPO5L0RCNXqhtiAC
sgqf6NWpXoc8i4JAqQDDeNqzhKo5T7Ke3wkwWHPCZyPR2eoyN++YVBcO16b21kD+
e5EDuQq3hnWDmDvKq3B/yQ85wQg/9xHjZyRFqFru1M6FGyhEOBAAUSYU8q4uzzt1
eoQjMsAu+f0PwSXAD79xF+2qeRTPWcwEW+Qdr+AEqN004Z2fekwr1lTxKtWfc4cc
iZptvKh2YxUBet85Vw1ueHFZjlsX+QOMjCKZwCI3L4xkAuUIo75D3FGQAFxK+cbD
a03QTe8FVJHTtux1CgeoL+HQfH0DzhDNRi16I44kTMa4FjtHDow48d+wczCGcqzy
bvEq3s72/b9lOj0t7v1rCmdiMkxvLv7jNtCPLO8+UzgQrYzZrA9/AlwvLidDBQeu
V0jb8JfuMfyqCTvWon+P5On+v5DtqcdRdNPD2rihkYot9rajnsG6UnKq5G8gIRe7
OQogeeadS29qM50g3o/mq9YAnj45PF3wvjXiixhsQPN/ok1Y7wololy7eYbsMnlc
4D3rRUbIwhpKpJySe7S//L1nRlkYQI3YL5IQBkbJRJgT5Apo5ofgc+cS5BMP21OE
yQLvDjcGbJRbz1l5gCtUGqryBl78d9941jPx52NUeBgdliU+GTsPgTKZbn834xWu
DtMEJCWQEiqGzm4Z3MZwZqbmlhJVbOobU94FX4bpUCpNX4HnJZpSdWyx2aI07MmE
pnzrSiEIiYJFfm/ETBDewk4ZXq9gdLRlfEhNH/jSldhQMk1OnVUAC1wIdGIpVnKx
lS0H4JkDKiaWWc5ea02HWndIRNt+uvF84m8XyErkLOzT20dj35qi73+VOAnRKVK/
licaCOMkQWYqTeoKJPMqJWGI/sVYVHKtORTVWTLbnYoc9igKqNczBk9SN9hmKmGe
PcV+xgx1vKigIpxRAYuCICUFavIOA6uRD9Us6gDm9bLlkjEqXmLRTOa3cmcZOFog
32CuvD21aLVhYMETtvSmd5PB05XDlHkHe297am3RIPz3F/hu3FP2Jmak8Lge7ReZ
f/j3dbX6vyZbVGBb3SiML+G/1Ga7FzZK6gQtLvMYq97Vui5LztksZWjadxROAQWc
3LysdtxAnIraE1+QiIxPjKZSFPY+Ck39YBLiOtSWMLnbwTso5AQMz9Ui5i1E/b0Z
Aqn2uIp822m6srKUQ9SSphq4YGBxeybUT+9xbnKcUnMV0++f1nDTRNV3V6R5HqeV
f9zXGcRS2FSLs34i6R2c16YfEDMLvW+3kNplrSoz6l1DhJYO8WqPqrlVW1gkmW48
GLAK78JjDegvjWMCTAI9PlbkVd0z1okedn+gfa4h2ivgygDR2Y7eWW+bskircDmn
DcIq7QOB6psWj9BFq8VRsl3A0SFUZyXWHozxUfNttAIgKFSrDUnSSmBgE6IucbhH
lCQQN1I4vod1e50/YekyJpJsflRRMPXwZ0aXBt3drlum9xaB7Kq+Hr5Edd85jTu6
jVCme2aoU4SFeM2GZhWq4tdhPRSBmThlmGdCW1IeppIcmm+6tPqd6QLNA6d1wuQb
b0u69wCxLEIzbQkNmf4AYadakKTu8n66WwnRjO85Rgh2dr9MyV0wZXGeZAsiJR8a
VjA/cizTBGq5rFjWLH/G+B7M7tYY9Z6vXCQXxkZISqPYn5CWVdqoUHPB+OtX38Wb
+g3GXU5sOXkrWW9BJZLjYnG8iCCRKC787nh0AcVZcaQ0qWpiMZf+Joa5mXq0HpM+
EUUPLaqhInWmsbQtNd4eOLfYkwhWFvBICWubp1MXHgEGKJQVkcb71w6U04n27bXt
NZIU5GDvOO/dfe9KIFFgg8REsrJaQYCWYfFH7fXOoOHNQbGEHLk9G55KLsWiYYSR
pS+Yd5EcmQUdn9U5LPNUACHMVNBNbcYxdWwGzcgN4vEhHOndesxUWlaCS4I+M1wB
a2tPzUgMkm3xTFvicE7Fx3MYPv45+RLLFINgGiST7kDbOdnk+MT0T/S0GOa4iIsl
dv/uBPjndv6D+pe4Eofy/FeAmwKsfDilAETPeGnShUizMppZGQluxTVs4NKx54GF
1IU8xB1etRgJju+1mfjcp0EP02OJIfQIhkBmLpiVHHm70lcYykIbvkOW2NdWUIxW
My74xnVEnQy0CZ2UP2LKbGZykJg/s0mRx+8G6FK+Hv15f+Y0k/W0z7U5EdTpEh31
0NNaF1ozl9b8Bt06X+FDeZ8IC4BfBJVCSVtHMm3Pw8wsHGs759vlFbWA8nA3J2R+
owN9FRpDyy1w9fvQv5PD/lXIy7PuCkcYyedU5/QIzOu5jNicN59RnsIpRFzaNZ9m
S7hIxMGoyBkiVhw/VNLa2Z1GzzZE8/nuZURfGXUmtqaew1z51kcl/yI4X26Y42k8
QaRIFu7FbQ/h9Z4y3tecxrW1Rw/sY0FeGFCueczv80Z8dd+4eHGvcQzUl+GKEMLB
SryCLDGAjRujhc1D8xYH+TzmIeC8cuf/U3QD0UEReYyx1GuTNidJbJIEld5tlfJU
I3MDYyq0r/JMYa+/wEePf3cG8DYIpMbMMg3QJFU25kkBnhtUJdsaJyBLT36sG9fj
mup7frEp16I/iIjZklgB72GvGEo8MZpovOeseZAKJSoyIa5HqVewG2T3hGV9YPjb
kR0urZsVI6IHMftNbqoQL9rznjHlfNnx7Y8i9Xg8oqLu8YZ4/gXMcTwV0IkXsr2C
0PbXFd05osVjGDaYznRS+dFdRrD4L4nYYf2c2RIbVNk5bSTt0FmBGKsnF6nQ6J4E
fEcEtLgL9CmbK36Pighbp2p4TvXClWdcTqT2sze/OnF18jNumW3c1vDyst2QXrmk
fsBLGKfK4n2MnPlOEVDcVgTscC6ZaXr3gJ8cXvjtTZAKrCQpZRRQm+5EB2n/0Vj9
tAkAJLxQCBSTFU9S9UCJ90/aYfHgXQf+dZ72vzT4d3Ft/oY7SQKQLaEXHuctFl4q
laT0265rv8z2WpyxwW/huNWpKMWivOtpjLPrbe6SLcG83QAtX7vY28WNACSIHnx2
NppdVGugpXDDakpy8lF8GL8FzIL0OrIXBpSWyEyxRBCxthuwcp1YQVslQbODouAJ
d6QBmooiVqDqtpYyQv3OklOee8SZ2IMIUikElaOq5F0dNQ9Gx904Ye4JubGJl7r/
l1WrKkWwVWFtDdoht5+IrtmwmqtR39BRYcdBCdHKuc8m1PFV4Q+d/AWPg0IQNS4v
ybaeKLNNtVeaJv02ncZWKpdkJtAEX32ikHmL4HsEIe7At8Viieu8TUu/aqJ6EXMz
QGKKzPFTHDG9uEYnMLs7ZarAX6W2iv4uf1+jwK2AhM7dSIogOuLMHwLGDQ3SbBq7
XOUm9VCfdMh2bnvSYirNl+UAAO6R4ywRjdVnnTOr/X4U/rURfcNMAquzAhHmGTj8
e3dqZA4tx80zI5VaGumnmy/xSXI3wcmOQzagneT0bInBFll1NsmisggHwuDcGr7F
mlefmfyY/rSiPEZUmM+BkIFp1LlsCC7233sX4VYrSXbUu2yBreqGvLnnU+hayLh9
Xd6ZoFvr0mdPFmo7BE2GezTV1UCbjc5hAAR8c2/+gQcQaK4iaWgXPo6rrZPXGYgT
IlVZP1eKMwSc9J0NhF/5cN/W8wKkSMlM+Xp8PtDmCo3uXM+dmCBnr7/VpJxa84WK
hior4GvVpZvhyLoxRJSZ8BTmK7nTZ3vDc2gUepxa2s+DC84QxfZF9uKLQWZg7psh
Eib4pPRj3B9uD1FeoUPgkxSgF8bh7SImQTMLNTLVIge7yjYMT1hbQcfOivTlxENK
Zn51gTxPPTq8zIyE+zK3DXVkKj8Au9z/VzD4ZoftOBeAsrfd2z2JoVzEZkoTS6Ag
6Dd8F2h1ZhnF7fMwp0K6Ci8qZerjLkTmjGUHYPrE5NPvPF4kmqiPloDiSjJlRa9C
TZ24kde4ZfT/I3YnhcS9IO7BLHDAS68JFkVM56kG9cgriVskuU1wW/sEXQckioc1
aj0aZvbqtfWUwM55HLcHxPgfsQa6YzA5adzGKQKsYSRXx0yuBCnt9qzb87fp1QOX
UCV9HLlyWMiqS4aTr2FOpeesSt2fKu2Jcn+JaZc0YycXn+Jvr9gjWdohQfARK6bu
WSNprmYyEQZLdLdbEP2pPYSWBxD9jcrcu3Ty7TOAdrzq31u6tFRLywuB9H1ELXqY
p+wgY1rCjjIW21dMU+vKMf5hna34j9kDKTmRFOpEwtbtIjd8sZPqfCymz8+C22iZ
IOes4fWTFhpIrU6wdS2hycLOPDveJujyrW/UWsj4m27EyJgzbOnwu8RTckEoy8w7
cKxVIeAlYS8n7IK2kjrTW3T2qhWMZhSKpioXDpPGVFh9Y+r5YzQSN8ZdwwXvDskv
G9FR2RV0yrLTc4N9EmxXdshJT7CQiuSfEqihoMpMcOJKhoT3tQWkmEh/OAN0hBmr
i4+HJkxQfAe5eQYmjp+ie0dOFTtGD6cvyNxfgGwwSAH5OKZF0v8bTwv8RF2PRkIO
u7B2NzlZBcHM6QfHJLq48vvmmmh5jHbdeFn8CXnAI0ZsLkTg/gv5nEJOURkHPGkj
rCuKUma86dAaxNC+Df2pZYT/hkVd2vkerN2mGGQ/rGTPSIxtCUncGZ7kFme2oZ33
VO+aG/VRjWu7Va0/AON7Uknfsi5VLNotXnICwq1LpqLx64QFfi0OvL4wOkcfQ0HC
U8O8mxsMaHsWUKROFuhab+1wv9fOc2DbhE4GA3GpdlR5AdSa4Qn7ZUhE/I+E5yxw
F1MvqOm6Rl8NE7dM328nygw/sEOpK+EPqnMsGYRw+jNgEWIgXj5P+M0hdtjM7i8k
SMXpJTjSrv4bjZux9ClzdZNGWBo3YcuiVvuKWNkj1gar5zhVxYEdpLroN6mT9Gss
lJS0s68kcIsg98GUFwVEXpoYthYd8cYtjsNH2VgbgjKLIxpPqlaHVKLhQqfgIRHx
fzs9zHTgdr0mmq0In7ZZQz5UTBR7aWFEBM66HnkSXC8qiriWFwj23i/ahHnOfHUK
hopm6ijXbMGdpQXOyjUPrOwnl/9CU+1PaXC/d98HWixDe1mZu9hIH2dOtoegjU4a
RIB6XeaqKm94D8dujEgZjWKKQK/mTwOsLpWY3bLwtWS93k4coLWm427SKyDFhb+y
+d4cKWdIVwnjOwz0it3WxhHKxyeQntZg2rLkoSyG4yhD23TUEgDpBKjh9G/+UvR5
I0/1Wlfh0qub9OHLL4kRwEOHMCvLgUkWcyw31FQIQ6LoZbEtg3R5QQ/HUkFHXisy
Bp2o0AmdC7tmMDMLUNk+shaQu3VldfTgmgssDDha5awW+EWnvMx+b5YowRfwB0ku
OSeCJoRWql+X5c556B0OQzL4PcCLoS/R/roybxGlKSrEA9kAoK7p9pbpLXrELiO4
RhbaiW+0Zzl2JY+Nv8AjizATQ91pYItl+ytkJbdQ4fgmOy3hqDxsS47MQUCIu4/S
yxLTcRa8LBVkLocsJoaNM1uWNQ4h5CVNoUMyS3xzpx+ICUZchfZPWD12/1QvHJrS
+tJwftx6jr1rttLpQm+5VHMBsOCNksPIWbZuoY5VnnL6dDAaxOmkpdiQR2UiUZjk
HX1+RvFGOlt6DURN8XS44N0Ax05bMIXhB5tVxKuJwVBTu5xxpXpYvyaJ/EkS2T6P
Iz9VvA4iaH7oOvD8H3bsFE/YKpHXpWQHCYM6ChnjBF6QK42hx1dSZu3ZznHybady
VA9OmRicpIzb3EHklsKEdXNdgt0mVLN0+5mi9f2XAuo0rD+TPiCmkuF2ptm2KOcf
SYXOs59ocRfWiYyifLPfe3xJHGoB2iaVxLngn2p7yAVd6ulLDa0ZqEtclg5RVnw1
3QL3DepcE/JV1hlpwsmRI+zGfsb3gnT3k0yoIyiA3ViewlmKizt0aOUobwJYUDZ4
uSkMJE8cAz1qDQTj/m5CiUCULmuQT91OjCw/6hvdRTaQVUSj3TN9R7xsLc1s1jjO
dEraGyhTjrIOXbA31jnKCoC8Llq9TLGEgsp6JqVjNryo8E0gC5esW44C1c0DZ+Fz
ROYR0F/jMDQAjntpjhj1O6nUYlN5n0Qa/Sk7dMFdvq8dyJ8DZktA4ksABycrhzpZ
x1424fVCxOMPmBxGXwMn3xkPXyVUj00AvSe55AzC/WFbeHzgSgJaoqhj0NbuNHK8
xykemizBXvT9COKoydMcHZSaH6S0Si+JZ6BUGajW/MGICCrxD3FiVWaYMxERhzPD
QNJE2ptOu6GGEazuZUD3RD56PlfWqeEgkv7EiJxCvGxrJfy+Rn0cZCBlzVESzFVY
f0Wwf5N+CPM52csuUFogr7T0AzH4Ioze6VIhrgmKqEnltduOjbRAT0bMnq61Uwng
3CcVvQnVxdHr0fJGi4sO2XD5C4SuSEyeig3QOS8RKJcgbnQsKQr9GSvur0c+ftIa
43t6QiqQwxTFKPpqgos36X2tRr9tm195XS8O9HNJ9NtsZOLH4IOqUYAPDhceCXhJ
2JJ6nl3DMW7xsFYs41iiLejD2h8eCOJr67/nPZrx+yKWjemh3MnOCY6n44o3h9c7
z9hIvBY2GMQ+P7xG8rVbq5v64jDdVWh0n60vMXNetsWRBP10e+8BYmLBjGYTJ6hN
wfDwGcfpSmVgVDumHToPfomhAi/AiNhGXkfuiUxncJPxMnqbJIkcnH/IP4bUA+Vr
hP8VdSY97bUeGGiPMywisBJhyzyttXkQ0doKUwwZMHAB/oa+nNm8OZ2eReRhONIE
Zxs9N68+ZEIP7iKm9ALTM4LQcgPoI7AraEWBoCMjAbYms6xnZ0HL/z2XV+v1kU/5
yiVIrdhES9jJkDUnOyL1k4UfB8ASLDwbUIJwRjp/bA1wYiCM02y2t1n8Lclse0F8
wvwQw1odsI5K89Ia/VeSCQbiFII9k4z3nxOyWGHxDzst+AXIzLByjSmxaurDqVuz
rL4pYlJsUvQN3FN0BPyh6y+nWLGgr7KOWKvHzhT0zp2I1hhA7ODe38i+l1IQr8Ln
gXKhdiO1WHNPQ83+8wyuWNrR1G4UHuucnLFGMmchoLyR74PYGTaPQWTNCOWL49xB
4eV+AG18EAyZWadJWBydmTZn5ixR8oo9y/s/2J2WNQFMdU/XPs4J7Hnn83BzUHJH
iIQhaHcnEK6/AQyIHd0xkZW2HfPPczywwkCnogCML2OEV8jHlUpxmFNrRa6+P71H
fwM73UmS9+QpTHtY32MByUApgyz+8Q8lNoUANnuiQ1ID5A5cHXs7nqsdXVGsTdF4
Fm7N6bq2xKF4HVxl75Uky6vDGKWIPmXc+GlBAkmqoWUpuGe3V0/7HioZMssWxiKT
1LsN58m+2TbbP1A7LrR7B5nyaKcVOI5p9IQmdeWASkk+1aZoWLwMdBp4cRt2jKih
sCTJRN+Qqym2E1TFFDEg5OAJn0TPEE3KwbRamTjmUqeVMaRDdRRgWh2DAqeewJB6
RnDSsBDnKXWIueSzOt0ccqNhx56y0+CfKmKyoKm0zdxTyXzTu7cxyxtOtCVEYaJ5
InAN/ZEBYh9uHymv10XE3Q7fdkTd8Nt6zpGJJ4B9K8jnCyMuFdjqLt3sRMGsODac
EHLhduZfzRAvvptGF4Mv09ogz9mCaK8APBLVwQ59s0WPHa2UHK9F5ch+ZgrlPBkb
BOVj6u5wDAnJTFVx+UI+L71FoF0Ix5RyG+gd+3isD6QVMPanmEK6qketSuXszVXi
XtdRBcHaCtlidiSyQ4FGxhyL5O879TpAMvy/+5zV5B+xY3gxFdWrV5Lxy+zd2NNw
SDje+0zJEJkBFkmzMBHFetuMU/x5KLthYK8LiwHS0JVdzHAZUei/y+/155k9nmU3
Z+OctGeviLGc7AUlvDtdZP9jzFvgtF3JoJnF2LqudOswv+aDrs5Xhk2kUKJWyI2b
+Aiqh6fLw/ICdG1ul7aZW4n6zr20eP2086QfM2IzdxgP9QijikE7Vozuf4KdpmWS
FgWGE70Oa00QDGKPZdatJlhrpWtGXjW+mrkZTRgp6snt04/DyAENP5eYwqQ82qFa
RzP5f3DMF5DrpMPan+NpPTQPG4MlDrnxrZNIzW1ayhleekvQbDdgKFvh6BDeVHDG
JuG0lfXb5Eb0JLTe2xalAI4MjrXGtRPLYiBIocjLe4JXt9S6zQlefafSH3AkpHJL
uIjDJ0FrfaQT4PLug+/V0HpYQzFPIkuJ6ipC3c6I3TFzmJDTpKjh+L+3Nw+e+suv
3ddG3aC2buO1+bTh6Yk2hsh//ztOZVOUKTWz+GFgjmdueorHc01IDEa5W2FOdiV8
33dXIG9DpZp9nwO0UkfTVWrla3Wz+D+seeGgeX78C1lnD3Kbvtj3+AyvTxb1QPTo
Uw+Maw+bZrJbSFgsYH1OAn/TkdG+iMtvShfVYLWv0GrX9hmA5+aFOqvBjSe3Aczm
2e2k1M+1/NlEtvjLGFUDoJ/F0i5pR+tPdKtZZpq4LMtkDIz/z9lqMe40NqNqgtwl
PMyYcDAh3aM5ze408sc+bChg///x/eMIdv311GNnQdfAR3xYn1Iyqg/kC0RaaLg+
9Y1L414X2sp8i06wSUaAmBRS7F9hPNrjkO9fAN4nxhl9Bos0Gtd3WOUXruP7FeKs
GHrparyRDqJFXMLJgUEM1phKMHmypFRKAzPfCe5V9zKgFgkW3NNK1yxgDZuZR0sv
/gocNeBapRaqccvwOFXSmjazA+3WxJQTYG13qeLctaXfyCcUYcV2qwCWuUaCkDiI
qV1mu2Q8x1NiuJBGX4SuYLn+oUYlN98N1M5poF6UQIjzy96qALpkA2XLR59sYJh6
b0+MzCOiAlebC4/CrfNP+vaA5kY10+tPixpUBlzvzKnazdhSv6eDNA2zsD4w2Bvm
pw1h8MXdl7SDjSRwmGnr/PVbVtscClV+bLjlLcZxFjgSlpyG22G2qsRgwFZq9eRY
jEllFJiKox90Y8QBj9ZxGzGjW72X/cN2rN4/wLbmS6MgSIkKCXKYsIrnjOXDjW1b
nh9z1Z0ZZPp+GTyBprIblicGwz39TtxJDI5yx7MDKOZn8xOLM6bdkND8PJWut3bS
1yQM5P0xPw3OklE3gVKV4POeO0SXoWUTD5LS4y+bLeayQAKLHPZ5Tu7NJONfZK3M
+t2ka9qnhyWtVj/OfwUwV0sK7svJykJPwrWRy1lUDyUzWIC+eq23lNwF8H/F0Jw4
cMe5Xt1SJysAN7VnXndVkrzXLSPD/x4qZSXLk3OwbSCPZQPAJs+MCyIUC+knNgfq
PN6fegKdQGpp+9pkCsfAqyPpS0esG4ZA0+yWTJ5JvqaCMIN/d32+l+NBQC16TcHv
+WKHXRqIgQbO0vtm1NuEBLVAtWJwIL9RshAEXIJCZWbYG2IzpBUf3ukxcf98Znkk
TrK6zU7lp8/O6j0btAXz8xHhMenDPrvyaGMCBYJHG2PZw25WsLiGMp648PtHEzc5
O3l7zQ589q7ZBj28uyNfYjyt+jBipK86+DqENeGVRjWfn2vmEPMElekcdqXrhw5b
qasS7nWuT28QWgB5JR8VY5ofShHufJuIF9af+3NPasj6uG2EGj1KKzAFRkJvuueL
eMUvKKg6brNJ+2rp/VQPQi34RU3b3ASF9yR+EjMPYPYCQbkshsCTrrDEgpg6Z+c+
ef7j6PUbAovpa7Kc108lquXVH1YX0owbn58gsoYUVq1+lmcHhmxF3SWsSaX+acbM
pYch3DCa+R2UD2MaU8W5spwdE+C1dJpvrf+YnB941TmElSe07FDHCkJsoTSbWfgB
XFO/IrkzCtKrcpUmsUlMBH8SiU1vwCaGBjjjVonh5DDpqpYt3LI3nft1tf6+I0OW
sND87N8Wxoi4olYPn9HPuRNCkwLybEtGEBDYvack907EH0dZNUCO1V4ckiy/S4KK
IEltIQiQUg6Q8Zv8QLwPWGmOh+9gE0+ZmBWtmx1PyXiBPBmF1jOzJ/9YY7Il1F2p
YfLP2aCizMsLeQ+ngVkM8Kwh9vAH/vuWOpOhE9CPFFTr0u3NEaK4vg/AWp3R2YO+
dRtFwKpw7IXxwhIqrhr+i0iaeSI8D83vGOmss0n2JX9fqbvbbNwff9LE9FeBLs8D
wstqd026flpd7dYRh+nDVVF+0UMIvIVJPE85nWrgDGGfmu5iwAfTuR31cEAMhfm7
RtWoX4P63D4VAkCGRL+Qh6UBtdyBVqdGj8ibd4tc2/VzMJxVgfrwInRcxeZKjsQW
H8Ol5M/xgpTF2/PU3f/X2BTud8GcNn952LTV55cGXFnnR/vQNkTAIYsrgN3m26PN
G+wYbHnjENOg9j1FKfuQBQRn5e7q1xqNKLfI7j+Zcm5LyYSbZ7K0QwIkal1dKM7a
G5UaPqqt7uitJjFR4XidOai3apr5B1N4xaoe3s0pSPRtN9aAFmnkYyCKwdYcb/oj
+9slj+nVI3ozxx1TykXfan2tJfhZegfeswv5ljgp5gvWY7rSWYP9gxn3Tf0D/1yD
h1KIlx/vuZgoEKVS0n3LuTis3SJueswY5717mBTlXTmx4oYrTLPHivebTdnqvjUM
gmamo4of9n+Idm4K/5+KxhWuqpxRqEqxStnCogUMp+IUzitmwQv44pHPWxr1VDT2
ec5JrjHNiVg+71GbRRQNS5htlLHmNbNZl+fF9qJD8OxScdH1YhxyaJ1fNDj0RUjA
BWL0DNj6Ep6u9cb5vAarAsXQjlICAbWqMPqklDOjF0ulYSxoNH1zwfBlMANA9gkr
iayq3iCQdJ1PFkiLEzEvKkMWCJHqhJBPtXI5IOZIaBWM1jAEJw+jqAKb6KKJHUG4
daKwCdLz19oz6hRlSo52V2XP1j+75qB/JXGWZhmQLfNKCPP23ak8n6vBUO6yDzfP
BQASafU1Wl+lhVAbiFZ7E1ElQRmzLLryFZywUOQSb2zcpfVpv8WCiWX3+fF13cLZ
xd7fz3iyo2qFxqUkuRzNB7yjOc3cPM5jCSHkvcdCAfMcgkdvr/oNcWRE4M9dchk8
sT60SRSqMUyWCm1V+ILg7FYaT01/CZ8CsoSxj1fxq8UM3dm3Qth3hNjDvHN7/rxq
6Dytc0VlaQj7npRc83DO2hFrXzHj9CE7TMP1uMK2hD7547Oii0DyvCeGoytf2dUW
wgoORcZnQobaNyz6o74g0Tcn78HUMTnuv9KSn91XNSQCxefvGj8WOAMHFNKvpzZV
HtYwU6ZiOEzJ2vczGHfyMn4Lkk14Xa6DB1AXl4bGw+sb7j9wLWw/1HYSXwzCcuXN
jz2aPAJvRqh1vadr3x0kY8UIvl5uqLPZNlHy+Bqxtm2VdlCr1fB8wasRIY7NRUR+
Yp3EQnZK0aEPXnYI2tBD/TgRsfiGvGnl1gdgPvh4onVziv066wZ3wWa1QUUfa1MM
LKm4BD9NrKlG3J4pDjP39Ao5qsyPFDi0IlTuOivOTpM1Uvftx2zok1A+59IQHVyr
fSbVXBqKvRUMQPUdZTQoZKVRKrZJnwe2tgsg/FiGg9PiK359zg0bauHrIa5UAQVa
M6oUCCWcU9pxGC0lmx2A1qjh3hxxZqMexHYF5HcwCo+2UqsTLmY0SMqV+hxBmxky
hIWRMRCAW1CPvTXHGwz4o9zSu541m56Rii1qeMIQz+0Tj8eYpk3xwjMm+3CrSNB6
9S8xjMqkE2li3r7T6ep60h6jio68yEV8BjUCYVsrBQ0LMb+bpFKOhzTEugIVTaY9
NQZwsFAsNZpRv//q/KeGy03SbGx/9xoo3KQWT1MwiM/FtBlaH4nLKG1yeT3baFFr
bfZmJCjpxTiphYPbkxo+YJAdlQ37X6vR69H1QEgOH+RWwIsRaEQop3yZJXo95uXm
hKwk9ocSzhK/eAZm1fXMOSkoqjGpSKJuSVpww5WshnmEmBRfhd+hDljiP2OFRVfn
y2Qok5dMW98w0fMlDkAJB+9nymvD1GB1dD6HTa64gnjAL5/wg+/vlRSUUvX8AEfA
Fadd9IX45au8yWRo4lPKofHa9hq3SMVyUvT9GY2Qi2H5An8Ovolr4LyRZsAkeYxV
rl3JMC9Mk1chMs1A20lQdsOLY5zVE9LqQhc1TIHzVN0Y9CAPNqTIBI679vHhURTG
3dPwkWsSkNNY/SUnD1o8kuNqxar1su3iRvSa5vbckEZI8cAAlWbMOv9emOC+cyca
OAyD6H9/TUCzLdJrkEeN/26XArihjhuuCmeXgCYdIuQ0FAMZN9A8qMi/ylkolBjE
HMbHUExuMN2g5UFT9NRmyQ8/ez9XqBfvKrYzvK3rFtUmF5rcX4lbkBTh9JZR6iJg
6BtGlIL+Js9XPruFWCGs1KqHv1Uo93JWpJtgWB0toZqVX4Ffbf6s6gccoH10Via1
CEmtuGIRSrdHKRAuUBy/3Z7rf96z5jMEo+ZPBLumkZ2FRb9rwPnoiA0STsDGmqve
xzp8cMVmLmmlcHzOz4XJqfzRPhoGKN0GcTJ/GAPMFx1j+54itLZo3wNNPlqFZ8ki
TFWMCaLx6t2KlD04/xtI3VAz5HIPRox4IqK9GXaQYIaZkxCllqDb13rhEZnOHQm9
xJ0iQFjv5Z+aaiWVqs9hRzy+zM74wAyuaYVGfmP+W8RSe53SyL8dy097FmNFjDND
7b7rEHBm135fUEr6KyoTmLjBKiCXX1NK1pZaUvcvoi1Lwy2gN+BbuPaF0B2XFV5G
rvDfCVXiFuYPubm760s2gg98iW0pgYKhRhsxIhz4+J/L+taXp6j8qLos2R3z/nFo
BNFe3begbz9gcPXf4LIGx8h//bZFzEL3kCfY6U4aHxGYDOdoqirsun9gTnrlpYnA
1lCfmClCilEAT2zKSFAt4EBhgrMjviel9GviUXOCgJnAY0GVRFAwFCgyK5+HkasU
KiR/YFz/EIj1LZc8Tt+PiCY9VXU7lHeLxc3drHug8rH+D4kKJSWLF4o6UXEsQqLC
6+TfU7TNCjqXkb7CmrrJWBGe7/I+6S9Pbs+figOW2shHEmjV+wekhXVKbeL2gCr6
jk79z/wXt2aaMEL0A+Vh77yrWSWSk03GtRzGCK25wDajQnTI3hOTd5/JKZNnGzeG
Ju04JXX58kb7w68wJhdueaiNxMvdt/jzda9hcpJenCdpNpYvcc9UUuMClXYwRtsS
a2sqRHiUb1vMDOChbd7xn6x0Ys21SMIWmvUOme9EmWoQ8KC6JsCRyyV+fdojkBwt
deh23qKjvECJIlk8OByNYEgx5fB6BCXUKTGF6EERUsP05zJKMc+eFOrNKVpMl/Hb
X9cIrCm8moVlw9MjfAHaLyukhJf/2hsxduDM7jxQI79xaaS2DKH93Qjvx6FDseV/
C72sxIPKrcioS3cHxYczfid1ST9GxB/O5UBS15QttELH59+bSckHHzn2As3SKy+B
aaoepyWzqTGC4M6pk/gcYsA78YOgTu53HenJZAj7NH1iDZqF0MgkyChPXi6vVzyL
+8seZ3vQh+ldvRwQz3pjiWbUvUgcft4Xx1WXd10nHYsKzkYhmdJtkux7eGiEI4VQ
wwjNtQA6lt3+BcnqVSk7VvxcQYzTbYRrBA2JcnDcj3EbkOnqAduyWoaX5XDcfmVh
5ZZc+32LjPsrfo+YOKtdaWCE0NwWPv0/JTzhvuQpYMuZeCoNSFx9dknHn/eA8ux+
KqdXEESV12/jwLvVuVBESIhKDWKcSlg+ziqwd8W/sNCeJFt2XDRP56djP6b6tzaM
ESIjSzbpZPNRZNPzUd7XhCpulONoBepyWYgDT0trUQUNyZxXIPWuC3HSXy1ewymQ
B/7KyOBcKuXaDMZ7ccbuqdAdpFxud+1I7G9KohsXIWKJLXg/RpNHGVHUQj8luKlQ
WQYPxCzzLjyBJoy/NrpfUPpdqQwYLXzKzg8UGx4ZvJOJ/ixtShkFGOj+ig2BX36E
qnhVI8l7Q435rrd01qbVcCYHrKZtXhn42HBfziGxHyP94Xb/4w3C7yiALSJvo/1W
YWXqeS1kosVFW3VRg4VmaJjOZJ4ocFZgLzFlnUrfSXqvhKKWT0nmZWR3h8AoLBcg
9i9Cm1ElxOikqxOhGfSCggcgKjC9QWIB+x9KJj6rw9eIgY9SVTOeG/mZb8rDrg9C
c6ORbGBuKvtCBxaIADgr9RsCWC9FquEJJ0HGHLpjoXoFh7tkfkYQBPt4wYD1N7+V
159xphQq9k4/V4FgZrgZVzzrXu7uDLiktURT6ZQF8QYUx8c/HgX6AfQ4UmcWluvi
pxNEPIPp0bSIUh5lvf/vS0h/uR1bln1QsTrJPX355e3G0h4UlFE/C7cnYjZiQaZc
fcor2cKs1uKKX3b7tZFrofHWW6h/fGJitgTe9/N2TDo/xjHRf+d5TiXF2nQLiRVM
yUfZeTZZbdE5F84p8ZAiPqjutraaArjmdQ/CO8Qoo+4fORrS7zlSC9ffDfCObWbz
TJVSywBi+qtKfkP6h9kBZH0Ip50nLE6DQnxNgBZjGiGqvUJbtN9iH91rKt/OX49B
9Drass/FuMcm7DJ60WztPBreofqUyJjTLcv3RI3NSbpPIJOlzIvkp97PdMdRfBSU
Ds0yFYVze7LcOA4zKPJFQD/c0rA9rMZ6XeQbldXs1BxIDUHdhKeimbIYJv/NSPhO
FleX8rlsofX4gCQEZDQxt++JI09c10pFU/P5eFekRyr+44oQo4oeadODmD62+HHI
ZNPXv6nHNH42GA7JFEHwgrx1HVASoOLPPmNy24RoF5Vy4BCOKEHwvCqzYFlni2fr
rB4ftQ3KzpBO72bEm3QhX/AQUcfQ1oSxM1dY9s8V+/1TZRBo7iw5lpIORFJm6rA1
WHx+fjdZdGtN2kKgKseIDRodioaagh0/nq24XHTy6V3is4Nucn+pjDldXOzMtWaI
6sybhblFdfRwRZ7OIma1QHwY1lZJmJEOxtkGQB88/3/BpTJmOZ8uOhMLW69d4Oys
5wWWocMFtdV8xLgoGQmBDpuNXpKlRfn+WdfMQWLzBODPqXe76xDiPwpk3iwZ99bL
WvTmSFYiqqjXzefpxNwgwM4c5Vm1yofdGA5sUQo7OpvVJxdKjxb3NRX7QLA6W8yk
UNwtv4h3XP3zB/ElFKHicl145b4uWmuHAuiyQsL5V9mrMIYs7m9cbw8UIRbOnt0F
6QebShhwhQQr21Vx+zEU5G3Z8QlVKieU9znxSMf7GMPvpazWCZj5gQ5jL5BLE63g
FK4jqil3a+tiJZpH7rKNwZR9BZeKNGGOLqvMtMlpFqFkznRMIy+fnKGRHZzMIhAy
0tpokwpdsyKKkchSjiq+yioeHI95pp2teb47z1NhNZ+J9ck9bk/KOo/oMrnQvuiN
rJdUGl91U5idkAtylF091XNguQPqCnuaKz87+oEG32NLz4xxVpauzv5eAd5pdiV8
omrVS12ZfzA31fVjWTdI/OYJnTqSfMASCAx6/8aOR26rkMnLSrFYKU3da/JdRMOm
SENNWzCzqYOU/SifnrWerhsBF/lCEX+cvUjhQcqPaRnCA7YY4ynXEp0KtMrNKlbd
t/ioPotp0GOToDwoOCCIMxejCDodSbBTFTF2hCovrTPocbdvTj5Ty1BW9BB7EsIM
uFgzxQttjrTsQGOd5PDO44DGJ8wU3xndJEH27us1VB9YJphunfLDjS8nPiJbtQ7Y
MbG9DvrJ76SFmBz9VYVGIEYB7H32hLVfKX/lPfcBEpmfmPixD6izAsNY61cXD38Q
oYEr59mDBQ61xQGfistwMpG7/AfhpP+ZQjhd0hkLP9P64imdovU7brHqRuYJmS6B
opiA63khlG/KdJCVM1jOSgXymaAiyqn52+kEIC8Nm+IATRD6YyPI/aoCDxFEF4QW
vRm7OY5KWnsNQlKOK95BoCZoWDfrLnTdiznMeFC6XXSjOI7K95jfFNqIf0z7qvC4
RkEIOV1gbY2BiKoSqlq8mFQJJsyQoSYXkvyo2cpk8OQPIUe3c9aIs8bpOqQ7xgBo
U7xjyDPz1OGOGJ1xH0JNEFPPgVxNnaNynEr78Ba4dn8I1WIgG1IQCYj4MWdsxP2a
0OdhL6nxe0oWgR8/HUSjWS/Jo86BC8DpQtA/tLvvfiUG4x6XzjctuCew/8/QTwlQ
yF28IAHitaYF1V6I8moRyLmkKHovZ/2O6EzWF4MgksQiDfU5NMPyLDGhZXJqH0Qp
eK9q+ngNE6uhvh3Xkea2pZf8AlwaZtO1CZhuOKcSXfkrgCM+gwANfES6bXpyg7BM
RnzqR3iCczAOEdcCuFvJPde8wreBVWtPJiOj2N8wLm45ZcLGyn5ZRXmMgd8L0UTp
Se+IY7NrkFrId0QSGLUFmXm95cAJnc1EXAU618n7gcPzOiIzaTKK7FnB1rtBg5cQ
qYhWobaL2xfJ65xZ4tnlXEwTTtZtjGbIJTiQ8e7NGZTDq+LtphBAPfkymEcA+/id
xVF+hcHnnKbLi089+MpC6xBd5cwzbo3nNKj7eBRnjyYLv5YxEKD6i6WxoMPjK9aV
dUeTZI4LL9unDaT9W9JMmWpoxDrdO9YszkX1aN1rZ9Uge+czD4rJ7F3euLKNjfYi
BiRhU9XA7iJPw8BLsYXAvO7FMZQvBeIONNdVsmqU3nxqvOmjhsRgKmUCeWg5DARV
+0EZD5RjBTpqN2pmJKxuHqYf3wxJuAKKLvu3os07QMtnU3gz7Tu+Id6gfwPWOe61
zhVRDENuZT2pUelKyqADPfkATYDSD5cSdIVLMGGa0RouKCfjetu5AwpjdO7p6Z6e
FpRJjzt7fseCCToMX3uKBJHcfTA4e2xgg7Is6C/Stb4pcc4dpJL6oTPBnvKLfn0/
78/KGtAR1uxNQD3wFP3qupAG6WaxdlUMZJJmbu7kRoX+dUvMhVNa4q6biKUGTt09
eL8q05MmkC4RCOTQTG/B6Im2Fm2/U6Y2phvMUDQ9RRihvDRFZv5iIsEBFp4QGBry
wIj1WjOovPllp7TEXvgsKhLhr6SiuHF+ckmHxOf7RG4kWUY+Zjuu07FVxIDIgfkv
oyj4ovLTvMpi0G/iRz57+jqcC0nAkOSg3Nge/nvLeRWt3jO4dskefwo7Rl42mGTI
v1NwfyxllQ0c9be7OnkYgW21deyWbj9zfo8FQZXULQM3AyVJgN27a448FXRxQ2I+
QK7ImsALuDdC3R78EkDoOtS+mtQXVt9kG9GRE/S6ZK1H/rw8hBru/UHN/80MnaC2
tD5coRGZ49Q4FBkjYR1GQxDSUT9gbU2cG3DM7MWUDt3WLyWMIMrginAGWf2fPm5J
PM31lCg5VvCLu4ybcZxB12XrqD5XNil1eFogL1b3YdoCawRI0IhjMfbbEi5rfB9F
81GdewrvZUA5dfPg+9CAGbQzjbg/ZbGrtiezqKuF1GCl+uy0eYT137M5AumdMcfp
/r/BbNQ3zkGWu/Msl+R04qdI6IDszvY11/+bzLowc0lB3GUrNwIgoaGI5AmrsZ+0
NbjUd3oadNuYsoTQ2zUIxgGOcgZHXkgO73RYqYg4OL9FgbZMuqvI5gLTc4fdQnV9
yC2UxlhGiAz/5arP2+VpT087P7cTvSIdJSgEeX+68Kbw7z9S0ED2//8z8sYAKzIa
vvLf1uxgnJUHE0eaxx04/+g9Jf6roy9143zWCMVRv5NyWARhHAWJ6IkYMQfDswuy
TW74irgIEw7lDc46CBoq+R5zYcjJl2RwjBX4R49JnIHQvBMA6yuzwtIpYfH0uafh
JF+YOy79rKr5gCeIMkssj12XofCLZiaRYYdnLPr2p7bt472LUzYpd3XT9yl8Nbmq
iKGNE50qF0kV+6nRc4Loo0utO6P/cjh1jG/VYqi0IaxbIUN0XeNNYraXIYOEo1wA
W0nvy9fTeMnfgAITsGk2sHdJsoiAmqlU1K3dd92u60mgjzK9Q7bMGV2+fmerR0DZ
IC3Fcmz4M/Y8Ac2ESYutS5x3yMTGdxoTdIjHFozC6uakPTSxcOE86sK1IVhDoOaS
LNdHgKI72uEpfcW8HFlwL2lo9qFe7e3rJmEIaTm9M8gPf4mJhqVY4rWV8Rr2TJqd
C6WLx9KRd9q4+H0GP5j3vzpr3+IMKSgHv17C5UIihwiqKoxqB4uPIBPc1sfrAl4/
KkkTW+lErqrXIwAQz8ZnUGlEw/kJQryXwkYVqnQAzQp8IYsqwU+YUKCts/pw4JeR
ac1F77/dDXuZesZEcM5GYSul5vhwkvF2qXImUAEUVHjp7rX+0DArsxQAvetBugtK
SitQXqOS/4XaMvYlk3RaTNybhKvs2kcmrU7s3Dfkhxng3kBqtHAyOl7yEVZXTcZ1
2eTJHeGIcvyhs875AurRhS0wAoXBAufSvwKzgLYKJH0ONLEv5qrg7wJgoKbW0UZ4
X89kLM2teMPpt7G6mzno0XtpvRIWqti5cHqdt3cDz6+20aK5BuRdOyN6O2rG0kdN
bUhfiDwMRzn2qRxZ7ZR3aYTrIZeYxvIp13BL+4EBBlkNeg22aRRIwFVCRpkmqjRO
cVbkJCLOHIclFzIWJtLV7dPn5WHbHPsuV+qiIBDOEo1AeEnK+bZL5Dn4P514FrSU
ZY35zlj/kj7hp8KPwmtHvBfxOZSoOOfsdvyV5zXyPK7zgSLxztF2sArw7aOgMNjj
R/1stOHBmxpGIXlWM7KOD7V5tuY7UlLhKre4kPP3SkWWzQoxunYBCmtE13uhMKYk
WeZHlcY4jg9HfBDqvgx61uJqnbsFf5k6o+uSoyEfVT6MsD3jBJUbnIlGHxMU/583
a4pHymastPX/rr/PcsDyzT9L3vykHdYiZg25iDdELGW1AHNnSN3gcLrIJYj8VkPB
xBecNyoAOq0Xzds3qyZQlUwgqQCLtkkIP8f1BShs6pK8XW9MH8raiq9tQtt+p3Uk
ITwJQuPFdopuFg4IU65Ae59uEJsUQ52YQc8YcigLg5sHveYD4ac1TVxGLJ8nyxlR
wAlCj9ulJYE835qSsXsOa8MzldVBgXteFqPiCsIk1gz/T8UWMMZWm0aVdeFOIyl7
PYFSOVtqEVEuSigH23qvmbZftIRZeMnNRUHciTd+aofWUw7z+p4NzLmFJxeSjLm6
zSiQtMeTdgF4P8LXk2lQfU3yw6T4lmqoPLxY4d0kscIehP6PZLA+pR7KQqufA9yh
7VWRRWoIVw+ZMKusnP01eL34VLQCKl79Bn8KHV0RFij7Uq00nehzTgdlJumW7M1V
vkdy0PAzXZrC1RbTiWHh9bn8KTRu0UBJgIJJywOk6dSphzyLTGFr7u34WOlkXSrX
f4xwHYykHO9WrDzefxEs7FWxazyJ0Co8Uld+Q6/M9yUANOhupxMYoIsWzHyyTXol
p/338DkYO36I1Gthuqz37oKnYaQZkzRO766nWgJn9wI0C7fXkxl3ZHmni41Bt1Au
e/00YI4hMQ6f8UD1gad+rn6oaFt6V2yAwiXy78kWwRxp6Qqfc86Lp05bbOfKqaRc
nKHW/JwzkaIoR3iQB802Zgdb8YIWWKCHIryy+INKE9Kxke+w69TO8gkVqzKxRYC3
50xGTKn1/olNOBN5PwVA8URkhEQj6EbxbKMn0SNqe9dFrrB5cTI288aLfNF8gs2d
XkeodF0ZIsOqc+sRhBfITP9ZE+gkBv7248v58M9zAaP67zH93cAfVDJfLwKR+qOf
LF6TkGRmPWbM55u2Z3LQZUz6TjlgwCg6b5GFRLoNw2USgo+La+ogcFawNTLMbwQP
dMA+e5raWspUBAEK+71z4tK8K1pxdxKwbO5Eix1WSY8cC74hhMnFoX2mFnZEkOIG
hHyZskeetmmnH0gqdHJffhYN4z9xkCSjkiNqKLkMjFJNhy3csHixrg9lPzBSEwDA
PsdCSaUve0QyCI0lLKxPR4BsjVPEsdSkMHiclaoZAX+J3z0uxb+b/0JmL+88MPQT
/I+bDRIcb9jyCihRXdqxK2Cb78/ZeFmxvSTGbtNlZrD7AQg3K8RFSz6LPo49IpLb
P4hfWrD9KhsDRM+CGj/3ZkvpovuY0QGbeHydmoOEb5rznaeYWfOlZ4IeWnQNu/U6
MUqJgjx5ifB0VbI+g7qdwHuyOESefsE/RpwVHGyJQgBr+/ISO+5t2f3XC90Zj0+6
v8tqtnE+Nvg0RD5NKR2q+0i0cKXeuR5ElJeQk0VLAZKkfCQqEwKxFKgMkBxsj3Al
gBUX1eOlKocov8FdTsWEsUGIwSvFYSkJdq2zZN4yxc2lKoSPtGwnA+OOiepD98iJ
lnj0PwiWGR+Q/2+0o7dhX8akT+s1/beO9yafTxqnWxfABFejGJG9tYGpqsrOqU11
wdomYsxdw6JxWkPFFjxfgNB7dryc79WoAfxNHeju6N8WISpCI08+fDHsNgUOKG42
FqwsA0rJQmgmgiHozBORyij+s6wV1iMsytWY3kYjDZIFGF6C0AqC8kCLwtmyGVoc
J/HnghHXCbJgjClxYZm9FLMPkurSN+9IRX3x7OWvIAetHcUovjtETtOL0kgGuRNO
6GBMMdqog9TtcyWPd7sDLmfKhYFT7mqxyc9w+dxS2o+t4Cxti4zHc5U0NY6d5bJ/
UmP4sstIYn8nX+R3Yp3BdfBMODzBgQ0Qls2oxqHWewRT79whaG+iE3f+mM4XorTd
0Dy6xJ3nvGFb2zt8fGj5Gfg71AEAPaG8hZ8f4slmQSMU+qKNiR7EqsiAKYQ2aaj4
CBm0XWLOCAP/0O+eY5yqviWRMvyIFGTmc4bEyNoW+69PVAG2c2KVNuQwtTioPwuA
yc6Ic3BmPUtuKXglBQo147O0HxLwm4IlkPv5s8g8hi3tIx37cwdpsV4eGBaSPzrk
6BathUBm5EYozeR2SilXY0K8APMED0H8BTGvAsaHEpk5vb9Sv/JpABwR/846YSOz
y2IOwEBufnwRWwPsntiKWWNZsm3EzmuLOvyzk8xCD5uAHX+4MrvIwPd5AsUCxS2i
MGfmoZQLoPXEIfH0uesi2p/xg5TuhKMl9n509CK19mVcxO0HL5o4dCqSlIVp87jL
f6Ug3qAXtToJwdy5gfthkwK5+j+UXbf0MOLe1V0RHBOjOf+sxrS8lxlM98XIUcfB
isccgqfpcZ3z2HMiZkaCSionWS17/iXanY73K9ggVgLnMLtAn4s3yiLu9CNh5Jwz
oWCMkiAJO5Y3nnvF/TWJD/jPoNWRb4OWID7+m6f/r2KnyD41p9tSbHNszn7x6PfW
xhJAixG2boQXzAVxjCUb8hEsYZD8CA6UhbLcwm+7dMEVyyRm7CQpgyPcv709me8z
cU5FWy47pBr8zyDC1oBnzJkwRH5uWtnIK8RRtwFV7fXg1bhsOzr7IknJPv9tNxGm
0dwcZ/9k/E0dWAcXjyAzXftaAW3Ns4YLrhlBqm8coDVnj5FOg9p4Ntfj3+2CWRBg
vDojduNbyG5eW47R8cl1WS7qutbwWuSG3K3Bbtd6uizIxZOo2DZffFKFfIc2kWPU
boBAvJCYdyt1PkMuc6gG09lM+1cgUdB0ZOoyKQSV6/oKOkEB3NX7stA8vQgsJ5m7
4g5fEYTsUYr3aOfvnCn3vZiRVjBvyOjWlmjreHpYlFf3EXY0K8Hz6pLd5Q5OHT//
aW54mm2WSyVdAcNG6keXwxVFsY+XDkVgR8Daxy4/ERFDR5hD9PVHLcODMkgDrmgC
pcomzAFgbGeGRYM7jHyOzTqmUspXE3w6sCeOIVmb2nVTxbTiw9dMny/3XayQalWO
efB1Ow6OCnLP9I703IXkgpWxL4cmM2oelcUZV8/yroMwXNbJG2AqdBrZUjZXR4CK
5Q+327Kn2vcx9kiGon8E5t+/zCCQCbRTEHeqqr4BPIqTn/hsRfvkly0QTmGtL9dP
38/A83nBMql9A93zzxfsbbPCQxvKMnxK2JT/mDcyrvUnkxUNj0USAZ0MtG310Jqa
wjCCCg8tmNjbPzu8Zvkbc9IfCxmRpcj8Est15FJzZay4RNcXBDessHIqaybmMvSK
VXLJ3F4D0i9+dwtEq066YixCowEGYQI4ZN+PZTg6VvIbg0wg/+mlskCY4vNUl99X
QpFHZGkGFOhzVKykKfwX+Cb0cbV9AVgJN0PBouzf78bjl1/xedsSGrziXTK36hb1
Ol5QRnCfCp5bdlMy4B6yCkFKzboGu/59PfXmg72TKgehB/cY05lSk25JO2jPRXQQ
m60DjozsHbXVRCvswxZAtp0FEY83t4F7a3Hx+kC8yb/91bCRgATuSua+Y7e1Anl4
NXe8bhGAK/MjH8V5EEBQpuSCBalDMMgx+5ooOX49nPxRlHMr0Y9bFxiTV6ytGhoD
Sj5RUXzQEYmsLAU6wcKzVA5Qw5ZKa8lwKHO9aQuaBdEKUB5yp9E4xe5cpzj8hzKY
sZIwQomX4PqRYhK9o/rd92yRAZCUxrt9eo0LhpZs/b/tkvI3zVJW1bGKoDFbke6W
XXeZs2bpc64f4REl5CDIgoZ71PXF1QcPaREkfIcvYd657eimj6vikHP7216d99H9
j/pbzR3KcM8Vi6NqX0LqlZamQky7/uX3Pj2UYHZJULMGBKQot1rFG65fh4dEKzSE
dorgQeaFpUzno8lNl9wYFHRQ0229XRfEWRi3eY72f9MTajbzNgFCcXtngY2h3k3/
Fnbwe0ZnWiIQDY8x5TKnPO9KZvaL32N3v/u8cyTjx/BuxCGGgrSh+8JQ7WzKeIW4
cyjxqszFAHbZ7L2r0MdX6SKL3ZrNKzYqYv4vjG7erZp4f7fJnQ906fWHhYHD0mwW
IB5t5xv8tV9kszHckiqZYvhy1nuwyXtVcLAnvV8bA4+lMsOPL+rcSUkgunlDaYYg
rMSHIR+XX3I9WtFfw+NhiQFn03enH/Y+YPNbhvJuZoCmBCC4bFnmbtJ+iBLGcBSe
02e2CzaWi3jSoAhmQGwNOi1uVL/ryMqVHkISHusXKhrH1ibflUjWo6x+R+pjpONp
7Qa46KyRjgOV2/jNyYxnjDd3GhmVY+pbBnXq5Kp7bFZVCaVqz2Vcke2Ps5Z4sC8Q
+sPqbgpzU2AkRsO22R1WrJmecFaA1AxXjLi28va73vk9J+r4MCjAsViOBpuJr1Uj
T9k2JGtcPViTBlVcbn1D/OzL6TMlsemHdQnv6SPdy+Qrqey6D76hsySTdX0TR94r
cm6SQhA0sOPwXh3PDKmairAYoly1pl9NyX+JCwp8ceNISIEh2Rtd/jbXlKxrZBT0
ez3+2paDSGZiATXgIE7KeOYVcQG4Xo593KgA9T6lTxBcV5hoEahB/oeHNwk5qK35
fDOKa+PgC3XIagpWQl5sqsrSNF/dbE6dEF9iqUmExlHCnv2N5pg8LaMGIPuTJn90
gN8g4ViwS/GjiN7leWDPbyiCxtG2TjBQ7v0CXjpT/Y8k/YiWjAG+E/Y9Qi8KTHiw
Ql643BcE5mNwTL8aosZL4zYRBUHXVlUt4WRi6cE6wjTmpxsimd2xzAf1yONa+0rE
Zc2X4ehDK+yYIQyfKkkPlC8nVuAdYdA1O1iri7gjcaETliH1vmSSSFtoGJiHl1WM
G05JrOBSpx5qjCkzrFuAR9ibdJBOC9p4pVpEGBT80uAfrXOlyj4gd5+5jPIu96P5
7NnxXAXpgqc1sbAThRM4VQuYTQj/nV1Nd6stglhU68nQ3bHlJgsUhhegbWW04hNq
3RGKC8HzMTPxGR6Y7jNLKxMaAhWbeQU32XrF+280A0IprSqf5+DTySaZdk6cmrg/
xuXMh+OHr5cQOq7Vh1zL6JG/rj4Ix4FZexKcewz+P0QgH0OeLCINYsgA2XGYQ2wo
mwEBf2vK56dE7EwJX/3aBhQo7/9WGPsRNPAvPKYeXgy6E2RFZef868eu0TpEPm1Q
Sg/n8TYrKzYiPplm10eysFuY1nVDDkxXFTYRl1DfWVFFV7qBjuSHhqDvKzzQ1MTz
UmO7zA/2RogfjYW3PevWmuhPxa0Qj97sFI3I9FA6VdIKrOmLc8zE7kQV0puTaBds
bpD5D7M5ZFT91JxrbmzA4YU5y/mu2VaCkKEnepAlBmgPkc37G2m40AxcI/8LLFLC
YWxMHCTA+aj3odiQ01A+PiJjrMeEWgUjF0D7HmGRjb1F1DjugysOmSp031lSkAR3
mTv82x9akXmR/aTturN0dFcLQzRtQL4tPezf6yay30NIgHDuEY9HSM8ho40I7RGs
oszLi1YxilUAkahmgXIwSBSyxS/Rxd4qUFZBRE53Qdf4rMl9wg3aZ0lGwSpMM+Ch
XJU7Fmu29neyrwgTw1h2u/Ru6jWb/Tv7na3GcIKXyjnu+HbDXr2BCXU7piniip8C
mnBRfu3L4EUUD08KBeUIm0QA5AvjaRVWQTA6rnXpmwxOJZ/1whq6LI+NRv6ceh1N
xZjJVo9HdKBkg+nqhrs0I+dx4ByTTzCBs/27xsRRkcxwnoNmz/Eoo9RbIzCAxMbU
uPiSZJz46/Q/n1blmKi3C1RvUYIk4UzBZFQ/Bw9KEd7YjaODTuL8FehxQGyvm/O2
M8jYTeoVf6fUvej9aTLhn5ztjEqqPPVP9AGKKGZO7NuyZctRB/e7V8Yc8HGze9aE
z9IhOV8rV73CFS5TD7ufuXdPrwyjgOfqLzOjmCfQXHeeZd5ytIJE1JriEkuGZYvu
T/srhRsPHcIjAidILe762MtI7dMq2DnpBT6px2uy+vwoiGgvZixDk4wxTfzDRb3G
GQgIlr9Icoi3OMli/IgfpW73hfqBOIOyGTXc4guLlsRQSr4DyefVwItvx7OM1Yaz
vPQq/+dezgwrp7aPE/hS9aZC5FyyI+x2tnRLLn/J5DV51+vxo5bGzVRJG87a9T0a
dAZ3dctlKVCIyNdUcckxfFMx8A4pK+YchWQq4/SHh3Wz/3GEOviW0v38+26PgrJg
CFdao6Il07rOZHYb9GEntMw+x0duI+SAI2zDmBJJjknLky319mVe1EN1xdN4dvcp
W8ZgaP9AIAHrRaNqJR46CL+obRGr6dJKBchY+U7kPm/p1FynAycP7+JktivIsyt7
lIgNsxrTXyOVSISEhcseY3XPKcDsPCw1OfmOnOjMlaJD165v9by8IALkbeiNBZLr
4LONikRdGGBp39XtzbQinQ+NQAZl4OEtKY7hGYQPbfVkVJwbh4i9ZVqyyh1Bdahb
O72Td0fcutQ5xnQR6h1UmcavHzh/NCAn3CDlx5Rfhv+m4VwLktXNqp3qZ+T3iMKN
a+iOqtx3+1ZnXZsD4IobFXgYezDIigM7tSLkExLuJrRAIX9dyJhb8W/WJVb70wgd
puPwAOHOxT57xCkYdM+g3+CdSP/CyKKlFcLsTBVC9v26a9/F5U2VbnCQ8DpiFhud
XMtZsx8GoGKqb3wY/lqDwkrgDZDsyWZGWLFnMtBaOTCq8uCbV4MugLiOmNfCE/tI
LdhiFeRiXMXKJnvRSSrwn2qakowASEVjGVTFtsXp8UsiUB5k0i5wwB8cR8feBa3P
UBz0HRjlmuGByonNA1nHBTbLnaCWTVc5/RnWbwn/zrvDClFvFplwOnfzwcAreL0n
BokL4sQouUBp8UUBFLtfx5g4n0ERvxpqVfkchiOehnKIoJIPgo96eLjanReAvjCL
lixLcHgZNCENagKfOwqMEU8Sc6j/ATWulJspiG60Uqfmcq6Fhl8FFIu9oAmNAFN/
j0H4VXfOEJtN5jUXGaf7gAqJEun+DYgMdH5qDIR7lhOTkn+4KL2uU/Rx/ZB484zQ
KEzUCdfcqtUYI7jy4rtXgP1YInKV/EBuHyQailnlhajy+88RnQIxc54deaDv0CSM
A+ChIicnnKz4txsNRzLm+WCohTAUXEsaRe7838qD1zPZxk08RZ/36AVT2sLLhfnF
ZN4ZszoelC/zWGTy0v5WNiO0lAVAnoVLGMg6UxqAa5jvEIBCiU+GZayhUGKKxZih
s8DyKXmQlq3ZAYuaPOArBKscy18F35k6iVedfAwcaxbZr5sAM6hxAylMSmGlOss7
SqJ1rngj3EYKnUYJZk5Pj1RB+XFRQTUar88PzwSJkfGSkVhdrsq2J5cz0/NmI+lc
R+ig4Lklk3nt5j9n+jGJyUVqHVu9MuAHCnZVyJUs8Qthly+/qaSqtUS3SFT8GW0c
BBnWghruQZvjYV1G0wQ5WnqD1VyR5HxHQfERn6T+9+JUpW3L6frn83q8phY5L+A0
hDsgfjopBelJt+p0KkZG37LrhPe4gsanTBE4ESUTryJ6Jp+tZlddAqs/2lpSCCEN
uvHVaSKFRXP5objtUsq4bNuaLp4MZUqVl0/5U/LriWyot+9HlVol6G/6/Zc5+Bap
fx7pmYd4dnslLRFsb80mhtrukv/ow73ct2JS6dm3AFoMAQxrJ3iKOvjF8w3ptvKm
Zvq7Fy7eUPItEOB8YRgyA5mqW9X6pWBaTC9WkqROTytXunFO4WgHXajIpt+THQ/Q
sjHyG7KYwjPbWhuuHWnlK2loSXra5JTOeFBjza4qaAKifn7BfoFIHqUMJ73VeQ6H
iYmXCJtVoW/RxelZL3DwGSCwMRhZyHu7RE9gDKgR2zEZ+lVMeFTuDAHKjNaI/8yI
LCcKwnbwuYiv9RVxkdRTfciCh9oS4l3gPO7UIt/AdSqi2EYvxQFJukGFBeHMd+ru
e3Q75SiEThnL0FEZEESjFwBOwuFN7yJx8MUX6grmXCdODy7oMgDJapfBKODAfqv9
9pb5+1tDDSwEXRCKBWxD6FCDpcZpFBMed5LMO6IZZKEUzcWmKuAnKlqtIidb4XGo
yVOvIUhJjAWZukN7JUolRy3JCKyZiQdJrdZrTnjziSHfa/MCWSK0r+yTxvr+Fw+T
SR76mLoipcWrpni2QDYBeznH8soyD3/J29vdlZc2HvwlLQCcM2dNVWt4b+Yc8awu
wXQfZAb6Xx7hSaqPrsAog7TADdODRiqcfkBCFFfU1NXDrwd+UW9mhHFZF+Nt0ztI
cNYVgTsRgDWDKkEIc5+88QOunfkKbKWq6wJ20ThPPlpacC8RHx0SpUZt2fpZRevt
RLvxGukVlmkz9cBIbK18+Q7jOK6//dmGX0kKCBeXm7omBMzKzgxl0YwLFgR9Hh6X
u4Rj6xwaVzG4ef9oiEMTDetcYTBoDILebC6YFswIHkpmgmc1C1Tk6BdJxLu0Oiia
3CDugQiYx1p9fLEKzrSTHiU03YuQWupm1P7fAgU942YfrqLaZ7HHkWaeB7aHa/o/
yD/yJRv6Z+h+4Qqx48gyW50YAz0+Q9waCK06pq+HnmymMDZIMUeYkOZ3ZhPZhZBv
Y3N49I5O/CCqjjiPOeDegR/QMHZ1JFx3JPVD9NziXGmoLo27XBK77ym6oBnV/A+S
D0V3oOgpfgvpo/nzIqH4k4RypOE7KFRwf6IrHAnz2ZEm25YundmpFktidNS8ZhPh
Pt3tgBGghCyVrEhm7Ju/H63Uo6k0WshRVWaSmw1hvtb6oMrsYP0Kmx8j51+ksoaU
9UE2H2mYe/RHzBH8dQIlOv5fs424XgVVT9U6uz3cfY9kik3hBqoV+efvb4b0glXT
Yiaqu6TFN0lJPW4TGZ8Y3r5MuPHR6JCuK0p+bBNm2sqVmIG6rFMDpscDlM5Xm4vH
KiU0WMl0ixCL5o3Ett8XV7w9O5DwzN9UiGbQDX52uavAezlnebjjqp78bhyPKgU3
Z/rrrs2AgDMGULztVD/JAQCoNV8IQVmLH2kSSllZO4TyhwfiCLOklqj/Kz8Wpuvj
kCHTACOC23h0T7LGt46PyQJmnBNE0tV9s9Ugig1eH+rG2KdTJ3OSBWg/ZbKn8K8j
MHjNV3NLj8bmnPB4wJXb6vmLtLLPmNzV93VRfikB3ZFWCMkLZ+mn/B1fm1n4xbhQ
KDeWI61RuL8iHEAhftDPXF2mfgDUdUraFk/XT8Y+CQ+/jQfbc/bfB7w+12tHUTQT
EH5QYrLam47X1ezN4xEbljp/TV5OE65FWeKxYQzbuFm8aDTEXG6Qoqsucu0hL/KS
doHbyCcOMcztsa2XaGZZj0kZLV4tJgxfQc8T3MEk5Qr5PEP9qMETVVwKiOg2/+ab
tpe5SQSA5Nncn/Zh/ZKkMM/Gje8GaSqOnjMn/vJqUvd5RNQ9DKmkfjBUSWG7zhHV
K/bu4Ys6Pwktu85rZqvNQgNd5RN8MyEdW6a0OEe2c0GYHRHIOvb23jn8Fzq8er/3
DGAFfTmaZPOsckGDMAIBirjZ5oVIi73YUNtQJT8u2pggoXiX7VgjraGSQtPkqCJ4
wh2r5bP3I5So9yGYd+y0nm60cCLTWDHxJW8MXA8NbgivXVUxPNtrjt34GlpO5t+R
3W2B0t8gXK+RWbhSJl4O7gN9D1+iofRtXFDKOujoEnnIBgVOj+JR69/ceDS1oZ5A
hf3skyDVlagYRJ+R1t9RWQNMnOcYpEfqgzNIIj/oh6wu6D9NYzSlbHD9nD/JmWtY
N2s3n6GOXPp5/CcU5uYuIdMGgDSilYlvHyhBtONvoN+VE4o24aMr2KUygS2Isdx6
sOtuIF/fMUPFqIBxntU0IFpoj6/KZZH8jJ1w7uPUtI11eVkkvbRfn4B+uBkPEJvb
rkECvTusFLmSYvZ2xe/RmXb/LVlYyvoLRMAT5JZP+gjXD0Spxnwbutpeh9cK3orj
t0Ijayz7Gy8eU1Wdg650mUYf5kAeTNioOec9wqQLpVtRFLuR2LFuk1jQcUCYMNZV
pd1HUvF93TLw7E2Xi9k6G6L/A6gCQ2Mn3XrpuZFLCpO+fvG2ByNO9p8hrs8eJbcb
slWaDFw5gfqM8hF8K/kOHBv5nk5jvGpWPcCnjDR7/+v9lpDjCzU1ixp2ExZdSD8e
vJzhNsfwCSAlDvUf5tXp6rNBoDioEVUtH4zzNtTE7SQlJdtRTtnnxjau+OhV1ypf
jLPgVIaeVO6FcP68azgUQL2+nZV48SSmH7ffK2sR/Un/Fy468hiMAM21bPz8eOx2
zJ1gzVRzMLTAZ2xVE6XZK12aNxxsCblgLu6NfHj+nkAPmYqSsZDq+eQkI47J9hZT
HAH/k2SU7WEuhjRW9D/2JR0V7YM1hbRQ4csS0rHcOaN2YeAC46E4KRF8HJRzF4Sm
HB0ReLW6VJUhUB6oZUxjBchWaHUGF8IesGKWntlKhIsck4Wl6uZURdOdxfaZqrc/
1WF3HIgPpW9FZ7V41UblbG7APewXrN9Tu6ION3VRjwTm/Y1SK4fXm0e9uJwZy28D
mf4M9BMTMhtoRjoq0A7H2KvOo/MsFFDUSKCZ9SK27YoXQRzvpMo2ht1glkE3/lfW
TURG76jjcGEL1lvDSvKkiHjsNdcunE9F1t1oNR5QRaL0SvJFnYluiV3kiS5PvlhE
/BvULzNYBst25731xNiaBDMiMe/vxY+zwclgoJ1OmO5cPeyEmKIEVnvpiyYHizzf
Qc/b5pc+GQs7LhW8WQ9U+rYl+fVRpWWR18IbsIkbOo2s/t7s/EIlynnDyjPIBRuE
41+CF/H4NtV3u75IMyYIZNIYK7nReaYTznUeYwOnh/gYOrwAyT9pvlo8zl7m9ATJ
xKVUkXEqfc82/kNEUNC0kBpkWUuIlPxsGXKgYQqt3P4ryLcQsCmiE+nSef1/orDP
BDxoIdKiwXAqzuooVZpEDKGwli1vxJIjqsJX2iyP+ZUhnGl+WscpWXP2MhwR6ktL
DOcNA3wsZq6js80ligTIvTHIF0UMf6gq6SXlWue9w1nSCvypQgm926r3Rw8O6rU8
cSodQaV41yY9788AxzHP9AJ+WH+yLUSwpBdwWfCUj9u3f/0SwSjVU4aov7v0+SDb
Hcbk/BnJG6KAjYdcscDyNeFGPEMyTube0dB00cgKc9bDnl1+Odawztr3c2jvtgYM
4Abcqbsob1GyP/63bHp1jjAVamietGESMBhLnwZssjmsAYJUsQV/QPMbvzOxZrN7
RIsiXTRbtPPwRrGwodnCWrRPpTJJs/k9YYB/NUskqu7YbsXzEMbzY763J89cgGvG
qC0TgE/WjQ+Ti5mJGk5TMQDvZW2DwM6QaMJHv9dwJc5IR6oNn1OvsJZvG5k2K22B
MAsuTXrHcPTR/3z1EfDjYS/v2SwRjDVdE/mHpcbe56T4U/7AGr05D02YO0t/Bpjc
u7bfISZyvhmg1g4leSEmwTeIQgZ7ekow+0PpgYMIRjUjFy4qOYzHxSCRQqLzaiaU
IyM0WxfcqrEHqp8GPGE6nn/fLKHgkeTHHSdxFM/VTHw4HPZTi4vyg2XjZnQDjb0S
Ut15ncqBpjCho1A1muVIEkwfdZku7B4piVoetgCn+wTeRbZi9Py3yOTSEqfvZoUg
pb93xEeqlNVUU/+bVVUgq2O6niH0lN/jjGiX0KQ76qLenCb5HQ0zE9t4BsAOgzja
m72cWe3OefF9KqNZyNk/Ls9LPHR2ZPwqlzST96RIzrehgv0373sji/y0UgOqxmRV
HS4pxMjMHTe5IKkPr/pZ3QU1ZKIndZEHZcF/b7nAKiqvTWrZQeOgZKFsKh0YNOYI
hzGMizDy0KlzOOfSTWNZ1IAWld04iGJtz01h3yjtvf+flnj+0oig8DeC5QwN8r84
+tFJ25XMxcEZF03qVEOi961DVJh1BLqBCN58ptVqNcAhuZuikjFTgbljJ6Bvk1fG
TzQGrI8JNiepUTKwLneD7D/U1UBbmm7DBXx0oc/Mr+6/3pBwSK90gpzrdEWKfFPc
KD1T86rwRhAMcoRLnTYijzUEHqEMn1SbwOlJkBr6mKZC+UuvOWU42M9v0O93U7Ue
uRm5gwDv8mtih5Zb9k5HIyaFYx9auREPpQjX22RkcDBe2jNa0a8rbgaTT4UUkh+T
OnVCjcUj2wM5NE7tiGatncpOPDG4xeIC3TRoG7qQKiXFDRG4bbQA7tX4w9tOqMIM
uVKhbwNQNtLw7jTVq85qcVqZKNQVHDQMCrgNq1s8I9FxWSa6+fmbRK4WSmIGmwdu
t6V6Z0iFcq6t3KPViNrCXmLTwaIzmenQbMwDzKrdkRxRMUY+wc+AiTqEEEShotx6
jVrzY6wigWwrj5+giaVbfeWvEW4N9549/JREbBJfWMKBP5TEvZ/4mcQySSLA0fj/
hequvH56upU6LFjWDc5ljkDEDTl6JX6pC93jGl35i9XvjuuHaqTo69PmmBlHHfYY
MwZJ5HYRsHFbF6uy6nCgKs8x75nb4S6Qditzy9TUijIILl/z4qN41aGUwRaiFO58
viWfFxFnSHawkR2RMp18CGDa1cN9K9GSxvL7qXhvfOt2rhJe0cgy+gHSjjQ1OjDi
X1sAcju5wDJ6EHPZYOUZZRC/8bq3KcOsplhejLVyeH8vhW0FDpU+kid6FJa2OcQB
jULPQtD9VyMm4wiT5/V9bpuU59oP9MqNAR8ay5KSPtQAoK7TypElUdHPCZLHVXR8
wXpwnIgT/DL4e1WWJzRsWH0iRun3N2NQ1TyFHUlNhofRzb5n1NF7XPTzN3ha6Z3E
kkudtCZvufUaJUIkdNN7OvzAmLbMaJ4b0HNMl7I/VvgZM7Mp0nbm3EivfQr3epxk
0IQQH205pSoCgJvLjhtdIc1tgqm3WsPPRHnnm0/VMB00LONPbRRFfgPZJQzUIsF7
kSahQttXEM7foMizodAQr9MpzJiPrXTdJPJjxKTPaV6ng2Fs+luAIlJ/pOiXtkl2
neheoQaY4mRuv6OCI1gzf9u7aAGisKvAgxmMfamPOvRDnOn1wUs2Q5q0KDczrLl8
gm6deAYkLlJq0714vJah3jcl7XZDX/myM7/9OzowFN/wJXM5dzm3BeI7SdDnFKXW
RJ7VIL9tKFpdiEDPhhKwo7XtJg84nmHxfpyOcPiT1NuQKQ52CejEdhhesrwgYWIy
HeYD0RaKJb6s05bJBdRd0owiVQOaXd/fUtaTtM3Ebk7d6FdWjgEWtMCSf+Lnm/zX
ymbX267haW/Mvf394MLf/LWC5zSxqIxsB3Isz5VtW/AgtjXXFleWffWi4/sRoopE
txO0+OtV44pFtvpOE4V4BoCKWjAeMmVk7GQVHNqSEVx8rXgrAPRa0D1TJUSGMF2M
fpYrLYcsZ1ztFr4WBJ0tz3SaTsAZfZ2b3ncw94vxEcAjAzHLjtR61DlUAFFipznT
rMqyB+oJ7UWy3xEG0bgjvBv7aIvm65Vfeflgi7bP28UGNrquFgniXDTEJakIHivs
BDj3cHLz8J2GoCJQt5KK6ny7iPl17A3tTxAVSl6qlMIsgXtiuRuwSJAPfN8FB1ey
k7elAfndq3mKqtlkve+fpTiGbC8WmtlgwIZHJyR5tEckz03WCLeB5pe7a9aCvEpY
Ka9WAZ2mJKljxfWajwiqqXWrjrj7DCRN647RwkOEW4MGL74iwaZtpp5pV+4Tikt/
BZliB3RzCIeTMwx4lze+gCJEESI1EkIU24hqC/JS8OPJGSNuqImVODZQniOW/kmh
lQbs+o76l4/pk3/Io1sNeENickxgqMPKpz0b9ouvSV3ALQQ+Xs9GwoEFRopFcLHq
lkiKw7aKGIfFplVFsopuKz0XecvJJbw0qqlfL86XWz9t2N7bHaw/OeQIkIRlFdXP
ICNH/eI3Lz8EzUPTDV0+C3YqtlJqF/XJ8Br+uRsnONfZLqB0ujIaaE4Gu0mfEMD9
H2+g8Dc2rI96/o+qqbxPyXjyjVIiJ/QUuZvvLNg69Y2fcpTKog5gmJNKe8Dk7dTW
4Xxo4foM4tTQavQLSgi/Hf7wH2zzl7ChIfpfPBRdDKth37zjEi0Inm3KvxxnZr3C
C7uHUzd7zfH11BLdhDt2fDoU0roUglTHSI7ULtQPPchrbUe6c0HC75ITo9r2/ecI
Z3velA1x5nwx31o3sNjl/3llquO4s3NOjGHt2zT9UWO1sNx+PzM1NMJyeehI3ssv
giBwa6qeMTyp/GD23A9eQVPYrGdl2wSVkaprgt9yS324hI9/cIt/Onwe69FNfL9G
oyh4OLXJ8C7FV0rTysJC2kAqqHDWeiZC1kAhpxTfnw0tK6Gac0dbbe+nFGtfkxpt
/as/5RpSOOFUNA9WLkamiJXjNdaF31J5qR7jp/JJ3UGBmwMfBeI2qtIZNaCcz84L
MA0JymMtj/gQwYM4+mlGaUxGnP8tAT7qxxYefp7dljqfVFos6yyep48fMNDWi0VV
gRQjUZXa3z5euCIb/BFP8zUlH7qgk0W4XRKEFvF3LfQ7tKXwQELitnw5oiPxaDIZ
O8OoI9OV9poWEG95QRh94HdHJeNMmu2ra/0tZdj0fLDfqdesDU12Y4PrVr61ytl0
bki22fYYYAe8q7Rc2OHCweNyL87WzeUevpxvbzQeBZpclnUntcbmCHz0vv3nyCAK
AGuo3tXl7aAyQjoc6ERvPgWRmyfs+Vhd9pCeQpQhWx6ZeMf/bCL379m31+hIXePw
VGLCRLGL8eTuIF1ZuTQKpp2Q86ROBD2JrnMwXmh3hTcr+uxFD7JXAupLiD/oNKqI
NblPk/x/uIvkELhdkmM5Vc4Bebs5oeIxaWMetHD9FEguJSQHFj1v93hBRbb43G8n
GyZ4/lgTB0K+WxZM0ctm22SMKqhCRcdl3BL88KQPVbISGiEVsFtXyLPu2jEq/rvT
cwLPF5j6BaCP2ClrRt1EeLb4TpkO0WXqWdvTmRuWU5xIEdxcSUD4SHiSY8I0/xEJ
roAEAAhsLCigUH/loYhpezKvQz+0GCmYo8FaUqXF//XfMLYyusT7oMfBeBmLqPYV
b217i0TSwImmXv5D8XB+50ilXV9aLPAROaCGe5pncsKIUnnqDB+7SJGe8GcNWbqS
ZV08LCKe1GFTRLi688jNPWAXpxNBnhakfGDVZoQZwHJgU31KeSss7WktOQRAJXfQ
pYNtVyKWZfrLmw98j8Iyi3gYadBsl8EaWQOqTQ8vsKirfnbL7VPrUs7t29+0XhsD
x7othYJPQmWdQDQgqqt2E0cZqZajB8rHFWxqri28WsBydLwiGxTBIT8ls5x8NRud
j3zCfnwsPoz/jYYSgwLd/1fG4BzHKU53MPeufQf2qoqx+LkdEwPU0ZJdAFTuWuS5
QpCClnkVTxwMzeYjwrfYW/VAJqF3Vj2F3I83nuXX3YtlLngEL4mHlRsaxXwm+OPC
YEFAJVY3lA/5kla9b4DB0NgSGzIfEBrpWwP7phzBFPzilU4+uvWiSPVF90bCPskj
M4AWk4VqsX4ePbYmEyWCWmz1geh0sAPjue12/pfoebw0o3fEyMiMdUcArygMmkpB
l6OXejv98iTiJw0o4Vhqa8GN3xSGCY3UM0FvpZKZFzXhKtO6fqzdxbVamkwR+b9m
pE4e+cqyTOV0EbRgKICw1DzyzkkhJDGB4yw7AI5V6p/w2EepAbZFfCUP+xDVrxu0
RJ0KO4i/XiE2Iki+KAhLghNLiZIrOF0N0ZlY5hpJKqBBI+F+By78tUdf875/TAUp
f+Gpu1izFIuugMCC1IftXB+ZQLXbqpZ65aiN4adzvs9B/0UUhRvP/Y8KPrGqsjN7
RRfRSwrMptN2RrULjmGaFp+kXQTzr6DcdBHtqCgyBNP+ie+0sy9ybk0vQlyAf+zQ
9fPZjM2i2WHGEYHtmREZVyN7qH+j04FAUVYPX2EPYAvioTJYqFBdq0p89gCr6o5r
BoC/vCvF0G32p88XrP48BRBwqMUJmKX3arYzLBMcvf2BqiytNX3E6UUexBdUgKVK
LjMi8bIgPwTdj+kCiRPA5E+WrmGbMn+FgusHqlgkCSeWNH3gn1k4H+N8TkKI0WPn
Oe0dTx2433iHg5ZctzsflTKx1HnbRaV5IzPh1sxYYyX2mMPyhtQ1bQF6YZeTWQkY
dgka41Ao3L2ftZr3lcQ2MxZjiGazpaCXKfqLD2JXMaP6YLu5eGxYMd7yb820QnnQ
92xH28Jy+SShLUs7mqSDyLwAskcNb01m4Cu7AObw0Gg033HeKPumsMuUvvQETBBS
EJLTSeB85pdpqWq7ZQ/9hyIbPzc0OwL2zu+oJ4Thw8pP1cfdhBpmPvIN8KRPk/9y
AI4JrAZ6KCD3SPsQsxbLkD8TT/SYdsocncL6L55AT54lzlQyc7Z+i8RZUMbajFYF
JsH+OZVzRblYxRhgmRwaLMNkIP2525WHUB7ceGIK1mEX9ED9KlEWSaG4crsAe5f8
nVqHhJLUmWaBeKVTCVomIsCvc/jjqf1z22pohDqDGC1jBaY9SuO8NHEjlwLhmkdZ
mWIn7PMVEqKR0wRFLXGJoF4fdFFbND9TI7xt2Jq2Dcpzj4i2mNA63Iu1egWH8Ska
vrQ+IXtAy/onsUwEg+N+OZjLJiAmDqFyQdpqoZSjrlYuqmECmfsegERJlOj8j+ID
oPGKqsVfmCLaoWoj6pAokE7+bzuINWvKT27l+8iITFGJHUsP5dJjWlZeu/yX8wC3
77kE9bEKwQ3Up/v8b/ida5c0VeZlR0E6THRLafmcfsb6gqHetmvYqz5ezWzP7Gsd
6AG48YsPi+pfYLVBXM7jASGXVgYzheRebd5J6pfr+mxM/TfH+z+detAlDWr1PVWU
XMx/LZKoL3AiLzdyUNJWsw+ZOWszuN1D1VNemwFWRzA1Awz5jh/PmPBuKRJNg+2c
TBd+qmVUow1BURG99eJn+Lr3mQFI511gNJr15HUpTq0fkjdPiTwDjrfnd+AChhVm
dfLBLL1oIKOKMODM1W+ufuHSXSsmq2Xa95D/dRR56RpCq2Mr658JfT8g3ZSWtBGb
xSQPP0qbX1nZhg15zSeRswrW5yYmhP54qXRgyN9uylBBPx34X5p/2A+uOaSbiSot
aluERSXmWVULur37XBZUZO9MmJlhQ1FWdGHQbY0hJJ3bXG3botMB3eYmIsLKpKcJ
mQ3JoSl59c1jkycogBhKWbGUs7tCmBIZDi3loJ2oNMaEnsxkXhYfukEhjUSQGOFo
RoCvaWyP0UZmsHTr8if/gv1DqZUKNXdOfRZ1vue6xesIAIlxBjbn77KyF2r3moFy
rmsuhw2Bc67RpqrBMGRWhXhLJKKEz66ZVIIBX1qfo6o19IO1Qx6jMzeXgFULup9m
8aVFJ8NUPJ1vZr6FD//rSQjHHGTbVtYz0N3W5jmPCw3PpEWB/CYWN7YJj+iw9tsF
793ThAtLNbvrul/ivC/JhBjUWP03UQa5IB+zivRAtmGLwxKyDBFpoh9zJWb5bb5R
r1fBCmTXO8fvsPSo6AvfLdSFl9tOYIoIwp0VMo8Nfb/8+ZFzRLzwGxGq2/wBqkoC
+Fq/i7T7BeU+K6wxtT6Bw/N4tBcLmyP2XALbYNH7ZKrXaWqaPBO3eE49kSMuDzHd
AUvuuxzgsVRZF3mJ+gjTJ+A8cqkv8LLv5FyIqVTRIsmNc65c4kTqezyoNnBSl4Wx
g3sdiyZrDQowQIuBdmdEbeR/nvkLThLFKmwWqGHRzFGGN8rlc9T2zG+PMgAiqrJg
xyNMIpBmMe6sigofYp0KWKH8XGAZwFLutiaRszqB33rbWw30ymD5gBsT4dFKnWGG
W1xujD7X3cNfrMaa3JP4efj/19S+Qmmq961M56lQIDuwZL9f8u5XxH7umaIJec8Q
NBDrkDdE1RyunVL+700rOG+oCGjLMQA1QBgzBshLZIMxAHS4ha+yvGgC4mYGmQTs
RJeaP5hT4hJjG/TXpwjSOTN+DLLkbmcJaRPkCnjS8EvGy+U7I8toPSf+iwZwTwdS
pJNydk+OzTD51adO2TdwtZpSh6PcnEGVpYsrVzAaMw8mFeKLKD4Iuqx5QUWr4lgf
KzdVtyfpadriWDWgg1mnETon4/osMPDMwg7FRTGNcRKkS+yrEHDUabYLg1eOolgZ
ZPSBLd7SJltkJh5TSe6VUfl47HciI+FGJuOyXA6udNuCc3TOCAVpzyZWZ0/v2fFb
/v/8MDurwL1ZAY6wTo7JOpxVJ9aOHKTmbgrGwQm1oTkekf/4Le6Q2MCP491qm3DB
MVbJ53Nr/97dZdo0XqeiGBbfbZeTSlScq2fVQkSO84myh5zP60mTWJTLXThFjJ+c
Yhy6K97h3f8wBRGaGqWvcrRUsaufe6i+Z3ctqsO0GrlTHB8LY92B/112lInqwckT
Bz/hqP5KQQb70Vuol1woTVhEDJXmH2s7wIHnRbSvCrQgrnGewfVI95uJoVSlJwPP
FaxTcpAM+kL6t5a97uWwKxncfS2W6TVzhNv5sSLH2nTrGOl1agb21NDbZhRT/oQm
6IK3StnVAo+btHog5wL2NKQ9GGCWrdn55tud88k5/XOMbk1eizblW/LruxzO++vE
46Ztnfc5DkVTUVrgYrHhP55Kj2HPr4EaHTX/C6pOuW3FS6JKGb/nMEcmIgsTS2vl
X0Hpx24KvasejGHhdMnM1UztEx7C5+6mH9U10GZRS6TVHQtfWhrex5EE6ZCxtBij
xS8tw5buGhs1vTIMFRYEMu/0XT7oInWhVVFVl8bOOpeiCJ+V3Be9Pu3kbSRZuNWy
rcrcPicHhs1zSe962s42qwtke1G86CTlXlonqueebyeSSMaG5UywviMX1rcyL0Fs
18jZVlzKIaCTO9gpKWwGAvJk9j010dGjbLBHJEzj7SrS9PTdePNERhelHzoqPQgY
bjaEVIt3OEdPP5mPSgahkqWAf+R/ccf//PnbXaYANAgnRk5AcYYAmr1df86sJiY7
MRQtA0vennhkwS1oCnOo8iEl1I0Cq2hg9u2AffOFuMj2ENzBip5wrksnPxuMZbEn
5N4doB2nVaXkJJzFaJ+IJreQ3L4OIEZmcQ69F0Su5+QDQZOvJK1ESeyRSefAerHh
Dq0Mne+rrFf7kkfnCOG7SwTq4bcCmOI1iWzXZ7sYK9WOtFhSgxlqw9inygkvYudX
yMfGAZQ0YH/gSvifMPKjL5yq07hJOSK82IOqmiLOs5jqpK5qi4aL07sR4S9o7oNd
v3u5GMr4yZBqyUoJRcIprWiLkQtlMJ884cHQZDFOPgwOF/kQaZNiJezUvkc2pbra
MenkxDtxgjzsQK2t3pB6r+y/ch9LwMrbIkYEjiKHuXjSzcORPCHjQ1aJbk0HcRkq
56He1Xc3TEG7WLiEVTQ8LqO1VmIGdOufZ9B6mrGumuGUphtMXhvhMF6bTX+Vo5n0
3ruC9A7wCooj5BMSHh0SogPHc/sGwKGiNHTTWwfA6h4NAvjndvMMk3Ch9XVK+ARa
MDAGdmL7kGk4URl1450rh3cYkyRdbs51PfRWT2fr/NozCfFIY010R+gOJhNDFyZe
gmaetLALqgQaocpZ/l5KX0dAvzcrcATY3nh2g3BfINrSVWk0Vivo064LvISrJ8si
WNbJQbJ4BmLH3vzM9K0UFCBYCufKv1uLZoUaPAJV1kXroDfnW74PiM16sSps63xe
fv8jZMhw/WB0PoRjivdit5aNJS+Ef/Zlz6CUKl/0aULrtP1t87m/uMBerhjR0z50
TtYxRrTQIu+7JRVFwn3ue8TfbIL3iky5AP46cdVVQeaQkddSK7aEoLcD7OAAsMUs
PPs99+7Lv4nRER0ZcXylmdU/o78xXq9g4LxQkjPMfpAdJ/k2g6vF4MvXNvjbwzou
2DYzWwTRctqk5fbtaqN77eIvOYL/ImfPjDA1qvRHaB6EbpSNvztphybHXUlM5V8G
6DHIYVH67Hjdn5f7PH8wxJ+WNOuLEzQKaMSiT6mVi4CccIg8DPG+6B7MdACDrXUn
5LXw2yfQNGWtZ02y4I4ZT0yNDlzFMsth37XLCl+nwerAB0JvAwa+Iir49P6Fh1wf
/XCcUGTt2Kxo82FMuBGs4jVDU4JS0P/mSz0j7o29XDnoTC85yf99IjGDXdcpT8Ro
6FSDCTQ4zbZDlDPSi9W/ajDYmRRinOOLdKe8jh47600AKE2f8z5xIG/egaicY56t
qYsRmJlguc0jY2sPv2dEdGnPfQeIyzed8WF3X3Rs4+9Nx/h7PLJoVnG585p1btME
gLs4oUry/ZULaRx9AJtLnHdpFJsGjzA7+7qdvjkFlmKf7FGKUJKkJ1FVXc2Yr40u
NcPEISSvItcc35Mv6hl03jp6OziHOI2fVN2luWsbh9Xz7jWB0ITFXSiZTINJC7dZ
me6YMA65+dkOa/vFsFEtfI2uROs8b/c3BZ2A3FXyeCAfoN3IDiVHyYYYeY2nhw5y
oLTfrKWBaiPN/2K2VWg3tTv3b71v2xp3MgnRGtvfxZnlbZCBCyR1dwiYQ5wb7Lxn
fmWD4HVhiDVYUT/M2h7ioxIYszBgGIXDm6nlN5rvZGdqQN0w3mu+nRtvWJeLMlUk
hRcZIGXr3toDGoOLZ4ZDUDPDW55hfssgbBMZcHLPWW7sSd9aaYmLB1bGC+fZHD+5
74Y4/DWKj25htBStmcYn28s64PP5sG/GPBIVsJbH2a7mHBfogm6ImhhC3W4tN8pp
RbUOSR1aY4xknUpDKH2cOGvYITxJPHiEGneJbpgV+gGgbIynIYJiE7bdh1sHEW97
56JUzACIUyz5Mbz8cIChw2aUc0bWX4dd6RKgpvPVmhCGGnsKPa4Pg+ZBSs407YzW
ryQz1G+ILkmGppNRhntrHYkq/3RSzk2WsN7VeBbqo5KdTGGGl1aL5FRQr1JMuza9
WytOuy4TgeF5zm4eQDTbDm9M0t80gzxWCDcNY+jvq5HWKZ/Nn4E4qVzs+0dSRm56
OwH7ySR9zpy3UvmdXoCd+4y1l+SSqty4zsd7W0BlehXmB6xSwvTQgIMdPsnmdn3Q
t/Z+iWPN/URhCmkWGMI9HGgV8mIc9nGSGufvBZ6pNUMd+5lxLC+xmilQtPyGLb+o
95nkTo+kDDIwYQFp6wrVM2o1tpYl/sbzElqN53MdI6apR6GEg4BwAkPS5v9URdMG
rGngb2VPFKQWELjmWrZvJ/VxZ6rjsCdnSEMEBaErsbYN1bxshYF/6Kr+/QaGBgcY
ujuw5RAEAtAh1FPygaaU2GDW1SHnchRkFtaviWo9MbLt1DDBJHMw9UcTXgwnHCbn
4gv+N1HGz+hXM64LC9NepUmFYo++lNsxbZUntTgN0zQogs6WlEprOnVbu6m8Q1l7
zbx7jorez5RBCseP1NVlx0/MBswpprFF2XW5PGHxT9Fhm066IkVEk3woYcg4c6U2
AFxnQuKcz+kqwIDrNh9I6HivgM7yaWYN91i4eQr5xCLMCvsFvaaCqOPohyawgeYz
DOn7UgeRnhobn1vdayF7gljjjqz9OIN9EotyYBXStPsNQXt1IzeITI0oTMglWINQ
DTCncl8REinpf/8KFl+KWx/mXO6AN6+SRzb3xhMlY3gzT3gniDLma8igVbnePF2E
Jxrsnvw1BqZ6Zz2glEZhKPsr4UtSKDQFN+GuLbtmf1bCP+Zgp4DaYmLnTboicwXZ
bCAPIn3MIV+wVRsxfm/lf2RixSvwgPKMJYmougFbK9jyOTrjgmphgOgPA3d6m6lr
ELz25NYTpiRLegrH2YMg25aUYqGG1KBgex6wAH0kV6dJTloZ//ets0MLb6afKTM6
rj4cPZm1GqSmvpqkzv6LY0s8B7hxvXpWGh6iHUk8U/bbiOC5zdmeaMoMaphHpulq
0pU4kxkmSiU1Qi+Mg3PziOvs3rz6QyD1mfcwpMR0tPF9SNJ4hIrw5RJ4jf2eVpA9
imH83O8lp06yL9q2+boX2Qwfl4wf5dtUba1gthiObPH0Z3zobUw6eKTrifv3DJqi
CCFM+hpEJi+Njz4IrkEV3I2FAgeyp7MW4lru2xrgRqEoB1Pkj9u/aHo8hq3LlsbQ
3wHrejtwD+SRylI5cZI9HcLmfpFkm8vbdN05xmi3ytdOcAvR+KKZ1l+n9aL4SAn3
pUsLZhRRB4j5GMGFGKFbgJRlfrwm8N3T0bKGto2q1D6HH0nXHRd4UQsF2VQFm0d8
1X4PSCK47R0fQePrE02tuuRx6pQK6vRhKRNxPn5Vl15Hyc37eWLz1vlk5TG1Usrd
mWV29OGdevoIte5eNnPkWfHOseucTaGmSXBjMNESsr59508DuYZGYA52SgBxZa0L
OVsBVoXciR9TqPtj24+lxYATJ/CfHT1h4+dmDq0fZ2PFKXoikMfe6iLJpf9TVhXP
zgraIxhyvhGbdOubXQhbjiW8nhXyFRjA6Z9ZaJitbYEB0B5DJKssr0cyUpyox1q6
Jq0wpCWu1nLHxuI6nfHzS+wMOFpVPkjVRG9H6civkJYxcT5/nAc4RNj2CuHwKKXe
M/nm1FwM/IhSyZgFTHsWIGg+MONDsKddAs71Q2XoOBXSAVx6IBhZf/qWViUltm9U
wNYSI4Yc8/BUVIZLUMMpoNx7oOG1/z0+7wAuCDj40RSJwCN64X43idn0btVyUUor
HR5HoBuKGPZFtoRkggOwCNiSElGbJtPvUDt3eUi5X1Ec7tsi90ToSRk21ELyxym3
K6UkRnbPf/W+mfKiQWg261w5cMMIkC7J8gpJu2X4ho0J/M8zXO+WBP+3JdM7xa8/
S2eotx+/Xth803/tbZqHsLE88OSZ2Ci9pggGZb1f5xyjv15HXZLRnBRjU36rlM+5
PFmQA3bTtcSkHhkp0mc2/IgbL8GMVfaNqjof1YSNtfBBnmES8Ah7ABmWv6V1JOXg
fxK9NjpccTaRdkEj58ayjazCot8ixGG10Xriek6eEj5GBz91VH4w6/DvfYBwbKqU
ZHUOwHe8f8/P+++gHGG+YZVO6JTpyoRL9LLEJGe9haG29V36FFmVTzciQDxEYQKw
DgP21lYwy54uToMvKWmxdcnCVVc0cNcIGiIHr8bF51U7uFTVSTR5lKR7DMmnWYp1
fAfFgBlzYjfbZCmpN8hQmAutV2eswh6EAWF+crafkey+3RenOMMFLWDx4H1llt15
x8fmCPwKfmzYF5v4Laz31d0eIYOgHH/zO1uVRCPmjf22HEKm7WVUImroW8xg/cqw
0DKmGv2WFRD7ZBeELXBsWJgz2/zShK+ymx4CA7klnBZnSxtMogaId+OnMtb1MQzy
fXaN0hPM3nV4oJrnJ8h+MD8U5+ncCwoFS4Ud9OGcFx2bUHITjDtg7pWMaHVbUXfX
oHtl60G8e5UiA58Rb7aM5NPU8SZlZ9KdtBV6TlP1Zy/oBrYp4JULp2EFjbOz82Zx
C785Ue0NtQHnTo+a36flCVtFEbX54C7oTDAODEAgngYGCslwps3TijMK/hyxcJWy
KqnbA87blJHGeEZ68L1Cr5Hk++nWBhHTg1Ufbk7+UmYNFweUjTF+BHjGntHCyVGC
e1hTnfrJ8PAWT993arMMlzuQZcxdO6I7kd/c09wPeObb/L3sK3QA3uJdStdRPyON
/QFkoDov3Tx+d5q5WpGESrtHOLeac0ShoOaCaHe+ipRoAkbnu9G66Ux+WYJVh3gM
4D5OLwnHJZbbrpZ4g1+JyViOYt7es8m9NRD88/QyCPkiTB1cl3kLSxt7Vrgesnrb
stX2eHyIBf1TLBdNq3xDbHOBCjEIu2q76TZ+IjXbbjsdnpe1a/QhV1Wh4qUAlmHr
IystWyGKfGV5bWG/z62cPjFOOmctRoqj+W8F0gG34jKsVjd8rrpVy6IA9ZQS/p4x
Pk3GGPZ/rwSStZS2vCRLqR+74Hup6dUnisqJqrtarcFTl9YCikTPFHI/1jt21z5B
nE4jqazflZVjmSj+9NbpwmffLlPCpieFl4n8D6sTElKUXaYBDrwRehYbtl5Nptrz
h7Hw7/qv2a5nbIyHJh65AKetCdtD/Ga4zlioIxGwxbmU8lQms0hexj1ugPZ8Bhdu
78gVEtnH94iB3IZSMulWIbUnGMrjbW8G9M4hr1EK+pf1YKlVho3zUOV8478yECEa
iNvqOc+t/qhWGOldmEcO53FdB8CPVGM85Y8eKX2VRckLn0nFtaG/+elPkQCs6jkk
glxr8Gw+nen0Wd/rhczGT3TlGpSw5DxDcwin5M5Qt5K/Y4BgG+duA+F5xz3GDaOT
/Ox5bxvxh2Wi5cqqzvRGBXtkKr71Usfw81vjzf91b2bTMdaMznnKV7KjdWCaxoyb
GhSLey5ftIiF1lUwhAfjfssDVNpGbHz0BawVgfN3fWn4phUrcfUJncrdwK16RN47
ss987GNCaQRwR49hA6zNOj8JPCmgwgw+wC9BkKakGgL6aXdietDzs60S/1rcmGc4
f+/FIprn4gGozwfeTY3tlWeFoSh3TO6x6iAQXLNe4CeRTcmYoOorRQhnHhEgVMdt
eLhf7GZUYWic0UutO8yea8yk17j+vLIkJtE1dRNyppm3Ns3/aJjrFVAh6cxfOvXJ
KQ/NU63rMw8y7T3ZG/NFrPsIP41ycqWct3TAnlWjWgoDFRBU+JQd5D+33Pdd6TAe
FgITQKS2G2SiFvazNxejcY2QdWCqZfCdq7IXoDiR1HwgQVLktQ9myE9jFSwmru5i
Ny4UtSLx1yLtgkswDlJwVt1+Q1arzBfVRh2U9ZQquLjsXgt5U9JPZUfu/2IsYM/w
EHqIl4G7FjMoABQ/lMUujATSOjJbJBnzPzSSUtmlvHn/CSZhsn+PIo1v3dNyNHmW
/V92J2jtR23w/Hydmdv7FVN2dsZWW9HJBJGvq4ROb6EQI7x8cpaimQeYGPNET9O8
aV9hOqBp0E+rbIr0KeLf8sdOX58sS8fqSFKpHiO1jjtQSqUq3DDCBaWFM+Q7zfwJ
xhPCZSnSNkRyIpOopOx+NFmXwrD1gWrVQU3BIZMk8LuFDgWzA9+cScKme3W3fZ2f
1ZiOohnagchNpBAaXvQTe9twv0k8doo+WpkNX3MwiZkPVM26w8eRpjmnOPseGyLC
ntsWCyTD85sfcSND/Sm+wXvxo1Lfb7P9c0+lAMK7mRmtGr2U+a/DOxirUZxIgV6S
at0VY1aaaorilVYutsBrZUsyK1AvUSEWUMkqreYW/DdbvPmz790od3+smD7nDe6E
kygVwZiJZqrGcPZWtj7v8+mCmppfHC9YWNfIjB1sWCvyaYUrb7CBN6gsRdKdAE0k
V7S2S+bZhmFdf5hm1ClS+HMEw/zsP4JkctuH9GvsJZb0I7X+T+BLIXuolRQMcdrP
LWqTsOgIwO8YWgcDo83HHe/PykHK8nMc/Cr8eCq4J3n4YT/WP3iLuTliULd+KygA
HZGPsEsFDI++fQXeMZeWQxCcux/KXC5+levQffkMfJlQSy+EP4wU2lsq/DJMUGRr
xPeyALI6CPNf3d8QdrIT/ViXukBG3qtJSdHsXiw6bxrqFJLOXKAqLYHYDxtR/aVV
v2U4ZJCn0J5nHsty7jT8X0rsx/wf10sgj/bYIopzyZuLfZW7Ev1BClNXxoMGhDMs
f/28aeehBOHnqThcE5lYGfxetiEWdxQ31TVxGDa4krb/fgPI8PhQZL8EL09hWTpA
UioUyqhjmDmuSbTVYN+VWbZa7GhhSdeivnvTA+drVRaFuG8Ks/dcT9R+wnFeikIG
Is+4RW0qPv0id3KZqKNowRdv1SiUQ3aEqOhnA4RdwV96nVULtcji/WwSijz+hhe0
99APn7VSeiAo14FW712fcr9XeNjrz9EtUNaubNeAmSH2cPuSYkIV7Gej3sIHxxkk
634XV6GTCFzuFGDARNvf+FOyTPOT3Q+Xlka/S0JnFs+Ad32Dbn7rSQFgBCoZ/GRW
L976XCPXHXcgYCGIU2lUd4o+zkJay4lwFrIL1wvKdRkjN0VHsXB4O07YGKFcppPn
7ce0UqEDUeMY9KWnKX/gM/bPWgXlUjYLxyB3g2mYkBN+ujzcWMNw1ZHeQTIqyiDn
maIcz982uQw+yS8wiBxxPNLNHIUyInkZwuBGrd2zID+c45SJsQV8HDdydJ4ysAe5
0znYCDBCR/TeN2aJXRu0/5Qci/0Et4F1k6C1j7oIcpBm9STjS+Nd7icTvV5zjsZK
zBOjgOJp40AjBxCGioBqy4+5lDnHYFMpj/eGRGD53vI1b9A0495uVhR7IJNztwzV
rAooYwkRJBiX1qpdy+mqsComysMFS9XfdZbwqyeqr//2ZAxU4eDQ+A5jF2y9dOds
pvOFgmoUnZT6OBTcGQWwPGCzssF9JlGh4PrjCrksu9Mp+XEppYIlnEcF4pnsgx2V
yLnhwKder28q+hk8zKylwJ4s/QC4W4UE4Mtzm6larFYz4qSCXruHr6Dy6qYsKtH5
t540fuOJcd8f3JKfTC0lesh+aFCzMtyrj4CVs3umCWjVn/kBhfFK4CWg4NbCAD6g
YEdoy9CrHIvJHnspw8VdFDULeLnG5v0rVf7mmSjrfCJZAowuPN80WvH8iuJ+4sWg
qO3i34MgieJN8/NWQLB7Cd1l9eo4HDlBgZNVr9LCCfJT5Tkb0U2bf8JhYKwrLt0c
BKBOcvsFlTSQSCzOw8yo5jmzribonYRILYh2HLS2pycKPZdo5njXqs8YSHrebDO/
CQDRI+mzHumVZItovFkw1sw6vmvCIJZ/RNOJMIJSBpC0QX4T5moCHTmkddkefmZx
7ZKs1NNc0DUv6gLEJBWx87+gaERx1PstxS/D/kOitrck+hgkQB5W79SzLuAueCPP
5Z/u3m0tM3h6MSel8+hIQgktbtl9w2zYYT/5YisnUJN4rDeNV3WNh2xS7LFGNR5h
IK2lDDsm+UUsCWUhd26DGLiJXUSF+Vsg0Kwzg1L3qJ09iItqg/ORmhlF+SJ8sLLa
6yi8JVG1qRZ87WPGbBaoOok3EwxwvTtX14RuOiRriKDBcvPZzXVsgRaZ1FJX38zx
T5GT9QTVcQpYexJGiSoUDXFFm7LAacTwUz+B2A8Lc3OyFIbYzQh1RHwgZCeEVgS0
+A/+nHzgsMmLiDW87UhRhwtVk4uwHZszvoAZj3rDe1fTBBh/2m7e7nG5TuDAifnm
Uw7TDc6slXtY3F6re/8PhRUDpswmQpv24wrPi8+1J9DlLzdh/OhKyvVy6boozsC/
XwUNd9y1JFfi9MAwMLpmHXvl+mpvmQmlg+42c9ORyKaxXswENgQFKr6iv9SkddyS
W+tWHauMNQcp7DI0GzFfdYkfov6RAygqX9X9+1sOid33vUvHKY7eZFmTxk7FIJ+7
9smQi03/l8wa5DRpyxuVotMcAZ0+bqQuKq7uOrgujgzAIQT0ame7pgRAKO3XRJvi
/hEgYRAetk23PxnDWS85xEChUXbhDIbQ0xhrWeGCW3EtrFuMLdV970mQwdRsL+4z
5m8yNfrmengMLVGIGrQyp0CFfxpp4AZEtXDgWlPlczvQA5oRtP5mHEE9jaKHq7Il
GFT6if2PlJ65fIsYM8JrIyMmM02QDb1FavfFBkaA+1YQBvKL09x5TxivRD6RVWfw
Uc6t1YxnvVh03r/Z+XuhL8iZ3ltFUOLp2tXXpRLH/aUAC/cJbdrfjIbH3eCf1ESV
zx6fKNLXaOcpON84YtTIlgr4K+D/q6ncok4OTsWGjzz4k7YRUwGMApphjArvIb46
Xb3iiNSkXjznrwjEVqBDJystpIFJNBvCZU1HmHm/L3MVWlCx76IeFhjOBdtdIbO8
tMCayWIpnh1rXO14R2zexx64mp/qYD5z1Pe0B3QMwP53ysBYeFQ5yeoLTq5q1m08
FnZk0WzFqvVwqrpSBU1XJQEI5sjYj8IgZlm9n1r2jYU+pP/RZWPAcLZDuc30mpY4
p5EcoVChA00wi+k0QBa3yi3yt5CEvB6+ILf0EyaLG30dQllrRPAYF2M0LV2rq8J0
aSPAWiL6e1obw+e52sU/lsjYRz/fM9YdvebJTd/wWCFJoL3FnlX/4nolhlhZ0YYK
yzC72YbLznO+MaPYhmCjtgBQp6WyLTwgnitq/ozKJnUA15WtRuOsIThah0PsdyC8
5G/ojRf/HA5+CbEWgzuGXStHlW5wKgCe20s0BJ+XiI/WsybhneqRjBcprrhP3fl0
U+/eUUis4e5RQTeSJ221KQxIQsTrS96Ls1+SWEn5jKcAgv8opw3sr0HHMUCQJp/l
cIldDRUUAY0dW4NoCIy/9mSy1Gp2Me7uBW9ARe61e2YgA9rG5y/By9AwnNqBHP9G
sjKntkzjj6HXidvWYScJjBL6DYtRC2VwPzeWp3OeZtmdt3KE1eRnTl576v0WSQkU
9BjjMoSMs3/k/bGJh6JklsTjX0ocO3hmHkqOGo0Fy1+8HblflFiPpi1WE/ltKS57
SZYgDcH9s91mBigXbzL+ATwoFgVJCm0dATtwrOqLTBU355EOXkf24zzueinJDO4d
HtJWt/xZ80AsSP3+SsH7EVb/LmVS97KwmiNHtCjO+r7VBr9MNyKYNmXw/fkRTgJn
x2blkyyVVzQGo9X/tyUxxtVq5TMm9sJLv/a7pY+z+5vQ4iiCRYqQjhWjkHMG3Is4
riNvKA71JLEZ1LdntHtmdoLGKVzMq5lfFV9XqwVidZagw0H+qmlHsSnUwK0FWj12
9dR2e72nKv6nXjA3ZpAL6v0RtyYP/r1gw/QuPDz/frcsnWvlv0SOpOeGOKFLr5KW
Szyb4RXSjQ31/XVa+1ewS5FMSVEoRqEbVnHklQJttEif0g5hulZi46C+2DKml9yy
wuaLUL5Wu4dQguuJKX32uUHADmT/lQsIymO9fo1fil7gZaz327CDGqlvOGOwty+T
eeOcYELRK4T6Y0N8y7UQaz9Wvbkzbxy0WfBq9a5fMMOhelDncZQdRc42xtVcr3D7
sCshF6pytvz6rTl8FhhbfVs80VuQPcagaM05CV5gw25tTfssUA6Qm1ZRXIUldiYO
NboFgQF4xsbhuxOTmYd2y35DEQvrbMjjK65nWTektgLhkCYwGlnhtRWaxnFAtt0C
Zt10gZf6ZD3BTogfuhuLhULO1EyQEo1i90jBEogDp8IOlsIgAnkuQkNqyPu1Esr+
+AZetTObcwGNOFOyGzufqMRE2h45mltyVc7v+R5xKFvtkA3UU0GHNGIzZPlPXu57
qGk3bUefqqprRhRzpq47z6U0ZXs1yDuWjtdx8GJnQnJUzCVs23xHfQCQh5RO6x3x
TN4+py2w+UHWk/D8FfAt3mGrCL/IF1HJDXJ7QQY8UKyY3rlCYYYnrSxHEieCDKOk
YUf2EpvyBymcj24AXuTgfbzDOnQ3lRf+wlrAouif1v/A97oUF0hwItukNun3t1ET
8yMhWecISn6i9zq+qfhzUesunrmwnD++VbMAQRATP4QR6rxhqVnIa5JbrWt/lVpl
EeS6nzJ91kD+kLLeRhizWIBtWmfSquf++bcgZwcj0TrRnTMvqFInbSMEO74QFr3O
2p5lfw39W47+odVUOcDIhFYvKGvl/EJY0ISLl6wJUTb6qWhvj+AihoCLiE4vr1Fz
8F93LXSREIMCIuCx/v+Vh1s25c7c5Ugziz3AP7yv2sCPqrNXauyeKcWsYvmxevxV
UfW64D8NMJ2LkOy1atteyreLkD5UIFtMR/48fQBL0GxuI3rHGXzGH++O6zVwuvWZ
BPBMtoYgTYYXaJFW9y764ZxaT+fSY55jAO1tKwd7EOK/uBvD/ZQrq9vXoWzg774N
Ptn9dohnXMVdDlNLNkGnQvA5xXvhTc7++VrNk+GPHYwyLx8gL7ip25+nKPIJijqX
yOw9HIsUfE7B06Pd8t+qdErkGiRRtepHHDVB/k4iP1emmZwFc8JvgTJ+GSyKETGh
W9FEaE5QdWyXNhNPC+th9Lpt21sCnack2hotsQo35lVYyfZoxPHveW8G039dM4am
IDsTw4bHx8pgTmDTebuu4FnGVU2UdBa7b7IMfhZ+QFJ4tT/iUC9hNd7zaiXjR4jt
HDTl2/UFSdimMMQmJOiUR7KFFwiQc6dCHUK04sKDR11d3wN3VBz/WoEPUl/e1XNK
vKAFX5guYMmxM88WRqtvho8+PYqnHy7Aza3sPjO3APQawRiFzecHv7bJr/cHkof3
52xocKG1rpddktKmBEqKA7joid0Nmc3urwdA2Ifg+4WJyTRuoEioqn/8p1K6JkXJ
8mVXrTrAVB0c1uJTMyzx8epNomCMMWbz7tD+AMQv5H+PTyzPB7R0IvxTCAC0XmUV
HU91KI/wVxOp/Y4r7sfJePPh9h+e0IaAvc4XRscHdt1+KFrzzN/hX12nSw+S0iU5
d3EZy1FArbXYqpaH3lNX0xp3vdhXTPQ6t7UJOpeSNbzzpVhwQEtguulSar4RfDkE
OtMO4QBgv9vm+S1kVW3d/abItgKtm9zq/gbFm/DlGZIVz7ha6YLL7OFzy950CCLH
Rjas8hzEMwTuu1hLOSHSNwAz1LT4a8654gKvry2+4ni2zntFtC5yd0RF7o3b8vuf
Z9sVk8GqRoX18u1mPutYOL5LkcTlKkPr3PuLhXY2GMYTlM3p51C5zVJnSzmhY3sn
UfJRpYtdPhri5+8PL4zbPjdD8JRPAPt2z0j1f0PsO0QoobYw0lxV8gnzfVVtn2Qt
5E4wiurEcDQNHM/40hOrBzwNbN2QyHzQiQXnxBvnrUd8WEAHknrT/+Rxmfo5yk9K
cIq3DCbU7Kk92AV10f5N11Q6ut8DAH+Ny+o+JGB+Jkj6jUKX6PiAjpAmrrE62CJJ
xb1aJyFFHI1pvNz/lTELSopoNClGBcGxLHNdXPEBEsYZPBhwQA9Y+75pdFNzn+aY
8Ib1MphFiRAOsteV6phdme+WmWOc8wv9knII9OK2tnAjivGyoxm465bAed8Fs35S
FawF5T6NSnXv/1q0+0OTIX9tJv0n8eIXgL2GEAt67eS3Dh2dGDPEnvYTvaGOmVIJ
jZqTZ6ixWti3tY2CGNjrImorm607PpLhiiS5RoFxgBnN/kG83xeuul+uDd6ED0WC
BpmahxfmcTJ7/cZvsc0EoNlp8j8F+UVlTUdqXV/AvEDlKTV/caKp4NRiQAKGRovG
jQNzzgp1lpbYPPoJU3ZCxFKxozAxUUuVggKHMcK72TUZkRe9W9g7ObsdHFwCjrl0
zN/RDYCClWJ2UfphDjm/SVx3LMcAu0gn8fENA7j0G9PKgtO98bYbM7px5LK7u3Gg
pewaqLaMm9suw2IqjeRWssmFyV5Jm0d3DH8iFwR9/KY+r+IzJfvXY2+qYqvyKSal
OjchFiAiA7FPeX5PZ466fHp0aMuZcb4t8T6ARZSxiWs4t6B7t/+hVwPmh9+ywBTv
CET2Dft6W34lduBv1bByIwgVHLzmHWHHE0pxUtlxs4nrkpjvGRHCEKd5pR+fADhD
yCp4fw9Nhvp+pVA0KPH58qpTk7Dei+hBUvrMyeVP4zxOoBcXEgObSWjCNYoAAqtG
Ykw/JbtAHL5OzmcgOMxxyrxmvz2X0V0H3Ham4kvnvMLYocjUh2F1eq2pm1ziSWG/
lHnHjFetfpfHVjF0mQptg8qllAdD99gmX9cq84fY3mcpFeEqZBmb2yCjbmTSpaJY
1wpc5bFatUqCcvwmDc5I2D9mJnsFaYAn9+msQzMGiqbk8QNZLI6Ag+BDINBDe/e8
Ir5uBy4OVi0H70/eozXgxi1sywknyTqKuBL8Xz33LH1ElctgWptaxmR7zGygkfYM
X/FmFkQU0b1VMybx7pj7HYLINT0EZ2nHIZA5x1/Xmnag9uBXdG6TMB50V4HJeNrx
XezxhDAtC5bFHfaJ9Eo5LRSevpoiY/NfQWsgkSzp/7uh+HDDO06ImffrgyINivp7
mZiH9v4pwQjsS6LNCYgqCAj8Xqjm19znvrBPEbvO90EHJ4at6uoZJ3wFA6g7DRUo
0QSr9xMmQxyNFi5tmSaWkVX2CfiUAAO/Vxq7Cxv0RQW5Dzbwsj041OD4Rn7qSMmM
eMLO+GwMsOC9PGTDPEJDmWVD9M2XiIeAQ246vp2gbA8hmCU4hepb8GZw7mU00B0h
p1inNqjQq6dKonkzV7QP5BrFTA9OsCrSFimOmU7DdlHrB/nxF90hOVZjtROrOrL4
mrBtOBt5qYtC6O0kj8eEtU9iwV3uHRdWJTQRMUnhc3t60EOqa2WULsGGrufnePm5
x1/UX+DfYfUYjq4hqPS7saIlX9HPMv87r69rUnO3379TlSEO23vSfZvj1EQlsFRk
aHqjgzruLR7CxSNbLOhiF55wGhSiBK/7utG6rlSSR2jbUkU53by5tQW0uhG53mZM
BhJC4A53/3k9L+D/joo8Wb37i3MtoQcYXrb56+sDJ2eBYi33W/bZt08D+s4XlETC
YmGo9GlcLoq/d2QUJlPkZodDWcMVOsdAJbKMv5tXbfitMqleVNtdvgTA4jjbfEcV
kUmPH+7Ihe0xxyl3+PSp8lr0wmyDcp6JP9OpfwqBUZQZVYPGVfOBlP08I1nA/2Jc
DPyT7HJ3zZ2tgvRCOisze2VoJVWanwfgCR5bkEQcKh/Dl2zazkEGYodl8UbTnQqe
HCnFZv7KRvBqkBeV7xnoe4rYtPUpqgGat3QBx1aF8+1b3uB5NhPYtpmKyJgdQEgB
MKvupafwV+7DwBzUouKtnvbJ5+8P667vv5k5sbB/OFgGmSBGdbPxCmJf8YMEi7YY
aFHQbgjsS0kjzR5OUG9EUQQIZ1DcXVIARXeFh8ymPgtq37t2Qkv4pVvGGDwCbRYQ
4R5B3aUvQxll2wbM3Xs1LnLWmNw8le2eFk1FP5EB1QBpio77YUB1qGAkcdHIgQhC
ju2fVJEE/QEd1EOmI3RExoA6G3Y7mWC/YiLovta4qKwTiIPRh22PqhhQQXgJvQ6Q
waUMgh1ppRibFeL80LPKfX8UmIBvlhHskop57MlglwgV2vakcLIcKldnYRvPgwKb
FchAWEUQAaW0a8EmPKJWsmipBKBZvEtpZ/rtHFDGXpJ1B8vy8DM9NPlbUJiGHZ06
GOrtX+x0WAnN0xTOHwWql+7rxvW6DqEmsAJbmk1t1CIpZk7IXkP7c1f9MFg6eulo
5ze1yh5uZHxK+LISLRLjJcF9jJDkOjHMiZSzBrjgyVz38rSWWen7eLPD2WZpFe3c
vuVGSFtlpTV/T75EBoCdA0g6AvIoCkKuNshp6CKjzCkAYFY2UhHN+XZNIQKXwxhs
rrILsyUgvQ42LglqDg3LK/CRjFsDTEMflpI1+vPBStU0Kg2Sn5x6eyMqsE3OXAId
oxkmCjS0heiqnfMaUByUrWCfw8TCO88uAARFXzS0wz/fGSrvd7Yv2CFsYnm4pz/q
UI3KauC+00Jv9ZbfHvCQcb4BInw7FESIFXnH+r9lOesc2GpJDdqlT5r0wO+4b7c7
x+ps5hMm+fdbVpfnFmK52pcKXDE7qDAZC448P1C1OJ2+74enkE7SYnXZh6aCdktv
j82OjBehc7lJ8so1iHot2+1LIqdVv0feoSwyczHC3S3dsdG2yaAUePDUy88YYUfG
6IpsF8iLPtP2Wf/sdTExdjk07edKZUDx2lxJGqF5slSuVGOpmNvbDzrmGsQphnZd
qj9UdOLHmUOwUg+M3Ts7geLqiVx5CeI7TzPkASoQD0v0s+XgMR57SwPP2YYAoX3y
EOmnTKvrT85Hutcn+7WyZH3GBq2Tj70sAV2hlAluVrezA0jhHEg7kxJ4m+j9IWHQ
NkLwGhKIbnw08KMzuGqSvRm/C99GfFIN4m86bk4F/A3XNl3rOAbncT1CXuT+DoAS
vEAjzaMZrSEE05PYqy9AGlsM0Nqwyj5NL7WFERESrrcGMXcDXLfUk3BK9khSzjRU
Ox6hg5glY+g3ooKK7n43Jho7oy5YCXP7/4m8Sdi9vBisPRv5Q1+cH0n9PuOSssOq
ca+VKX4g4aWaa37r0e0eNk9EuekkghRICHghZPwz5PDKk/AlXU4tmg3HWYuSniY8
lapzF27hFWXyih/4P/1zYoEWe5ZULt9+336kpk0l0pwejbIPCVrZ1dkdsrEvjbHt
hlzd6BcfPDf0q9JApQWG0+8s0+lc10rwzCvNqqqvGH2rb06Jr15pltKqwpfryAcW
gwtlqhQSKtpMXMCQAT1YEEOaYoRMImuDEwZlSsck8aKUqkBgcS57kr3GBvy+Vzjt
ZYJnYS/PGi6O2wf+r/77BATWF8hoov+imXqO0l1Ai4Xc9ojR6Z7LfvNJZZCdOUHG
Niz6O9LHMg4VwSiKbH2DQ1sd2WVSo/jnsQQltQRWmKLv9vQ9JohINcuhkOZalNrD
aAyZnDC37MUI8xZTe2R/67mfSBBzFCU6ykQFMoilxDFKCvs3AodAL5afDnMBFtTh
d4qlj532RPI2q2BSa8NZF3HAitUzOlJPdVbl1VZAqI+VmF56bJBWcpNXlEXhj/VG
h8jbHYxuUx+R/aOrp0PEHVO/lhr8m4PIXN1knW/hVZFZ1GawWD7iGKFCu/8WJq8I
m195UP7OAm7X5m7ebLmZpb6U3+qNQ6sKbwHzcYFBoy9VB2sMC9sz/qjvwzxY8yfS
yD697l9HklfyTumgUE8lGf3m0wbB6AVGfxoKt/2WrZFPigUMtLL68kYVDy6pvRAG
DhUL/SZdVeqQwiP3accvNGtqLyq9PuIOKu4C8QjgU7xf0+9jOjEfgaEMuRQagbAu
2Ez1QFGY7zBG5BHnU4i20zbUA33FGzxx6DTVbq49thXL0tzfe71lCX1gH+eGwMB6
tjhT/TlEVZC53n2asPRhBT+eKgXYEOvpIzPrbt1COzbb0n7nsNBBxSWMo0Ku1pha
5vlLk1ZD4KMs08I/c3vEuQL5zouciEgeagO1KGRQfBGKjB4djciAmpfs3LHjVMFn
c34XpAqWrXR8uuN1LXTkSyujl7HWYrqShcALNHHLVhcogcizbl1xWHQ+fjYLKI8f
zmxGm9RzGTQdE5pJta6iDPzu3ceOOxEf5mVxNke19ecSjmxtv50SobprXYrV7mMO
qktMTgsFc0jLexF1O9vpi3EuZWvYKJ8kblr4++M6RWthANL4/YDMdMGeT9Q2jJl2
c2C3BAjE7MY6SmpOpwFda2VWuR33vNuFzA35gwxzK2t78IaEr5n44BiT/QnoJWmv
haQ1fX1VodJ7J6AB3jHsyqDxopC3Inp2H/PLAxvjQURDFVGHugXveewhgZf3wsFb
iZz0pGhEtrSOlmlwpshCEi3zac0DyJRCKlLRNlNq0SU8W5kxcBSi7afEzZy+x4IL
G3or9gzx7KesGEPSMHQt1GR76xPU313KW50z+xqjvkOfDIA9uaY4/3Nr0Sob27dV
CbyBou9a9CwUC43cNzSYulIbBfaf5LPKkmi+eUOLx+F8q9cv3J3JmzrW/sUt2h5L
E+E3cZyeFmrpQB1GzDZ0o6d2XwN4mOVhhWJdnWaZKr5TKrh+3kMPMb7mGoTV/KOD
FDFIfElAxSR8EMbhHz5t8/L0yautTeNB/i7WkwD1hooesET8PKaGmdd2g8yMRS9i
iOYwnU0BloabloUf/1wGs7ZaiGkKnKIvMXFua2hLhBKn7N0/HUBW3uPboBP7zyUI
A650XbmwT7UAe9qLAE0EoWRcxtK5LXxtzcFFa6qpWOwgKaZ8JMiz3DpIdA2isVnG
+6znO9Bz/R/wQRugO8fw9ngxZYL/4nibvo7LOuypSQ0cLGZxYwcybUHRyWFxSKwK
3uhPcy0Gy/BJiE04ol4j7lEHBXqnW1a1f4CKnquQjxbA2J9mSh37toOnGGD75bxm
rBGVP/ry8MnsM9xSqVuJ7CcAWzGMLgkSW44ieKRQ3cLj08JW67gFkiBQniTvtGnH
bIWRyQukTYYDVHVrXPw324qMdmepLAWKoMBvHumj5AnAJ6WSMWCCX8sqThTVUJ8/
TBu2Rcmf3Vsm2/D4xy11fxR3S8uCoEzm7rwng+kqYxH15Gy9eSqWXdQbdhk6SfGV
doSReZlPri7SjvrodWK8bR2V6xQ9/asWoIS2l554nQL6T2N1qU4Xvf3mxV8ME+Kh
cuDvXx1Y2Ejh3gQXh+IZXEuJfwVinhm9nghYHdkvDtZanMJt3EUt7JTSZdYG08+b
dK/wefMPc79YBtnTqyHb9LAiFWKda4dOmfEDmElMSScrnNmFivehDLdiqTnhVfhV
eQCPv/UUxxWPCCfrCWYJ+2DK2LJzzxaIZhcN0dfOfxvsomsYsvoOneNnuki2lD3B
U4CiU+saPec2uJY+phveTtbvCaXIbqUTcjRJrFO6EpPSbyH57/gnq2hO6a+RlMnd
1gEQWXTEGuALQpCTjVJImK30Swfa09Fr6fUpVvzpdAqpnfMy8lxn1+5UbbBCHMlG
UTznbRnm7VDFDhc/A1rDZrMC2pyo8EbhDvIaPapfgZ2NJx99y5MLEzFtvWaZgVil
STuxRquwk33LOlfog43AfamG+UX9gUTGwCj5knuyZN7KqQua/rfcmXF0egIfwSd+
N/+N1hG7v1R9snKmIOR2ZplykquA8d/YAjwK4iXu+8cEAWU0qATR+7gEkzKke0vr
eT/EcXU+uFkAHjLc4EPfZRYtiZBA71/3GB3U665ihUJc/vyWcsubM9l00JBrzK9z
YROb4EuB7DyBGzFb54p2iNNgJws7P6uNdpuEC/VtjfN+Dgc1Wjkp6zdTz91MQGMq
v5Aktmntgs/ixmfFFKz9XfrpEm+Fc46+E07VlOjlCZAGgpOng+R9kTIFc0KguTeb
GSFQgW/QAttxV2YuT+jtWEXaq9B3bdxSPVlix6kPRCUnQflhaey5ZHlBsctWhqh+
xrg5sZrnw3D8HgRj31sKG/oY3DQdtJLWH1irQ/oK8QZY2u4gCvrm54DiMCVsjr2F
wQwf0F8tXTri3W7WmXd5lHmfVWv7LkLp5u2rHTcB7e/R5j1r7V2jXgIm08t4hFLA
6NqQ/xew/IGTiobbXDztM2h6BTE9rD07+0IyoGcGCrrFXTXr9aKre6+A5PiLV/+U
nVi3TR+kSZLoIDdWdiQpi0FalzKJHvZxkLiAucDMo7d0hugVEyLXYu4NAwkJ+WjB
Vw3oHVGSVcGTBtjrAk0mo//snVAlgXotvWblKSUjuxcO1NV79ADqZFVp9UY+LTPz
2G3Nn4fJ93kyTYn2xZMhtHxZMS5fSC98YQHlcRJpzEdEO69CQJzcZ1+bj9oTKQQI
QjYi8nX1wCPfvX4kwwoviQ9cAEkbwZ61kdO5tTvxjB2Wu1BSa1CHYzMDx+04Lywv
oyUhB6gqQGRfzAq4ypF3oekvefhzjFD9RuO5E7Arq1R4pmrE2tY6idMvonUqNrSQ
+cgTcX3jFgxiBabBIcJRETFsCv4mvgwSUaZsJdLcZXdx3bEPFqQ955lQVuNspD2a
3oIPYgppnG9QP4gq6KjhmhvhIjqKtqWJ908AI0i/+DV3wkgWl/sny93B5caz6jzh
Lk8ocjRCXvqV/oK6Isevm9+3bvUSIj1Bed+AUreUJxAaTk4K4ta98ehs+PdIllLn
Qo+ssExUZm3NPq/sJG53DMtd2LR5Bht7y/PtlZBClEe4qGTDRO0typfkNsBZ/TLu
EqI72YJPiu/QzBZu7ph+OGveNCfzzUgQbYvMPgBb98IsQMh6hMU3N9dWcuwnETZy
9eIG226OTtMOHDIipXYyV3dp9kPoolAtuNDtvH9IDqioXHDU0b1ZwLJVBcXlUUw9
89VI0O503DvsKgGVROhj3NBCbYzPqSWY1PQZbdKTu2JN+KJw8RQzGn7qYCLiLCxm
iJU/YTuMzfc6WMeKKtCsLn7rFdzFoQWQ2aYPpUwp6KeNT3llRYBXoJQbmIUQr8xc
HG4pB+KGQcFnhgRmRkQWOlAy6NsTNsDaIG0wCq1SwXYde1cfmfjyDCLCr8BHszSy
/+f5KcvBX0ZpL6QXsdzkMBx6R2+Bsbo6Xdyymrnlpl+XWIlQtSY8YbnCkRMKlVgu
i1QW37fTOoQ+/zmVhZOYE7KaeDhQv2p4zJsNx9xdbEuirp/jUHZFIaeybAzoQCU2
l4D7iP0LFglAQUI8mrj8XAmZFxLQV3ptOwQaSghkvoyqZJgbJexwKd+parSzl2JX
hX7fSRsUcv3xw8tlJGBij+/Tab3RZjt0LlkcGnzYucMQ6q/XYhLg7kdVM2lqe2w+
k+d6I7Su6J/PSAYwdlNqZczAbhEult9XfImv4QGsxkbrlJk8K7gUzvgSkiN+CtJc
QwKKS5S9cSB8rv4lIALPARDzI9twiD+a6srjPyULFKhU/FGtGzdR+ssobJdJi9Oz
9u583SdXm/qh6bCoZiJwLM3YU05lYNb1/strrNn1uTmvTx9jk385OnTUT4/CuYzH
j1DCu5X5VQQVU3/Q49I5lyva6dSgZmKSSc9kHevdyJb/4nlEn5nsd3obj3VVbuv6
89c6qGXktr+8LdcXpIQ3Oq62dzjJNPuhyeL5gCH+m5C3MLRvkeWn7o+Rm1RLYrhO
wpTXKuXHLejvsWWZDj9KIM1PGQpCE6aE+chXpPKYO1FapX3sntlMEVdt6Sdd2Rgx
l+LL+yUgdEtXnp6MaElCuV0r1/tR3wsindO7EM61Fu54Y8kFTEYOMYO9mVr09tkA
5kpIrgmGyATDE2agmd55dNzc4O66bz2dnmenPEKCUAT/8aL6Z2Sxdw1DuC+N+/uN
Zo/6ho1wxGUQ9E31mo69OnzXJITEVMPYcCxQ5y/XA3A92wi5jXC5DzkXtPl2K1w9
khhL7cdUXziIy74i1JpPBj6VwfLWHxEXNBjfXWFCZEdwxLX8bkMkJacON0NeLq6x
KnC5iH9HSq7C6bc0y6Sfg5+nWA8eY+IMb2wTMCZMnTYvupUs+YCE3EMjpl+n2s0+
fA6CAKPMKj+Uq/t3uop5C+//bsov29RgkdtyTkomD4+KGGgLWe/gwWdbtPQF59e7
MwvnMP/5Gp3mtcqDCP4jMMMLnoAbbsREio7MAHovcBZxzXEFfwYHMfnZXa7zpQII
otbcI39FRkusspB/T5JtrtU9if03VcNSlt6ehMVcY85HD5iljLF3/lYfuzE8+Jmd
62TZBkt8VpCIOeTLwqwLskmIdBzYuURyOJw6gh1wRkEvV0Pt87vWhq1o/PyOzLxL
YVpDxGidWtmr+2P3RM1IWOv4RfRNUXfon0vIXpzkJ43EEZbpT3cyyAdg4UAEUZma
lEfTn1cPSoDxyulghtqXgCYJSWwmFVoFerOZdwTxBtgn+V9ZbiFwmQhaCa3fJ7+X
G/5EHFnJG+D1ipiXW4srwGbrQ8fXhJCDc2aij4kbvgrckW4+lQT+TvtibxFLFtue
u8S4VDKWr0XB9t5g7iwxet/ZQH12ZYrpLacu9kTsCfpd+tBWdrUHecNL2WG2BisD
onfiTSgLIFSJ6ob2+3dsLVBiB68E0xuuukkgn8niuvMLFoVISBcBGCjpclvJsp9K
tWV6V51XgQujzt2coN16QnJauHGXuikE39zxVSjMGTid2EACLiDqc8aYwSGNq1ud
3RFWAg9XcrCKfi1P/6rWRvZqwfqr2v7rnSoxHV2MsgV6lFYloMvWnXbVDYrGNe0+
YVjouiXdFqxw69R0vbvYRsqj/gB7KO+3BqQf1IpyXRBJ5NlRaBPXvfUY7bL3w6V8
q7R0uJW2mCGpiqO7SXuAeoGf/hqBbmkw0p/Ophpdz3QeF/52kuoc8uo57krroKtS
C478q94tx67Gc9Ygx1D8+zzSY2HNaBLhibPXHici8qar6xuZLu63lwXaYR94P1RA
pSp0BNZldvcxYcVTrU8KRIcgBOoKn4fB2gYFlQm1MEZeZP2T/pHgrWuz30+GakcF
XlMVPrcDcG1gaYVl6gxoDXWmWVsx10SyCRtjIWp4ddbrSRKX44XTftFg4lXuur+x
aYN7GkE5r9Er/t0VfExBS50B4IXOg/1P4dEjhl7HE1yvEzBZ4K+lrr77KuoFVDtc
v0ec+GBgExf71d+2xPu0kcf/uZg7N2Ajwa4C0o0oTYZ2r7UDpoHY+EbHtJ1+1GIA
3QbUbN61A+GjTkiUKZbBC4WYw2HKLXg3bWAGiQYRNVlL2y8U6TfM4HWTli+/37Gf
s7xfYqUqju5rxbFeeRT6pEkVXadRouRoIKqF8TZEtIkehIS7qfz6d9I86xioc1fi
50MO/+JmGn/+WhLtX7YYN6kuWguaebmD+Oj7KzUTgsCzz93x+5SxraFvkCcSoW9Y
50aWkgkcw3gmLVNq0VncDq3iwQfE9l96snf9dp0nrSxMdZQyc6ZCR5Y0r4DCNhg+
rHSr88mvCeEyWjkSLm4En6XwnMf18gm6aNO9OnTA8nZ0xjLjbp/M+QQ4j40wTUo0
F8lLzgstvJFlhkmOlX0crsb4QP6mUiIsjUHIxmjeZ93OE6RVI92drs5SIEu5KAUB
Th6cd48/qbuaahMq5eHxmdSL6eA2iUb0pOTFkYX3UTLcMhUdd3fjdY5krZZxC8DF
UX/oN40TYxWKDjY+GmQ6Cn5h80WbjfGWYjWVjRzmLXT4zV8U0tS47dEmbozDla2Y
c2y8IPwIcGjcdSUUZbHUycL0aHAv41CULnTE7QLIaMxA8f6RoQYWYDI50MQjXyRY
/aFIKrx43lvUbTxMa6zTB8FOs+SIObN/xk0/vHQm/762rG+2xi1gMu0UmKunwZ4m
fYYmIveO/joElXu2+ZrkmCE+zUiNs7vC1pXG8m3GcOPRiuL6TPVfTBbltXNMwJ1r
zAM6dgX+d4M4ZAHPCPs6Jg6kz9u+314+IqF1m9syAi1aeOlmUgjLGt+T2qlPDRKc
vsuS7Y3ej6iNI6vBA2/VGTO913GUmaL43Nk+l0J/dIfJwT/ro2bViJEBprHeeG42
U/zG02hGeQGmLiKho5Nf7aQFPimdUxRx6X6phhbq8DrB3kJ3loyjcJLHRBuhi4Ed
6K8t22y162tO8mKiKrNrWtVXasxq5Tv/0tSjdJuAIn7Ar3zPBMoCDKnt7j/PlkVN
I+X86AemquB6FkuXJ2hhgnf96BnjKEN77783aT7X7XMGu+GZKOeaq5vg84jVA5e6
g3uJcNeBvKLvuo7tnohCvVqjEjSicDCiCfUijXtWnsncA5Y+iA7wZEtWo9CYH7/f
gMNTk/z1c0Zzq0LCGkowHxv5RIxvldyHJEFnJ03ESTTk7+LoNKksjRcF0/z9Grq0
X4kTDyeYh0sGYL8dI1FCFaA2lLpesnDJA/XCz9nPuz2VgfQ0c6fOVK9Z1dPLwYK0
n1etk7LVzo8aMRoJCT4UtcbW+RXx+RU9xkHOIIFV/EazBaa2QTFGDA0XpdpkFcvc
LKYx0AbRn1CerXL1qhMbtDdsEsPJTgYRthxgySZLvsdy0+DkXgGEcGUKofN2Qlbb
97QRGMVFM55emgKigrock+/ZqwVy+eAV/hXtMNUEEMc/U3JJw2bKbTu5+RyorCMZ
N7oA0NOepfsZURsaRTaZchuZMO/KZpMxd34o72jp3CiTIB3Uxhi/OR9PeSbMnmed
k4yEvaT3SckD8GN9idVvC1BP4Ef9EhMAIpQmwrRNQgiMIo2ePzuU6uDG11ApJl5z
RaNUiqVCRBIyUW3vzAVBbFVufOK4lDyDu+hg+m15VNaIpQcPYR3F/8BCa+9uNEFm
ZvxZi5TkE+zZLCSlApFAAOMcU4X7379eWjKN5SScEhaMA9Ewes661IbXRABcVsn6
1SXeg/YnPJFzvtmeSbfIO12Qs3jDa47g0ED/hKs0deiPtCVA4fJEEydEkaIiHjmF
dEALNGxvLn0f9HU/mtmH46bVZFbAgT9B0BWyk9zG7Q0orYz151aMP9wUBil6kzJr
f4VkFnpjZZ2gFEOTAmSdyExvKfyEtUeO04wVu+FfPN8l/VEVgrCYPJGRXMdHJW/1
znf3BUsm4bzCz7YFbOmloGsqzKHMYtTXQVQHDpLFx0yqmcj3UCQirdRVR8E4MZGe
epCPT4zO6A5Uec2TKIeYsaBX2pswVDa4+O86UCmZUR6eTdzb+czWr0UuhkvEDK8M
HX4v97F4B7E+I9wq2/mfXUIsBL5pA798i/Av7lD1z+CCvmXbV3CRSt+sDvE/n/dO
zSFdqJQCehcI8HJxk+hUOqrHjuJNGPkcXeTgPluR0CzU+bEtNG20Bb+2EzUmXQFb
6XDKya0k4nty0ov+J0iSzRNpnSMHk7zOBMzeEL2zqQFPA4Ta25zPWSmTZlkdQ3Lm
T0wAPoXl9IDuorXMZcoxnUc+bjbstM33qKrOYFDiIjyDqLF/VZ+KfGdHIFeSlf7J
Mv52vRK8RMEUq6oT0xfo10RtX2ixz1UoBOq6JUWUjLajW8QuibuCzoI0RIZATiN8
bsaY/q9nqY16Al+q8iClXRU4kXLlfh1AtW+GXNUN+c734jO3/FrBGqMrRcD0g7xf
4P2FWbl3uWN+40lu2gbSoySNNsradqeoHx4HteU6lXoUtoR7T5e9gEjb2voeDu4B
mAd/20Ny1WCxw3W8ZAz2kv/lR8cjVexvp7pCBX6fYSqIhBGDOy+D3OA2J9ZIWklj
GcnGhMJP+ZJRj9K5LRoej6FcwN6FGV6zxgYEjkdKm0PIeVYwIQBWnd1+wbrmBFX/
ojhn9XWhnx/HHYw+wt9klC8dk8xQjN3sUSimOwPymQ4h4IkWzyMEsB9XaS7cJmkT
Zi2HXWDYErx00wMuoSQ2RlLvmH0mOhsKj/SoiwnRzGQlTITnkFHtAeIGTKVr4N5x
FWAIhPI0ZDbgLfEH+3T5zUdexIa59J3aAunv3HjyN3jV7DmzSUG3PMKYsA6abPj7
cBHG+B5Fa076aZo8oVtt2bbNB4BU0V+FYwhuiT6GsXnunKkKtEsNLVODAm23mhvb
DD9kcM3/XecBN0BYOammhEfXQEpJpi6mNjZfNpkvwvJeKvyI+hkSmXZbAKV8Fiuc
MYFtCvqjd8rzvzkrjTQe41Xh3k/jgww/RMaK4lRO5/rK6FpPviiEXebnQ6OPNWea
TS0wf1wTQv319Ilsb6OFbu9JRlfJ0DxKIQpDilWT2Yy51R27E7UYceTuAzExhMhx
ZveQdoMhQu2N/kMdxrMdvV1Ja6rCnqFohNzmNgJoQC/atOV9mjtcaiAE80Nnb9ii
JZGXmF+jkVvn1zIrqolu0QBjKKBylTWBxzECvug8x9OjqaFR18G54wuVv2bV+BhL
RaUHUXtj0Um4Oizf+Z5YmviyoGl++Frh9HYj4U4szI6++76Pk339eh4NulGO+Pdm
J9gRQEub3ywuUseK0j1ZXe1DF+bmFpJiaBMDz+z+2m5RXClgq+ltnL6s+Bz4tKvP
W0zyU4rEcU++IclC3hYcRcQUUeaZL7F5KyKSkvycjjILVPFG1X7+R1hh+XaTXG1R
Ox5ZBr+qDfHTzPaK0zJHu+7Sb5AL+ieF9pzoFMAm059gTx80Z4H7FnrLcFFajShd
Vbu2/fnZYbJjHaQ0n8sop9SCDy8VVfobIXmnrYVFZRKKc7dNdbvbfbIUB/KKZUsx
7UbsxKSvrw4XgrAdpbGFZ/CAqIga/PTl2vTPXQaxOyI61N+ZmkooHopa9RYCpznT
sG6uTumZ5zWLEgh5uPVGg1YtKL8Gy8NXNcs1HiqpRIPGLWZXRSx9Z7GJlUKCg0At
Zh5c/FKgbgxgqvU824xZFXTFFBw8BG2csiL8EtukUYAI7ed33MS8v/NW5WzV/Tyf
HiUcUwH7kHs14V2GngLWqTc1o08twbtxzwDxx5qZ7X0OiHR8Lvx//Ho9CHs1g6gD
hwcBmsp/x/ff3d+6rsxeywcB3rZce+VbzUIAT6g2d7zQ6/i4AtQYEdaX4wNpI5Qd
vaWsb4bvoYRC4kzjLuzAdE2Xen25jRdF31L6/6zSsoTdYQ01WpWW3dZ57aLmwluz
wQ02AJd6WLbkU65DSmvPXr6U0GaUElONuNw+hySphrX8UKt1hNQgaA+ksGeP99xc
y4k0sbmy+1PlmldJtyTYMtImjxiHDJY+qXzk+5q8NsrQfgP8AdnyjKyf7Yl6tlVQ
+0tCbj7fp1K9scBznZRitxRHqxtdd1UsIbTpTDqjfSwmSkYiUjsrBEstKW7EIbAU
oehxifLXaYkvAhvxsF4YFfIOJ0HjIeI5580kRF1mWcLocEuWt+KcND2C5iLWdsP+
PzlpQdjK3tpaWoV0teCTZoReHPVP1+aiRGrN3ZfqvTZ4IVd+IEpEbwDX17POWlpD
btBij1IOzJGXni+vvcA53rV5PpcCdKIX//Mu3MMGAdWJXEcUTLqNVbzShkfsu88l
+01liBY0+bpu7WcCwaY2vKmo03OMITBTAok8x68brXRSbg869NUU6HXWnWXLLZ4u
tv7uJK6UyXdHesoHOurcU+LYMgReu3gNcxeC2+2hvdKM+v9Iov1Lo0F0OSPL4txl
J0acPbmn/JJvxepMy57w+/rI6NH40np/yK/NhE9fmU1lLmLfEgQ4LRPYS5kIREkr
qeFTmA87PSNpGEw+3k2Kk+J/ECpLec3h56P+F848/B+bkDWdQBsh184+e//IVr1T
1AhGQJmty2O0/evuB8dSIRPAhMM5UayGgI/gxRfLpHjWWk54wVAlm0pKVkuixPZJ
Pwu987i20NTPCKmzx3GmRlWSS6NPRq3prFQoEWdtizFMa+fXHxsYFZAzLmU2Uj/6
uNxq7Js+wQz2ujphxiBWaZNbNTxDNj45R3xZfS/izhuSECaTWZnHw14ghpNc3vqW
GJS8Z0QtgbchmqI6vEO8rAALJOlPHbjWLYoXFzAR+ev6iKsALo7JosfJPZKEg6TV
ZzXvRWOqUP55A9DH1Ku+7sX5bNpsq4zesOA3QfW0OM0ijxVzylVpqcrMzw6QfTh/
CLcFeTBORaOrf87ZlREqhqKWisSdKP3lPajONlPUCb3corKLOI78t3litIp5AKll
SGaSSNzLz9cQgx78ZuT+jcdFbnlJ9Tl0DYLHCZUsTC/9Ioghbps5LbL7jbbCoklM
oZArczB7S5P7JwVlpvVy4KeYcUJuDbW+El4dcvfc7UIn/roe3PUU+k2/cDZ2alyo
YJFv8q3AC6t/yz+UhkoxbCEzvlULssXMV7rPpfAIBllWom8+lThnjqLGRo4w0ypM
0tJ+7Xqru3IC6X3Y9dJqXrmodYWGThNge1t8wetVlni/fzgWAy05EmZLX4OeZhE4
1fJLEP1CJ35foHkfebQ2cLMew0m2lKZuHXUhdprFo1psfcVjkHjSTHx/aqoGw8tI
Hno1iAqUB1OmtLhxw9428Snu5A1/MLmixaUGMry1/xk/rSUHKyEFk7tQBM4J9u9l
Jwtx2YDrdsRW9Fw/cv5ffa3W9N1l4bcX4PgqpUwCFhrA3368FQo5Bl1ToUXwlNgL
zWyRsbOeo6SIH0cEvKmYVzmEU61dX0KChVtJyh4Ek9DNIwwKerNIuNdf3iCMkevd
JF+UEK0udFGUYiwiMnJ1P5b6v4IKn3FsCv3HggszsUzRVS1A8RABs2ZS96/lBsEz
KZmpgVn6QbkRwSEt3pJwhDbA84/nq8GV8yzcV5L6rmV3fmxjjZH0GjAcyJPkP5Jf
HVHJB3cH+uWaov2t2bnzwLpLjcoaJlU/jw+ehMv9ve28kophyH/L/raU1s/+xdPS
SAOex5og7x9zklqWXTjPAHgVbYykXvfSt7/UuLnim5whurrxPmhDVXYThizdqyjE
L7OdVDuy/hsdeD5jx3O2pgVZJDq/DSgrka64EprVRtiODKl2KZDczEGsHJ38wO8m
B/wQjAZmkbawPg79E/fh++dKUsXmYsf1J3aL2qlrHWk8tXDsFt9blpj+lXOHtO9Z
lnAiHkr9OIt0Ft84TU0gePNFleqh7R8Qliwn3ZOa3iOxjZVPOQi5zu04QTu6w9BS
CPmLZbYbzUEhVRN/RhIYkowB0Q7zk5uq/eOXLybTLWHMuSTBT2UPhLolvaoxWQB6
369Is5eZ5hxexmKN1WskM7cft1xtfA21yEY2zTWf75Z6uY9eCp9rIVDmNNeMJIo6
PCTGQzLMF2Sy5547uREuZ+F4IgYsoTSFVBSg4R8iWkIFFcZA6FpseBY0VISXM/by
5CLO8krE7xM1TG6tIC+B7KIhn03z4lq/xOOQKh678K3nS/0Fq/3ejl7NkL+TuMEp
tmTlCfDsY4az9XGkTuSw4oCrofejMS+ngSrc141i9bcJNpUMxGD+Ye3Ow50SSvLq
jwUvpE5sM86+kFyj3Cr/Vdxi9U/sPYEVM8glO4B/BOyaX/C9TL2/ShC1S7SdS9R1
rXpzWMDad19mif4JWFOTFScIO3uZV9OmJz9euimMIEGfJnQoM8TRep3vlikeiaoV
wX2c/oHR0z6U0GLIVnpW8tGj8DgtFfMD+kQzoZxMRj5qwOnXjhZ89E8Y1r2X8n2O
FgF9V7urm/0SQRw6b7RWOvXgj1uknBaQBYELTqVeQLYEf4MzyNgBXgrsMXIj75YN
zXGOy8oCUn34JlAbDL/dRn/uQIy8JWHL5fBDNiKTWvAU0K6LFhoD+evWS7j4TKV+
PX7sCQXm3DPMdaUBZvriAJOpmliumuDWaNcUEl57g/4gelPvLjogGFCz73JCxW08
eWNvaj1eCXx+/9LPUv/b7ojQIhgQhaNXbyNnfk4vwi3H7A2dao831hChuZ/XSeWU
DfQxp4KRd1jw7aGZiMkKmHUMDcC5jlasQ0h3feOy/kXynDBSjVyVr5DD2dXoyBAN
9gHBvJAe1dX169xSz/ZkxgbqKjBU/1NH8foIt2GcFC1ydx5+I0ZkcyjyWlZM2P97
Krb++HVZJOQn6zI7KMlCBGQmeM6dqRZA7hXnXyO9/n/GKVgTwBA/rs00wy0aE8Zp
DGuXrW17M6GQKsXL+oANoAxlfzwokAeP+6qXERorJJ0LpdBcfMq81y7O4QGb9cgx
S+djRLmIUCJTlCzX7iiGRQsrfvSJhjYDgBRu12LUyjkSt7LwHNsnvDS1d4nLL8Dt
2sWdWW/w1OS+lXHxyRMMFssPxtRy0qXT6DTKpEsxfOFEZuOKuXMH0UtRywS1D7Ke
NnoZqbvFCUZzXwqxzyIG8VdfZDbuVzJ4bFp/zOMVxuGbBHo1vLAp7NubelbOVDBV
06bIW/a1Qol1pqJyWit4jZ5vuaV0t0MdHGt4QooDXNFhSqvY5sp/CWuCpitvA7iO
5J/LQB1yVmeRTFcODY4Fr/4Ajzr5/ouW6NQEp36p/anWEd39SX4d6tfuX8MObASG
QOhVgUtXjF6yOYJ3dpgtvLuXW6n0A9AZc0rta8PRYcMkC3a9J/FjgXvzrFRZFFOX
T0G98WZ8UYxITgJQfAiuptYu9ZA8m7l4BWuO+arqwcadjcxYQmcW4mEElps9ZpDY
xPN2CrRgq4r7rV3LPUtsfjCLM5AKPBlIBKrTFLrlc0bcLNnJg2XlRLQ8Pp1OtmIR
a24AiTXiDDCpbIgoy1ILWhwnijteAW2NvTSN8DWCpR1YuDpJB6jF9b2IiqPgaJb5
Qv+kPNIVu/TnNUTEmpL3XHTq0PJ8X0txbHimnu68PhMkBxyKsEHMopgj0hqk1wrz
tSnG/zMesKIfzJ82r/glEQoGvrP4ZldT1p212XAlOoqH9N7vJ+726pVnmq0zEbE2
IP9+so81nvb3ZwdVgaN5VIKnHlbj2CJZr9fp+VwwY/paj5mMM0jetAZlebWAchDT
3sELc8JsqEHBEVcagTDJ6+9GFVxzVP0vbwp31/sRny0M3QY+AcjV0sk0UvypdLzE
XIp9avy96bz5mrWG3mUlU9CvMMZp9CzOPS1OlCJqEjGIEfQrvCPb4fCdu10mix6+
mQZfnfEiT+hlM5zWA7yG8aPWQwR7SpYLDDUlC+tj2a7AsOfaJeEO0TKsZBcP2GFX
Z+CA07W8P8G/MIZz5BjSFohyDh/1O4zIwDe30iR9u7gaoavwoqzetOdbsAnyUv7R
Wk8QdpgZjGQ++FiWZYGG7c2u06UQ/vPMTIrW+LbnqEJ9kTSzy/CIMmHHQwWnkCVs
3GhpnSM2g7YniFdSpyARK50e/GNU6gXUQpww28A3Ogbu11ZTcSoXdzSHIL62rCxx
eXctEELi56B3eI8ehqCP2J5tEy/ChoJVVoDZnzWnbjwM2mLwhOS9UP1OMUpcQ0vF
8zJcpHkc+ftX37xW6Jz3VdU6ZhV6SrbLTKJh14cewcoMgVKBDVaGLZEtowFv6Rjx
iTbpxxIZnOCcEha7qvg+qH110yeizQjZJgZ9A6qza9RSwuMWUg4rqZQbqBsbNvW0
8802jvHg28MVGhiyYR/0t6JmmV6j5EmJ408n0DA4nSDeflw679xs1bNcJy0VrdaT
Ic+ODnLhtHaTe+A6ATRWbWSIc5JBIfjvC1Qs5xNc+BVDD5yOtjCD8tMMBkL7OiHR
VlVTR2wmY42iE77cXqHx3OM6skFbeEN7JsLzaoojDCbmUQLdYAIF+2PdKjz6XgHG
Y3sLem68D6AHfQIRuwMZNLNzAQJ/Lt66Ssf9xMOJCsaa47ch/FmZUS9xM69JGX68
EXqaY/QC1/hrankse/uGPFxqxl+Hzt7eOYa+2eJcBA8WhsQKGcgkoyWjGs7R+ofK
Hqd8bb4sKtI9EBY1kFXyWW0o0GBI5nAi/6cCx08reoQXXKVLeASSjbLBudLOT15+
oYswquwW5Pw2ntJuVHupcAOvTHmlGIK+belZVYKOHjUdZXsv7PEFKngYXQWPsFsh
CMK1mTXlUa/IEWpazWFD5+ErzFB3JE3iOjIer5bsRF1ApMXTApjc1NJzfhho2wcR
7rDXODvik7vF/2RK2kDEn+1xDZXctcA5srA2AbF/BZrqmUVFWz6YCnHltBdY8PT+
xS/zYW3aPL7Oh1Xukw0XMZo/7mCLASet0KXPlnbCqiXcSDD3pkNHM7n5tL3F1Dp3
QLJSvjGyfjSCFNg5I4tYdiGaMdhXfZ3ldWHu5wsT5sDNNzrwTYOf7AS6BjkhFJ0J
KExCfOGydzsTfbfNiUQaKT8Z8TY7EyrwIdXv6dr7zUTB0xzx4mUt711ydiltvcYz
DT+9G4Vn9uPboroiXS/5mmVBRGO1xAu/LRnV96Qz2fuDCkHyZpV8BttH3DQMASOb
MuSHlvgWwXQ6dJ+v2CFTLaw+5phEjP/KctBcEjHxQIzpv2TAvrNEbPhyTMCqqdsE
P9nrJTufISYP3Yh0GW7OiPCKfsq9OfsqlJ+cixq3SsZYbxrbhaosXJIJE+5VOfmJ
W9YfCDZ8Atf74mDgJDwwFwjvXdk6Firgg5W34ydtMoj/9Joo2ZwVUvTNABcYNY/1
M0MpwOuSfTEC3vCiqzs/6eF6irY7pUBqYmHL9eRORlv6wZILHXqq5g0owVLi3JLv
vVyC5wTzDf/uEUjaRmU00smTBFC7Un0gksz5WkKwnPnDdD/A2Hdc8f8uR6cjKEi/
UWDdb5lF1TMXlPG/MyHdQQMHqN8JeqaTiZJnOeFVokFsXIQ7MocyHECjOITCUBLk
8Mso1WpEiQPHMM81uQ0dqmwOuEFOHJAHdyhqdF37Gd4x05yNJsoANGEhAkLzSad9
Xx2taAvVBnZug6WmEqSCchGrTXvF+ChmUvdcy/gFAkosyKD8PNx/cL5i6YOlfvWI
9wMExzXJUMKAiXy9uNscg5eww68QCJ3tBd2k4V+G0wWvvgnDuGd3IEGAJ7lN4pVi
HdasY8Cpm6MOcHg1+5g43q75det4lRPwYc3CYV00Ujgv4WirBI0fmmPJ5APeK9AK
rj3X7yr2313ocJTfHQWlKO9dTVD40GSCL6D0S5yN+UwPyuqo7BQfCj+HkWn+BIFK
Tk0hhgv2QkTR1daT9MJs3Of7vBJJXUYTkvc5wvfL5j7//nggzzLy2xTd2/2hheLX
2s1yGpgJ3bca1lIcaK1dMRT71IRiFIzFa0SPTg9o+8jMBPJv62ANEST5Q/wawoIY
TWwWxyZvlBziqtPYon284+DSd3/7H+XLxQ22FljXPR4JOk7yTqw8glaI8Z1cBa7t
ZuUnufHbwS7cdNBVtqNU+2z1TA/x4/vl/+iGF4Pn8poaGJJhSXU/W/mWC2r3H8xe
cuxR+XBjXMDpb9GZjoIKIFqLmk3K888VlN7mKdBMvz1KGFketff4twagqqIuvEJV
ZMJ+QuQMZNnD9rPR0MuCbdJ10O43526HuIkIsgFYPbIMq9Y+vHJ1G0RXnkd9Fuuz
wM9i30nulgUTSCX3pQaY7V5Qu3rCFPKyS5uVTn3bz4DDy6OtBWC4iPV2QLqwlx5F
5QozVVco6Pvyxe/CPn79nC5KOUz6vEwOq6tiD4xyQy1R16pW8POWLxDgHmEay1zR
rhtLgLL0lNSzRERgVMxL6sVaNJN94EG6kdwAfu2BQHn8sOHeQqOlegHTfFvyyO3V
6+gZ8baDybHNdHWzxAj1q3i2882T8SP6J3atUKsOZ73kEYeF6N/FdhS7OHj5uVla
NDnZLnhTDq79Mp+2dIwcBNhZXyE+dcXumiiJzgAdHucERTl8C7b0cOK4qXtVP2kT
aHwbW0l8XaIII6gtxS6TqhWZVgzPZ4lnXqflf0XpX1SE24E+hP3YgH0TOyCS7Rad
kR1OB24TAdap+JdzoG5oEzUrokHqYWojAK9IROuuXgimveLeO+F98+fckmWLYg1Q
1zw6R19BaBsSXLLJLpoNu7osAnl22lBy/FgWJBn6AGVBocA5hkxfXmZc4DQIZhfN
jBy4MN/cBduVFSltH2Wh4xcg6lDV16gOPV1AFoKg4fVdsv/g3QZbm/9KQmaK+OzC
v/5od7QECYvEMzPpMVrq8f96eIklIcAb6otxQ1yjQWOGpUQtoJ/K+EkCnkGjJZ1S
CAlACDlrhZJbARBoKc8QX8jOEADOjqtO7XGCax6vm0EBUAxXk6nmZWG5n4nGW486
WBQVvNMcRSUTTHXKlY82o02LgEXq0lTOhUc523ijqM7GXOCkaG5cxAS+frhZLzUv
XQ/ALkNjRt8SgHK8wOkaUdzA7WTEd3exTl5yNYwDSNi9o2rsp5HOi1mzsx6mHnd3
7DdwdV917oedmjCgMN9kwzZ82Ij+xaimGmySsuO89UpL/MChbalVU7GpSThwwDYD
spsuUEwgFMlB7CVKTcZmOhJs5AAPz1ytzE/uzr2jZz8lwQBgcAYterKCqMPOUh5d
oJBKiTDPlr3u/qx7+lLiXuMPpoGpbksdrbqKwdB7XD9YvPvHFXJhZJ/3MsmqbKi/
94a2VIsig9b88ECMiVE1zoHELW1No41B/YXnUxQuq5M2Ek0xSldCifWiJL8QV2H3
YZKz+dppoihv77uF22u7lNy6BM9SHl6N0Lc+4KjmobyInPRwym1CJDNgyCcO4i8x
xP5WyWNRjHjoMuvjI5+0+upiubYJChJ3wcUgxuWy/VnGPizlnEVyu/br+HwrprkG
ZyfgA7ZVDmBb6FaOmVH13PUKXjt8HLp4UDIL1w0C6R0CvvQJYPFWgbhe2MIDN7k0
QJ1lVwae56c2L42jaZu039g0TxuYcQuJfr+0QslSHKP4buuCbNCIkYXYPkrxxS+F
NVy4jjx2C4OCm5P2THREz1gfpvvLljKxT04eALJWq0oxtXbAKxnaCRgEbvSuBe46
APR/5YoMfg6+NVd/j0B8EBiNFvU55MQd1CJ0Df6LhD4vTSiO3VoVx1Q8jmPzHbs+
tp7BTlfum5doH9EMJoTQugraEUfZgJCeW/I24RbCAR2DQ8urkrA4W8898SptRGvs
fggEWzPXjAkbAAxhlOBkPYK4V4K+cWBBGPVa1cHMZnuKo4lS4uvNgqgbV9arsVxJ
iSkjUNb8/Pxb085gCgWWoRwmsiEJcyZFWOczt4pxR50m0uu6O9TjTTRu/Yo1SxUu
SAadBbULc9lFclx9nrB5D4D1mkYJV5BEGpz12Fm4ZolxIU9GctO2VQh8ga5cFurF
S6zzB904FGx0HjNHcnqZgFjkv8txzaoGR3aIanGzweTVwW+chNtV+jvTeDbKDqUi
iciBIv94ABy6aTbTe8ZQwmjHYSk8AT1Ise0oBItT2dBb9xkzXCfNIlOU8tCesxUp
PSS//0m/Zf8w0dwVGS1684gtL1HDtBN3OP/oEDxfripRoz/7v6jPMFaXO8gAS9cA
s9oSADIUA8qRCey5S8/0yVXYIwJpz2yzt59FRhZjvtT1IYqqk9gyIyX+hQchKgrY
xfaCu2oYiZnPEtdYookJ+GCMDjUqbmKXqfzf4VyMXuSnjKcl1K9vkzwCEGnB9Ued
V8JStDQ8VLwDl58ioPrwf/bHhopB1uBtzADGHLTdGQQL46zwdynPRnYEDbr7Njj3
OTeKZjsRWL0CXwPJPQBrMM+V19ZqWELEWK6Bt69C0Q4TvGryBkthSX+1eWxw1x1C
VEbB7ne6Xw1ir69qobYhKQfVwULMJooKHpPaIws4OyEejjfRzvjR5rJvOgvl2a/b
WTO8oGowuFpJSdSe3y4gPpu/0nrjqdRQjsD9sspwfGucCzBpzvEmeslt011v4gex
eWjfFDTG6GInc9VJrpJtqlXSCBJrFdjxeKt4FKFZlRYg9FNCnSzfbv5M3brTlgYK
48Q80wKLQiq+F6fFmt4LHzplUxc/1hhKP5zkqpF8Bn0XwlYdUMPo13P7TAD/ekN4
KWy8J9N8ON6AYNkF5nYbajYK54qUlpRls7jdD2WYRyc0c7OMiQeDvtg+KtvlfK6B
IPZBVZwqoqkFqNdF09oGdQI/A3gBhQbJYusS1/hDQfft7EiPAfDAwfRrRqGp2rmq
vu47P4QmJLBGpuroseVV3SojrCm7lsNQTgIlMQUanVqK11agkgYFCMxsqy7l3ZW7
q3rCnq8ajEhe+X59yT0IXSwyd6kJon5wPbeeHyZQdkZKzBBZDsc4x/LW7S30freX
VHL4jrjlqzRfM+9o6tuFSQfVDWbT3jt1EBNZ2++SF5p/RIW+Eb9OLcJRyWcqvWQm
X8+23gb4/8aHkqSIN6lT6nDhhsbOf68LHeNTQVHXOKJs9Jm1DofREQNZ3Yyo7Gjy
TFDi3Ph0tgojhFdEOqyM4mAFlRngQ3G1Ms7XJNtdRioGOyA+pl9tqZm6X5YNgTd2
h/2kxWtqMphPs8aYyc6HE2WB+dg6AX7IL54Lg0XihR93DzuEMaCK7pruHqveDkN7
cm/e3inn0GyDVpiN3z6NINuspksj5WBssVpXOeKykHfnAV25+iUCA3R9o14vTz3D
AZQ6ZcX7UNQMpeQObLUxs1e6q6XDOhhgxu8emklWfhh956VPLRU3ZnQoNmdjI8XX
Ij0177EDVPyphaA1aJNKQfVphKWKzNn4gKovAm44SvK8mivdI/NRUMdfRgFOn6Em
/TSf1m7jy4hOKqZxt2GgXsYf3MTuK3Jn2hCLA/snzczZGTybMbU4d5xZyQlGlJfV
OCz39S8MRzf23dLrv/Us3P+B2s5KmvAZqCZdfNVno7Ya+++Qio04cJOUYO9y0VL6
ORT19aR78m4YT7xExv9e6c6X2KY/7Nthcq+mrDfir25wCwmwb3ZAJEyNRtxITjpK
ZMbl1XojS8MZ2PbuAEyhcsQxAr8IgLSK2NnGzxla/cdl3eSMtuVnLhm/yaz+UYTk
1x6zOeRw81xKRyE9YXWaChPpOGPbldW7qjOKVOPj5HVn8E7N0aiyEUyzhbLYOLG4
G0Qkypc7hv5u5VZYoW6lVbacPaksgiwrRQFh7lmvUuniTPFUTGfAhbAOzQnnQsJm
4uXgdMGPJ9QSXL9Nj5owZjH+CtWlYRq7xQrclAEMAGcNjBXzY9eL50SYh35c0VWW
ZgnNuHecJvuD/wiYn6ygZjUyVRBKdeLGo6Sq7XXcfQ0xwj0SHZtqNe8XcK3b2l/A
sbvIBHvCV0qIyG5ijRwzLAhYXVQKzZJoTNpggZGzpje20i83wSWDXcX/1rww6tVu
74XGoRy/TfG/dTD1qxIGGBpKjUOGf9YsHNcunJyfiklqlfrIpL1mpVJWQRR6D008
1AzfI8b19yqvPrZLW3CDIsFc7YGgLSueKbSYDbWlyzhgOkFgc+MR4e8+wtPvbOl4
jicWlE6YOGkz3mlzNVjsfr22+PG8l+HFyg7hhGYIi/xFHT9zcRirMhyLVj+twFsZ
wZXc66Xro1jpHzt0tAYiqmZwyHhOVIvrrFvjmeCXvZ2uqki3Dag8xFjBWBbz0xkk
jesish4GniBv4XE/mtMx20IZw07+u4OMMRN/MpvdGZOjGLYkmtZGMGvMp/eIZXe3
0cXDqcDkuWqiwNhtjZbcGkEPJ9+E4inhcBH0Agstklm8RPMu60wZTzr2t8Qmdcoh
b0rV+QwIfSbmgZex73bco4Id6B36PdsAzz+iUVYRtlBKhU3FHoDrA36dD5CorXIR
bnqAWE6zvATxbHpQk2ZtExrR+84+rw1zuVo+dPMUBVi85qRNQ2hJe6irKakuL+RX
ozJSOHxpzISMFrov6QLm8yHansH2ohDG3rvrd8QJTEj0TCoHZSvu7Jibhs8W2nGp
Hgnf5gBf/XAyqFKEb/bDdRsoi6HhRBNHcGGmeK8tgV4e1DMFz6IR2kLFQM1AyeoJ
pJF31pjVEeqN30XyTr9hr/d4qCkOI5EPStgQZTh9JL55GJcLJDfXfRpBlboMx2wC
yeA1nlANRzf/q1Si1lM48WsxE1ye5zqGrh2q4s+Qv2kI+T3IvcG6JM6fUjVU9tIm
UU5ZDRCQYqUxgDHQLpNBFVzWTNtO2uyqeu9yfodFkBEYz1DAJosC7TrSiIW8U6hr
q73tcrruqVG+3wjb1lL5LDtz92Y4XT1fYe5DKJ4kwjZM2PTy+vtu8umgvpUqinbs
lGsM0ixV7Iz91+8NBblwQoSKbroD8zJQGatY4vkXA7qWk/QgqwwiipSGBSGliDcH
fmN6ty3+AEUHm6nfc6xTBEjJX5kbCCe5XBfJgJLpOPfFkfBO71MV87WHaCfWVQWK
du1NRRsur26l3QmWIfrJWVIvM4oEh1I5rA50KW7LvyDc7Il/SL26kT+kxJnWuFcM
heTIKJjbEN6pXffwYdIGoseO49oRT09N7Aq5yOf/wggGMs24eZ5qVhqKrdfMr1KY
WKhAidcDq0Eu/K8iI6B9AGxeTLs1StS+/G12rCb5CCSdUarYVL/TefvxExK9Q9NX
rLM1QbvWX2v+fXAzEw6egmirRLs2/113heso2Coo/s9nCWBx0PS/8PPGKyDq9R8w
sn6J1n89fgZ820sDJMc1bDCE1QF1TPnczFbOZ8N+g66pijcoc13KzpBaXZTqAp7+
ZNJ7mCY0wfG7DsUXT6OxO1O87qKQwUueYk8fDoQkpF2xyZXMcukuj0/jzkY/AUUL
2StHLXlU4L1MsTXkfVGQ9MAP85y0xnVlFiBYN4wJiEk/wbJZr1EAk1R5KyU5HJjn
/7HQwvLrVKhcT1aXuex/aNPpp1z3yK7Sm4DWVasu+RDZdw6do/8Ud/EWyui7Zck/
9mm9wTZFRznvp9067rr7daGh4vk5fJ+0OvFJ7oRxQ2LTlqwL7oAstbfsiimJbbm9
5JkNAY5hk9SgKuCKMA9k8O/z3jfY6ektgc3np9junRWnKg2l+n7WgnN/EybSqtOL
laeguJq7xGlrS9ShRaC5QvQ30qurtQ1dbBAkYrUsmEl8n5M+pkUW6Oa4DOKDtFq3
uu9q3KrVemC2bTkXnD0/AK27cXvDBe4GbOMiUPQrAUAK9aVSYpBtK9gWfaVs91zq
ZbuCrdA54BiJNeBhyiRT/jKTu64IcjpZ/pxNOUnesYf+MPbmJ8RLPxHgVyuRX3ey
g0KSYsfBpTWiHJhUOTjuYhq/jEuG0iBNSHyh1KrJiYh4AlND55Kk4zokURxKaXPA
1HDrWbEYYbguKLUu8V0pvwmRyKbHlJZnqVMc+ZS8kH2VOEPOMnvd5Ix/uXuxasrx
fZdiG4JSAs4CCfULmYcj9wiSDC5YJpkBAuVCWNViDK4gc3n4nWYYSVTAzw+437Dl
5TgFhp0TQzgbqrYAum2fwSi0JYNb9TzRyrwpKXJiVVcEbscRzfF11NpLtUWpEZTS
LZGk+9Oat8jA96SkBxSMgUvD9YIaMi8gmkVZ0/1zcD2oIipLAQzygeHxgUqSYXTd
1imtcdTDY81SJJWV5f6QF2bpdycJBlvqFATf92e0B09yhJPSyEbrJaJrzsV5oODo
FyGga0PW0z1E9rnH1g2/QPAxPy1AaWDycIwtMe0h3mURLE8pFPnRMjzDlDy9BdLa
ybf5EYdHV/eUhgTpu8TRrQHOaT0HZJyk8ROFuyM/FrmBQJMPW5WDODfR3qVAVulQ
bE/6ekJ7zOdo/Nk3iA2nxPu5Y5SZauG2nhyHiPr5gysHszfmZnVH8MPNrbZ7+dym
ehlrrNVwbj+z5xrry99Xxyo4p4ggWMJrnAR71ih0bban+zOyopsIQr4RBBzJilIT
Io3vIlt47ULMNcSNXQjxETGTpWQPKfTjgfqfSgRmL5j7+8qFz9FKJR21HjM1wDQ0
M1dhzDi4cE34U2E7Ua2hpnJqoZhy3wDprAw1FY7Bqof6GX2SO4Fug8UY5ujmEFJY
n//Po+rkaOaD3FNA9HvT3wNQGYBQ8+1MdgrWV10vmvyDnzu2w5sd/Zqv/xjf37cq
7lYdXhiJe6ay6sDSzMIVWxBsHGsMbanxZm0ALx5QJCOvZHxE4EdKkw28o/VzP7RG
sJ5KujoQB9/bsoflebXO04ptuN6WJqnZYCQrUIMNpufYSraJZKdBzFKPOXTfJHIZ
/0IvimNXbcQSG2cShlQ5J0AhUk2NsGZ7kRP5eGmn4F7/13rWh854nqpcQZYxD+4H
cPWVKhx8Hu3EhZSdAGdfUBoSss0fNF6JurEID65a/aLnp1VPZQ3Q8yHVp+/HAOdi
S5AbNFCKnS1j8vmhxia6G9mCKj8X2xz7UEQMcxlFM59mYru3rguT9BBu/rZDdo0L
Xn6C3sAYp1XPs2esfaeB861Bgm+QOemHEfyWxjyEu0Ih9B47X9mYLZ6Kk03m2+5B
0s4VibDufUUarPio2BXYhP/TrPMlCAY7XnA8xUjtSytJBXJ81k7apoAvMFPdu2S/
7yEPvmEHfey1wFde/BxW8Ds1k0+EaxZWQKsnG6wG9XHwdPDZ4WLo+E0vVV4yNsGH
i/POOqD93w7PYTbb0045VE9t8GJTRGMUUCbz3d+XM2ZkNYXcCHANEp55u6JGtGtJ
6ygaT5byD9ECAV9baZrNXz/EDN5wmrN+c/qO91QUhJ9f8P8sJK/alNa0FE/+Lics
dMKJawz6phs7izxJBp7NkuetOJ/Wkg+XVPlsNDKxCGKrzSRMnQfo88H6pIi49gOS
CKR3M2n4WhoWTelV8HBBj2CM6aSHrIYVmqUVTefNeThYrdgO/SI3sL812o4hbzlF
/W2SJJejMcin1tMkIVOH13wzJ5RBKP3cqVshHBF3gfAYKh9/HG0loXKe5IIjt/HO
3BzdGnjOq5oGwx76KtyzK0rL74NB9HaweoIx2bSM2+rB6ohlPAx92dR55U2wz6Am
xOctfUSWaPqGWP/stuIoVVU9a3YgxGocb6Pt8UjX/ECpDfHt7y+Pe2X4TJTxwznn
iq7pkii8RCQ51iaUHt1A9G4RT/XPdbP5yacQd7f7RC3WwLoCpomiqgaHheymYC2+
ppbzSLHnxREQ1GH2zPE0VK9R6PbFjfTsxLHW37MfB/u9550iCqVO/y/Ouc1iTOlo
c3PA/FUewG1AR6T7ejFqbQP8qicLISN2gmyWzjvxTNOf52Kn4IBfxK6V9XEB1Y6e
toGsQLWsDZxuD/MEWq2H6Bqu7uukNjVqfmYJm8XFergonwHp6+j/NjFfQSoGPKJ4
Qy8d97GJciB4qA/I8PWx9i5fwMwLUXbN/h0kv/7mYAxpegydqEH+Ihe+NY1IxWW1
6C1IEQUVVXFpzll3/r8aWMkxHFLoDn5w7zjQnb2j03ODG9y5akHoPk+fnzalKFPp
SUORnRfojTG8yx5AzMfAG44My0ruGEWGKgi9Hr8IpTBG6QoX4iI0LuPh7C9DGxZ0
P4ao3AnWJg8sd5qCMqlUe/GsUIc1T3OLoFFkutkDAg53O6tvFGUKr1LN9QLBzkIF
VxmwSzMNWy/RbmFtPjKf5kGJXFynZQp6vg8dumS/+294aGcwPdJlMFleX/RYyHH5
ZYCsguyoFhyu5jLWmlA8DsSbLup2TvlNKdSrv/CBHM6fIeHAqqIVI9BirP55JTIz
3n73PmxykvHVIC5zind2tXRf1P7bfC6V+g4lUuVWl/SKLFiI8wymVuXNW2L3klWP
LIlwq1h9AuvC5mRlcFvxmjJ/0t4GLTJaBFQMjNOlDme+JUpbpBZ9nw9e6rUrMmCg
nRebPttZ5NtHZY+KbRR+aIovBBBSmaF8Wykj6hlgEtqJwr7qqeU4C3evAEHl5M5M
iDX5ZWoEqsGLb2H7e/J8sPPo4tPeT6a14yi0bjZNaWBzrLUHle/z7Mxt8smS10DU
/eyDdoTDaA0e1ocs7DnTVOBdycMxrrlQKPIey3pO/iHdZlg3day+AtbSOmoDPLWz
xJT/WnNR9Mjfauyhdj68OWSYMGtxy8eJqiXlfNyE06WzDKFZRApfyJhYWv+UCRit
n3ldNY3SnwQBs4zlRxN/uzvQuEwhPPqGvRgFg/8lyiay49TQN2m0DJCvFd9sUfAQ
yomyHX+7/3+WHaKejaG+Rm3iOm17j3Iwba52k6e4K/AE8TdYnsRC3NR6BmYma0S3
cKjbvgGP6L9uF0qlJD1G3ITW7pAFD1ZgI8wtygCOA0UytCU0h8dm01dEVyi8weNs
JjpCxZQXTK0mbCE0/xyoyvlbC0nobf6PWOfWXQfSEX2ybMFkDYupH+EIUJQgURLg
ZqdtTEuMRRCJQgHXP3bcFNtyIrmXYOaoO6XcrVaxW37P7TzlhQVxkUjDCPurYra/
j1xEbhIR/ld33oscCrONYJfbtrLbtKmHwg+au7N5l3gi99CqYsN/bCci15JM534D
5rtsKa74OUcJkDfftQnOGE7IlLaeTUeLrSbAgDgJsWkq0Pu5+pCgS+q6ahq7s4o2
GwCmwvUeJCaB4PMDj3WTPkZ5nFvvJZ3kIoLWtKdpgmZDL7Wm00+D+8cFgZAwjWrB
1/G8BnAYPbrMAe/UUEUpo1TBYO6uM34oWsotaunwyww6Pm7N9R9fSY2mS6qvii9k
YvSPt8xgBKzy69mzweGlalqRDc0BYbboSgk6uSpNAs4/XuUL9B8k665WIzmrz/Ru
PJhSMgCKDuWApVbd3r3fdIlEvz3WA0xZlUyBbeB4IrZUtsmcd88hj6a+B4AlCvxZ
iUKTwOm/Nv6hT90q9yWWkXF4sHpB0wxCqFR+rOXEDh/B2+IqHd69xicEw7IZTw5n
oKWbMnfWInBLT20peVPFgI7eZTxr75QIqMR0OqEIYdW++NvaYUYUJYdyx3cD/cpU
9By353lpml9z2E5JSteP4JA8ZECJA90bA+RY1O0iYBA2uJpl+dyh9U8iChMTdYpL
o9bCICSVFg73qOYkgjGTkUFZx+j/mAY9vf9hHoahfj+l6QLNcV3N5hJeXTL9Mxdi
zJFLDgTrYw7zTysS6/3NxhzvhleeE7wrXA9lw6SR1dqcbFpfbwAtGNyd5GvSKox6
Qa8Heoqn4QrPkZDwdkyAXlp6np+weC5o9jF3LmQgStAu4llHB+C5NiuZ233q7A2s
ZCqNz1oxQ+eqzfRmDpC+UxXaOiqSBhxkrSzC/7lE0loq0DMqM9Xk0i1+Q1HYJFaA
SNRDOJx5Hlw552aj3NJBX5X47Hfg9xHqmKk1a0+pSshZGAFPUqLCrd7hqhWsytSx
l0n73DApIh3Xf6Eid9Yvmh2Yft45NRc8e1L1RmOz84zXt0EjHGPSNYvdfgGAKaAd
5DpDgvMSJJf7aUFNw8G8dGfPaTpV+K/MF1fTR5fjZexaZo6o1aot+nZp55ZTldgU
QnuTYs+0OPn3DmVlEdjtaKDVnajgIv3O5S7DwvtmgEECxJ5KUob8UUsYQhRd+Y6/
jvy2qsI9UIRHDtpMkIIpNPyhzGCES4pN8rOfBu+ofxvrM8LW40IXbHGebe3thkO8
aSj3K1KO5bNVeQ+pwgccsnptFGxiEdEvjUenIljk1fiUXqQ5xcn6rTReYY1Kd0Tr
7s2nSrifuSP3rCWormINmM2xrhJTIK2Abm7rScL2MlwW7s35+RbNFA/aRsomxfYc
dQ2U2+Yocs6jcPmg4CbY4AnvTqSoLRgRrY8N0CK6nie4a1vW8HrMGHfSmXOhFLAO
EGaurcJvKhV59zEscsWJRMC7xPAq8FjcyWgJ/OUkeItMjcTW1xfK2kp0lrRV80KI
b6NrZQG0jsNtTRkegjMhHbaVT3nkv3VqjcWhktDPdRP8y8x3c7RYU2kteqYi1lRm
GnuaT4j5B8cUu5uKCMF7OmB0BfwAVEuE74AFtDN9J6D1XYCcqGeUDz0/l3uDZ+hv
269BcEkbOdkxgVn5ee4t+ygj9Ll2mpEv9zyWPDBEpxueVf8F2G9nPdN4srX3CW9a
NFmDjGADtG1oJxO9bz9HMjc1BvNBU4SJwWhA+ZHx5jXi7VD7XxV/zwBYwJqRIpB7
/AVxI6tDWfzPzB17Gcxc6mj2pfpoyd/4IAsQtt+03i/0XfKOPRF+UCdiN5nsfhhX
hC03tKOsgW9R+6XLx8CWrEpsw00t59Us0C2QF7eQOD2mPEA5EzBkCUNYF43WLpJR
Dz9Grt6Tqwj/REA1GGd6FZc8tvATka3UM+tfWeCwAeHOC+BEKsJZ3NKdCHrqlwCc
gJpi9vBPFqIGraOvVE3E75ksrwysgLK3+cyLlNtmXjAhwWHJcFbMMjB7ti+2tPag
8bG/uzZ3swxNs/PPL3c/VYE5TbcWdiUgzkt5VVRVoNp/1wGXPYxWYw5O0uv2Xw27
yF2LSLi7Latzlx3UT/0KtGO0KlY3VBawq69Wo3d1U5hc49wXbMeCcsCOe0tYeZUz
CXSiJu3dJWuTQQlFAYUc/ej+t6w4/TPgsSUlayXd2Hwu1nEJgjR5FbV7cL4feHdX
DUafcFkQE3syw5YTM8uNALCPPLDdrwUW71Zc9bSYIqG0KCXqn3GDy6iBsmyEH7/t
w36wmsRIiBoLnoYOSrD3exrBqnKnOfhU60gK6oM4aQFqTMm8WkJGjA27IS+a/H/B
sGTCw8bmryLY91PTMJwcj4cA+6rMguczLFsHXRMCG5y/JU4estvWyXEwcAzkw6Wt
8eNmAiOraRxPLIeYh0B1oWlRGgInwuakHx5FGAU/BJ+cnzidzXaVW50FZz/U0YsR
5G+P6hhzHhHoUooJj78SSFHpIRGXg3xt/GwWxzzSllcVvugcvKhw+sSPE8tYMzMa
fe3i7LzIALqAEpujD17U1pMK+1z35tGwKOgIz2aB6WE6n4GCdS362EXvdY1pWvLs
L/8wwY9Hq2FIjW7dJBlSeeEQHrLr4JUUTnuiwD7WAaeYtR/L2p1XERit8QOvNu1o
lRb1ivDcR8VQABVvCWKtTARz0StN5/2GD64weMn470cjT5OMVFaS2u5KCIL3HGYX
TpDv4AkkWbHtvMVRKkxqM19XinaES/JyvjLGicfoA2DWdkTkEnqxQzJaWGeAZvqA
U9+HKSRRTMEIar/ZsAMSyTTrMn2DhQ+F5W2iqnUMH0gK5L+AOSd9bt1zuTZ9PZlF
uSS1KsBUvZ7r9BOY0aOQgn+qwO0lKIhUpPTZIX4zuwOF3QXMaJLhkdVadu7J0C/u
BqYNMrJw4872/Eq0O5oCNPtOiKJvQUNIiHvqjr8ynPKiZ08kfzi4crQuzHgjMJk5
i/IFHmYSY4Hq3Cl6aTb4VbzBahDLspwfYhKkYzg32XH4QpZ/V/AMrnmXV8l3Lapp
Qu+PCm2P+Mk7+1BI34AG4ro/aMqdNH84mE7+mL0k4HgiOirLPeDnsh20QBAL42dA
S9eNNqPhkW5FxDJ8Dh7agpRjhfBMTCGntmdLx5Onxzb95tRRQMU6oY4NDl+HCMc5
4f2nx3TM96nj+eoOQ0CknsSC8mtv7aKOYzWtW2l15fUiJCeOqmae4jCgAahDm9wa
R15LFU/c0LbnPIzdamQlBIvkazT/h34AS290Mq9/Gnse1eRG2o5Mw+Lt/O0OtICK
o3q34G2jXt3yMsD9oiiiGclb6/GjOWCdnH8nvF4j+f4TtOw3C5TSRzmvpPR4vXtg
tRvd73r8B6lVKRqYQqU6IYj9XtywI2PXoEcQ5IB32EmsANqqNJWsGVWVFfbdRvtI
2mTPFngx2DlPw3j+OkKN3pkAbjYyJyBHBca0cBOY4Kwtr1yX+PQvB8k1xVa4B3z0
+jHdh2jGizQgwlFGoAklEn2qvy7b2mhhrCKv9JzVJ1AuyHMroBkGE8RZuFNcVKt1
SDvGybwky4T5TtBbRXFOtUT/sM334s47LLHHdKp4h/3rHwjCON07AN9HfPu5AUdr
GkrtrrB6/c50GkY4suT88mRLmrsnMAvvNzFqsnjxRcNSmaIkS+SUBdnamQva32b2
BmD331TM7uetj3Xd/XcfDMNIthoq6VNxWc06ELuCx+zqYTCaZTmQqUA3Aj4Sh4iF
AnLNWSijSfTpyiK8otzYaI40WikNWoWd1hbHtGN5LtXx9OnuiB95Cu5W5yV0HMyZ
0gf4a9gvksQFV+0QZXBkdxCv+EhXhD/3BNBdne63iBxMebZPOwHY0Pv/jzk7Pl4D
+9hC+P0hemqyhzCXe8lPbARNa+n2E/4A39qnETJdKLvx5Nwo++M/kJZftTMBHSvy
a+V2TkHMhwLz1gAENdCm26iylvPBHhtP6sc06PMtMXgZ66ZaFVWchIC9neU5i/eG
Zx0FC8Gg/x3r4MOxoYn2E9fBZSZuEMvC6feUwo9hAtDmahSHesgztqwsWH3ihP6F
XWMBeGjdzKbX73q3BEoASTF/05f+uEr0rsuGXmMwK8vKssyBRz1AGLkHgtU9t5lv
RuhLTCV7fio4cqqRkx3plykDbnE3VRgoiJjSMDlZx4IjlupaO9XgCkqrIAJwa69P
KVvDTjQ/Bq5eCk8iCkJArAAUm4qQ7Qf+kwfzeNKpbd1DH9DuYE4lj1rK2LMS2dCy
otqhxXGMKkU0LW2RFI6yUU+aQKkZpbEHn8ew8Bx5ByaY/PGrKWUd8kU7IJ0uimqL
+TZSABLsW15vnaeF7u0wF/i8ohIrohycsYpM0KxZmr6gRS2D1L5DJsduRfcuE4Td
z125ODKYE4KVVqHuXnnoiPRT3DPI0aXokYnPr7vN82xUK7uBkqUOTLd2RuC52BD8
6p0m92JBoahHpVaeEIu4c0XmoC0cxGw1+zMe0hbAO+D8mmmk4ODwX26m3OBA7mOz
8TQjBY1pZy8inDUJqJIVuEOpHmr+bYL0G+Bztl7gYCmR4xj/TOrKQKVt2vT2bjaI
/mSuSWgv0fsjVB6CURyM187pQZw+nwJoLU7UL1rkLWAaxW6tcC88PCYh2+ALgu5F
UfIuLoWye87LPGbviwGK/3eBca7sJWQ6Lu2oD70hLtimCQWDsPsX1Rhee2wJwooR
EfLAAQIGf9TMJZZ/EdH0ybbPh1eqU3V3lLQXhG/voCdWYMEg2PqqSvOJv1TIxw+j
VRRxok+8o1F4BcuARl84UXmvuq0PX4cfaply5FplvgPUhjGA3cdhf+iC8W+g6r1f
uDliRffQZB5HN+jpqOXtygBXVR5fRagwFDciYXtUqnT+iUqYwJ4vof35ep9pYT96
NcFT4cqntc99zs3j07YvYRzBDvNlTEnzpyIAp5cjaP2UT+TE7dND/gQyMS0AVRis
PIENC0K7P7drhJJGWjltGlvU8VUAYW9B0bxCzOl6b0cgBpM9NKzC0JuSI5nPSY6i
Jz0m3worA5Li98oRMjtc3Y4yQCS5qhrNWRvXzelinZjVGdg6Oehd2esuzpKTSLE3
EWX/fRsbF1V6Q3fM2sXc/w1BhTKugdD2WXSz7QBm4tn+xnTpUFB11n3FKoISaWI6
h+W14ThlKPZRoG76ctV5OLnhGfrdge3NX/DsoHGskKDUOkDtvkGsOe8rQp8MdGWo
z5AZ+gE2P9fzj02K/4sxn7XLPsfvdAv2PTtsm9Bk0XabsAl4PuFsPjhOizyNq4zp
gK37e53eJKITRKoenaEkVUKfp4yadHyDNEbRXpzWKYucFHzD/+MEZ7o7W4qnano7
1vv2YuJc+jbaVErt1o//nrfwY49CeeoJIzUWE7d986+Zp4XzzIPP7mSliZWkM5la
ixf45BkB31Kx4/6VgYTADkFY+UIFILnGDTTBz1ZL3nsjBF/dONTX3TbEWOIVgIa1
+7WZmkODNMlRIXDU9SoHWsZBck2vBFETjaAqvGrqlUHxK6UsqTcR6H/VdPAmoFxw
50S7YV/8ruft7wfKtA2XNSAmg5ZCH8x0NzLViN24s/SY9TWLMdTBEr+KpYI85Ecq
0Y1zvgJVg9/bQDTMKaaztowsjyaGFIWxJuPSs61H+YUyJe+TbPklNF5L9Lib4Ijl
e00H4byHmXtLaDbCv6wxfxuA914JrMrOCMrriqfi/cn9ckfsvVpBeqal+rznp5ni
CjarQfSsSc/76J0WBJEUfgMg5+0UHemC/C8FQjL02ikSQmsM2bpnhBybuUEWsF7Z
Ap2nSuG2zpDNfz5ZUcq+Nq9Cb1TiM/XyaY/wwWbhfTqbOOGcyFGgpey+0+qB1md3
VMLVGPz7/itr3sjjE/dTxOQC1DpE0kfMh1jckuUZNw8evg8DvgSfAUdGLU8Ep1Jh
8XcVPN2NPHb1iMEZr6UGSz8T5MsnyOCgmBNSSHRjp00Iv5xSwNt+kYOf4Miw5Mmi
pk5/m0wtrrNB92x96diX5MwpsTQ53SVZNB0rbYM2sk/rFteeL44wWIJXqw6xIGKw
7Fn7PGMGZIQh2wu8QqpKJgwUFkfQmSAeL4lsUfXn6oGlUBLrb/s/VhgH862FlsZJ
glL2Sgtv0WvEY0rRhGY/czP53g1DETROjmS5/Haziy/AAgXvyEvD52UxQrgRGYNT
tz1mneL9lDWteh6p9auYRkG5Qsl4GnaIKyFHFNdE71y5iXmF0+aY9mrp/e27lEcd
5zBMRsoloUKJswaWmE1D7VUj3ecbiNGKUql8k6k+7tdOJqzFxjIL7H86d0zxSJBV
40eUrhinm09mISjDlqxamM8364wq7WaGaLr6MYq1hddJL7rtJGGOwRUK2zL6OZET
09d++cOuFbf9hU+dtzxHpbI6NdZWiLpOpSEhDkW0qSTOkCWY8jsdQy7c9mwhoHOy
Yt8YLocydOGgCdy6OxWkgnoBWtGZc5OKMq8/OiKWnGFAhnFkhhIHMG32dK+ghYNj
99I9F7+PclEyGubhyjh167xq7u/TzimTtxrgleexI9RdYacIZ3/iSfvvNRzHlyPN
2IJ8lUrbcJ0aEUltWrr5axQ/vXhQswojlObQXQSDEPWiVWjACe3GJ/42HpEU+7Fl
YhIUWd0B1oc5mvMOjSW86ZoeOcP9vmtio7IsUo3XVpE7kbRUh2WSN3I6wEgcSik9
xEnryR5Gyk5k7WsS+5/JrHSwUOlL+PSR/yvr4/3gBDkNGLV1WYQr7Bps6WGa1hZQ
Xn8DkC9jcD7XRYhKj0+pEHLaSdhUiub3VtdJmW+mKN1fSPLIiLWaqXvAMOBmneOU
G0i4tD5Ug9NtIAUhChlqIG06+8Q9iK4SVUiU7sf20a7xv2O4wrXhi3ifzjYv1FGk
zFkAOfLLIpLa0A2tQfxP/RAxxZUvyww8utPNNaDoaECNo7HYsJUaS0GRpdAwpcf8
pMq4lBAsbZMuntjhVNoPfdndIUZB3vSueIN8bCZeeq3ris8oZyHsQs3XLhZsOmxt
Ua5DFIT8i2Bgk3fZdBWudbOkB/JRMkeRb65UvKX0op48mDYArbNipHu/xwoBt3Y0
6m68eO6GyLzf8BJyneesWXAfXyK1FbQ/8CwsTmiWOn27IV13Bp/k+T+TFmRsQSLV
dC6XUVkX4B+0fd8uzB5GYD77fbZGf6geqATpXJWQhUfCwkGf3QRSwTqdg8vQO+mJ
qcaZQKML/YiHw55b8CPRI0s/tFV9vrz77NnNrJvSMDv3E/qOH30DI+DAQ4RK2Y6x
ierxdvztH//dZ2aOQnOVC7logUGIEoDmI8kwI7ldQSxNqNsNk3QN7FJcGWfEhY/k
pK76YOcn1/0ZX/KQSayrWqKcLe3qRMqZdOFcDnxtNpAV+qLOzXEPWIJbAxAYB0/p
Yuj9PNr6G/h1/jmBfSVgsH8t85vIWMWe2SAb3Dl1auITUy+z/VxU8izvf+G+O3wD
82kcITx9dLEY7koOpSjdXdf0eJ425gk74FtKX48LzF0J2weR2rVCcuQgGa6Tq85n
VsvxDkhivy02yNcq9+N283abbiRmeulB6UjwnhWBcpKY4qdpMaSEmpixlsBY/PAl
mHJpVxgS5MSS5jxo4AXBt8yGrPpLCBwmfRhBEyFLUxq7cAftb4OL+v4OP92gHqyS
7hwy+E8Q4840ACeDXBBcfZZwg5Hwhfv4L41tAL2n9cTp/0ntRbMpzsR0PvdwPYQy
UcpJxzoTEh24ZkEzzltN6mrpct9NcFYWVSxT7mefFphnb72rQnSUtMat5phptuEb
gqg5w+bGTPHx6HTTHVg8AiVHJKBlGVn9b2FC5x5ymMfgrbf7vuO8TNRzelzWj00Y
+1s1M3JKJUYa5dIh+pjrE7R0o6S7yOQv0+UUxBaUHA1VMcmZSX9hSczzPpzPd4Fi
m6HesOYJ+s5gfwGX1IoAJLmvR5SH1IaDdvPvVHx+9F5utopj48qa/GRIuKL6Bfj8
sEz3jOOQquWtbMgm3uMmISBDoakCq+5krH4bSLtOhN8RhSMFvBKhx4NFBdw1VQqk
C2jHCsL70AJCOB/lX8xMHaChfoRdmeAktWHP8xwwgCrGSb3Yo3Fpvz/rNLMSKHfX
eu3PcAqhPnMKy6efXx9yHiQjTxuGC4QJh4tO1KTzzThWvFKJLdG0SRGrYuWWAD0P
dfaVVQkbf4ZQIlQuImza6TOXMkux5UPS3vDWGZ6JRzBkyOws1b62WYYQYyfoidwl
+2AfRITnL4GDcwIaVsO9CODHTohgoojDVHrrhEGmxn7EQIqsjKax4vcc7ivXtyH/
1aBZ+j99g8A5O4f6gNASN+NIhvP8BrMmrjor2+RBJEndtj+wGFvAIS8b8HiBgITm
dWCehEVFKNSQCD0gWnGBbcxKyFEVuRDj0kHaWRJiOBWMc62ddOF2N8GbNuA6dRdV
Yt8GhsXrjuNQQvmkenHpnRHbIygij2S+gKNP9d1o5ABU1XRVHTrPdrxBsQ1c7a4E
mwMtCqks/2FDNRHfWCGCTeDO0zJZWhxSgwftR3FBy1nVI81kKWGQ+tVQWHs794hm
xI+0Ye7qTnnzIsSyCTJ3XTGXey2esqjR6mjGirjC+10DKw/xxRPqEDOdlxU926BP
u730uF8vlc34Y7qG5/tWCvBTFO4RdJTQ5V7jf+Vf0t6/9hW8sRzG2oBPC6DbHehJ
m0Ubouihuhqtto+28LNzS5ukdIBxjTbBZyPOZlCVII6rmcvTDcAEadTKK4vpfP7s
yXWe355GzauASOpYuEjQjvVgkJC2OqZsrXm+JJjXTBmITUmUe4NgDHexwJFNEOF5
hIepztfO+GNXqTaA2Y0Am3tSaShDXr+WZ0cNeJd/BN/QLuCz9gmAh6EMNeinDP9L
yJczUh2txIWypUTR49wlKRpFv5cnoj97vjVNrgOIAz84XQ14niSpGBYwkUeO0ma2
bAUkk+t9V2QBVKu3Q7WdVJ5Lx+TjjyO3zTI5l4R/DUzaR06kEVFilc3C9hwCCY4a
5h1mtUYKbvtTLBPnZuwS4A4TlEdo9InKniSIbDlOKUDMbGaXm/HuLJMah6Xrtk7U
o2aRpyO1spBcMERXUeAiF5F70vO2jltDg1yKyny+JUNItwS8IB4tf49jCb/6W07t
PlHBKpC1ix0qPxOSooRpxUrbXGxpnJNrQ87CKgjnDvgoUdGtmPEoRsdv2Z4oHnV3
2aI26JrkqrCDMnKz9t0P0+utY3mM6f44ZLl909U47N0PAgTyiDul4NplFfAiP6F0
yA4j5TOlA4pX3H1WfjjILKL2jyp7NUDm6MqPF9ssb0TkWv0CIf0wQze43YBPXImO
V3hEQLYW9xHV5SVlA/FeIic/bdFtlDbOtm0C1ZTPpOB/Eur7M3vFbkmCB0+iJr3C
ZvC9Tx2/Kp8Pqa1jDDcKJu9wlzd/bxmIbBbiUCytf8/zdZYVOA4i8Li5BtEP2xOH
2K1mhxcWbswwgpcC3RSIu3VvLtcMh+anPbjWIpbHaoEFoqyMiLr+1m5uU4lAblCh
YxpPOGCN8JyrvS5BUPxbW0B6d+vbAOcjaWFBCk+tBcdSXyb9+psRBo3jk0KESTQ9
9jkDrNA0GcF4sH7fgoh1I8ijP2rbrA3cWRzx1a4Jr3nT+Me9Rf0eW9UW3dwm/6CX
w3/GwS/oppaAE+vdzULop1K0eNFZBmdynPvjJddAn7H7oDorA6//CNiiHE1Iezrz
cDUlVp5zB4JZ5aNT4T+a1oU/SSCpotY4emOalzgfG6sybMdyLQuNDhLTcg05QjYu
zf7eC4iCwi4/GOk3DVd3SHd3hqcOyWAxcO3PJzk85RHZd2rQbdg6uw1qTVlrUv/Q
bNUaInlT66RHjaQZshJlhRnEqYs35f4i1mLlZu09kLA8tx6fS5i9SUk7Scx+gkDF
J5JoYVXZwU49qgp2AqlzxLYyOs0FQ+poMLZklk2mZE8qMx2tEpwiYg4pQAbPGef3
4IEAZ1YCtqtIIXYWFyPtUa+QFKbBMKbWmgdNxSoboKEKMz7H5E1dQsS9AkOkKMBV
OAtXYJxv0hMDLkhzNqkJom3PLGtfUYfgU/P3xPiNUO5yvv9xpbETmwEdc/7mV1wU
Zpl5vj6yzH8m6sGwLQ2/B3kwxF0vMG2bz8Sixso0FstSmZ+I3uipYWa/u6mBSkvS
0NGB8ECupQPa9G/5k8RV/hyCNnk2M9o6cmhea9GabPuLrSu/R39JoPMXyEc1y1kk
sDx6yFexj2gGJ6D9Zu28ysyyTOJ95IuqD3mTyxPnyef2zeYWxKFFyMDKw29xfgHF
KxvsWr6IwQjkFwJKjGjdtGViRlDmwXElAz19AD225WE5hHOTt55jv9/DivVtWFzn
S2Fvme4YKtpFiNzFrD1VmPOkUMTN5Nln2KVy6f7JWX8zNfuDGuyTbRSR7wUnRPMz
IW+uMB7dfVv2bVGEe9KBeETXKoBKppkD4Y6vjml+l2vOnV3wSkeX1Bdan1bxM/qp
+jdaavmbTmTXSTpnrZ2dXnaCFTXf15ZMj2/enaeHVnOhY3Jx6By2KrJz2WCSXG3m
uV6urft2L/ARCZazV2dQCm4YJkkc8AuNgf6Uc7aNEVQGTCCgzqPyj0Qv0wsaoVd/
UIA5KXCPC03aaace8loiE3WESdm63cJjJqWl/khNvicAt6tm6Qpp73YAWuZChjxC
Nr9nuwe04B25pMMO1K3kpmnI8N5xfdQAt+tqDK78HYzWyjq0EWyGBbo/un2J7/kh
UVWZn+3Jgvq07IeUldwOZbGpRfnMHSHVcxCQJQa8a4wdIyk469M3nnmVBxDdTRap
aONRw4QBdkMcHCubDsNUWCClOPjXgc4S8Pb1LtBDjVl97aeA9fl7KQxvhRmnfikn
FGTTryRfpVLXxl4RgxEuiWWbkGc6LMH/5D2etoXhkYAYnevj5/VLwIaT+L9uiZkO
OHdx6eh52+6sfBC3ngrIlqD0ihP65d65jfBndlu7iBX8gL4QsnZSCUNQyw4ICrRb
65OU6J3FVt95g6NYujo9gMitIUDZ2Cg3oZ0fjvRvEWJC8nKHr6QVOtWWuzUFKwYu
9NJMQcsj+PcnLR0tUvTVEKFEEM72qjO8CkmO26FUvP5oVmOviNCFIRfzA7XGmfnl
EjWYFXYCV1ujWsjnx7KqYkbEzo/YJ5tnCdIXJjQyy5e1GYDeBsj0H3r1ai2IwIPj
vZiqiwkigzTFXG90lJutGMxyddbX8pAtqwPMUYL76eHLulnMxjIn3AruNAXtAINe
LVhm5cnSejGcKSF9NhVZAzNyz3/ml7HbD5b2biGsXSINq7aDcWAanbaRJzZdKiDK
96CJNiibu3uS6BqhtMrQv8W3KxL0eVc8MmsE5WeMRdAFxXoOQeo92E5Vjkb4sfya
npk/dWXzMPzD6Fxqdgfng+mcRW0ik8MEYbMeAOawIoU8XCBecX6IRNu2pT92Vo/3
U7gcV+S+DJ23RlqL1aso46ODInYLDRYuAjvWof5gjgTl7PxaaoZphB534QqEpWwE
fF7BZh7nfgefL4HOpxliaFeaYDQUhBkvioZZ3QXA2327Jmat2kZSwBF/TvqwK2K9
Rf5MnHzbJAq7oZYFreAOzsVpoObJQxGaGGok2E5RaFKqZnwIp45UoezU4lgsBnYy
VH64cWFk6R15nZ6NPa0ecem7jaxJPOc1a7/g1G+skIsZy7i3qVQuYdMQb9dTaOhI
RLpiDyCYdZ617wjae3MhP4BfAKVy7/HtbbTGVnkdkugq630mPtAMCh8g854S4GmH
VgCh4xZfcG3Ve4xsR73VO+cdfx5+yz8agx66qIDtppMSpl+TeIIxEQYXLNiqh0cZ
Vu66V/WxOQMWRyrF21RdsgB3Sbh/lG4+cY8LymQcGIr3wOVQKqURu/JWVkBpg9n0
zPd6zSyZGWhDkPIF8MKwKPWW16b/Yerp2lJo7isGDiSvIHT0086BwL6UdD8Mx9ld
Cq0Q39DnylDd2ko1lb3l43cYstg+nz7BdyGRVdljm94LKe8xkDMYCbs1HHLlgAuc
fPo7kGalh5mB1oD62U001wLx2rk1jWKOYGo02TZgNOF5VsgrE5Tn5AIN/wdJLig6
3kj0c7umIQWXPfBe0TLE2XWRk1aXj2aoLS2hKewFuT9UgvoqAOWqAIH4X5E1nw87
2Hyw76KsE0oQID4qI4o7EW54Mt74u94MGC5r352WSdLuz1pW2O7MA09zT6490ThZ
tneEnNXjYZ1bq+KOtsHk1GH+8uzde3yauPxvNpQIaOG5edg8QaF9R0ffnhQA1e96
OFIbNgl50OXfRwG/0FfMt+qAFMxyBaKTrYTCnjGcpHpy1C78rhyBZAVkYDp0MG05
WzoizzUEr9pVfnk67YnXodkX9xe/k2dgQvewCrx9S/IsGfxAKLAe2F22JEO4GEdp
psW6h6AQQeFj9+Oui6DRwGCYs5uyj0HInh10GtpHz2imcUONHy8Q6yqD+fVHHS5R
Xh0r8OIuFEb2XYDg+0jsKtTg9/YUvx/6GuC/L9yt7SIoNQX1j2giqpUnq4QQ4Ukh
d/V6UNlmFJO9ym2or+RkGTqiIWaVFiTuRpJyJjpwDktjghU2q9If/wNDOIr5DL4W
ZFPNzOY/TC3BNhZJOWF84kjckpQBKx1aUk0jAW1S3n3P0AewSCmmm42L0E2isDeg
Ll5uF+OuNm/BVHVz2f7v2VgJq69123J1s1dAS4otllMYAvUlfyEJtzFO4rpiokYt
Tc3aY8U7iczIuKnrgl8eFQs7jHQxDbDfpB1++VXmmM9wla1+qB4wh/Cqg4sH1RiV
lFOrkSc/Bdp4R4egh4Gvz7N1LHVebGZcJi6WYgwXCW7SoTirPFa+4jxm620zGYic
eix5HkIIfIXJWjKlMXX2WSpZ2v2w0GdLzJXihSw5I9tu2RYKA0n1LdfUXjxWScq0
Wwo+Vo7I7VOlG+KgMUac97jCoQlgPeGAeX0Wjl0kxG9SeUjvVaG1Cwe1BU1iBLsm
qjr8+4IYKTX96pbBEIrpJDYsvAAJta7HdgM4L7AZllazLjlCRsuB2INXhW1pop0h
0W7yoe/bB120HdHv0QTO5cLqsWjLcdZRI70+WbejXRTeS1p04fkzkonVXpFR0ceZ
jH4N4EoWJMy0/ZGdpi46oT1S59/jTl2gGxcaZzCKbSzY5LHc9l/w5ePaSUJ4yK4D
poN9sC5LO6CpvfsTx8bSe1g5QdZ6GTMQbbjJ0STd73CLP9Tl3r5WOr09yeNN7vIV
zFaIoOONDFZb+G4KPyuCGpV3t3fNzfVUroERLAFQTRehGIRI+wMzWswuLGtoBhzP
4gwLWrko0dS2fwjRU5VGzD+vyPZ9uMCOTmPkbQFxwUE+XaWxh3veaNNkyxV89Z8u
74YUyjmiYAtwricpHmTr1AQjee45x780exe95XFjo+qsB0qVxksb5/9Dg+HimB3W
IgoOPNnBCY+pZXIcJ4J/qVurEblcwFqSTOZbX/m2gNFfd1SdKRfsp9hEE/S2TPgN
xkNddEjhGPRUr496SqcFzFwQqGYu7n0nBE+O6O0peo0mmrgM9pC/VuSjlx9BeAOf
kISyC3jxG1YU9YrUHj22+23nh23mBUo8ojX1pwFJe7OKa+lLGDkvAqWbnmIQei3o
tG4B4RsZF+NHOaB7NBGUoiv75ZlqmTozNN1RVHyYFinZiAjyOk8P9KePjxQMJblZ
BxWkrr/KEfcRA9m/X3jPlOzqSUuXNaARSwkzem8uy37OEgWHKiNQ+226STnUWNXN
xVfdx1guuSeMSMWtI5Fs1ZjtuzMSMXpOtD+O7FSEYmkKZwlETkGK2ReAuHbmtFWQ
FdzrA80r18HywVcuQEKCUdwnv5gC3bm80geQ3Q9b+FJZ+qPjds2HYhcB7NlJPqWV
wuKtQStCvJ6UN84vCvLrb8pu8cRRPmDtXLlDDZDYoz0gYGEB9Zmm51JORrQgdy01
z4lp54DxmaHutwZnl+NMqpo8KH4hzqYh3qm9iOyii1LWPKoSA59PIq3HCUn3rqGU
OFA1Xe0r4ujnmi5vfW8Yg1ex0x2T8vVW6+QtpSTCEQZpyRejgQPOL6zj8kWc2tek
3qAIrVEKll0N6VoKPMITb7Adr7S9lL2Z840kf+YFWk4ZaIsmSjt1r2xzxKewoSCw
P6ms7Ax4142FPX2Xin8HT/s5dAKVw/OSxtRASsRQD1Zo/wwCU/LA55YlBmdPMoVW
vz5vPfo1TLTC5rBDBDD3/0bcQ+kBrSLoaQGWtoEUCu+tjm5sGqhe+UkR7b0nQUsH
rf2YEXGvz0r/S91I1EKkwKMVwnOrBhQGyCBTtQeetV/FQp7xL1QXEEgCHcjIQfBM
6yxRFV0geEljuH1xAp3LBdA5ivsOR1mow4drYZwi91GYRUsD5bGmqJJV9u29ZlKx
+wbg4l5WaTB807O4+dBulZgxxLUh1EUx5l738uwt9tvC0MRxXK3goDjBCz7sMRpE
C50PBfmpDSGFh/8C0F1lqcj0yJ37aFXjF/aZVA50mXbW5Gy86nhipNLF2tsAUJa8
fJ9tWWaD3jT5plgwLlkmIH2a1xMG1VbwwhLta1iNrhIdGqqqbIsapvO7d8+HyDHu
xU6sp4YdTkT6vusCDfvPshN5OVsqUsdl8vVRx5m1KFGO6UoABAYPleLPRbXGXXRI
kbHejnV1CXn0rL+BzOey1ua9YvKHswtIwfBt6qxyQc9kVAcNwPwN/o9s/aL5QgFn
siTKsfQU/tqNI2ZZungZfMBnvmfXQeWOtBkhO+EPcxpII1Qd3uEX6a+bUQ8jVNe3
gbrU3ih0mfUEbOkqv3P9EWm0jhWNt+PlI01yfc7s9qOPDEqPgHk9fY/KpNl5EC+P
i0NNikViFsJ+hLwdUdxR6Eme0t4fZ8HUTEHuKODVBv2nTRhLD97PYqv0LsONYesS
QVXNLakbL41sv5BQbwZHng2UWkWavrItHtePXOCbsvdyE+HlldTUxTaTeC4VSB24
8Hb5NeMyMzy7sdyL9SgKayz6bHipn3eYKXlrPppnxNd1AAyYqccEA8TuCJDohab2
qufp1QnXwaJeZ+/EhwALFGhrYJ5CFEqvdPIHFCLGoKCdz4gkM4Sl9WztVZOLA7Fq
R1CBuBR8RkmVQ193u2Q1yZLL7v4UDkaZf5DS1BQr5rJIm6l99dcq9as8PzrcWnY/
Ml4SdBauQ82BDwqvio2CpJkjO8J80lc9Vxcffad8FcSSJebcD7TszG/zqYdwHKiJ
p78YckhNiuAmEv/TRRgDzqPeU20T2rK04NtaR+DA95UiAG/zClKE6KtoCzSdKY+n
/V+7MriajE8YSJzkcsL4pM/cbWyh5iwp/KHEmnOdMAE/e8bYNwhBLA9n22CLlhcW
PysO2R87EyKSv1544QriYwl0YWthREZvP1vSDMsQT2co2t9dqBB3Q2rE7JqwsY/c
mQFCHxdPJSJVc3Yk0jpTFl+o7Kk2sNtvZ2zDmGljS3TYuIMS9fow2Vc1ALM0dBi5
kDsesllhigLFG+xH9CA0MslUNmFN+77wwuMzM73T5pW/NfComNABCuYWm76Pg20B
UXgbpLN+2mrDjsKe+o2MQlpNVAHnF/6JdykuSzqpYlB+J74520q3YlO9BwmtU8jw
yvFygLfHBdN/1Z9vNDsvD2/1EA6JjBm0EpsALXvQub4hg1kpuT2CKTj03hLmovae
huiwLs5irvbh8RFnv5nutUWdGyF+MPeku0D1Z6vrBs53VNyLtzP/ME5La9ESMtZ/
YesK0G8iwOROGXz6K3oRTDRhf7K93FzuLEQnRMIwfDXpqxAIhvc0ip/5HhiZyZ1r
CQDU+/P3jwlG2QudkcUTMy9UOax7JegGXf4oTKBTUGIJ3HZA7lULkrMSKs8egbFj
c7U0C+aXZXal2w5Fs3Mn23enFhT/JwuFKpbjhxwgpN7OXGbCqK+BGpZF7JNp1q9v
LyO8RP3wJSjlYSTUyqODvf8xt9ufFfOPLkX6fVJP31hTJri+EFisY5jTto1eeaZX
u1i3q+n8mEWOXKdOegL5z2pa0LZCWPqk0n8/VB0lMziqnGPOFV2ztEu3PrI0TMbG
fQCBMfjpRo9JFkw+92EjVh7qcEGu1dbJ8z6HImpo13CsY9GgrJyjrUafx/IjSYoj
uqt4DqVN47kBgY5u0vkYKsNxFlN58jnbfAm//j3oY3ECxkrrHUPtkNXphWCE5t9u
eYlbmBQ6BlQhTLeZ6n4PNtV+MZZCX/yPejWTc3UMsNfEMeugMITwNe0cu+J0ccQV
I33rmt3S2c+Z0mmgtS45YLFUu/h/ex6rYRTsYP3U4xzhtD9rjwvfKI0enFP1Szv5
t1JoltYC3wytIREWddc3VrLgnOiuTxcuqwMVFL5MrVrtPuiUBfrYCGQXUJlLMwOc
naupq6GrVvg/syBluUygU24DuymwDxkE9+PPWHlXXUTQIz8TstNE3wK6lSjcy2r9
6sngSivg6Zd8tz2hxjEN6XZT+TDtUTgtW7ifq+sjZYwm86DsMsP7Iz5csYjkAQgD
tMgYimiN7zzCor6w+ews4S4CrgyPtfrbCTDS/O4Q33X5T9xXdPMFsVRoJmt8f9MF
HPT8bUywHFPG+u8Losq8XeGg3UB/dH5kBH017dwIwbPto3FTiQYbI8i5V1umMIZ6
4vqj8HiS1KtSf5704HVILqAOQOaDMg4G21CrPbVXepRf522JR59HjLqtq+361mqS
qq3agAXoxApBv1B/LOmeJvI9vN0P06SEU4QPiYRe7dgk+02xrk25ay8szym2QbUj
VBZB1fDBQtaiuSFA9X/qk0Bst+LSj4L3oJ8DcIM3JtE8JDa5C/NSMLu1xhLnDC9w
TH83QhTIoPNxMUiYOvysePACYLWRwsPcQtyaqbNETyjYM8nhFLJokiXXe5i6nDVm
cNzmzol93NP1NRWryx/S7FbtznFVMnyKXpPNeOuGz3hD8k4d0BvyAaedNyX1/hWY
2fpcXszcP0BySH+aNJhFAev409s65uo4iLXPFR0ZeNdhQ1ozsijGCHucxUjvk5qO
sdnW/VyGXQ1au18W0IxJ5IebUsT6G7BNeQ6h1CzQ1GnnHGsBMOAl4j14xtDwww7Z
55Jj7lSaBR0upUNjtuJdVxdDIHWUjdSmWSCPORXVynzOJASq6q8D5viWhiCrG3Qr
m8SHskXeQsHI7IdUym85MGHQRd0vw7YP7BO0avLhtDMeSwU2JA757LrSieeTuPG8
ZG5LQHsB4C40tyahPRlelEtmAZVuD8yQcLyS97cc5mG2BgizJKPArFpogVx32/QM
OF0B6pFvVz06IS7Lga++yp6fKMRCdpj40v58FqAT7WV5w3T8II+5Ks8qgNCJJpji
zL00iPR1Me09JtJncRIonb5lpjzn6b+Ll2HkP0ZnSitGIkLnjyUgFS7jIp8xxUyA
j7nB0kiNhpUV5srfq79AWkMMT//qku1yGq3mSebtblKV2Hkyry++rMJS5PVaOejW
FfFWmbG9mz4CHckcsn+U4SzY3asp8kOKhii5Pk1HgCqtk6H73QBkmyvtaKsotGgx
KdkL5z5Q/u3rUn/lteJUum27xbWns3N/BF8cM9NWSyZIU+8i7aGhntJ+oXoN6tcc
TnU21OutXV2yAlv5x+Y9OTjt99l/RDQ1W9ZI5DZa+YoRryaQK92GXRwpn0wB3LGH
hS/GaUId2vkYx0figzYh+yDJVjS7sh+MDOdZoajal8LXZtxgV7f6VIzlq4sGQV8k
MP1UWmx5c0UTtc8HyL2BrH7reJKtLTtz3h494LxT88M3t/wE54Gf2BmaKL4Sq/dO
t5/Fg9IQ+GRwAwgOry6kqIYSqinaocfheATRJnudvQrdDYpWry4FQ7y+J/3Q06Wj
uMfVTZbA1C08asf4ts56BgHgxX2ZMgEJ8dRK2CSXocHfxOsnwIaL5f7opfnr7Y8u
O7RbLpQlKRW5jiJDbsHPYoMCZCYVc9LqAhGbgrGhNXsO6qUFxNKSoWOY14hlU0Aj
V5BXDYyR7QbNRauB7KJuaNrCeN2JeJbgEvF6DqmYUyBWQWw+Nkktqt63Pp0O5Cvd
bQW5WNRPhkkg/TVyqSrrV2P3utVzay5vCcqbHADs0XZIinkAq7dSOtqwLNLR230k
EO9jIJtJARa0cQsefDv2hMRu62DkhGMuP+rgfEqVcBnhsjvjnhp7ZgzQ7/0FD6F9
BQlKjAX/qeQAp9cw83SGc0tsklgQuEUJN8OiL8umFoUJ7a21OpH0egurFVU2IV1A
xmwwvgaMpQIE2tRo2fE4YzeqANxmdhPb1Cdgv3b+Qa0U4PuWX72j6v4fTygrlQaF
m6v9B+a2UJqqY6K2YzZlqo5zo6xU73DL6ABgyxQN+1Ouf86gMeq4XSnQgE2eoDpk
zjgTVwAMCWJRf4v/tuMojloVIzMvIOh+v4lEQbUE+W3MKcYw0O5ERqtzcefBF1fG
Zdo/vzaIalKkbSOM3OlNfFOd39nWm7R/rhkwbJ35eV6TMu1EkzuD4a3gUnMxjxq0
8yh156Ib4OfVx0NrQLpoSFKKYVmGFpehmQdxLJbiPkryd49Y1WRx9KBfclw+03Jp
/u4MWMcLeJ6lq7HUVLuxgRmWvxNdPM9Ryvlwe3DqBM8Vs/IDyskCeGo3Ri14QdAn
pSvPSrJ/W+5az5iv38XIV7jKXE7s0tez0yY00KOnfVIx4BNRHwnRtvOsqY90Z6fc
TgiLrs+FbcUDpbh9sCoTB8MPL7vw9J+J60+Bb7uzUIehCMWD40YF1PsY7rkuw/vt
+9D9njl8oMeudG4n6E9rOkmtw3ZvMBJrgO1tQYFRPQSm8+rFGtuRtYUY7kzX+ZyC
dGdiAeJx0cvcqPjmoDLrmLoh7f22l7SF1Nn7UcRKwBLfa+Zohiak02OdmMiBWjJB
msHLpxC4k+kIwgy4eHahExLX31o4IYVaSI52koG/wVKTsbojJptS4b4Vv3dprhih
k5IV873vXjWG16Trx/xbaVL85DBNeDCzo2BqEZywfqLQ9M2tWP+LILeBheFTTl0p
5/zKrVvDkLbV3VhIYAxMt6ZovM09VH1NIXe2e3YOmLcElgN+we1dPumZoT0suvg0
c5bnQ5BUUyytvLKgFf8oQlb7XB3DdG3b2N9DpdFXTWmrH7JKkgTJ1mN7T3/hcsCe
3c+lEYghiFnAQIzbRfMJZ2DA2Hm6aeGtflqBgvRRb6T44Og8LKRDPicnDG/Ua8z6
BpBOCRkX04AFPNGQQyp/GDKUAoiLythDOylY6ZkkFI5uFKqSYg2yrKS6AmNrUiBV
DUMF6CDlBbyJrnRMVg3cZGNlbu7qJEHYk4qR3mlR5SWaCdTJ0KX2Des9H6PXElRM
WnAKO3nzUuZ0HNs5k/gX0OYfL0ZzhLW2Wx6/3tLJgJlyPXvkNVAjJBW6Rw+wLMvk
ykOkiL0M0ouHYZLNtoEvqBVAS8ApzGIoO2YOW7od7D0tGu63mfmt0wC0a42xAYQe
Y6vNzWgXNFQIyj8Lgi3CF7mAsPFWFubCV3drkaMZRXBdsCFSEEE95yygFZTD1rLg
TARoG52sGO6p+L4rp11BgcdNVsjqIZp1Sy1SNoLuwoipw+7iMxC2mHsLJJWAaLw4
MpLzHn4DWXHwKPCKpAdGNVWAwxxAh6/3Gw7o0khew0g8O7zguxkBFEzY9wt7ECty
ZAIAKIRvG/kITeNiSxwKeFw46DKEzvGOvadgMv0quaC5F7JURb0jWNJCrDaqKOn8
cogzGAElDQWU7I7qzcRpNDBHter5Tc6l/RiZKBjwGqQcFRm9CtMYB9n3ob0xQ3li
oMWq+g95+cYYsn87ZaR2PNk8fDn9oAR0reUuC5XALguW8vH4cmeL0EfzLg6qexA8
ui72tFo+96nkI0SJjuIdvXuNAgdd/G28aJeFa4qxvvHz/MJAiweR7OeJOXlwoTjp
t9Lme5rnMnvjJa4AKxya9J39qv7sPgp9J9Lcu9gHIJd1czlybbGQOAj+LRDyGEa8
HOf4jl1NLl8apeT+gRWHCXpZ6fp6ZPxya9g/noGrkQcdkLXe2wnabhUt7D3fhGvO
svxPpLdTJ9+jgnTxWwQ7mbUTLceo2zgS1itgQ6UCcvt/eMR/JC96p0ZCaGCGLyaZ
vhtqQin1sdhm5YwdfTj6cwmaBD33OQ/ByGslL9l6hjCHyDWAR6n/bxGqAb+gUI83
/ebkXWLAYhgdsDdrUKuyybPVa1G8708YANGb8DNbmXxDSevL1Q9QmgmQdm86E2h+
tl2BEqFPsJ8o17fcgcRxbFyOg5ox8Sne+dvkGYp/xmjZLL1LNAE+B0CcKGIQgugd
LMaTcGGABLLZ+JjgQLnfdm/jp4qZXY4k64fl4QbaiAcJXFi5JDLD9D6K9rE2oF2N
hvQU7hEpEERzTDsbVxjlNcn91BFIzrrMX73WtgaJudCxjj84GhedYkSIWVMmz0pr
yP+LlXNXpBxaTgYPnkn+ZdD7xDOtg+NQrr5M2LqTUg5EgOi7R3w2ZxOEl/dUQB66
kN99je6CIiGI37fK/vvvT67IGzD5x6w1oadESvf6qrNCQEjfOCm86K9azmyCwMD2
3okk2RTb7CKqOSrfa+VqkbirjTXcYRuFriiRJgPcIWbDfzquWwqEtFOkBgZZCGO6
XwQR/xSlkKMuWZIJxn+eKDuPvvMnmZnZ6ZM7vDK28u36yPnCUKAJDYV8GJJE/WF4
zmX1vusAIh2bitrMbFolkh+s8+x3j3ZqOjh/0z8zAN5cM2Co+Y3K3fYzlzNVMIYh
+mFpzEoO+75fNd8umShGgvqVH7lz0dgEIKk5cSI718KzSMEvhm0jimPtWy5xIuCI
VvBYRl1Esfi8pWYQEoBcdPJI+24rhn5lY2KqMg899g7DPJ6zDWTSqYkN+deQEGjT
j6EnFXZ7nJyC0w76n1+QvJ5D7aHNIJJZ2uMToaMkrXW9dy3ZfHeub8amLf2MIK63
sykHFZkWVFsytfISjt+XHd8xTbBW3BH+/flCbvH+l9w8bA++uzzUImWtBrDFhF31
xmA8mKova56WzmNA6R3Qpy16x9N48ObHiKmjETCaRfgkkTv3sEWDDJ1y0jJaV6pw
BkLLZULhx2F5T0+igyN+T1x8Bf8e9dd80iRoKf+7mLnH06Ami33vdda1uJXnPu8d
zuNJqO71FE6CaiU4YDPGKvv6VKA1InQT6zi/4Jwpig9P3psHT+yzu8lrbqX3NIT5
q0Hng3VFEI3MWjymC8qkBUovZuy3ZGnjoCJS9I8xN+bRRUx1/HWC+2FjXfn+wRE8
unbSssP5jhQcw0f89TK4R3NFcK0R/c+g19r179X0H+Cvk2xDbKNIAhLr3JuehK6h
TjUizER2EuAbGRAGpetUZncwzQC4nnbwo3yxSPW40i9WgAXw6uW887W9zTFj4OBB
zKN+brkWtHGPe9riKQTwktuJPFbhNJDX6cd8sRHF1FGqhszRdqS2F3MI9Rn8BIad
JdPnkJrFOF3F4goS4G8TvGeFbG81dJ7iCuZxJuA8Pq6El3+IhPoQLR/5cwkoGhfu
ytsc4CbU5mnuSQLELWdLMTmvd1uDSkEoGBHLrA8hGrg8qj/7u/9eoe5yGrJDz3gF
CrrAs9yWf+pSbNdQMRqzUcyEDvv3S892l/jzQPUU04yL3cYyq5jWkoMgU5pLwxYm
eY772kzNCzW4UptU+dHzV3lplLOoBrz528pRh7CXnPNhCLyMwqL6WR0cAZIJi7GI
dlupgNJPwkjQo8CzPNcAi5Lq/rn0RCcSX6eKtMCbx1srxHb0QnaH1zpr4TK0wk0U
FfPrJcrcTRWBjPVbCF/W1xYJmmrOq9T/iL+ZK9EL4mkB3JZtPkN1hD5aJE49lRPI
gaDPO9PgeRqgGYUcGnMJxhJ5PL/n9d8q+eN2Tmcr4ijAL+QvXjz0cbFTHdudOwZb
U4nfsx1BSIh7pqlcMA1RQh/cihNnOV4ahe8xnQ+FfyTtZ/KYAVLCCbrI9VuuwRUQ
uEac1Ulgn4YDoljOMq+HfOk3xN5vvpz5qtvI+8cd837KW9glQuUh3lBmAPeBAGi6
JsHqHtNpI75q9VEpY4wcyTOZaDg5UV2l9Usr1XNFOqWV92FxiDvkbbpN42fxVeUg
2wTLRNaF1JQLg/qbsKA5PUJ6c99hOjFqyaXIouJf+yaWS325XQPXdx04/ydPncMS
0r2Fl5PI4i5v6KCd7+OFjceXzV9tIQOyNfybFwcVSWdPt44wYv+ddet3FuU7J7Lj
5EybRvqkHxsqGpy1XE+U3p7+aHZLNCLML3hLa7qxTnlzTKB4JtWz5vLfg3emOavb
n8fJrnVEXTu5ah/zbyeHxL4vSr/fnNsKfvmyECsa+W4SBHCiEVtjI5OSfT6xftG2
N39XEzGODB4ZHNyE8u4FdPAx1jYC7vQUiHF48gIb1/FZKAB//owJffobEg8a2s7v
SNxsBqkT4fkffmdLb8vokjVS2t1Blbe8P1OnJ/adEqvkD0lPBzxbWoo+A2B8/mh5
qSVpWtx8L+O+SSLSDRpsSgiDfxiCy5ls/MEHP+z3CIk+D27YWN1TN8QHEzMzhlbg
1Bz1hvY04pRoN2GIV0YsQ9ds1G/bvJxIfb2VVAZJ7sxFJy/KBw4fGOtrVNyI0r/p
nV9J3p377P5T3gRhKY6no2aQCaGzi46H7N+JVTRKEzwdvHWRwJIJGCt8b9j+/KBS
cdYi3+xc+WIpBPxN8mEzJvm4j1SpGm2qCXudgYRfqFt0RNYbIA5RwIuKCRt85yjb
CK2SXiGqGacV3EJIpq6i24F2j0AJ1iwa7XutHqvpcmUHbvFlZgqrnWC0yKkLv+3W
8L8f1m2xogwJudt9amvBVwzSCOxpyBvhix9lEejHD6x/toGdUEjwSnNRlMOud9o9
OmXFwywZp8Lt0TZXuswtCuKl/cjcG+worKOlD1UMyQvXak+whR3/vqvPNM0Na7NH
5E0wNYV9Wmg8cBmFYtnq8yKLkkDdWLW3sl5l4qcMXRUjZPhoz75z6/+N1rvhWGs3
g3y8uiAzsGo1leEQwjpQ0CEZ0ZLGi+TJlQsBfjhu8owqrEl1PoYjXZBA+rHbenmQ
/TpBq9qKVQwJx9p32dajSf8Y0INfJBkaITMbyy0Ga9h3FFnX9mvu6EolHDFPVgxT
0WBNKoWCDY9P6L5Svs5DswJJcFE+qSUOzLPYzcFpeMJkRRt4FVgJJyL6oulrAzqW
liaT5MDe8fX2P/Bx6VqLo3R8Vox1b88dZr+5c5DBQSTAOY0nNCSN++gB0jbYX1Yw
T/A+0cAryzKbFgy+ge7RyX8/5EI26dNBREEndFZN6Z/P82JSz8/46wVV/DmGzFyl
S6bFLcEffenM6Tf5nMD7edVwHOBP+VbM+0T0lB9fLygR7j1JKT58BRYG+NqYsMMW
EfTmN3AirFzBB8f0FTHRjzuBwLF0zJMp+aGQSGybJ1URUYlV3HM/3EaO6UIqrwwU
t1UREquHZt+CaNK1QnaUxT0dsorP2hdHXJE5WU6eYYV+HmOr1XRcWKJVRupZgnET
/c2X/dFML2OdX8mMSEcA4di8OjNvVR0RrdJNK6dQMWJTTMZQKxvxMhmJCJmP3Kkm
2RoryLBr5iLhysw3WXIGce5IMY30LQkcpUrpc2OHfjk3tprnq5J6mxfefjKJKu+r
d5D0GiP6eDd8HekIYa1ZR8hFPUJD3sEzrrVEHX9EcTLnomFI2mOH0feRIZI5RlEM
7XORc0oxX6glV1DmfdVG+++/HrpUec4iWp0D1OvV0OXw7hCp05xeFKH/bZjhJYNU
Wphg6I8wRT0MjngbcIT4bj2/6T6AWdBHTIUT0Wr2A1sfHWXRCsMq4YxfqQBgJexS
6Uw9bXNviLxf47Cp3QMNNG0jI7JbUlFcRjoKyWx1NNHD1GYamaIXwhsQV1qJQ1WE
EorQ015rgi/gTaLcC/WhDGOzSCiELHE71EU2vlkgmn0Ly+6HQirvFKdL45N9lfYR
7HHf2zl3gdtKj6LVcRkfVByd2oP974pXpznRd0aAp1JR52Ji32HCgTOYZ0WflzJM
PVJRYgS002srH0HB5dBvoReaE8dYYUm9lturxc5LaQ2CF9676lzaISlJPv+EvShO
BavpJbBvzHtmfxLN0XI0QsXs1GpTs/YCRGSGbPrVidPlqCtqnftNkS2he6jG2D+I
mvi4EIF0ZLmTJJuxDzuC/YU4dVu18Batw2zAvOX8PaQ/uw5udCT0CZraFgveuhPa
3nQbYcqYvcPpc2uwV9W3jcJuwn6ZtDN8aVqt8Nhzq+gqystTOmK+ejJiepcK65zt
TCqDrIsC+Ors3c3W42X0bEDgXiVw/60ihTPM1ZnZu/EkhyYOn1MrRQKUdjUWM28R
snBaEOhC5QFUjP3MsKvkkOt/5ST9YqdqX0FJWp2ylPkmBWRsFZqZdeo1CF0H4z37
XN/B9mg9sB/xzfHMKLMYMANZf353dY/62+FClZB5faP9e/XiSd+xJwABtmzq1Cck
v4lqpBpQN4Rd4Xw6jZqFFzo6ZYuBx0cZz4KFeTeKQ7E8EmW6DthrrQ7xGoEQW1Y+
YEhBG9M6Q08tzsMFuiszKvzWDHaXt6WFCUJ/PWJVfMpVKhULIlxsfmJo2BsxI3/q
KzBeGee4YMyZP9v0x9qScli59PGUjl2b/Sa9LqINXKyWraIGZ/2UPQan5ipWkqul
hUY6GIJfeB36z+poFCA6hvvMpYJdZN3hOABPyrimPTzslpOZBzJ/FtVAKqaldLPx
ked1A85riqiouf/6ooIVKQ5WSPdiP/t96/D9LzZVVCAC3n2d23AbSpSxlXAr5lsw
j3KojiaUrL3vFvqqfsWMTnp+PSw5ZnHVNNrMuX0fVjF0dxF5MHUhSZ37yCVVzd9j
LCgsMt9Ck8dAiZKzqKICW7cXZjZbdluVDxAoTIWiNMYNZeLlXN5xa4Xkoxz9hvzB
fTNiVXHmde1mgARlCDVtx9xvMHA+xdewWL1OmRY40dM0rvH10rVGvuEqUb3IQmdi
mTNh62wHrqa+y/JwJFtnyDZvTUt8aCqODTXitLIj2ltcFFPEE++ns6Tf+hLaWrdR
esce62kMKhRryqlb93OQn9QQD22XbBscoDvFT0g/6tqhgln/Tj/131zqweVyWsP3
Hxs804ZVdD/pUd0b4AflpcyZW0s6Cq/KFvx1FLxZAdaqSAq7SMR0s9HMpkg+fpKf
rzA5/3uaCsJv5zK/G5XEMr1D+3M0p0Qd0a5KjcizeBNeksVPb4Ao0h7f1gD6MMwl
UodhUZ+hSH9tof/duWS09j3OwfL+aELRIRtEabpKiL2UNROpIhte3WGWXd0uaoFp
bayqjNcOTlldvP2H3YZ/MbFfi9epxvKJjGEpZLLIOKjp9U860CjlvuvO5WzNV4d9
IfUfDQtvXRjPdVFmR/xqQc5sJcaUX2OTrl89QQ9tcwYb3fK9aXINHwLv/Cfv3nKx
e39XdDt4hcl7ZWrW9u9IWeNyrelm7aFvyKEZnKrYKBP/UGxs+JYsGps6rrNYxzbf
SIEh2tMW/vjKCF2btqDEs1e6TyMiS5OraY2kzr8C23sid8I0SIIlWhu38V+axxaN
xbJJtVoTyMGNZLKtfUv0G1tujOTMvlSnXas1a1lazOcF7f5zm6jdW/UlASXjwyPm
nym3rViq+TVV8B5E9SCh/3cte9zMXm0FJPnEZnIWHuYmrelcBJYbbj5bZKwdaWsy
JgyUlLuqZW2hpX11f+rQQwGX8X3SIm8JAhLCTtWC5f42vt9IwlK9XlUuxOTKVM84
db9VqVBjg+eE3t4/EgPkFrcqaEOH/sRFhg6uGaq2F25pMqbUmTpOYF1ZXTiLSTpl
txfZzf3yhslWOT86QCkdOXBxpnn3Pun6a0ZDsVeRhSMLipKd8nE+HBhoWUV4urvJ
0+6SaEv3l0uEqOJxcRPGWfK5xhBctEMIxXQl5qCr5inNWO6DnLtE0EeLegPCa77R
QNNWbkzaHfNU/vBfVUTly24GyZSOML9Mr4T+LuX3nGS4xP8JeAnJgTQIRJdFc6nn
q2HyNrmjFND/JvznbBO3zLL9C0vH5merq4TAs0q9QnA2M4v7pLSu6Q+vASJks6PE
DN79UvnugC9gCqvjkBvw5c5rv5hm+IharIY6GUCajrJvjVB62Pqg/A+xU0lxgaKR
0pNFIHQfu+yLEnFeaFpeq5bMOHGverGJeiNN5/mDsC1oymuNJKBLxGgTbtP7MmUx
TFnpAJ1sNgvlFJqCvgsKkTAr+so++Ye34YXRTCle663t60hPsTRUutmE1RzcPlfo
EitYHk6ccyr/5qxcQuuzcF5Piq5U5phUkKboAeanJ9wDry/gLJNsh2zYA9zpKUgt
wRimdK9bHT2Pcr5h2X5UcqseJtx+BJWerfKi12SjhA/jTln0KeiPSQ8UWBZj2xEL
5IcO94omX46LxxdDEHrxvDJjJFSPKFKmsDfM99ayEsoGa6k1hP/IReNBGfZ8YwUS
sMnTalsgW416/ibk9oUL1Oa9QqRXa1hCbRIa6u0uKditW9gy9A94I/03aELCzq7a
CqoBWY5rer3g31QvjaUTW3mTFJroZvpNL8sK0sB59o7pqc7YrSoV2/vj5wqJ1/dh
g6CNNJMwyJQbjP+hUbUIfNeo5S1/jJ/wKIMuYe0F92Y8P4CMSk9KGKCB+t6I+Dsn
VU86GUWceAhsLHS8bHgWfIsarLxfOOFc7iaGjuwk6WTqgQk5jF0zCTOLfhPKafVa
ptPdilNZsbm3IETNmufqURNyPrH3QTvOuarp1SFJxuUZaswxGL1octdx9RwhUDSI
l5BvWYX0ovYLi7EEq2XcjtChZJJHr/eioM0EVhKXzr+VI1dkRUb9Bz97uJJhHhuO
GAn5kGiAVW2W5pYfX9Pu7nuha6BWce4sCPH5m7Lc5+OCQCiA6VKBeG/Pim188dDO
8mK19vdKrKmSBW5WIjhkgETnLwt/R4dgMbFYCPE9VE6Bx16ID3KJin0YLFDkby+Q
qZwxRAJ6Ci6Yc8Cssl+DWsjUx67HA0DEq4y2NjzgN0y8j7snSSktUQNK/Kqx19Sl
qPlJrWUz1CFBY+91PEI3Y/Y4s/m72wztFcq36OWYztJNZSnXonI7cIYFrz3CEkcH
9vmxLjpSLyIyBNCY2a1hLfc4skgTycx/VIZ2jR+66SWn4iYzX8jrU2m63LO5BGx3
tvDieymN7rbYC3WUiqJqLq1ChAj0MF/XCNVlcs+GxKIt0sWCeQoG6xmFh2pUpEKf
hL0xwhAbZr0JmJM4q9KGnV53v7sXpFuKvmYEpw3nhGZYP1p9IC1tA2v3ryivAH3Z
UTXNOpdnlu9BulpI23lmAl2Jbr4HaraAuThssbPWgWAy8yDWWzQlrPtvyfYzZW1x
9sl2Nt057IWqGN1mEkIZy2YDnZfPjMU25NqyYi+B+2W1ubb1KQ3UCJV7H1tQozMg
+oJEva1Jte/QxYlPbp54ERECyp76cCXJfFjxRqQL4c1VV3pftCwtZud4ABB4UEdN
u7zxVTf+ws8oegbz8JoWY00zKbxXFTG+mwDsicWP/YQZ+krWwRFnfQh3WaFT0jwv
hoVx0dbjK3rgNwhqsGNnYGDcLDUfhbSjzrYZkNEZe9PTGU6Dvi6m1J7muNsvAZqH
bG+PnG4Vu5poJl6nyiVMGVBhgYAWyNjSQpCIvE/jZxQcxfPbemoABV/fkM3g3eBf
4HDn12ubLA3rt80JwLZIjc6FMeWTmAirOhcdiDP1khcB+9Qi0OT4lvDT+Xv6L01N
9P+7eymu0cIwv3EAhoK6jJXOplJShZxYZ9ElhbJAeFgvMrnADAn6VBS6/dry8CMJ
GK/Ueidumky9x0fbXN7HkDvBaCznpNt0tplzVBjfN0xPZO0B2SGLkWQP7O50wdft
7vYrgG6y5kCu6NdPcRIPUz0+++w20S7976VHGLso0LHWq7yJeM71KI0j7kRnlHTJ
VEsNB8SBtG/yrbHnFdHXs/kmGmFlSssVXMHJbNIs/Wl7TjBlLU5Sq2T3zSf4V6HM
E9r76RfH9VovbZ6iU5ZowDeVxnYTPHW2SYrkG3ZVQolG23EjmPS11S6bL5+1GLms
UXZ9jr+R0mDM3M1n8QCHTUltt711p/fOD4Ttq1bBXl8xgFHh0sVeYzFovNTh5K2w
Np0eL7Z6KnSX4HzHijQkej8sn6AL8x9sNLOAK2Squ+f/pcguKHwKGv3dA0jMPxIi
5mJ+A+Zug7f7TFVswcG8ZR1AurCexQP5C/UOlgIqcHEu8jcd8pkYzZjPGjG7oKJu
DqONwvrtoHCTo/0ZUWRcopgrrfPQ/SxlzUyNfjlg87OdOFFv/AcRvXki3TLFpWtI
AgrcjjYBTIRVXL/mG9+xn7FO0EyPSVwbjgyNo2LYRD9414QT/8DLfqjZyFX6Fl/L
AsQFAE1IClBNfCt8tMG9b6hqUbIAJ0HPpBbrELUUwB2dikVb3qi8ZYpziow8+p9V
jpb026KYYdhLihXF4G6czsXiUavwAjN2rbTuI3DAKyUZm27lESecfziZDeaASCtU
pVOFIjmK044YFx5oUUb0ojUkaQxaJHl6JlJXBUmhGsZhMe5/WpGj/Ascf0wcNZXh
B9YSH+0xzyASoGY6qXvOn2utAFIfh/roJZuxjne2u8HKQJpBlYhZYlysdwsq32Ay
qLv82Ig0jGJ3q86P1eDmwiX5N40XuKs/MPJHl7xo30Giz6C4Os+qXScy/tHiFie7
VAkXPWh6zoh3RVgzoatmtsEj3wboqlOUo2w6bA+TsNZKWGbXzMtYYKBrEUbtv4yG
mLzSVXjDiweTaKvnAuPFfFMRjuhHi1+hrj5+M+bLYHB73dBLrJmtUlgpTjIbr0dk
RysERz1IJUsUk/ATqH7OqDZICGaaXQC7ajLUu8293eYcQnYh+5Iaf61C92F0THv2
vxigRK36aNY54QKVRLYOWUeC5jFoOMKh4OTDOyTTL5hptEdV2Xl/MZSqX+/J+4j9
J6M9I1NfDX57GMkxGHYx/4ordp73I8Vl35HWExImeeN3TwT3xaSd6SXS1JAXYixM
Gz8Y5/3OG6eaIsTfDgFyFt1X+e/HzVEa0fo4Qx/o5GCtoeSJDVUjX9r/pIoOig+5
QVtBNyQ7KgMYCa51By9dwYeQdTcx34Ni1iSi7QcYyXr7utONDJPLDmeDqoeg7zzy
t0CwpUgLCkQCBaDDInWdYgtgr8eOisQYwvnm62q5IMhA7Ipw+ttJn/VXJhhvcIEd
fsSQfyUbkV7AMhv36MB6BpmQC0ZtzEAUyurrhbIAIMNdCtm9njyNrBw9zLGqB71j
nag2t4qTEJaQNSLYMjf27cpbGd8hCKq72Fw/O8iD5ZU30DJk+rLuDruxky1y90XT
9sElSGzTi/IGTJajl5yI1AgUI9nxeMPTOqnSCm5nmnZJfGtZvwb2KFEfdY2pMvX5
swdincfwFbB0u3OVLX/XCxjlEY/lYFkknUrsUqvZJIO/mh6OeFLThdmkEMO1s/b4
RiKzmpybjm8Uaw+s3G68t9/xdWTe4rY8f1SiICowNwAUOgYsgFzczklI47Kc2lW9
qGTBDkOFfKvS9OZC1uDWHOseTh5SpgXKxBcltUxguCul0A2tqqHdF2AbQKP1zSqa
1033vCaSxPy1nKEJBSbYX8gwpXfsjY3wrkmma6bPDEG4YwNys7ALxlL+lKrE1PRQ
pEJHn/yBgKQUyWCPPdIVYjSXsFMJPYVS4rrfDAoex8e4WceE1adp129lYH4/ar42
kuq4Vy0kDDFEWv5hfvGTJ2Z+931hModJVP5Wd4lWwdweFp/JU3JNm77y7eYHds7H
irPFYmaWrrq3WT1T42xZ6qoLILjKN/7V4/gr7M2aO2AIDx4WwjepJKSPhDENPCpb
etWGwc9fEST170NFXRpTwuvID3KEgJzntQqUzfnqht9vBB6YuryNWaACWSGO7Q/X
bjvj4oo2/Zvwzjlfvo0R71KP06aEM/vzgo64PESChX4sVJk8XGulz7UscFLOIEfJ
6hOevlmYQQuDDzzTTONzZyc4iONjMlJLSYuWmls71GX1v5n5FpIfY9c9cnP9XANA
ZpylyCRtjZjJfYB7hYCyEKfABfyvK8sluP+P3u8iZekxtDYGCRiljlmmwNtHvi5L
EcYrTDj3KmiNECN++NEY0B1JLluKA+zQC5iVdIuXF9Fo3VurLaCux40y7XVTK5zo
6KOz3dutRTkqHiIQdMuFVAMVjkhIX1O5oquO4ObLp3qy/qSnyqcKFDeQd6tZpjKo
hzMg+ilh8Wsa1rN5tcUryBYRGJSoVmaYMGn2LUmBgtzypB4moqt9FTSGCInjyz7s
/8rL4mO7sFWL+9xnzmAdbvDerwxrQOz66ErVgMFcHRscrLTRh75sPm5fVCTs9i/f
UVEfS+FJjEM6x7vB4hLOprzVGr2K+BgpaZhSZFzIm3ZpTWgofqE4ykYKZWSz+Z76
looZtXsDnM7n0XSf3SU5SvavqE2NT4WL2NfLMQRSe4VbKb4xGTWSsmB18rANBTZq
MfM/DeUQhJYu76u3iPaTCG9dvUnQMWeNwzPph3+CmIfCvP0LdvMU3NlftqzYTF9c
hl8ePiPOSHMLVhCEtZF6dmtajLH51YEisvf2sYTAovBMQ0neYwYYjmW+3ehEl6Ab
vwB9X2m7exJx+RT0iI1e6oK1/1WJbhFP6J5WH595zeWKWLHWWDWP5/j7Woubo8nK
YPqAMBEJVj/u9J69tHE0dlDSpOQHosYEREnVgjbYrdXZwNZ6Qm1To8iCDief3LWH
z78PDWw1f7qQWzEi2GAjE+BLSGlUcEiPY1ZpTh3G7r4IVA2zKWf1Sn8189V6KuPA
2IkDSpeZXsTy0CtkVnn5kvMAy1Myg/jtkjvcfq4ljcRejwYbfZk8aISni9TgeeZz
GstuoVt+3eygvtZC0larpH4pkdh9Y2QHyjYrAm/ITK0Eg1rRNH+gILClzQZsiRDY
h9/4034L9jRcIywpUQhgrM/xALAdm3EXWe6g8gn9cApk3VvMAduBiosY0CPSB0rg
W4lvvbGi6Mkgw61EBTap2BL/1baIhPd1Q2i318NXuQYQM252bBQUldDdPq/WZEvR
aNteBDzg9vSKC5bvhrVSFHyz46b40vJByPq9cCYz0zmoZfZY9xYWI07Y2Frh1Hua
kflSxKs+NSgn1ZOjym25aB/lT6IhxY4Fp239pcszKCaiFoYbomWF+ahDfVpWcav/
QQd+mrIcC/+x3ZZUnSZQTVrGA8b2WEkuPJ1uMfuRGeCS3eVaPouXASI3CbaLySzP
K2MR3ndVTwHjdLAnEBzeLQEulSQxoAGamu/sfP+hSSo9IIwxkeVRkL/49pgsAbXc
a9Hz30jBLfVgJMJul3+UZgqdPBWD4Q+emVOAd4Z+ZyVciu3gqzUyJASb7qAafEfL
yMpZbJcq7ZnaBMrfr4iKBfOTo22Lby4+lskT19bSPH2KLhz+Jq4NBEN61kDEWuHK
hz5G8QmHR3tSA4SVBIfPGct8VmmRGllDVwzQ+cQrYG95cu1fV1hvJJEzwYhx19A8
Lgbu7d0z5q7noEFwkyx0KZd95mXMyvpxwrRzbuUmMeS26qGQNsSynsSEHPOSXGMM
zt8brVZbsDWjl9dPHwlRjyPeWqhjGVwVFjiaHqCyrqyqveZKaQHCII37/zqa17Jl
7ny9IHWPfenVZZP/UWe7sToPSCFrt/0dONgSasn+mj0PEmEVUfdSjVLTxeqEpr87
UZYxNznlpATxwPsvQtYHDHo1by1H5re+flo9rbfd3jxFHW4/z0bUvOK7jCabCsly
XAvaUWWbWyM5N6G0ptCbfv5+5PhYxZCmv9Ip3avzdXsF/KuNbtET76/Jv6OoCPUN
SwGfsChT31WyhNuS8HQu/ByCL+tLCfOeCLqXgIUC5jnMUi1SINvrPRKOXPawzsKI
df7VsYPIY30IjB6ne6gVhM41uGIfTKLQ19l4SOqz1X0thGIH6F3OcOFg7o17zVrq
628Kj9ptOuUDdg50u+HjKe327VOxjoC/7ei85G7gtdDAFahdlwq5bJAtxgpkQBVB
VMATmS2SYsyPw7LQzNYOu4lWLPtqTNcC+svoOAazqzbfNGPgYqrM9W0E3qybUvk3
xo4h6TVOPu+/bdggnz3ycz6bsbJtzWBMTNc8DcIKpCKkR2DQnUp/ooFxhA+V3o0Q
/KV0xWJYCvwjdQ4k5wtffBY0VzW6oiqvIba5LZEs1RafXOHjYXrzTobteQY0rP13
/WMG5ftgRF2Oy1H0QfXNQB+NZqowq1WrZXKfvrHRd5v1RzYnGBTLlkzNmCYiYYUx
m9eMGSIs73JfexRBwRq04TlPJQ3M0aBWhefyyQj7m1Jdf/ucULJEr6N1m/UPYQ18
QgtfaE7ig9WqC8fF3lJvQxiXqpY3L2ArEB99sFEu1UjdAwUi8HqjALBDDdWTtoPj
zeFeDbYuat0heKQblc4wWzlrjfWTu+IJ5YVu/BcH1Ax8Ak0+uoPhOGwYgmk3kGFC
XZCdBUIHFvjvDHumDhX6cPGHtqm8XZ3175vw+E6SkifpN3au0FTW9PPcFaPrHUVF
n0VIRB19rpn6TQeUMcf6TBxVeR2jrzRpXCnrwzlQuG4C7pzFdN1CdD2PomCX15qI
itnVKtRZJqRgO0pYQyeW6tdwXbzkfz7wnaytyCKysTYUKyV1hVOoxqGlXGGKXhp1
ZEViXEaW3Y0qxteJ4ZgzvK2APEKnTTW3WPNLbQg6SpKd6mLhpU6BgyL5Ah/owUsy
vPvY4E2ntdlT1rgWG/YxiUEZcBuTjA6AxDSpJD6oDDW71a7d9kXxJcXXlKMO/Ofm
xfiDgfTDMi2DRIdxM/RxRIIFj8l4x+sebJ1zwg8jhXScsHTFPrvnnYd6dLo/udxj
z7ypCtXPWIqql5FjnggSMnkJa0DWW917LtQp18LVXQnqNIxuH0whmNTRhOLgegcr
IpLmNSni70SDsIQLSxQcmgpuUANU0dXeDXeSDASXe6RLoeaTsCnHwEbb1PBy1xJI
OtbCBoWCkOakxQ1em6Fi7uYiF0yXK2M/Ji49nWodJRmAJaXqIBP/0IU1H2lM9n3H
jUCFV4dyyoGxIdDVcbNUwcS8niqoFdrJ22qV5DEqCifux+nkhlINXX7PFkA0IjJb
Sn8AB1MMIJTTEXpCfVuRy/AeOqu9bFV6ZYyp2mLQcgFNmZzPN9qnQ2bclb+pZFUg
TriOr9fnLit/4AQiLF7anLWXJlDwVOBHWBCOzx29q2tZDeX36zxfnKMEruCv6Shb
U61KU/uMoEeOb+onGBDe+5+Dt52fRzdimnR17D/hYyHvR77+Bbn29+wzHO8WrJfd
u/WAUOrFlhqbRCaYlJSaD/ViRNpZAa639tyvLiJ/IloV+DcaS1LRtJ2EkEMCMnq5
6mADgnsnaHfraKgCFP29KutKZhghHwRYiDmw3oJZ0A3G4G6Hf7fOShH5VIYn+fBN
FPdipWcqiiRgDUXh8gxyrZlkHCcnrgX62BBrAhqeoOWLh8RJI5tn9WOfkeJsxrmi
3JvKhy6Z95lXlaapQA2CrrRD43ulrGMkqTlc5sHK/H5Z7K+wouvhEb1wR87MYu/z
d3DXiHZHo5GkGrOxpa6xa96BAydqtT1hyeYNt0tkJS/uDYWnVcvO1Z6oB2zUioxU
fSyTqH8jJLd/hjYT80FqHLMlclYogiQefJRTFMziOuML3eol5eU5XpMmT7QbOe1S
unbMfheBDZbwN2KwB8a90jRWRZ1mEK9e7qTEvVdsv8eHmVFWHG9l5lBbI3JXoR/R
nCTHf+f/Pmod+oHdrs465IwdSbzXPL2tkARalhgQ/ePSNcxt4Fmrkw+SipP2x4uI
a2b2mej0bQv/oDepVfZGAKotqO8epG/JxJFj1bAG0A0x2Hp4APiaaQLXBK2Au46H
Qz95HHo2LMzpJ7oXUJrhYfmznZXFWITFEuR5Wg9+oaEwcc6sbuzpLWHxpGQFwX/2
Jhf6ldJJi79192ckd5u352bMYjtkVV6eIYk2G5DAOFhB5MO66eV0/mw3NSEuRuFV
TehtJcQDRGbwRB7FaLnm+8UhXgwQVjDpqlYUPoQsDvcSMatlBdmA0ws4mOE79Cyg
aX1JmOGTEyN+gg3M/WZoPn4csbysV2eed2NvwSqoVEY+7xVbLKU3dN9HPGruIJB9
8ZkhN+jkzGmWktf5KjkIJJdBd51D82Q0q7ujlPBP/+9wlAdMhMKX8Ieq5oNhXHO+
dbPT+ReX0pU8+wKjRqs99SMJHNH5KOQR2NutZP2w/sntPCXnYy0x8AR5ZKRIciSj
gVTHE/qzFmVvYrnb4sD4ShA9FYDNwa5UmVHNsijpBQhL4g65fvIK3TePMrwLKC+R
f44/BLACdamfa1ghMcfxyA5wba4KFMvZsZ1AGFsJIZOQFcGRAXUsfBppFbD9MPSn
jLghP1/5R/2Ne5f9/mzoXVW6f8IrvzmUy3kjocy9nVHUPb8vdJw4bwB0XQABvnsz
HKPoOJDDF5CQdiW8c4Tw2lfD02d2LZOE4WHzsT9O+OLsJ4gAyVjVE+N7t34Ekjd3
7muq+mX7TqDRPy8znHqGJF0VoKoAVAKlA6YFoMtkgyqpbldbLiLWAaVPbdJnKCLd
8kzKNEua+x1aKkJTMyT4WdxvXPUXZWU+a36uFtn2aXHa8XqVS9VLCYBFLdWibfW8
gYjMf/tEmu36tm4XfMHIl/8FQtSb7uA3yL6gWwBZl/qb8gD0FJwG0sWy1U7/P3vD
6NozqU0l8XqOQosFob3jeSyXip9mJqnaYN4Qpvkbl4Lr0NIgLI8UNyQ1h6+JCivL
2OPU3xQ6xeqd8FKI4q1eBelPY4C/Fadx8ThAAUXfKqbdc+wazvlV3E3if+d/tJMA
rC5HBNvW96HHOV496CQEXlFShFFPigmG0uG6986piZAs72OWT0YfG5DiA9Py3D9o
LpuxccxUIC5ljT9b1IXGP/PQ9BjNRyHhXv1jNK+Tb82NwaraGBIQqN7MqNcvHIKJ
J2+JFuejO30wbnBeo928zjhKln7zKP80HcVdogyRi7RfJy7lGaGX1ODtSq4aZT6x
NdlKQblKidyortE9NHw5HHzJ/+0ko1JNWspg+BoNg1u1dvEwwmDPAz8nPPX9UGsc
/lUNJw/Z32Nyyu2GoVsKqcWrhq/t/19AcI5QeKqZ3f8EJQh4Nf9NywKR9imEDfCn
tSjzbsVvUNCcwB7ruI+t78gmqbpJZ/Zn9FfgE7aYIJv1kPSxpuUreMxbeKen6xj9
z3LVFN7sgJD7Wei2dOdZxheAXahC4Whp8xUpKCJHgIV4SPBtR3D4D3LD09Txnt9A
CfEG5WLfwbf8cd7l74SU+8T3GDavJyPQRm5RTV5wn6oDOP79QIO7tI7P2LFa+PDY
gG0NLzFZqIlvWNXJ2q9tu5lJv7ZEXgVyV+QAq713N1f3g08eglQuWtpGY4uUf9D9
39YzWsTElQ9D17RNnk0NvaFEvcHKqTBUepxth0YTGIBGFNaceRc+gNveTRZ3af4M
rLr757ekEL1eJwUpYqVn2PiH1YB31QOh3+rKqvHngn/a3slt8quiuHJZwBQ2cPKz
YmXJmzFMZ+C2NJRF9S1HoWndspMIly2VJ7H/fnXGiorUArsu44WJqsvkx9EWExji
+kLxMwjZN8tq9QTRvbJuWSzkP27OZ0KLL+9C73WpYjo3Cx65WjW87o4g0RxFCjO8
D5TisY8G7ZZSgXprgDKsbvtHGKS3LJOuFiAdgVjWJu3GFFVaVuWrmn9zzno0fGFt
1ZDVjwyklOd0Yg0eFdq89JoAhpAIwyB+yoyqhNbA0W/obZNAnK0CrpH/kFbR34as
NrCoqJPnTonConVZiGgUt5xgroxHtA1qp9mESosJaRBrMpBokboBhR5J7UG/4D0N
Lza5ji2yBzQwqZ/j1qZ14IJZDu5xsS0AUsCUMNZFee8Zb6eq+Jo4ZpADmZRA/ncw
A31zUQ62ic5HQy/381b2a2gT023ZuBr2MPktyP/eP20vssb8ioSfPLrroJ0dwxgE
ymJJxQZgJOgYW3b/QhdX9KK9/y7xGurxnOatxIYG1cxTG2+pj22jslvmLzedNSWV
q+eilb9kXbpNkXZY2vf7ZjKAeg2iqNgCN8XEHMvVxgtGgWlJ/6CGRtEsMM+cMV0R
RIAYPsCmb9NLsfiYKiiSBYEy9OWINXxmPOPQ/MhiUk99S4Bk43sVj3gdc7Jwh1WX
aO+0pbyjfzEddg5XNg/SCKnCS7RMfUpzlNrlYK4Sok6AniDbtlhBnQDTmgGFZFTU
c5mXKIZmTzrJwlO5FzgHyj7350YnB5/HaD8+7R56e5RiLik5RP+tB+XTpf3utY2G
jJnRzOQjuQeqXIBOnoVYZdfejmp70PkfJXB1aPDczNCjbbqtvUz0kO3CCO9ANrhf
Zyudf1vexLHG9oOap0mrcJ0B/LKIu/a1N3iIpWNnfbrcRSuUDYqptRDbEMT5f+rZ
xNqmlP3LvBktNJoiVlH9lzl3e6GO1gdbXWqIkELOF1qnG/2kwWz95qPfw8ROkx/7
w49Hmwwm71253Rv8B19pPHp+ZUmS0e5irEYRKFEswN7/gNLT/3PSY1r0V0oOtaxq
8Hyi5X/V6pKMoOc8c3DLk/Sma6Umv+/5NVFFKrrcoEPcF+1Eya9mufskDOEERkLC
2OsbDpd62Tsb8gVmiCH1thcQ0cKYMcOzsB77HbEzwKIx7RZneVzg/9AM9NUe9NM6
V8Zl7U/hqmTIM3HHOJlV6PV48FyjundpjlTwTMAJaBQgVCu0WvCmRyIxra93dRDL
QyXOyl/LejoxTD4d+E9mYfk1Vwg1f8VHVOAOQZsmvW401Zm5/Af3Q4yLM405Dl7S
2QNJKLJ7QNNs7hiZfNFujbk4bvWKkNoIoQL9yG2cm+YX0seHMVr6gwqed5ZmbSS7
1NZarQcsxy++JLlHXyrpbYsGeGwPCkt00UWsafVFi1sxWlUhax/i/kFpPjN9G6rx
2IWEUR4CgQrL8sLtQQgdSuLfakbv8fk3fnAlePUL4375IqzVY11Q9PE2Xdxjhtsg
7+X9BUFAo+swCH7djWV7S2aywWUxXE8VgYkLThW22RrheNFjLWtvSG+54I92yC+V
1ZQpJDTrJ11x9Dx5eE0DlwEc+nl1MbZFk3K+04dyteLID2AIm0L0F8ZyQjSccplY
f+XumvbWumpf75kdFZmjX4y0YXyvy3VcednFkavZ1XLYyW4PKYqLmvRuO3ehG6db
ruwNeyXpZx4dn8K0XanRTCS9bGazekZce5cDtPs/IVMbIMwDIFN8fmDbk/+I6pet
QmlqeImSJL2ahmRf0ccTA5qqKjuV1x+GM3xMk3IX7Fs18NAC2B3D/gGvDgJguvJc
csMRHAEzTdK01nITYRidlzp1Ztcib7dAaycXXC4/5fOAOcHzszee9cXgARN4pT1X
D+OmVhwsdMFYcRoYE+cC5LqI/5rjDVaHArAqjY66KEOMQAnfCrgTCPnzCamnt28q
8cH/nWD/E8sp45RqDj/AmiaXTbQg9dR9KKrZa0Xox6Q2/tCAUmCvT4voOJJBsE11
WyHW+mRq7itjMzcVcU6uMlTySMQzLn7zImR9j75TmkJTwUI47oA2SyXd3lxW4Af8
2ivNWQQdyB8jpLVn3rgQJ0UCfvdVxWkdSGXokDIaVfm4gXMuNOvA0DRFwg0prvgg
0iG+SXMWRuZ1VXBNbjcPf9EOTpig9YKVhgwejaUyH4jT7cQTA2lK5jLaN4WmInxw
y22FsJKmnvPK2cpChfCLCvYALATG/L8CRokstHZqtuTG2fIYz55Rkdw1ukMBvCJw
QHmCZOFApUDvkHoawSgIZda0QgPTDwkR20lRIc1fu92hcOmDXOhgRI0etJXSMu0E
lOAXmBPw3Wte/vN8aSqOl9gqdk6MRX5uDAmvK0q92NfVGMZ1a3JBuT9QphqERfVl
1T7lxCJKJbEYrQzSRkEBQGJxZIqUhUxQ9Hl8T8aa2wxAxOMlmOSkr+O6JJn+iT1z
Skgh3FEJLa8GBRV/io5Rwu6JURLqxhTPPb2aU96t3gvBsJuEpiUvO8CYkX5iK1IX
rXrZ9YncCT/hI6HnLBjHxlig0251A57qPUrQttwG89owjHSjo38itaVH3OsSKcfE
ivycJd+RRbjhZMDVVNC2ZWOFOHBpNva3umyZG+JDhHsEx6ici/Lm6bf9FgB2z1g9
D1b3zqOgRcI8+xb3y9fOVLeTY4MUKNgiR7x56cD72VM1IYAzp8XgWohtHD+9qjUV
sx0wxbya7HrLGH+L0E2OMIERYfZLf5DOz8AQXUQ+w999VxyNYfvBftKx+1L/VV4D
OsI8auPBVO543LNaS2DQw77dNxcV8XKKencEOfS8wGVJT/SSI3bxa/iRLzfebKsK
IcrR+FeKlRZfXqrjgEDShSKkbiKNheH+2jBAxAb4iIdCdR4oP2A0qMW7xFSjSHz1
l/RBLhBAwvQnN5Gp5U2eqQCwR2wIiL5AJuIn2Hv0NgXxUqw4WeWOW2bTNMfjUFfM
cg3mvsJTs5G+OC0voY/lGcGRlSsqoh+SjPfNcGUUpd+53tFQiaKsVmGrLmHSuN/j
K+MX3lNY4mphdl6S1TEEBmEnV715j0UPCeoCC0Br/VIzbx2vSfnbcINGDl+07ChQ
6GwFlsOPmQmjipuRQS7P17vTA7m05Rpn81dYnTZDdJdbKls0uZ8xNUmO7xRHZi9T
LBdMWCfjbL+0Hpumy1iJkWK+vStxuuV1T9oAW5AUmji5ciqQ3/qletbBjN65V9dH
gjwq31e3bKa5V5H7IzVm1Ee9CfYsrk36vRal4DVoky0Wh7F6LKg8zOZiF8AkKGOI
u/Hl8SLUrq1k7BXpZe+H4nnBHg/dPTl4diWfrGImkXPnuJEZNFmCLU+qVRXht31c
MHEmLe4hej5i3jOqJPGuTsIg5JIvVy5wRi0Q8CUoh74yTj1nSjNe8xSaqc42+FfW
Zn2IYnS2gplK4SbmX7iRBVsBwv6XH+cL/tzmxfJjFgcym8muG66cdCdmXTPb3jZi
XbzdckyB6PUXHWJ0FHLQZj7HvHuE6scal5izNED6lmu2WroeGlUsWm9aW3aESmG/
iMqwXHZ0fhP7M32i47hN9FL/H7ybJgcynivCrYjdIJSkDCWkWeYvtJiiWhwb73B9
VbuRUn2hgFK7cWqQqAjhuAyJul6fdZbRIup342hL37wBlNEWNYpkv55dOgQyEICj
e57nrasclvrCuYre2kIA9oqCr1+w9lLw9EIWpMr+KM3GLB7MSqTFFTPk4B0CcrnC
yAor3xGZUx8/i4rTt3Npl0Y38jxvPkLu1o73T/uN/7GnJscyBnNDK7gt79CIvzxw
jiRSqb/jdR0yqY4atTsPYWWJhoXcP6UhQK/8h3zIAFIuBSUwtQ2jHKfcNMj7A2oa
ypLJMxNBhQ6NtrLIqrToo+ThO1KrTj7XrVSkam7vHk++NY1lNppuRY96CmGmBxbo
SKeU4Yvb2FLfPruhS+9/WWurdSddPjkx+FiXt285gBqI9wIzxNCvTzMJymMKZx8u
jvCpk7QLl+TBBfy9E1fuPGSuxDf6P1cU6YpKy4WuLgYGfc+99U0ipr+hh8mb02Vo
A68JlmYmvD+RR0jSbm+JVdYySFAHIhyw6UVs85xogxLTbOOba/l69LXGZ46MHQTR
lNbyS6SKHLDbSA4YHRJZf8QrkSTIMCXhLEf/24y64lqxEui3b0ky77fYl6LSPd6g
3LbnsOQKsJtbpzxjNMUF40P6/m/vpFQN01CGdrPuSHttDlu1TCj237MSeSe3792M
cdZc8P0OUstPDCnwtjHnbZZnk2yLBJNSMdrFlStNVIywLwaW5Q2Ohi7Zm83gAKXp
PHSu9VAVvZMXTcWV1Gq7hQTzD3//vPJFY9BndKvofVRk9P8sc7WpJF2NojZ5uEY0
85jqnp+k66Qar801PkKrDqYQPiDtlHwFdp/7TsNwBVtbxRC66Aw6MoL8Q5iSveeZ
SG8hHBZDqV4bQGwcBZj1TzyfU1bzzosuOwEe8L894SFlqqH2w87NOEpGNuK3hSFC
4S/6sPqLgVgISo9ACRw22x8Z7PbnGUfzeqThWjJ5HpMu7AMyzUfd+LgB4jVBGafT
YJ+L6DhVjthqY4rBTnA0FkL+d+jks4N337fzZVhG1F+00PuMqkDeK2LfLFTHZpPt
5IsLdCe5dFKOlqj/hoWnDS3s+rlcbIxCR3849baDufGj4WY+paPtI8UWRgqeFBIL
TJExrEZYxCLpAx2Qqj8m8DQFIsq+aRys6t9Aoyd0uZXkQF0/thhB7RevuMFwW69y
zQ6aT/nIcN00obVISpVA7z5QApAmiNjc8bBHAdfLUjikhc9BZ78BPtYj8gYTzFra
MpZO2LXGeRFZRh3kbDJwtNkeLBTsODOxcm8LV7kgh6Wxc1DeqaEmp43GgnXBgGQv
Iz2Cuu1geY1a0c4ZuIs1p5uWbXo3sNXa1S86Q/CCknC9wuDTApYXFq5K5UjUDV2X
fYwOL8iyiV/VO20B5ikjodQ7+oXza429yW9uNb3MyU1s6PJwnpWfWejusq3DEyi2
QpkV0BebcZQ8k3hdX/4dE5MHN7wBaAcaejRnIUFyf0ruhquzv12/06yLvgW8EKkt
zMzTcOOkXsvRGgLrkncI0hkReDg4wgH0Xqj0Xui81UN9hsDw1fM29GagAtivodFT
FKsfwWNbndBdYz83d2X2SvHdGNKHYJTlyimg9sHiUX1D7md4R70TGuaeDl7+EagQ
v96zuQIdJ+/C5XspCmnThWR4JF/SOi6Q0aleQPkntCsFDVSWn/fL6RZ4L1u+A++c
kJEZ/tkVbVpxeMr2VfTyy2O36NrUUSv0aihYUCZyblUtgqjkm6vloo3gNo83U6Ct
aKJxC9ZR0zFIC++/ExyzxotY2/E6/CwnZEZqtVwn26zOUI+thC5/puJdtEeN1dkb
JIJPFM8zqjmh9LvBlwQSSnQquW2zvu/g3CutlWouYtkDUOlxjksrP5j0LeKGAe6r
2g4bCznT/9OSMM0eY3W/s1VUdLskEPNzPbMRP6ppSRXjJv3jyX4g8KZ+9W7NQLK4
oLrDDbRAdv7sVeJKyHwBWmvArgix+rUbH6sBNcY0Xo5Klc6kWGgbpS3qcQr3++Ww
ahOUsSrffPejQ/v62JvpUDkuFsySzVBadwozk8Z+wEqhqYwbh3AvzWdfTe5U8aXf
MsZNgQxTPSR+hVRUwadHKnR1o6nleGGlgUOmfmpp/LEQcgGQSjZh7aeNSO0gweQS
heP5NmftryKhdd+JR2T4cqbSgXvE1JZsLNGK/QBqD7gggN9eijwXorkOqqpCvOw7
Ik6FzEvtDGprIkd4HKqCsWaxmdWKSGs0P5V7loVbK2gIKZOUS/kHNrUjVK+/TDpT
FSqTbZfpB/BpZnljKZ3NSalghbNZ78BVJO5UY/sV+2Ib7uE/8uKYt5w0mlhtGhMZ
46qmjJ2o3Pvn5Ljmexh5j1K6py3apS4UouugZ4B/PtorudicCiDhpj2pETaf5rPZ
lH9XxTstEnLGRlRSTWsLgheihxHNRpsklM1bomtUU0sUVeDZkhO9JdJHj5Yj8cEL
o6gqKWinl4lrNMJKkP8usRqhjBs9AbLnhJpQanc1GSyoS4RiJlVQ/mZpNIx+uUt2
Xckv7TVJxJNtRIIbyW9Jf+r1gav2+ya5jHtAxKudowc5drhokSZyTsmDcva5hJhc
Ek4iPZ7pcTmaGrc+/SvyUGjx8feSOpWgzVme88Jx74SQ71EePweeXDUa0PgGKwuS
iPdKSodsYqN4/Zz4rdhflz6BZDaFV3m4nD5DTVR0ZvfAmvna1gypCxGXT9tH0VhB
nw/fhAoYDsqOGuiYAb2AImxhKnljcbWo1xUr6ZbnG7lcCUz5ZVa02J2uVTE58j8E
JSzFLIwJ6uwaIu+tFhl2P8B7/0qf3UyH1XroZwYsu0JXkLMgVp47l7gL3sCUjbvV
LjJV0e3Ct+txf/geDt13EHFptDoYMxVliwrayyfOF8OiiOesD4BUSCrSdZ8j2vkv
9MYYAaJMzzgYboW1EsWC51OTa1WkOxAnNXllQ/wGBeESV5EqpfCt2i59KbBNWw1w
ehfoVZXY5Q+6kK1X6FhklVGez8UNuwzlyqUoHhiSTthepyHPZXsvwROfL1IHLdre
ryomOMLLL/qd9qLFtHadcd2nKq7HEy7d91gwJmQ9jRKRTNC3MbBBdcdJhdyckZJ3
pB0M3ETFZ+rK5M0LJCaWA8XzyKy3da9O38eNC1XxHZhKwJMWwkKfmGq8xGTcnsO0
TBOc4jExKaCjlzNxT+Gi4Vj/sG+30PtJFjMQJQbsURVmQK+Bvs7h2qctcOtuit+S
1IzDlHNabP1+2atCQWWbSQoTDG1JiGRJ3B0KE5uQPoVtd9OxcNEdE6fadDEQ7A69
o647rVk1lFPcc4fNAR13DNA6IL1HSS8h1+OenC/MaBPiNs//KbH3FyDDWYu3QFkn
ecFbCZgIRqHyUQ2uZbWxQLsfx3akLpu20OIx7MN5Bj5O398BWkUXJohU/em2vTIt
RKTXKCxfWPgB9eczTOL7DxW7ULm020zIo68uHJz4xUSzMs/s6lP7VPNcRxcU6NNJ
kGgqQL5TfQHd38/FvOnjou3dv0JNjbQpin5lIJ7Yup/3eCRknLYLnJf2mRRTIhbh
aQclBDbqLkqyEMhkb1aF0bBJRxW4/WDA2xWgd5E+CpmEx3gxoamgO7AS7OGs/NWI
Duy733xTfSMoPsTMqziv8SHzY1qEsYF56L/oU5lOkcp8Op7Oraqy2ea5rsxnAexr
QZAaJeImY11U6U4b4RPVb4/idA1i8Mgcg8QsuWyihzksp/MPb3EmTshsOP8KJXt1
SYxPE0zp7oH0+tpC3FR9JWccSVvtOcXv8HsXRDM9nN1ylDd6ytDnUGB2Db3Uw8uU
Xq3aXzE2fEd8fYRN6IjbLalhfhptEihVRMa05zOumn2eH6iOTJAMVw//aaHpZa1m
JTamNqIYa/CC8zA4EbNseQrB7EWOLmhAdAscAJ4hG0hk52bJ2zdpiGXnCI1GQuI5
Ye5lBL3eIB3/QhvQRJgU07eY1p3GzW2VaqCiWWeiWuvv2VrQT9idEATQuY356JcF
qcalluNsTgQATYRF4Wg04JBHDLdt47VUh+a/LOM4DnUqO0+cF/4RcjDEUsgHWhfg
XHfzuFCnY3fo/GVCgnYHYZIhYwzxAg5xvUkCSsgx28YLxTMTnV8o8q7IZLhNRwPf
bCFhbv4RROt8u7uqatMwNMT4VP4V40GKPTjKBQOncn72QlGxzHQSXdMRX2biR/yO
N8qDIoDfVWpUQgxNoI0Y8CSPKBfrhZdGESMYNjik0HPm8ERJutpoqEMkWX5dWLJ5
m1zm64VQC0SOeEnA8LpViXPiv4kTBCpjO5IYdk5pj2yD/vKEPMa4itjVjtrr+bk6
ETzV95mtSke5ucjaONj8R3rArAl1iKA5Tt2+SW9gQKm/lR68bBnnOJUrv89cxeXV
DCEN2g5RDOrL7ttuJYvlY8/Td8rEPziOrVQBz3RMckuvsHEp/3cOJdR/tab7YRyk
Lwav5ndlMgS1f+BjqoSFEPVN40dY6QcXYk346iyWSMu2w0l1pzYsPwFHfBpVfOTh
NGmfEmE+tfaMo6096vcB4L51H4B0iPjNpEzwo2W+Gm+d0CDVAiYrnp/VFZc/JWY1
iOtulTaVj3YWid/LnWcrWFcJQKN0hSg9/05ieZLvTSYFc4Pftev1IeftY1wI3/wx
XwcPbl4RiLXDNrDUk4f56Xsnap56SCgJgdlHUNZHNWVeW36IqGa+oDVT663mnbMF
66Ml03K1125MRJtYTIXe3eVcT7I+5WGiQ1JZwn2WKqPGsvtgtHBkMLM6cXsR1q00
MtOBQOqHm8GTevBM7BMncbCpyBp39hSwZe/cI6/FdyVWm+u6AgKQi247hWTDYKrC
Z5sZs3PW7RXn4mjTbe3C7bKKNn4RNdIC6AAiOkSUE8j45j4kKH7Qd4qwSzQnkTh5
vPzFkOZpyi0wXD8tKSvHnA30zif5yw9mo+kt/Ia0oDry55PS/7UCH0hD8onjlo7E
mFkT1xkp9z9MhYhFCcMFWEHNS7hyo25/Wrd0/3v1UZCVKn9IRbytySNFlU4+uld/
s9dGhCTjb9xd0plCqU3fbdZZ7vmzrJglwyjnELDcRAXbuukqdDxXsyJ6qED3Zn7E
6+cqpubvAhaY9o1IOv9CcXsuc3dMIqLg8fSws7R86iPH3Un4/CzM3XuN4e/w3LSn
O0ihF5uO4AwVAKzd/xmTNGid930NBkLTHVeDGNP+I9pSAcuvX3vVaf4tx8kMJ3pi
vEcLWfQ/H8jo3yC5dOgy9DkP6Ow5XN6zzCVQJcIzYv0iFnayvD8JlqQ1jRYbKfZT
DHjo6FBeS9clXDOi3OA+0ZvzIreaFrlQOTPDyX3AKogayz9UWwTcpRrUKy7wlI/Y
kja3SVT5SotO/yuov7+FzcKbPqexX8uwVyqPWpK4Y5xmxMbFQUqF5YSVQPmD7SW1
Ah41vO+s8OPdPk8MmCrek9RByiU4RkvAHFgzZx6c6sfDu9WKE0runqeJDe8D6Jtc
cs/G42Oje4tiT0V+ga/f8UJVf75X5Oxs36LswcOMqwdRXFnxXNj5lr4xCOXDdMLZ
UPqr4bgBwImQf7Is1UoBkB4+uYAgMDdPiXgF3e4B9qxt/8bnEUpMfKb6WqUdb0dh
jDovzVd5+IRZI1EK5/cCBaRqMTGHwoHY/u5r/M5RpBn4mzyjhVEedmiFo3vlqEYe
1kITiaTvZNMU+Ziif3naZ6gST6TTALLBLi1qkWFpug3uM5xgvnKNum236DM+mDla
zl0k3fwe5RFt8WXpkZa6hrh6nOCiQnH6VYT1k8us56X9gg26xcyg9kBLzQaNg3qR
DFrqd0KENXBjM9wPZDwHOsGz6p+QKh5bXmkq1fpyZUDTiHFdPevAURzLd8+izJuD
kh9u8PKH3EK1V1g/4nSnXyPBPQLUgI9ympl6u0sVcrV/FaVWkSAvbXKxdPF3dMHi
VyRxDQQ2ONhQh95ISyxN9PwoOPnuZd+hPe6l54zK2x290G1tU8PcBLAGSF+YkDTN
8vP0MfkWVoBYdjoJPWxOu22WCgPPEWysHzMl4p7d5LLjIpnkAh6ZFSvU0N2VpPN4
LlXZB6IvyDzEe32bS8vNSdQEMqQlKQz5oiBonGbBp4FhFfhkqNZmIt020z5WZn9d
VPoiDvoFnSyVJYyFmn/ozGe3CysFLGiNucw0emxv3r6XmkmK/fNYKlfcoU246RpG
isBzMsILsy8/fTUzI6T04UZOIywnxpJOWOkRHcmD0W5p3TAygCDznZ/4efNj+3w2
fS9CiVE67WhWrvGB/y1464Ba4Ih/v2VmWvUtRrNQNO7FIGWfe/NnW9a7vnVPSSNi
RGHSdAru5MGLnptH965ymwSJ/1FcAJ2JojsR+QdG0vWTOSCGmVFpwdjLtrbtbynt
XD6tZ29Vw5Iyak9WO+EHtrGEpn8ypbBtLkKYipUtCvmbZJQZ0k/uR1Yf7gUGvkGx
7xawr9XeEP8XoWDLOEVLPsqw4TUq6m1ancNmVTw7J/7Y/uqEnIZ7zLs9W6zOo3Lj
+zgUVm8poVTJ0ddXshsDZMzAofelhowXMabhydWsHz9TPsP9eEqGhLG13ivTB7cd
lp++NI5WF0gUbx2r1o/6nqzo2oy3m3HjzzgdNcvd5PhKpx40ESMZvh6xc/E2JKOb
apKFUvEc87QT+mYDA15GtNnoXz91erHYFwmzvo7TvBHXsmWiVCZy1F8KemjjG5BR
8dTFURMjILWtopG7DivBes+rppAAljh2UX0cIOW1AUXv/5prYXneB17/7kVjAbN7
Fq/ocxReF9mV4MX8x+0xZ6S4UzW7OD+ft29p6NevTGYvUWHu5BpF4ceQVseLm8qc
yIjdhc43udzuSLiDsCmQB650HeQ+Dy74f8V9R3CHAfH3A05S/4TE+XiUiA0ES0Kn
7Yv2howMZs5fNTHmZHCEg3nNGCZVrQt/YOuY+G2UgMvcMu2YYogQeaWBXtJpfBFI
/WUFJWnFB7knsXG1ATX9VK8/GSNBlGRVx32ANFVLhxLGWOHujb3wBhj53/V07aPg
W7I8bm7gbQWXVDGjTo4IvFQoUuk2Mq+2Sy2EoDaR2wHPapFpuKKQ0vU7Tk1drMFo
awL1shlP4Ubk1dI+bJhKYeEC7P1hsMcxx5zQq3LCJ5tOfbS7WdECRzMtiAHzLbm5
mdE5PDrKIhU7hsPtNGoOwP+PCMgf0hbkxQK/eUhntZgTRVlqlob9E9vYsLsw9Qhw
QcEKMy6XRZ86BX4MQ7Ipy3Ke48Pudg/1/UYHlfEd1VLGIyxBHBtpZWOwZrh0/wSj
gMK7ruhM5XOSLoURs974kCNYRket11kOxKWymb9eEBe00LhBoV4HV5Bt5xv4/iNR
q1OE7S5BqquVGGB/1OhYXCnC6/JS95gaAXJgO7EG9ni4NkoDSNnFEY0EwAnh+VRe
QqIUvFizkluab4ifIdTj930jUbXlf0qZy/udiUUXM6KWzqp5L9LBpW8lQTBV5e3Q
P64RGpxHoJxDfw4CbaZVqKcjqqU/fZN9dbwIrybDTe6AXZTR4slYl+WMIhn1l+3z
XibZ5IATpDC7fYV9itpY7F5jj3hLJyyu+3J1Slkm/1H5X1bVvuYaIJq4YQ5fZcqb
7CXD177ywG+mwzsjXFOfNg+kGGUAvLXWqfA68F5wh0ZR3JNT/Wlrc65WZdczJha6
DnesjGd0DvtOqdzsaTAlTpyMG01G8u/pU1/aVQkIc5E2m+AIOjrlnIdDnxiI9GeC
j5F8bFsyMVPKeLnWtoy/bWTwlIwI1PdEKnzPgjOQbCULnUI/UFGtqSho0D0eyln3
6tm0dE9bWceZn/PEDo/ptRJ/r/AgpkM2Nxunsfgwo4L/bKBd+DM/UHmS1kOPRiDL
HbDUQBw+sLYoyQcCpuiErs/XJ6NY7lNsF7h8VkG1molyU1YALC7D5gmE3P/tcexS
K6hibd6xDt5z9d5yBedZORcHkv2d+nnEfkNOBF4IOwREICRwbki5GVqJ2JjFgCLG
oZ4fh0bY7zwdT+ra6Rnh5k5Kgo+LSETa7OGVa8mMm0IbfZbD9UIel1sYtIGpbq/7
WPEg9bx24qywsS5fTIOTnmEsVeIiDl9gGReIEnzxFFfmG4oNKmK/RrruhV8ZTquf
TBkMbGB66bGYpdDGsuy1KPqYSIZAWuYZ6ULlf8V1jrbXdOI4WFxEsFYIItVHbqTk
/5P3DcSfoUR1LkH4ctw0O21OC3K3SEPOJS8DatQrizb6UZ7HLwFCWfPHny1vQQkh
qmVsHW1uQKbC7u2uj009buJNyZrKpuD52pn2u4nKr5430rG00Obya4rFDY1BnwlB
9F4uLRhQAzbkUclGPtpO5ueesitGikiwC6skIu2jdacT8GVxZwknULTPyKDB5j/a
yVZpWs/kCKvzlym3BsEuWA/d8JDSmf+B/Y2Ryx1NqeGf3yIgVs4937pWzHWAvumx
6n9nnHaUw9Wcnd1Sxxx/MvI4Z4uRL7cS/r5euq9mBzVppfQFS0KFHPc0ZH7AFPNi
skufQP1+9QwsjixKNW+v9VRlpufp/QPAdz0GwKMVl33jF+QpWsKi9N3pqxBHmGMb
u3JWFuX4kiV3ICfTrwnKXHadF+JmEJwLoodI+G14ZkYTYaw1w/gY2VKYqFJ+beuZ
rXI8JZ5MDjA1yIHayrc2JDKy+SBfoh5m5AJeS+xZnPiPfplRUfqPrLP+dU75DXoL
8R13odOqI6GRAhb4s/S7BNmiOjiDQuelcJ4EqnFdNNcwRGKYduF485tJw6gp2/Hx
8xw810xefZgkLjPxV7m5KG433y5oTiAvaooUFG1Efnsm48pWH5pLTXnchnrxv4Tk
/GoLJXU1L7FBKInMl/tYtTfujRNqhEl4KhC8IxE1pnuqVwcoOvrDAN/8KR8CcCvz
OMBQIdUDGDoVVZ1narhc3MD39ejJaHDPQw9S98aODJrFwzYv9TfgSGZXGFRDKY/t
O269Fzp08GquAHs1YuF4mJzSyHpgqeKOjKZG3LFnuuL2RkiE3wxCJetDq/B6Wwqo
X3zY73Y0vb+TwdCCBxF96iM0ixSthSlA/6zwru/Lv2nVQbuuMJkNj7+RZHSr1+pv
Kd3PusuRhONFhXxVE2TZ39Wu/OQb4sV+Pm9ZUXE5v7C6NG7FkWKkiTCJOtnc80O4
cgqd3m+VFh+6sIrmNUM/zaFomc/0l2Jql7FVofP7qATTURvoQZtB/NqxA2MEzJUh
Yf/wWmpNRU0od3RaZQECjmL1p2zKjihBC3Y11VkzultYdkyIpBPTmHJpc3HxFE5t
0lIJqg4u8hMEk4IqH5HZqs7FDPW9EGarH5qxRA0ozSkpDcaDrLlJ/diYl2YFrcre
dJWxplc2+GSEcnDrrEi5KonhkNkzn92Zwxazy7QqtAntb6RvwXFyJjyiSYis6H2h
Rn3dYNta7Y88xR8J5uSOvIg2e8iZEgxbKIltR6XoTRBEKOvnutR9KKlP6IuKechW
Z1FZ80wiytblv1qTBuemO2hODHquZrS/yxjWOh4oLpRrv58cvRgMKMnEaieUSziV
BSS67gjxmKiZoX8JdJgrVorRnd27KlImEQ83U+AeWnYaSRBet/QIYs2I1E7xisne
kj+l20VVrxpuGOuiFFo9hItnIphjgmejnwUYqTsBzn9Fpxbrik5JjGirlyia2Xmk
cxZ9WKwpDG9N1NMVigXPaDonYwcsjZZwfMDZ8CRymUTFHd5muZAXlUyVoFcwzZ+0
Aj3hNulvWBxScm7kwg3zttyNqa3pdGUb+xjO3CRYxMYs/CqF94RXgNNZHanVqsdz
UVgwj5A56KR0+5P3S3GY0P+vIaS7SI+Zcceve1x3CWBmEHdRCK2EZY6AxKFmagG5
nyF8s51655YJwZKj4V4vykDGDUjWwDpQPMqOSpw17uVa5d/deEtgPsKBX4xkNg0a
IK0x9JoJ8Nhs90g+xOl6Y8nGCBweLQKAz5yjXZZ7/HEcHdXmSxvIlvU5etI+cMEx
GBmVAoEhs20d1xczus1kI4A8dMyxG3S4Q4DYlbacDnwI7Fn+wQMOFg2YQFPccmXr
mJ8dw9mqo1JVBRF3gFd27tY/uGU0LAw26z2lAxE6y3I/uTdBvvsDoTixDru8pi2z
9IfiuHFoVnH9bRh9CSO2prcW+rn1Ze5FT7ROekCbGsiCBIgLZCmh6+lxdgeDHg7t
187N2i6D0I8DIj15Kj2dycpXgiFXYOZJ02SE0nGzVgYhAvE5PoB73LxUb4IJOY5S
ma1CoBIJWBMF+vK4Gl0QnzEcijq0+4TFlApu0Z2T0p4YICII59HrgaxUBrDcowHO
ifrIIduxr/vObj5uy28RUzMjZHsJCnLq/TkAKwT7xBHJQziQVv1s+VkP3CZKK1jX
d7NBu6bMZSbaPBUyZlzcUjhnkGGi/XqCjST6EB3uIvPwKpZsD2gfcCGgk5gQ4TxX
gmubENOm9akL9LQYAKywGb6gxiyXq9xAmle5RMAC3mLL+b6yHwCvM6EYnlTfsQv1
WVyH5I+1YMT3KC8DlhHHPFJjaxuwdKiIG7l+8ti44lsAsgCx/ccZAIBHnAeLOvvP
N1WehHLqDNUheQw7m90+1FN9mmzlVvVPZrr/zbXTdn5hncrG6gyQ/wKWwFy8PfxU
9jiY7V78X5kAv8U3YXkuw+d4qr9CmDwJOj0qgWbp0gBQLO8whvoQKxytNR+B+nE2
iZnuCaf8v3wM7WyrnihBlxRAMRditdemQMKAOfqN3FR5NBq3fAV3EHwgyKWMcdxc
J6czmXx3HePp4dMtNkHIYW0nVCNF/21UaNWdBYTRelpqPfhM3d/Z/LijUX8CZTL8
tSqdjvEIMx8JoXiFvglYAj0b2nlJkjSeopR1Ib+RnRO4SYiraQBdGgPM5Sl+z2J+
UqsL8pj7AEhOWa20BGakFgJ7LCvnllKkzh2Xcdh99EUNnRHEhFAomP9ukKiKdB1D
oLOQxc4C+fMXpx34YJU1vK6WoaARVdgzk18UCR4l2VRyHyk7S8WhQehg4z7RITo5
Q+uP9sJYU0deT5BJ7guYR42bwmpDLkFfnxmq31nHvd1hhhQeUsNs9O60NtCBlxK4
hCLkR/FD63c4QFw0L7HXUhkUr+lAGhhg07y+HPDqjKLoEPc4wiWzFCsQdg1QL7we
DW8+N1Y2apQXKH2E0My/H+kdL5GXAegEFuj3zBaHzXunsQZco5Lvk0AZ6Bu5mMe2
xgwGm+gj2d3345Qo4O64VET9QOR/35pL79Hij8DU/ngkCwdF84W+GHzf6oqvb4gG
Z2bssNquE8fZ/fCL6/FO8x3qIpDAQEJJPdO1CaSyBzs2DwFjCLSjI26UHTBzyElT
ehZ3yoVPoQ6c4ks4q+YGBITq8tSt8j2RNhUwwxMMX/MMrkHlqyMIyWx6J/WKMwA3
ZsDPwqTAQscT7l+ssmsHx/+DSBU/nXXpw6gw0LWzMfC0uTBZJrjVZstp8lAypTWc
GVTErzPhidMAjXkmiFGWLTzy54q72Yz7WYnrK0Ux6odXYCagoU1nM8mF5zKJ/lLW
0qogfxGk2H68iUKFF0UH/2jN9mPvgGZHJ31BlKBKrTuJX5D4tko7TOs11CBuq0hL
VTT6DwjXJkUdYL8f5F1MK68gyfE26GMj4Q2HoEAmDumKW5RODkZxzqiDrdSEG0Uv
+HE7o4lqS4h0uANDGAInA8LvCLdFGzGCeCmpYJ4z+qi9G6nu8P5YiBKPJW/bS3zd
54EO8OtTXjsqIsSB49CCcXhpoxYJTEfwefNsyDlB9snR6D2i3fbBsdnq/qgHLF/Z
PI4zAZttjsqIcsG7mZs8BOhaffUHNaN8VAjRvuhj12tDWtp9a8Svdm1r1Slz8HSM
goqi6vgFtoQasOHAb+jn841GLfIsIbwpNz0ufplBeDNnI9V0lfsRSewb3LMgFLbb
sExx9EMlTwuDlWxglf8pf3BCXwGAFduxjWvWbobhGAh5Qa9NmjIPcm+TrXy5cEV0
8AoOde0E09Y5vqMGPWMaH+xsVKl0PYUQzdlxRVq3oQJua1oLyPJ1PziWr/TT6J8c
nLSVHEhFgtoAIPL+BzMvuxxV+7WdAk25QqU9wlSdPjJCHldMTtmvFB9MUWA2SQkQ
DyCccRofs7ntD+QpzFm5mrQs9DwRRczMJmTfSqLfYM8eWhU6n5wKjjXaOhcyi1/c
fePqTEkgW2zXHURDBfHo6vvJAui9Mvcayyrp0TL234d6j/+HCVeTELMpXzm2iVG3
YdPHfITBhGGgT3dvgSSA8bV8KxBhQibAGeWgiB7SGtIDPSmwdmri0nXd2ewnLbJi
odzQ4oqyLHRLh/jKXTKdv/zBMnA0dflkUjoVL1PWBHJnqa2hR8c5UASpMYvbJbUw
DSf0nkGc6n3m7HaHCNLSfnGKmbMGLsfwpSKRa0gLAs9tChaM5QvlBS763K9YRWaZ
BboBlK+hrSOMMojWz7vBJ/6fC9py7QmOixulX/TuSairjgF+XxO+Y/DanI9cP1SP
W6jPc+hFF1qvDUaizbec2GE81RAtTCdrpbsQ2XaRQmYY8pPzm8lJQrxWUPLlRG10
FifgfsyZSZ1s4VSIbm0WAi93IKJWGkCSKJ1npZp9vuzg0IPNcqoQ57L7VZg8NBzH
Q5KqtswyW+IkH9XUHCJPLOhlZDfcI+apeH+Q9XoSbJB+eXSUEoonDokdDqMaR+Pv
pq1cTtipEJVBMTyuOB2hWusdcB4tGBsIs9V/EnZaQ8YAL8+YMgXjqaJ0tPg6rGB5
3w5AS68jRZqrFE0i2h4gbEoL0wA1QgmneI/S0TWizOpI9Z7iitD1/Ia4CDHJ/VhK
iie2erkfWwo4Qd0h8b1+TKXUBhOd1jB3wzPjwMrylSXUZUDqeZOpLSMP6+840Ex5
a22lSSA5T8H6oTVx7lXDcV/gkWbOvtHKlVXdfdr5HHE3Jo74XL4drnTOUtxjS2vF
FskSNiVYBEar276LnopnklxZjBfQH9oVjDxK3BwkqgNDgQtThTmVixxWf0UOTSOg
Ax6eIEVDDTQMpD+K9GTlid5L0ygsjMYjq4ZpMwgGbPrf146aBPbowyxDN9+WEwQQ
8eep4A3CMVuqu0B0s8lrdxgB16271qaIkaqNjXPupB1IuQr1q9psXof+rENOsVHj
oQPJGMMKhLFiwtvFjkfasnwa/zTFV/UldXKWw15ybFycc3T36Cnmrea00NJ19/wW
mmnFiO3Mj1RW7wT8zDzFnMu3O2lNplM6k0MPgvW+jSUGHhv46sghx6BXRk5i0g+1
qGJPZ3Qd4f1mxRPupPzKMincnPHDMTWzf4K8dQkoAZU7j1EdvgSe4NfP/4HQt+K9
GycD1c2DYORXTXF8HQ0ev14K259eCq9n87r3RBUajALATQVS/TfcoQec6gC+EYvx
bBYZu0d9hMbAHqqMmjni4d+b9NY41Pe52RWMmLWFO6n8Lnyesh1547di3jtN+PnA
hkcFy9mHvF/y5E9Oeompiog40GyTW6Dxo1l2tPaKI8xA7UkxEtKYL00Q6om82Lxv
H24Lb+YHSVrK4YuXI546lRjvK1PjcC2pYQb8H7ROWV9NM3VPsxTJUqTAvyk+poS0
s41qjiNwobd/HwyyTKCXH0d1UAWFpaUkhdU+87SVDfDAwkHZf2OMo19mxuBHg8Kc
PQZ8a3j/Udc845h++MFisdqiQ+ptiMtBEkQnIaOx5D85fhTg4eUdi11xWsikJyxw
SqjLtQ7Nfsgy1wFi3Coc77twsh1ktw8Mv4867n5goXGAoexNL1KSG7MnMum9l60k
SwAj3u/g+BQMyZugaII07Kn7Mszk59dMT2/l1wavrsHdryInOk2WmpJH47ecyaou
EInVKeMAUEbUw2FYaNDenfJx/8EF1XepPRN3fljSWNy81Ddxbgik0l7hd6iRhBda
z6xnxbVJjgoZkHCNn5oi5MJLD+rz4R4MHvCnvMY36Vv/P+H3wbzYMRPXvsQSlIRp
WX0DDMGKMIEV4WPjchO5njLQlIirNjjruncWjZXHGdFt3+GBpL1TxHENKW2jZS1O
8QtVFfkjWjsVJUOa9L16EPv/1yvEXJLWMIiWUgstv7GPIDjmQhMocAMTTNLhUAaw
67D5gIIer5vtFxFhsPP5hpKAPxOni/yqk/TISeoMjhHbjHZOrvHtSwR9mnQd5VLL
gdwCAKXle8qW8RkyYMcX1+Bss5KQcjPZjv+lKmQx28psKI+2oZSrcdE3dnaImrhB
Q0n5YbXwcjLpDOQhTTo7Hu6AtdI2itc45vjua3o/X98xkYbSpaV32j41+EYy42oL
nquT3f/VJbqWfr/oN3fXX44UStYhlXV5KQJAXsQOoXK4TkflYWRctXiyLpG1xJQB
AjGuPGIBzVdLnUX6rlf/J19MP/UgmlaXAEwdDXBehzIFwfGcILa4yTWjXgrKDP1X
BMmKQHc7LpV4BFv5HebPuefxyUHtMmSDwETxJqCR19ibRvfhrkyJFGEgxbimCLV+
LtwW3qXz0qLWVl2/OkRXiagjopJs+yNjuiR1jTTtUy0/d2vrMcWvFkP6AmHmNDPP
5c5+0XDnECeXjj+WUpDzrsU7nFNevp2kxzjghDcqbGyFWE/VlqJLx3eVnm5fEJ16
ZU3aFBi07XJPJmJCtegRKZz39+FKRiiWgzEzqL4IKlbg/rGonKAeB4xznzeURkca
vRC1AA8xtE5IDqbTSrvn9VlhUcu0QsryFQuY83qmXXvjjMJ5sEK6sHI5KMZzxhLe
rV6JjU12nIYKVUWPdPzLXCnF/JaTbQe7RZLxYFgAeQB9vEZ7PSLXN4QnrIILcgBo
Hsc8KxbHh0q1RSLdZyyIcGPC7iVyetXyIKcOuGccQ4/JDG2DtqchNiF069OpH+vW
KCoVlFLJTldHL3P7mqy42JVaR4djR/fzWIUwueNB7g1k1uQ7aReMLRVszFwaRYfH
Z54z5R7EX3J5q0HkZKsckCYcuw/Z5JN+yG4jh49Zqzo2bJFLxfD8+KGVRI3OUbNp
w18yzZiD665vcyGdb27EQtgnhTum5eWzc5DfaRCSBy0Bs9y1szVEgcCXaVRSSOeR
ageTzJqwIV4JU4NeqU/RdgxfSqA22rMsy/cWULluaL+Xv5DDaOTNrVsQVsgocG03
OAVJWoT8rN9Y00/o/lDCmEjJx6r+DGbFKg7AZwwCUJZsKxI3NpVxoith2Nnbt0we
5JlsQSJJPv508nMQPBfzvBfsNBN5dgqv82D3Q4NpyKPz1R8ez1dHXRk79VFGetKa
9dOUKZ+XGsCRKII49vP7UuiqjzF2xZ6yTK/7e7F0IVOg5Q8mi6WWcLbbLuyQExGc
h37F3WQVgNhgOv3/CBbsc+R2+K9fHlcZlXfRZrp65x7um4lo5OaYroGvkCaB/9JE
SZv4ZondVaRiTQmfFGtzfmWvQwgBaDXx9ju7a0x6iEmg97cR5+YRWa/Xz/74QepM
I/2dCAp0fnhbr/08OMcQ9BPBRfBO7uwE5qpO0vKi038imVnWFUdF56a+paCMJvZA
AlSYsAIpXUaU8v/wyp6v+zk50j+JPPyHsftXsrEc+XD/dLn6KCG8nRhz2POms6om
vM2zL7m/BNOgvJuXCHBBUqthNIDq77PQsb7qyzYn5LyCwBjjxc93XhNw1uej54le
MXvYEEljvST+7Ntfr1BTTElnFodqny6IoRQ/lxSot3dNudr/tALPNCcVH4RcmjT7
tqy5OuAVnt/0v3bCvRdRc2gttsFBNuT6PkqB+SvjtQnKA2794e50sEVglN3q4J1b
iRZVc7udcQTTAfX8tHMOkOwu8UYkIsoKLrtWJzoeZ9ANDGd3gm1N3O6P9biP+1gb
5P7c/lNn0Qw11XlqIRFmHYTOedMaHqxj2Rfsqo5pkog2t8GiO6jVBIpRVtomK6u5
LJYQGjnTcLQd+PbSUxveQ+rxPCQ+wKXjLKUgyRxALTAI3D8zzfc9zAtaH7KkG7/o
giZLwInFrV7ot78A7LWuIJy+3ybFAUeAbixs4boLhyqKs/Z7hkxu41rizFYixroz
Fga96YpOTR9SqAg9rfsUIA7IAH87WQ5OwkFVITpZNHCxE2Xht62snzjihvaIBw7p
F/lnsXA21diCOIVyNPF2B9L2Ew/AsfGd4Zaf+t3wjVh5+rZbWqxHSEV8GA2Vv/2t
RJB+dWAoJZbudPs930cLyd/KuPNuII9N7e0qk95rIgLT323dBwRzWdvpstce66/I
RFEecIB0UINo/6mS5b/tlnUlHCKwB5A3GzH/mo6gDssBqW5ufxa5dzTMSXy4IgoJ
Vt0zt4/2ieJBICbzZ7myL+TlOMdeU/pC44dKTfMNSAaKEqo4PvBmlrd9WtsIt8W7
ZX9mKVxaJRiNGTDd7jpfZSZmGqk22CMEyZWj6YHIaSc0vfGHi3W1HpWJ4GDFu/Ut
Wx1nOxV+hUqG8Q9OgcdFh1VPY7+3VTosOgUGuCb3oIwpmMCLhlDnY23XA6rNBREh
RuCJ4xDo67fOpPXIar7hNBNMKmDn8mpD2H9BP/2RI+2LbfYUNMFz2UVEN4FEEAwU
ONYfRjwJuEcNSz4/7II8KqJalPH9U/fLra0FoZIpErx/hacBlkkSWjGdNidx+EfC
zhmJfzeKfPWJpippH3whrL+r6Owkj33YZk/86IZ4/rC4MpzoQUrnWkh7PSJnEk//
62xFsoCN1YBhxrOBhN59wrs+njjp2JdZbxgG/8+cHhMxFKHhDLfBtkZXOnGrHcAR
aN5hhsWRb1t1O3D2dEu0cN8pcCDAsDtLpbvLVmgIbYJvrR/SL4huKvlNUds+Bro2
RUfCUF5XAUkWzPRQzkKhUCTp59EqSvtkB3vtUCvR3YlSFuEZ2qiSwiBVpUGPC/R5
IzOSzqiCCrzylfh+VBpzb9Ox/g8kOfRQIRNO0dI7AULt8igiehi44V8RKo1iP2bg
b48HA+MBHh6MAml3lbtNlVUtcYpbIEWROmwebdGgkj0X+Kf1j3c5/a++GTSKTiJj
NxGcmpR6ud6naTHhzs5Foptq+Sghl907mgvUY0YHcaEyXYzY0ki5c6KtkK/KaFvD
rDWiuaH8UztJvtrepLKgDqlCjEAh3QWkbG34WuYW6GqsyRPRmei4KFTE3YHUvzhR
jR/gGz2JwfB2k+fsfum3N7q6KAopdRD4X6pHYeEEVFFI96bMiEVgS1tpsMo1TaHB
BEsRNf0rgxyh9rAu8XuekdIJyTKmkOZzp+oIdis6DeJYsOrj7XMeCov4Wmp56At5
pqTN0/8ndSjrvTQ8elebuBBrpzhImoJG3DEJBwYR4ItWWucBQEcGBPm+eF0KAkyL
jQu6JQEtGi6ZiNfYlWco6V8a85LzeLx7J+oAS/6EZt/yUEQw0Fx3qla6Vb70G2VU
1Rl6eZdmr7yW6h7w8e2dSMrxW06FS5kN4k3UPpbqgUJEG06gshS+SAlw8PodOfUL
QKccp9u8unlyd8LdHs07y2RMzT8AVD1pNLzNyiq6zVcm2n/gcTJ7v6cfOWMa/Ifn
aOppmPlnqStpJWJO+YZIGCXtb52KRGt22K3IY+lQpmYgLxvC3igNIN8as4wMse/B
XMjAZ9csAmj6j0iecI9DiGXv5wxFSPiesvTbrnT4ylPwTgQ9k1qfvsg04LRGOMPq
CyMcTgVhpO0wlMbiWFDS1L/eC7aGVZ+Vsu8N9aparME8IN3b3cAmGDPyreJ4aB2J
MnCWth9DLdGgMfw5w9GzQyFCkG4OC55oxZUM2PAb61lMEHT6b20cCFqGX9YaWqoB
htP+eFnP9cD0AGnBvcaYunMSC5NI/76DgADUcnIXSNhTSmKlHPpZpwNBWXeTQvTf
+OZwa6s3srfLyVYq4JfU+qjGBixGYd1lIsjWH9KgYL0a7BqVgImKT18eXxCOZWaE
2eQp9K71CnrA6C4vDARyDp3DiXFoBMiq6N8xsNBlDBlS1dXqiOhhB1T6kl7Zd8jt
Njwnjd+I480g/a7b2WKB6oJW0QZh+ymglL8J3CU0NVio6nFrRFH+BCBBx6N5ta+N
TVtUK7E+PZCoAWXpHCBRo5dhuKCEIL4LUEmwwhcRd6UQMsZiHXtSuaI1KaGSfRfu
PLk4YPgafc56oQkCfYfVVkRPNsccyZ5qPIRR4ejHjSl5wK2VU8eEqYdl8c8NCAz3
qWj35xrd+cWaUqv8i2JwvxC0NT+Vwd8q9NT3+0bKvDEOgU3pjbdCZ/Xy6JPlEXlK
fTjeFE08hFQ/ygX7jIMcyFkLalhOSwLCQBo+AvJAYmbmMQHuN4rN3Q/RCwXO+pE6
rXfhFAe8yHNwMaPzy5Edc1cxAdlwSC+4hvwntBMkATNbhCA54MoK9gngi0wZcvAh
sK7E/iaEjdqsnq7kmh79ItSkKQ7o4AsUtO/gmFkCt5BV279A9g5f74ewrrrlsB3x
Fl79h0lLcGkcOXg8yJSc/71xMb3Hq4S105kz9YXY9KR5JCz43u3RxMLTOoC2f+D/
S6BKzMD3Q0u7j668S1KY2e9XYHWyOgEKlE4l7ix1BiSTHQw421nHkviCEewk/AOK
VrjLzt2eeyk8Q6NE75VEbd/4LP5Pki8yNe5w3b7Vdb8dp2hz7TpBy1y8+SwUfDgC
ffBuw0aYOAZ47dQBosO2wG/eKUlEUn0DirRzgVRRhn7RzjdHHZEgZjpMzyTXOxPq
oKXf3JH7zNADBBjg6mnSHtft+l46RwNnWrohiltB84DUfx1mCIMYApATitvJEPEq
5jU9QKATJgpK32mNgCE9CubiAeHH1c2/JaniJ06O7fwjXgRHBQVhc65xspzEs3xw
W4JFMVZL9aw9zNXhTIi8dbKZqdstIjfmCQnltc9nOIPkX0y9UwsU8OZQez5WN+og
WnfrmasKOJuveauyvlcNo4g/2heW9CvZMUo8LQvUDBzCR/uAmOaEB1pBq49pkX5T
ZjxGr1ifxHdUfkCLcTJTD11FG15OF/z5hzUm6oHhlYYbT2HXZzXx0rp8+DsPxYdN
f+z5Gv+O2xWFeeXz8UkGqn7LeXI4f45+wK/W2ATA5aCz3MJH4RUcHBiJvu9yvmcP
xKG1RZ+PURFlcT4npV2Y9MS3bjkrN51ih0iK+uZqhbDVb/0G420hroQfBbYkJ9ae
lIEphimmwBFgyG8vNGqZJNA+BkqNznKBXAVAbOQkym45JckEvLIzjmwf7tdlBzsj
jiZ4f+c8Kzbyza7+D5WPF17Gr85IKy3dMcqrCFWD3m9Oyjz986dG2cI2f0mQb+5d
LwgCzwDC2Mm4k/lNQ9J5W0yQymOnF2NYVE3bj2bIxNWX0mwJ6BaAp8B848cHirxN
ZGFyU2n4tBUPBkqLLM9oKris4huLU287a6qai1C84pVKPxCDMbnjA6rIEyYAoOx3
MQzS5zcpbsqzKG+wSQNVnU6r720fR7f17YtjpfsfIpCbAWWdyzYppfRl4uL0vrTA
g0tqQL1WtnNhcIeiaSqTUYRgr8z38smF6Wg998/2OHNvjHBt79Pjkn+qjpRVSAXN
RnxkJUS975ImJnI3WLrnghGArFEr0COr35hFsKmDt1VVS328h6dox53KlthDK7Fj
p+4VPuzXKpznCw945o6qrgqMidpApYOebKcue0tn7By3YyywOdPy4f4YvohAePo/
pgsjoiFc/AF0L564FAVhAW4y4Ujh98nNngaOHvRteuUayPjvkQbpVjsnqJpiA03A
/YxhyXAi9/R/1D9wFRTr9cl6F/OdmyNIl/NYM9lCiU0PlnCdCwUdxtpchTWPR3Ao
cNb5ZLTD9vKIQUVODAat5YXNdUPfFihm+E3Qg8XCzjYrygH0/VwPvknCWYOwJi3e
qPHle4SWBYdYWxPkPabqQ0yERxvVVpMrxXBrLeOYOGDSnp3cwZOakz2GV2PbPnzE
hIsfUYdpoZCVISbtZpVnCkzVB12i+X9926S4gLhw6l9JJvRefQ+BgZ/zKX/EC0Db
n9B5fR0kqUL5/l5/ghNABRsJz4BVTqlk5rdW9d4fqTDk5iMQXRaKcE9SYtf4JStC
r91NZH+9PqumHHSNkZCwADkcNetM2g+obeHANfeIzVaHQAL1THilt4QtEtyXbhs2
IAe4NlopdZTWkSGaGIUHVsDo2OxmhoUkD9f6RJUCWL163fFuN9R4wx0zSPcLMzFj
oybN86dkas8Gl4oMQbQ4IIocvAogepY2/29iWqfgIkLL0/udbNfLQ19UAOkSjndo
LyYU0e6S2TiBlum0rB2+iL5lUaEuS2BJxfnJO/I4nrdVf+7paA0OR1+sSSOZKmvA
08rJIAZy3ivh9xGQnAT8OVjkEBIdR+HntwQg+Eel4793HmgZyRsoAhttEC2+Ftbg
fhTOoda8wOLrEZtLnOwI73DfsiyhZ9iPIQZdjnZ8+YEzCpeLuKyhf13e3uah1dAE
r0XtYZGyLQXe3AIMbHT/TINx4NO3UvxRMCmGFXPeNBkHz1L/VuYaKMnJtcEeoamN
smXPhXpQRgnc780SJl2reoxXm8jS7Jd24mtdc6HoWi2f7EkvLcG1RDDTizYHAf0i
WIsQtx73PZn5DtFV2X0LVR6kyjwr+QmSXOqeFlsKJb4OIY7VJvW3gOjQ59nDb4o9
Hvst606C55IvKLZZ8F2oE8Fl+MXs4goskjwoi4WpWcmfHUE/EjaOxCmSG5GVENTF
mioZNnDbutctbc5382maBIqCrBInpA7iGCeLoVcTjg0nW15I2jxqaaXn20Es6fG9
C8AigJbuHkICZ8BEOC3p5pN47cYxcS1zyKo2mE5Gt3rzLWSDZrYmqDW+2W2OqUff
U6/5ODnn5wpbRY6+RJsmkmHsQQVZ00msZ6HsSx5UO++ANssDsMkal1jhrPhsO/6Q
pGuMrPq1XMx7kdDiLtY/ZXPTPS7qC8z3iF4gm+s7R42yVK7YnjIFdHBEHQZ04pTZ
aqmcj1pOfc7CEp6EMrTyQ9H30xN1/rdefUYa6hT7+xqMavd6uiOBihzcnxFQf2Vg
GBav4gJEka/Pbhria+mfSCaPzfAUcZ6HU3bNdZSk73/VgFNRZHA6aJLosmjvkoAo
o/BjTGqihGQqKFYSCjeclep5IHlTJf9O4eGgh5RFwCisSBIeh6EN3VfP5EtD7TfO
aYEVRG/a7/INWvp23wcEGjw0Sy/zkiPvAsTEoJUj2N4uCEWJ4GdFteXDrl0SXHDA
vFqQ5DWG6SnJ4g9D/AFLh55EK4Gjbq9CTE+5/oDbYK0f9TiixfS/o9GnJRuUuGDI
sfKmhRqDaIYOe4/2Ui5AxcwRNBV+PuXULPkqm0JBQrmZX2PaqDHuxbZasfvrza0g
DzuoZgOnpER5HScCmwZvoFXNMPjuW/mkyB+KXFg9ebM7iNElGdtRLGmfcHFPdUJL
aaJafSylHas8R5JuLBXi964UTLhLELkgAMc/WxRralzZfaSN4F0o+SugMlE68Yur
2EyIDfyCei+Ty+USJBw/aF5YNTZY6ycGBrh8gZk8fDa/9JJ5QcKAw7JVOIxo4jv9
FgtzdXa7Cw+U/+9rQfDnvzgjPPpRQFeD/ttcarjhU75dXcZy9j6xjK+v23SaruBX
TJfSSCCAhJxL+T/gOSVdvo9zvyKKHG0aVLPfplNPk72o0FAImzgnepZc6Lp0SwHz
DRPpkxC9SVBIpWokmGSwUd7UW8uoefRQidH8LSyFwIzdC9GuM6cjUObz9T7DQnEE
Ll1aDTAF/+noyYnJpo1IdLCCwfcstVdQCMhlRsgmIZ2o85Up1xygVW/Xia2IJ7IN
4Nfqcx+yWp9AP3DxRTB6/tmS97f9zLnQ4CG2yop91WLNVDjV8GJ9mPzEXDuZY969
tOciRvWD/vslcN6qg2PYnyY4ga72H38fsk026XbfZaHrNvoHPBTqJ+/UEQ3rpG+I
1NlSbxK/otA3dTbrQYYYSLt20wtolJ/zmpixaGyCwK85U0Zjvg3XX421WPjml2gu
dD5d7Uc3Ff5/U7XvXrY32EG+KowUBje6FwHHvsykCiQdKvXbImxRtp5fLthyor+E
CLmES/d1GdGo8mkAn97q7ua/gQ/a24fNDCyHHRQI499fm/ACIW/9tDgj1c5rin/p
CaRXguEI5fAoPHA4c4FK9382u6F8dckmaufURz5T9kAPbfbZWGDHodmcLpS07SPw
EnoSdCsloRGJan25V2Z7iCW4oupa/WVlQP2yP+eYzPyTO8K0SjEiTUDHpliq9LHX
EtF2OU6+wN5fyrj1HC63DKWAHd3HFAHfga0D0iQBnE0xVGaf4pmz1+ingQ2sdepk
k6Fd4TYqsECNb+bTyK+4UHksfJu4u7CTsxfvisv8MOZ2SNHuUvAL5txH2Van/Gvm
cW4D5aVlavWLVLVMSYlZzBvWEWTCfK2kp9E74FQlySKuOPlMHG12sz0fRRXpjvW0
/cRU45qzxQXhK7A0HDseMcBIIzxdpOAy9wCnm/6rNZWsy6OZludaj5qzy1VxxPYA
P0Q9iGg7avRiaD1L3wNVLoAIVlvqNshXPILQt2957EGqczpCtBTWMq0tP43KVAyH
QVVUYmJYCLE2UeBOAEivZtq+AYOZkyOJohIvgk+W+AY/1RnyzhMJH49EDpWmzL6t
VnKcaBoyTTPnFtPcV8UqQgiOz7NIfq/R2MoufCGubTBGtsHgb3oxG6lK2sshqH2q
B8pjgMXmXpohHWC6E5R4LMLHQ64vSLMAQs3bsR8uce0ZUgRLLGUrOCylAj952tTe
xeh5emRht0cBe0VNvMBQQWVcW1zNgfIF6Kz2iVm81vlliGRci9oduE0s8r5sngwg
6GENOlRhXfyxBcD8hTOHIvRR4JSUr0xErT4jZxKpe07rBbLFUB+u83hCK4W/Oj52
gni+QVtCWWik0Qg2ji5K3iirAAVXnjLgssbT+GCnd6SO60iMhEADkLegfxYCuGFr
5k31U9obT0KcelqMEPLwyBplwR1e3p0wONhzdIgKuGX8d8DvQgSu7mZvAw34QwbQ
Nr0U+fXL0rPQGOu0lN3qpwFTWtk2m8GPaPh9Fmi2fHHnM3YlCYLLEekPsj0n+xyS
p41ZhaE/3xJfwd4zhdwWYFiqELDuefxf1YN1k1VMCl79Nb3IOBs6Rr37vdeLJxpX
6D0U0D6yNHkEThaV6yGDB8RLrm6jbYH99hhJ7SfDFPwIkyyVkjPxOdNJEW+EFE/L
SqA1f81+wKcPB9BgU1P+quiq4bVA/ZaFx+qiM7VyTzpooinM/24cS6dutisjuyBk
LVhWS3bpIXWSgWNuRVW6ISv3B9lFzmJgy2TCgNc/GCIc87/+qjPzIOcwg5uh2EgP
h6U7fH6NC+SsP4ufnBKXCX0Mu10Z3hUBQ7rOOWDvogmg4K23lRDYtkWWLMakDkHL
rDQGrJx9R2X6o7v4ywpR7Dk+Egou4EM0yoRyWM0PC/a8guX66LobBTm6NQUWb51A
fIWOUREsiELSAVG5050L5Nbk31eXY5d3WOExBc4np+pvg1Bd6XcnDsZuuuyS+GGJ
cKXEqfrHEbU14htje4v/rW0ZkWQoEDExBUfYFWyLzJgFE1fjULA7FUeDJJ7/JS+Y
cJmgjYbEGz72HHPIXLKXQtHsYOH7e+JVOAC1SzWCYXpA5T1TabEmNKe0ia84bmWO
5sgo6Ws/8B1hGSeV7bBjMOx4Kcl2K1vUBKf/u6AYnEK1xbIXVdAp8Ni1aHTHPRuP
5fEqkGMMkkUyyw5Z5jHCbzU9pIpyr3NEvc+YLn5083pvbbobzYja8gOp6VbuLgJv
Rs2aDyBJmlTy9QYog66l7szkCoQrWe/IG0wll/F6FFJl0yqoL8LJ1d00mVj3WwRE
kdInP/wWyTwUAgdlGAqi3j2xnJXrxc1+qjsjYmsNRKtjvj7EH30i+olg0S2bwrvU
3ykugPmHxEnGtgzcyqG+WPk6x6eXr2C3d+bQoeZuLOo5zlXs16SvwizwAtB5+45O
H+mGXKonYxANw5oV24CkFehe7UKzvRVJNDgHfPSZTe/TZyLoLr8Fz3vasJbeTCsV
iuPnIewabvaxqQfWxg0nhJDqVf/gdIFr+p58gTS8J3XAAAJm4tAZVnkWiNuDQUYj
d/UPdRidMdu8yStavvKLEUBqCdQ8+r2Hr34OA5lf5mIp7luXgeSg5m28drVtPW7c
LMJWl52vT5b4hBgKyGrDh3VQZ+L+8Ow+LdkN533Yo4DGiDHs499ax5I6gHcIG6RC
rieeV4kPibQl2KhWDtBwSE9D+QG7SDJiJYIomraX/b5dDk+Z2qS2FVEcDP04fumG
1GIsZQgVb8EZ8xrkO7mBrKYoLsVievuh1g5nXYbJsiosuKTpOHWyqJGOc+gCYOCK
+PP88ZzHnp+jOQYgrFAmpgCXx76JrY3qcAA/RS4CWYF6zrbafkduVZJzYg25b612
rhqJHKTENZfS1kdBmPCdZP4xq6iWU6hCh8hmRmlWJiRJANSZ0HCaHO7ICh9Srnsz
S+BqhzlzvHJP1E1i4M+fC/s8mjIoyPKytW+dau3qz9e7QNoYT1HMD8Z+ANBFsdKz
eXxrXzNLHxMMyhlwBUltu1KrQqVQapTRU0Q4kED7IwnA0tbOemNwtVkoZIxWACU5
nwC0HjdcTkLD4GBkwI1i33xpx5IFosyMH0OcBqOQI7hGkW4zzYutAre0ugWyIuyw
khIWzY6a7Am7Dekb+6WXhUZN2/kV9xuSWfYCW24Ag7Vhwk18uN3AR+PWnCrOSSAy
n2mFrUC2JWNqG3z8BB5N9mTa5ER3InO3dvc574uANZY4/oPb0MTBlMNqS6OI00fM
fAujLvQKThRykVgYr8EvnMq2FLJvz0+MsFzwvhWRmL/WsJ+MAnBfu3s++3unhx4/
wcteqkBXNVEWUS6bWJDpl3Am5vLF5UK732h095y9RN3wmp3i8lviR9M2NURT2b8A
l2Sc4PaG7J0gcRUG3wp/XhHuCo/dSYlnqqJyA4YC8N2HJ7QaqMs3kJT4zx+oUIUp
sgWQdcowhhg7K1HvFGPMLfG6Vge+0FKPehT1S+q+x7H67DDrqR/Puzlyzb4+vAzq
YSlfc/sf61bdp5TMFOKtYYLv6ipP3wqBMxJCY28hEdAWoZePsGb9TVPxdtCstZ01
IX6/DfjcoQPa9IJVLa9IygGWJoQtYp3sXhhZ/Lbcuyo14UcKAYPolgyEI6vYQif9
11peCxucWBlh8t5yc6n6iUj7pHxXVOAfSjxFNVaQw2Ivr76CLUlpa86x5jtn5AVw
iXBIK7aiQpriGoytwsJJ1ygr4YDUW2mKgh+b36Fs4XEo53xpqj3hTw5IrK2PcXL0
C10peaaP4zUWv3METyaJOHWqWOKulNKgZehG9o3H4Pjs8rrgVQJyBGtDIn/Ovtwo
+ngSDi+Bt/cNPSbH+kOEmhlfr4YZpb1Tv5uqVyMvaPPHmP8UXaFJWMLoGME8i6rJ
JLyu4mpUD3oNNbfv0zXCwE10Wn+EZ0Qo37If3bGfw2wltzqzeheMc43Dx+KcEag6
REQCJC3WL2CdkAGe7PoETvWIlfZLVA488JUPzfBn9VY6WB/jAxReX39EbMOvkE89
Pll36XWDtyhjl9e4Hk68pPDCTv6C87OEiuLeBTsgQEIsgG3xil4bg34ym50aX2zD
UeZVNZjFJKdbxGO4C7+vuKcbySApiBSPN1/57nJz/5ujACYMwFu17bDmYp5Ktdd7
fJpNE94pFLgnGrvQvQzFqUHHzsSeCm5HsTkflStzy08fnarHwIpgqOKBpvuEaCOs
9//k8h12onkSXBjXVEtgTDOQzxVLmxMJHggOWP11dvNukxS9yDn7bfmMbP7a/Cgy
9sv7ZI8LpsPwu+aro4idtKuaZ9OQ6Tcd+UaAj8A0dTcrXkIRBxPLH14Pq3mQWir3
zXDo2MnWnyKCHw4y5rukNWyLehIPFrliimQ6MMPyq5z/vNEjSHqC2pOWHRNUuiWz
abrGTVHDLco9cljE83iDE3ihpEK4DuTJM27u7CHrJPt9y0aC5hedURvl+rAUSBYL
lR4vNjXKZ/X++mZVKo+aPwRsKwcLfoD6fmmKBnNf0eXrvFPeYKvr/qccJErtxd0n
N11r4p7UfDxYUleDVfviTgtMJpzXrXOGqu5NShJFx/TuhHJxCg+EpFYhawXOmCqQ
rd8WJkWJwgrcoaIHoiFiBJ5aRGhiLoGQs9DZYIWEpNHC83ya44e0i5mkF1zmWZV+
1XoR3qKrw0ukYQt8LrZmWsaOkBo6XAV99NOWcoeXgq0TpEC5lXZiXEKnuMCsRafT
Q7gdvucN5KNysZn+gXnpvonyxqHfcTUv3JoGUXYRYv4XNAJyl7U46X4lbgcH9mvR
2BBZ/0VadoJpoZEJR7jPil0V+FeSUrnN7FSYPrDz5MMNm2gdX42iFKX/vfwfb6Mx
7d41haes/vbiskKKQ1SGScNsDz3qm3GYLp09uifjnS/akJD2nukaqcPOEpZ1OLIv
yWsI3oh+VE/VFz/zs+S2/T2TusVDC6XZ3YJrP3timE3hJpKubkb7oZ6nlkr/Zsvt
xzOcqcDFuvp4Bu4E9cqhggI0Q2ccdJp+W5xF6vaSyt4PujzTx7g1n5FaWjIx/suZ
gAcgdHE3DZZlsElpe1yigZ90BSt88ITAQ4sv2UCH7xjIOIKEgp1BFDH5JrobGdAg
s9aoJYF2QSf9eOtn/aBjL23OdT8ZuL+92fXHzskAfQ8JqYoYkYr2hiK/v0+1uxZM
wRagi8WCF2mhPJc4efnikwbqnBgT0kxaV6bPX9SOSgeyOp2NHiSuXOXCwnxY7Vkf
Iw4Al1JV2JrOLCsfx0C7LlShuSjskGDpaHOhljOesAMWeq2dPAprugoiR4FcGULW
RvG2v47rDp4EdL7d9sa1MRaOAcEdCzdSLHXBbQS3Z7R6n5Nfd11Z/C1Vq6S0ihUK
QR58k0fPrKrS7UAGiaWHWJcOgpvp5cNwKxG1BnQWBZnplhcoaitCFPdG4q70oAJ/
NaT3UYw+uVj+oquRgFELQwBwzckQmNjPeCGpxC7jniEEvJHaaBSBWQMoYKA66DAX
oWgkt7aYB8puZr/gVw4+xr+oHeaM07uewaS9RUiZ17NL7BX53MdOAI5gUecSSOt9
l8VTUiOV6V7+JTmpf3OumWktMKsTm4zJOqozbMbqe0bYn0O7I8urAhxnt9HUnTLk
V5TS27fyyo/GP6eXaG1UqoUUOrmVEEbhVb5yNI0CNl1PosHSZZoPLGl9fzS3i1nu
A9j4Z39WLQDVndK3q6nTSL+Ki9bUxVFVPrUxZ6NEwSMVRJOZRvWkPED4YWiAaKvg
P3uEP6tNoTyNSiCjNtG6S/FcdP430grwZjz/bhMFaALJTzQ7AuaNsZo4EMXVUC5c
m0cNdntvuGfQ5j/cvXXwxcwuZITRP6Lls4oyGSeapKQ5pnZ1piqnhYgDdqVcO7Sb
W+F4hvJl3IRGyKIhDeFjnbkjTYgUswNJrAxMV9pfFvaTzJ3vkJIKJdCUCA31LIT7
BgK0TNZsMzE+GZ8Il2dVzPG/UUS+40gKu39g3bBAqRH6VPb5xbZ7O551olXxSWhP
+h6iP5KKJKGzn1LYkug8GZO/zvPaMZ9Iw93CH6b6LSXUECBOC9TbxpM6HDu6dMjL
iA9PcOKBXcR1XU4B351maIpntdxw/upP3yiOCXB34JVWFrzEdVFojSNsnSQ8M4yv
rZW7padKkKLiiE1ANnQrf/g7q7i6MHJiSnR/e1Y9jv3/0QoCRa7CcyOgmtVsHOfX
TMEzGf/GVAmwW+vB55w5gMhzhdrVSwJnXl+7LG8eGnYMvUXD4uJdAiXQ0I7qxTOo
t0MzBcWi2Rw+5wOwkCAkIqaGCiyxfBIRdK0NVFxxWWdJeAcb/FVX7t7dA9pAHrcZ
aw9oM8d6FqoremuMKLwzjEFfMfi8me6U9yRjdYDpZ8kih215HKIm+jIIAK9GYYK3
jbkOSjEXWQJp0GwP0oidEQtX/P4vsNA4JXzKOIKUpDscSVMJ/mNqlQcd6rNGHjWM
HOzBEugoBzX5uoeqoaezXripH69AEewbqrqqzXkawSDcsjn8M+RWKKtfJ0TqlFxS
UEtBKOkMkK6pIFKwAZ4++Hy2aATCXwXtfTXgyETcvTkchxtDsE0Bhxw9Aw2sc7jv
KOj1iZqQJLCIX3Or+JclxDTYYL4rVOkJ3uqTIolhPzq8M5BRBwLpeSrhQVcvTsKS
aavaYVysSDkBHubxt1vNoK61TAZ9iCsPVsGRxb8PrO5eI3aQOq7RgifZ6+zkKXtz
bJz+YoJBa19ntge3XqajqOkF78NMBMPVLhLCe0nBwg9JUdphHWE+NVk96GTuWbbb
0iyJCoFb3N47KpjkTOFkTHEDs+y3HOC/y/UOji+3nC1DchJCblTaoitaK8VC3dI9
e0Og7uwc8y6j8Vrl1DMF68y9JqjxoM39xKb6vjT4kMuY8UKlG6ptMWtfuic7UCVS
cO3WbLNFgMRYUBIAr3yYvn1e8EBWkJu+MldB/ORXGqIpdGxSfm3XuIObzgQ3AtIt
e3ydevtEpLXBP39V/uaWR+qnbCC2iLIAy5aMLPVDORZohIkY3haCRJ2P1k9PR6sW
yE2ylbQeVrsntupFBb0rV4bt6F5ViNBwmtIM7Tod+xTqh+/Id85jHtfHSpWZVFHy
AdLAllk2UOUJrVr/XoQTowbQz9PaRlBYMcZk4H4ByDV5z3+AbwdKnED9mvgm02Dk
0o1NfDMI8jiheRkDLSIkPUKEWKH/9sUEpKy6aX7kyuCefv9e16NN5+gKBnRoB6EH
I/t3LJTfSCRtNk+jHeSIYETOaXlxh1Tpu4WPRu6Zqb8zMnYFrvWbNdId+CW9hi/M
Ak2zcYKpiAWup+X2UkNO6q1zn5hxo0v3BIW/mJpi08pTmLibkkkcTw2+VxBCmE6C
VHCGDBv71ieQqk/CcE6Clqaf105jA4doeHvkc3L4yEtRgQ1oVaxepaNnYrkAvpDW
gKAjg5J5AdqCEWKNtCxz0mu94Pmvt5WnZyvq9LWPRK7Q8Bt3peFJl2KdtDjvb0yv
seGHTuQv8+4+et1SkQNvhZyBGlhHaN+4478h2X+f8RjkNP/Fbvjk0ihPpO2iyapj
RINjBVFnBKHJQPy8L3jGPn3uwWP8hN4qrpJayt0uWer5gJca0Y1JgSkRcedaLMJA
z1q+odqKANW+S7xasfkufBaYIMTNOm+3agbiAus9YiAW8AuQPyuqcV3JJuJZ+Scy
bHgPkWFDotPcrh+ic49oqoJh52eBFSKbYOsyczsF+GoC5MjeM5oUo/dOjGBxXwwl
xHOnb/MV9HlYPD7P+dvQq7XDzB1mPnHMroZHfRdzBWkD/z+HCrvnl/rWxvXy+pxh
Y8o5t9cDE1yrJ2bd54YqyJqeMcfkUMcPO1QLvXm3iSySmBlUzWrxYvHNvcSYfkBM
z0paMhQquwXUokIMCRCihMrc/leDbfquLSbL5nHAaxMZYBb4mxr6Frmp4nqz+dx8
6VewTnmQXTwF1o5RCs5a3wMGZaTESUU5Tqc5UTJEZ3xTRYWpIoLSGYo8avludM9s
KFz+mKwuoZePgxiTkZHTLCkkIX5AmkZXBTmC3uy6Q1kqf0z6gIM046BBeIweLK1L
2fuRqHcJZW3tT3a+8UzM0DZymL1JQPFSSxTtYSaUtJMKYbn/ig+2ECxKUuWxWN59
okjeFpIBj3n7IedBJcmIttK5WWv7hwtjcFmlPy13RzAlugec2oFsLVei9zFl+pNS
bXkICU7CFsjIzZ1zqOtQcEm6yx/bFy9DWjANyJajIWojU0Cl6Ww196Mclxf8yUxI
WKuHnp8KY7Gjd8iXkKRCkYq7/qkTyZx6gJyHleS2FSq2qA0cG1lBFPBKikHpoSz1
O9yh666NTgnkX6DPHCbQphp7fcSLb64YfCP4V6fW6mEbu0HA/5CeH9w1Th7vRJIV
MsEmfQwhT0r+SH9kceiWgR/tR/Jx7j5+i92OvKB3YVDFlnmkK1Ax0pWqaRBDHtam
KgSXPijBFn44U/CvSV3/tcIoB1yfm2r4k7jaMyFzaH+ITOXzC0x01YudAMfzJW90
IfFlaQOKQ01dWVv6t/iFGT6pxIHADiTy9U90oOkc3rdMkRk1XwdCm4Y9+PTYD5bN
AczrLG4TKsBxOYmEf3kQgsYuBKWfTT2orfdeLfuFK8P5Q2/S2khPV6BAiYTfnXY7
/oEShaNBcYLl130bZYqybujLzbfwruBdZnuczisnGEdMNTeDJF7LEtVVmDZLw4sU
9fIHRJXnkgBwzOvHfWrbKyXItqn+HTl3L6AjXThkdffA9IIXlscXFDObrxjFsSo0
pSKL6NsVri/kTgVba4BQfejDXVQaPU3IHIGDv8TwPLScncQ3dzUDbD1LuWfg0AHh
sb+iz8XWNACKr5HCx1quBKg2MTG+A/15RtZhR9PM3jBgHwz4l6pmC49xqBprmt9e
dYDeu0bSJprU0OPVP6cCvGHe+JROqwQo60TFGgmDgwtspffx2qnncivDWpENkupX
DPHH6B8NcYW7Yl5ZVmJo7LsBrd8WJ9d5kkVawohIjG25CklXdcYS6j/a7RZuuLDP
Izyz5y8cezEaQ+5s07/GMZnVcjMgwhz5/aSzJQ3y6Up9ymuW1A29ab9iPxOGN0r8
aH0HBdJXXxea0whZJCq6y5grNYX0QjLMr07URAqgf5JhP5b3RP4iM/CHYqR8zh6t
DESjL2uLAr0b/ZTeDwKLpoxa3Yslz+nmviI+CXsM4r1R8OuvHrIFrEcUPSeJbJtI
Tk4SPjnX8SrZfuDwebJilshoCnxtP06R8UvCrm3HxRai/bZ9Kj0NVJ0XjID6BrvN
PHGk/uyNl6vy3/fB/g7pB/eO/V9Chv3tiTRr+mGMpef4AdsHutqAK9QbHPnyA9mQ
Z9C0C7yFFKhGyyfPbJPU1nFy9dmWDTo9I/iPEUiHMKg9JOH2lPzeLr5CJW5K9grR
j/f5kEnlZ/A70KY0/xY+EduFQRK6LtiroMg5HKhoVQ5cB767Of+0LprOGJTdTJ61
Y0cxZVl9aC3ktDpFnMM9NBBTewccCsF8lDIHlLUxLOm/AcNX/R64MOf5ScE6aiUU
4bWgl+ueBEmkasAZmTsVfyrkpJ6OBkEOpQz86zx4Z3ZOug+T50S4geGcgUugqgrq
KCM1ha1o2GwvnfhfQSi1LdV7C2tH6EjJ68pP+ft6HHVrA8GFBVwIzZc7STpbjokG
B74BXFd3Gkk0UmqxSMSCQ3u7moq8zT+bX0bHbJOJ71be9gWtssvrFBZNb86/dIFF
l89Y1mmFRVDLa5GMeSipp87a+RsQ7/P9wAf8T4VizKmUaQjX2517b6VbGBzM2dvP
7X8sgT32gR8hbBkJ26FZ93ayaF+5MDvBujjYBEY6852icB8qKXu3w2H3deqnDAjh
2fXz2Zyw0OC74sBWJ1g9EN36HLRpKCgFxHODe+VuXfr2li9ZBfUkBGj+vpt/oDy1
vAfCiwAdM4WSOEyWI2vYLcyfT1sR2sHkPGVga/T50QQm4fa7SeQiw3LbzaqPo1if
RDnfcYPwtDFEbEHOC12IZDasZqS0I9fDfOat1kWQYhP3qEBmquCSM6uFGzWUQN6K
wZ8to0kz1EQQfvYV8fJPOuiTzO115v0aMANVtoIODJFneoZtmqVJhKb+o8+sgQE/
aO3H/Ti9auZCmxnR3aOk5fmFksubklzEVQ2JjGKADJmOWKvhvusNEvgX57bwBoyY
3x0lI2WgROy/uE2yHS4Xes6RyuTJgNtLQ9wBXX8KcRjUlIFnze6rFz5mayv9MVDF
W153MWb92DY7H84J3mefdJluXjy/hxRlOX53CgDtDgbh2Y88ZGTmPE1HLO5rarr1
C1zGnWXZ2t8kp6oFl3NF8hM9bJeCGLirDYoiDp3AJ27sd0rrpVhEBw1rW90F8Iji
pZBGy9wk+m5hzrqEh9vo8dQQ9pc7c5G1grvBsZNLYW1vLR42cM98eGRJHnSTThbE
NQ7RQKnT0uplpJ4KgLY9kmGtNfCPnivWshL6h1AUiCjqmn1BOBQd5H/KXMr3gPpp
rd4qlI8THX0qN0xjxz35kg7nPgEzPhxw3IpaqLzoQjAwMwc3i2qaKvO/ktTHofS6
TRMy6iyBJEybe84K5ImJvkgtCKUOydRTI3vQbKmc6JH0TJTmnDlsseF3jl9wav3V
AxQMlM+/Mu41Or8x+r75I27HijiPS0aTtBL1phmltVxuyUOv3Scn+42ovCH+XDIR
Xa0NDluoxf9F9KJYpGLRjHeAwR0LFaX573bQviZsEcegpuR93w5Ho0GxiwTOUeoX
BPIXpk3zItYoydSi+ntztKpUvACDM1WIodyxBIjD1nbZBwE8G3mKMHuygOWlRUxB
mDiTnu4xebf5cWCHg07q6MZ7cs7/k91+lSx49/xFu7Zd71LF1ofKVFcVkbjc9vkW
cBxalcgMvncvVXoAXzLPF6EeW8nP1mtO1FLrXSzvDxgVQ4lp8aUya5VCjeM1jmuM
D0LzjSdxBGuReqWKCju74tg0/NXWfize3DhgR3hWUoSEqZ49LelJ/TE373Hi//Pg
ySDQ45VCKFjE+hjkjWcdthL+mIryFHQVOk7KnHBr+O5ShLNG4LmmSkFq+M5psEcB
7xVUaSaD2n2RRC0Tdfo4iMPnbjmo7/Y/Kmmm7noj6GGNRyjmU7z3mkFeyjHLRqwa
iH/5dNHRwpuq0ggH2bgGtKS/DpBKn1TOZD1zZ6/Tu7hQ0pYW/DLBKt3Mh4KHYZps
I9ei1JVboJQUYlLgZHFbgvG6REWDRVNdofD9cKtWD6C1VB6aMCdjaZdr5E+HyQsz
eQIDiXhpFwQNG9KSL/iaHMQgfoO3+u79qNSbWvPVkRQpA5CCpBqi2rkXwXuX42zO
3k0ZujzgCbzg9vo/krbUoLHPjqxaWPN7pTcW8B4um+trQs1pwhAlOTPR80ZQOwt3
24GalQuaCQjRf+cqAiukMDe087HTOJsxBxEtsZZaVdoxU3EtTRqoyd25bwDZLKGy
V5fp8ZFIoCY9g4EOABW+KusPv15Vu1l6GerP31qr1scaCpkHQpDWAdIT62BAPQN0
qcRQTiAa0gd1XgXq8FH9fIcOSd4wl8DBp1iSiuXfY/Im4ye7vPROdaOXz6irFa52
bM9jXsO+boklLmnE/JE49ojM5CdalR7gs2Rr+YGbz1U4ehpyj5tPwWCCroU1+w/5
cU5pLdGA7gKQAmR8OMoTNQaIsQw/hTwPrko5wpnQ9wzynOkDPbQJ/WLK++g34xQU
7K4Z0rzpsC13eFoScFEy/5skO2xoxs8OmIGjxyqkvRiLJyFK0jtHQ9iW9hqzXW8l
0PF3PCLAE/YuKpoK/AoVnUQ1pkU75werJfRkXRAnNSB/d72Vh6rHfDLcp94+D7JY
fiDgWC8WW3ETT4sUStCCGLvtab1DP5nk86bowJl5f+qhQKPHXHV28+kjYI2N+66L
jJ8tBv6qhp6oj5PpGIXBTtGZMad3Hc3DTf127CrlodWHpmF+DZpTJU0NK36I8sNm
JJocA5mySCxxjPfiKWmujLAr1EaANqy6MtmCnuPWHXs7fsvyKV9A4zoWWzC9EoEf
05Gk95WKttGRxZwBLIZXUaQqeW9pknVzkbs3+3v8qc5H1wqpDhPxULmn07GNz+y6
431uwa09aXt2lAfZl2FfSm0iIgtneoanOOydYqa2GGOA426qqDW5nGMRWsU+54/E
Gp9Wov0lSgDzNZ/Ln9QWbhjmEU/npbrhwYYy0ScDmNErVPmIqq00Fc8W9YOHMjEp
7oUiw3eNjmp6f+qOFlc0zEoI9xALzhgHorA4UKSi016IA1mZw6lMxHtBwZNfgHyE
rFL0FA6xkH6/UMtNmIiF0YpdKtFngU5Z6rDU+vZkWQkKFzTAeEY2qKAlnOC4TFIP
KiaQlmTgfHiKKAGGvvlZPBvCyilV//tsgmM2QsTL59ePnqL6E2ONG9aQWebz5YBH
hhWtMOKgruprtW9Ssl+ek0TOeUwlOmH8p0vMXoJKn6pvLsmtloJNJaQqcdHDCjSw
0Rsl8Pf+yrkbh4SECWMyNPqpXP72GLyiUAb+k8yNjJKX3bqyV+FrGguAHPBIA8fO
j/BELK/51K1w85evibXy0OPdmqz7vQDOwwyjpNhb0U8l3ByDB6/Qh3h3vNnEc/d2
HMaHcMKjNLt0AYFKRSmhhIfVOj1PoHtLQiZW+owHLAvFFQX9vKnUbTY4wXT7E2dd
SKi8ytIO1TFUF5M2I+gPTOduRqUQQsxDK9e/fpQOTUbDGtBLBX9YctUjLBssORtt
Nibl6d34Iq804laACDc2gF5cN+AFQChqog0vtWjku/cxDCD6NGDjmXHmGjC0Ftvc
anpbuHhXMY3gCgX4ojDS/zYHJd+iwUv96oxingK75IKYfQ1V8Eh64ukaFAsckumb
zlxVdHa/oWx0mPXEL9T1pLLvG0VIKUuOJXwGOKjJazBVsZ3M/SPnX1zQVgk7kXlw
M3FmGBOv3mdGkm7Z0TN2W2gpOBOBE03P2+PrN0D/jQyoUNF7ePCOgmhHGxJMvl+z
WVgKBut9drY8a2MbVjeXoaer3tId5bK4PtSyWgAx2Sf5JTtXV/sYYElBTyF3Ta19
tEZ+RKDe9q3P7I81UcC73uVHL42Yqbq6phYvJHXyrcv+AdBLUheFBWoUbC21jVn6
aA34v5VpPJUc1ED67CavsQjKXb7icYkMPbqKJUQhYB4TA17rY6yfBr6Hz8mnZvjE
mWEDl13CoZvQqGAW6PzKQpZLfKwJkxqi34vWOfGENzD8pyBIJ+CzREcD4ym953FR
Q1M1IPqYNUvzptWfyfJp7PUDFKdiQcnYcDTo3OyzRI/gr5lDUKrAt9tFkXHOGEhD
rq1WTCLpqT3RUBl6KkuFgCCmQY2zGjr0KJ2u0u139DjjbrWJ6SJbs8NIO5D/bWJu
f2qe6SwCknnENVPQPECVa/7Slk9/OiwJlJHr2UuyA31hqZnUg+pKPgULJ20xJKMB
Ajv7J3rn8sTyx2f1rKizqO+A+zaWHixIMbDtqBh9tv6cJq0Ce+Ocoq1GvHTQyJBo
+eAxgwcewzQ8OMIYYwsrxjUcwYoQWfRAeddr1Be7hfzH7PDRCdc74lywIVNab+KH
btcrMO+QAPqPr2woCKxZ8N/NvOT3QleyHl3yl7y0PXqMxChTj1cv+sK/p0TUyfc7
X4KEKGL9VLspvCuyGZ55SDISWR3YGOx3Gr5cBEGmVjkvTI7p9p5ADslqE8Z2Fvao
N7k7TgCEzzwc9sZ+yZ6PzzpB322U0c9zVxEd/5jzqJZmXxETLVS6vs9bhDl9brKr
id7vk5WMUxsKqK+wE5RiuAfFjlHff0MdabfwCb32RB3mSwey7NMUVIMd1wE61auN
L8Q/UyPCR8gYKbwFkV8N8MLErapTVcbO8ioiXiRTHuekKREP813cIv9bLB6nMr0m
QvbyUI0+/+vr8MX3KKoWa6IxMOBlLJ3n5pUbTmmj+X4pqI1JW42fLNNTfrfcqCzE
S2OH5m+Rhvgx2gcIjGJ1LXb1L21noJJDrkyr2WC14QSPdQ8KIf6NfEDzqazq36/d
RxsticSAZoWPNHKpIzExj+h+4fzFilPOC6XB4iTuKBIm5CsGVz62O3nbxSKD9G9y
gYIWYWmmJY1/lEd6SFesw2AGZs3zhDkExgXaVHSW48yZjz4H95h1bwXltvqhD6f6
g406OeCheYQlXsf3RLtyb+Esv/GyaBshirL3dV+mR9auFsfKVNvD4Mgj0+7APcpn
I39hncQZy38J3itgDwEs4mv+d3ORhJU1CgYVYQRnDk/xIiGdvQ1JWOU6l1mht7PU
iUFKfL3RAxYllkLDQBRFVnX92GRX/WZozxaCeObSOy6IN5lpTGrviou6VuvRUOx8
cPWpLK7F/jML7Jg4i49S2cZkGb1REMXilcbUF4AvFIXcE4DQNJWwMhv88eRdsULi
raIJtLe+uNVh0IgnubVgF/+5AVX/jMJs0VhmY9o0vJruBgD1xzeE53FRmwRtubw+
Kx8Zv9NLkmlMb7qnMGZsscwg3V19vkw4ClEsFf4762MHQxM/sPwOkMBaxoahz/Oe
nbtNh7cJf4APjwX2RWUYYcqYWTT2nxu4lfD7Gsq6HCSgvad0bOkNdYCzIX7LPKdu
kBF32/8Wp5d2owmPcoDGyJOwloaNjnF7JNfu+mrl+row4XgEpvc01sVhKG7hDWfT
0zxqJhCg3mBywnFDYqhl4QM/bhZ8BoroZ854KNGSymlMMX8TbHv1zv6plztxeBzu
E1zWS7C2LjbbJYe+tphYrTmLwEOZQNqRY3GpHVRQKUuDyHQSwWcxAtOsyVRqqvho
PI+EEAHlgonUSGOOkEbXXMe+XpAunw0A8yuLKSzusZPoCEFfdIebL8FkrS9U1oDh
hoKExEXYmmr9PqC0e4jltCsLPg/O3h0bbf2xur9ILkn8AoC4kAyPTtwIiIAPWKYX
ollz+n1yx5SUoYfZ9AUqrz8AcVFBWr82OZRHiIMwOZAEaq5uzmq+1lHHCPGDW7Tk
dI8+P4AcIq2KK9TvOa2gPNkaWj4Su/c4+okkmwK6UyR+XiT9muHypf+aH8GEdGH9
Sfzw18YLrqW3FzyA7CgQA6+Wf4jRwd3o39wSTAPjN/u+iqOdwMSZ5F958rzjSt2x
Re7dfFqWVkEiMx/YVqOPKequ2dwZ6AmST8rKFQpkSCZ2XdYicvIsEoHkitHcPAmI
PyXaCeC7UiNqJ6zaim2Zdxg4DSpjRNdyzxOJN6YetsWpUeKOV7FIVbgY3ClsUG4H
D1qFw2kIhtjr/t3zQwiaBRbRRcqaNY0VcKNJ6453K8+gKzcw05ev6JfV2Wmgcdv0
K0TAkiET7HZAv6iQPfrDmer3cIRF+bvwRxC/xXeKVpChbqz5bVzGQQWXMrUTWHWq
mPxCPPSYSTJEciF/9WIYFmg8AAjmtVGFARG2tG4dbPo/gcE70+OwuoWWFEuVCXdg
S+nPTCPAfnc1c8Z4TiqPSebNA/sBZI08/YvG+I+uI0ytWvabhO2/KFXr5SLU+Cbu
VIv7FFnzVWtYvx1a4SXJQezZbvQmlFleABlvtbPvFXV6RlqMTQYM9tOT5ifpiq6k
UVmoUm4iMEIKRPgYmgEL4K/7B2e41O2gtJg5Vpbw+syrhvkrSCKHLorOZZYWjOF7
ND6j7Wp/RfZZa93khnisQSbS/YqeX9z2pDNrjK3cMmwivOCbKeubtdi7qrk0RIKt
YJeSwCxJli7YKZodAxSsWPOju8UqE9syilWTH4eFWJXfVMcEbjZ3SEUz6qDb7ldz
M9Sh9xvQpo4L9BVcjiO7q0+ZQMWLqC9Bku98nC2wWRwKqspHPEb+fbeyzVu8q8Xl
BUql5bXH/+0VzV9ScelyrHeVnMqcpVR0Ri13zhsDm8d8WkI7fzPTjjTXQtGxAnyE
paLHU4xtKzJ9rDZFBluAUMyCi8EaoWWN+JgcqPte3JucUvZsqIsyKEnmq+Y1wEjY
w9Aq0IOLVvag1Rw/HoCsPZtUpEfZFjR60x8g4t00zBpDaY9+U6GshWV8KsXg763i
ROHlKmF9/xyxnY2gpiJPC+PjCPqBrqbuoTCzY3byj16j6TgzHwv657Hz2DtXAJot
mVPWrRffSlvRa6A/nFMOFFeOO9/w1dAorWRybOkXW1aEx/KU+kpAqqicSMTyuZ8q
jhxoqFsHDm42EgVyOyGaPnp8sSHeBLiExNrO0dxrIpKkVt9lKRnVxwnX5yPMX9BJ
E2+fBqghqMpaaAF0H6uvpt12+ErrAH2y1Exl++zDuYBUIxhobSVCd72GLTcErX7F
Ieg+zM+CKTjZnhKudH/c/Ogd9PAzgbEi2vmZdPrREJgHGlg8z8m5L33XeF9jknI+
eGY62u8vSudSFH6TyC5jkCNLTei9cWx4E+nSnjJpWsVRTQkvuK6zHsl4Uz4u4WSc
h1KEIUJSkcUUJNuMAjE/dq8sor8p5z9zhBmRHE7Ft7THVfjF27CNFjNvyv7qiNZv
RUYc5g2A6l2BtT7ATa+T82F19ktA5YqvAJsIk2pkPvGrjwe407rgVW/qdrwHW0lR
Ms66iZBdmB5jw3jlXsPWsjW8ZAhass+B1F2qn//DTvR/onso3aI/llnNFnUczF0F
sxiU7rM2zhlmAdTc7voG4GIpbHgDSmsuCOoWFc0BKLnTNihC6Mc1lA5yHOzrKS9N
maJLw/vtDce6y1ZR6RAVx83flg046EE8AAbw5t2BSXeHQCcyyzsLa2It0fdHrNQF
jxREdFD/ELorkzQXXZrAxyBSXXNzB5AaYASxez9US3O2a+14mUdcTe3lyjqTw6pI
/JKxKc7AdrfwA6qu82ZSspGPakrv5ejvt9Ie4huPeTu+vNH6cgSXapcXZKekAkBb
dYbvVWwXK86klzTuIxPZj6ACISp9ocVfjRO0h2wKv6NefZuiyJGAl/T+asCIw/93
hyFy9r4p+9wbwYbtfMg8BaKkRipHwesDkQXqavneGPTG3zd+IjXLrjwcRQZEWhaI
iI6HU2HhkyXWOyO39R5rBo3nso1+axjTWGLWcsE50apU7feiY9ZL5ZB2PQ3vr+fl
fNJoqRFnfiq1x5k08281cWaVbsSRIfQGjI+z0k4QAhremjnoJ4x0JYjfHWiRMEZf
c9ETS7td8qZ799trlTvHVQV4mg0UU15gajbBOeIdQxwlE9oH+82z0jRY0t9Rspb7
VB0KvV32NxxSURRL/9xfxTvSgLWUC1lUDtR1vXGJAKYvoaDJstixdoBOeGct08kW
uRiH3ONj7vM8KH4oyqie/ePSibqH0MqpaiLDvSM0DnbhvnX5v1/k5f2KalsZAfEw
Cib1syEv5RngRqRCuvz+mBNDimWblOcyRcmogYEWzME68qEWNf3YwjeNrIj+aLUi
ytcrUWSY1YZX4tAB0AXy7G2d5s4f6XROrPgejCvN++8Er7jK1YaYps1HSpT9VZRi
c0aiNEIHan3Ca6P7mKCFUgsMs+cofulIh6H3CYaMN79ci20APyIR3v+wCorqbnVH
ZHdpFgeKQS+tpbrhWel50JG0ZCaFuw75FASmgFqZONkOSLwuARRW8xm2gb+PrCJo
vIxTV28QEbGKJMGv0Bsn9T7AYqa2sR4IxFecf8qDkAdLX8gk++wkxIIkieuIAERJ
OHMg4Ft7Yb2liCaBF0Td0AVixLSB+KO9f1RZBDL2qYbuCdEZFgAK6+VwTeRo5sen
GCcej544QomxxBLY0KXwig5VjCa0VVs2HDiHeByeCS1y9Kkk5XCBTUX6EV+xDNlc
s3pBeNvE1eV1VKxLMUNA4gJgUOhRv3liRTNf7EDbtN8fkOXtrUbvguQ7azgGaT2U
i66xeK7KIjBKqkaRWUi7K8KYEQTGZLjBS6PdyHVviMqgo4XDIhCrY4xQJMWLoMne
TaJWY7CULFqMvp5Yq1puyxgVeyQLqkjugkYIZ7KcBzchsFWCa0XWKpXK2uAJ+mh6
8ic7oRQ8jqiaDjQkgW9FjR+beT9ezbLrGm6eLQG7SNvhw42obBiHzqtmsOxo5ns4
67Vw8jRjCJ+uUvl/ezraCgMYMewcfaTADK0A5GQkATUmoINQec/N1GHPLSN5U1Oi
T+CVd6MGgY4L4H2hPCCttP80PjUhMXFBZE4m34H4RKhcS74a/KaQeYIyadwkLO6Z
rN9k4D8iyU4P/3VquuWcQTquMt8uJ6snNc/fFuuxDiO6OgVfUjtDlpOEdM2LFBdz
dykbyY2TT/rVVUuwVNgfB0D4weNgLm3ADToVR1gDLp0Zj9XO2mxlejAdMpql9wOI
qLVDAgAnw6ohPULo/bd0AbhJrtEOCEKyYW0qtEGaAV5dqt5s3neqN+6apq7ct8Ha
T+bbWNudxahdGeN3vw5nfeKMNSpCFp0i8rteyKu960Vg0H9qa6e8+ZDN9RtAO7Y9
n9fqXoDRl8qnFNFGrEm9OwYeT3KkU4DXgzcjJn/hhveYlpJaNDejvOs56DYghRPJ
9FV8IVHgiiC+K6gEvy6uJpRQSNvMigZ2596DMTJCAw2+WyYnmCmfgGaGjVoeRnP8
/jhPsHWRr/CILo4inMnEHW8TreFUGZ5QLo3UhLKOqz5jeqlCiEoFrgAlIh/IO7FI
SDuwkSbmhyHaShpxNKyfYP7ZwC3zxD7VIYuQasZMnpvGQYuflOdiYXVvQTegFOVF
a3X4uEVRN8eR8ZFDfKBryB7l/tgFpMiaB0FtsWFhjBN1dLds+cVOqZTKFZpiFIkc
enxy/EWqHq17KBmnFP1x+FTY87lHoanxJEQ5lFbHaDm9WMTvlHCQc9FvZdkB4o7m
PT4wuVX6z5TJR3iXjbIXQprF5yDsjz8vOTpsM37r4LS6Qc7mP0Q4O27RjulpRFyK
WRuIAdMLHNWUjl8eRHrrrQC2eL5JvYrwyFDodWG0Kd0qj7hFbXD5XMOpNgudmRIT
8gFw3eQok/GhSTiaE17QxYIiYempe88EoLSv0EzVBscnBrgwkptE2O2bj3az3RJn
9bRL5bmyYzWxodmfQc6VTqnfUoedaZOxEbZJqBPOkWZYfG1uA5J+TGfCLrxJPYE1
5q+X1O1ofDGwPajvmJsMNL1KKvWyoG/OKZddd2jn7+uvwcC2Pz+hbdRi/FZDDNLH
ZxhWlu1ttM9iBw8NOkGfY4P/2iTiJhHMBleWhvmIiRrIkKS+lTjnxkQnedQtahe9
izJC9WxfL3tDVAoyXJcCHb6hGr8y7L+aD/topK7kjiv4VmwpRsoo3hYbPRdaJfCw
JMss3uh74SUCcNqXOKceBlt/FjERHUOmkQnOhHh633DVsTl5KgrKV1gGHpWT3YmI
KIn4QL4lbjUdNSSVYzq/jsfAydQsDsYLN0xPNamUQ3deYXsNDKFDvQsrMNMVCL3e
hgMZj7UjKeZsfKfNRVzKPYP9KYmGJ5XyP8j6Q++Ve7lEXM/LiWDxDz9blvobZVI6
56cYoo3bs9sZXn3fSX+JBuhJwcqpqYNSd1j4cScUQDMbisxVbsCeHT2g2YcPn537
dSCxo3JtJjZvYrYbqsuwNBHZ0bHkK5D6VJtqRq0moActaUPyHXuFEJK4lYwSpQ3N
3ERxcYBNytcnA8O3kO/Db1EiFD4ZskFL5JPslaDu3+Ej8hSwSrGkMaRnrVIP+3o8
D/1E6yFs+kRua1G3OerIi+ZqEz0k5K1s6LnoVSNIXHMunVroi0yJJ2IN1mZgS07a
4UwQ6Dbsuiic/dlJMPUTAiRqXyX+Ytrdgi/eImubvX7S+/fKcPMF+4VhXuMQJ1O1
yvq8fDyeiWkia1rjgjaLECGSIESPTN6HCh+h+5INrG5cl5kgLtb71hrNsjN8F9R6
FZBzjvqR9MTOgW+LyPugqK1SOh3GqrjMq0rIzA4ZHH6oDkusoOv8L2H6htX7/kR8
Kej1zenTiUS8iMl2wvSdHYbQiJ9lSb2SMguQ5i2mwx4B5/MNsrJEyyBCVoEKNUl0
M5tlxiPBp4AmU+0mFW7oCb0Wgzugg8PT6CEHbUR1yJmx//d04bF5uVQilv6Kzmm7
ILkNqpmYsI3sy4ocsc+edZICyjbntmS8qkTjtDHsQWKGXKk6tV9lByxxz69ePrx6
T/hZxH76YcNvo9nmYBQ6XBKlTl17MGmKuDD22lAgobN+mg+0vgD+PvYDhvysgU3S
dtawdxo0pk7eLwEfYXWC/WU2D8Mio9bgN9QZZKWSRP9Q9DPNconvIx2x08MZ774C
kQ5WPGzI1ULq/wpvAC8n9fbkJ/xDAwVjLhVwXKSIxyfrlRW3foNK9KRWkfk2xDsP
xKAsip41kefH29lnsQCbI1xL5yVH94Qx4pSWQjFvhfdvA3aP/bL1dMKlkdznbDnw
1h+bgyk3GHCLXUUnUrfztKOipKeGZDU6rCD1txPqj8N3wRm6NNxe9VB0G0YpWTm5
SiiiCDsQwKyXjfKHplGnKFwkZmtvM0UaOdVCsbsi/eQziBaMRp3BmHy6Hg3QeinG
i1sMJGsdmZkJ3bD+vGgY7QXqYtNp9fjCoqSTsnuZ+ZrY+34YvE0lZaN3J95Hon6z
6nJMn52s5raYFQ80Uyx+gLq8Z3Df8Gclqh8EdRNTTteEBPNTcbgYBelp57nNntWy
AxkFCHsQyzLAB3hpD9Ng6PiBGVzeKKdE+D9G/hVHhhcRwK06yDbD2kMjxI+jsnay
rWDqYiZ52+mNdfllgpCjHrZTADt2dFGo8YtYAqKfxV85iMNdgAJ+IIB2aJ/DYKPo
/wP9qOYllJZ+IgoIeYiXK953AD17SLtEG3dZl6LXyAlIEPYTXzegMt6qCeahtokg
ejAIfdhw+JRZ5TIFhKnmRPnBqWizx7G1njD/1TJDfKx/lNjD9+VOIzOLI8+pahHe
twTJchhVSSjCDCyjRvfUd60O/aqV5+PujiUExAcA4OCaunUvpMw52FOWj2Hh/WtK
9fLByQBvZ2p2808EYQqVivHzRcjQiYP9zYi65Xda6dA/4nPJI3Sul12G3cr4hf8N
P1exOtfwoIVZofKv/mH1JjZCxM7YWWieYQ6qPWt5Rj5HkOHeD2xnxOTxaK134rrA
4ddEf7ONdZ+ilxD7aJ9xbF0q0g10HhZKqRBXBWnY1E+amtHV3ZSlcX8M3hWUuReT
Ep6IQp0kx41jSUVLT2teTQiD/QK4rkrALkc/sDk8zlFnbnKMxQxDJO3yVLeQ1ZpT
lilCd/uhIO7Ces3gip9lRNrvrNktDYke0T4iwvXI4iokCDAZbNxaJj4Ec1w+K816
wEBMHsNbD2iPB+o9Zvnvn1pOmZJM0v2I9zQgT1eqSUf5PH1o6Xjp/SprP5SecqRT
f1KwZHKyoU0F3go122WF3A8dhsI5NrV99gOapnJcG0S4Wyaj3sXPNJ/zFKaqEU5i
HL/nfyJZod5Q3Rb4ECkS/1y0aLH7cGCQ2XXRZz2N1bwdMGZJO3lw5cTeot0MLglQ
/mvHGcH2lojMevPmsEkeLhc2aLjYBTAJy8B1KjhQfRDLDNkwlUG5mxBP2p5STv3Z
Lb/+dwLWWWfDzCpbrI9c40oTehXjdX59XA0PvqIKs1O+zsYLA1dbWtWE7UHIUANr
4n34m3F+EQcsgkGLVoq/06xDf/XEv6PFWch7Kqi/zmsxKlJ0auxs9n0wvETBf1s6
73rIFk66iYvF/V896QVUJL1duxh+0ieVG33l0fFAJ5nNzXruiv5ekv2x6OR0GiUy
yZTudmrLhFCcLAhCUhJg3UoK37l/Hks2HO4I4J1OFEv1+kUA0SatzZJ97zviIH45
x7CJrcNb65xVkiMjeikB6HCtDwYhMqWyuqBm/FfunOQFuMWdIBmmpOCVCzwYYzXd
0eSjXRPOPxSjuCo25WDuI6grgeoniKi/kR6LwS/GAmaiGT6kvBoQvjeXeQt90SgD
y9SoxdFsWzO/Iz2AMG25f4RSBnEVcO1nMouspUIXytxZR8YdLK8+as4CfdPxSCrr
tCDtM3RYcSm8XdgzVyaKuHhMpdy0g5LnMytkd534vm41Pl1hlONJKQ2Bo5lb5S/F
DEZeZNe2Knpu2sNfcp6TebBk1lSBi4v1bWWSz1JCb/M4yj/BN1c44DUmDmOitmS6
G8mq+Rzk5s4PT8I26RA1S45D/BLPehCts57eVvlVnHDtpv4e6QMkcSEQL4Fv/cWs
ihULTGdzDUFw7quN8oZnguX4Ci0odUhPyO+SVhMtUVk5JAjtCOlfp9ZG+juvVUht
xliaaJItaVfxzyp1+lm7wvvj6G3pCeBzxHeFsKJ30xN5D4bUXziQ4y42xX1d3+oT
X2Hqg7rvgUeJ5HNhIRIYLfOtsyfa/Cgbm8D6RktzQ+BtCElvsoKGJE+Ky0wEo9+L
Z+1ngOj7q1BqiS1NGwpbMgVWJ4LyRjuSaJZP0nSjq9HcpQIN1SpJPf3YiCMSQTDz
HsdCipTKuC4wb5vU0ja5ATyNXd8FbveA4XplOy9++7fCh50nm3ipBxzJlIMkD48Q
e7PPqDVckT117dZoVb/9Gmn45bzy0LocBcGa0UmnsutzQrJmdTvO3S5JsiNepK+V
VVb0Wd5+b4uySBncVu26zQEWuhGDnyD9JlO07B5cWKQoOfZqsjrIpYX6XCfkC7hz
W5T6+e3JZizkblHEkea1aGpj96eZv9cHxLnug0V12qfzmzPs4BgFbOUybHcx0vGD
9bjkjAZSQkyCryIoKC1CWG+hn8As+eBsPowiVo2BbHHqyPFsZV1l2BUozJZGbSx+
aGGEi3Lg1591swRZ1XJMOQolgZRQgsh19wPsWGgLHhvNwxbBmrcTgD74UZmIdKwr
rdfS5FBsLV9+jXSSKy+8+v00GhP/hHqgSoIfw5VKKT5DsnWscmhKyYDRtZIX4mBn
qmTtf2BXGvk9HMjdRkHBOKYEhpcLg/n25+Kc+Lo4MwXejUqy/5JNgdbHStu9Nef2
VJ7VN0FTQvIrtvsH7QjQm8XikbkbuZLATwAUd4aioNQYhXLjGaOnesrgQBoqkgLn
1jbEUtWyhmdODoGQiej7F3jUQJBa/HsUR1u0/ohxEBeeIKG8aXU6DwEryrMv42ZF
kh/i4vAdDdE05FAJalSxTnd84IkYITGz9DFjUD1X8l6fRKEbYpkN1DMBF/StbR7L
wVup5fXjEsfvL6m303oXR24ANY4w6OnTr18jR1fRX0vvj4GPzGeNpuk1RDxlM4JL
+iErHk7xhB79eoxsLkaNuFfFBeKUFyefzf6qkVshvaWY3LIv/UAih98G8twoUHL6
kkwYKRB2hSe8trdwURuiBvSfBd/M9Yu7k3Ej50sutb+GEBGez3RGzAgWdnvh3SGm
FlqJmoY3pki2j9DM0OYhMmlX61kVeLYd5Px8KvDf/9tCU63z800A6S1q30Dt5jne
X2Pqi0xJgoGP0D/UDQoxL1n0rYAJNiE71o0YMgwNhCnhabTlGwKjtO8Fqf6jH2Je
M/etoYiZHVVQ3arJ1UxjF1cwr/ktL9aBFcTgmxA20iICGS2rltTuu8q5R1HM1Y4I
JbsLxTgmY3r8Th/YHCUrnw3S7nS8fTzwVnbOTO66LOBrP3IlUW6Y2X6nVvn4s9mi
VurN9ADrBO+g6UXaXPu58sZoltA0b3uaOkGReiKYpEeHZs0Y+oDt3e/CqEF65Rw8
dwbJcOVPx8PqIDwoMVkHMsVZSYeOEUlCiWXZF2FAAzMQtmHqQ95Butdgxqu4zffJ
Be3gAvSk4T5eWSc46hAC8kPvWO/oViKcB/iY1sMXyGNAUUmgEDAK/fMUzQkMDnXq
rlt+ShJUu4jB1WAQM3RCDic6RIUp0Rx9qN/L7GTbKUKZldK9VjYJY1sqt5vKA4te
lsBRc4eXXESUhGBcpVO2hz1HiIjgKZClhNnzL8aPU0Zwifdy0TgTwRBHYX/enoCn
jW74bBSM56ZC5gp+KjSGc2UykYjlq4hALc3lM3gxonMQ5HMR4q0CDF716/9CGPnm
y/tYyDCKlimjZH/aaGXXZ9Di+EpEucu18CILaB5ZdaUgnh0BPSzWC+J7jWGqRGHQ
T3emVWZIuDJ3+j1YxtzL8+GkowP5g9t+d2hO525IuHwyc32Y3ZZPRZZ8HOBvhH0i
TAekK+rECDhcYUsXzb9QXtkpeMrjmimLNGSCvoxSMKQb5Qr7b0tDDzyFw47F3F1g
zX2VxuqycXk1KLkEVtB7HyhWE3DA4MFoUxlbQuqT/vE/fAoGByJzA5uCnEH7mwkJ
yvPd01FLEnpC7hFAnE1mjgHPMBMqgdnsZt1JZFWJDPmD10ZsSjc1+Km2NnuSZi5/
wYnu99e6IRP/rkqb+WWLTZE+iGyJGVvSEd5L78pwxn7y5qz4HeAvkNLojdpZhrK/
mGX2oyjCWnVm/rH6B/LovJogixTkSXcXqPrb8RmMMWi47DyYOGgu72ZcJgNr70Tj
drADtl8KeEE7lcQu7XWVn5vwMwSHnhns4OB06ZPu3U84kuIZVt90asUrpqc1nJA/
SySSz3s/xVl+BwNbCW8VLs9HbHOzVCxHps0M5lE9Baiy9zTPXyVHop9VzbJC4we3
Ihc04rl6JDJCIs9Z2utcJ7caJZujMw00cH2Ns+XtE2uyHIb2FUAfcSj4QSZCEZ9/
MrQ6YpkeF5O5Z1o8E8w8WQ8YRVrwFvllcyIfLIdb/0FI3vJ9+VXN4AffD5Q44ESt
U0D3FlxKOotPwsXtp1LHNVXtxiWgCD2YsSXyc2FB4QypKxhVtSP0x/ce2UZVzBTC
9jmesR3B6C0pfp/3b9Vg5Uky0ox6/vpiBmHK6vvYavvT0TLOXAVZTCtTI4skzA97
jZxHOIZhBfR1PFVtQIx9QVpP5ekRi2YqlzlFVwwowJR0hABHcQ98ygWgfx7qdCKo
E+sZShtp4/M+mbUPVF1BFPOImPUYPhHuq7mgEVlHlJtcYhwRX3CjyWkjWCCy3lUV
3hnzVbP2bMNFwiRonXtUid8+lY/BaMCapozek3vWbmWnfoXHqcFJMQKv9QZrEdKa
QzNZgFScOfuDImEqJo5//lNVYWv/e9QdBQ0yiwjl7nk5P/BM3xaqEqjM6dIhIE1N
8jcjU6MJmOguHQWnZNIKxX5W4/KCiXsdkul4gVuyGWPCcJFHsESArDf6NZYbJm+J
+yW2/NWgFHfrLaPOuFRalqqz2/zH+/kvLWfv6Ll0UX/js+WpKgo8NSqFU5VemRkD
f0xKL4Nrw/MeH8IbAw87knFmUtEpYz+pbLfMUcB3LqZ7kWVuN0dtIabo4q8sEjEH
WP/2auRknGlQwqihn2JsHlfwuQk0nduBCzRwrSajSGnReS6BRbethWAMJnsiAdyL
RT2ZjvsqQang+o64isuTI3knY04we0ntP5jZmCPThtR1CdE6haijzFteFq0/a2hc
kndAp6g5XjM2jXEfusos0NCF39staep+FQp2+ylKVM6d/Phg2J0zF5k/3/6TcCxM
Q+92J7EOIGA/igj5JloIJ9dVXGcj83LNtOv/yzZAfxoBdjg379O72pg1+I0zvBNz
AIjZd5k2CcatbvEkCXKiOyhsP0BiNoZhn7xfYNaKPF0fe3XefmpiWUSwiTvC/ggA
ptzSYpjwQNN3HDzSX1N392q/Xx6mKDK5wtVcg1rANCKPGkCuInV10nas2u4o64v4
odpqqUSkta5mHHklUq1uN8jx5o84FeqUwCZCd7AC8LBsFhOlnqpN3F/Ye+eiVoFw
JgBAD3cmqE9bPG+SxDShss/v9kKwxKETi59pU94JlekOgKYqrLw42qaQ5eNTu9IU
2ibEEo9o8sUzFX8Y40AvsDhaQXay2PjfIKxwLdvYk+X3bA83nDLmswGQk8b6eUaZ
i1rOZKO2ggEaV0AjTqc59sCSLVPz5cjNZfqcWTdE9XYy5cEjmZQWnU+Jz9ENlcfJ
n4KEq7mnsI/SOwZTdIoWJfOJbSiHppbp2UWxvj1IWj5lifS7UfLoJ9oo8aFALZ31
xe1AN6YeZ/YW/km2/by2Kvb3PbBd3sr6rTjuiV6qXR2VPjoYmuJ24IHxQqWX5saM
CirfVOpYQ+baoVlXCGaZ9xFqKYaiWDDEDqB7qRabz2LYGdjFG9Mz60PX7xKEd/9O
XNGbFCzU7HxaLMKCpWeqObC2fjPnpFHpOfhHdB8hWPgqn4Io/1URb+yRrYgKM2Sr
a7e0ewqU+y38EVTea4/T8UeO5lILhNHnE4GSBTRBlXv48e9ii7Goor6WYYBbAik6
xV8oHzymDx6/xqmYZ2zxHuH3SXw2mPg5+FNWrdM0lDhNOfyMTM35feplFq5fAL5T
psM4eWIUDLA3tTQlt7rEnrWhxhJmFEQCVeDOi50ZtgCuh4ODMrxJcrvc2zcRtWIg
kzQeRMgEAdPe2cXKuVzPrui8iuPJ33cfKtz0vMeSAh91JHLXDcEHKUXqP2M9jvTG
zazHAwvcVFnEdJ0/rnM6ckngZ09VoGRYZdM08G34ihfvHEa0QPGPEW5/v5cINr5x
mQBNDhQ1y5wzNT3avCRlsbTrI320MP/cdXRZxwchYGW8somEd3Stv85O9JjxtpEb
4H4V2d5ZgFktduVVIycByt4+8NowBgutcU+Ka1j4k7Zr7JCV0GDRsqzQIJs+e64N
R/pmA3HUfZAmr2xrpPpap9PVB+VKZEJ7N9HPl2NL0GWHuJ52//Rn5LPmyeJ+CbIy
i2gCKQm+m+yIjmWToGgj/JeZMCeDYTawb4K1yc+2x7TU2KUrO3j85kM3CXHrfGvZ
QStXMorJB8/9GxaNPxPyWQsAHUXV1ExEDEy+vat3JIR+VCk/nkOjFHusq/K50ohs
cJwwtxqMVT/klbBPhHjC+OL07YxKTM6xluELqIasSs1Cx7nRfkZVL4SXBK6YerTe
9rVJar4itjz7ZHMLHSV49WUQpBO0j5IPc4SLJRxsGN7umoGwNJkhqbTw9/8ZJsOZ
L5TGO+R8LldbbSybzP8E9SoFE9DA8lJU2RxQ8PXMBy6jSnAILgvd2L+2mO4tsLv8
dV98+hm5w4DwB4Or4cNHG7JD/MRF6hedlEOFn+XzQikCHTBXvb2zejQyCW8O0ciY
RDT4eSMguTMdtJeg4YWPPD8IsNqjvZgDlDDbByIfUp6BNNBGyB21fbtQyj8szc+v
E3Q1B/PvDpmR9H3ahnRyxls38CNzo8EjABBZzODdLN2aM96/e0UTO2Tp7b0uC3bg
CaZGM122N0jleKRW+XMOuGKvSre9uF8JESACydXnG2qGAS2CPscVDzRBk9GsIbA3
h1Cf8XwdZhYCXLj5h/ZTv8i/bGiqAsoD1+BvHKftQwamBlmBkF+V1xMlVraGGfBr
/aGGK9n8xlGf/KTHvW2E8UYK4d/Q796NBbt9ywpAOKisWkyK5/6SrsoJClLLtIBa
GGcjOTKyC8NjjuDPIrqd8viEQJgUZ7vWPI0cLulwM90M5iHej0iix7jfwwYGM25p
OKi3wBi/tymk4xwbTQh2/n/LT09GHersDouVW5ZLRyb26aTLOcVij/OaH1p33QB2
M2SsWatcAw3q03jHbG6CnTUmh2eahZJibUoFnPE+SZ7P0Kz1cFDgPH67pZVL930O
pthVR2zQP7x0T/ovBvOlGqrMv0HOpZl1AJoKPSvFfKEFzwfXxttqMSsdoYysmrC3
h2uhtpZMlLn6RG+er6xWN+DrTz5nEDSKZcr9o0PdTVx7vFNofSI83v5C7FbRWmI3
fQ+D7ngcaw+EWx4a70AeT1cZZ2QjczTDZAdQJzNmWe1wZYkvR8JrXWrshBn9+BFR
6lD0adwQ/GjKY7GzlbyPmXsO8LMGwGFj0Jv0qYvKtU3fYuwcvRVx7jAJGNkwSMr2
78aT5WyVXpVZ1GpEGOM4pvN5r5k9M52WL0uDiJeBIW9r3+ig52gbv+5BnGBJCeF0
wGoPdhGCmiu6VHLgg/hRXGCZRZgQ7WvEAAd/6Dzk80bi4rvcu5w/5ETfugXtGhqc
eZEprQjbJ9tmOHw4domDakY/2wMg27pUMEPgU/aNPYzsloAqO4M4FhbDh9qy5sV6
pXMz69rjrztYl+Rwwy/GOKyp54zu/VE5VxI9y3JydBZM/djQf8qZVi0Ylb22m4/T
CbHVCp2CwslRfJU2VfBDa2dFWQYNU/Oqygyr/foh6PxmzY3komCYNs606LNOJspn
+PCcuScjQszBDAzEYfozXWQMRFJZU5hdt4BQlTddJi7FAx98/lHZyLBVsDS2930V
V5OOUXQvjkdeMMRBMDVwOq/zYirsukieGxy3axynhGNYc+3DtjTq9S/I0Ql91CMo
UF5rDP0Z788/KrVLx/ce9+5I/gLvrHe/K64H3wK7h5dSaoiIDTnxoJWQcf9nTi5S
kLpqlKRtvJL7d3JTYYl6520pzUC8SHOe1QljcnqExpkFaJCRKScCPsMGy8cWQQoa
wyViJ8XjBjZVLaRgIQPYL2YZBE0Er9JtCk/xeloCOYyFe8vQFRNk0QBZpwgikpa1
cI2OFCMkCcLXrS+dgzZPihXzwafc4Sb+Ih796URcbTS4OdtCB45XFlGEmR1a5yeJ
DOokznX5bWlJf1swc6UwWCkTzR5jw5qZoJo053SNJDkgECepbYxojnCe4u4OxOXO
1W6/wn4jXCot9JUHnUpHpf30jv8bU5zM0QQw30hE9heDQuPvKcDj6Y921EBj/Po3
g4ZrgamuE9Q8VOTGz0xKPxEBQCp/yUxTuOU1FAsp6sNS/St1HdBJHi9Lebv9DL5j
k8RlP0x7sYDF0Tin3Dkac3cFq0R1a5c8bb7E9ibdQ1FXn6NN0HU8b36L0Ri/+Vwh
7ndNK4vOw8dS+rVED+xRscxof+QQc4Kl9Kb86Ykxzvyga6D9IT1+0gSHyFy5mVRg
xxVFT7ViIc+11/9D+qrNW18oiSuubqRN8ylpgBmecGm9EMki1hLtVDqojnKVvRNV
vmfE+zhfQgXVWLjfZINcLTLfwEQ664enBWnG0PCmQGCvJLVFVQshU/z3YKmcEtWX
KZ4WkhNgUQUXG/b+cQZ5H6Z40WUcwMotdjRvAtJ755DFySZwMG0GZVgnNwEwuqzh
KqKS9wn9xqSfxQ5LFpP1mXIf9UOpzJ+aAO6UH6ArqpqWonmCiDPo/6qw58mbIudA
T+F3miUKgGKusAYOaF/XbXu3xwQ4bY1vmLNALneJs6oc7S9SEIXqUhq4728O2Sub
vh96tfTulIxO/Eo8tu3ANMeWJlAQGGoiry4IYXXIXkzgY2yJXbvfELyU2PknctI9
gVcjB0bXtE7Vi67gGEFzVGzflF3N9kLkN3UpzfIRDtMorIJ62GJZc6a4b0mywUj/
kjhJhbprhKC3dR4Ja47/G2MS2K+i6pTe451OeX2HoiTqVE6Jx0ISUnKBv7c7cy5m
WV3uZQhfvxmj4l9InVOJMFUjRZc7izNhjlyZ36Ha64KAdHEV4KzfmrJzykJZzwd7
th9+vRFiQ/l5sIXWvFgVunfiskD6PIMpl1oZLjaypC/e2bI5ubn+DdM1aqOXnWu3
TI94t6+NXrrQasDmw1crc0+htYHEpcm+PjaFyeKiCbKOnp71+TcrRe9PuFEmu8YO
VjuK06iBkra+skgTvxV+pvRByzAoobvi2sAO75pvkeCud1xyVuEHdORhm6BrQIHa
eGdpOB+iSvecsoLLeaBca9Rp1n932W2oq/vFCecYliwrXzVQLIM2vxKuKRpn75hv
p9xSc7Ipxl3s9Rjs30oph3UX1DUWs+ctsSWCMn7Ttg1+ANSJkgAmEsqkLLlx2GKN
x+R3lRO2RIc1CMmfyyYBs1SSILNmtNTYmpM4XBG9LhoD8t2ZBjyDwnK09OFC/LeT
qyQYa8HSuueUdw9vdttiJ2Vbo/MGyxebTJWzm2Dp2Lm0UhdTYKNMEJ/u485Nz92O
VVb2SoI69o4mICUxaNrsrbPLrffDALGsly5q6QSG0UZpYMgX05Y9a5dkbZF7bjTv
WzNsUgShAmSEHPCJU9xYpbUAPOuXahCKAhOF6s8ea0n9Uj/qT8ZCr3t2PQZ4jptX
fzCeb3V5EVZeuFqqr0Of6Y5skjMltCv1KYObCdocc/YoL5PtvH+YsdezWB8jEmML
3CjQshhE31Lb4Mfmwli0ooa7EdtKaTx5Q+eXIPPLQ3OmKa16Dft7AVMCVS17WGK4
qH+lr+mvh3/QEkQr7pmbUulxXUZLGC+AXVvMhWOrvy7l0PtNUfjdOyxhJG6EBCRK
5KHsCRYT4B0elIKiymr4L7BhUEEM99FPaFj4f0JsZ+6OI55hFI1/lHK5hhcH8SSV
LRBTbYHFuan1gEMqRBfcHssbsuXO0qaTyR0oA4VTakETWHefHD//Q+F8jHKEfIk5
mCULUEH5Ej2hOALC2o6e25tDbTSHvZ4M7FLJH4FrsEgyzS/bisxUXtiH4n9oPJnN
lweBgfCh42HS4hISzgRcpWiY33q2SvVPOITIuxZ8Rb7PEz/hqXlrWtOiXDWzog0u
bkQPxqOEi7PqXACD9qR7wqWUZXKfS6pkZ5PAqTHKfK6kD5gFrs0JrHx0XbsQffkH
vbeI4BVs6gtjSBtwjV86W73y8FFzgJMjlTTK0gRalZn+M9c71uCUJp/MG1w2pAc0
UIN7uF1geHGrVW7CEoTN9NAXgTama3t768POCzXnj3IJuuD0g0Y6gCvu2oqC4bZb
NdQr5+Mvr2N6WRrgwDH8jJnXZEcVTkrHbbuzJ0DGqoFU6lmPaGy81vXJ5K36cIMp
1uIYB2FfrwCwVLjEyOEJCIGqigBRSVz7oYbEgyv7XnLvKllrSoBt6N7TF7kVZ4j/
/XRZBMOsH00+23WGsOrVhCswm0yJ02e11kgg+U2j/inrcA8SckuWcDUnFKDPAJEZ
zrbcGKn4StjtvTZpTDeZxmGmBlZ6msogwyxtoqL7UUJtmHdByOV8IHARBmP8ZNFZ
JoRSqp0KTwfR7lzUlhnLIvG40NDz8FqTsfEeVbcSw1xKerWg2pru8lzT1dBGd65z
OA6TCVDLZcKNrQViIdadL2vLySpyQBTQx9deob2x1DV6oq6zhFf0T8AAIoaTZ0uc
P+6PODSWYjqAfKbc1ezbv6He3jU0HdUEkIn5AK0Jn/JaZOVbJ5AuNvJzUgKqfixA
iucPCgpGNEyUJOKE+tQrtImjin0chIfdLxGlzhQKmUUXdUbaVxZSa2D3fn69VUMr
jCn1T1r4AaNw/2pyHEsTuZVmO2YCNk5gnw8ZEuj1vagez14mNpV7o5f/QTf/aiAu
aRuJ23vhXIpvCm+vmnljiz53wBX03NzNuwjshsmwJJ1+HIZhsy81RfpExiYXro7Q
/zB8slEXo7MR4xkvyih+LNnCGpUs1FLjyE702a8YFhuWVAot+nP1VIevivg8sPxX
/lccwtgh+jUOGbCmDula+01c0PNnkNL56FHkvHGHcN5ZtyWFdqIOQ3+pgX7gDp0G
YkwLMytWgSvy60beAEELZTSyI06hPVF2XfAkA9uxk8yNUqRDqrEPEr7Z26U9uFu9
KEKaVwDkY+SMnemC4NUI0QfBxO+I6luEF0A/qXGg3L+8xp4jIomevmQH3vHIyEjO
hnEga+VWqm5k03GPbC5cqDJx61Xpp5MQ/7uldhu1Pn0uERpoD/4WDkVAAtJzsnA2
/MWBvzJohlC5PMMXqBWtvqM8iW+6E9Fz2ivjSuOL5rRQPK/Z2vel4u7TkZcaOaN/
cNp2f4EFwC6ukcoVFdkPS3WL2gLYrV5hRlLcloSDT9JkglJvdAEQp2CzeeOBEW/Y
MUfM0lBiif/ny0SLdacsKVri/W19zMOrySUKaeWUPiH7VBaHw2hQbltCo9/xpMan
erzaRL9JbaedIYjMV8Q+nAYTjQ99n18Kwp+kPpj4pCgzsK1bW2epeh0xyCNtNhn9
TrWytzMhv+Xctxyqv1tHOXdnf6OWoWQaEAo19L/MfOFvQNycUomxVZVtza3Pa835
yWOTw9m/WV0GOPP7LUXAC6oo/yA6ihlfUHRu9xwYF5LMlSv1JMoNaZrPdg6wblN6
w6KmxcjHLh28pBsYye3yNZ63Wr33ya4cWk5B2TZVs35KQXomr09ALS2axYuJxiDu
o7q0Gp3tFgXQFpRh4nHmYEo8Z7V2a8DQBIYOtwJeWe0s5osAAKaY/jvxcxj8U0ZD
WBgvLqd3yp9KMLkif+RHUOpJaJuSciOT9u0ysG3KxFnjwKL7J5WEef3kZWWkk3o8
hHFRVk+xTujHsPP451+iNddHJDR8xeubsOFc8n3hBErsUbDFv8vGaAVxsP3zh20P
vUybtSMeIvW8ce8DIqI2vEEQdljXGDznrv8EK78ti5iJR/x/yLRkDq9rD2B7THlT
G0e+IKs3yd0vMqEMjL8sUMbC9/SpPV5qhL5vUbCpLlNQ88BKZl5BEGEsMcZ8O+Oc
8jA/yjH0THEdWB2JaHfy/UlZa+EYIzwYM0kYtog+gLSJXty2vvRBhjmIH9fSXQi1
hA9IUVeYSMrH9XIi/O/emJU7ozMeWLdMWEbDmSyTiAxXllurXqMlBuppljBs3FCZ
8I1tINA/8RNcI0esf1TFCs5uEbjpQiqkMrmowTmUMQ7ONev1UsOQRQZ4nRjXOhU7
Cmz7FbxxL5SU3J3MThUhtkrSxXXMSDKLcqaVum/xfnxARM2c76VaZMDUnO2JDgbx
UKXCTFN1CgPMa2WXPxx4I0yghtqioI2ouCStkdMYyX6ATEd1cghfIugXfHYYTCb0
cR0WM5HAQFCOJDBtO5bCp0Z0EJhNkGIr0eA+zIjF8XPatgw3C5BAH8p95XivZfS8
Vs9gkOcHoO46Kwuz9Wu3/uYgMqjK1IsRx6MRYqaeG6uSoZW4/1eRmNImZXHVBa5z
UIHAQjsPhpaPZUyPmGapXODC2Dr64+CmgFucNWFhHw9qWa4hCRLzqjL3dwtdmHGO
QGSXS3Mu0vDSkyjW6VKY+1IdklpP6t0Kh+KRnQkOz7bplmE93Y81HnfEl1E/gHYK
70JCbBXR33ApycmZ0S2ui5Bbl/mnHVOeEDWTtZN8aWPvpjobYHINiB2ked0LzSU9
LE2nhEfPeDstZ+4y2rIKMdgnM7LpDwQW9Edug9g/9zH/0tNsbOwMa2Qa7ypKNvuY
/QE9UouaS1MUam0x9RSK2hyqopuRjjNqJCKxBHe3UjXmiiyyAioYOubUV9hWXXJq
iazZB08c87M2Pm2I456Z9lUqse76I8ZRg2K205HEguHFqS+v6FoYw+ogYoS01gJM
XG4szzpMOH0v27TtS1H2WbcvsCd87A+pYprPvi1AVhxDzx1kuWhxPPTIJY4fy/Kc
FPcOxMmBYg3MPCahSp+qGfo/draG4u/1pyd/D1KR8GUmDFwH712I1z+2SvPv+pbZ
lK4uh82Jk6DT7f5BPKDnpVByVo/yJ27iI/Yg/oB/Zn4sJscolrfYeSXD2CAOM10T
1+fjCar4ad77mnq8IRWfbWapk/czqjdmxH1+qgSwpiEzsNFUasVzD4vRq9eixSNF
3m02w5B6h7LcexlzY1hD6yTZHcBNtNCs/sM5Iz9evkBvnD6rX8bs+Opztxwj+54l
4D3bMgy7IUZ8b/QzGnDVdiBfMOY8+4/1CuofD6TE6ov7A892Euvr/VP8mYcQuYYQ
++bJ+ibXUfx4/E2Ny181vtrU9zR0j29ubML20FoBUU0hMVv1GHKrTDshvyISJKZd
u470W8n2P+Nn+XM6pfZHv/R8XVDOwv0NehtPD1bf9vyKI5n3EM2fkTZLHfmF0BXt
m9nF9o0mw1FercLhrZueP0Asn/0hh4WZ9vYD5NLVDfUYR1fQ72/OsmTYLMtoLi99
WUfaMU6ldDWrZeDRzqbVQV1/fKtdZYZwKB1OEW9nfsT8hVgkZM2sgWINSI9eF6dU
TfYOZ+nxUv8UJN156kWjpzEPOA2xvNUKD/1gDhQKDPCtUirKTObY3Q1YW9fcx/IH
+jHrAbzakBFafubtHrGBcBxZ3yB/RhwF0MnzxsO99kZk+l6b6U+TmM62xNbl31U0
UW/aBn56ymPlBv7Ts3PQ+LCIVk7CJTWzEeHikfj0zCqVn5kelJxzIUtuqXdbj6OT
4aMZv+x0FGEde/kQpjlA6Ms0RTfjcNguB8DjgXniIy3tHql3CkO9lUfq21VC6Br0
nvcJ0nHlehpHYs8nWHbBgTpPq7focFb7Wr1lk7YSi+mr6g/duxIk9mSGunB7LAl7
ncdoIE/cpi4Z12RnifIq0sd7n0NfhrBa1tiMiI+GIhGMSN5fXZJJoXdEVBY9DgDM
YHtfove0bKbeYTXUrZRxJ/rdVaoRbE/H4lA5puioS527MAtrLTbR4I+gPKSshbJg
An+JYixVDL0EHAWkNTv8w0ur63z1qPia6tdvsZNao62cZHFDEB4vOz7ruBMmo+BA
Zg/UaGSl88Jr/UOCIqZ/CywWcPixYJIPzsraEInrolDrqldOqJK6B+lDyvwgBLlM
G/vvx6aTIniqbzAIJZMmq9wsT2+6EdiQ8Kbf870aUp9NyrrieD23zTaLcsrq0q06
yUjE1x0djGQfC2zNdHjxY1ghblIiITlmtkcpJdhoZM7D+IQ1kQO7/YwwnZx4DyBw
QuVTycmsB+T85OcIFGRySE9xyYhfQ+uUkdNKfKMy5VPa5CwRt7+sFlZBy6lQJFu5
0xJKlCZkS1skq36KIYH0JQVI9K1xzfEBe+CUM1R4Y80Myx54zs/ksPVLnDi8236g
FoxrRONeLqOGGEaRVUKeecKCyhLi/86mCnVHyxB/YEy9j9wGUXqvILVSxvywoOle
bPYnBDs5qvk9KeFW8CjGqtYZ5T8r8/ZQk0PYYqmsoqC4yo0WeeRM9741ORaF69Db
5jrWENLBGM9/QOPOylMMZJCAf3EMDHyYMuJeak1DyG26MadCvUpIJpF/4Lj2iQNQ
7aHwnbXCReuEzvMZ6Hz6XU8VhUVQaDZi+w1e+ynPiMayTsvZpfkDVQizoWtTqZ62
zDW9itK3CdaAhbinSC1V/048TJkn9FX88G+0wT9R+IPVGO/lCZkRWS7xHhmw9QGA
f7g+WEPByW9Znxr3dk905p9mQiIDw54hyjnFHIpCS2LC4qIWVpp6jWOyNjb6ONHV
qHHsZ7R5rx7mWCEpJqsQuSeZbylbbmoDUyCdqeidWIdCCoURBGNCfgpBfZDD4Hp2
snN7WmlQcE95Xg773mS/GOYO2MGsVrX4kI1GJaHmPO8LVhaKF+3bYuLntNwypYz6
M76CKcYcWIVB0XDhiOK1ngAZMeC8j6IGlY4u+Ue0vnsFZVuN0+WvsTZ8jbpnRnxa
WqvMCr0wo65i+xVKFO8O/U+T5W9ckMtHmFfoeWIYDa0MVfuRuJN3EFdTFUbvpXhx
BhS2MMGjb0sXvu7/jnzh7C2rokve8IQiiWR8CK3/TNiH5MH40bNNrFAn9UvTPJn6
dQjgUobrpPw0KZFGIZt7M7rlQ6dudbQVovMKRdlXc9/mQS9PvqO9fb31HsBqv6C1
8wSMvOHEwoXIBpCb3aEWqsHX6hGueXKPSZAAUUPihYs7XtWVORQIpoB8TpjcTmwd
tH90EwnzBXPRPVus8PfVYOBQMyEDKzOQaRTCuvjSj726kEXLjHgfTlk5GKPe+Ame
Bb+TGHID/sqWZYcHLj+vtsdzST6lrgVfLBesgGeV1pUYCz7KFgJD+gaceEsAgJC1
D5BU/oh8fnuaL+bRl+H8J0+MgjzT/A5vLYstffCfHgzFNX1PNVCfcfnpk/TtDCvC
ryNCrVTwlZAfY+1wzv4ScspCF+KSwgvch2m2PnJjl+BJFbJvK6xnhZBHQbpDhT7y
q9fgcjpQP0xOOnZV6ldawqpTBAih/NZ+W4/chz1PCnYs0BIobQOxvPzDNdywOyrg
9zWgyy8/TLBuKWSlITm8aWw/BnZnRJ37BbaU7X25wo6u6OM1XfDFDlJk+DGHhaHl
NSvs5GZcKEgkEEdDxgq6VrBCYrkjZLalKo24riETNP1WwWKJxB8UT0BuTiq7cLcb
f5WIy5T38zxfXaOkOAJfJE0gv5M0SSgYbROCcH1tUOTUcKHDiJAxuBc2OCstciHy
gck1gWZV90AzcxVqZNbRL0jKrSk9wOvNJaUuXLnzGqF8klNtztSmFFnEyJSFJwFj
U9+8lkjobNt1iKJyG4K0hIAixAJfVIVNhzJqOfmzbHw0CpgYq5fNtW9/pVbK3L4w
+pbNrPXytjQubCCVGGjMat/j/36HuzY0qe3JSlyvFdvhD1ci0PkPKsz2PrdASdTF
NdiPeYUSoC8OYl3WN9wmsNtn5vedG4b1HLSHZaIJ1OjfYBvbiLpRJSgRKwekMUuB
1zNhppgVUsV5CyzQB5AcnbCrUPcNaZzhyjoFPbeT/KLxF6K6HhQ47M3rh05lVMEF
8VjzUNYd+cfed5IbqUi3oWqc+yWj9fEigsiNsxzjJhokQZu5eNnsidd+urMHnlz1
TRzIvHc0ek/Tlrhm0CeicJGRuJpcAxWKq5QAhvWiVNurcwa8gOg3jS58qu4nMRe2
vszFX19JH7jPPv/4yFx06koPJRfxapOcijwqdiuT+jiwNLU8XLGnKO359uNnAfN5
o/fkn+yQTgOxzhys01K7hJK89GM+1+wTHY8kBYZCcG6lVawp/wa9F/RMb4XcH9Nl
HcgNtI+gSVasG/gnhpf7BtSN0WLy9z1YyJVUtcE/WQ01xHZaoWRc84xr/LI0muZj
N9msVNt0y6B9gGItK4YTujuBd1q6vRje+grsO9nV0ulK6MM5pOfQavjgROElPRFd
pv/MkF8BMuqP3Nr8UrXF7tOWjgoyZGgWbodNfdJJonwPOT9bi86OTPp4u3iP4Lpk
AR/6rhID8Mrhx2c2E8BpkMYkSTM+o1ugIRuNRGY0Ya3nHJ57zdRxrD4vLqlkfrjJ
u/6eAYckKSyMWa6KNIPlvHeOsfAXqe7ckBPj3A66pOgwFVvEXmFiztJlcv/FQ0nB
GaAvkdpmOzRszoBL9l0IsrO86RQL0WHbf0+TcFFvYgoWoG9NrZGtp5MH4NjNcLXo
SSBTMoG/Yb/u62eXXaK5/aNYqEEA7IMsTlQqc0S9vCwqjw5mGXm62Fd2ERHzVVEN
R4On6tNa+IP0g+j2gHQHupnqxcnuIjSUOpHfaFHBB/oypVD2inY1f3dYXJir6mu2
xtigpBPK+S+iVjUpUhOMr3A0FCNVCs1IUz7gV+4sfpOwzoxz6/aI6C1F174h6X7e
ejwSiXxXCYkvuh5fnrBXJk7vbZpZok/sHZoFHTiNcib//wBcZlti+6TgkFqoG8AH
ePLXfWuhkPoZmGkUCrTZ3PDuRfAKreciU40ONFPqTBjF5GeqPl3y2fHffpJuqiYq
ppCi7sFSOaVdnGC6f96l64dDk2rW1hO8MT1NPhlL7nWcgxRxBYf6oTKjhqAF9e7Z
Hs7HW5rvfO/FzmhSMb3U4AOkufPQlRJSNY2ytDO5U2xYgtKlxTlQYUGO+oeILbGS
wBMFX9Ud3H5y+5McmlbLWf9LegUfBS9WfXSXXYbH3RgT1/HU+Mv7t4y8Q8EB3Pdj
mqMrEvpSIEqJA5GPkkoG/9lHzL7MrchonqlYyFgX6eTKYSODNjQXnKiTm46uauG8
h5yrG5Y3SqpqKUr2vEy0ZLfjl/9O0wrNI3Co1s8bsss9wa4EOtSNtEp8KjmzOkdx
rph4wQtvwgG2bpns/rqSiDyALsT/GSsoWGnggaWvv9T0HKtuaMAfN7Iuolg10NIz
tBBHDzOnhqFV/8cmRn0XpmqofG7F1SSzLv2IgL5e8uW68ZOdtSRyNcZ++0tk9i4j
T68Ft4xtkmBH06rEIx9FezSu30RpiYX5jLMsDeXubnwH1SDS980JghGB7h2C/TzJ
7cnbjDhPHeGE9NTBgZ813AprokwaA/3w/FRYSzPAXleM02XPszxzxFo503cwBmg5
PQ50j+p6cdcHR24CXG81R4G1O5ZTJLyAcos4vVZMV5CYwCIzxkoOSclBZ+stAe8P
QLmF5PndNajysCNkclAo80QEPNiio46cGUvL37Ir9zGqnetiG1bfJat1gapEN9UT
Cfd5kNsQrGi9s+yt0LE/jf0cdd1E4KODXWNyGnLgPSJw4mqGW2KHd/z7kdFdRJVQ
fOHL1wjbo/DV00a9XaE4TjvPZP20sgdcW0cGE4dQwHfsK/uT/KOnsyE7S7Y3lELx
VMCrcNiYN8syeWpEdgTLqQFlYKjdysQWrLcp73C8x85sgwLv9d3MlKTcg05/syda
PwuXve4OBg2yes7ExoGHkLOgdfG4V7RWlg2tpAjcMhN/vHsU4eD40JsNBEZ6hhMx
52Z8Ypu7BrYQ6JHwUqpCyZKe9afw7jamNwQMoeEkiCp6qmMEeaDggOsNd6PVPS4t
6jE4E5bWyrMY5SN0g64HCRCZafXsnT05zAxIMe9+TuoceQYIZdj7MKpQ7QBByO/g
0fgKa9G007VOb7rk1IQm5SU0ifJMUjT7x0YHsG7mU+l02ros3xKl1O6TMIryv8+1
isUmkqjOBpz3nrSRrQGln24MLKBI+XJuekgrpYAi543/qV7u0WhRmCOEeWekfHZf
K0la3VVNpYaT1EXoU1p4WFooh8Q2pBHxlHpbZnAbwFQLR1KDlfnPEwAodwteVY84
kDOfu1ZUA4etbSQjAvP0+viH1Rf+rJQ43f+AJGeMGz6+c5LfirnobPR0lDGL8aPV
/hRbBmefAHd5X8siAvxd5IL/hEiZ1nsnL0m4/ojhL6vfEYnpYXyA/Kqzcl3hhOoO
I3kdJ+wMs3KRXzqMtVSDeAWDxEfUZWLRp/1NA271txJwMqM2ydPMZPPq0tS4Ad4r
/HbzWdZeTY3OHTMFaUy1c77Q2W+h0rNzE/a288lUQIIxf0ErCcTufuo51dk5zTjA
fNRKsFrHRS7Yo/Icrq6jLbHf6yBqjo8ZlUyLehY1xYpohz9cku7+LS4Gjzf5KQls
yb7o3QDqai9KdRcf0wqjq+UVwNg2n36GaksVTGCgjuep6C1vSkxM40A3MN/XUVOl
jp0aBiKkkMHSF0VmDprXFV9MIzH1zbicWL5DQCK2XE0mhbNLqeEByRkrn76fm0DZ
lI5OwmS4t2w4yAQNAHngwpWgynK7zJF3oblmaf08oORo7rKMDSVgRNC1A/dEk1Iz
JXUk7baMyIoMDAQPKinyR0Nq/xY8D2j7+pYJDqmDu2Gklf9RmKGAgl/KionglZ01
NRd5ycqsSxeoLOdlLRBAaf/wwQKKavvhSOJuf0aoIfdDyNvB32pYPANErp1CSZPV
HoqYbeAcCqvmqGsJ/KSu0GFILOnaCJHntzE1nIMxC+1+P/9+M7hxCgih+0FYqsBg
ZyBVRi6ZMkVq7v6EDApZf10X8GTCy7Stj9QBT2NJrHA6BsKXGPvCv7j+g97VJ0a2
XOY/WLv6ccxcBl8OlwIoSgWIrIw8nRiXI3I7zdDvsai3s6c/kLc8GMaVqX9rVxA9
ZMT40XzEl6loCmMqXndlcjDhI0QBJ/thqpObE9xluLfY6br2vaRDyFOJLBD4lvp0
m7dH2mUPWzSw2mkcAew9ts0gVqeeDXn2uRKzSEcnbnEUTXCCRMuHvdTyR9BcB3SO
FGbQmekkYM5amzDek+xDOT3SaDNBwdp+KY+hd0PzBMSVSuF0WNXcS1i1YBnc2CO1
yZx0BeWjNIaQE8XE0i567TyL7NLTDBJrQKll0n5WVQdUVvbXY5oCu6nOJ+xjoY6u
7ZTa+VrUb3FEhM/v0FuSSeMPTduz+Z8UajMnJVr3lKbtCLevoa2hsj4mDw+KTXd3
oMx7UBJ8yWRd10we16H1ZlFEMdAWAL/gHPZDqlc5MYdS5ub9/PLnpBhuGbTWL/Cj
r2J+P0jpNakLRzYign/GDCBW5DcnNfrQstBijXuWeIK7a9UlcqWTBX2Oue2OOAqN
zNGsFLYESDLUxF6CstL3uvT+qEDr1iX4qXAzZgIr9rGYewc1z4BBbEKV3wu1IefL
JQR/ki7LOt9+eV5c4irSJczqkT7a3hvil6qdsOucELfxvAAwd7wRVj+sje7tAxMo
W1bEjKzDEWouB/w1UWtFbyuNa09T+mK7EG5/eO6gXJDI+pLv3oIavn7Yy3eW7nfl
0vpKH2QQ3NzXodjCKwjeTVtig8qtF2AB+Ex7/adaAWq/yZI68nSMIn3g29yTgZAN
T3IeSXr3HmDE1dapSAfWQmfislE+ETEWHTKLqa59iFOYqKK3kTIUiwmI/O5FZoiM
WsVBgEy0e5xreq2IjVv07uCaBgnALMD8t24XSMZBpYvX7K2ZFp1cSv0fhy0DMwfz
GOHRB/PjBenO+9xi2RIgbYs+jJ7gArmGmyY9da+pB8Oj7chy6yIlklciIwAFgQYd
KZllkh1rs+zx+e/klFVywr1cUpl1D8FRPNV4y8qx/nDKjyND2qLs5SHtN17z7SgY
kVdmuSZ/w+LOSRshU/gobvKMu/tLOoxtU2FeRVSM6tRfj2ur2JvsFw8tWESeaWup
wu1iBYPk7+Pw9a3D5/PBg9+6y9grDRhTyFCZDaD4a+mUlh+4qrYmZWl99FDFq7sL
RuUJgwlVjjVnMzqaGGiVT8Pj2qxbWGElMenu75xHSi/ka/PfGsS4IN+PIH8E4wsu
Ncs0sH2YRFpxcDQXduo13EEFCE8kgt4IJVWhP3Ig7MA92DOwv56eLSbN3kBW5Esq
WJ2JxTZlbC/MtnWQv23Ijushev2vfjrXs6WFv+mpOk3tmIjRplfQrgYLcNv8VyIr
eWbYNqEgR7qc7igd2VkBWpHgH+Mg5S0LDTPbQGDEYUiqlqmDzWKEMCfGW3WEQliW
MnFSHgpiQHp5Cujn2LzNYZsWeOYkmjzrvGin3A1GMFDz/U1ahQJfSe3GJlNptCSc
jtxckoMAMSfdQAu9pXxZl6YrYDWrdRtwntDiIxrkmTP3ZZ3XKRVNOH6Ay+xFHbEn
qIP5Q3BBLO9avasKGPTm0HGMDubqFb0H9OnQCLcJQDb79/vqzmjPWSW6m7VcsZx8
Drb3n3F4wTnjW83YZmXxZvRxIKjLBcVj4yGMNfTRnjHVP6IUccn6RRkDkfwcYj5l
QH7yFfX5HOHPbejMK/UXo9L6jVRC6x4OwiRIQfRYPK0y9cqVtdsyNFvcn4XCwCkf
Njk5/yQsmgyqIbvJLH3BT5HpgLxHqC9l6fiIj8gSXI4qAewC1AS+KTdl9+HYcI37
xNRhoBBA4KO7Z/Pdm4RKCKlALs4c5tE27eUaMH4TqLxxHxP9TwG/EqFcKgiu2ejI
G2rvU+hWfyHflSZtmzULKErQmS+rjb3C+n5BqWjlvb8sts3/y3/MFxkNTsO00nLQ
tojrDp5ujc8INXzUrpTnR4/ewa/kf5Fsfe+n0BqWf2MiXMiYX5PECCGQenKAcro9
EpLBUBACfcZGHYbhfz5pqnJ8+a2F4Sk5Kcj0y0wP/n8EoRt2Bo8+IeVPKMRk7MUO
6mVcwLFqnVdD/ChK0v/CszmjVnJ+k53s8+lNGwJyEhC4ips5bh/cTLtZXhjgXplL
wbJKPQqO8SeVSIKvmE8K+UI4L/hN7NgpN4Ukg7+Z2yVzw3T0hx7IxNoa6UQjL2/S
EAVpRW2SCRQ8NI53H57pP05leJKctjCAt+FrUYzfBq+WyNyQKdbYT9jVq1nBdI1G
j2y2dBlRNgdjp78JPCDJs7zWFcFCH0YMPCJFtcEapRWU2IbZRC/LNg7+M0203yuV
jPtDxAYSCjaW+GoJtKqrzApmHJDsLQdD6+8l4CpclU3N9AGXsWiJytt7qDn0ZKjr
8hnGF9R75+UzKW4H+Vg87N85nkPY3IjBb/rT86z2UaTx79UHPKLZ+j5ZoBFWCc3O
Xd69u7EajHNFpcvYEKF1+raVkkskeNhkMypeqwkvwICe2Jxws3Z7C3BbDQcRJxch
7xHE3nqsguOTGjegpUcRxulX13KmrcdJauLqze7CFtoF8ZCOrMc0/EhbvNpddM/8
tKLO2WHysBG06gqWQv96H0pmwabgG8Je5tcoEVOu/mYNfvEe1dpVsUmC8kZvlVAL
cMcT9KO6Wz9LI2KhsNG5yxT4BAt2D6u64rWe5ynygRK0x/81Lbxa/x3jCvXptFp0
Hocx+zISvkmigW6ms+0PG5+ap5dpWMDuIEhMvzuiBBldz+qGeFSFYtjIF6ch16/Y
z5FZuL7dDmrhUrGT75VScZpwA2D4de/B45DFEQGZSsJro9KqB64q9a58lugySuad
JnFmS6D7Nq35lV43FNKEBLTZu3dJA3d9A3X3PJGrXRzOPK4/RAqpOQ2DGkZOgXMZ
I58W22ajOi09TAoatVX95Xh5mqn9SyfCDBEHKNDXf4WgMzu8X/ZXCx+V3iY7dxzK
lKrYSLfuDflnjS8JID4vL6lKQiqvLcnwAAePUCd4Uz8zhCeuPqOxt9x5iRSJf/c5
wrLn7fXvkYak7ON1iI+DjZ6Sr92m+68Du68CbBPGb207qA82RVOgRvW6qb+WyEsC
akKnE0QvVl++wt6M5YKAnEiAa9BFwjD/Qdsz0iE71PPjWBWTgMWILLcS+aT0Jot3
HzNzEBL2cqBPiFlsftlqE+nq5f85wuy9g9VcagLfA7e2uLuWDTaj5I8smeAz7OWU
My4jLPsDvLM/tzCHa2NGYXLLKhw1yLutZ8UjRn1bZTR2pquHA4DoFabURX1vGrxG
Jmuh1x96WSsFXYc+b0hobADpBmb9e+K7ZEKukqveDL1uLVUP5XQL+8izBZRhPgf2
h13HKf8pXKHN3PsAVtzMHAzReNpB14rm/Fy7dOPzvp9B1LG9vEwKcM8oLoSHSNpz
zowxRGhIj2El+3eMDKwa99MmsiUIAqLsGhkJMSKPEmDJ7vHsdvyngBHRBizE/EIG
h+p+z5OWL5JEpRJjvV2k1M6mf9G924mPcQZJP1TDn2dTkd9Vs/zO/IT2f06u9/gQ
G2hqJu9ERxTu+63BuLDvAUJLCFITiHo6qgcuqY0Nx+mEQTEBbkCNSTp6GApWYTU8
Uv/3mv0atlE5YuYZ+gyTtT1j/rsCFCUT57w46d4cHE6uYeiaoDVi7ORZsQKptCi6
nfq1f+dUq3UZlyF6uPUVSbs4dJhHfM4Xy6tVPt9VS3uvMYYy3Jz/zGIdWT6p5QmD
zoqKNcESs/BGDMib1eM0Q5BNw3YlmDXhJerl2xOtmvgFSDlYC5AkM+egbry/LNzm
MSnGy+9jWYbFehVQolNJQGq5NSRRbTgzQf+BdquYB7BSgqsCBgVVXJoZmdCgtR9O
ioHY/rceQctKouCtPOi0OuUHwn549rOAG60ducpKqRDNg4gvXfGK+4LrBzc+oIwW
hQVXoGha3coVfAwlhVuguH9q8sSjfVsNQKIwfZRK3Lk8Jjt8lHEyM+VEupf6F6Ga
MlCeXAPH5z7Wajfo/HgOSa0xfgGZlMz7tUqPo+aLH4r48kkbjkaZ+eEAsOxiMHO5
zWkh8eFEMk87f4yHfEAEeKf4qXzXGJK06JkhlXPxPGPOfwsRBOTh4gczBOh7G+fD
CHj26K4JvfpFnERMLpURVwGJdWBERZo3h+tx1YOkDHp51Fhgnob0JFD0NVAz1j9s
7S4so7ANK85IoSPxmdtyFr6RuLJpweRWlwtv2f6v4Mj0L8zV6oEejIwxP73R/GJr
EZk5uFFxSD3DNpq5bseGsQkh5j4CXm8uvrZ89x/w7au35Dcntc8FQHPlpM86iJWq
fAYJEQAGD0cMgmog8TjJUCiq7Q0b90MtnKmmveWt0jBULl3o0e9YZ9CsXcquIHmn
AKNEJ+XWa7xfTgI+BaMqxvbDUgKcg1JMs0z207g4np4aUMMSg/H60edNfpq+x9k3
W7S03ojG0qAeOsGBFKL3urT/VE3fSStmoiLYDdiyJmxufcFAJq6sCLzJI4aRuEQi
kaycFlWn1riXvpERvWg7KxVrE83AdLndxNBLjkuVnYun4QeRWGlsW7j3QkaVnLJS
8KBaM8uTGiZwahRLjAlWVhZfDQONqqp2Dqws/TUoNAmdA0sRDiKxa14qEgaqUtLq
XrqmKIQ1YGvU0hY+ODFJC60jc9yJ16XU/WEIrEdklU7cz1+GiSPzz1j2bKx0evLb
Xpgea5BQUQv/+VcbnSgElB+Tb/JiS1MoNr7TU2UOYMRxrjnbg9uMG2XjqBqeCBix
ZzICJBOQAgPpuZBv4y65yWO7jWLGYIY+mt7vqwhPnTrdx/V2ioYcMVdL1ua6vuzg
a0IfRYkuAEvYmE57Jef4kpUOAUwXVoa1dAZ5MDhMbPpaHm+dQwyXlcU/Y1IJMp6f
7TzGyVK41u949fnL0kKBAf7BRz4iy4TqPWdy6oP2FhETSZHDFQ90slwTxRz6c85D
/50RElTzdvuBuwW2aRCK1pu8kXyKef7Rm0EbTaLc1T9kODnKi/Fy17MaYz4cp3if
AJgQZiPKWM51gZaxdaueuWI7IkHDMoFL9GNmLFn9llMD5YVrcVYsdmYZZZbFpNMT
jg3DSAwstU2MpaNRX9dvPbjcpStNWMELAZcL527WDSel/rAhVLIZCOzCLJ+q8lAh
jB3QC2WU2EvzZZsOY2gQVOTguGHRi0AvsjuMOzXKYv0KTUkx5ZlwqiqSNXDEfHAD
zN1P2M9Yo7e/yCX6SDtiZCiJKGTvwmnfZQ5WXAqBNKNKTjgq3GV1Q8n1xtZlLLqs
Ki4jMdpp+hhqptAGGEZHAWeUa56d41OVapnhpn6ESHQiZt+1FPuqyNNKBx8HppeZ
JayLBFvOMphcFmfaavVlgdrQZSNEi8IDR6QFu9UiAPR0kMyBouEMcIDjMmZUOYqr
7Db7J3pKWBB/F8JT71rIx8EZ6obd6L5HTruwlVg9bJC29Vrcoa5KI7EFDZ1pqjCg
rFFwugy4oTwnkCYEQqspzh1azMdTPz5m4MmEF33plAL245QfKA1uRR/LXpHw6lYU
Y3TY3P/zjXHLIHhJFoQaz2dPRGOSxPSbmMmn6TdQk2Agso2owf6syY1xodTJ3ePZ
vkq3g9/Lj6+EAYJ0Tg51ha/srrrVVjI7WM309UT7CW7mrj2W7jY7RaltmGtXW0q5
JTTBAZ7EGPCCzc2NQKZ4NAiVjTjqUZe9E2NW/XsBt+OA/D51lObWRiMJZkjQMP22
2+dtt529J7Vuvr7CyGKng79oLhGBTJzEHaqPYOkbvLKFcm9QVYRXSW3ry8KUy8XK
FY6eJv34JMTxJnwwa9oh6yHzGCpLyPEKq0J5Lby0xHDVl8GmuaruPLX5KXsQvio6
RHKcyxMqVoP1Q+X+0G4fAjUhV+kM34I4ty6ChezHmAUvMqj/1rKqagyUa9nErFZm
BZ0xj7Uf0GZ3GrJjg6NfdesD/zGxfnD1QbgrrcXNAq2g9VGYKbpFzdgsFMg8O1Qf
WoJQthCDo3soHhnXLfJXuHwT+H3Ok5DlmGUNnhqTU7+5p/ITN25HRocDyQRowhM8
hAYICFhEBjV+uSYNVUb1GCe+sIi2ZBF1kmGXpqE5idnmscQYINqjA/zW9B33E+Rh
zKKY8L7tAVhLpGrziDBY6rbTx5iOmyDSBo0TT7z6fJySO339GByGLKJaYCWD11m8
QOmX7skQ3ZVwo6zoLJvlUQE2q8zoXs50jupfMXsxniNo7fV6qLTHZH8EYb53o9Um
pVzxbC5xCsLCBWnLaZx3lkuEdQrKpllhseqLTf6uiM8lZBSs64pGt4OTpIbIRI5X
VHmC6PuR0hMwCtwRe2A0vUCg+unId63QTfLgtfX0gVWYKWcBN2axUauIuwnEMUaj
k2MLjDpQ+pxOrAdDPfzU4RDFmbYpYY98KB3l679lsJclXUZMCv1WsYdUf5KPGsyD
fyOahw0CqNxk659FvRcONBlM8Q4Z4WP+qODsvK+N6WR10NX8tYWniqmg8LQZkbfZ
aO7og14B0MWQQDNAbW2/gQJiRSHI4vuW3t57XKTpjHtzCedEEcJaKl5yRGf2ZkiB
4yoMD8dY7Ev2BYSusEcxYgVJdWwUVhDBfm1YjlCPzFwGx5P9uTg8Z9wxTbl+gHGr
Yznnhh1sR6mZMWCO2JNRp8qDTuRoO8ZLA8SMCHEnqtTWttdUYLYd87zf3udb2DpK
DXRDW34dJ9GCJQsFLQOtXG2gRIjMkyIDf0uqaAj1S2vv3/wUZVX750ozM1lYJCv3
hF+PDZJIuMoiZTmGdV7GAngbq/NcE3DziLmKFo5LEomTh5o1GpvgI8jGDWXLlx5W
M8H3rHlOmiA2pJTJVK4Re5QhLQROnkY8iJCERnruJbnBut3D1mry3tIlESaLktwX
g/hpw9ZLsQMlxMkTjiFg5NiFdfX9c1KFnVWzqtHtACw/z48XaObelZAyxWjiiT04
C5kc5W/yfOqq67cGvBCqKhaKbYuJ1VZL1EbF3UiSv2RfWignsfQWsJQII/5rwx6J
/X/2QCs5Zp8Bzx13wIz40MwGseEE25vi+yT9cqZ5Di9zPCf0zVkx6j0C1otO6zNp
tQtIYQsKhA6Wvo01NpGMMfNAbZBSBEO0y8VP5hJ7Ao3IJhFQ2WvD0yn3cjnY1NCS
8gPUkJpx28pInWhycuv3h2HxLwgNibtLKab6iFniLqBwCQxe/rbSDmahe3yoHMFZ
xwPX3Aab0Azfpk6SUNKERmQtHsqY466pbB3pdHYH9D7MCPZKeXuiTU3jBe1A8VHD
PcbpyhcsBG4XsgpJJhMqWIApeZSzilKjmCwdAVRY/VafL4KSB/GkH84sYBgHXtW7
MGEvTmrqe4N304uCZ24ZpP+hQrVUN8Ng6UgCSRgpBQLHUYm83JKVPpW8vk0+n3G9
QA9xNRlvwouBAOpKYOYrJdH4ascN4zMstmp/28EZ8Ius+vg4HbS3tOaRu8ty25Ft
12LQr0go6c39G5y9Oz0UsazcxWKWZYhFuFeZq3OvI/El7YLTPi09M4aJ4NXOV4bh
Me+uBvPqmHWiXBl2M5zg9XarGhpAD0XfFffBFUZwH55nbX0D4wxH0oWiT9FdDtHX
uCEoLw2io4wnjD+IDZAJZ7JfEPSiGly0OPMvIgE6lE4UzVQXrvdqS3hDACqsCT/D
fSHSV3V0/ZC/06MKXreQmT4SF5gQgJmU9OrBMQBX+R5ld7zgRPc0fOrhkO3VK72+
zLgnzp/W5KhJvHBpLcchL1wFUaGVwxWZCgCuCBiJawcnEm4YymenBidtIhW9Nghl
zJCsJtuVnHbTcOtNixAhUH/YxfkAN2puerc6E6HvmTKAxZ6QrD1KOLAcdiLBHdEz
yaVNXdW+4vDoLnkwWp8PhYcggzKWpKhNnotfzHOQicHbMGm/9oXnQkAjt7RsUv4n
U5E3/YcI+YU8Grgzi8Y/TVVXazEP7i4d//vcgaQ7SxpUQYfgS+czLvI0fKWkOSiP
Ew9ry9WtYu1a9ayiAgzXf0i0I0/ZsmGixlkxwMS51r+CblV9BnmdipNHiIdL/wyi
bLR3QSanvXCpTT6VCLzGSzT3IXII26WfZg3MKUAstekEMYpu/WjiWmPDOJHeL9ob
KwlDvouk8/W+gmGKtY28RaTrnEDPCJOi6J7YV5UoVmes4IIYX/EO33db1lnM7Joo
r3DYpjpMz4NKU6qU1fFRRJmRHTFDfZgcxpwvbLpHKlqORUOZneysllmBrOFgmwIv
qGQIyfUBMzpJSaRyuq7ZUh6TU2OeTj48ohVMoH8mg/xmSUvBK1jy+7pmQRp1MUWg
Y3cjtZDJ2jrm+somX+DFjkTb1uO7JVALvFTo0QkzYm0+n2YKRSvBbqQBbOGE/2o4
jRmOnZ95NFKYvFVwlGq+a/QQ/+xO7UP29q2dsxSjtJSA2aekyMIP/LgDumWKv/Qu
tTajrFXkjJwXOmqZJv6c9trk5KVpHz93rFvGHTGrI1QOi3fg69JD3FNhXl3dwYy2
/Hytv3WJhwZpOQI8IdH/O7bmgJj34gbU9QFCoSX4+rZfWKG3vZIfWnTX+Z2mmHnn
ZltvLXyF7kie2awPfhXj0zJhL76tp6XyZi3tDZnL90hEmbbIBvr3nWUUKJTeUD/+
vUdd4zAoGcm2lAAtPuOyk3prgAXS3Pj4EtmLsf2PP2Sgu0novzgGqGStOmgI67cU
qkKHEmflLa+Ew2jQZYy3p+00B8U6OukYxmiryHxI8BgCrA6gmIGGX45dPp825sTh
e2IfeljKyp05gaoC5+eYTteMicrf7wnhZDz01HN900NEhDRk7tNal0NQxqDZNPtV
VQrlG8tKoo59ZNcgRoY3s5W+EQrjjFyU1bSza6QZdbZ6LUWWoHBdRivmAA/A/bgn
DRKcNV9K1MWGJL5JQJoMbzigW60uTNwWqqfqwMxDH8VGLEJK/DZSSYhTX+k9Vda+
TillEBA9rkxGRax8uovEzQvoGToPWTPknooEQcHggAYHAGGGPSEa0jcM4X2S/3d/
rPgvaQN6Mo5p0trFKaodYik4CZBBYfugbfUbGrRUctsjhnZZUXmyz9pgBGmYy2h4
NaWE5IDjsZ2/l2z1JfQ9b2P9bMBq6FCNDfuaRv9Tz1bOCWgrGB6plt6IWrbMU7ke
4KiBcErFvCNNDI9gPV5ZrakVkgI/09FAxhkIDTjA+horOOocsdqteKIp6w1Bmjvh
Q3SeNmDaOECYCFn58RJRp/y9n5lfqXNexgxylArG91q9ae9FyyCh6eZ68I0w0D4w
EMGVtKPktDKU6eQhTxNCxPdVrwKKf2WYT3nzRkMlOBHXUNB9lRusNvzQ+jm1xo/q
RFA7Lu+t+9ST64tFne4Gur+beDh4QW0eHIkUaQsShjh3/+3RCkh6uICFpthbo16M
97yXyyD6nON9xEJswLIWZE/adS8j0fqc4Qtpsxc5U5DYDk2DsI6DyP2DZi8r1rcN
O+w/CEQRiouIEnpAx01pizHzzqBmGZN3YL8KnHqB2KvQ3in5AuIMnGgPJzjYKbzu
ED2pnsMd/hCUS5WKYcGBdVFeBQOl1Nc+gHNVwmULKmmUfe63+mdsVBImbq1gv6kU
IbfKSKmGCioOcjZ8cgBmq+xt9XOaq3Nh+4Fj62J5oPfVTNdYbbpWhwsZuOx9j8jO
o1veJ1xlznRWaMjZemKw7tozple/OMdvwWO8qLy/uyCu1wuJN0zgCFsc8o0E7Kuk
cAnNjj8JNFgJHzRn7E7BjGtN2owUxF89h0qpWEbEs/wvsQrySpx34+NCfDelcLw/
MfJMEFq1ZQ0u/R0APqOdF2XcAQI1UPb9HAbomT00N5OzNUclmelvh2uznb4D93jf
VOdVow3ochGXXQh0YI1T8ANOJDqwQM6GJozTgJwjoBQgNdbwLB/J8Yj4Q1r4fq3U
VstD1HDRBf3gpubLzoJPxcrC90SELanEDWk64txTS96ZL5gmKS+84Kvy0ziVjdT6
CB/gDBn8FgER7LRcwKoqvva5ECtqVemS1G163Sphh/427x/mNy71fUtLrCJXBcvQ
CnJHjOiAkyCqvfKLXhdzjfBOtSWdDb7bTSE+6/SF0n+X8A4fmexLauSbAzfF9saH
Jfj2mMGAaI5EGam/vFcz9dtXIwKRW8LYEISiLm/YI/j/p7AuBOYdhrIvaVoi6QJ+
uv0kRZLvdtWl7YGCdjlgwUmfDPnjWBN/tJp57/G+JjJu1RxvgEQqw9oz1AlEmh1S
a3VB+2k6XTJTCVYUevXt+SNl1eb5SDifcSfo6zcVxF1aO/UBVKMt3Ik3ni0ADgfM
BpfdjS27Sc0Q7ynRThGGahB1G9HA2nYOAYjpUz4CJLbfxRAMRiBoQBSo4RJZIKXh
q+KkXscoiqCNL3GeGnHYnB/kS3hb7I+J6Nl3yl39LtxS+SI7H7rK1/hmFodiizmH
KOnAK/yyDmvYVuqEaOp2POCA4SEdWduwdGd1uwMAM3Mcos4lwD811rVR+08bcZmO
aR5fVfB/sHxhpqqUeq9lr3Bn8NXDQ2XRK7Pp1BviTMe/nKUnjcwtCTwts/45lJAA
jsiG0pKBD6wr6I1z6vHCBgeUKOgLE6KlK3AV1HEDpec4V5nWao5O0NqDXM6DNFg0
i5g5xiLXNiyyNvJcBP9W9si+VJOvfMVsUPcH3e3Am77g0G8HpqBEbKGTeOJnAqlj
BLcRVcCfb5xYXT7yYckGFEDPtP4Sho2AOAtfb3x6SNxdp/ZglyooQbdvS4W9rBLU
GWKp7YJfnGApp6wbx0UpJ4ZIfbsaiq1UNUqQd5SZ5ErfcnUBn/0iPm3zSLurJbg9
rPusSzd69EbeX74AklZbEkVVc4IsLjyveJB191NWKr6oywgZOwHqCo2hSuTvAe1U
/OsZMKsAyTvYAhQcGbk7IfajN9plIqzRhyXzGxkVf8cr502hi/UlJcBQm5aPRT7r
bWq2f27z6AfgRipiSgPkNySfCel4QEgJy5MdREGlNbSvsyvpQYPnH/oCyCKA46fy
DfwUMK+sXsaKd/V9wZfXwk063ZfIQrv7CGqJEMrEYQa8t3OhZfzd/JZUJBPQEWxk
Tbl31/KD/lRWm8Av3qujW8+CfQ/wjX2S5WEvPZvMNBVDa4eLCi3sWCT2X3ArTgVQ
KBA6zyP2lqNTruZaoVX+hIUfu7cVKos2Jjf+9q7z4WoiwkgjuCPjJGn8m6PzMiFc
k0F22EP0ewozVIjg17oQ2UtcIRyFJ7VaE3e1pIwPxC2jSAw/kqhGUtacIfP1bjnE
H/6rMJQnoP6RNpJ4hmyHq9GBVJXXu4e/KOQmOnGlTQeAc+vvjYI/3TRwM/5Ymk7t
k2JikFpTh2YyyOfd+vPKtWfAwZzVSRZ6i2YCMa23PiYVxgtaL1R3ProPQEfScT1J
r4vTBpMA7XDh9JWW/cUOHpkN+Bs3DK8P9EzhAfqCVegJjHRWobTruyekQ41In2Q1
KRTSqv6hcozVJWmvsjZmifj2kCE3T74+u4NUeUsA2Q/Augmd6KE0ez8RZlwQqAk/
kQR+j6b52xlBc6INOJ5DffnmxrWWR47D3qiTMqp2ewmonlT9Yk0Ej8ffYpNEtAia
qlNQ/oLc1587ZFEvZTiKUM/CvjueyhyWa2pRg7MCaCKun/yGfoaQ6yFbEcVFe2+8
Xj0BibrN8IrUHWZPE3dunxyTNQdifZ6nqFdaqI9XSNcuSwLWcKJLrEa3ZlbcxYPH
t4LFsRK6T8i2zI0wff5JkJx9mxLIMrqtTWU7d7qSThI2SV7ehExux/sKfp5Bf1M5
7D9nhUWy1/Td7nOQMioYzseWFXR5SPtz6yxTrR3aM3SDzQw7bfobScfhz9QZ0YVh
m41sI+CAdU3ijsvL1GOq/cZUzPIsg9yoccVVt0ryVD4XKr2ygenwpRctaQ6hkcBO
LqZnapQGQMAJnzs5nTDCl3JdTYEc8ncY123Glo308ubFPOBsiu7awTEbBageqkH3
+Km4Z9GAYsCwK6hHFxO5erkFR+dnjbD4HEY/ky29rFp4U+JwGWFWlnQI2xGWqWd6
dGzwKS+hONST4liPqrcB0w/1zpCSKvq3wF53mZtjDcy9IYa50M5Wbh2wwCbMUBuI
tNWskLZV6ptTd4BepJ8uL8XUma3zRsiJATomJSfXywC3ouf8IMl4OYY8ilLKdvaM
Gdq8hx7SLiMvJGFdQvKu4DWnoGke79FyeSVhGs9IMUBSmRTV+GQyTrXJejpM003a
Mo6K/0v7GhO+XSySyLZlMl/kKA4PwlzFfkxzjQyGYsXevOSI2oaQnUD6qjnb+/+K
NU0ZwyNT+QuuksvVlX2GyRQKlQ9WUrb3093Z2F5LtQj/sK2Yn97OEk07QpVcGjAX
kGqalh1HxNoftlvqVnXCDSRnP+KVD/CDmDd7oZfB6zIX3OnCn0SjX6wT+6/OWdty
WmqGxygA6w2wwtsYgOvZCTzLkvZ3PWZB/jYImSJg5sRW2ylCYARN6JzXU6ciOCt4
hTHtNTfGuyzrb6zt8lI1l9Jh08qCCzsn18GhaJ580jk/qv/cjD7BqwQKxiChevw2
9Dz2bUvr5H/RSJSbNAC6RD/+79myhf6eh11wZBL0YqzgF8scLD/elx5gB3rw9Bp+
JUabzQa0nmeNToCyVttllAPvpPJP4lIg2XjR7FvHRijnOe4+bj/Ku1cx+0mJjnWD
8R2DRVjx1StXTB5QJqXiCbkrir2ycJMIv1ToR6EFBLCvZRGZbKDTTTNXGMMpjqyS
NRmte9ImNBNow+7KHSUpJ0q8G9bfMbzA7xNjYhBrhWIhQ9yRkFs1IXROKWhHrIzH
3jmBZP1BruCpQ3wa4RAUxnMXmZnfIVQU5LVBk8diFAotI3NFBZhSsTyiT3fQARYo
PCmm5JHFwJdPqnkZdmHcUQc7nWygxqtWD0ivrE5u3N/u2jk2ohXiWoXAXYJvXVuQ
8UuX1yxZ8s+neUEAOZ+b6CbOhmSdx6g8Zr53BILrUqBwqLrckVnwoFnpGuQLWZm8
eXfjcqV+beRSAyAkkPiMc1GmzZNs1NAD5Qs2smjjgfmjhJoTBJ598WCusk4JcatS
zBJs7+Sm9kFPwfjC0/yJxmXsR+3GK9jjE5xfccWkDKIV3/GO9tj+K/lX2KX5LMNp
xKuytRf3duflokoCyLdS9petwNF1Xegvu1tHrQ8CJ6Uhn4fJEzDrEzbZDSw34God
L886ByLY18O9XfecHywpXE9YI5Dh4/sh97i78he0GnuxkVuh6YkFUConxakewS+Q
bXQuCE0Har6xIU5Ei3BLLreFHttKHVY/J1ksmJULOUNEyLJ9jq8Gb3L98BRieKoq
HRrV3Y/TKJP2O0QY4ScIanoHoYQt9XDaBLQwNArX3oqBm6pa6kucMD+60YoKM/y8
hIJHaCr8KdtQWHW3XWgpe82c1IPwDeTwyy0I5TCo6wFngXPYKU161pAdYDdfHF6a
Ow6fVtVa/xWR7vglEDrLtup2MtkbpXEeN47mcnWOxZKGy/Ztb7WqaCK898ECOPg+
mybbdvOJnUC9QB1nlRD52wHWhcwzp8RmhV49M/LHGTvJmSusmm1u5FLqRRYKu4tl
+GOi1DoB9lzc2kL0tuToYBLrLWAYDGv+DRhDrMvIJGhVgnBHDdVw7ehfmY0pI0r4
Ve4OnwbG796mMwgeO9gT7pTR7vdusD3xQbU3U0YC1gtbLNtbckwuMlUUTvN9AiNn
N6tEzeeNHoUsbiAcylgo2PwcI67/cpHBjJFhlCChnjFcJyb7GxszTTEJ3mPK901N
5w2xlqL5sKmjAhDc6s4z37+rBYXepPQzQrC+3B1b3UEuyQT2AJKg5GVismEUDU+h
KRtnvRSIvb458D2n2Hy8a4cEntedN9tMiPgv0883tKeT2HXlofrjgsSM5eY2Zfp7
sg0UqWx/xQvW+b72NqQP9S6Lo4AD04lomTin3xhykNVIFXYZa81NCrwVezOn2x54
9n+NVkp6jK3078eo/4Sprdm4tUuRTgN+esPbqBMnbmeNMcLwvtnDC3Fv31coRzAF
9ZeHEUAgdZFrXmhUKW2XWVzhPbx+e0DTCWFQT0fce2H2P0yZfLwcg07fju3lTVwA
Pw/4yN2g07HxgfxslsX2ACQozDALNHH5r4aRA8MKHYHIAzJqHRDaRekI6Pk3X1UQ
k2Kv01MeidJlDaWmrcVJuVodgRg0Lg9L/gBVXMKEaBo3dKvBuWASm5xKyDb8LYVC
7PFXYAkyXWjDNk3DX039hLl/Yp74oF63odL8SExu1EV7nawOX0nU5/+fgXy5zabs
UahRfAeiKQ2dx/tD7Xh2I95DltKU2Z0PznLom0jKhF50dJhvWhtNI+intwmMmPoQ
QrKnH5lEl2OWHaoqhzPACisaMktks4wq2nb+1yTnSWQwNv5Jk5BA3kLz9ZavJNgd
TEVAtSkxp36aSoQaWwqtzh7BdwanvjUBvqfKbI0wzWRsSvq1BxCn3hr0K2PnBItU
yDIV6ZPF2aa/lQzOiZEKaaaSG9P2cVgm8AlbEfQJC/vNOlsMUpeVygMomuSVrsQ2
xlldpZlA9zCDBSL3kxX8e2fSBtUyINeDK82hpSM5DJSa/DZSjHgB4qRi5ssks+R6
Y3FYMTnoKjYUOtd12rHXXRD/ScEEc+jmRGIOOnl0JqzurRD3vUI+8POb5Bpd0QVZ
G/p07veclJ9Bct14D6H5xs4hS0oeJ/LZ47kqZspcoGaXND9Z6xwPm4vRYBNx7VH4
BNB2kanMQmapp3FjedS6n+NHqhxCQeeOPj8yN9H780X9sUllh6m/WXaLWrhZ0aDw
rKwH3OBKStfwtR7Rsvbjl62XOYyk8TnxZCfna8FOKgx2QbU6J8mtzmM4mr1ww/+G
68XG01DGl/QwXkZHmLRZFckG4FVr91DsdxY7u49JrwsLU5cUU4zs3WS1wjWEud9H
UJNaXt/2HYZzs3EA/EsCvkm91ZctqYOlVC/xJvCl/xzV1YTtNgnAHs6jGkfW4KnZ
oZDkAhBr6BBOuEO/ZDYo3/FbYSyJgmZmW4vNmOwQJxCSjXOb5Cg9XQgahAz43AbA
Fap96NkFOPyMDkA2KwcktVP60o7FGiIikCbTdGrmOIm2JMY5TP9uY53hga1V52RF
jDuTC+YzVGq4MgYZiU5NPqpxzZ7B/hhsHqNkglY5+WYckciGn5hMkDKQ0W69G4Rj
AjwTJaDvUxEdoDTRoGkeLxclFPVgTfMcONPXiQ/AAeb5CDjAimPnuvxpYf2Rjh7Y
KIoTmcMBFRzrYJL1oTy91vQ2mI+YZeUa2DoB99ofFakHeOCtVge2PFl9xJ/5nR4J
5aDDNjGUK06PJe4R+oKs04ejBhEw9eWgO6NfBliRM/ej2r3oX+lRsIaHaBQlQkPV
KIFxQbTc2G0SuHUV5CnFeFCyKt3iOV/Sf1UQmDKO41xWM7OZxT7hsqLT5TW7cMA0
MvPnpXzyX2t7sS1iUJo95jZ+pfr6LjuQz3AqxLA7B5O3b9bUNI+RF9kzSGKNPh8k
BZA8uiLvNUdMjFMKLDx9hvus010TaMKG19f9gUEGemK+qI6vS0PboRWT4fvvMGmo
zCvNMvpWTJZEaQEpUD8dLK8nvUgu2TFKdrc8qHT2Jg1qhqhGSYbNa0Y8FDNej2lf
BM5EEkB5og6+dbjlZKDKKE1fW//smAB+SEqqbtxVomXuhO9qiz3o2JOq5GYRGwAm
Sog2Uk1TEIU1YG5gqfuGoDA9xmTJBWvT2MeTIWRYo2JdfAatAo7JyuAd7FdEC5+7
fJuys4TPIdqbXtzH2nIepjyQ0gRK9icuI57chxVNhxL8ty6OH/1Gs6GOK8p8e0nS
dM+qLNoEnDuVMkLJAIL56shHFV4/cK1dDpr7MlDpXpAvhZ2fnreYDX7krLiOegK4
Eve6Ht78M/K5lnvtNOxpFKGfEuWGvfrNwiIYcS3A28+Zjfs9wW5QYabuoltS41GX
ZNGG2V2ybNM3G+S9zO9W8rMfkovv+siO7CHdHPbue8ysGkymHqGXO8eCuvN2qYTW
GOoeH/TqezJVh/ExEXrurdFTijooIIhRELIUCnX3Mxfmx/wlbUfAmlDvXYwsxTY+
LAnzE+ZXq8I36LdYgbzGQIP5JkWcf/RgVCysJ5r9BEXa9m9oZsm9xtmLW3E8OtzL
We9SpHbFOhcSt0XU9SSp/+exTMa8ul2UenbqRZKpCaP98d/b2PRcG4Ebg5hAkhtE
YEbRAwy8iQjfmskDVDBt7dDiMxIzRxwbhuSPZGoCVrDA3yvHG/UonWFAVdme06bK
oI51EwSiV0EPH4C9tKaQT3FawE2kseNHIIptjmivqkg4E8slQ7xv83by1Dq19zcB
KtqQMHbuhlVNuPD1ZUCjVWygdz9SbrVmFga1Bo0/UTHnefdCF8MROWOHB0kGF7HT
ry35mML5Gyjom8X/Y9NmZaDVO4cqu0hRkTs3d4zWseQGVKjp82nGhCYULUim7yNE
FtlHi8hW7c6j4wZoTL8vFBN/9ZOOs+shmHNll7TEEVK24wTsRi3pBpgTs3KSwF6Q
b3wc1l/firq+Jn6MgGgNwHHLW6ye8uKlSc33hR6LqJ93bBIdXgmZGUZkJjB2j1iL
1AkGu1eNGNsjXokvNzQFLzUtwQ/7xW+TQU7TgeiuKQ5sQxGx2IsnxXrUcz9cnXTr
96RmKfqVHrGpereNUiQVsqCmNMGxOAMP9gI9T5+PD/29UwS9fA67/44Tn8pDbkLm
5s63b7g3mA5M4Gn2v5kZvNoKtUVZ7tBoFvVMlHTSWFVQdyj8Cc8mYK7ZVFEQjsfV
IHOz5OEQtIxm/3wuYWlhW9M8lzlnxmV7z06NG7DY2FP8ssTm7lAaIe1pfkH63JeE
UYWxPR982Xp5nN6P6vAUNnrOQZ7Kzo5d7zjwvNhQVCh3WU2ffiWaEy5ulrVxA+up
uB6vcg8KB0MFdDZVO3iIANVHp8A/RbDgn/N7oFg+6R3f5VNV0wmCVscLx/YImYiu
D2adZ6/zQcIUTG9yr6tG9am7wBmxRMS3IIyMJivKNhQkmfuN8wGL7IQFozHu8sCD
vyco06vxjaGlXTAwgzzfCAk8O0Y6mGChYSQFCYoF7aYck++zGKlEGv64/uhU+7Ln
Ig1ajCTNMFJPsEtMd9Qu88XYug/sq0qZLI3g7NqhN1WX30nNqqKqNlG+G8xN1AsS
2obG3mPbTyzLNBXUfTBMg8w9Q1m3JZYxag5vnYdCrWk6Kz3NlOTOohBGAADJ/0XL
sxGsgotTkuTDGDjlQO3awr2ZYgtve5et9mekpNi5NB/Plrvjw71qwuJsGlPqzboq
aPeiphMe5de7LiKGSCE+K8fX54gKIN3fhpkM20CLXaJvIeb5mSELMsM4cMakOTZb
yxAA3SFic/w5tkMg1M1YTb9lztpdITjWerSdRuI+T4Qj2b5Cj+VdfLQ5ZnZwnxtn
sEZ9TN0Y6hAgVxdFbg0b7S/bhL32oBq27dCpGFTzlOmdfOg7cdZiiLUAPGfJ1f7G
qntAxPV0+edd0dJB9iGxujVtsvKcrf3ZMRtulbPxYPvwI7x5QzDcrZQB6n+9K33K
rkfLKORhuFdt9vThBFKBYiIIB7xCgrlSmLgn6JetHJa1VrFmqK5Da4IfwLQrAcs4
RsY8p1a7A9Tl872QlW8PfUMR6pfjs1wZfTwbU4bmNsEpl8cE2a2Mu+7aA5nJ83K+
WDsjVN+dgj2l6jO3EkFLjSzA29kuNxOREg6QSCLDDcmmPx4uQrpW68L43EilRHDv
GniM1kI0b/kXENYqmpE6kzQnrXJ7nPuCIjIJHjS6GCQ3XeWih9DNymoMU/SP3u8j
AF3dL0Lw55ERFO7xK+m45esvzh3evBWKGvzRCbmn6EQn3Yoe005yi2l5A5vEynqK
+TzDeXXVnZCiQyFz6XbaInM0J22CATxZZaWJJv5ecWWZrV3+8ahKy7l/Q/I1sxhm
SeRUhfecHqiwiW4wD4Co1lgb9ZQVs8xKcgscXP+d8sSwJu6RJA3wS6dhFijThbaY
y1hz87jRBF9NQNxKi37rhok2uUbnmFhm6V1QUUuhA35nFB3NSJFtyodrUAZu0G1y
7kMNnjZ8D5PUZTThNtRWvsE6nZFK8OACnABm9xs8v28JCzLKeOeUGZX9K9n2rRve
2511+d9QezjgXPfAylC+RECCRAu5Sw+YFm3pfqXSyMlWfjwEAFogHTpdHpN4UHCU
bOdPseS+cv//R2IgTlG/lBRdyt9vJWnx3p7vJJi9OtQ2Ife972DQkpiw/dyjxZsb
V2GwsXiZhBJfp9bC7P1knsYCKtZG+Qjo2M/jppa2ZLDLp+09x616yaYsddNB/Dgo
n+qSCe6xzHXAvOpCm1czGueKT4Fway31qIKRcCu6THxM8O6XsJ2/sHA0Qh1oOGY9
syJ2JbkYiD9pfgk9axDFx3sB6fZtA3sjmRVI/upqrTt/di+1ZBNHcUB8oSIH5MeP
gWB7yUWh59rV1vrYoaDJC/I0yb8h3SB6I1PYqbutKOzP6A0enCOQWQpOmb0nIFe5
JapPTP3UOzkX8B+jAvMWBPdXto2BsWMuL3o12K1QvUKzVAd78AOZoA9XqUXnA3ew
ukGdoTWshG/GXMCcVe0EzzY5khnUNS19Lp4bVVK7VFm87X4dtILmHnB/Uv5SVSCy
ERfe41bqN6zmZsfUh3xmukajBU9kuI0EXD3sbOGaAFawADW7uW3XrCATexYcbKg/
dWTDtS/M4up1tP/c/QMS1X3D4whbbXgNBST3V/AKf7nIIeOrmLGbn6mTpVvlCdHZ
NV5eEXnxASQBWypK4gATALyQ5YVcSLDClOwTNkY/y96jz1MhrKcwfY95+9mQKu5A
ViXfJydWv3K3zMGORByWVS4i3RUwLiGU8R7PvY28jPpEnY2m8dpWn0/UWvobT2Xm
KMguDoq8V36nUdakvK5J62dDyn15jnqsF0KhVcLCiSUo3N9aXD3gah8TLs0Asw84
gjmnM84lO9Aqyq/Bbw1i9pt6Z9n2UOTeDhhYUXY8p4ilGoxzggRwz8KB6xEyZyjP
aBciWblV7FkwSvRX7R8MepoG4oyRm17dhmJlXGL/JC6MI0aD11p+N4BoD/HnQYtF
oShq67crMHtO7eZpUWm7QC7CwZfDZOEsOvAEAV+gFfhK3RSU5d/JaBQi63LhfEET
wwrNgQbM3TsnHb9ianQBmbg1UCni8ggNnkbxPbL4FRzQa6M5PQsTBELjABo/3mrm
y3b//y6pbLuF7p/9HbKSEIJp3b8XD4Qptr2Yn3qzX/Y62gEjfVixn2wg8plVwhsd
sTjQJJtqcE/hC0iJHOk0dxnb/+c6DbFmD8Fb3/L8jVW2ThPMStL4G0VWpmAmhjfY
QpUt0NqgK1075+/Y2U3Ic2acB3xMvCQ4IUNp4Opj3yEe2kd3ZLjlk93VArh8HL01
8SWZm+7G1TCR2kLxnWlaDH7xbGpM2IFswfQxoWCSK53d6yxvVb4vChsR+HwbnuvK
3B97CokzmSG/1XBYT4Jf4MAZl5urg0afcp7llnd0XbQ9uU5ZQXNXPluXoSzB/OGO
XKzfG2qkUEPgnfDioKFSEXdEZdjHZgCXTYmieEJsJZozCZJnOLm6inw8To0Hxbtb
SgfxcpGaXqaONqpjqStqkHolWlbku66bV1g3gG5olRsceKK2JNw6Ib6L71Y2hjeV
T/9e9UVHunnl5AkPQ6/+X14oFkz1ut4jEMpKJFJ1Zn9JLG+KQRniH6zq/XUzA9CL
6I9W6LtYsuY3jU1lxLvtESCS98B9ecbYRkFc+Z68os+m09mkY6sWTp98UH4l4/ZD
i7tV/gw/V5Eo7icUhsJM8WIAMMn7tP7BITpi5tK0lFg6oi8VdUClo33PF+vpuTj2
3WmvvXOGhrwjf2gybDg7ogdhhyhrec7FVcN+oKtIbz7RWTMWTp2cOugO0X4+7YW0
GjacCGpjG0Ce6cQw3SeClm2jeJ0nSOAwYaTpKUf+BVgDLfgoZpKpi1k9T5VXET9t
6/5dnQiaDxznzb+03RXGVFAvTR3nXcCtC9C6Af2mxhxtTZfXX2xFd5z8m30N71Nt
OM60v+DATjdk0Efk2JQdyI4YuflwmPKpn5ljVXoABr7MkIMbkSTLJKtAovLqcIcB
ZYueTFQBmNzwF32U4WrkfKyePhiq9a3jduD7OkSCbuD8Iy/bn62DxH0DGdGM9pll
0T5+pK3gUReW/1trpQsap7oBexz4zMW3ZFkjqSEr73j1cIw6zTdnDTs7jdsrFLk/
iJylATQ4ml3mo6Uqn24r4+oGW6e+psUZ8WyLTt/fIT2OinXLAcFLNb8HgoZNGlSI
kYMusfknmPBonkD7fRE+GciPl4SkYFF3Cjc4E5rI13GKGunxivDXMts6GKrnxYs8
RTXcyFtxfh44x9wRhVz/5t9g4bkeJwHeteoJ48iNswLNdKLK7WdNs8ImlvkP5NHz
aNrD9Hx2DrNutktdaxTXfrAjVa8lTXt3vOuoMS7uC7f2CGkdM3bIjyAIkCbRRJOY
Ht8GLAXVZYS+b48q7nhzeJpeZQsVAQ79Uhi4a625CIHLMv3nmtKpKBiVbq+/MWBL
3XP+uRL0rCfgo0eHrDYPj0MdUPFNojLCekPGKpSirHmmwPirC5rR0HlKz8dJuHW5
uclyXxTcwe8+ULUtxs8bDprIC3J0r6zdYek2H/aPMnlLRJ40usmzE85FcbHWapnC
5Sky2vtO68BbO9kJQvlgFVC127aGNx/s4DwEFMiNKnxGqjdfZe6AjccuAoXSTXO6
xFOavPDRvd3wxXOaPNjO20ePZdUgKgfktS8W3C+xBemG5MxCZzE6QvdSuUfBWuiB
rVxG7qSvDIVKIEwxnL+/WrvcYBGEpECtaw96gNempLkl0kTeLnaGowsn/8pRL7rg
h/iMacCncoGKE1tBNNj3MxmBR0tzLFzLyv9utDihdRCybWagWrXSL7LsZ7HMWk2z
E9KDw/2SqGvEDdcUDPDVU+VrT21fNp98MQkAY92mLNZkl/TbiquLe80Sq6Wep1Q7
8zKNCHVOYVyIZ/KNJQN+exERU3DcJkaDkaKTGHoDR9cgUsMHErY8qgrPbBRz9er1
vtGgtN0FAuiae17En3RxVvbvO+nx9Qr9EJaQIhjRiazPfkAh2fuUXVV0bLkhsAZn
qaM8x0KSGfm+b23lUGxR8mHWNt/7I13lYPP+YOnHdgDgaiLRjhSDlvBObyU+7wjd
HR0hI1S8/b7JpGqIatqTF12zE9pt0NUv84Dii6iowOmRB2VZ1PNLfwYhH86XKGrc
YwnVxUgjFEsncIOlIffle5yjNsbeHpwa7YnXYlnb9TA7OQgoxMa2wh7te59VJ+5K
YLoLu/fmTBx+/X6/IoeC+sH7+B5f9qX0R4XZW7MXvHBpBkossjSaiYJrZxo1XSXp
FzYqJTukM23PtO9V8PBjfckey3SsAgf1cz+u6Rtlll47b24hEkw3UYrRcZKFEyd7
1Muj/Ro4WtrO4geEfPgx+vS9zkFcf+hL4XXHfIZ1Kp7jVuek8EbVUSc4VeirTm3T
Iv8STlT0dmgqLIFr1H9HI3xVq8y5n8vNiutIB/b3n5Gn4RW6ThS+Pg5G+3TMd1WD
xkrTdd0CBUUc5bFnBWleumOpsrkO71sYfvW8IDQ5qEQ5jrCNckZAm4z0WzQWuodz
cV/0cwI2k5dnMGALnwQ2h/7XByAEV/gI84/DDm7/DcCYfOIxvQLlU/BC9yRpLEO+
iYW6e00n6vTMYaxpr1OjE/xcPOi1AP9XQfn7A2NGeq7yxD1/YflPorWFWb2YEp/9
DwhPF9mW3RjN0cUBlijqEjJ+fvgMIrxr58UTlwuzZx2tgOgTwBKYJjBhUnhONtGf
k5O40z5hY9/oFaG8fQ3ZuzVYQcK0/ks7vBE0IgVQ6mtsXAqru1EEKe/i9AnKYC+V
wTPl8RPauvsXQf4ueSAtqklz0FzrKAbgqrQ/8KPLwJQZOMqEMIfy/XdF3SRlJ8ld
SlAiZRQf7mo1LXLnO39kTqiRsPyNfvXe9xWDcBEGPusYp/wLdi18GYSxIz/bk5gr
62tiAgyvja2Pq1abWtVnEAMiOT6SU4CQBcha4b+7ha+v5TsS6+9BElihE/zjd9b6
ks6qdobH3qvoT7RWvBJ2kGmXMLof+cMTzG26U/rIMHO8Ce9cBYR8X3WcMhaM2l7o
m9vjBSXkrG+kZkfwsMfkRAfHzR5Car59ufjlM5fMLzolg5M0IOCgAoQ0alxtINMM
ap17j1PtrR2eh8RUzLnLK5YS3vVs0IGEDCKtw1RIaZfBqmNNPi1wdBbipYCbX25Q
V6Ill8vPWVvMpQHHvqluqQJEmpRCDEUEWBYBBRAoBD4FotInGEK9ul70pFqwVpxy
MTw24faJLkjd/D3W2MDRwfscmGFylHmqf0KkpLdENgrYqCtGcw1KN6F9mOoqQBLH
R0xikTLIzX8zkAygot7skgLEehYVlND/ZdtxsCzd9sbnUmKd7arJ9gpkgwUYsi0i
FzC08pM2ZmUgfFVEyfLbIRTr1RN2b5vQhulKRJ2CUv352XV+TBkgg+PA66BO+C/G
hTkohYuStk39Q2oHIl7StF7PN4kDOJf818UYtaHhW675RKNmucUhTbJvEMSWuVfN
qJ2AOYqtDcOU6XVbJqEnsFYzcOj7Vhryg4kCkR/I8tLTkYYqdi+vOy5WMZonlR18
6aTCX+6Zzy2krc5spTqFoSc8+J0XYzZmjRyJq6RBDZkZ4pkVZQvW/KjgNyNSaxO3
F43hbzqyAduLqPagwMdNCb8Akc29HDbp+SfsW5HVSZ77AF2KymImT1BiSQxn5LKz
2o/n2tbVsZoCV130JKTwWhOcBWrnBS37YxICpGwUsmc1PlwMJjtpIuFGvI4kL4Jm
i1kzNKzXQtg71k0Zsa7PvLGkHz3Oo0+TAX7v0vBHWJct7CmJKyD+ngNvqSOfbQv/
09guPhrysHBWPbhZzfO1fTCjADLM9+NuvRhYxo/T4ALooi8IF/a3AXnaGWF35Q20
gN69FZtli0/kKI231ACbWhZ32a6SDs3MVDEAH9L5BbIX+roD89YjvVrzsNHJ7Mvg
YhDxrXp0QrMcEXtct/pq9x1lLfOPws2zhUlmPlA6GE2QLjottEs3PmxFn5Ukbtns
ppeocw0XnsSB07bWHZuc7ej0TSEgl12SxH4tx12p4dCq6Tt/B8iysFmde/s7Jwzd
uLAZDaXpRt1Er4dwo5so4uHAEn+zENAEMSFBQy5TIgoaDe+GJz+J7tPsamgsRKgC
wcub7QXO0wMvDtzxVpfOK0/XS8S7dePQ97H17FIV1r/kqSllRicu3+nmvobcFNId
bfwmvccZodEF4sg/3mZIQjQ1J2U8uSjfYYzoLHO9oURTVePAkMugCtQ2QQzSl4uu
45bRkpajGEkM92njmVykRq+1Z8ZhZ8i5ZNweIpsJa5vnvUeIPjpHdLj22tHkqxV8
kNXFMYkeiqoCK/VbSkzmr1ZMC1WzOBKGUj3oN3eGatgZkjbcveg2P0Zih10o2xl5
B5RW5cjE5Yjy0eLMnligKXAf3Q6F9eKm2ZjWEgcg3rdKh/mftlRyYHanc55+azQD
xFdRdGm3pJlBo5RxBBRoE/sKcQgk0kGl6bcHTEJX4N+nQZ7yfKbkHirpny2qGSjH
mrHop555L6PFY5t9PoImM4gC4BgS7UCz9AF0Wx00RkrfoJcUvjETJDYobXZWaVnZ
katzfu2fxAsr1HLNJs53NU+G2WmSDErJUQ0l583UrbcWRbkc+mSHMOtn4nG8SNAN
PXFfjxOMAvuEDaspszO+gU5ZCJnhKZa+Dz161CpIJyAqqqgY54io/LHVjV+rCuZo
7aiHcldoaNtqchq1VIFull7s+wFq+O4RHQ0L73mDoyXOj10tSAB0wRSiU0wmdjod
guA8fCbbtErbPI0ZSucA4kHQ2Q+qKlwddK4CKPiQTCtS66o0fTBn1V3W3ZymmGpv
eUOJVgNfXlwSkrffa4Dr+l6ytnNP48CZ2I/0pVdecG4s18v1U49AobNaIKgy+emX
esrIwY6ll84k2fk5IR7Kv9Y+8nGGKppejEsIQnIU43kvbqiO4gTA4XjKMGjKBtqm
2IQlt5ChBjLBgLy5zzkZznclNOS3sy813VbjV+SoOWFJpWB0A3zgrNe+H/6OmliS
Hch0I6SZLf1YkvNzE4zpw5QXazw4X3RkJQiMKrzzqF1pM0S5V885p6+MbtOzkQak
8T2sT4ejUzCfV9ifZo4D64+3hfKlGt5YvplsKOui7cxdoLlPJWntJMaEP2ftTcSA
+vtczVF4qo5pCQPHm+iKq317goCPVwm8fxOnxYipOVHk7F5Iu1LqpvUeSbSFRbij
qc+oVaWEQ989BMAykbf7rqPhNnx6jT+ERgdAieimPP+VQ3211fpPIVKn5Z+tV8Ie
oNGwtYMK/99O6rBdg9eG+Xedk8zx5Xh4ETq8iR/9xXJuf2uoF1zkyL6VZhJ63iNb
pdd0UspjrInVDNXSVwY1LVNI1vJNAVM867qHZfvnzqEo41rCj/zF2lqE3n9SVFtf
aFzj7YkXVGwnJq7vVRKoocy38yb66rLvxcuj2evQYEPbu45VZ4w9i7yHERbMpDzj
6rfeU8a8CRLjn1SHejkE5hHxPzRVd91rQ7EveNpeXkRjD6ExehuglfUTdwDnAH5F
/tRQqBYrMfBjf70tEmpgS+wfTytdkNX1jKzGYAMrCE7fkucfXfGjxryy+7M97x4R
VLnyS0N+sKy78e4lXXcreJYhfqhJYkABCmxzeqiX6/57YoUy1KGXHBp7hVZ4Jgrm
q6vW+sKQKnZdowlC0vrOpO5NX9d3Gv2W3MFHLMB+popuBmWiYOpxDW9OuDGi4xHo
8Tq2fZSbyj7KUVHFm591Zcrd8i1HXOSeV3m1LGy9VpSqS3q61O0CEIIvbdF53XXV
I3QDvmRUI4pRPKMKIi3ieN+fKLiNfoyOLkBfLMEeYPtcGIt2FRBL3S4QEPZN/VpH
cL11RrynsE/9pSdtTxO7g53REOL75DuxJDBBEuMZphqqlSfue+8Ld+Zhkb/IdrZY
+kCgz54rU8ZryoOgtvojNoO+asSQOXuescszzKwdNYrrVAfW0MHOUbs3TdG9MHHa
9dzdOhu/399EBET9Q8Ps9n9Cubj5DRqM3f8PnaseORWgoF5IC75veIO9iqrMrrR8
14z7bcDGlrSs8hb89wC4UjWGoT/TaoyZBWOeo93Jr9dlTLCUKG+Om+AfT9i3XFxX
OS/AOdZw8gG7Ot8Xv/waeJF3XUG/Td9VbIkhC6okGufB8RjG7/wQYGjDwyTbGwo5
SyUPPg48SroU3WQKBuGsSBfGeB4sHsgPxg87QZwwNbqxZmWZS1nHNCaYzkvFEE4j
hqtUWDoqMcx4ZJEW3kEFJs4G1bLBshnWppu8CwqJgp7OOue30pwr3H3IZYqz92cY
uHG95b/87/8qxg4tq/8SA4RqiaSssDipMss43uVUzM7Q+4vVsB/pgFcpDEl6ybma
WB1opFXAznsE/06f2UxPfmwEXewpXqk/7ixgfG3RS4xfjx8eFKUzeSf1Uhkmb3GT
flM96rjMFRrbpxrwZQOiiuOfyo5D/TSyYUMVTEtacxNyk9S1zQL0YwsmDJw+wKp2
Gtdh/SMnwuIXiWP5Ibo+ZrkX0RI5DY3LbHFQ5UA/qnO9KXwCfL3F8lJPVUqqTWD9
0j1+kKTWINDOoaoquyY3FqQv3bKeKoAVeKu2wmQfRMYdAc4TSEr5YvuUR48ZWMzT
3Qwyaj0vHBQuoJpxPTPxA6Zgk7RaLQ9H2eul49ElLydjXO0lqNORunufZJdZ9oSw
BbeG36GwxbdbwAL8NmzpoV6hkJVkGvvZq1hafm3XlHHW2lFXzxzB+ZIh2d5lZ102
9Qzk9NeyIPFGzptLIPvL6MIcj8qJrbgPJBBjnAGp0Mp8QV+Aa9UHJ4uEeCuA0StW
9cNd6WLA+gzYSvdzlkItAwv5FempOqpc4jarOyqrozByQRS2fsEzSSp0791mY7k7
DhaexS7QAAmJYGQNjAZSydC2txO/kBps/ekpOVQGUCFYbEPdnI/Be0x5MRmMX1ZD
Zkgnejev21wig3rTpzBfSqu2Zh0FaUgMZ5eyNkpzSVYB3pMUuIhSEoYEfgvxlVSl
2jFlHSWxYWsSFlU91bnVZzjrRpeJ5nHEzj8XrH3yepkdTmUEGR12EDLyAtc95EGq
VXeVFLZ5Sf1IVohpJ+Z5ORZE0hAvlqL/6HLVOXT7h/ASWNpfsT0ZFJpaN4N3Gq2q
iTVm3pmdaCD0qJj5Z2A/KISCCO/9vkTK8Ej82EFiqNfI+IxlVr/fJgZqIcAxe8RY
VDo3GGtuZGu7sWZcjKiHbUy+IYk5+4G6QaWgdenUuRe2Oip/8wk+2H4Fo92OH/0c
/xXnB4ObS59vsefoJWBVWsMYOtBI5xd08FczUdiVpJ6/NQ2V6W8Kex5C7j/jERvs
uYBL779EDhfeRAzM/6Bv2+GHQzOG8kf2xJj1hEy5yrJQBGPKKD9pE434rhO38oiU
EcxM7Qb2dE4hW0kIN39/pw5b6FYBU+2Ay5qUwUOMn3ZqvByCUvtY4Qw85eKKuvmg
seAB3ZfZPwOTEVnW3xZgyDF3jUiP26zpIVeeZ4iQi0XP+myMNLLRpKlTDAaw3f3i
EGUPZOu5GZnfIaO8iutzUNKvvS+3O7budttHaiZK6Io5z+9r6mA1MSnzoAh2qHsc
7c31k22J1GCwvPSyxgaFAwWc1Eo7ns3zawZatRsePlKCJGeX712luRiMjQw4vC7Z
/Win0TgDI6jwaxYvpBtcsgAAfWiidXKAhUOd1o8L8eyk9btOcrtB48s799wijiru
0rnJBZtKOEI/Q/jv/lvojxN3p1ykyfInPLh5hrT7P+4PVlJ1HOwDPIkzBVxhFOGu
td+5IJRrvW7/X7JUquQ5xz0DmOjQbHRY8EbSiuhY2wt6X9hoiC22Ht9aF5Zyldcj
I1J0mt9Z3u9IeYjS+t8nyf+CKokjNRUpPQihrDfDi1kffd2A+mbyt77CUGn5w9JN
03VOcssmkt2RY6cNrt2sLXT8nbASYLsCTXqAp3/QPQJ8ah0z+bh4SDTizPoBnpW1
RpNDqlzmZY5ffefJVUU7yxC93ZDoDezy8OHcrMdRdz/DwxZxlHXaMLb6zSpHDFeo
kpP5NwgPRlDqTvvSCUh60cz2DD2XisOxopgD+TwG7iNOTHEq8hfppON9oLhrf0Tf
JxBFZjM+a/7ywh0l2ePrfctgpRYeqS5geSZOgyOOAft2IX4KQPzDa1opxbmjbHbw
kU//KMUvt7tKFUnrK5MIZyUd7SeZASEPUCvhk/erWCuWruAyh0KZe7W0xMOp7egk
3kcLLRZjmYBHKohR+XMMPI9OiUOQ4GLoc9oqAi+92L5/BTsLp/KavtUobH0t9/PA
YFZgjiF4g7S3pUvpvKoI+/knnJ0PKbmzfG3fI3xP3546j4HuT6/ZxcbS1WRH9saW
gVnnw7e/fs/3JD+XNgTIsFo0ezLcvFIvnaS+MiAeK6nUY37QAtuR73GeBZspZA87
NoJ+XphVpd4LkGTHP97taMrnQedbHvLsu1FVBuh1BgB4/KOhx5sqEP/2AShtceWS
ItF4EwgxOf6YKNvaWbZQBzTJKbSQS+CRfmQGF1f6Oc6+68Oyc9kFN/8OUz6xds4y
jhDinbbwbCix3nHk3NfwODRfhZFDwDcy41uPgEBx2xhUmqCBQs9IPx2IEPtkjYnJ
c4LI3NsSMvyadqaiiUYcsybXyZey6tgH6KBwnUUhnzYzlRi3EK9UwOhCz+wQX97n
Iqg9mxZkz64ccngqsGdhIkX8VgtFJIANrrKkGbUp3WLU22xo1rwu+pHE9sAjJHzp
Pt+zf5zE2NPIRtWxSDQgrqIS1xErFqVl92VITfnlQD+UOx/9p0XfDm3c+H0LjNeu
Iq9nLgBnROR50pmlm07vyTUOGgsbbdhwgpo8oI3K7TqThQJGwEsKsQRFEYkQ7M0+
oEZ7o4eAGjAJiDD6jP5TUPSR5e3F1zGVBIKZ33H+7EG81OJsmMsSpmLNHPZCKyvx
MmHMAfdu6rBWb5JHXK3Vd4KLC6bb620eWui3fTbv4isAg/OJnuUopHrWWUZOSlNh
M49DOdPMe+b01YLXi0/zUrdybMxThXzjcNAj8LZmfiWljpur19rw7SgVlxS6J1iH
pW1VoHTdPRB0aQ6vBAWrJb9nK7/nRNykz5VuDXdFo9ymdWMAQ86HpkOuf2a8HLFv
v+XATUTtF4+BuCHCqkxHKQ1ImJTeWMabhqkcByk3gC9BVZc74i/lySimiFypcA/r
2XROWtDS4wF+7a2oyWPMW8xKwbxg7whCy/nkSch8rIdjOHUkrt17PCz8uyDr/XiZ
Cfj7rCsaGm65T5bG6PQkcKSPRcccEW7gouQD3K3KqkRtxznHkVmCHG6IxTGd3Fch
7LJc8hQz8csKhOGOxy5LHep8E438z55uhl+ycfH2LUSfK73u6VJWsVzJpRWyqWzP
vUWtuN507arg0al9kxjWY3VbbHguKFmsWTyyc2EhpK43A/UL5iJqgngVhxA1a8i8
QcL5bif0x9m/kl+pGdqwRYz2dFr5D2KeUZnWh0OehH0Qib/CqUhuCywm7Mv2oklI
EKtm7K0t6uy2jARZG+zIRHPgOLJh8MOqEqVWWpqeEjfD2rGs7TQQGfHlusJSoXox
RKQhr31tkVs/hJMNEDLMJeULM7LgzbpT9w/3mr82C49Ge7WmAWpgFyJCoUi0a5bc
KMLfXuNh7DQgl1KZcVCYRg2g8EBuY1rimA3Y22RquG7gNSfehz40UohihUG5QJdA
RSZpMWKrEolnWdRhtGY7xdlnDKclQX9QZ/LLSaCBsUqAEjuW4PSU2oiSIs2ipKeL
Xms1YnmCgCQNjSnDAyeJwFqb5vAn2hf+nO0TKc0yZDBraWCBIhoQs19ne3GeGSxf
YmxcJUTkVABgTJkZQByuq+RIhbvsvsxPsnP470Da/YzZBOQMtHQBXqsclaTCfRwt
aOw2oxmVSNmuTlX3PpUhv8gRXJD7zdiBMuHen2Wzr6Ja5HWTFHNkr5fCSx1mR6FC
cOVmJiaQqfajZqjXYLPg3sHiM/Y5/dbsz8WWEXxj2ACsemEcYf98Z4dlwbGNDUGt
mvDlWm49bGECzuy/ZB5tVkYNrRlLHWTiWPdOGjYO4ac7V4wEa5whpjI2/nPDp6V7
rAlsrr1aVU9D5zIi632lsYDdF4Wl19HO+u7itpmQh84wQisz4amqjGyuXUvTdmyt
vOedyK5t/ChXczuIz7nUxABy2T12TzW3YIfUYKLXQFED81H1q33i4GlQSdIaDkOR
xl+we54CdhIimwFyayj/yghjGTavCbxfyvqWIYeUms1n+lGHvHpkHvJwjpdPyhpV
PxSqMnJPxOFBwhJPzixwIRhWaCpQTsm885JZk2pC17t10B56FmDjRT1r0TomCFR6
LXf2/jRjAgNW0rQbMqi3ZwSEc4Nfj7R6GTCowDQLz750D9QPUVsd38RvebqOzgug
Q7bW3zBNulghfzsy60Ne+3XrpmQX+h880x3C27azmoOyo2uvADc4geJ+A4i7RWWn
mk5Xre3aVsvWeaAnFFrDfYAiVXmOSJGY6Bobz5tfu2LJ2Mxxdvb6AV4IfbQFoPUf
+F53RreBJWTvMqLabL4qfIYMxGwF7qasMwxiu173fy0IXChRhDc1sgGk/X45ereI
KuFzmiOALKADAnzuThnD9l9zoYDiT3E0hy2Uxbef3sio/jF0iE3uPJhAVmbtahao
lsnzxkpSrNLxqBfllZuORm8jXULADfsl/EFwuVj+PLGDcLfOTI6kCesi8YPAGMzy
k5ZtOVaSRcHOZJL40qZGwKNCg7JB+Zpov9FbTty4EYGXt8ojr9m3+rrUGsGPW0jx
HjHE7i2tC+d4JHuH7s4EOa1/dTMrDmksDqog3+cN2ad4FXflk2SO/cWn+AEnQAdF
YmW5zWADli7LRVCDCtC6kLVdWCYJBnAsgNQSiByk+DdhUW5fUJKQ+2FSu3vs9xtp
tuGmLMngk/QYJUV/aPeQeNg9t4xa5pO67SVhNNWYZXpwZt0UALwlZpMifM8PNClu
vBzQV3pJzUD+vWbragn44GsldHBt3291AuI6V/LMDpB8ybJ1V6jfyMlQM68nNZ71
bP18kTO2QSZzXXY/44k2kVnCdLIedASZPRTbsJNEpifYRpCCvrN6S1l+woKBZQkw
qZAoSgl3iiw7vpREN9g/PZ3glhgEmRaDc9TJ7dPSnlZ5K+YwzPiPyZdk9DWLRM5x
8mocnLNDL2mQom3YJG3IR5sg2UrHR+Q9vj7yREmmGI+4RQdnn4q0R3RqW+rFgRFe
AyGA6Pe9xq0iv7LzVgNGqpHLQ8HyqbpZ4Dal8Do5Fmo0sgMAA409Fgk1OpVvygIg
QjOwg6iBPXJJQC4JItTUbLCkNHaacWYDW0hCNfO6OKSdOmZErZEPhgiOUPg8gJoW
zo9bI0a00zt5avCbJiYTaOeUAp2F6zNV8VM/tBsqtn8NXjPrdF+/viCTFYVZCcfZ
Gk4ySMKu0va4QicIsYG7G2Ys5jEcEiyxuD5lRtlpYmhU6U3eBCPSIXj7mF3Ys/WI
4mmM4/xuRdCrzFtm8WHtBaaLStzE1KjTGHlqg4EX/4GUT8vHc3AZ1OUxxMZJXNSh
56FhnoLXLejOjpe0RvlBdFZB3Bae7VvcewP2E+zY6lAHqnZeWRRYeTBK81Bgj+Ky
rpSiOpwLDnycG/yJWGzLwHFoGPR28rEJvQi2lqFyM87ij6hk1jNUwUH1RNXOV/W1
PV6VPyZmEYtVFU6+6uMcwEaGZm744T9uVgVdaaQ398ImvXcu5riKpukHmJAUSUyq
hBuQyQozBPjqZwqJJtNx7gm6WU0zi5IuVvh7landL3U01pbZ5Es403jzY16JiYGi
oD68iqIbKSkdvbwLxRNoldCUUewVyityZCGC+ZMhOPYgWE0vMob9+LRc7XiU5Z/P
4EOrm/EHbsoS7ZVuHP3TH4212bMJnxjYrh932+Dj3y42U7QF6YOR8wYzvv0DLwW+
cD6AXep192GhCbhim0wKX0y0Lmm/qAwMynQfASR3tj+RlPPsskfieVT5mQJdk2nS
CDLG4//XfBsXSU7JheCzimCYv5SaW+FlJFZ75wWzvUjMaibPHukGEbtZ1DwKDhWM
MSdqJSpJImmmvX8gP2kmpP4Di6mj/RwY6vq4QOPf2lkg3gD6zx39OTKa55eaL1q+
cY6lpU9v17q7mfikbsLbc1Hh665RuAFBhceuAikrO0RVcJAP5NfmPsk0d35cTi9r
e/IHHJ1txAH5Vv0BgNtJH/94mRXExiuK56FM1m2fwedDl7d/9DWd0wFnXy1Yfg1A
EoM/CssL3YDFyooWFtYbYb/o8sWRlpGVbsb1M+dcgpNDwh6z+5cvW6JG+HFwMhOC
xm9Vh1sqPgKjJ3XgVgwHTMR9oKveyieC1+nqxRhv+5S5dIvU2NfpJ4PMd8psEQiG
h2MnKCT6J0P1o9XU6E8Jf8QgfLUUf2oCoFRm3qXqXajrw8euffbsap+Z+4GdYxcn
6JEKeqTs6dXmVk8LKHcKWr8MkaFvhccHATwO4H9NukoucZjNHGnmRuMa4+WA5jtC
6MNhpbNs23galKx/+QVPcWEhS6SaH1+Obx5dJA/4MN7hGWunVl7X0TsVS50LkrJZ
0PzO0RcoQpFCQ56JnsSo85uwk9yF639eEA3G5alGrz4/+c20IKjjOc79j7jXOvQt
UFB9k47uL58Y5Nw/6eTEpoeUFBnitI+gTADwt5ukoQ2AOjcxriGs0h98uphbHGpF
yeCIp//RRlcCfEOMO2TGUgIve8XOhf/XODmSGgt2pDRCjycb9gPoJj2ekNo3wIMM
8upsh3KeYld+nsIJ7zLFNyqtRNAniOkXeaKi5L7/q3D9EsOYfG/Beut+uzSgsjrF
HF01cHu2hrJQqMuCwiJz5s6oGWRMCNc14k3SkBL+LVMqqPcjTNSDqv+7qcdeOAMK
t89YshRrXiGNNQAbVsI3kmnBJvoH+leVRl9I+4zYbIUhdxFn64Q5lc8ZZ3PPpnWN
ywcro4vvqKFBOSFgvhlNj6fRc+Ez/FidLJdPNfSCjpC2PyB5i/DuhzYWfEXQuF7v
xGq6LpGwNRqJNkWe087G5qBIdMcOktga5ssgpqXOFFiXhzvy0annLHeI5X6NSdiN
ZnEsWO9KRnzrHqubkgK+MOI3+P1DKWC1wBNX5+kmROoLohxWTyvT4Ndp1zG/rAUS
HPTFRdy3mGpvexj93uBy4JBb3iRZi1FI2/kvS555WLefSqPSacKKojWLY/WkSdIj
KYMA3u2BhtwM8LtTC5yZnzn5CWXMLr7rVvtXw9PZV36G+ZWITNKuvTLRFNWGA8HP
WSiwH8FFbu0FjhwJS0CxZHyv2XTaCe77lpVZsdpDNBXCb6c+r7hEs4VpF/2RM7aH
4ozOeL+ifW4wpakTHaggYio/yr2F0E+KrRrsbVShbcsRU1CTNBzBOdkpvNg10Hbq
2XRkRFRggm9GV30yxrjZ7s9SNuXMLctHdB+yCdFdku3MRN23kiRn01VAtxkWomR5
x/kRHHn8zvv1l08h0leg8+REA2Ou6Ng07ReaTCU0tbr947LQ2WM4Fg068ne7zk8Z
Qgf+7rfBYwFFrtkvm7xU3ymYflkhhq/Qy9GsiYkjnXiHs1mDKWeX96s2TLJSQJjI
u5OWWUjgfw0seUIXDf3WvmSEru8Q53Ypi5s+yetb7+tB5TRr+AcNbOCXPI+C/TRt
Ks+hB1XQhfkDeJXGHY7bHd2Uu6xDbKU2JIORZ30CqBVEYwyZkD76aWD1mA/9zoog
5HYw1Ws3KqkXIfH9pfE+qMMHcFyOXlFvuXe+uaUDHqYRuK+oYl/ZUGTLpZlpxJRt
VvgJH/E7jo5wNgGO1vNq99Cvf52h9cjl68FHvbQ7oVZtmhGC+KNMm0vczanIx3U0
oWZK2G5h7kXqXLYSMeFZWLvpS94lOjqJz26kQGVOsaHSFUgDJsneQqb9VLZt/iNz
AVZRKIknBCqfiDB8OC2JwDtKbUa79Xy0O4WHEMrV3v2nTXqE8mNq870m4i2pkPjN
7FYepqRg8GFDrOKd3MzunjeNPNSFlCev06UamgPHEigqW8xs26XY6yoAPO+PbOVT
nMzTZrGJyWJ5FLo9wW506zJizJ8INfwnL+uhKz0+oFqxzByij6T2HgCNssH3nbtg
XzgQHQzRmVhD2eytndzN9Fk2LVWjlKzv5E7fU6rNT3E25GwrViVZAY5MkrLR0g5C
Rm0uYn9em0WAiVQAXu1WQMl1DfMKcgS9zywkZKWJVU0m6wS072F3iRJf1VnkYcCd
MaDA+oMPiVreonEhcAvg8OSaL2NsjdIQTxXh1DHJ7H2mn4WgcnmkwJQWvYilniUp
57xBUlJx88XxG+bXUiBOqXHF+QfXNbaqNBIrVN5PtY/xeB8EeXqCKIxm5aijp2rV
49f7b+8NoJUnPIz1GMYGs4yYw5gv3hC3MgWo9Pa2wsgDV7Mm/KyYwS6QIAVyA3X2
H01ATAkQM/2PXh7ezHKVlnLgzIaL+7u6McVZFOt1xxbThJyFnLi7nOFHON1FAsUQ
zAw6Tbv4xya6MJ67ba5mT60uMMZI3D81XccS2wyIzNHGEw4FRESlA+qLmYemU+ap
fJfZjetNIot512qZ8wosV7cVY4+0E6pMjq1n9L953rExkTqAR78tLcAQUfETC1Ku
aVhX7zEwSax7R2FacwwK9l9XkChczXqC040DT3ZArKhPBuG4y92dzXbaAU/aKtPA
0KEVWeCFmFAFlX0HItnhgERSXHIRUFhiF4h+jHN72kFM6+hmHQi9/tjHaVro6aCY
NQsYHAFEoJx2sDb4FZhZeQJjMxW170HgRybQC47aWwVS9t0Z1yv7vRzyf1RMUMpT
q7lGk4fw4dxj4qq+rHNKD/5a9UG0/EjjZ59fYp6fyHn2WuptERxvSleEW5yjoNEK
DZrX+lR+eEOhGrwBRZLQgHxQW4R0Q4S8yVa3+yjl+JYcsyOUUTq+EFy/dLv6E5+S
bplK3Nxhhfaj5/QVhVDGVoL5U6hGnyfqnuij/biKhhuOV2Ehu6lY53O7yHR+LBVD
975Jn4UmKflMeLwSKXv1+UGAXr+/Q2ju2XFroLRJTPjHzG+nsVnNEriysVpwOIQ6
QbNB4/SENo6rTtuGu6pcdlpJmWbvo/KGzF00DO2kLX1sDBvhiK7g2n8szH30cVFy
XgSJcxYHcMmC013o/hMJGQzNMq+gApBL5FCnTZJqhwasenVUJV2XWKGEkkdo7WhX
Ef0+n+kEunkTUs8qkLnv0i/fJNqslNpnMxfwBMuqifVWdCfzRDQqOPfepSiEYwWi
GA6vKtTdu2g+w6CA+2x7k8WvZMeQoSJ1T+OdVE1WMw//27+sL8AzocHgtznB+xkk
wKAJJ70BjxS5latGu9vWV0+XDK6cjxUmQgOprTGwuhJ+dl0uBQvg6ozwfPU7CEMw
y7RknBJ6v5FhprU/GsPPRKQLd+hsToK+oTN2Dz4oIL3Rt2OPzIF155qn4O+RZktI
b/e4APpT+gGeloycjpe1TJ1HKbuxylit/xmTgc0Xb7RvWH3DQDogKpcFilIy80Ht
SzFX9HOn3TmCbTxCEFHgBigrptHkOkSQnYqWSFPGzmEDs27okWD0VMjoAGKEAHnw
sy3ToyyC3pPZ57ssUB6mqUoiP+wzSq90xc4DOzXgiPzwROQPf2vQ2yrzogPIZx6Y
AIbRwIumN2cd1sxlZi5DznHLVeW119Axl/4jPLU4miNOWe5FZUSdBcFS1/CG5Gs1
YdWs86QhwnOAaxYSmgbyn9KSD+ppXJutPUSfvLkOkH5MIj5ZUdiKxJFIJW92bgwp
K86LmUVxFkUQVydrGUxvB9N6Nv7b5+bmEB35l5QPB6ZKqNmcAR8gD9ry3Kfl/J2M
TAyaai8/SAwAG4tPmRZq47ne3VXZS01U+794k48ejoiYNf3HYwwYHWMBk6LsCt6p
UDE3ZhWTPgw6RyrXd8FmEcnFSOxil1mQKW/7oT9WQBBiKtvlgQgxDNbMHMqb+QXP
JDC8FAtCcYUoAqhx2ZMV/SCJLU/7svcUjJb/QNPK/Lv8NXuA0tiaE0fKdrGuWfg8
8+G1Cq+XTp76gLZth26UmDic/+mo6Gb7K68MSmpqcMJC/b85m7uv+/+2wGb+GyHe
ACPdRB2iqarak3YDEunBIKmfX75qcBiBnn9efmhLdSkiR5UyYc/6r43Efx4Dc5Qw
RHE8xM81MCqu4l0c7EUE60DRMQZBh82VGOea9QsFN8wUdW5hpC4Zp3SOv4l6/MKG
O+CHAoLrzHYiLaQWY/e8Fbk+YqoTTYeEBk/vDEzeTSqSFL/agJjpJBIxOUQcHxy4
D1f9vPhmau5v+MfLQjIhc237uklR53/vdfxeWZy6kJNokacEkrNBdQMVNQWfMc1m
SPf3L8+8RhEXU4myhbr7q54Fi8iS69RY0n1aaRZuhJEq0MCVxy5SI3mxJwM3ZYTk
Qh0NH47RA1Iz+enDSceEp5wKEV2xs8xIiWYH/iwXoEZDZOYShgGP+FpOzUGqAoVQ
M2/RBGijeN53jxsl4+VKFipvfbXTFXf+/qYsMjCsxC6NPn3+fIRp/5Ea8bhLrkqi
oAkFhmAIxPAAZkA4cud7I1HgjsUWWW35jFjILgJWDL8c04TqXMlZwmb1RxCBgnwc
DHwI8mtQ6bEuPN6u5vzixQ/6sE29YGY0J72aY/2eKrzj2YOLQPXKw4EbRNLNTLy2
HLPU/2Rt1RYMn/5oDB5ive7F5W0Q+6YlDOdPJSBTxIkkdn+znyoULnSsfJu2k/KC
xUW4mj951xXVUNWf3wja2lVw93dhbWmH71zYUqdGHpOlPn40E0BoxAzzXrA7Oss6
9k9wnIQIcHh+fjUbFJM2VM3FZ0wmIohzc/26ZwObV8U1SnefRbjavOsugSSukGOf
ggAddCCUyJmt/1wWvS9kvxmhEVkkOaQT3SFshm0zR40AHMHjfhjnW54KiVhF7rgB
1SQ4EB4kLh/lLyvk3wOLMKKEjSKh59hB1BcbhDrmZ38rHcD1DgBa8P+qPemR0p7b
zvN/RKFtqwkVFEt9kaU1PJFwsvNZBMjDR5S31aRc5ss/Cn/9dXo2K5cvLIinGyWB
QIgxuMkEdxbxK3txF2EY50gx81cWMy6/SR4AXf7vrFLzbT3w0d1uYHr0AFfmi6fE
YVn94d53AvI6FqVly4749YBp5+39ISCrGq7bnzU5IMZH8vhpKCN7E1fJ2cLceD/n
HyoBtRSmq8W3v0NeCzAZedrqTVgpzUXLyQZuK5u0G6STwovhnTl3HpBRigtfB4yK
/5hs50L394hz0eYlBrGrOsIBjlzUEjssSjf5H48qP6QqSHkoSmd5WWpr6ZO5ZrTp
JHP98AEgJS8u3CUZhbOvJUZefmd4IDeGDTeQmbuj2mJMj+LBWRJz4W7C9qDi9uNw
/Z5VBKR3Sv7cd3z79MOy2PPScrm/5U4R9SSuWHHP+C7keBCAk2eSDICUDbS29A4C
p/AcB9LkOW7vLqFHqrcKACfWWq2GHGzZGUPNCDeUzyXHpGx7d57/twDIV9+UKhDe
5Q20hMXB8VBDb32bE2Nc1VzG0KjIcI1TE7FybNCsD3sIpjTx9ML9NLX72cl9SRqc
8XsD/iOlwxWHEl9Spaxov7RxnpXlecA9JiKGA+hWEjKY1FYIXafLRHhUzOSvxPgG
K2z61oRDJHzYFNIULI8Rh560u7UEho4r6B69lfWWY7519Ob9DnrebM5NmRoNxUvO
YRnfVP/+7nKNDrkCBIeUUiHcTSkXJZsqzotJ+IOcoDoT1R6NUhNJBuGEPit7znta
u/kEWJZ/U+8/lA9CShWdYSP7Of0T5bm3udczzTZTkVv9ZmW4/ilNLZiySZIq+Kl5
lVgK3Gcg+lYP0XeQrPE7ySzEUd+QOyGITdrwPSuqQn4jx1D0DV7g6nYxTx/mu1eY
NZakson5W+lwRvXwzSI3SAlfqiTqnP4BqD/7/hEUwfaTCw86/cvdzbJH67rzttd2
YfQq+JM5GEdXc63ZSUAiyKk/ex5zIWRXgeyNXy3O/5Wb8YsqcOoy2vU5teqbTj1y
yWh71vfevHPKwWTpYrZHVJWLSsUmf0PZRIj4RXNC9xZ9Ot5SVrjWACv2czBg8Kn/
eoMsg4XnX8SkDkW4c2yGtl4Mp1ffBUwZuj51KLKQTox5+pz29VYtwl/1hfDhaJBK
7zmu9mHn8jvPN7oce3SakBqGIsJDqsQKJIhLXZujEwmuMjkBr/q8o83Wt1KExtjG
HZRUNmpb2L5EDHXiTte+yWSjS+CZ6Jm2EcOU7h4zg0znWd9OKo7sFW6A17/Oad9q
/mlw/+dIiJeoE1bCEk/z2xtsoDjcUjokFlEE/JJG2gAqz8jh9l5rsNWMZ6zkqtE2
cfRy3LGWySG2Sf1/ssofx1Xudz4zHjddGDAv0YtXmgEWxOMso2nfY3Vh32n+jqHi
11+yfuibX6nQFEK2BzX+bFx8K/hrbRZJVXP3Np7HN1zJY+wW6IdzGFgpHuFu3MFu
C70ixey56AHfoDCc8XrT4ADyyj1howR4BJ7cbeup9P61vOEqoG+yMv0lAA9pS+KU
8CJ2whDtRKAFhNabzqk3RPIsPDnTEWd4KYFWVRlmRtgQRpLLno6AKXJtQdeo6VjJ
1H3YkjoqZ2+W/U8Zmqj88yrBEWwkbLIQG3F1+wgk54stTsgv/85YPIPL6SlbCBk8
CQpm5wBFWq9AyXgEtL9RJY0dwbc355YhXJ1rDdOQPmgsO/BamSuswAE/l2WWF6LH
0e8MuXbJanjBMRgkAH+p7Ac3+te7BY/4/iygLxaEMX6q0+Fjnb4CNyKXOXmmyMMq
ZXf9tMnR6wV4Q6BwqbIHK+rsnN9f0NThzymnrrun5tBMs3+R9fLlQ5PfZTVA4RS0
itVmPHgbXQjOM1dUIHzC/VGCm+TJ53O8ANA/4J/9gW6EYAwLPIBdPohriXIEYAJT
w5GI/y2R2wJZnnYCtTcL7RWlbIeA5HTPZfIYQeqCWN5FW7bISxRi4N3dyxO/LDRA
Un3aYKn6XcC9ntJ9PynpdrgH+7zcoSryoTz/NHFq2uCNAmLT8ZUWFGtey01mKATe
gm032Km8KaVilwNL5ER+GQTgWSXueClY5MHApShWV8V1Da4gQDhK1FLARZZfyrmu
OJpkzYX+2Dzi2ky0WMaKhXYmw4Gx3iW7/PQsDmaiVYLldrlmCcwCuGrU6fEvKskl
3xl8GfE31I1yvXtabzEhPSvl3HA9on459OzBBzks6f6Dub25v0GGwgyRLt4Etv3F
iFLlYh1d1tYIYD2qDlDTW/wq5rvzYWuU3f6rpe6tr+CQBAJw9UZ3dEJJy+wLETjv
hwRQFJSwzqXc5rsVVzX9NR92TA75UvcWyY7EzeEe0zQfTE/akOQ3hfNxFGukGScN
kdnXZR0VeRt9OBrBofPh1x2IGmYefyXKImmq69vkRMp2xyvGpmwDqegHQDm+AxjT
yKZrtIEEFdvQuASTRWiiobY/39tfHEmgvUeCnlvSFka4FpttHieKKsaC76kfSFaA
ZkjFSQ+tOoyPViVUvlBZT11OkSE+TKsyfFQh2XyO1dkI1miIfAUfKw+sCQawVJtW
Zxif2QHhjvmrOnYXH392iTpRQrE5AQJD2Rk2TI9wgetoDhOjOCrPt5GW50WuLe0z
KCNkvraXDjuEmMOISj/826TwWijJDosf0nL00s1mZ1CgxkotNNYZRlKGj6G1vHLf
Sgatd0CDWdEMSa+DdXneNG8ttAhd60aHswKCoVIB+wijbcZVB0jViMAw7gsG2MnF
Zz48N6OHbvqAfUjKVM6KeqDQzsiA9OJL5PES8XTWDXJ9kEUn+KRpQ4X861YlhWla
lZ0rNFWD+NexUFK/GrlPPYFdQ/ab1iHmniMQQj3JC0qWcCZ7MsSqUD5zfgYtmguU
YzOHWyWw7rWuUz3vjyaveYHhuns8qdCmumh7cZE4Ba+dkAOD1+1NxiLUsDzVO633
qnwi11y8Ijvw5fikcXEuM0VdcRPxIzn/kvPKb0EfDGuMUHyjXOL3jpmbm4VoNw07
QNqSAVKDzQphoi1Ii6BlGjj9y32Q7lt6CJExxZO+UaWnchMOT/Zk8yDZlZIzXDgs
0mMak3tQzaZWUnIUZ54ocyytq0AXZhrm8RwJAZ8ko9gOMXBBAr3xpnsbtP9IoXbn
uaCQyXT0CzthvvKNeuBfj210s7hTUz2VqPEXrnCQk6FwSK419UjrjKRNIzvbRU3c
i9CH9Tli2QL535Q4ULbxBo5nwad1P3T9cXnvzP1mECTLbl6b4yHvapwyafLSXvjZ
bIy7Sdi9Pc/SbHJdlJxYlVj3q19P8qcT+qRF1n9HdoqhaWqGZwciIv3gIopjkRhi
ZmaT8duvDfKf74qseX+n7Lg8aE2CNGkvQYRmDgvY+zm9VzGEr9Zxyz7soz7ykcNz
fIII5B4s+sPqMMfGP26tiMlzXmPScmhQa2UJmQcIZezu+QE0lUzP/ucJNeW+vQV4
2os6jXzsBpGizMwWLvzSoWUpIbiW7A0sCcNdXyJZwLlRnkvOHEoPzMZl577zPa1D
8j6M3VfPqOpfMd5mtaleU/fsFPjfRcnFB7yuQCHcbnn7EzoGHndLnBi9lxTlsOKt
mcYHLfK89PWzKmx/s8/jovWpkvvUQhp2z2Wf8gm1+7/JI5Ce8ziTARqAZmZBWanz
a2A7wYYe5+AhWH9iXO4PxPVev3ol3Zh+pXDON5ehowCEXpLUQ2QGIIIEB1CIgus7
Pqo3qSvxBvJiWsQqFv3ALS9j9ixzvFaXnAyeswCDQXO3KCwmkwPEgW0eQj4i+WRX
w5qssZl3iKX9ZELLBkZrO6vixdBHUVGlPj+/ucJSLAJemmzO3Fdb3u7ozb+OzSWE
6P77qGxVMijQeIXkGfF6LwPIlyxpl2LNh6d0mtEPHAEMKcNEymENW/WJiodwM9NP
Yqqap8yn0E3aXWSJA7rUYmVsLUR6wAu/aOtTxJQzH+18Ri2+UvS8eBi8AJ+Tfs40
rspVBR4sAKbZFtl7XAHQ3xeGFEjG34lbj+HyZcMneVmB1m024J6Ve6WhEnzSyhC+
avM9qOXj0Br2enrxej/ZBfvf+EYHPRNqJYekQeQN2c+7H3ml9RVp5NAnuU+IFLJP
tDegv8+HpWnLNE3FVWoy/Xxu1ndufaK1HZygLppgplbp8sNfHNgE7mIAAPDqQ7bo
gBib6ZrgzCPq79CpByWHXmwF8f3JT4glp06tBZk89P/SVxb4SuCRdDrvYMk5mFuC
O4AoF4nq0upZ75j29Q79L7lSMZuipVLDLfFMxa/JcTRY/8WqyDQVTc/etnxHLOz1
1pp/G0+kie8zABRdWuJ+bpniRuv5qqRaqKS31LLJ4tZUapBS+aUAdwfJHSjdCRlH
mAqJgwkOD+gHPGK7i/IPmaTRoRuhrRTXQWZ8ouylhZm2PekXIn442kCABswxNtcp
7m0shKdZg7UYZHAv2+rnWwo5n7rJwdJisP9R2sx8PTrcz19wjjulyArbBlpuJceC
d8KVYYV9+kNtEqykO9a01F28rpRvwK9f3QAhoiNwpDxEVODpntJUR/L1e8hLyzfr
VDdVhgaLVBW3OsNGL0Mzy8pgAzfMVbfV5Ok+ENl7q0Rut32xz5XCriLslUB6kZSw
gku0sUffDkViC9LeyooLtkWXIgUeWUABWlD4ie1CHEFmW0DmsEM4pB3R9M2x1ikP
9yZdFt5GS9DxN3eEYDAxs6vDq1P/fYHgX7YWWUnplrR9IM1IypuiwZ98pmoLI5zj
JWbGws3HSWt/a0auKRIS1e3Mg23OLA7F0LWntyUKtESTnYy5Jn8UFsALhlo2WsGI
ROGFh2CTJ963Zrzx3tW+5Q/9I9kzj5FKZvXcjRETl87MZsHuLUvJKXD/DkUQjOds
VS3ZjHpAnf2nidwF3IeAHhpivfK/JN72ZVbxZGLc1KCphLrmbigzuzmNL7LLGzB3
hs9TgudiMk38yScGrf3KLTzO7di0UtzTFPScukRS97HLfRS14q2aw9uVESqS+tk4
TvC+A35e+XVVMg+YyvnhyaXnbUVb7M6RAnTrv7GltEr30lsI0Fywi3sYqOt2elSF
ARsrQGzds9RhWf8/ALkLEuHfoxZvXhOLaBqC/lyhjGNNRpsCe/J7OJes9jfRl6bP
Ibh964dnJCFFgnSOu0pUupCZ7ANzQpB12eglGobKWdIssYnD/zSwbupAq0Sv7jzj
VMbnH4exdB84pVi0HuBv0KTjw4JzbgqEmWc9mL2MzBZXohzVrCJOvNJ/JNIxYCnq
K/+lZT/T0gjgIZ+ZqFU/96y2Rm2cjkBmv21c+1wigA1HP68CFumk4R/u/o/0ToR7
oUgDosEuSNrQqL7YIfZ5k92dKxFWwBzr2KtsGTPH2Gzrj3VssFMBjc/RSpZpEOwg
mhNiOrAEGe4cUnsSsBsGIxLn3LUGwIj5WsMiE1ms4jI2pQ8BsiOW0WudiPG1LYtd
AHiQ3dwdF7EUNo4tI25RO7igFPR4LNr7cDub8PHrFsGABTvMf63QIL8mkEiImzwH
eAtMiX1QlnDWfrkWaTIJ53wdc7acGIFRQQxLTOykTplhQvhnJmJz30YB8XS22cXN
2vOndvinsLVQUy6zDLVNHfDs6FTDXPJ4TIta/F+QGDKbMfmQuoEpOm5FhSq0g6Ak
Ofy4+QP1/m3MeR8Cs51c3rGJ3DqCeyWhDADLZEPSO9VTOn6ih1pSlgRtl0i6mAwP
2tAV3avqPyEqRwegY9O7L8jsmIfU9NXhhlBC/vo96945J9D0FRRXWI7RNRX8xpB+
Vd1AOC9QbQGZqz4JuA8PFYXyyqX1KAL4SqULzIRlGU7I3ieN4klrMt+9kOe8bIt6
UjzDUNTYVoKp02PFlwDCfqFgFCPKonZIZ2byyuAIr5famEaOOvYQCAU5OUtFyP6U
wvt/zEM3+W9nZmIxuZzL/zAf4i7zA2qlHfnwvCep0zkCeSiACA8sYjkBY05Gbnh6
JdtJUpeItCGquB2YYSXYxrX/xYPVvuJx4MyMJc0NuklpOthYzmiDTQbThD3TUbsC
n5e8cF9DGgiGqNgrSYQT6Y1JPZIFvhYxzhInrRqX3uhpwtwrKFIZPK3+didvbTH8
og3aSinqwtGx84M85jUGFSE7s/9bjXI/un2wgY5xaw7bI59YryqKViYMm+MjT71w
KKcgOnk2w6lqQkx8GWXRJFryc2Ij/sobmVVAIJFsg68bNL0BwLV+sMTSWhTCNLQW
i2gaPbr1HEaRpYaEG9ggAuxkEqK5RRizQrg3poCgA/3hgrXHIfK4fqYhFfqH3aZ9
0klJCO7rlDdG3B3k/us1fLpbg+etnT11F3oqw/UlMwAOqhF3Gzrw0jgVoO0X/XOf
cnLPyFEiJ9XDgzvbHdvdDkddsdeY6TRfKlH3yCBzp1jB3ORu2DXTfvwq5yNhAWdB
on0VcySiGxWV0JsJnr0ofZ3oEcHOZAYca2c/DtDUJOrau4yfNaeIYHhjvfVQK9Ic
am4EQdEgglSGMU2PNAqokfxK+sBW6UC9liZNShxYJW9oJdO/4amix4YHO+gwJXOQ
HQTLfgTtOEts/LF3G+ylFWcHKyZ8hqEhIqDJxCrE5eEDfGJqPq9s81kFw20Ubne4
R023q39hU1AdXxSWgHzZ85k1sLMi8Im0abQY111XgSQU5cwIN5wfZY21OWQR+CDq
4hgq0HEP5TeXMkiS+QdoUuh/wlqYcM1nKIM1TEuvULPAMsLNOkGWUzZdAkVHhL7z
3vU3TNTyJo7zyRM9D0Aa12edGr5Iu3xMabU7mw7Qcx1ztZ5jfXnwlrDFCAJlwmfh
QfFK/njoW6TiQfvaO6O9EXB1V/rS/P5Ux9l0d5z2gwBziBG4Wi1KJAWQljEeL3ys
Bzh4YN2SBp/6pMvaJAD7owxF90YhzSIqb8tnMManmNUa2VHNeTgTG2eCcNPfunz3
qizCHuvfCNFjoiEwLY+XVw4vL4f+q5TV9g0+jvRAXSZIden3tF4hhXwR1KEuBHQE
MxSZR3zmhr5L20sSvbpz0Vg5muPYSgoPHkylISW56cBzJ2evF+SoX4eY5VOgewmd
SeBJVpv7cS9iKdwk/mPIpLSB7qjraLDqCReOv1KeLOK1tvAGdnwQ1cKEQZ+O+XMy
gSCExcw7eMIXVv3s6Piae7fDBPvZ2trkk5mintzpaXqh99hRQ1HZ7c2b2rCdl35j
61K5tVgYzyEWUC0UzmpCCjmfb20/VOBz39iZLV595DUQbeRrIxKrdrZLe75zH0g7
nBqSqfiI0u+tVTplq54WABEnJ2nRwruFCmSEjBA567vXzu2LjWyufFcceYQjyqjW
YcCP/wRp930grCIMKIal33WTLCHBRpYo0xmIZbGqdLxKsS0ofnlipi/6NatJKY5N
umlU6e70LGgXO+lGA4HlqGnF1xWM3aBudssWcmm5F5jed4lfRFxEOorulWqljtFI
f2k3rOasZaBppGZG6E/Fke2sz+l4A1DLxltVQ6Jepf45kx+RsNZHPWqF4/B255RS
xRj6sw24Dp454COWN3e367ue8Z90r7kBn/6e+Mzmoozs++YUHFYj0ftjZ+FCoAlQ
iGO8Vsx1IFTmopVHcyufgEJsn8WFeZiCdaZX/5o+TvTRnIp/9PeRn+QJqVlVBLMa
1z1mxzZ4ekPqkwoOvg/uO7ax/TggIuEAsTSA5ZioJSuhZ6/tu/Z2h67nm75685XQ
xL/4wSt1Jq78NB4y2usFiYtXNhjYPi5oS/cbXXL5pCAcnMGMyZ1/TmnzmoCTy6dg
p2UMgK9buYae14L5ibuyHiQthu2eDr8eLr+jExCNxTdOgXrFzourmaI/L6ROyfnq
el6eSL6PcVbcweygRsDLqyN+iaA/cR0YWno/pN+xIi05knXSFt5If6w8r6TjnXwn
gYWxj1oALppZfMpyFu8O39UU/MA04P17AWfVDrC+lwIU96i8NQ3mmYnejwaHYVlY
SmuI+jFwKmJfElWS243TnvjpzezhN/QxVkYAVn1wFqtL3Z46Nq2XcXDNCpdke10w
rYCRpUdqCZMSk23iJRkoYD9vO2dVDiaKEAnyc51k8/ukfc56r6osvPb+V+jbYhP+
g7OguqJMjLi9UqMsTLZEIhj+FjaTXhnT4v1b1gtDtJyKGGhYAJ/OMb0myccFDAeM
tlLBNVibZaDZTZAvt+kEcWU2wJInabN3ZaDOb/2YdXG+tTZnPK7ZQASVt0asOoBj
PrQgMPhCD47zJReHM8OtOJeI/NU7+8EgQv4ILZcyDGnXOQSGuPtB16PPsQuk1Lfj
eLGpP++RR1yMjY4j4hz9S5NQNJRjPH8e2h+Z2UyNwGI+uQdx2t5SPz5/Aa9m4sbJ
jGMTrsuCXgJ5i3B+Sz7b/RkO2nvDGHjo2MwmxdqYBPD8m4LJIBlG8Lhi2WxR9c7G
KvNZIk7rBpS3h741wVKhF8hFLWRosXmbY2Gsm4qDwEoKoqVAPy+PQFWHbET/HQEw
gt5DltU6NRhvKjHwTjL8o3NH4t0C5hMymZ/kO3FWT3WqDXOjKVO359XuWyPoHbYw
RP+t4qJU6fxxG7g7U9XA7+Lx8espmIQdy/3YLiRHuHpR6/UZATXV8T91Ebs/O5eh
SMB6aPvJt3aUypUuD1jwiUcI7WQ+ois5i3IsjYF3TbsPEc/561qN1Vx6AKjPQG4/
BheWT0ETv3fw9xZu5N621K6NV4GP/K+hc6BxSeOk2yVRg2kJpJUmD4Bg0ETUKFml
mex2eenipS2kC6p+tfxLsUFPC07PomEpgJk1crmAnpjxPAxsZJ+7p+PuNNh6exS3
55O+s2WaLE945UsIicQ+s0DWrCRy3G0EZIjPNztof5cXWz1vm/BSXt0+dYiiLaIj
gV8wbtQVXvbkPFsIoBeurGWcxEe/YgqKO+Tqs68DnoYgWUugTHDcGaGmlBEDjhlD
UM8uEYj0tLzl0wKi7uk1gNC9H7UG0CMGMSdWFkDeou/wqZsIIMmdMTemP4+mSfEg
kA4AQ9dA5tPBuOdQklCbh/n2dSj2zKNBBoT746J/S8I/+OK771DqvpYNHRPuy5Zb
gy7Ty3zW7FKe9ebx2+IYeSD0qyXPBETTRkhExlyPyXZzQqsgElKhSp3+q8QN53Lg
WpMGMxWY6j/vRQ+0+rWnCm4fW7qwGTc0T9ggA8sQ1JYGW8bmFl2sliz70EjH33iJ
KRi/Tf+UZqsUXtm3ZvG8AEPWQjeVu8JKheIeJnNUhu4LkHOphNHzLMca5M+hq3fR
zZBOobnJUpbM+hLJ5skumfg8B63thJXCIjbLzemhqg/G4YTvsKsh0FARC0NAN2xX
3Sa9SO+RnDqT65WjO3EVnKs86g2lBrcZmEmXPOhPixcFi0XwgDGkEkTLVUYTpQWp
swT5mfeuaqkByEHbQ982j3eP9+gWKwnQDeloGPVRvr6Fc3jEgNC7zvBOMPDYVUNK
py0T0TowmIJ0UTZS+88oeMC732j6aWT7s4eQXjkYpYHF9AuEgz6QYo12NbVefWXp
P46PjZKPcCcXCpgpvb3YufurSpqqBUwgZV3JuOKcFwiDJSBmJQf8akHlWywB0D+i
2FKQK1GyzC81K9BJhpThW0LsRtMUVBppuFHSf5/FhK45csVBel+nKhHhQGjoMj3u
M824PpmYbr91IID80RugJ8uGDSFN3ltTHpJWhSBejSeLxA+Zi9gcTLMo2ZNzHJuV
nj2wRM+8msysusAQmUBjNywL6suw2s1cV6Ii98Y52fQMGFyFZBof07ewiaUI26Gd
1Px2S2I5wd6L5gmuFZA4Jerpv6XXsumWi6D8m1pzU9PA3mP6LHz91y0HHpqXgE2/
fjNLlMcW1zj02tMN6Wi4NNoR74p5ZO+1bxMnDfNjzAorRinnzCqufsCM6z9YxJgx
Cp3XdZk22ZWIlaoUXSgQzGpW2dQJD0eeDExLhInYs8z8EwZPJOMKVvtMsSR5WssW
gl2XOIZd81Ej/l6niuRPeY/5i1R6yzr37EpDENE8WsnV1ODM5VmwLijucU4QtnqS
9bK/etYrAahbU63I+Q4S4QPJVWxrix54YkqmZH5HyK1jCPPcrbiRs/V81yBJkPnS
Zmw7ynsGQ6XhVFyxmVgSFVRez+3yl6n+qnKmpFQG9mjSyZUAKOBCM/PnyAzL0DBn
rmkE0JIpd8WbaEyp4iEc47yJZxyFuKvi34wBfPlo1xHdHeDQgNl0zxLl+45yFj41
3Fjgjss+xCSKs1cO531GVF4ho1MRVmufyUZsjnJOeMxgISxT0i5K6TlMNIxiWl9l
v3Ave2ssJqYjEmFurry4/pOqGBIdbKxN5XQCnQES3XZlW9tpDzsPe4JKSdBdOytH
ysvcHKRIkFu6pI4luS/kQJ0y0uf7PyFPgBPDUkzyHKjQoEulVnS8iLRAZxdqsapa
DVsHxd5LpRIaaQ1wmbepeFv+6/Tch+0GzhiVqcqJf13RXz5Tgsk/Xolc1p9292sn
LychUtN3AMIKhxqfR/4hSvRFQ0CdOxZwwdv2lST1Uz753RI/ifLZsBLRQEInawy+
nNPLd+Euctkdcz4TCIbsNNH27d7Q0GH347cYonBZcZlYYBVuFpPSayBYbvdH0rRy
cXQ7Phk0aPl1xLCVbaK+/qVMc9Udn5eTrium62O/CHU7X46phOC4LXoxRckLjZhK
iHWuhcpHMD6SHGlEhgpUxHqF7ht5wLmGc0fMnR9QGg3i0skidwcYpxZ83EcCBPlt
PAs+/oBuG7klgqWLWA+OFWNkNPO+HlJ+sFVSDSVVhf4yVKjkgBkvg82vNMr4TAvT
Nk4Sx/lwzuxmoz7UZQLgwTLn3Fq1xlX8BbFNpDanZZWZNns4g3KKWIkMCc2ACFvY
AVDeNmvaoq8hN19dLjv4/+fN86wVL8tUVP+fk0aV0IYa3BRP9V+H8LlGpoalUmDm
sQdbIiPQcGg5hSZCSfnsWLD5M61NXpNTQLPceRcz9Vrv2Nyxu+Jz07eT1YAkDtI8
IZoqvTR6sfLWaTOSiogf2S7SP3QLoUnceyJSglYe16YbTTh0f0GFDvtx5TpT1G5u
aD4RrPq6jG8UbuPxr78VywlcAHKzGzLv2tQQOyyyxT4htgzsW0/TZ5YaLb91a1hb
GmUnvKDNykKfIo0paYcJBFjsfKq3R2OL4F32nXn0u40of9w/166WOT3tUzfS0KhY
n9cIOx/kXVQC7lVncSABzWwodlOZhHqN/9GSyLokQBkNif3rYF2/pCud3Xnbu5cS
x/0c6ifGyglnGXLamcGOaewV7sJijsCICuThVzXV346rYmKKse+Wrng4+4YT9qzK
EcgZ/VCmNam2+kauDsVtxQbX7hIsBYCMeNzcoM59Q3uEZfUmqLVq6QUdaZvxYNAO
Ew1+rZvJuo12SJq9wqnPwdvbZa2wkXdB6hcRem7+nor9Y+Tbe71s0YRIn64S+lM4
fX6yoNnIuFo/ssDKv7Q4SUzHB9b3OoCprl2odRojExN4OrJPiMMJaW5GzLDNxLdf
8DFFJTlIGCNWRz7dxwJPLSHTR/kT4Ua6TgVWkhydqUOkFxGnAbK1dsjy2RDngpNR
V9u2hXGXXwxabAznosfX/PjWUDvJi7TnEwSUe1iDrssY/xU7ALSpUrewywU2zW34
CJI52AB/q63Nza+sei9SEzaf4tGGR5WHKqvf7bueVDr1TJlkM1Gv+qNOexSLbThm
GUn7noXOmeI/ZKKjgh3RMEuhDJ2YIXyx7mWkjwBCqriEl/bGByRh1reJAiv7Ub+J
6XKCjaHirGFEvA5VLwNqPDuV/0rH7QuAnwaSzd/tslgzvze67ZjwHSPjof3pHTG9
KPRcvXnlQL/Dhii46iRzC1Q1syHj97IOi6ka/GvjE9T3jpTcwV01rD8B6ksBFSnX
CRkRhfdrn8mGqPiBEnNg4JfJySy//b/T0A1IshXR07h0BDdU53R5LBS1/WJF+hox
1e2gepa0UtamtlIrxnDrG3Z3sJ4oJ5F4p4uvGdyq7sk1dPtw98VJR3druqby20vo
pBhXFkma1EL/1ENuSLmNmc2yruhaDwZ2u9f8zRTn41KroZ7+gatxX2GGjrZToMny
65ur5thmXvB/LRdC79XzhWgRXSzJ1+q5sBjOpYlgA6plmIgEd7pbvZyGN3Tacl54
XNQVxwpkhgfsG7wbAApPEXh1gqcVjyxldhyrnvD3E0Wf1k46ZeCdzfTO2Te40CXx
KtgGOYwVBUgzQdEeC5rL9LlzDLCiNAtmU0vur36pw34uOSm/cLOQ93GZX6E9fqDt
XZwm+xXrymDqQkd9sgNkrDrOJKMYqOkBoig4ZTQziIwpt8Fw/Rinj6FQ0jVX9+Qm
Bmamwj1jXxnSsi8VtEihYDIs13dBtXIOZJP9UMIfqKC3okShA66vQhLtXHBBHFzZ
QYmBNub4yD8Skq+5N75Ay3DIGKKINzDZmndIK5/awwNTAE3MiVZ/vqg2Daw7IEsu
8X04vhVF2ImRYdTkQWKsMskn72NG2kSTac+uQ+xqcl8xaUuJmFWcXx8h5DA9In8+
lyYNqGuA8zy3FIgWBTuI7tW63/3Vw9V0w8zB9XUPGvAsdMEattHcAAVu/ZdChrnv
RMIPQSKXnBpmuL2HglPP62QX75Zb6YGNqLIDCTf1uZQDxERjwWP/RTNccPf40vDa
Pi3AZhMnB+0GIVvtXe3K3kMvOfn6GUICnyxr7zwmOAyoDi2vcUHChqZZfoVdehQy
mi0Mu4r37cGJ+VNydNm+/hrXBqcCcTjMfnHIIcEuJyKp/ZhYLZWq3uWcYr5MXCoM
Cvywe+l7Avv7ZON9EaH1IwSW6B6w78JmQVZmXCFTVP+mFVhglQazuHDqXcjXSMrm
va7fnVKNqSxiHTLVoKwfI/OTnroPPJiNenlNBaRDCyhFZflQhdQpO5krVCzAwL2x
SxOpMKOUeIA70WpJ8v8uJS2qb5lUgVxYBYIc35XQKh1FttXzwPMYofebV5z55WWo
6E8PXKu2gwI7U2lTksUc3lNY4XfTVBN0e1ttoUKtO1ONrna4r7GdKAKjZUrdFmT1
RL9QClsshUzvKzsE6jpzslHpOxGqXcVZ03lTPgNM7uJl4dYqPilZp1gmoOUPAMiy
PlxL65naF53kPW0/ehieTGUJ7z5UXKJiG/Dme8GBnR45uod9tkkdZ6+qTErA3oqC
dNqooqh/uZa1qYttg5VBNarrPZCE264NwkuNB2ZaeTrd38RWwBu7BOuPUK4j3z0h
SRpYUpeTtTItkNP7421BuBFRxQJxaNDNpLe/5B/DNbltrGbKBLieJvkgfBNf2OGC
A27EJKGq0/idzK+Zplt1xjcfOl0Fo4eYqG3qZTEftoUukMnitzQLd6lL5+DvxH8Y
2ksnEbZSGQcIJ6dboCq5Y+yaigeAk1XT0wvi0g6keaMaEOQcMrvz6vslV/jPYqFD
9YF1QE79UmKL0xBSdlF3BdhuHUA5zEYknisb4jHtg0v2EZqeaNRZpRN54KyNcACQ
PRG7BDwYK6OrswbDwQFvWVy5kNQ0Wtmd0TgJGkDRooqrFrQs4EpQo51DmNaB3pWZ
ILtiWEfJhqo3DaXTO6e8A4PRuvVGoOlVBNoVkKSGk4g3j+f7JG+4JoZoBR1pKVes
pcgJ6JCgZpxSUxtDmR7fPAODW/bwPNPMkizGZCsmUQxALwKhYmXfWJEkl7m7BuNs
GSlNG9lCXa3/XGUVJ/ONAvFvhFCdtZ0tTtwheLD0N4tAq51c0cPzTXyukCgmOZ/C
nLyOcSwETrl/zghoUivrCsY+2Jr5MeaHgV1hBr/hwPobnJb3R2EjJ9bg6b7tWC7N
AD3szzUrbV1XapbrwXg5YFQfgDQyz69zvlyb4Cn7L4WuSsKqNpWwdt7W8rAAHgdB
XIhoOIVq9hx4QECS+Rq4909xWfOxDyAPRXllr9/jkVM78ln7D6xBR8B3qbcL8YFi
BJhaJURsDZfXNDupcgi50Wc2TvcR2KP8qdZ502+B93FSgH36/TVWepNJJpOTTT3d
drlKoRshdaiz6jVZm86dLy6caNwvYO/n4uzdvKDx6l9x5TXrCr5yK+0spmGp+LLO
bmdkhGGHrorM/cAkrbdCesl2xAEa+fL5t4EoRZWgsSEXTbt7LcsMsWdRF4q1ck+5
BeZwsXiwqOP26VCCXQmOGcGQC0jdX1x7odCxS9TG43PBieOEnjp5Ov35mkoiOQ5d
8Y8REozH9G6bjlPDAX+j3k97JPVmIxS3svFlyqr4Cr381BAquSSFR3HLGa4uj2PK
XfCaTnAjdORxNrEC6/DfPTi0BktGgbeW6lqE+Ncv0V55VIbD3K9byFllafMoShaG
9ZvNAIC9sbAbkYcZbH2Ttg/Y+H2j3G+VHzdRJFklYMyqO7gP8A0DIG4yCy4L+D6h
/hhqNzYL4naSxX1lMjFRyuo+UBMBK3aXypHiTTxyX3sW82SKVdOBUb6nouCO/cZd
uIAy3tjC35s18/qWCHnGfsmUo7KAeaItpYO06fYjaDYVuxNTMGbeQ1y6QGHC6HYp
UJ+sk241a/UUEWfk9klL+PYkNpmp//wUDlKJor7ZbhhxgJBdv9ofPqJeUL7lGcw+
SVbE59zNJsKiu2+dAfjTFXGi3ThxsHsx77K3Of3AqkeAeF+BBCPPbf2S1v4Tmj3P
zPV3B/2Glnu6VjGUgRL7waPX+8KlEwRpcQHghXmRsNGFDevXvMYmZLQb54qaNtQx
jestWJWFhtRxQDrByfQiOIZsapOO5GDohs4SyQtwD+2P6TJIMrQHFn6n5P19ru0q
iPnLIW/HS8lqi1ojPMxc4jDvK7Up3f+87jb2p4yOjuEcxXFwUmcH0yWQ2nVgL8zy
KlXLUbYIcyuybqbcUqnAZOJotB3tAUkfDv1TExm+Ww3pWYdV5ZvAKA7FhWgb/U1w
AgQrkv9uLS4Yf/KpFdqGoYwjo46OG/7nkpNV0KRR+vizvuGptKjRl5y/2xpPuNGC
cghvQcxXv9XBnKvbZ0RuWJhXHk+Pp5S0AAnbeYBtc2v8oKCAqXVv0+TTjV1FZb3M
MgK4zQ1KPz5jubtid1T/2DbhylycELN+AufqfyJrzIjEpMS9STme43PltC+zvRXK
IAelSIcMvkzwH6//xjke9f93mjC3ZV33wTTJ9ll5MKOXkb/pd9IeXaUk7cUqkpw+
1eXeCa3d+EfnmR+wsffpEScUckSIdZHd+CqGPfAsrdVmXa880IiKoLj7z/eBesNb
9AKoAOF6umQvohmre9RyN/5EZEwCT3R6MctN5WV2wiz+IiFxyLePw+U11+IG0blz
TVaGOnd+LNf3O2/A30msWr7EVZcPn5gejgB+c8E+VyFocItWBj9G52VEMCw5bsb3
JjiU14Lip6aoS9VA5330T6rCn5vLAQBLMk5fyQ5kFdfx7u0soorR3LXinSrxMMTu
/aKMnxdElIHLfFddfVLmWowFSmUevk8uOPjj2u1tL98zU8daefSxaDcV/n3A2Mxk
fGJrzy9KflgqFuS4X6AHmfpEqC1Le5EqFvuxY92Tybiq04iyKkykruXy3vs/HD5M
x2GmpBPFpuaDnNJf7oUdxGwPxxuYbsx1g3J8hEqTVrtn18Eh0qD+k9i3/bag6jua
7meVoVNfdwMn871tUT2mD/M0sp+sMxqMjq3AygB0/JoMvp91EH3cDZTSYtAX6jwp
LOeYfIS/fFykRNNBx2BQOJAESPfho6vv0J4RJVYLFN7qEwftq81eqO5lJyhaiWuo
CmW3uJxb487wp+zdyTXV2Ws4vl9whjwmQuFO8xvz+oLo5Fabsn2oSYmGnU4iah4Q
6TgmlrKxbGr2cRk+nUOShqWIfqoo0XIt5fwVQZ8ydT8ONFy5v0RS085A/4X2N1Ss
Gv753POWa98vmQWyMrojwBChswogNiO6xcw8RRuy4+svv52l/5eIZHBmpgcl0arG
/xTL5moLvHvQ6S+Aa7tQewCTWIPN62XBJ0oT8J7+ARBtZxzMuLnLkiRjzLTGxCLU
JzaEBY7/X1kV0bYlYTpvEW9/ci8eQWi+OJaWPOr+IExMGks57HSMldItK65qNcZ3
NUjCAjyZbPT2PiBJwWgMDz1R5uDKycU11XrF9dHU2xv4h32BnjZ8QdK59UCZSzZr
ZjPP0FTIeBhqiW33vRv2rEsvn+8PP3yiOGJEOsOhTsIiURFDnZyE+jf2UV4QhkQ0
NK6oFzVbgl86ZJbjeiEdaGzCbmqyBJRPoU2SkYqWjED02LBkCM1il2UP0G0uojiu
Zb8AEJGdVx7cmXvOhPGE/u++de9TDzdaJK/7e8YJG8rpWYKbN4SZvzdLTri42jw9
bLA/U/p5t7W4p6r9yJj+/dFb6E37pHcGHvr+T4yueDJb2LJe4JmlcyFioyzL873e
vRV33XhpMjd6tZTrhPSrqNyMS26GSxJj8P14qgW1bJyaR5ST8hoFzdrRPdY/h56T
8msoVptB9sLIJjJZksvdli/bnK1wVYUjXMEURGBVdD7Gj5r3LEAg9OY645VDbKDd
2tJEhnnNv85WVw+K1qUdSmGq45mDyICQ2dgutbZqzwOOGwdonB5qroFyNHbn3f90
7UPGCTY6VTVxGYAaF3CPJEnTwpwy6uk9EcFVq3VfUSSNunqNYUVLrncqOJ8+ifPE
sI5yD/mJgRVsZZn9I/asc7xAUbU555pudfo7ErqW5Lrid92tYeRKwDkVBGKqVW49
+p8a9Foq4HSohf4Yo6zs9iLe2yKTjjDLWk3ZtE6wGU2/XGZvrysIGD+r5WfWyUAF
dECIE7eFgUT3KSxsD1t8HQCb+qU3GwCYLrQMMca0ufo9qZTotUDF1yPrt2OM3EPp
YJ6DizlhglUaKjK7c7uCBUWkjrGa1X7wOzlyDDiccLBzmjjf7MGFyu4FLjmlvfFH
Wa2UnmLGZ9y+Rj4o4eJhHuZ1ydvujx9JsTFlQNdj1ITMQvEMtX9E13AHp952iTPQ
mloYIJKJJw1OAzxnCE7U+eoOJv9jc5QFdQbAXARuM1JDZtKTwkF5fWyMKrcMrUUL
bOcaGEv/pIG0Ryo89MLDMgdaSN2aDCyIm/uCNImqTwz94gMemfOQx8MkbcJnTujO
Z/UIh+VrxozvqiftW/ajkTpeIAIYjfuIWezxCiEMM4ewd8Wfrn9ldyvcUdgGiV0Z
o/q+hJcRbdUZUujai+yyqiiS6mZGXYPpumBOF6EJUWzLYhLs6m6m/fXV96PMlfBb
h4+8Js4/+dgGO1IoxxuNw80fiNrUEZ0A9PSJoqbQ6+Zr5TiTgINqv73ilxIkarPL
25H1JTTYEcjxfx/JT6OpcBJ1Fspe+LqTmjjt8ceCOdwWGuAqChmXBVm/Xgldx4Q8
zryFns0hM3TdDS+GizIk3ZfI3SoMvRfYRqNCybO5xWijtSpXnrbEspuTWe87KFnP
7Gg3P/O0/I39gXBNjId+NiM4FXAxyzS+oPPWjeYqTMzDvHfFDgRDI+pncWM9OxuO
lI3LwcyzNLc8M9MoCC2Wd1RyjdeX0kD02OPcCPUgURJx3hpkeRXGFKN1z9NUR4v+
PsL+PW9jpz/IGlDZZ6aQxLFo9QgnIb/HMgKXrcGWQj+UsZCiYlVuaPqeaSDay7M1
NjfdiAApDZteX4QxDf2VwUo8w2XcYfvdDfGbqBkqQ1rnQiCviDR0o4Zc8lRC7xrg
DaN49S5Bi8IrUzrsgP3Zz+mKAc85q3pNSIsn7t82ijkqqQ9qJDViZ0Oj1w1RYyDX
lVnAg5Uvx5+VfhzWkyOIjuBG5gj8evj3CikQ5gwWO5FsIIBCEOp8l1E4pVB/6M9S
dKKX6/tyT6Gtv5scZFdAp4ssx4zprj20FmpmFBhpTSd+Xoq4giL2Ky6XiHQ+fcRP
HvqbWVac8iuOJCqAYMTmwIH3M8UViXhsggROfqiLYBfOXOomiOLumRICUGVeUCv3
4UAzzbqtuo2olbZ9hLf14ZLDivcKqPnez5YQMRPmST01npFVuLEdTZC0HNIGGFt2
cTJlzt+NcmR8CTlF6s7HcHfXl0ymWLResvs7rwIsmzOexNnfDPdx/6pqE2m4zKez
/xxMcOxccXL04qaXj/NYDQzWoPoHVEbbq2zO6pz3xsiFdZHx+wfasS0hbPzhn1Fk
V13gMae7ccF4zSxH1msfOrUW0jOL9iNP7C0n1+PHVCDZE5R4co3AWtHNXxnZ3eHU
U+J0ziVfur2Eo/fetZpSvzKRAjtfJEKiaYQjc1RqcrQvEMbD21K5+WHxAfSDE9UF
LGRgKltNl1AZaAu+pubgbTjEwvLsLEYg9QrI6LfRy1UuufgCCRsoa+/og42oAQd3
bIHNzjKreUKZvjoE86R5Gp46wL/GFTC29v1cbXOCAorjy5C08AVzI5aC4WvpIils
K1ymdvVMlD6BIgiGbsyF3xO+TpxZlbfo91a5lVpI2Vt3FCsxdYLa72K2mOW91pd0
D/VvX4Ab1ZGuej0wDHKWUNyufo82c53YXKT/aTdYO7KjuGP2symZHUFefvzNJlwt
ir3KO9n9qtcAo0o9uLQ8TXDhngwOjD98tcWroSvclLALEKjuICYtNqY1eI/JyZZZ
wM8n62mw0dyzLNOqQy5LnawTwcmsPzCpfNKWi+rC1i8AOLj04nDv0cC0IkCzFozr
pPNmu46Pv+BmEg1YjNFX+dPDWHDDKCF+kp7me/HgbsT8Lmgoq5GnDL3ayk4q7Pgy
3QMAopBNVOYoX7UHjZDZGLt5x6/6lKCh5Vt/pwps8ZgyW7lEJjDA+I8g/KgcCVU/
TnoN5VA4mc2q1KAMopF5n1XprLYemE3cSAB//UJYN3blj+n6xs+QP6zvYae23jt7
FCDvxAWsKRb+B8oUh03tS/bYRh2XOVjk2IktCBx/8vb0rLwaEgyeGndxFRkEI2oP
dBxcUmgKNZJ8yTv8+jdll+V+BcLvRwB1qS/pBn0uOXGgBiCdZd19EMyyvl+woLvI
yzXFg0EXaO09hSHezelgu63Sj2zGbfWlGoXUBiLmhthpgmCHteSLlvzL+FVjj+tR
r0FbsAlbklb+0EXi9zIyfLvvLNo28WXW42ToK6BUBHNFwXyuhyq5WBahOUqUkB0g
NPoc2ImCN4uakTok4Fu+3c1dQXPtW7fgDATcStplN7IxQcMmW+7uro2dqkWQXTdi
/RaWC3iCLmXpT5p/aNR/mwR43WBodO3zQ8pOUFT3aPlQ89ubFTtPUT6DSgBjWLjY
R3KX3OOxyyRBs/EaWy89dQ0kPn2/AnStI0duEKAqTAGpGvPEjecOVn2Bj1Sf94Xf
DAwxmiTxl2SjI+A6eI2MBLgo/eZyJHFFRBm0Th/tuHJnC107bSRIDfE6+0ZGjbmp
RMNBQFmx6JoyvWVavX4lEWz9uot5wn9OGj1SuOV/J8znoz/5jEcwpmHHj7Thox1a
dlXmez8MTBllEqhMOLa6tHfr6PQJnZ5a1n3Go+DgQy/Cl+ZMUDGzGu3iGQ1QC1PH
YpR0PRLl8j4PO+w6DOANuNiDrUNf15WgLtTvmYv2Wk7VL6voIVh6QsnaLy7lH0+N
o7GKMCcUMet1JSR0EK/Zst7KM338tk+1v37CmZDeplREbtD9zJQKT6AqqwHxfZmj
MA2pXh2KY+nqtkrQmWfAMuv/6ecVO43B7lpzzcEl3RfgplBb1NmQza6llX4q6VpE
EXSw4EoF4fOj5mS86Hpduq+I1UaY7gw/82lTf69wbPXstJdmSF45Ewy6DYdWAw6d
Q3KGyfmpI1G+X8tGNRg7M1tsOBU+S2YK7FFu02DNTf1n3KKRK7GealeurNWsccye
WrjQwZ0OrHrubUJMc0W0a2F25zEuEF+HIa52Sj/XhWaZXL59Gedy3Bzn0dH/CYh8
tX7NsGhY85xZaOJAtNzsGEhmVMuOlMb0HuO9IjDYF36HAlONPS5yWcAzCx3GQGCq
siZJF/qaFBZ2/PFdtusOtGQrfU/ANvLP+viZMgPVQBs7Gb8kNVzPlTPUZMaSEXLe
BceZESgxdVTc+6eyib+hF/7FX6F3/U86S4fPq/heJk0xYm5hGO0539CjrWe94sW+
WGt0OS0WfJ0k6WCZv+3mUkFBhtTmdaJFNhKnrJ1BG03HkA8dqbd74QmLCJJ7Eukr
kHqR/kGZDL7JVNsuTecvmqVgTODPwpXmYna438OXFSAU12RQpA3Zgjhpf0vYw5lz
sQr85/PBj+s3g0JnzdxlVfGDIE/UIuET5RWSvD4mVpkvlC8zcQYwAaxzZ2trHy0Z
DnxVOwAS8Gu1uRTUsYMZZ6rtXzahUqLWadW4LUGshQPDaXC9tIQKJhF0pbHR/8xd
jQ81SEG0Mxrwu0qwiIPNBpCDfb8oG8eKsE7jpUrrXJ0kKpd2EEwkjtGUpQ6eLU13
+mkD+P4+SAyNWCGBRklgwAwiPiFjGMrMUpwQf/kh4JdjKw/PE1sUyIC9HfXc2YuE
wCfgYfg6leo4fEJtK+crpL0xrYLP1NF/z9WmN1n3NwhY0vaYUqWl/XYCH6WtPQO6
lTBJ+WnQaSaaQIt/LVR6NoEWybPiPr+9pD1pwpN7eM+1HVZrKx87QupJ3et1j9yY
wevXyH2XvVTucTktLq6tN/nDUj7j30XO7KoABlH9YDi+cazDT8y8GAj0AhMy0TNZ
wnWQDbI9Qxi6x5DIAfpMGEMK7nSAc8SmuxdW+RvQpBSLmJAcIKDtQTjYRrNeGNhC
WesfEa7w36ChUeW08OdpGT1jCP3VRuzkPx3JTqY41pHqrnwKxVfkOspaMqwhFSgt
DvwQhf+hGS4MPsopTqyQrWDf0zOX1aG3vqqWCB8wGTbO0wFnMu0ZeLpx5IOmnq3J
Yo2JkkDCf3eIxnCgfvvcN+7nUhSDyt/sGeXtaNFn7+Da3Q5/Cz3TPvbxTvEV1GdP
gLR9tuvYBsi5bg2WVL5LQLbIPOC+uIjDlR+Dy4DH6/jYbIh9R4FA2qro4fOYhCj1
EU6avAHBxZolkuJ3P9E5BUWnekDHnozUlOEYGJVH22Q2OluMxXUa8OzYib68JgvT
sx7t3hAGfG8ekUQsdGM9mwEoEoR7COfUBDfIOiV+wBZMz8a6jxyWTP0o7lrfbbGc
kZV5wcTX/QGQtC73ZpaofrrW7Jl1ybchhS7DC2xt+8w8FQ+iQ0wEEbAFK439LK3L
xPwP7WmX2WqjjucwEtv7YmpO/eiB5vRCsq4D6PKLKfPX6bpM79jMpZHxVtDhjWdV
Ekg7l7pZRMafegUMcwp9bqblpXJDnfKC1mno9mmuk0JD0FPA1P/kN0DvJETAm2NM
XZoudXkYQ5wU667iErCRSc+3pcH0lrDewa2xJUO5AkgsL5oRdTrDULKCUudYbQxS
gyz01GCkmW00zAaG8jNwqcdxDc9LgJzvv52Ji0EFOpAMguv2kZN4qmeGGYLf+hY/
6FDi+FXBsSnWjQ+5ZJR+tOPD9F40iwOqNdSDWjj+LV432AtPX+J0huqBPtRbcrjP
v44VyklK3MdoSqOlfq120X6dsrGjSphFkeKJFP5xdF7VPVeVgLVu+LiXn433nRgd
vt5FJQ/2nC2bm9/UH/+0cIaZxWPnF42fbeztY+wQxSev9EdiRne9n9qg93gQqDcV
TcUKlpFat4GHAV/T3voN7Sy/ySBT/OJfLu+dFLyNVG4ueldF0GqLofyscHO6lhRv
j3tp79BKOv72vKtbkmJ0welAHD82Y6v1CEzgv/XXy3kV1fPO/U1FMJ4iQwekQd8Y
Z4eLaM8RZFo+5j5RO6vC0xQ6K/LxIy9p7Q9FosV+JuiEtPj4QLLnrHwCh0DAqcV2
fEPrVCJglqFCuzYeXas/kzmiIzR85DIsuNekv9hniJ0P63cjJLda7eCvdXX7z+vA
LSOpka+4mfXSJ9m9VX7ZffOZ4LAgQQH3HRb684C5Tu705zdNMFDbOfQQssuL1MKG
IwgJKUBdULTcsevR5W/Ugs7FrROXpfPKqOOhCfF66Dn93jekgGmJKLjvbz6r9ANv
HI08pq2Tp9PbcAMCQwtbAyKFrMP5EuMLgUegrWKDVKVAs5iR1phhpRet9XUqWkKB
VfgpWqaPgunYvUcMbdT2yxcXyTZ+Un1s+Ef7UqExHCuWYxSgEkJVwJHoZU4aB5b3
7NjjmsmvnFrCdTjKXL11CFRGburlfwRcxImYdsSY2udYdZEOYMsToufdjywkeEns
dC6xiUC26MwSMRw4VPQQW78Gp5hsN7H3mZGUqxVHuJOduDx662HzDIl8NC1Vu5Z/
wrByFLPyC/cwIuT835YDTQDb4uGodK2ILC01ThXyVY4aAKeSayhMNYi5y7T3JYfP
SBpcIAzCiPjuM8fHuWwJupQLiNxKteCC1hFhzDSRbD4qVpYIyPA83lJEVrX0p/Ju
N97F5jgOOXUKGIWuHuvkc3NENXIxa0eeEJUNZ1I5KQs+MH9BHPMwh8/myXo6NI/Y
WtJIM01bEiwBsK1PCBFdXEToqdATDu2lsP15y/qBco6JRJyrafUpFIptTdZzhzJ7
ClbBI7GMtHGEVNtaACrSSg5QIvaYMpJCVHh0umj1fX/hZClbaDUePk7OCj3JNix7
Ox7iaS0F7Uh0uKyYBnpGZbuhsw1V8BCv1jzDh+v3s8bSufi1rjkKF+XY19NrygE+
6/QE9jnVjW/QvfBQgzyIYP7Pqh4KOgv7B4yKLjTSfzRsZeTAyOXcCSq8Z+Zb0iSl
UWmEx4xvdJynJ64IZRHO909o+lV7GxDhGwn1ctGs2bVMT/OzB4h69cRRh+i48rVA
WJ6d3ku2rOQlaZp7dRFzxLPCjw7p5dz74VYjlDIolsBtqZCbsnrU3SMVu9Hs4Xrs
nSfk2bNHS1fpcrxTeY3YcpmYqtz7owoVB2EzpRYC9+58MA11CyAGQGTO2qOMjNvp
Hqgigo2hgpwIuvvYau0yYZAte1sDVY24NY6wJ4um1FwwL8eHCy346VuvulY6IykC
2Ado9lPFsjO86ZZCXhVJYgwnM5GvSfzGQYNksKmgVOjeO7sAlZOzFyb2u4ZF+rWJ
HP108oisHqyy9p553amNsonPqBZGkWW+vqENHn4RwuCVv18H86nBGSUSVfvBYMod
2sOB667UHx/2g1ggzTQyimunUdOkumk+1xW2AsczbeZXYBt3nPtI0g/zqgIIhYue
WuZxxnXmdOqL3Oe4sg4MScUoXlEdGSeytFqGKbJgbUbAAY43ZoZmqKJkpbFnWWOI
I/MntUs9BGFJmsOkKc4JH3elyxn/oCSk78waKSNVTlVHSFTNle8PoJ6WMS/VumCO
GjSZjYsjteO1zKqDMlAUrWm/89RewYQAq32MVqu9wqd1gQ0sgX1VusxbjERkF3nK
+BuDtRSlMhtTh/4XUnWouhhdauclM1RrnQc5cJQiViYLC7wHa7lWX2FniSH7zWiq
fGNpq21PjgeQw22B0IgCgmykBIXUu4Pgy8Wvmqb2wOeGtXChjhH2A/itgEYlD7T3
cKqVqB/AcuzQvGmHBrU856eKpOCVPZCRM0nl1reaPtylFYksZJTMxTOm6ghdDjeg
nYqya8Ukx7sPPj6Q/EOWDaUXSQLs06Z6bath1ESVG8a6il4pivvSGEzBwKXAeLJP
hN4fxphXE2zVEVREP+KpG+SBeReyAhGl9qFl3dSQT3Lc1Ebun4DQt/1HszmvoyKf
dNmpLc9HVj+BMLWxFbPKuTXp4rEkY1NfSyCUPBu6mjvqVYVqwMx83P4aYdYJMf/i
qc7GDqo8XS117AgOxJWazzRbBA9tfNUAitcIsCZ7FQX/U3HZ436cb0L0/UIvaOAw
i1xfkba1TyX9PINskwEHLbEaSegBkdZNdJFBYbXTPFcbLb+7cpzEDO1vRzzte3Ye
2RDSVPpOXkYAaPgQKqCR0nVmqgYpmW64fWfvRRBI7sZTDTg9BFiYNCyZ6dOMcceg
4TbJaz1QUG/kRlUdbrZcaA4f6flQUenmnT1SkKxcBW2bRPirVHEISii2imAL+cRS
dgIwLHBTHG2hKqMQoMB9B3YIoYCJNx149iML09/3WRkYXUQ0WcaGFL7cEKLosAnf
jHCNjeD3xs/3LNdi8Emi6Y0xb71WtWU/77Ed5uGB8wFRX8EwsF/RTQGvaBVrghw2
v+e6falzLANsb3nAOGyf18w4Lg6csBY3hU3tmVltjRyi84YLJ8PGLCAkMCcECuc9
F7uW7CLlOoudpnfaesmO5e/PQBxJ2deamcQRgVAFWSgC5zQee0lDT4rlngZOIwhY
sEj4S32NfP/iQJKyH25p5yXDV9unbdfHajZQCzQHvReDWuX+J4V12TK3Dy8T5jhn
Z/iwzywikOG28N1WYPBSNUDwhOjptpWqisweeDAVfZi/uijoRPGfOA1lhh8p4cRI
u6/p+vZgzdvDEFGjDZxPNYgUwa/SCy6lP4e9QOB7WQImKaIK56eBbfSjTkAFRy41
b1nsO3jayCYJ8PMt0fenNjso9XHgnBn81yCHlgZoOq6J1+T9OL/kWNUIcSaRoNBG
SCGT5lrJsUHZSl+YoNlYq9/hbbt7qkSLBwtxraIhwjotsnnSED/nuBj0JJTdy6+f
3x/7IwsahnD4xHxHkhbIuIA9n65Az/hWy8pEtvyGFwUkRkN9XTfLS26qV1Cd0dR2
Hi8cFFAvOo9XwjZMZuhgDKts0amI13tfKfXSsCdQdV2gpScFQvpUJtbZ/RfyWLet
YpCZMTZzeHPupmXEbFx2GiPq3alH7XYUL0obScFQ3/2S5a+c2CRjsFXzp6KfMu0Y
RPWEzIqOkxeyU6KNeFR8igIb7kxozuhG66CETDyGRtjDeGVnzCDUubzsdczk8pW9
z5KqhS+zsR0TXAQVYOAmcsjN0d7jN6RtgtzgVdrmnqWy5Wf5fgzJYntM4YMMCBDA
NtVnUUAzPe3c9fMAEf7SmKhpAffLqVffdS74Yx2rDjQ+/5f6/EMbHOYuHUIFcMW3
HjSinYmdq5jRm+KT+7kEiNP8rE7ergH4bwRqCUcsEKcDLI8cA3sl4vL4SybVWkke
+6DzpUQWO6PzwlXzlObTnfH4SVaCwaxpbVuLWiznpnApBjXg6PEKJ6eXCmWG6KXj
OaX13LgEB4gOFZZK6W4hYoJWH+/zRGPRILtHfUuyPYj32RqnauE1Dl/cdJ3/t7LZ
6yn93DAt4LBLiSh8Il+eQ+j4k8GBTqf9eu0mHecSpOt7AIqs9lLAe8kJKfhNorny
9RXwIiqqeRh1up91BfH6a3dkiNOaMGwuJys8Dci2AINU7j7yYIDD6hHP7RLF5lgN
OmWtxb56EIOUlmvHlc0ckClxNKcCoKfL9hcmj1Q9sTJ0dzSZOM2LZlaoO/fmiRH9
KTS5QlhHFZZfjW+1FLGxO9rpKMDjxEzD/ot5ZUiFivU8TlRwLwG1kqHHK7PQ1wCs
up+Jlc51pNlgsnN7EI5S9aV53pdCXbz4OOUTIDlEq3YCQID2t2JxpP9ZNFE5RV2q
4trMsu2/3Zp8MOc6TrwK6UDo9bPDGLgwEHJY1NXWO6uNkJwcBGdw20srqxVYZv15
t9MxHmKqZcTRkRe61TNdV4y4Ef0mi+/ZhZ5Y8t1bHhp9LtL8llXA2E9O4W4enqsf
meFMPgivAoLMhpFk3ro/IplUD/y0H2FIYy4LjRi/Ew7IvoimJwtUKaee0pHR19NY
nfauIcb8zAmR2t0Jywo7zZCENqjMB/jP6cAkud0kjQIBZrzcPQx5o+bEgi+YPlhS
/eGazgGxY3YY0dtdUxLwaA3NzSflEDnPUQITsLQ7a0x7xbMBBKXNBz+5NhzkwFDf
BXki89FtE4sO4OURz7aEl1zZOQw0GJNo5dy4n3j5B8A8bt312g1RdUFdwd4rOeJc
+UqwyVeioPe7FiSfOqEIhGVOyUul0VSQrolD4GV/m3UfkfjHMJ7uQhIzz7dK+rwZ
/SWtG1JWHuEqMSJak+Yx9XPe1121os9Kajt3lOv22Yciz58GyQiO4Ns8r9rQAK2Q
LBSVpHzKPY9KADP+V6zufX/HjMcxs4o8OdYkeFolF3fAlYphRSatX2Fn+TvzWzJX
ZjUq0sCDTzo9n6v9L/TX4WTLhQMdlf16MygoOYCFazMx45yTEAatmN7DzJljVPgD
j/RLzs1TRUxWkt8eDdBzm9F8mgSO3zIZ9cKySHAo5oYHu65WDR1h/dg9afWOhy2k
B8xwTjXJxATzFpsz4SVTvxVRiQsNgnlgKV3mi/j4dkCaAfhwgzI+FgVxdR40IFU9
Zm7ou1M52gruTi9cpD8BRC1/m8EbP2nwsH0rfRchQXs8R32C21Q93xZIT4pwuGQw
pGYZHo5nES5Uv2N5ngLjWCkE8DKE8gaEPgUX/TeHs0B6qALKAux2jFN9klQ9UdWV
ZlnDvgrwD8iixcSthNWUsYb3l0DhOabITvXgZODyW1N69t2JjovwUkCWpoxEr2S1
8Mo7R4ujS2jCuVqEcon+gJkFFYXiFYdzobOY7CcwkZAG/6OxMm2ZV/p5SvYXUiT0
h27H64iOkZBa5Rrje3HHLyF7GOQ9YnMpEGnxa0baAXVu9neB6zIzBEuvzJ3X9265
88JzeNg9Bc1JV3Lca6uRdSSzkK9NZg3m8j0NwbsSZjk9E3SXCdDO2FyBzVQQp0fz
4yLbtY4JpAeVUKwxPxEQuhhXDuohTRv9J+m9jsjKr+P/SbSTyDAC9OL2fRD71Toz
i/dpWVxhJ3J3Iclulsrh2yqjtICHXRdZSSj+eo/fuYb/1n0KiGmjmWNS4zNX70o/
7bXoOYmDjRzRuEcnWKm7M8YQOMaCq1ehaO2bKituA5BKZC3RT5Bn8JS2/Qfd7J7T
aIBGBmpFqm/d8Kd0+blAbjCfs7JpMO5OUhjYq7fOWEZpzZZzcYyuyrLAj0z3uH09
qfHMt9G7KOBQKmaKzsJlt497vAVUfHolzJJpX3W/9ZisH4wjESKBU/vyyzI6qW8D
+P3uxVqdEpxqIgwlb9WpG1nLAm/WhyP8ZW6yk4/h44eOA7DsyqL5sq+cYuhLGCgi
vJlt55K9FmY5nJSV0xaF7IQRK/1s3xgx3du7u9PS+BA5y19P4TU5YHDqMKMEUz2M
Vf3x65mepn9mNhfTHF6tCqdI3KLR3SNqS5ozvsKbXb2f/e723gpceO3JvkuqHpZZ
G2Upob9sbGKwYGcqg6jcQ0VFg0OJIo27BGwmIb0wgliHs0dbCFYEOYlz9X1uahZK
FA2wOZiTj95ice93sdWYqsCiRRCwaN7iKNVuD0Ogk0S+CLlKku5YQZyw39Nt/ZXv
4EY3MmK20KBt/vBXEgyk+mA2mlVpDT+f+zeakxf89BGFGTEtIBn3OrJUCIaDZHy5
xaFS1haGjvpm/uyafqMvVsN68hshfmbJVsol+eny6HT5sTnFxXQ2N8F6mswymqL2
HAknW6A9zNmwGNZb1slY4X4FKCE7Anio7DYioyyj1uGbjpRjKOPhKqT6AzWTZJpr
VyVfVXtlMgWynzQG+Bxeoi/jZHg/T6HiJISpZkPDzmdPkSkycLlt/20D4OojfZoB
T5P7j3Ang243kSgtOowJijY7Klp1VrDpvFEuNZYavydF5dpGAE2ZAG9ORe77+/h2
eePoZ6NdMyIhhbTMB+rpIPwPhukCuSwpuuLoxcmEopKvFYs+SVX8QLXs5SgnJIN1
+MgiDKaJ48tHvO0Fovr5Ires5fvIvrdqt1dBQNYqDYipTs+Q5QZS87ABhAaGIGKu
OO7YqImc4O1aEJUgx3226hHrZcZDIGEd+0fMHRB7/U5Wsw2M/V0MDwvYALClTmbo
LBLWPU/HGFUndApBM5XKvwkuY+RuCHesVYR2KRNmnNFzJpqTHolq8luMQ903iePX
+tTl48bKnhvjBTKFEgOJHkdTujhtYJizeWrJ4DGBszo8kwDh9PpLPvp0T1ZIcJtC
YqU27wDKxn2jU1jnesfy73OU3hKDbITCiwK2p4f8+HISjSauUZvwVw6yqhsFrw89
zPGao2Gs3PClyiyDIyKi+60rNgGE/RvkaVWwKoBToWeC78QGR4/bdCMlBt6+DDt+
NZn4tYCpy5S34BTRFyhkE356b1cHRW6nUimxWp0Cd5C88UVt7NO3mDE0Wm0zU7JA
z7JNJI1n2VM8zO0Fu6GzXdv39vYkLTrrlrEhK9rXccT8ehGQjOK4Po097eUTTCk9
wkrfA9JfuR7jgIE8oUxUXF5GvZ+ivMmoAsApX4vS9Bi2U6are7KL5hClDoQtuWlW
/ZenAEdZEY/Z5/eGt12PFNoxCu4V8XzUIh02wsMRJka6oLacPUVLRJp96gZFXYCV
qCM/jH5l9qTgv6FuPvPB/isXz5T3RputjE8rNwUiXsxpICftt/h5fhp8YwByfkyQ
2zz8Fu8JrqN51Rli5oWV0Em1tZLRiAeNp8KEVhoPPnxIPpA9NhES2dt0pkTK39VE
PLq4uKfUBWqUM7wHgJMbGyplPzUBvEqm3XDGEARQpOPo+oEuY1uNFPN3IdxyaG3T
7IXfatgc+hJUCOika12vSbObpNf9y/pVHi4MTH/84aqpsrqy0uAJrAuZ2AgR91dX
4JC8R8zYtoYluY5uC8veKxJKrbTOUG4KG0tVF184cbpqYKpm1vLq5w4DcVRTgrkt
gGO+gEwwMAzCE8UVAhkfgVo1Suv7+7UcwvGH1iHcGEY65ekk9rP2F+75mInlrqR2
yoJVj0bAC3GsuGrWfQkW0xaBSTevyUeq3D6/C/SRnU+4vXitGwiSs+2o7v0X/B6P
f6A2dg4ZD3j66UW90uz1nfx7hOW+o66eCsZnaKTqNxOjjHgSbR1LoTnuheF11Jin
zuLNnlyrGRw9yplLQv0bC2NDmBJNa1K6wbd5whWLOPSnHGaHMdaIbcwEXQTF7wpA
mO1p5nBal+jizBz4jsboG+0oFjkLbJ/l3yfggTjnAj/kbAsWpaSOMHwjUwECvXSC
b8rt3B0PyQI9t4OMQ+HTxuzqI6fIF6j3KYq1DumSWPMqh8d0xsRs6I9Bd1COWFG2
hvwE/h6aHvL8cXAjh+8hbzQWxBRf52P+3+5/ViGy+FoZieqVbbLf0YCpQzZKp1t7
fwITgamKk3neK2XK5ufdOdK+c5cxR1e08mOAJ0gyG9psY8RTXvdTqcieKSFEEKHH
zJgYwx+ONSAXuOdYVZnz/zT4iqa50VV0DoEoYGDbA32yl2+7jVjHodzZLnxSMm+m
31Le0TjrUbmtm0EfOdLYNRPq2sLarpYHNP+2IW7+tc9P0jFQkGQOsdol0YRq7Mpm
d2G975DZIAd7kTaPgP8+TYTpVIdiT10IZxfBT1L0V0OPDPpEfVruHVbSmZjGBv+e
jWwvYsKu6RSE6wzJtwdmZx6qhRVaesfb4SlHdcKzRT227e5/pDUp3BrvJQThDc4B
HRAICuBJUqRpiDhEh+IqQ2cgAtbNsNLhMTqNRhFlbt6sDuC+bV4j3MELfmyb9sh6
T65eST/hSWIHCeAaU8pfE6PkVc/VVaTeZ9bRwHR8R6pEbv42j+yDAIO6efDVaAS2
pnv8b2J/F0hLBni7XwhmS2oP9MeWCPMM6P5XxNJWZY26pv9K5mUvDu+hFGzHAcoH
Tilp5RTw2g3ksCo0/Szx9SlU5JwRGLb2f8fkBx5/kRcXN+q3hkigUBu9dkFRD7/J
8b3xnYuY8jgpqEbFrXcMbeaTFFi2sx7OGaidcm8ojySoWPIW4n6cqKfZ4rtrCe4c
82AQ4jafHkQk/DXivnoo9JPWyiBpEpPKpRi2CY3P15jsI/0R8kExxr9WHAc8Z9DI
nhPwn9+49UCbjKdT9n2kM9tZhE5bFAi/I5iznHKw3KSoa9VVClu5hNRWorzQJmtv
xxsf66zI/vCefuTnOb8aMLs1031S9Bnip1SszflvpLyivKAK257qlkByEa9HFSX+
0J+feygTv1bv81rEtBxe5gUUuobr+F3GkeC6UTwZK9D3HLOhTG5IolXZJipuKTcT
XDV784rdqM9igz4qePdCj1XorohvgVHbJ2j2vcj4cxlMvf/ARk8ETJPqw3UQbDkk
d3y+OZen6HvFCe5tq7HJybmnGQG3yrR9Dv3xI7+SDNV3LkHpSsTQmRytspKvGhzZ
QXkbBj85duPGISmAVlKzlO8M7OgbVB8KFYbmb0v3dnpKOyG/oO8FxJDSV+r842yq
Wmc9iNtC21r/yJaajpznRsPu6SIZ4UYZIY3uTmS33fsPiOO7MXDSYrco9OAjvd1R
hhx4FJ3XJh+/dVM8TfpDe4gL+Er0BLZgDrRj4X/yqdnBw9Oe5O6BklNUKJ6qNlyF
whvN1FeqjGGMn7Vud+Kummwv9s0sH0xWXzNCv2wpd+xDaimvHEIkwArxvvaRkccN
gv8cxxXyznwSLMFBbh1rCtL9iHsIry/2zIG4UYy3ye/lWWxZwnFXk/e/J1h2B344
x0rQGcKQEu5cvTwPuJyB7+IJZNjbjr9JhfFr0FkdkOWsK8B5ExaeIzqpcYgps6Y4
h96c0FHD0YC68Ebgz0USB0e9hD4QkJRcg6FXO3G7uQmCpW/cwUk3u6nqiGGJEwHK
UBGc9Fz7ERX17KrHws6qJA83aiovyietw2HDILS9UPVOU/FvZcGZvP8+EYtyAux4
K7VM8kjTN/KvIEVxT1KIJ3qojIePYTQxPI6kUDUW8cYaiI8MxUvgPzWLmFbn3aIc
o0XA8LIQdV+GaLyOPYjrHCkXRMMGmoM1P7Mqe+3B+uo3elBgBWQ2PYknIrhSdBTJ
XqlyiYwS12w2v2UoUX1AmC6woqKYpFprQCuLGgp82ldd3x4HlYwxucbf91ug+SOX
hrk8dPvE0818RlLbZootao6EJ5TvIr3as0u8k7lAE6sbLucT2VhT5sKO9iDdiSVt
UiBNgIW3nKJZH7Q+D458YOvZH0AoGC2myvZVOI3af+2rjZRuD0xLUOonaw9U9uTK
Akvu0cfmgsmK8Z7Li+NZT/c2IDs1zOtBKVYkxVdykkcy+ZmDwjl+7yHDKSCXjFUN
7uEcDslzaqkpgcffnzgHgDImaBQ4IFPCdNZ4IpizTOVS707bZdfvpbF+Ey2+YZfM
C2jeHH8LRy9vb5m1YSee1sSokld+8OuKwbKY1bl2gY4dASZCVJGkGx9VPOOpALdO
OCjZN4Opw/FMz7hNTfSP4tUqMagiddOkhA8PvyEx+MjRpdxhAc2Tl5VzW/5ae94E
JPbZM2vcGE2bq/MWTgzyopsqe6N5t6m3OG0EbfhTp/5GcdS17/x+M7vgbEW0/cpk
/DvYjGEhwXALogfWqWV51CvQekjpFrpR2D6sMXyfSY13CRyOTg4s4ouNeXbECyDT
W26AUjuqFXfrAkJyLD/+p2ca2ejEZl61gaqM813tjHbjG9UxFs+NoLEQMvKmoFS7
SZtFVpcWh7pY7SkfvfR3+lJLoBl4STez+mHns4FFYN9i0xHYuh/5wOqQLyX3MWQM
VxMj8u0ORRiUKEPibGM15vLg9r/qm6OlUMZI3Vxo9q6Y7r/bSAAhJqI9FEjIrNGY
Dw35kEpJ6ztuOARx34rLX+6sZlX+xEx4HeUIGTKn5LMOQGReEMLIc+HXaW/FPWCn
3Ro7geZb8yLRqhWHUa+8V1Z+T9+wse5X9fELduTWr7wyfd1MKUOVHKEbN+Z890xS
FzVYRfOo0Nmn3TkrWvTLUogFcIstwPD+ly/YPb4CPn7eiluuVXr3yQ+0D1igvL5i
nhEeFEwEFSDQXW6/YsMFGiLpKiZYsnWoYj6bTVFD10BEg/cZzPCvXSOEIAg8ubY7
pBkd0s2FxSS9g+mahHWdqXzZkMcbY9DqX/Hgf43+M+vKEuvhlE42+nJGVOObreBz
AWMaZ3pZqQazGlKchh6RSITHP1wQQassfwdO1QXmpTMYHmSqxsWjmmx/jZJUZlpx
/qfX699nXNY9Qwi0Ppo8zmoksNiTUub0j4052UYN4TCEJP7PxPO75RsufS9at3kF
IUMnDOwliN4Fe8b8Y8Qtl646uASy3G8lWBaAe7pDg+MXtCOEuLL72DGCixTIA/Ma
ZM+GE/cRxiLJwoaOlrwYv1gpqqQjrd3T2vgrkGVBUYpEvU8xPsqpIb8/I51LNUbw
v8Jh1BXf1ppLLwyfjQvgPcM4EUzbD2bIJ6W8aMX/wKuP5jfBWzspHMB6LULSOmJl
ORtUumrll3fZHO+4MW41Z2xYNiFO26TWMP2rVkyl9vKR/Ve7mao4OKLS3rAVMov8
VYdeKmnAsoUwcqDaPG+danQu+Vr0+fHR+ZxywrXDQEw/geF+iEOnC+VkoYBgCP0R
PSdq2/mgSiOfocX6Wu1NKw9QXoieTfut1Tmp3h5tQEpnW4B/Qk8Prq6MSOYLTSuq
cITi/FO6Ui6Yia1R9x2k0JASnLNKi9xiAvHCQcDixoFi4Fehi31qqdCWGLvhtR0J
/cLFy/MVzb2FrrJqISx/NC3IXwUX6wm9GFXKqr7Sgrd8lC3enyNjCmqcR4lfFGDC
BcSZ97vkmZOi1B8lwDPFV+IJ8dLkX/gN5MpdM65OanloMsS0zb2rb3mo/hEtzbZ+
DaPysG6RVhcsPnCQ425vQbvPaPAr7wCZDjDtPgGpaJq2LDuAktFk2/x1mcNKsdet
5j7NSq/01MvsQt7xOPR++NXRQilCesujT/sqlkIgE8io9TE2azBj2RwiUaytgFWZ
F8YzcfL5tiZjBiCKeJ2qDxfDp8eTe5biJ+TW/DySfAhwyjOOC54K/IhJO+/dCZG4
LifWRYkoW2YP81aV5wtaJLhPH51Tqw+XZ0iWk7oXncOvRTzj3WKtj2bEs9QZzbCT
/16NE6rwIDPvIM7gqV27umftuKvEQNfTN0d2XpfDsz/e9QpjOcmag1LnjmEj+UH0
+EO1f3YfGoVDQklJmJErXluRhebA6EAup1TJAEUBCVIeNyrQQ6l4XD72nEK2IMTw
mJZqK12WtHMnjFgggCmUKxVE3+gLe8nd0KEzVgOs8XVvPdEqBo8tPH9aLmc2OAZK
yJ39RUVu6ptgXvr1x3ZvvgruPOTwFe/Fs2mhks5++K/HwRKsx68BT1HDGcg8OmdF
8JK2B5XCreRNulexMdSru/ceyVCCAa75wxvHx5prECZ434xB1bUqIkLkM/4tzxQ9
6jnlLEFUvM2ppI3sykaW2W9iq26+r4lFRxErs66+smr7bnYKiFsxP3+IdgVfWxcu
YfJfEU0vUTRPqiehw6jpBfFX5c44MvriYKi7+8MVdMETUofhEGbxt9AO6FS+48FM
tb7gMeXWzZBBPY4AWFPJk0BL1iZ9J2N6IP2ZZeoQx2/gGdtY6fkJzR5YfffLXqS2
fx88ZHmnn7oUSZE5TQtLMv8Z5SeOjHX1gf2Uq0af+FBXVxxqLbLlU6yWDwPrA1GQ
9CAhWrNGOXAxp7iiYO4cF9nqL+fC5FWKZCWFOshAaFks8Amku3jzqKiU3uVsBkUd
QfCZi46oQqdYRc3/Cin7Vs4yXUbQDnUvm5mnPGQkbWKssrdHIwSDDmf9UsBQm7Br
AU1yxRFKOsuQvvGyjaQlY3Vaexzj8zwN0VlyY8ht6UKM39njugL7EkutNkoqv1hn
CpH7bKd48F/RpzLB/EF8/VJkNiegkeXLyxZiE8Gvo4QFSTQeUN6Qwm/xYlwnrRcw
NVajqc+Vl8cDwrFBe8pcL/n7KVAtsiMEcY2VY5LxFFNjw347Z4vDhCi+KegkYguV
NGqooVZAx/iN7bmTOkzXvMRIjvRe3X5l5ujBjTByN/5MmVqXxDSo8e09FT4Ndhij
mPh5eQzEVev/cupvxxJQF7vVVzRrhrJq6Lt55aneubnS4cXrH4iNkTIQ3xUMN/16
gib+8GVg3O6JzWOaTW6UEAgoHmrxVFv8R2pAyJUcqmJzSBVXDztnv4k0O1+ulbR2
r+HdD03yY6u20SMhAuiayuAycd6RIIABmsvCjMJNN1yyz8V0bfeIwXvHFSUiizHb
wnWHrg+LvxAeSrRyWZLyCqqJGGzQZpmr4CSe5wEbbM/4uEZ5cq+p1eP+bZTe8bKG
no+kQyeEmtQhK/IKUsiGah4xQueJMINY/g8uMDdOtJR2BgvGrrVWIc9DYhJrG3Tj
icdNq4hXgebQxe+KKo0enuCqdjQ38yAemDAo4r6RP0byBeyHvw2avHfu/rZk7Su0
N/Rd7E0kQYSmUx7iXYPDIQ/Mi8lwTBQjSG5eWUyGyHHiSHYKSuHBlwTwgslIIDVl
asRym3zdnWTVqBJ1slssfcFGr+Xslpe+yGqjhCLc2ZoVUiRLH33pwz0r/CtS4lio
CLCzBWHbSCxrP7M6gasJQPCl9uS/mjoVcDFneXAkQs23t8SyzuPKKQ5iNO67D5eU
t9lhrHbR+MyvIHJ9om98YPlTj0MmRePF4QLWZuFLpgj1VMjSCT3x6sfQhDt/vA5J
0QNRjHt9XXR94IHwv8NsyrYUGRybl+Wl+h5XqPa19qwHOm5Zyda4vlRcoNnXAIhW
D2VemKHTs6ZNerXn6S85NG7DaePFVtYCAS/AkQ7fDJtGU9AhqaY3rqizIFdDC51y
z0mH+eE3KRuW+fomLxcgxIVujYnIkxnWJqplBS+E3YD2q8ru9Y1Guftjr7VFKZJQ
a6lLAbZIfieb3JlpgliAmknUtqP9KQHc+du6Tom7lGMjwqkHmz4LLePr8xIO7a8V
D7+NHWZkdXQ36wM1jKnacOIPHOTjr9Yh+vLCxlpX7XtPwNrGExqwzhKqZhw+9vHQ
Q7cIFN5rcRpk+6Vz+Tho/9780HMjUXBpfBptO2AQ6hczVoH96z4CZQR1TfSDr0zr
SyjFWP+GEkgZSK5N8+wUfanKzOtIYD05B84w7izrSXjuXi4iZrihPvohBRvP+UeC
8rRXmCVt6tyPK1PJa0BJr+3OtD7ZEZ/cb3s5zazni/70GTtF2xd/wiMLtIqyEbB2
tgrnFQ6SabxZ3yjPGxJgjEUp6RAUXNjpthlgfzZ7H7Hzun2wDz+zahjYO0oKT523
Gn3U8NvOQAYJiflkoNgmuZ0WKir88reByR9mYgeySV/ONR0YneuG5jxyY66gm7Hk
08WtChfuFjfz4QnDq1Jp+diQ4qqce/6QQGVCFV0vhR7MmIecY4Y6JD3oFqSIKAlW
4cq2w4/wAAnS3nSKwjOFpEiXE4gZ3KTdo/mZwdId0ABLt0bWwOGn8ydg8MgsVCig
oKflueRJ4f230AV/qW5wuXDMRiGAEfpjEUt5q3mvJQDltZZjJhG5S7KqBYSKdKG3
w6oTl91UqU5WsIAXUrs0t8KeDF0cq3w3BYdRj0Eq+NZhFJ1xfMI791QbC1YlhZZu
6xBSqyR/kJCJo5VROv0Dr4Hnd3Rv4X7cruryfT3ls/CUezzjrq15bFs+3oMORrtn
BB7YpHyYuik7eTI/bwr1HGGawaMFJlVcPNh9CVPf2Q2TAth8hT8qh9rmpxWC49p0
BhsP4ubokblDVrdj8XDHkPWnVKjnFmdmy4U/rQzsZjLH+ejeHDFZ08F7DffWXiVV
CUYnmnK805Yi7exZLNZH/jcyLORRNo75+c4l7/TwkXPJzxuOKReHEZgKgLQqseeX
VKdmt5F1ZIjoGkDBnbQuaw9wX29ZCR46JzFzXYfCR7yAmF8+sufF5R8bW3Wyr3Jz
eAbiPJsBmC5Pko/BLirhX1OMNcAxR5Mn5ldL2iXVXxyNsONXyecZYoy6QmbIqTfO
YjlJnlbZgncfJ+IaRySeVHucjXLhgpbOnll9S/en2yIOZ35J4HVP8ebfYTlqLvv6
IOFrSwWyQgWZEhi37qcvuZP1wDGAoz1sMoCUwdkzpE2sRSKEWtnytJ4RRc9ICIi+
KN56DcPqkPqXetpZs2nCbhuRFZcU5XUGFeJxI84d1vB5OYO0atAK++yaZ7o/pZKh
8suqQGfxT6hlHR+3I8opHhAzrv+kwwt9hu3hHtpd09ntt1eiSGPpC49+Xe/wBnWR
nsACorV0/Rcj5cT4/W8LZx78xzRXpGcACo48y1ql54MaNd3nVZlTqlVEcyjLtgwB
jO11zC9pYZMNVB062Ue0+esZ1TE+LFUqDPYC9/fYEY98wAOIwbKNTXrb8/rU2w2+
F/B5TRIDlAnNr9tJKBGnrJY36qvvN9/KD9twAjRvfZ+Fl8hg+1E7aN5e19zuoGAS
Jte8JGaAvqOIaSUzItEFDk0M4QDbNGQn3qGLcxZt8VtMJXroKWycO5RHHTAWUcxP
31T+1SkyjLwH6TPYzmoCU+ejForNonEl6LGpyTxnwBPSy5Z32HweluAM8yd3BNJ6
IZXA0HGDqaxPEhENZDshYBzw1Eo+psQUqqZU/0EmyORz82txFyBmQiH7VemVSo0u
jZ1IbF6q99WBn3CT6Au8m4ZTgFryMF0OTrxTvNXA7Zi6Ph6wXxRd+4UF9aXP/xUL
4pPO39we1XIPbpjt+JKzhc1b1CqWre9O/WFO6YbIsX8Iu3z804HpDUz3fvY0rBI9
EqqE4DZrPCIZpqV64P13N0OHfewokdQB5Vr0PUpreElhbz+hzHETxAVlERiiSCYC
1PO9GP1JUItwOkKRwUaisH81n38rHphGMBsl6ijrQu4re2VGhpXOgnHKMwaXSbO/
cisFjHEljiELxRdbfM/i6YkIzXAUpEOihv1dBznhLXH2dhnswaMdjVqIHu2frhYI
V+d/cO2HpRe+/wLNT5FArfxTk3Cxmf4Lkl73IId1xk31me2fuhWwWOIfcO/9Z1NQ
/bMW1Zoae96FgqKrZkeHxjIcplfz+lPC8Ak8FhiNJDea2S1mO2uAaG5LmQufoHox
fDQKFaS18MTlKiCyzsebR+xbKmqEdyAbcRXM0Gwibfo9K9tDdJVyH1zV5oB14EOH
ZcIUrlSZJGFTS/faFibDzC1FjG22CLjHAPrY8fWVRoe1tsnSv0SedNQ5518epP5r
Vl7D0ki439NJz/17aPeLQ8zoDGb0RwKQMFHK5o+/CYU32BMcgv5hCBWKjXhjS5/s
tEUNVRDgy3ZDP6c97bjCeir2SKUbD0fjmK6PaD4yjMJI11c9zdLz3Rhed1j7poOE
nZ/A1P0bEsUoVZik2iVFGlsrNQKwKcougze3MdrWgay9+6WwpokBgT7+URQRnUyD
681uJt03fU2u4l2fkGlX7cdIgxLXla35tsaFOsBjrLHyZzP5cn6U2rXgDqcMcf1V
4GRSEZQfpqw8puLLbTSwkVIXAPRRWk33ZWVEPoP2/l/JBOSaylE6rLY/yOJlltEG
BsbNHHWKd39jgMP3Ew9lJSeF3AdeKMJ92VAtB6qdT/YFqAImFKDKNWmMSOUDEC1X
Iwt7Mp9RGfeo6QoiviC8rDwOd2rbbB4KPkOP6ZoNxmJVo1bmVwpqyA8bDN64apht
MtH6oWq/FnUDsahBR0PsL7IwFTKtCEAKC6LLN+StShWfH5Pfol0VSYYudkicqsu2
WpNmYhVaxKTJHAxYiZRX27RM1Cvg/rJuDDrTch/gMwkL/HXpErwZLoV8PsQfNjQG
MPevtAEOlWoqvgS7jyxgfFcVnv1dGXrl2o7f1zT7XMkAYKgy3E4Kim3+12Qlcqfr
25XptUblOlTJeZB+fK5nfKWBgb0rJK7cut7V8L+KeX72Ar16bXEgn5PjEP5Zd3wI
yxsxxCMpdnsMREE12s1bgO8W1YGiLaPvodJMYvDel8saRikyMC7qA6IRFVs2XRXP
6AtNcWLpLWUU1oA8A/rtvpgYxbLAdGK7QYKe58MJJvllKREBXqmYTXUYNcqbFhd0
ZQVMg7jAzdqOkblnrBYu8PYpwOIpAe3suR9btHAXdVZJUlxt4uDnF0ZcM54UGsye
Aj48xuUyvuy+C52n7REhzRMRr24FFHBXLJ6VFIX7lQitJEuRQS3ucDYaeFD88HJM
KO5GJtLvX20DglET4WLgd7QdKMAMpGInICYDJGjZTQ9jFNes5asS84kIPDN00tSD
ifFpuueEnYUrCzBjiaGh/wZ/SPSWcY5gTLRW2mL6FDFHGRwuZG4CTWS7dDsRDOfU
VTNhrV328Dh71PY0qdLdkV5np+jPSdod5H2qT7ZITulhxhDNLAAC9xhkU71G8PjO
Q5QDlCWw1e3hO0bCVwZLvi6mcr08Fm8VjqCuxIPGwBrff1B8W+gvHpKGTnu0ORWV
3ddHH/pvK3W18GHl25xkD1Rtj/0/E9BJRnYdWDyCJgjwI02IhrEsch0RpRAARDAz
nSOJMJPU9RIpulbCExydguKHI2nMroq7PZiqEpbdfJgHndInUYxipILk+V2Jn0+a
wTiA+S6eOjPSnCKMGxAKb2sJRO0eICl5U5BHbCaAroaGXw5d5cy7wUkTVekrr3V2
Ev9Ii4Qd8E0EZowayE9Lh9yM7Q8YMQlSN9Uf75Ptjhsec4yFo7SpcClCjudrJnyT
YDwcvXybidmc7VymQvuI4Yfr2Ngs7sQjmd+b0CwVQsAneQlmPNXZ1ajSfK2e81HA
vvzA5+s747FqJbrJgVMlkLXe3SlVZcqIaJbPKsJssZxb9gBpMDIeaKP5WVe1cvNB
u7RSaUYvV/GaBSGer4uba4DJpQ+LLnv7V6HPeWOfoy7WjqJRaMiXCenPDjfxeZyg
5Kis+Q0jnPXYvmpm/1ZQqUkFwWGWblSQUNKc80a+DBhQixDxCIJ5jqUXJW3icTNf
SSYbTQju2IVniGXm/9IiSY/pOflQgxjEbcgBv85ljxtfaRsFyn/d4YaO0Aohu+3R
oL1yoE2+jpttV7qLR3j9A+Q5TpzR24FealMDaVwBcSJO59D3/TcbhsYk/oL+CSh/
t59aTCh4xHSx15IWGa9RlEexw9uRzQ2KpfP1wbPY27kGZ8yexo3+hMKR6Epa3Qcz
VnRTzOvgF85Q6KzXdBScO4XkycQaBIgqNE/V7Yjne1cq+s2U2l9r7jwXHkqajIdL
yU4rB0v9E2Lkt0CZ96DM8dAdbkRQxAIhvncKSmrM44A0QaQdxECeYhYjPO4fRIwh
Hoe/Ba8FQRRi7S/kbDy7QB2BD/UHdC8Xme+bG+pxICkzkfjB54oFrc+prRUiEa7V
iTb19Vz6QyXMzfwJ6/bHceFRy2AsV81UW/z+06DeF2cPSqUaIpyHty3LUnXXpAdY
39Q/KIXJgcBmYxksnbd3EIle81oiT3N2mEvAaoHsL86vHVgRXvMAAIccUJ9VJT1f
/BTKLGkI5i2b4ubP0ft0JkBA2DvDmBfZ6qyecxmiOYWcLelKBJ/wi5JUhhfE/2Ie
kpzQLl7OzjUWd4ZmId+WkEkwA1DBEZQZiyHZEGJtPAR//4FX353df/mUXRgnOmfg
Co5C+7wZvhUvhm9+wTEU6+wqV1cUTn9Zt3hnGIW6QOlTsObuxwXd8GtSKsRJog/h
/yG48OYQ463/Zp2Po4LkrbEbLYvojGN6bcBYP4q2VdYStXr6zDA7YguEkPXriuFQ
On0zuPP3o9nCxmrAsR0y0EMAHCMg8hwhqtoJfVE9qjAjjA3mwftHAwTDC3nGL8sa
/P+HDNdhvKyFaa2ak0rZwCnzYTrd0SkV3n/dOKjkEDegr7qEyKxA8vLn2ZrGf1Nl
d3ifJEbxmlV9+G+SX9RdzsWmvbMgCddKvh5QfOljVbhUfQOC9RrtaRKbwdcoF5oE
TcKu2wUGIhxudlZ3pbZoENqn+wWSkJFrq5hnhte4IBys9BgudeZk8vqPiaTpfaPU
pmCKa2w9BGrNAhW1gtBHLA4TvoXgIdR6M5Jie1+2RDvVa68Zz543OdqTFRw2tIba
qq3vxtdHO1PxjNOQvbUOpCYkQSFPe4pwl5G7KvtVZzp1G/VabRf4bLpbdhqIgnrh
aSjGGWio8b55THf7pfeijIewHxoQZrdX9MHDZ2uy/YBnMqUf8mO6epilFZ625REH
MTD5ejG8ETcIHVFCFgT8X/oSp4V0wMsZ6H+y/H4VgNeMRnNSOLNnUTFbHnq3Zl1t
X5bzd92bxP/gx1oMsHWIk517r2mtKnMSPCwLxx2BsCACLzLY6ueOkvi17mvIzmch
+fOeTPGMG5JIcHbTqAFLz+ZC+aCSitDC8EySFXi8ZhOiUfq1uZTQu1Rpffm+Io9T
YfAzV/d9eNtNhMfr3tBoU37EOux6KEbCUkcNbHKbyqJO28p4QGCyMVhRewXs1d62
FT4qPk1dzmyf/+u819RwReoptxSDW5Qi9JlpU15KaCGLTKHgWPpyAhZHpwnUiXwz
1R5Jh2fgAnnKd5CkJHLIe5daWglRr7z7H8HQcMwfwGl5J/PzamXT4y8l8MCNXGNX
Gft8hM/dXE8mS8He0zYitMyNnLyxvZNLol55tYkVOu/HtPh55RWJpuF0UXVnpN3m
8jIgyd9GQyqUa7/VdeKh/miS07qYZL+hmZzl7EVM6G4jbNFw+dXD9A4Og7FAbW1j
DpyUrBawfnKWQzdGrzL1UQc2XUy6yZO3mk8gtXkxANUd+VJEu441KZBkrKWkyVsW
Lgit5EGx+GuFqHKVMMF2BHGu6Y/KJ3FQgi3r7DvXNdVB7eR28K/x0FfB7UdITatj
fFxrFEQNxBCV6n2eU5uXp9222fckbF4W/DRifyBrLYaCPZYlZaudoDvBKH/THvaU
siDc1oA5aCL5xGdDScHr6EKnx8Huwn7TgQ/C0s0idePgB+avcW225+LtJd9X1wMM
dvcmT+F5Z6VRKSgDd75AJ3UYmSOl6kQaX55o2nAc4FnyR15r3nnBP2o53uoJQ/nI
gRmLwcIc8NO9RpO6A7NXXygRJUxYZG5UMIW7jxUMInMSvZedtQQHBuSI9FFTpUT5
13ZOHL6NDFvUHhXpM1m8XSSLxovIjeh9l6PStFXqaAvUNR3U/h/A/a5OXmKtMKs4
kLziSPZjaAEBPIPnkOKMM+u0i8RhvTqEEzFJW+T0hqp01HBV9Xw70iSQIEMqtEq4
q7INMU8vk1F9TUTg4V5TZqGBLESWZUGWy3olEO5KmP7L/SDUkp4F2BSqUQHatcEJ
jOjo84mhiB2RVr2uZqW8Xj5V1FqzZja2FprrIeWwRC2zgE85oRY8osHmZSLqfXDD
VFLsupM/oAVGYFjTUqxODZln7CEL5boB8Xhq7hBvHAj10+DUQZhHxcuXx2kuw1Qp
0cpTcLWElYuumNU+5Vn8VVY9LdJV1nrY+eoqZ7ObT0L98V8eNPjI2AxF3YkwhHWV
0+JQTh2QIxvZ3Vls/vzdGYu2rgiaE9e5o6cABm/YZq6qYlV/VCbyWZWBclsqT8ZZ
7B+PgfrwmH8rfQiqwgCXYcZfFbH+iHiSr7eE7DfiOp1syClbUnz7Hbs8zXRt+vu0
G7wmJxJQxPXp1/BdzqSv+XJ9LEn0P0Euf778Y7jpVEzMwl7IDWLeE8Fj/7MVbwXr
Limb9A9YvaBHbjAWKlz07FuW0sJHW8hYAWlVSaWTVlipV1i/VmW7KH4ewQQ6VsZj
cEue7QTJV8MrG92COCprLQdn1lprc4ozNTksRe5IGijUQQISzA+X6TyyjRikNNKZ
iZCVPTmpRY+mJO8tsSi8pmMkX7IrUJ9zujS6bmAxX3NjNUTQmThaqZVNeaRLy1lY
7Ep0pOqk/dlHS/qGboS4qg01ybzTqvu8NzTEDYifewDDDnGfZtCmiM5YH0QVPgTX
kY4sgFyOFvbdjUvfY9wsRLHNTTOgL2XNTIqtIoNWEh04ZcVeQt0kVoKsltDHYeal
6E+Fw0FMMyM/XW3LfD0heSbJR/Z5jb+qXPTArrdTWlr5qTudB/Qj5xls+3KSMBzJ
jAKzMqOqtEsqccVeKZdgk4pwNtv0xxLOUouiEVQ7w9n+gD+9OtOEv22POE/i3Ikw
mamMMDXdMrXJqQBvL4lvm1CsuoaadQ6EOmSquqtK6k/ISMTMLaWH3TnPKnv1H+2x
CgN8cEIFMSKfg0VQmZJq8M1T82rpf9+kW8D4Kr3J1Wm2dJFkRtfvI/TRz3tHq7yI
nLUpEqjBJB4Hwar914YWxLtVrUD5HPfDS8LaA9havJ8Ztq8WQb620IFXhDu439n/
4glSoQfDd5m0KanBjkAK0Jh4s+HMsiZCuW0AlbKQ+P2jnz+P1SwxeABl/XWfsIih
Ae06wXXd4Ku2X7A51RAVWYlUb5XeBJ9E/6JQWScZx8D+DBpqq7H7aFsFBXZSUX0l
y99I3BkpYHEzLTtjwidc6LVkUtRP6WD+DmkU5KXWpZXhOwXNJUxFbTjwQuMZDdUz
Oecpmbd9vFEay5nNuZcVskvf8tgAF8FhsoHpqX1z6rut9D/sKmkbT4VVN205wGIt
G5giO7RTkbxdis94my2d0SBMoImrXl+qK9e9NDEMz0KAyHNLz0nd4yAb9Kuaqu5e
0KNBDPWcgAm8bjZyzL8msR4kaaPKzE0sHvVVmwKCdFwon3hVWQq0H2z9KuIUHNMO
fT2CiTOj/jGldgjy68LRJ/actE5mRjuLbdQwj5XMwvaReDCVyvSvs7LcA6JejnIL
Edf89kBNW0a8ALFJI5CZJ1IZMagjlI9kcceBmpIcsjQBs3S2aJ0w/zggFrnZ+4oS
wJQOwxnsaXy36Cg4UjlddyMmPtUlNmimj+n99mifcQd1gdrRbi5VRLgkgo8XXPR2
q0PYedSo98/3GSJbxloizv2QamW/rz+2HI0vQ38mSxzIX2EWjJk1mX4YNS9tbAjJ
O2oQ+ILxXlhff51Mk+OEJQuxF01LfftwUHd6MhzRhMgTVh1cQNG/SfFAaBYU4jVW
bwwKj9P1D9WlswOJt83MHqTPhxYAWzaJQAt1sEiuKGr3E97JqSlwHzj3nSQ7BG9T
r8YALyJPrcyu8MgOQjH8UyOEqGayvLSSZYAi2c7n0cCrS6sk/6uoYbkJLNJU45xR
Ay3bfksjslYxSdB7nuzk9dSNP35BSSRRusiR9OXVxBKgrkGY0Tf8TmtVMxs/ecIt
YSnV+mihERK+VsyycJLqOTfeB5al5Towgk4DaEwwzPs/GG8EuVcBKTOE0pvGtbYx
6uuG6m2PhzpvTqe5y4FnqRtDv9kYn0enWlZydZ844kDyYMFJ918RjQVWV5hwqVvw
5YwsrEyryyX1qAmLLy8INrhfIq5C2AaMQkvNoRd1nNCPM4vsRqCzjTP6oo9OlVe5
aQF2sskMMZZYX/kHg51Dt0Hxe2h/BtRxSsz23h7nCHV61cXIkGelT77i9RPduWgR
Q4GBwhIiDgje1HPucaKLGCL+DDkEi/QPH+tdB2R9W4IFOzDeYmODpuiBU7MHdSTI
kGHck258EfkJTFWZRbKkkj+Kh0zOAF52bX8PZ3tblCvGWaEnF2ngLtnN10FTeYiB
m7cnGJtCvj88PqCx8CEyCW8foYHI/a9gy52vQPLSgcRIC/WEjVGqflwqyw61cGo+
wQZp8qzHBRqWQVI+TP0DykgWPmtF2da2dkfimRGcLNcABMWNJ7aRTiqJrd8BBnZm
9iBpEwIoUCh95pZwIm/DygVZsVwmKddB/1WdVkWauQbzgLSxwo9/t/dBTtNObiuy
h7lIbYdcSidD0aBBkRBDgQp4J7JwItx/MQbSDjpKvdTLU10s5OoGGaN5kC4bVP54
CMaIb0CHkeKTLPzMBBPeNRdCgf164IVzIcpxOgoeA6uwFac9KmDAw3pkF4J/7opI
NjZEMEzdjpQ3iKA5T8pzXvuI05gSHDIeHrkzP3Flb6aLRt7rFrfL5G6FLEx31xjD
JD7VmGpLn87Z/XIVzo7i81PlcyMonU8SbF2GAvfFu3terxNVX8zKYSzGkb7yYDF7
a+AgZYrVAsGP8n0U2hmgB9wAhjNDYCHAc8IjK5bLNXzWqpFxND0LwOF+CCpnOlTT
vOwEz9KT2U6ixSjfWSLOSP3GZTAqSs0XG7GlZdxVLZ62bTFZwZ0fb1t1AmzJpAxK
3P6oE/Kw2oKG4GG4GgGjte6TshcttV6yTEK2vmanldSzID1FhX8UxPogWa+nLAXZ
rq5hsVGwZLGhpmmOoOjbyjVZHkmtINtjhTd0KRo9NMWlPuB6ghNSETuvpXDv8AsU
WwZX0OCqVk1c1wPp9Zlpp4Y6hCMS49oR1RiVWclBu5zJMsRFjFZi2OMxiR9NF24U
hIr+Rc5tIexSq7j5zG4tVq2coC6kXZ7sG8oJPVCpRXCqDU8HQ1H3tUntFNh5bryT
rEU+XWwN9U3ZmnXPkhBj2Ig442pOcA8xYs1SBouxNvSIaUhXeW4w1fO1j/ax/ysZ
Cc1I4GVf0EZjlH846zpCeRC7M6Q0dx3dIH9DIRC26chbXEE1OfIQrDdOt5AHyJVu
tLN97Ggj8o+tiUaIFr1nTmByXvPAvZHMtmCX3ui7FYFlZo4TUEwC9VSmEnA1SN5t
O9PkbfLj9rGNvff6mAaTkYdh69hWQYUO80wfiSnb0mVWAHzgluPJZzWso6+/02V9
/k2FShhqzKoka6Qu/tu4wVPilu/G3UI4X+R2MuilgrtVLn48SUg+S5W0KPcL+I8E
jQY/P8e8l7yb9V7K0WP8o49O0C49KDdZJeXnGllAYrFm1476Zc4T+jzK0a7I0iQu
RamuMy6ENY3b36ruQjey0mf7RYg3QWr4AWQu9N+E8NPDb8EYUWq1gJHVdmnjeTwB
GxTraWMqW6rQQKeUOcaZ45uR4KdZPakLnPdAZPCNOD1UNpWfCPy7EFTucCjPJ8yG
S6SIMG4PkFH4fm8wmtjxXYmRB4nZSwdP2kAKZX0zxNqirBL8w59lS+7kOnfT9dte
LayiSterXnU5BsOZrXu6VS82pbCkU0LnABTT4kkLsfSa0p8iRqwQMIxVTOEwfd+L
benaSP9b/Cf6svue3x/8OFRmzj6C0kpSfEcl5RxpZNbaGcCxlKV6SR/x9OYgun/U
8JeQQjJhWuU9uY1rBZ2amLlkw+/9dm1nj3xaA3MaJVMCU3V3Atk93Q/aAqdguUJO
IoMfL2PNGCcp0W04lpwr1vcCHkMumISzybR7Z77hBdhy8DOYMQpoHyUPN6yqncdi
1a7sOOXstyASvwoxojj8vO+CSpvxGMkM8FUKbQC8UfPmkbFObFSRM2dmjlZFkeIm
Xk/ZjVku2/t457+awy+MmUgPqRWk5QOSTwioaNJe/f1SoIwFJ8OkBBqJyTiQPiDA
bLFdbskCpwSfDX68fDe/w3X1fZ5ce9brHP9ClQVGawUkSzutquoq7qP5V9bqXdk5
2ow/XJK0da7JmiPCVk9xaM2LwfWWYWknvnp/aKbRJBK+32EaWck1AAd1KiORPDkb
su1UmAUvD2fJj5tWoYCoxKjqM5ppDEp8aUTFOgFS0HBzrbeqVSXMPOpIea7VV3+7
9wYYAidIiO3QQPALpaSwWEHci3sc+pmeBYvvlE+G1gsZvdNZ4eqqwZQ+FXMLidod
uVWDzuGjPBxp1GszPd8YsuvCxV3b0VNvMUhl03K7s6wDC6Bm2DilwH5mdXcDrwt8
zwMfGoPyLy7jISNWswH0+54fIlvGfRDdulWLg4h5kdUMitnNdcJqTr8qh9gfybBw
y3X1OLY9S6UskRYI4JJRJOunAvs020QRMxO2LvsYvRvKfTnMKfSaNx8NlL+MEcaF
rJGQCEv4+cgQshR+x2AVRl17/rzXIH6/hFxjgrXHXfcDmjxFlqZ/mF2S0CSvhWtu
HL9cxYG5GvMqoGs82wGzNUPzHzjJkQOyOQtqy0mpG9ph6iQXzKPHkIdhvAaJSfx0
kWg0Z03IFt53tn/LJo7+XCBXj2BCKEq1D5GkxYJBD3ReMiWEP645ZJU+OPRabcWN
j2/UgNyPN7USawaR9M+Jtzv4IoCYjtjwsGv09otU1jT748JtfXr7nKuSJPsXK5kd
LGVNQcuuF6Q5DxylgO51oFEDmJO4ba5dK6S5rrge6w0/+0cYq0fZYOc3rTnz1kMo
+E3lVTO7TULu8ZY67Zwfj3T+k3og+9WxyatBg5+UuhIoxUq0G6DllCmJ/wnNgrGh
oB5OaliokGkgTScyZJn8aQ5iYe351pKZF7u5E1h5VydHtwuVWxaWdyu8YujLPwZF
6bTmO9JLDADeHRLTUKE9cvIdpZwhWiCtrwnI4f3dpOt+20c5NRJ7is+1xF2RCw0l
jLYCmxwVMWn41jsJyVAKNgsyTnPnXwcwqzKIolaT9DP5HdW0TTgXwVkVl9PmtWEp
44YyyYKgUHWIdXiVqOwC0JELhQNvAjL6IM8LsDhJ8SJOJ3rC+LQrgzBeTXP1k6Ih
he1AzHelXcIVpfi6rqe31b4KmkpJCSlFIXxWJIWQTQrPXTjZ9Bk3D9xBoEWisR1h
z9BsFzagu0dO80zw+aW22+Bk62HpzxZ9btIH6NXZwOP+rAT9BNfKOROhREG3dEOJ
qtgsKPrDa2qWnkxRvhv2+CdwVkELosBxTNm+U/01Un3M6u7fzfyuBgXwGcqRhYnA
OVjADMjGP9jEtv6zgR1jXErismUxuA6EP5uowTLn7+EKYvN8plykHyd5UAUfwIso
7xvGOXyVnc7vvxjd2hwdSGEybVDlQji8F9JEezRyCNKF0ZuO0Z4AzJfPOKvga04z
lj4T7glyu7+5SW4jPauT7JoRyaE4qibM0xZ7i6eNivJ3uPsA+NMZ57/5yqt9Ogb0
h+vxSwD7Oj33GmTS/Salkqkyep+qUmX+OOrUI6EyfvX6ycdAQQHhKJRJjU9D/baT
yTZtmy+rhQdSBl+Pivex1djMHVq69Yx8l7KhqsKqbGhNNA7ceyovShoTOnxvFCj8
DRSqYcVeqTSLJzNBEp31V9zWSa180W3rLrenABgBPj7IJpE1rNaPNPWrRjIDltqo
IX25dmPvZrrZAOyDIQIhc/D5BdBBpQylQ3Lbi7Lr+AvUq1bo0jRXrBE+SqYbI8xq
LHpnUNGfv7Cbu/5D3riKPfYJMcCZckPUoSSzG+6/2k1J51FN4EIehmzSN+chqxs7
Ovo9tDprFbS20lcx7M6rTyhJVitV6aFnzKdx6LlktebJUmWoQ2hHPudpgypf5b1+
q7pe46vhcXAMH1T0C6qhEa/70bK37cNzU3/PSuJOzZDG2tPQnmF8nqgZ+i1SNZ22
IbxpyS6z1RZxvpB8m+SEH1JQStlZCfanY0JUQq/DVjOjmXxCIZBy+nj27Ru3SPpY
NnZetqtTSZ3FYEMYz/MKs5ki1dBPpipzshoELTil80I2uf+NdAUSk3zgco26C+Hm
jO3mpLhq2Cv47N1ZoNsWc3h4i3wrRQkC1tElBcFjrl3SMgEN2HGqqq76Tf4RRTR8
E/WYmVtA//IDfnEA8axyabvOipPLAq72onpD0qYtYTZYXleiO8dAgDus4kDGIVVz
u7SFoXDrTreZ+2WVJ8Nw7sWgrvOt4M+W7877P0n0eo2qHBipsizqQZUaWTxDB6IR
f108Wuy99L1np8mxjOAB/yeeGmnxkf1FbNnlTMHdKPjQBEQNa95rfJj+3cLzG/VQ
cVWfqnKpCCYOh9V0j65G9xKstbTr8fD1p1tcycpnZMRi45wN8fHio21lamU5XkKm
6hHTjYdBetpOByQFF1VItAuFCg9QbizZUe2tcmt1Lm9GZNgft7jFJOy3XQFwqoxX
ncg+UFdrkJCY/8igBEnhHORmrhatbE+gX4K2WEVsfDUxa9RIKfSZ1o9zqWZbI6Qm
MxlhhkMOphwIfGxdWND4E9pOyCzOx6lPt/fFFlI8iuxpksaR/E282av48g4XEdYk
ksOFspf4nA9lSjsFasKgbBaZCKm7SftXav05882lWMXTgwnIVYQyDDbpDLqp/VJe
UJF8zmn5MMEu8YivpGE3MaImUKkjmJ2wevah3ra1/OxA2tYuUuhBxsfPRNIeQywv
ZIGPCzkiVjkSP2fYF/vZiHGhpSWosTZMVnEirRLiyqOBtGNGSJl5WN9dFkMMh0gj
0KBW1eOmDmXiA6sJVh2HZpwgDj8YeqbR50COOssXR5iH2DonJR76tP7e6jEpdjYN
ROpH/1dVIUd8W3ZF6RqLI7X5ZQYwmgYzJB2K+62zm/tQXunWCmbkrlShlzRaX4hl
ESddWej9j//uNItGdyBVPMticWMqKBMiD5MHQUVRJ047z4QFn/Sk+kw8jvlxmfRW
MBv3HGuLYd2Ai7BywNT8ECqgcH1Gce421AFIWqzQ5OJ2o0TMxHubzCOlhhwLviwZ
86Oj1IzqJyhaXn6gqOsC9/HSHiCAiTK5cQ8eDoZ+cbgpGG6KHXVXpPydWr03FutP
NoWVKrJy4m4/mBlk0jDfkGTkkveLoTooGf9zsC/RU3GxsPK6/8rrmItOTsSJ1fOM
LfxBnx4VpHTvJAnXGu/D5czJcJKxCjLe+EibyBXvKGRXNHv6IenypHiru92342/V
H1fCSlrYyhko3CUnNuX/xexMWH/cdSWuEjT03tUUL/aFJgFpzoCfoJncpzk4+b4f
Xy/UYkb2aqEENzs3LRWAZuJyntNFlHgVHTXKi4GxpgcUWwgGMZCTkFXjCVa1/JIl
sDrVnpWoZ37+8ldlGR+g0YfmM8MdTM9wo9BMDeLniKw6BveTUvfbpi5E72DJV6pi
skQUZNyK6i02O2S34Onu+BoST1R5SToyQm07o3DjHrZzf80Y4GPMDY8ZdsccyBlV
Dwnxm+R+KaDbfj712aGBnQ8/yO2MkITfTmP7wG0j6XFT1sPRm+mLnmnbR+di1X5u
KSob9azRji6WTOI/uPf7whPijZ7okhrASdJ5CNz320E5OgHbSYicf232rgBqek2o
JWXIbS9Z2mnEDrKzJxL6FdjBLOsZS8d1NTelk/KkRl+rrLbOukev3/Im2lnliLSM
u1DC2B1oyqaGPk826vUlVbhesCAHIV4AsaHQBnU9yyiJXiY6hHhhEDmghVxzgwVq
+M09R1uBzVjEOxC6PPTmv+w8Pf+nNRCmstoAqcYW1iuT5jjYPD/QaNYkHYdbWwjb
9ZKcrBk2aWU3hhxFoBoCsmAUNPKK3HJ86nd6bHayFx0ZBJGNWnlknbkuV9OA+UsA
zLKDTKimKKCeBLGcO3cXNky/bw1WfqxhOSx02wIUbFe42XPhCJO9TzbJu0V0AYpH
9tdcARqFS8tIuF/v45zIgbsdnhU9qIYu9zFrI0BBSdWG5a6Bp6kA58iugsoOoR6o
ZMXwAfue0XOCtHvafxWSgk3LLUS5VLd0S3I9Dtv5aXLWVfd2+A2zJCZykPAC4KN8
T8eXYznPTNH/JI/MdXVyhVkK9qhwYMA0gJpsdnA98Lu5ycnoMzULhdGjIEpHtdmS
Lb+U2c1qFqLpITBe2vrKERrEMfhYf+vaZxOY027tjNNfd3lwxbo61Msl04grn/tv
Y9YT0dJm73XyDuHTsKC9Ydu06UtZfmR2UHeTtyqQMNIaqzuGcqx2QxeVUr5FoAPs
6HO19SSq/c92i1oPfn4LDu0uH3N8nJktnKICOkcooQTgno9ylH08tlC7kjpWbSvj
JsJFRfe0jmLtHaveTNyPai6PUJUKTOfRILC0EmCCki0J9pK2T2oUGCJMEo6SJ9uM
aYJQkKZ2JdKIX0l6LQvb/eNNdPh8RYqpDEwk5wB89ueYr7R61/UEUk08dpUe/At8
Gn/baJjfnud+ESQgXTzUBoSSj+IeEzIf2p216JTeNqfEu6Ntl8lS1PI6AZ1BcZHa
dhq20WmdeD4rmiLaHLCnK4mNmk69CfHG0ZAQLLqCnxR7XerHl/H37kILC9tEW821
KRaaF4GRdiAZ6MPkyzKypZcR1cCzImInbrOFm3Pj0zGgOyHMpUHUBWgGYjC4g3aw
WKjUDIC06WbQoWLoMMNDyXA+RobUMHYQuqQuJlnZVq+vyFxvfH+H8GsLK03QojZv
JIDNXvS8BWVoRpD8voJKXOxqg8+7h9oLqFHqhaKfloWtWYxQQblunMpr7MXxqYpq
poveblHsrNu5PNbibPC/AP6Kb3uaxJq+WiDaWseljCJnqBOEr9WMKKGpar5svQOZ
DJErB7Mfgpcc4JAw6TXanSzwQATT+OPenRXX7eUXKeSz1mTcSrr1eDpRpmlb5KwF
7Qh5MI73W9JUxs/6S3lH3+Ii98rR/vIh7cFv1CzgnhwxVlJ42yfWAoh263pNk7eX
uiz65x7r8Fkk+5p2iye+J3v7BOAAKQhIH98fK6CLGXA5Yb9WYkjXrQ7UcC3jZKjA
eXhjFwwKdbMRylD/4meN/3JA3STYqLVg3nb62uy9EovmqqSsI5wH53fwC014yHGW
MaDl5XkLqoRjZSWHChzFkhsI/8A9QIzj/XI58tVQA1cvxfb0Cf/nwbodlRO7Le6r
dL18iQASLBgm/JMKUd7h7TeEgoMHyvK+Hp7FlgkknKWFHAwj5OA5HqYsnPwq9JZb
Wglnk3Jx6ZFXg6ha9LAWWek+H/USc8FS94nIbDEAa6r37F/pUnJZkxFOx6zMa6GQ
1L/MVZv3gnS6Tu53vJ+aml9UR9uty8Ykj4wsxUbgJiM9qET88Td/7TwmzILTg/fs
ApV+48L1KkqAD7pkimF3W8kv14dTwQH1jqbcygDsrAhxLIm2jjJRtPKOFv5F0z6X
be76Jr8iwyOYqUAhjcqzNTq1nGsaMrQZsZwkTMHBVT4JRzQWI4ipmm2/qkzMHKyx
CTnewbwyddUu/tHYWLrxJdKa9MniZ24ngEY2Et0jOXYdBk+gECU9qhPUe7nnIbEJ
NBr6AvPyVoTjQUHZH7MS3tw57kkpdNT5q+wbu4sUha/lsh6HT6v6t85ken9Tu+ci
5FQJ/KXgXvxSRWw9NE7/0Cg8jjZnI1zi+ffqNT4VN56g6CUzfv3LT7IxGXQVG5kf
QZkcwu7682aTqDO6I+y0k/RNMEbUaq5VmGBv7Pep7jxfyqXQJdrRuE1tkQBcl3b0
agbqpny4S1MFMI/CgMHMsY0sDJBfTKeeRDgJuci7HYn2Z1Qz0uc1ZUesUg2914GZ
8gp50Xdw343UK7kGXT+EFwkDVWaeOAvctEzGxg+oDaEo7MEMRCdCSs1YeChbIx7N
K0mnrW0tR+KmN7SPSOFrvZx0N94qjwmV+UxF+HMNwJ03Fnp7chHNyk03ntRZyOl2
xHccmWWPO8yY8ZnQY5XyTkVB10oUNdrilPbMlW1knbUW1cnhdSEeN7Ut7q2gB+ek
3lPDhDxd56U1lWP2CdanLVksJzYw1kPjoTuuXSztz/N806pdJxjNe90E6qLWPS7I
qlBudgo8aYdN/7afoocTm9bzvGUJA7AUubyPilDkxSOQ3lBfSxGyUKUdV9dKOSDd
m4W6m7T+luRAvRT8Pg3RlUokG8/7Gt2K+W+Ipqci6JFxEHWdfrBN+hhuL4/3qbOZ
jz1cpYKv0UaO5yVhaZ2Q50DCkOHxMnqJGu61h1PnoSKXY0122WIhmPEl+mF1tVjc
1HAaU53eMaOwEfxAhTVZFHHmK8ASzCePgnPJeThHg01CWwY3HnzjW8BjxesjQkTB
jsvgFnz4rO3Dp3I9c+PWu+2qLK0xu4jnMjDuIW1KUA8ogJHn7+iuwaXA1jOgvPUp
w3hb0rGf4lMWxSynStSFNNaE+VvhGCE5lHRf5nzm75C6RWE7GMc1OQdFwdTaPyzf
XTK71JySoE9+UnrE08y8wFOJm+Z2kGTjrmgtt7JsO2GGsvPvjqdrTTWeOBTkDvU5
UqDpvdYIhtktsm7Aa+9BSMpYSYfH6nWFmtlgXGO5KBCUMHlJjJvy2/q7WoS/Tdce
ZL3+lEBbSlc0AgFkf/X+/bx+bXgxFOp4b7KDybwUmGJu34z9uvAH6aTQv0IsTQ8a
bGi82zvI4c60Ln4PTZ8e5p/7acr8njhRalAGi+FSXR2ZqxmFsZoY4Jc/TSSXuuuU
rhOrgIfIoYFHIc2DHP5ykOyfnV9czSUozfz4k+uOFXHd42iY0PK4G1IdDJrhXDyl
VF7eyZZSMV9lY5p2qW2Q0zpgnlMJirJsBoUrANAg0VCWDl8GgoSBS7s3QldBM8ii
K3Qc8/5PfoCw4rdYyrxe6+lSx+0PWPtO/Q51WdhAp+H2uyTRZRJI5JQoL2WoCJQY
gwWTCfBiC3E/VMHi2gEZUut2RlKIKYqnzDHSyhCk5CtaXL0FTWbJaPgHHxpIcI0Y
jhL4XPoeFEj1s7O8FEG72hlrGJ1sUM5kv52PYO3LIoFFwyFhCLM9BnwYzvwuId8I
/q3bmgMOV7QkEVeTCnvZZh+4qnBsvQklsSTrBvYUzpCdMVByBS1WSxeCkl50CdiK
5vG/+oyEWxDnGCAQw6J/x9jS89iGdBeX8j81NeR5LgEjXX9p0mDEg/DOF2o3YlNC
ffhI4vpb/1FIGsr5ZOG9H6H5BY0T1E4iHz5MJ4WNI4zpGyANXUfFOW+Vr/c0p8k6
aFFkqhfz+iv+Pm3S1nZJtJcih6/zUbTe6yndy/H5Tat4cX+9uTQAv6QsWxeB2Ovh
kIiguqOEGNcCMKIBVDvXYlOrAep1MMjl4iT2HYQkFPjt/UWgNokPmDeXfyCZxYlm
vJkwE3Zc9ksauZftpTxMkxNIXwbKfXTk2QgdqCBPn0+sXEYuzF9657FG6LtMm80Y
xv0FOZRqSH+z/wv3Hrln2Sy9depwhSTE3g+65eqafWKQioaIFRYLSHvVlV9cyu5P
+1pn60VnU1NIMpp9UVEaK53HnHFL4lxP7lrCf+ZhoX43/Mktdrzegmij6bsux2Ug
clPcSEiH3uQ+M549PL7IBGM/19xJytSu+JFYIZ1l7nsRBkYYZWDfUWlWiufNS98t
HoDSEzqk8pICdR//TcLq2z/6pzQqPCTAIIaiPwSou4Y7SOLkEGElFr5Ndjbrqmmq
svPF6sEKHUrlJZwdQprpc/lvmtkA7EzM/hqg5Yhjz8MEuU3huhY70VWX8YyQX37Y
e4PKG2lux4Jpq6eiSBLlEQDYwXkQ8/h+Hww9nOppH6iydVzEr2XkFB9NDQ+xbqX3
MscRKlCuQVU+7Z4oknLvHQXzqOMtgxqIpkqQytDAbJSChKW397MUJEyZsgfaQWIo
S/RWrQ/6I8Ui0xpYUa+vyTsZXp9x6lWlaBkshP2rWRXu2hi7RC42PnCO3hsBNSLJ
N41oV4fy3FazGpN9cKLupxORQDI29cV9Q4IkGUDkFEXVI4wGfRgqfvTU/Bk5PZ84
GifVI3GsjYyz5c8NgfYoH5Umlx/qHHRlegFKVowap4nOT/xDQ+ELBa4o/tRfbyYs
cXYyoUFT6Uy23yR/nsyNJX1yFK4utZtvAd/2bHeaTNFK2SjNSMBWMH8G6vsxjFuf
XkilNtbQUewyzjKVqF5hQbxieoZi5mFAXGm4HLfUKARj+LZytQeYMXdnq2X6wfhP
6Wbbj1XBJKPXMNuGhZmQhusqn3X4FIUFtSXG55KSZIP/BWBb5PK/la4qpBh31F+S
3iGgBC4Y0+jid/tnsLnIzQ5T/bUBi036OxVDzpbupGsS7FhmNPF5+eHo92l2qjHB
O9jdC7Ogi4w7s7y/GNdtsiVUtAuQ8jtW3o7O1zZTxaJb1OHaPunEftWEih7KsSpI
vSKYnQFh3rWDQOi+CIKi0cn1QA2WMjYf04PpR6hlk6Cxb4WcRTOMcBa09kf7hTHP
lONoVCSxDVIv+Vz63/vavYyTkkw5+MAf7JYp90wdCWaPaN7OV3g3XvICWycuRquE
yTiNymK3QQVxHXcde9TBhy2N65I8ypDhG7ElmuZNujg+o6iZ6nHZ0ugBFVB0YxCA
t9Na/rXxtAKSMIicKBfV/gggPMg+fvLqvEV4x4xYBcXn1yobs5vSCv1AdkE2h/Nx
FE2Z4BHcnBXYhjlhB6DvP4iKAuUb4FilsRXwXJEvOKd1eX58IPMioOTagZzeO3MQ
zvQXPuL0wFKu5ZJJsRKt3Rb+wZxPE6Y1n3B3GnrT0dLa/5JE+n54z4to9gwc9hiE
EUtJdasyAKoNbuPEnRrYJB0DU6C6SlBRKe107m+E9PvubXi9Uuszww2YyvKH95O+
l0Baz4/+HNJ9i8DPSngDlqReAbMGL3CufOQcBnQVqk8YCMBIYSOIMKq5onqbyjpl
O6c3v5LRAKbSFaJt3ju8DBqUiK/p+POE27aja+9Q9AEllxXVNEEkx/r0d7krART6
xc6ew21tFJYafbIs7BNp4hvQsyp0kLj63Z9EiM2NK755HQfMqsmTh0q6dWt8oCa3
M2DnlMXFQxo230JGbnm51Q23Nh1OJUzFe6GKZW/YhJabDNkNuZ7GlDB94RzklSt7
uojfwtLlbF3h5mnLP3IIv0WV5t108LyRH/rpLif3kXWPvbohv7ACnznL0PLRnXp1
HLK3yjozjYZ753bEzScCH7yQnO2w6hwgYWzZtNFbUKHu7g8v2+LfLChkaHPhF8Xn
TRLWVHlYpysGjm/tUTf4k34eTkghuj0czuvpuA5bdbKrcHJ22UA+it302EjBfZbC
xCA+W/Y2M8zVSLds0edMTwLoKEQ84R5qDE+enLdOquxiRzJMFP1/H+BR10WtR4gT
32DVKjZAw3DlGqUqTP0juRfyDpKwtu3oIUpRU8MdI4384gq5rSCfMnoGzAEjRP5c
7dukNQV1Lqgc4JBMUIG8UMnhzywm9yvNaxVuIkmMj8kj6Xu88Bu9roy6VY3J6dsV
sSwKlizP2r+9GtV266uG2gIqjeH1EOs713y0iX04C6ya27VTVWXpAuXEzzR5ONWM
0aFtUGLp8IdqDNfdR/biQc0tN0ccMLOWdhoSa0rF1mmH50Tdf7VMEKj8jipqFzis
4DsCmmDywCRD6jijDMGlSI7jbyHfXP17Pg83oNBBoWF8LrvlWYJsUyJDxPI6t6KY
1ysIWSDyCWxkdU4Jhj1XynS7jcLWgs54k9OW1qUKHZ7BiX6DkzWW8JVdzZHQPJq1
c9yqL0DKr1O8JzIORbQjbMraYJtNVET3Vxm0e/7x6WnPy08UqVmHuwMqeoev+t9i
GEH4cvIGXNb17Sv8KlmNP8d+iiq0laKag7N0Wl3MAY+CRoolIWV8jaLdApUuxBLP
BSrd2N/zrTGp5eyGfzB75Ihsb4JBPcpdeV394ljL5xwrVhSnCgosUpG12auiINtu
yni6kuQM+Nx04mIXYmi+3+QLKHwA4ELVK0+mc6kgeGoNPrBJ4C+4cXPWuNGlUOl7
rU7h0BnhcwZe+MBJl/ZT3iLWzA4/Jt7c3H1rCc6AMfnQYCnvUhdERPCKoy3uJnhE
pBzFFMMv5qR97txJ9UPaw64v2iSwId2SmuXCNFgBzvDOyYATqNebvge5G0pwPrMC
U3RKsBobhk89fWIvEfKazeNpYpDaER8dGDcXx/Hh5rihOh3O9eb0lEdc0fMaqjfa
gxPp1iVgPlmilNksYGCj0qwqupEihXaoDvfT96E59t0JTNp64FT3jWLD0JA0fy2H
RuAoG81YQOGjVtayCl2jEJhQRUMacjiDRTxsW4hUAzyTaRrml0czZIhFRWwAo4Us
33i82bjNiVnNA3vcCxW4JM4IrpqqRhkiTkCXaqA4uzIh5POh3//i9vEZK2K2dyuh
vspOZflnKWwDCX+N4wYgYmx+yfW2ZL7Mcmx/yTYnLk/felPNEthvoQF/eiMro0Bi
ZCCvVOQyd5UmKqr4Qaavpep34CfrfhoyeMJi+Fwk5f714RKZKQ2OzH5xrzqt8rcj
yj7GSGVOlGMwVzN3q7PaAcYb9c/6+jxLo1ef1n86P4aQH01pM6e8FDVRY7iVnTBK
uWorpRC1pm1iQaZN7xpBc00NPTr+U9TYqBgF85PQuHtkiNTTv2Cn63K8xeSNdO47
CklqRQSdl9GvCR+o2R+yHDDKzyMqfkidMG+g5MiGiEgzT3lA8zmLNCo2YK4umjGq
r8QTkDloSTITbGeVxEedVZqIrjU+e2bKbMP/tPzERtjTGG59DnU03lZVPA2ruEV3
/EKeNNb15uOSZPLi5vFLRUhr99vxuCiZ9uiaJCw0/JVcpWRcR1GYOvcEAYqKrgL8
Ib+Xt03mkDNopxc5I16/VZ1RRyl6D8eOnSj3muM7oH/V02xS+XcyNa/ZU1EIpk60
wLnW1bEf2lRCyX6bTWLVYNa9LAlvbwOi4hw3zRie4czsw4Rukgb1ZRpDbhK0TiOO
tix+k3w84MRFdwLpu4cYHJOHBFAjzthczyGUzdW5mJcKrY7nknH7Eo3vmMZbQzA+
iQSiCIW5CE/N1xoms6xrMgWnquu93lnngqKrKDiHyP7MfEAHja+equ1ZbNzDIqOr
RDq6IkcDxG0ZYHv4FVb47ZXWrDmUq05qkDnkEAOcvqcJOOIgzf4d0nte40jUsOGW
HtRaZqJ0at8hwXAW9XZ9RpbEXCxg+zJROY+gPx/VEcC2JnR0xNrKaWiP34o3SALM
XKUMCYEsITRZw4K6ZByhFEjYhM/uPF6S3lm4ep0O6kESAYuzD2h2iptqAUOgYc4d
CV7Pue6lZXplquVetQrYEycFz+uxEEQpSL3szqt/yoLC9jt7ManTXlwkFxkn6cNJ
l6vf7IWdizy+Ls5chLOJjhCH/rLqWQ9PWOWlN5XIO0axbDMg0z5HX1epw1RrhyuZ
eJRgbnj+DnAqbQVmATbSpEoqcaA8t5p0RGfmcGy5Y6w4TNm4gDme3tUcMs+OORtn
hPcPI/GUdUeTS3HlqN//gnPIgBUiV7mPf/5Jxl40u3dsUO9l/5+/p3XFBTNjb5EV
t7QvGYrFUXQotXDQeBnk48zi7kwlbncRpWtV06a8WyjrF+oEo5JZM7DgTwrWTxlN
+iYizxFbhyKgFnK+uihruNbNETvMfq9Cy49ql06B9JOWUa3MQQWYbCTGnNTjYJI9
apbQ7tBW2Hu9BKDkBUviavQaIVu+plyXjI5bJI12vCtpyQwOEX+8QhLti/b7De6e
CYjv2LjrESS2EcU9PZlKLBbEI5gHnbMuTR0X4SyJc8X+X6cz3oElpU5ml9dBHZIb
rmUTHDW7H+kmKBYn+TSwYNjEBoghv1FfmONLbOAqN52zI+cdHzNB3zHcOdVcCYc5
Mtc2CJ6amF5LrgDlvoYV9VRTWOer2KXaTzLDl1W8Yl0DzOzRFpmRQgnB2U6t945j
uuYFqS2mtsWK69FLX5wsY9ir9bnrYMQBogQ1qktEyutSc5OiUdPDBQAz+XxQYdCJ
Wzf2ht8o9GzmaKoqEPm0xB7rX3aOmR8xZBFDyKWsu+L5dZiAjxAN6rXul78vpje+
BzKsROMCpG48y6EYWxExGkdDbwHajF0LDwGXX2EqmAR4NsNtS9AqquZvuAzEf37L
6mntwmMPyJMY/LPFi2b5dBLdcZaKUPxLG4Mb3Leaj3/L/cLRK/pAJVXCdaI0E+Sb
vIRnjfjvVZsRunQJO51IM+/eWqCeRm8C3nrQF/7cFKVu37JPJdEGMYWd/n6QmSQL
GBsmO1tCCLIgfYBEZAm2PB5+66YLVo7+keK9acz183Xr+qFikqauyBt+Y12cVb4O
wJNd6jquL5Czo0eGiZ0fyM8ln1tU2Wy4tyxCxsXI2+kI5c6r6ci6XQOM4FWvN1df
264YnJAvLDweLZeRmpAXfOjIDT0X4nCGnT5GEPCBYJJb/GMtQwmoW6DCeWYwpzgD
kocDQIL3lxf9jHbe2Edy/ZRZC+F/6XJTgwNYpagBwXV7OaXsrs3HaK12uikUWYDz
IMYfQCEPyn3W4wn+OtXtktbq9VON6FlzjAho8iCQJaIVaK6TiOyo7DjVV2R6ixJU
h7pI/GW2d3ObRPk6ILYQg20d/Yp7rUUEgCkcCJJ5xF0qyPW2AcEVREPW4k2XbqCx
vyeBHwdXRQWDAgDoJCPH4nANPb61Q4hlvZtIOrd8lyU44hWNJpmAVV5hvcIzcpcW
hlUOsmMTY8ws56zNzV0Jkw53YLEpgARimBTVpA+FgfdqO7KGHJN0gr8WQGdySVvT
f5lTCs3kvHuQFiKQL3BzjSvVedvuvFrwShP9xhbZiV/4OKhhXsqisuE/EW1XixJr
RDxgKuPWKMhOCp1Eb1ormRtxdqZDYUshHW29COzCcTUjU8/JU05Nfz34N6NQRpbU
rDoAk/qxSry/lSgb/qnZLi1WFK64M+lYJ5d0aoqWKhRmEMAYp21mxMR+ULxqKFPP
8ieYX7F+q4FWARaXi5DleRDaWyqYXDnzn0JFjcrIaTaNyMeWhrBXP7dJ+eytd71/
J+4jZbBIk2bFJTxUMUxIslefUNdtlI0dflN+DVwErVFNUmxF1o7opZ7MykuylHVb
X13E2ikspP6XSKqWV8QRec3e3Y0Up1XPBl1lqDNwOPTwDO39B2oNy98N0rkv47SG
5HH2qQvmSFIXuCCVDPw8Deyc6MggSNZ9dhB14aKoYJiI6MPuKVmuwODWRhOC7fCO
cwG3ntMgDLoe6L0q4d6wkHxgV96JkPDgPXvjJtFvZ8rC9ogcrZ25L0Do2Nr2hoEl
kWYS0dbMMnio5Ps2cB7Cag1+hmyjnFRpdIOFAT9idMi8EYmYG/i+dKyV+13y6/Xn
ypciVff5ENvb1Y984NDM9QEeJ02XM+Oq4Hgy9+gw2z0+jUvWwYsOiaeTMofg6Pwf
opmvlTa7oFg/cOjDLKWS1VOa5oqL+asSrAONofF3enZlKJerEmUUa72GhEiZuGCt
48uA5s8HzXa+fTiZWHpAtxgCDcUbkmtlDsT3X//+vVdsxDjSLJjJ1xfIWBEZFpcs
cuomug1syta0bzFDJJszR4Zhi5jcpbm5XPRSHbPdzH5uo1UaMTCWYp96GOvjMdUN
GOlKLEbh0Zy0MPEoR8sHPPpwDX9bndoWIddxqq3jtukU+/ERYLWmknlZcLE6HVtE
ozj6QQqMb/hYZ9IBxxNjU3vnXbAmj7j3CkVTmXUeJUYSOcaX/4PrQ5EtRLdNsxlb
RTZe2OJNTYHTkLbmqtwDpqiz0K1n6f6/ylgVCetQHehg3i6DraOMOH/oER6kgGAP
iY92U4HbKm5mlfBIur/LSB3iNtzETSr7jrUGJVMC3Bq/IXxnfZ0q5ffvDpSJq6x7
lAWmxpIEhORkfdTgaU1zc+0jp4TEBIV4fyZ+d1qig3AeYEjeSyDS/3GtoPedNXmG
wohwbiFZGD1bZwAKFfzKfg9xEDaP9SNvpTS2G4DFWZdbZOzDs8ZCIgsbObmAjEjp
DZVZ4/7+yxHbfHHAV/HWn1XkbMBPsAIaokiZq20xaOgvKNyjBfvQAHtIqW8AUzMD
FddCbiJTQfya1Qqov8FSij62GPm77gQi2gORpp4yPFhymmXs1WB3OS8l8AHIKGkG
llmXOB4Ir3nDg1cninC77ld6YQ3DWBiJVZBzoqPt+bc3iCmm5UYYZayfMKXgEwWO
Gpuu78+9SZqVBbDIwILHO+ic4ZNSH3/3c8nHDIYt9Wk8bqZhaxf8KQGBaKM74dVR
mrM+TUc+qn6H0IHfv/yIsDb+AFTzP0Eu1hKr3h1/zsTvQi19eMWnioKEl6Bw2vJ1
cwnPxEM8VFJMEuG3ateJYWGEYxZLF/rA5O5zwiWzIO1jqJkQII5dnh6RC+dQU/k5
unraF13qFobkpwIdNPy+JozoPAzC4BOfRiPySEUKFFeInB7tChzAMEqELJojVqXE
aZuFEETPuiJ6Du/rgkTkyeOHSnwjt+vsVF+SIej4HTe/yG3BwPiYO88F8/V4CiEP
XHrDcGT+evQ72Cja87xeJNquPkJKMzyPDALWUqzhyhrF4EjUiqiqtpsqLjPIk3IU
aOX5bvM5JSgLFxpDX04tfOjIe06rP8leJz4AmmdvV8rDXr1oMmQ+KY0iHXbIawVu
xzpwW3Dw+NauVm7X3Olqs6rv1Ewa3FjWvZQ5P4cmYli05TjIZ3xopYsw0WKddWBA
510dSKbcGlOO8v9wht6Xu3vmN8ko9QpArA810g4DtS2ZyN7uHdifmVrUzBNymnKx
TuuXgQCqzvOGzJApoFZ4NQ7Krm8BTRJAJaEPWHRhkBElgD4MmB+sr+02k31fJ0sO
aHFnkfG7orCmijjFf28RtikbtDXBGSBWhZEUK65x20umj4A/plhzmm11gt5mepBA
K4FfuqClAttD3X4Ut7Z/PpD8Rdh3msasWHwGwxoSukPw0w0PxgEsUgGTlD1/wnUN
HJ5sPT+Ktw8tvn5K7PsMuAE3cIKwKB9XfG8jop3KPZ6lAeVW4FRzP84EiETiSXRh
Nf5Xc63z+1EC+p43BdaXYxA3v4nYizuR9gTuBNloaqr6UX5a9Dvx99xwnohBFxmo
kejpmDi4UhSFQ4hAhHWIjurDA8Ba5IWfgGDTa45Znbk2/PFajAk5QrnJVdaExtO8
8Yk3tJ23X1zr4l3NTdfEHVR2tQ0lccbF+cIgxooCbS+/f4X1A5GSuozDkhe90KHK
PrrE3QPI9i8JSN5rnMrUbbqY1WbeH0jxoIJ0yg1BEvCvn2vgCl6R86gHsAuMxzZR
Iyeh2OH/4NmAUnlwVfI9fP2Gg+Js96Ar1Rv4/nrzl7Ac8c8Y+YBEcv9xCX3AVicn
etb+5wLplxSeaN7HU5bElMgSdyal7tMEHLi5Rd1mOLYV6TDRnFtZJe7d7BNJFuZx
0E4vUs2MUKePoFjA5TccJ6WJa8C8cOTY3C8h4IKioe2BPgaRcZpAddsWD5tl6G9Z
NF/TL6OPT7wurHMl2rHJD9I1CHL/iTJ0+NkSJ8zAv4XP9o3PX8NONzgvjx3D1qV1
yCujw+ACldOpkarRq8a6xnoqH3T3KoNWHRQu92+RwtZ8+ROejo6AmN19K48KdXOK
T9VdFJk/Z/Gk+uDofZ2dfjBrD/5W4wAvBYjOBWzoiC+CCsHRhMDLPKi9PbPEXj4k
a8QK6ujaNX3GyS0u/Xf3O31erJivLSj/ur9xbCfkL8p/X0OBYOlsIRzrMeoeYInW
Q7xnNi9XHrgAF6o8OjuXq4XW0VxuzMkl3Pbv3x6AXQh2k1bEdpDpOUooP//8su06
ENN0pjMH9SYkML3ChYY4SIqK4RoyGNrV9XhF5l+4Ac5z4WP/K7jmd3T+JjwVCh+B
UcTpzOuR5MRRPx3qRccrlcYkZsmEYfz98B+wt13KLTay8BgxeyXY4KUYY35H4/Bq
X3lYjSORf8zGHkcVlQGbqhe6cDyQKjrGcbffAsCb7+3cTRpBAanAKWGGYch8pwcl
o59I3K4+VjVjVFcy+m0qtxg5nwRlgi+FlJlJgLmeySZDf6GUsj+ncJyzgLpc6a+W
n8E0fgred8I/aL69Ol+zrlc4go0OtbsH+UMsHd052hFKAO2hPQhkLH0KFq/okUWC
Nnd0p8U/8JrzJGFYLKlrFvZOhzl+k8pbN4vI25GLlMjhRIBVNVHMlg0STwnXW+6x
7Fc6c1+rS4TK8NeeI1+w9f+cHnXUzoeGtGybgS83uLdoYVV9QbJWnGhhEsKzh3OF
S0es9T4+smRJaBPTsBmHODuB1j/Sz1hX7YKbCzzC/iMtplXEIAaKS9AFcPml1YeT
WroYiqI40L0f+E3LIco478ZKkNuJYN1SLl3gFjMsY/QbH9OBWn28WrtLYQeIDRQZ
K15Bzt23AZmiCOq9uuIesMk6daSwZaMnLBKkexa+XH/iFwqifBqH17ADxm+HcGI5
Wvq0BjeD8vVZip8x6GWQe1fdnTpRswULCZ8ChrVw8RFpztoJ8ajS2rzSqr+J+l7N
8W2+fLMtbqrdc7yNvC/wSMHl7fNlwWXqlYgYTaRyh/jCR8OqSw58MWaNUAFzon7c
0XknL1u5n0kAH2YE+wcOBv+WsWIXqFesb0b/DfvxGwGaK+CAPZsrkvgrCg/pdASW
/DNPSPd/2AJavctcU+B8oweaGZSgSCIZ5NICzuVmnQtjrnQRBD9TPGFdkM6fyOIX
1jSIqyTmiUPUaiN/9DHFvJXmqso5sp3TENaoWwJaHG2xeW02KQ75/+LBLFURj4mw
sb618sWoCjI+VlV3Cx8WMQGMZvoxjm4yRKRqkBL1lUoiktBaxHeJldDMGsa7gfF/
EzdZf5o7dvFPd0RoiMqHKX7xgee4TxKvxKViqtNrUOLEn3Wm+NVZ4IRWDA4MQ8Yb
EkrjEXg3tJPkY7TnN0BCqq6MTb3fGzeY7TnVphBWNPljTYRMZdbZxjiv6C/JDP0f
szKz+DsoqCvTjrcACQPMZy7kdsZHHgqb78ZQqMzw1nfg7ikAGCaZZ51yHMVdpo/s
RxKXo6LFSNN9nPX5VaFrubBpXpz9u3yzMH2NtwrKD+BN6LHyaemMygaooG2a4pLh
qESONKVwbQbhN5K2S+0BVupFbGQQPnAWrkQjqtuulqjzXbL1z8P77uqDqp5OPpxy
fDxED47RfmRrcxCXkC6wAQVfCso0L+ERSXUyuQRPQ+YE2a323efaPSVenqJJt/rb
653Ty6Yz1rzRMDkpHJrNj3oA72DGwlSk/HE1+UuGQlapIf/AbkQDumlNLlUS4i56
cFxzb7t+zc6NM5u4fiQtou12BT9FWhOQfGI36OVWajjNAJFNOjH9J/8sZPL7nxPT
KMuhpMf89SzLw3cjIF1vUzGd12t862sdXwuIDyEARsN4Z40UfiTtX5BGLS8EDMjO
GYsOgioYavDoUlVhKmFgSYd0sUggi4APA6xzqW8e67oX3E9++3MLFhuP4W91P9pO
aA/3sgzY7lBoSouXY4wV+1TDCij9t1k0zj4PAfLrs4O0KuGylOMHVsDPpjeWER8t
421sQ76UAgGUjzjYilRcLXWYxrWn7rs665p5le+AojPzsz81DCE9RQNpQDKdFnGT
pwlkKMDPI2YHb9rUXNlJt4aOF+r2KM5sHrh5PfhN3MeVdNKz7okkCvZbgb3T1Sli
0WMBnc3AzXA4OrKXmgM2lPuHURpGtvyl5gDDKZXYOuLxCUhol0GuFBztHOr213Qk
JWy6zqG/8hi5TRtwMhY2mW2WgxZNm3Tiu3ZMsJPAk5T9M1ZW3m+5nnsbr2pmxnGh
1JEDCHz7y8543qwrvDvAX3o35XtJTKTGEermkIMjFnRKp8N5qyFMstySuhnRgR5a
yWduzXKKdnOqT8vBnBLtfZqh7tcvoO/AtbuZlmywX5xmdQWfgiDF9KKfxFrXSihL
w/SRHDkvD3Q8W5ov35i/pW+O9BXgWBPR5X1UmMwmOEcj3YMYOkyoupXCAnHw3+RT
Ii2OMHifSuKAGxoTBqtCX7N634weFKdj8I4No2+vGHYyyLnRPGq8bmPRKMsOY6rh
0aeafCsV1CQmxv9O5APsrJ77AGq5xoVA5YtDl9vj0OWs+4WxhcH+WycSEYvwMc0r
1bVRLeAQqfOushKydKHncbNjI8bZ+T2sh0+vgSdoICl2I1Ga2ofIf8cLgjstAmWe
FzoWQpwMWQZdOFSMRFIiK6qRuq861rpVGRbMdepXBtoP9Y4FAF9WOGsnDdB0Yr/+
ISd483FeNuBpiDtI8GUDu5MkBiXVoeJn5T9JiqX0eNCj4zmnJxzOMvq0E/DXEynS
vivFR1d2CcwD6tsksy1OvSqeZV5rPRD5/NzGOu48+t5pz28OTkYj64esKYnMkLTN
kQrbTprFX4sJAMcjXAsfUF0n9PqylCNx+F4X1+KtTqUii3vfC85B28K7HVRnXlHm
Bq5Brmdst4qI1f6OUzq57LB8ZxPSa8q6BIYFJUe43EyMvtmNmG5jJ+0QXrbVfi1k
syzfCALfvAP6GYrPi5IkQLwyD6mfFKOJI4UCYRVwLDf92OuTGGr5Se8Egy/uCtMs
S2TRTZJlDzJpvJUgj684c5V92ub/mKMB4ST9ccifmREsUb2PcNVVd4qTKlbsTeGg
LdguOlxKooffj3J86qoE4oFgQzy1wFk6en+Uw4uqTyUpX6NFT4/zFZ+Jassj11z0
GPteSjUavb13GwoDN0Q9ioEVuqpb1fToZQn5/MrpjgwrtWzZBVqnbGMmV8X5YB5v
G/5BDp6ChcebzrP49K7hXgkAD0ivFOCJKNXFjJB/LbcFHWciDvIA5arqu/3f1al3
cDBdANCKi6avF2TGNnsGWFxBb4lxfUKGb7NTbA2DpBwlbAfPa9J6CqZ97+SMak+U
VOXKfc5fa86WxIYRoI2fjiVDaw/nBScct8mdWY5xQgW7NmqpCn9O4sDICO6PTp82
hmpoa3N26l04hNNsnabGbr1p8OZXB81KIgGh5dTlUhuyTJnrRdookmH4lEwj3BE5
kGNS1+HJVP8OzW37VCV3IcC5WoosGwOrmHHtVpgmU1vjqAO88ngJjdXT7TXho9p9
dszKysTSpbGXaFfFHG25EzA/SBNFA7Uj3hWv5pYpOYzRaZGtlGEjDveJaZSdIKtH
xRaaoaSFZAEuEmqodgPuHiO01YPgPn/a2ZqxFlpc8501WeNgznKvhYmCnHr9aZJr
uAfr3h+hJtXM/E1XQtJSaRiHqhO4E+n+zkwQLT0Nx1MddcLXXoh9/Lwj65HqnqCS
xRwEBGQyV0Bv3OuPP1figrU/ceksBvA7HoNErs0uQ1eOXY1JFCjmgHI0vd4RUydi
mCagLX6MaBYEQVF0x9cNitOxI0mZ4XMiAUiHn7GSB2J1JND2SKIx2Pti8w/nCAzS
rBhZViuUgA+m8+eMyLuNaj2X2MNJ93Xv8mPJ/AQb3iy3H82qQ4WJdZLYvIkHPVrM
EbvODjRrKZynS55r+58wGXjxpq0NA24paYyjKKuvAOO1nlIwaih2cfdAZaHNN42E
d3C5nOdzW1OlMLoqlsppTezczPFWnmAvvmKxARH+jpYOPkwhPCUJh4gggsHnUujm
iyBw8EGyr51TtIVDkLJV67ENTeX3vJ8NE3TfV5yXFurLR5uzrDSXzQgJmOPoP6L0
tTce3xuWx7na52/xpbDoIRyNfcMoa9cDLbT9bpGzaaEN5LWF0mkA5F32dGGm1wR+
/RG54twvbzxst+26r7AL6pCqgACpqR1ZPZN9nDS0wz7EQzJJCDzmQVL7gMW+TdMO
LJ28tM7FYEpaj6uV1HntPOHt/+19wnckger13Lk/J4dd/iY5P3UPmp2hOLZAq89/
xc14C3gJPNTgSFs5EtvIeyRXafEwMKrU8oyyzCioWHffvHhx+Yno207vZxelqqsR
fCjcYvn0aGqZPHq9b+jcr5GH3fFfD6OkHFGj5OfNvfWakFMyTyvD7uOAjGLK75qN
n67cSk2mup/yLSRZgjKYsrlBhWbnJRdWOC0RWqjCdyuv9PFygxBV/HU9Uew8iGZ3
QkMwpeVytw4ZfECRv0EExB3tOXGNQad9qUnf71ayIjCoIavyDVlGx+tj4k8ki7re
kpLYmID+YVU5DrvQ+341cS4kK+aOIzbgmgGK2JM1Oy1DUt50O5lO4aPxIaJrYLX9
Ff9Hl4et9zbEiv6m0Pq66rP2BJj38dicICY5p+N7lqygk/hm14rgX2o+7tLnyasd
VZ7DYEJF7cX9S2pFcEl1RATQS1gp9Mi5sKKv838mxW1gAO+xEKPbPKwm+bSYEk+e
QpWyzre2Sz8VQ0+y3rAl5voqXiO/clnzOpeBEq6MPZBOs/poIzj/fptjrhWJ/oLX
uLrQUf9dLa828PSvJtsnWC9+zMEGdULvvve4K+jsjr0rDpbNfP3C/+cQ+5XwFmZ3
mmXh5GMy4u4gH4Rkp59pnxczx/IkcNn+jlu7cHuZvqOaTzLiNJ9xjqx8aLSO47JD
g5rXFTrTUbXf08dK6NRCJCxHQFUOz6/mQDjVyxvwQ/d3nx5CaOE4ed7bqNRXpm6+
8j7B4uFVOcy45FnuKpltn7k9Mw7j487AR+NDbis4OnAnL5BgErGcWC6+S8aay45c
0rG4IPHPusmtteEb61EefHGpTi/8d+Ivxpbzuw8Apq2b8/fRrlJ5iEcUKBxSFSgl
RsIuOkuKwKsI7TUHqtMRz6GcP7AI0EO1SLoOdCfFR2gQ0XkFAWXPXyjETXcWP4/d
aavianNuVz6hAwSYcI9gF2eyruK2U9rlTt8wWFil9hyVti0aMg4e2QACo+ohQzFj
oLpPLO4K+3z02CFdyPOvDPNzOEVAMPXvKmqhj5TM9J6wBZlQ6s96QczO5FRHX1Bt
lTI8/PAi4uTUOsYH8fFkDMQtI0v1o/piHIFSJmWd7Dn2VhN6OSg1dWuEQfIpObj8
riGnvHdrR/jhyUqxKM+NtdeLt7CmrvhNmzcA6uSDoMPAu3uwL3qemjXmFD9NshJ7
Ta0mL4AXS+hal++XQPqye269rppkhxsDl0az8DqndTLEPZ8YviLg3xl3z2hvE+A1
EpLJTtDce3slSvLeJCXhjN9xEgEMvnbq1zLn/r191ZwimZnjbCV1IhJLdi1ZsGwx
ERvcvJYrZWlTs+2kE4fxSAkaH+SQe5NCuOfHX5t7q3VlO77ocMyuBgKzdPnmp29h
oAdM4c0QA7m//EadQSbyJyyfR3Jbhu0k0aM6kB/tyZGbEE6LFAtKmJOxYO8//pyE
YocoNvYSiIEMmN3VOqjopDZ4ExFidtHNpHU3Dnqhx7hgSX9blimQON9VpFHMmOhQ
8HOCaY8uoDBaLNZpUY3hihE4fqPB+PCdGA2GCokPZfeUAHUscUJfIiTzGQclE5RH
HqgJUo9yS1fIDFl6ji54l0upbNNXe1NUXVXuLJJDdpV8bWsx7hvleTrtSho+gBHd
7NnYEAEAxty/0FWbjR9WH9o6uxY19Ml+q7xuI8uKgE+9b8Keiptx8VAjix+LNlNj
0nTsO/hLPp7D39lZeWcOoc1ey26oePUC3p1LSXCx9OT4QLYACZAJUJ/7Hmftwe8S
/xQbLx3hiZPL2ZBWM13afZHDK2Ovid3yHVStRxqt5PyGqlW6bAC+F4jEB3wvYHNX
nUZbGIRo+gcXYoBdSRDOp7n23xFjwcNYYIVfgi8tI92XMz9ZF6c5mqsoNCkSWKY1
UyY7YmRkluEjzKs/v7cTt2Gn5mTiYSAt63yp3GrDPGO6EzWczphA9VVi0A4ZjbLY
gZcHTUFObYCG0n1vWznQvSEI3cyyKBi8e3N2btFF74lrXr0JMDp5Ox7aMl0CZFi0
LxziAoSmNuOExCGFUVfjyNpCoX5ygJftcMrzrHUywhqg/o00NYtT89MBSwtQXi7N
Cvd1qkxsBI+uQQUeTx6qZqDh5NXx68TFFBBRftotJN0FImFKcqi1+zlU4VvvYpsF
vEoaWmSoxrcIC7HpKSk5hc5fn+gqm4NV8HdPTB6PjNedIsWpsTAciazFLveZkvc9
0qnIgcEPp5nFIvYwcdhcQ0r6aioR6b+XMkC/CAavdyILpMs5cZE4d6guLZ/sF2mL
qAk0+H8z+E68nEoMjdzmvuveEDty/duz3OVl0KOl1JrxFA9DEFW1gEVVI8YSjkvr
s4C60Y11hCvkE2KmxOblzgbj5mHTkgygiBB8kA2PYG8kF9su+9esg6IuJN9BG84y
JQGwy5iDvBUMw+PaqXnRMXSASK9Z1e45IUdB/gtJqAmdW8jllcYAC2V942uRF1vT
jleFgurC6tiddBSW4RqxmKoXLINdxxjMG6RlFUTFVc3HriqLIYgZnTM4/lfZhhC5
Tkl0g/gczSJ3qLP6SjJyoN8ve59GtpcxhS/pfor+VSbzcSMPsVkTVyFPN2r+hjJM
Q3H94lS0YMUZf+o02vjDR9SU3ElIpn708oZnS6gZz+nnonbI2SrJX84FBtr5Wvwd
xMxX7uqhB7a3M+UJQi0XO/7kqSKOA8J7vdWsDSIn1u6nxotcHWYsGEeBHTLNYZrx
tpa+esLkTdv7YVwOm/Mtp9QrnEjCbF2qNMdrt0BmUTFHnI8vJL9tGcGvi1rTzEgu
4FlBgjb7RZdYCNMZ1bMVSFLApnJI5FJqAxcKghF3r7JZ1PrMNP9zp6HXa2IVBREe
cPmEfHjYJA9jVIi93y5Vcu+F/3u14ZTv8FsfMb4BVyx0jW8sqfwUe3L92Qkyza6a
zUesoVqLl9GqXAcwziz/nem+T7593izzCaeR7ojCRwkUHrMyojjo64hAeUZ4/Wp6
o0NPHuJbXrlabAi+Sx7D6ixWvsVnIfu5cSvRFIwpgcEbGYEEPOzTd54L1wrTD81Y
jZuVjzce9azy2ohOP5DRDNvDkXcLLl0VbVHS72r1CTkGWCR7aEY6v1/gIa2XoQw7
FqnbKY85VUPWoHzb4DkXygZ8kMdBMnQM45G+8zuaa8Hh2gOCS+NWzYEbfuSG50Dv
ABNFZErcLWmwNCO0jtQP4odT7PJ+eeDyIMOLZ1cLVtfUuGTFjAv0gQzw3U8rQ0Z9
cFkxoZjRGFVnzpWGRpLnxS7TPfOk9ZWlm+CD7q+3r8lQA7vUvzKhEBUieGZmd+h5
N+mA+SyW5tVvoY+cBraK524C+xyaS0zGVtKSu77RyaAmMZrEqJsDgSycVfEa0Nuk
RaUo4zplBHPUSz5EJ68fKWTYIA01cI00ShibbQ0WKEU/PhrjTar/LafGEvSOqL7K
EdCLmOmlrHx2ejzx7s7uqOKmGHBrjHlN/XLc3iL/we9o7lnnxcazHoB77EFejpQU
kayDl5/I0NP9ZoOqkb9KvRDpvEAnteBo2kdmWmDyVVbiGl9HJTC32fy/Wkg97Dqo
zWDR8rkePXNUXngI91ZH6seeKyq+NA4ydmE+lcRxIuHfa75TXubkfHklMPl9ZZyl
Db2oMgXEZoKr2dUpBPCpb+ODZh/oMe8qomA5a4KKgOp5FsxqyV2FPGN5hUSCEl68
yQ5ISdRbnOlmZwmhd9HGOBlCUXQA6gr5J91nW+DWutQHJjKeO/380ZdhVIy4e0Cv
3ML6vG4Jj4d0EwfPcogzNm94vx7odW3n4hMmzzwz/g5T4GKMWakqyryQO5GqHz58
f71vzfU8C3YiG6rGnvbVRn1IZKcoDefGdrwfFOrq0EZMS0tWmP/zm+QSbI5UPfvt
JOfgvTzxBv/miWKt0W+4JpHJCO9E0AW8514y7hHF2JGOKkN9Wpg5e/97cdzipQE8
lYATiwueI8ngdTt8leXaYC5qIiEpIU4G8b6XFPRxl20n5szeaK3najSletg7ehS6
0xOtL6m00wa9liMvXIhGA0VWpJdh+DXbpXj5wRB8zP+E/TRUoFW2qhLmGPhlToYr
oc9IZ53lX9pf5rv8el+0oLkh2rYblzZ/u2vIHc0Gwbjy1JaYYDLrN+3dfzeoeIFr
gCaDQYKdCrorxbAgaxaKPXiYiqQbaMe9Zf4hbt+6k55F5LehM3WTM7X7gn/zmvUa
I31nkBIdWbhKhZk44iQTiFlQyI4t3m7WTk+fNOmVmHASprzGC8EvklkIvzr4bjOS
htIm3ZCYjXldt4VSC0TUDFhTEN8Wg9dLrFI+15FhSXVhD/bJHq+RHe179Z0KWU7w
OA68fRhw+NkaJSKddGmUs0o7hx7LPcZN5AV6nAAiY9CgR0yk+FX+bwgbwZuswCXj
8aYmFr69a51t/FhcVTS54324o6/zo3hZrjytlpcX5ZC05Rg0pvVfC7+vFL1FVe0u
ADZ0PuyxvA/6qEAG3w3LG2tB0DR9AoAN9deB6V13Lm21eFsfOghNC6vwDRrjJC8/
+90xxNK4Whq3lBVACAhnYCqsxHx0lTLWGWP+7f+QNZXE+0zIP9hfdQ62prUh6KUv
fpijLK4xxukhhvpDC9JLJXe+onjxKHKVciWZxI/8HF5ZtVd4rIV4vBWOVnUU5egD
yp4gGpNv9YSVdBr0UIpyi6QDfJZzLrPF02wCbDVOlDmEYkPZqCLkr5OoO/KEWbnH
mdq3Ge2KpQr62ZSnLJ8/VRgmBO0yTJstKOcdQhDP4JdCJosGUMyGSBM9qX25SIci
wjgGI3bomP/onKZ1yTheUTHucRuVwn+7A/SOS3Cauxkkf9jypzU1xYkYQ1Kr+4wb
AvC1Jh59bn8ObEN77Ii1Qu0bDJRgji3PTifPuO9IcZWXt/Ru5FBCY+U5uuuDLPud
m1GOAbU2jIqqZye2XXxyCyzi2JvjVLr5nhsiflHTU73o1+8oPI0TVNhkwUSBvU4J
v8y9IaSd7B1CV2jfnPevwxmMEEmFXz1KuwvPiJmnSSLoxeEL9+2x6rNaAvvRdT7V
jK8EB4lp24M/a5ilsRtUmwEPuesh+D5NM17cSVOCY4AUzGeQvU5i6yUqQRntDv87
l9PGd523moN7uVyZACnIIjSoEzd9MOrFxM6Zd/aksxebhuaNPGkSwxRRW6Tndf//
7VWHqHZqdvMVBJ126vMQb7IB+eIeBb1+2NIK0r5BMlCbXAlj/qRixUuhgjBQachd
wXfsAg223CvuKOVtcPKLiNQbGeoiZ+B/Xhw1x/N2JLuIu0LTRgd43eTAHK+cQOhF
cJMV7AKUwZn1Z/SRiCUXHfs+rMHW6Y0C5RooQC1zoILjfA0uaKRL1d1st9UmRU4g
8ieVMZwI8fyD0/cUsizKYs4VDKZbrONsiaVRVxPpgChEIjEPduS5m/wtoeIl+2tm
zM0OT1iWuLihTjZlGt4Zxy0eNjzeSn9/0LP24tvxIdSzx6PTGsgb835ccuW4dyqw
s9EOb6BbqLX7cwuPc4+riaUcm/IaVrlQZXJvR1hvERgNLDSG8GEWdGUPfIU5KFXQ
QIWY1z1OGunnmxHQSNuv+aZXEgb3ASJZYINVZPoGtHuezAEmIIxKs+IxZIZHcNmF
K1Jd4cgc2T5rBZkrFCeDwn1U+vFxlE0gS2VPUImSXhMglQWiuT474Um0XM/zdR00
jlLcGFg/RujlehDdP7F+w7jVGWDTMcMmlLudWFakWT3d2UlQ7wkOwDwWWQunNonv
iWa2PL9vFSsWteeF8pbRepa3eWLq7twA9kAtI8SBCPQyDult2BO6270aSV4S5rti
Y0QMtF6Quf1L0aOdVB9jcW+ZvdaiMiaBX//C/tej5HHYMMnVPc6grKWs3wPVhoo1
pFhZ/cNIndXk3dtwk4d2NIPba6uEYF1ujFC7FdINnUuC0JP5B48t5CkVzHf6ybYo
Ky3HIu0sgqEH6Jvj527yHT4o/N0QzKVig1d8mJZG411n/MqCtoSvy210ZqN86qcw
xr2ZTSW3DtFOnFLJ2IKVssLWvVCwUwcOEMS6SyPDxORy7Sda93HqhavAszMxYf4F
f6GayWZLs6neTNI89MRUPMjmVEtDGoiJTbh8FzF8MTh+9H2zTvz3pIi1ObNuX1N+
UqGoxrg4i8lA3ojpgLf2cPiK3J7ZkBNWrp6uOBOmGI1k6woJOyavcHi6AN5yQ8I7
lIuMweRwKOcRZcLUWQyI4DJmB9AM+3VkekVyrp7yWrkbK5k8Gx/sB1DUZ+VHPsu8
/4i8PRA03t9Hy22FFeurf0I6RLl/KqabdINODX8tqFhdIXbIuVvbp7VIxrFJ1fOr
9fDzqJhQhHUIcthr/vbffTnj8oJAvM4y3sYQXb6kQ0H52A8yLfoOKuLtBp02j+iL
vJRvD45XVaha4I8gyr/Bi3igUY4zqUmEMqahIfklOGJezcu6gMBB9wlXpJWMlJem
ZRiwJhJTRDyoMcwdfS5kofM5SYQYDaBOeKWtOQd5XA75F8MKXMhjA7up7dfhbsak
rfivCOIiK7rhurtG+Ie1VLqVFZ375WNfXlq6qKbCp2b56ioPLMH0xsZVmHN21LpT
9DYtV1DO1hsZ4Yy6jiDnmDuBUnVZpZtToDjSRarxarNtBSziPkVabwl/+WIXhzre
0HxKi7gJ+VXguhOcX12zEXqO4itpIPwDBCTMIX2PZQSabynvflgqp5q78WNe1HZC
DmystUrLaOnrj4E2fuOgupR4uBs+yAAfyXelr00a71x9OH/i0az3/5ZKRipjw4K+
aQ+DEz1tQjVbIwROxF5F4Wppu/dh//RXbvZdDFpT/hfJkHWWKdlza8Gzx5sDCOOv
X4IVIIJ5Wn3A24fZycOxR6Y1E9uB9TYRFoVJPdq5/k1BjZtQDDrblgLIyp5hqlXA
ikzYcqvObBUL9ZfeRDtWWn3a4MH/VYJt5tHzA/3D57eXBh1imgKNkvJUYT8UBTZw
OOZ/xaDnyScWKLLXDlpOPpMgET+Fkc9ak8gWo0dlLvZ6ej9HEEjESC7ZuLojWBt/
MRLAyqvuYymVz2pFkvkXKT3ba6xhQGUZI+JuKNk/JCQPIi+nQJPPVwlB4VDxSXhi
LcuOv0WDmG+Lr4cr6sQoteOcxSM9Z3poU4Bj+DEZIfINDKFV1nbCB5p/4iGB3b+3
PIDtzV2feoqqQny5te6cYa2hPHAb1NbfHXRAKMOo0IOwKUkApp/lVx+UhKhFI7zo
2yLZFvdkNYeG3OHnobDDyfYMWDQyKSJnpMWLOWeQLLzaQwei+FZ1oBNiXQNEohXp
0EBAlG4oFOwWbiZ9dD090iiCwwspnfF+xNklfMPkh3hSKEWXZNb5XRfW5gBDXVll
tuJA6rk3tT9PXLHQGjMjqBGw3MBWHuS8ffOWekDE3zp5gkvILW4WStMWBW3cnQho
VW9Io1GecktG2OoAUJ0Y3SId8FHye2oMciDpi0EG7IvhVN0LrhOAQeJMdRv3jM09
EBJnci/82KzgBJYxYCINcDGesLW1IXcO/hf+xGi3hNV6HIjVhPrJF159k+Ash0n5
0YIYZxGoyCgCmbVqVambrpQ2Pw7K7IciueymuMn8Two8TCBlbby6Vc1pAv33BJM6
Kpsc4SkDuzWaf+15Zx6W3QBuOyxO/JEh4mAXvjiJv2BO9Jorn9QbW/vd/I/47oAy
+ZmbWXZd0GhRWCAqZPzDafF+lt2B6NbP4Y7BXChgGUJ4mZG+isPMTNmMaIK0XVJ5
yXTBstY5WZnOoTocoG2EuHSyCNHwUQgMiExzWmh3UgopZkiKWVamrR6QwaGVv0we
s7NbKtw+4Zj7zgr0yd81SGFZNJAqrd7j3GNCjY8breEJjoWZxxRIImgzWRc8D8cA
0eUwlobPtYSXeGhuXikAa8eSQquZEVtmakvhvK/nu8gB656yJ6XNjAYlANka5OmW
A9xc0GL/EPdI9Fvudt/4Liq06yREPCzs47W25p2HZNNkMYonDZXGhXvmZ7k9Khlh
rMx3cgpomWkTZclkuS+f7PE49JUwnNcwOG1jFFi4BUcZlJY22W1f4UF5+7l3c+6C
Y6YMuvbfcLGs+UZZdwdESzJMJhebaYES8Z4BtSn21u2YhnQJce9Oc7QlKJYsApgk
MIBsgJZULEpKBDQLWWCBmrGgBzEvAKOYO4tCKo+bvKf83ofYLVWCxB61dUzifa+n
q5XRI8nUC3erf+dOLZHe5TerihB4EkdlMScQy6rNS3zD52f/fd1Q+9/2iPZQZA4Z
wiLsWLZIWR9UC6PRA3LU7yN8Mgjxx7ov0fH0XM1GgiaQgvGhUnljlWZ7kxocRcw9
SC+Py4QVFObhXfe/HVuqu5CJqEP04x2HgPrs+9fXtsCTHP9Y4BQSYwmHrRsv/igN
We15+3+yzKix7dMy9vGoNSP3drCCxSzlQ/gT/iZBTZce/kp4pA4mPOU5c+JvOQ4J
kQPjiav171ofFpwU6hA7oTYjvh2SsiDJ0o9b3Kls/qYAXqN+RSqDhm19nQ/1Uh5s
0rH3bNXgPXYSw7C3dbCx88jYFx3QBIAP8GumExr3krhxjeG88W7/ZnwwlsE3gGIB
VJGt6hLd5NwuKVSKLUmSo5Nx8+Tf2sUrm+rUGAe2JlxSzovmDPYa6y1xo6OgZH0r
REoFBCCyTfpyFN17oP43aB5EVyE33YsKNUYxKuseQOEp9onaiwh4uHGu9fNY7+zn
t7NdQHJCARmiAYjY585iLRn3vzTH+68ltaxWmvb27m+UmKP1ceMtou0nV4dQYgNh
VWb4FesroFyhqwsHFoTMwBWTLrFs+aJ3GyWdm40S1s0Dn7ZHwr7iwuZUVVVGfdU5
Eaz7eHaEyfsPAShlVxqj/5glx9+NrdxY3H09hZvgsfdeSQ2771ZYKX7r7YPx31s0
7XMh89aM1w2G/8SD+bIaC5s8gIhUpiISZbyvhW0S70cnJnKIlQL81LAdwmuoa/fJ
DWJyar7Pu3zRFkaSBR+Y+UbxJgZ1xDYnoBCyIz7VGtUwRcl8tgh+dX1awGYp+6jC
VC7Ym03/11iaZqJ9fOvEuoCxvuXXbcEIYYsnJpWCQT8EB2Q+Ox+VdGCv8LW2Z2SJ
QcTIZ3gs1+VnXWg4paKsLVUV5NjqxM0YhWsqmJ/Hwxhkl/HBWM+IbnI7PGe4/mnZ
+VzWAsaujSL2qmaRKZ+hG7PlfCI+bpl2rkvAPWtYyQwvcwcoKOdg50/oqP9jqVuw
cc21zBedssdCCj9D5TWLRtXkh3ZtqySYrZnlGJwuVJiLECyiUvcP7FYpbP17/yZ9
gSLPE5X4XmhGYbwi28ovKuBCYYSsoWCZqrzndITGBXf1+ARBMynLxSQrZXLljYNh
Y4Wi0rc0x9cOf/6rmXD6/Bh1cTe8iDxZbESMVjkXJSubVzDyPQdpm1YVPq1ElG3U
nnY5+GBUxEbkc6xxzTRv9VuR1V1IFamhQ3r9Gq/Ld1yhHQCopCBklh6xmnL1Q93j
zm28dJUKbKY4ah0oakXbnKiVlR690QSEuMxLnKUKy9sMvraUG4f4Zkq77snlcbx7
OqPp/aediy0So3d9bLXwKNunWvHBeNKN48IKZ2H3Sz1wN0uxOWCrkXCLGvnn8pDs
JpIouUMFh2fJWrKs4p/YavxSAnjMlKN6lcXkiYd1I40tts+TDsF4fB40oBz7YBTu
plwm+/Y88e/5DE+KXWQXsLsCVyanxPjEF8UgUIy31n9bcfPQB1gt3OoV8xkvV0ub
r0xI+hk/3NY9i6Md4umQPMcXUZS7+N+0rvnd0Dtutg5hPggmLs+ZwObOUd8q3Y4F
Ntapa4iz2C7Ncrj6TD8AaVSTXR2V40VuO8Ty0EEKJ6wd4T1W56zKuPjMFURPnW68
QawEXU4G/JKC0JfTa0SqAFs4VQF4HtOU4gzYP0LoWOsTkK7h5i/7URl1X47T8Dmz
Mb8l3FzlmKn02qwHKYGEsZe0pDS1fhy5S4GcNoqNovCmwj6vMxHbon3599G2UA3r
Z1RcL7B789v2ERoZsJNk2J0eZ4KrtVWcWbzDNCvyPPVggujtwLECrqsPGR1roygk
hvLKCPYW32SJxVxxS4MhYuXRW6TbsduawW3NgG7KmKrsvycYqEcS1165y29U3/V4
qvGuQzb5RHnH8BDuRe6A25KZK6lvhSJsjr/OV3lmJLYGe27E56kq3GziKW56WJtt
xgd8tVSISn3/ElPUwkv2GWJpJQpQNa4O8SQd/UglzOfobKFUst6bGub1N0HRs36A
nRYFw7vYAA5d59AB8yOyXWMZl3rh5tsMNunmt+8T+nLBVJwN7bH9hQFFEZq8jjl9
zLgEqjl/ponR8XXeE8Mcq6Vgan9mi7wvIpYi89ibOu4EsHU2JnCXdY0HKnFXYpX7
fybKQ1nYy970AV3V00Nhv/U/VjDeDUgUD0Mr8WFGDoyf+2B686gJHKeVE3grvlrD
xRqMwEBhTJBF4Bihw8CbmOUW9JHAR3Bay+GJpeff/Rgee6vHpw33o3WXDe/xPO17
qWnndwkJngrkz8lvP658JuANxTw8OPHqB+AjAIRT233APHoTEfAI1OCPq+RGN4t5
NxsjYVc6AlL4/Y9nDM6lR0syVuOqilWbOm1rNkMMVm/SqTfgf41V54r6miLhHBYz
sLKU/YMS22IKajERsuz6vhyBIEaM5AYon2T1/n4Y2zP/ZODqWqxRmUdHuVj5bYKK
C3QWqhElgv4DVfC6Gs9SEjm82gf55aaGeB7OazkWktw+19e416NParAL2HBIoNJ0
HdeXJcqaK8PvO60etEXHKiAGIQg4FOntIw2lRQgaOiA616FPVw9pal1SCOZXALAm
nqh2aJ8HNnIj6Z2LNn1cseGBtwcp6MT7oUo3xoJgi+9rAWZK4PNAj4bSpHtzVC/h
CjSW/PBGZrca44qdAiOF+hAwVfJkHzLREAuJ6A/lNcme0vKcAaJkjtgCD+UOwHcP
2hw6tzZ15kQrC2oVQIq9nv56LU7/ysjk04KXjW+XZa/VQP64fsRtUU+yDNPqy+e8
OR/j60iuWw/drT9Rw+htlLovUElyksAVSJab5DKs3AIaBPc6xWGMyWfl5pJ9Jp3s
4lkwROQy27ct5RYA8u2iZZriNuCPyQUVTHWoHRkUmrPVfG5BufpnIA30/2upGF4X
Sdd6CYuWT4g9kMukIVM8KPxoNcWOxh2JlOW2bE0ZSzfHUwKfAMw11s6hXAd2GprL
N21ZRWKnYidgDGcNjD4oiua3yTd+tSpFESdDN9MHWWzWviNvBfAn54fz1FhZpHAz
Ul+keqPK9pb4/JyhKBCRi512ISBPLSIUGWFdBf2dLVjtyKYwV8ztGC/O0j6PbQhM
YBebfyhdQdWjd8y/Sjwn0HE3+gqRcUyOHOSljzNr5Yt8vAohXK6ZfZ/N2b+N1Mym
NCBsfaRq0pIfCQFimXM7UIg9BlDW6H6Zy4yIFbfNlc1AOn6UvcqG99dChWuxGhuK
ZZ0V0ZatVcqpHvTDDFTKfxXY1GrDz/aXJ+OY9KpiFdjZO6Z23STiobaAVLSGQQwu
EuML5unFU5WyZXfaLbCg40h6HTeLzb6RetzOBMmIRJQVc5NEY8aSzdL+30b5qOwg
Tb4Yhqu3QXt7+9jIrLx8bam00UhCMR3FsQa0cclv/XPCWUKrwM2SO4pXs5PoT1V/
iF29uxuiYlMrd5mQS79DFWIfR2X+h4Ricz49v/tJWX7lvwJXDQgMRTVPEa8gORp1
0dIGjZhH1/p+3VtcS4PVVvcI6n7hsddXsrjAvPs+bHgTZFjAdevBLg43XAdN6fRm
8CuTmZbGSV6tZlHfZa/w1xfck3K2K4LzS7sNnFlfT5ntZReRD5cDDos1bAK5Bfqt
Ao+xMqAIPCDK5TGS7cx1mYWuM1Ah54FhB6I+JEkulg5R6xdpLR+S15aBpIv2we0N
TtHCRNuUbqyEXDjJSBsb2RaIC8XdSKxt7WvPnz7B5/P2XttvoBLzreP8VfA0VRbb
fDFif6pXqiOi6NlnvwiBO60x5sjAosrVuMT/IhqGisxxjBeaUK0U/MxQibZzL4RU
S87j6vtp8b2lfmvkM8x+rCcQAP6AsjZzMsdm8dl23Dz/7kzmxOyA6KOUCLuKmY9a
IeLNn39OJbAhhUBlMYxbqNWcyBfCTIwKHhiY0tY2MqZi0WU2G098E8Suzv7gIVt1
iggs7myuR5cKXslrEGJFH6eN2YaHhEeZN86q+s0noMTJWVEKkAjbS51HA98uhP5r
bycOdrggqFlE3Sj3mjZn3UzVcUyn++ZdHMAQUIie0Vt8XYiNnA8B3DkxEeFzr7Q4
l1Ird8K5xkQYPwz9Vropr3VFuZTAJRjia3R3C1IcJztOM37voEzVn59vrABbZhQk
NZQf1JeFlmwYH/9opw0opAIOvPq+Pox1lF9W1Fl/c25b45tGDQqOhEin2EhW0HRa
YazFvgDB90wHHTJ2RGeqZVTSvpmBfwJWie7qzyp5H1/vTH9FR4jS33m1IxdmhTmH
thtioNJRpyOWAIvkLZQZT3BuDo1pNL5FFo8j8oVnqeG8aW0kqU68f9BFNCISRUmd
4kpzi9yKqQQbYrSxjnclOHPGolKp73ShIBYaPzAatHXfUj8KR7fOBPiKfT9aDr8U
pEXMNNwClG4bXnOFbnv8VkxoX3Ib9pCAMhiTWczDuCY/PzoX3a/klNDDG9jVsJu6
skn7BebsBTUBJgQ87hHmchxMnl88crE2MNDUyvEPPeRagH+Pdl9Isy2djHO8hFCv
ytnMKVld6SDt7PTj8yRTFzD38tky+7XMdMVyP62JwQznCDvdATSeY+duo6z5/zy9
15N2adBx44vraXgJOAtThg4BZ4uNVr/2Ca8S81RCsLVUff86UQtDnIdQUD8uXqaO
kUpbhmR3H3t02S9KtrAdtamTOBSCXfhK2DYuSdG5+zMuUtvRAY0a7vJPKx4gFMq/
zGNkwDmNCRpf2cCaroEdYWqUYdp9zX58SWlWdWUionjQn6Ib2Fsp1PxG8ryqiiRu
Rg7eOVUgb9/0iqrItTlzF+3t4KqjsnVMmD5LkqeAyMyzSaWSDqBvLO3PD4MghW/U
hCMlZzgOqZ2U2kxlochqVWrLyvlqJ7ofAgFWk4ZXAEjhC6W8iYM9OW2BBlekXMql
hOSrN13OlcwFN/nrES8fHMzpZ73ALk13JhEqF1R9xnxMg9oXi08/fSTD939s//5A
NiCLLejpQ7X9DnYM/eUtsXY1mvoBiGPuijUzPTTP397YVq5NpqXCxEKqOny/gXI1
FeK6D7Loq60mi7WVL3JDs72c8xOheSEatnD217LYRIVnu4s0jyYNMWwixYXUgSI7
0SI3RikOnIPjPlFZOJhZw4FVddUvx7H/UrVNwDVnU+CvT0r6VJ9jtyYu2RDOJqxs
uQa1xX0enOBCLhHk3K2P56SPI+D9SNVLvSrg18vR3w+JX0lbRMUM20AzfXpFJseB
ZehqIthvIWSCYlVja81qC03SpLh5XGuJcczsuQQjEGFUeIj5y8YbsmgEeAJL3VxB
xLrCEK7zpSQ/O1mG/5UI726wBkmb4JtDATTNKUfjeGi/V98Y8ZlRnjxN7h1LyTt5
1JUv6Sfd5sYAh/ig8jxFrjeBi4qQNgkQR+aHvSPWZsiSTtwIFw3ABd+8+YMPTKrY
8txBYcRKym5d+C/UzHaFksKJBbVIfaP6orkfVXzJDKU/sUFKa+oxTgf8m9COOsTL
AI/HvQuByeD+zk14c1HuaempzhNAUe3nHypM8MxW1SrXOxlJYTwvfFC22l1mtADe
czwrtyp30lujd3HJ6/q4K5/6f7RjzU6sA5yhgo+hOX61ouOUyHBAaZwcKN5KE/Id
QU0mWc8zWLMp+g6vTqzpQRjefzXNX8KwlAIH52xJ1awtBIW9KTb5BTMIr2fFhNhn
wo96Ts3VHRjMhoDkK+UrkzuEZ9FvFVWVpntnOBdfAVW8TGG74gTDGCrkaimD0d9S
qdmBpTJsSOai1Vtjz7cqD8qem+//p9U50hbOj5mkcM2ucSwqCsCVQBRvRP5YEnUx
+wccVZxaeQkDE3ac0MC0RDKqMax/xcOlESk+TuHUCgXz2nZhWRhe/Ojz7Xh4jcd9
T6o2k5Pq5GFXr10GCG9VI+KvBCw+wSzoeup7PUMvo50rIhyjm2It3ka3t3kRhdpE
lb7F7mT5f3s6/ZlOSTEXRZMll7uyMVXy0SykUo1dQc+x1NJcuSBYWST/Ip6fERa9
TZMQu/V7zmXBikwUi6AqBth7n9iCyrFlZxCRK/7JrYIcyY7LR4TYyOU0odcViOKq
8yOz+/aaLusQVl/b8GmQN4bvmzyGrcPiwMQO6Wnxo00yuMkeF7C4/ZBJn81zYJEP
Uus/POYBcUTNgqtXyCmWLnfFWziGgqA91LgFLPxM9VqT4LCd46uEW+922n2/rho5
v/uiVlW3yqb5UWrJUUpeLtzf3NBYRlWX76GdolVDlc7G+Fup7USboQSEztrDmxz3
+APhtZksiGjIdK4o7XAMSnjx3eiDcR+hZrQoMytugoSmIrVLxYIInBWHmKzEmzRd
xvJueP5/tNK6KNlBfWPiY2Y4Qy4dkSLW7a9L4fmkbH862RMD6u4oOIqKZElgTCIT
kRG/OhIlnbaAsDJ/QIj96hzHEp7yDwnox6fqIgaex/8w0q0hLiRVB6OeFBrYDVIE
nXkGNlC16OswFspJI560lBTNA9HMGMm5ebbyr6ybOvB+hR03cRil0VfmLM4hgdei
VMGOUpqCNFeDqTgjBFojyjgHw/1jabZa594B+wldKR4NMLvU0rRMa3hOT5jL9K44
66lBAKYReuAJMqmfo6fmK02R0L9goqEOLvND0Tpdi4pIGG3GMhW60NnkDdzQhv/e
zq9MUKIIdBNZr9fvC3dm9vFOHN1irrmbvVy6HFLm5byrioK7d+W+Z05vL9FgnGpT
T724VHYU8Xidgtw2QFwj4lIDoC01HjDosudN4YaKDpZLJwbANyez7g3J8ZgK1FEQ
bhBrdNpjZXa+F5PQeCEZbOmv6NCUD++kk3elaxqxed78iUNaAagsVJSYG4GEPA9H
C7THoBdZ8fxB79p51VVhTg7wkHypoR4x9GjPCRPz8ToOeIhFIzgOjNCKF+UtbrWy
sWKbevcLAqVFhlaTZJy60YIoOWcXUCJlv2lw3ORIYQS3HfIU0eQ3K83KU3nAs34V
eTntQEH7ymhlvA0hl2TD/CK3NaA7XWIAaBzFiuy9l72ags9SNKMNLOHAaMyYCUfd
1cD2Y2/pRdSLnsv/zyRbkQ01pgnNSrZBkjh4PQ37YYU+Zlb6jSE2go4dw/qjOXiL
hXd+OWGa3DK5ncnboAaAoBgUVTk0T8mC9wdhwJ2Josgjm+yvUDdSXkxyYQZXKlla
t8T20ilB3K4OozUmXUXKmWDqDVvREGWDgxo7ByRDRSubQAifYfDmMgM0IzG3ISp8
kuiuu6amcaXlz6G+Wf5Xy2RqkWiDLMRhjIKKf6rBnJ7IkK5OkNpeo1C6SUj3+vFj
SpCsRclJV/reWVz2AGjFZNVYeofK7K6nAAPo60KbTSapyjPtWj0ANAgyw16mNsDw
8MF9Ig5DU3pIOwe3H7bZbk/pDpyvwOeRciO/IJeDu9pv3UwjS6ZpQIpIv306Nykv
AxZI8pw+JswneZSCcXjaWHrLOHyFtXYT1299GXNA4uEF7aIarBfvNIUFCGO7wPFb
Jzs3mybmRHnOhFyF4d1fMAxmpA5BXNDG/mvLVB2PoydfBotNJLHlFAhEFQ7nw2N1
mVaP7GKab/o+nDOFXXpU6NQHTrxwnsFnX77fNOVugUJu7iKZWs+lTyHPwYqf6ag9
7807peJEowweKwRu7Spko/vQ73TPXJCiblbGY4H5GWPaDzY6Lo3d2Um/LI2IqwK4
LEhDx1nWNAF6MW8HQG2HE4recgjfAn2U0krqkQggCbPRF17m3jHEp6yRJg1ZY6OT
I+r44JbdqZYi8JTrx9DAuEU3WEUV+kAGYdVHnz6A2USZqu3REFWITMgRREfKRVDn
/kS+OfDzzbEAbF9ANkmX1jn3K0Jvd4b5eIUsq4kxkdC4ugFXBDgO2tmzqd8iKuKd
zKnBBBa9vgG+GbNbelG1X3l1U3y9/ZhILQwKc7gkXXPCvvQnTrOHH6dHJwgbxMw7
vRcDAt8u9spxOatNVkH8sE+cwPPFpVgsRgprb8I7WnT6NqAIwEK/j1jvmVZI/V3W
wHhTK+9xNxvthZMeFUKVKtaupCjMl7cZ6C2g00Vycawmc6f3rHYsH1CvvoI5HhgR
zebTZJvAu7rMlCsuNMupaU3160RWzzfOKsgZT0U/P++RmnLr5HbqjN2Uaho6kUDL
7i32pshYF9J5UJhAuyqddbboEBSLG4Du1I7WFiZFo/REXbyhAPMxt8goeKZEEX0h
/p0LkHYT0WX8CoD/dnT4u9QjkMuGi3NzfuwYSMgA4oZ7vGVEPKCSo31aW9Xax5Jb
T0o77mnkIjiH5pU/g3zn5DNe3JLKJcleQOqV9VWFONOsYGLUrLJcfhI397zw3cxb
mNjScDm9AHzWKFe6r+K/NTJYdZLNr5/WmSh0hYpMYIN7SElOVgBhffNQ8/yD80zn
K6sD7Ox4xc1yfZSt+mlhlXSmuHHgWpxwW9pEGcQkianlYg6Cscinr2OIodTRal4C
PVr3OwJE/cY0kNoOs8YM8jVM7fh6CipeSFH5dQArytDI9QEW0X6aytL3s7hGMLot
LoVJiWXH/oOygtYahDvjt5eCaOD4ERqp6ZWLPaKPMX2WCzExMH16TjunL4W41eUq
HiNQLrCHXP2Mc7j6A/6FoZSW7IybI3kITSMt7OYE8HCwsw7S+SOSyEPMcYnn4OYQ
8y3Efo3kjq8I695rDh+nw+mJZ9+uBbMzpkedBawG0M62DUoj4fujrNnM9xonu+jm
ys5xvaove3gAtNGDO09RhurN1M9LW3v6sWrh5sNe4waYNkDnOS3eERU8ezoHLuJg
Rv24hjRuKU+dSdw/RgZeMnmFPtee8Qy922GkNfFRgu6UGik2GcPz/D8Gk0R3Es/i
pEqSANiNXiZ6QL9ovm8qWKs+OwuR571Hn9Sf/6towcoHrSOaHDKJPiM3BuWAsxed
zupk3a4XQ5JzBOmKlZqlvsDlVFIaWm40768rZcJ8e7WloitbZfWetq1fmH+tePeT
lb1JYhoINLnLOMPi+aPJXdSLJLkLKxVkgmgNpgGwVk3gcd9x1RxyRwxJoqMBd31V
F7olw1YGYScW9bBloHG43iRkdJm5g3Ig98ZvfbqUSmbUm6zGtkexm8v2iARDc1TQ
ee3g0uBNNdYMFcTlUCURAknoIeNcxB4XfJ4i1OBNaXZ7jZxuUof56gEWA4F7yKV0
CUlbnvP8xRJVu6XcqwtTuaPkTeQkpUMhYgeMQMUe2J3bHGW+fC8bduJqCbTDYpoL
RcSq8T0UIrxUiECVNoIvvfQe4JT2AF5y53HxHwKA6TJTTB1XKKhU6pwkTMjYjhUf
E4N3SyQZwzgvWzJbfFKy9GR4z+Khvw6y9YugVg26Ex5tLVsL/Vx1vrz/5Kz+6n8z
eOqaAebWNa7cqzNclXTpCNo50/4uTEuLwNAdPNfkoXwHx3PnVsp0aTtc9csgDyzq
tDVEenJAiRDV/ZzEUMaYxSZvDA9MFr1bOVuMJ8MuTSW0pl+iH96ewPTitnZ+9YO2
EZvCVHwq+Vt5da08BgiKDRBmSEfa9bfV6TMNhN1Mu+kWHEJW/OE9EE7LnxsN3mBW
2tK/8KCG2Z+Vxr69T2Ttt0wsZ6CpPllhOj/tPp5ySBHBPb2DUHS7gXOJ28QpIMDm
C9cbKC8qXMwfsXVjzBIhi3Bjsr0aiq8INVOYjQuWMNj16x3J1t2Rauw66j5NBe5T
unjckjRLCv70tbwqtjNxWdTioit4BNvFHHhrhzTxQ34JXhAToSyIg91BytbpLVmr
EH2VA6+/tnlGeD8demKYFpXRj02BE3aj7VOCL0b6daNXbCcndUjeqEyq65lNktHW
L4XNuxSYw8VpV+MngSun8VZWJiHolPYuqLMpaI0zyiY0UU0FNuQ/zf/s3grslpW0
3Vherx6BLJ/mMIjcdkeopxIIFNPQdSBUOe4TKMOkoAxKC3qy/OZQQbCwpTxJFo0a
c6rVZeXnB3eq0SZmXERmJ1TrBFU9/G2BpPgIqDUmRYzQbC41svOj44tc0bg3K1hI
e1zkxV1S8v65yUJg8jtoJZGcS8wAqvNdzO0BWkg0iS7/ZvurenncXddb7i2VUOu6
3AQse6OwnsnbrPGOLGLy/StKN4yVRPuoTliPCT36Gtj+/gResG9iNf4fMPgY2PRV
hQVDA2HDeJ1m9LUiM5Crut5G1uasrRER4EteN8OynZs/QcM40zaULhjXhFpTh/Ll
F7N6YRViRtAJy4pXgJBiKqEV+nyXWTahWTjRnXFbgJUYXZa0H6u1VtFJIh0bF3UY
3JJMjQEdz33Sz+aR350NHHkKJ9akuPYM5TYDKeFj1VDY03LU/2fbIzmIh0b4B3bd
D0YHYEP9cx0KzAJXog6jgvIREsMgPY1zVUUYnqaDUIOg+E7Y1O2aoMbL6Ym5BQ2E
NX1eNYgAKmen/14JRUXwtdICuVQG1KOyWuRamehIZAUP+g+CE/8SSboPPItjkhZs
oy7q51NIS5YbuS/dvlSd6/GwFHKiE2FnSIW0/Rm6Ct+n61pXFfmC8Yy7yvTNE7zV
jP8lR30f+OfjLJoQDeqkuR8a+OhUjv2MPbIEkGP7onTRXfyfmCI7KEgtGU7rY7pH
5VdEZgsH85P1PAJwwGxnRXNyXFvGmywP6L/Uud6t0loHQJ36HwFfJeoWUhJSvlln
PG89m9liARONM4GajpSR6r2LJZQYhIUM6EjuwWco/wGTX5JFfC+uAicBY4rcWisK
PiSAf9vuQe5LVew186ncIVNQhuuN/i8+sv3QACto5tnIiwiZoi/9L1I0RenVob5k
Q08S6/3jE+x1gCUzC9tZ5gp66XPkbMMOdjvHh6RSzWdf8NSjX0OYAsEtsrJu4Qid
TMPJtFCF9bj4eBrSSn7ZrUqm294Wo7+wJAYqVGAN/MFv2iSulxmc9TUrgb1qdgGq
zNFq2KYCbHUOCE5LJqfuE/QGeG0VguwFvNmoJkRJc6cb4GUur1zAN/b4aCaeON0u
LgZr/dKGNs0CVAXHdq2E4Tuq+cGpR6Gc0r9gd2dDosljsnPF1lCzRwFyoK2Wsrd1
19m0CStVO4WjqMkJQ6WvR/8eb8N/LWwqxIYXB6F73Jyke2uULhS5foGxp7KLw54w
Fup+eJF/96cf6T+lbl0X2lRyvgbwnyPxSTQ7s5nVC40lbAwogwwiSjxnOaPjpyCp
2Pbc3mkGpQbVni8zUvQH+PZwHMz4FtvwvHv+rH1vJWGsz9EeukaRuk+JalfN/1bG
6XUu27OeOrWUeYsxgmf1NnS/B0uPvApZCXW7v3r+b3wXyKdG5iRqFUzff4sFgXz7
PkVIW9e65INxUaiVYnWzNPYgqWw5jVGuv69BL3X30yAsVTb3wvMjybDPx5Z60sba
gBkM/IojEQ4b4v6TinxsiVPJXpzxkTqGjGuZqqJtB49pPRJ/rRK6aqjs4N9lwySl
C04P1Y3cP/9Dx/zsBmu198qa48Yr0HDJ1YA3vCRvHvKDamHQr75lncYPUL3/MX+P
ahvIQibHXLoUXc1kuP52s365+OzcgRCkT3BMw+7i7n6QZw4VzrR2qfjSBByJl2q6
q9BwPDIZZJKLIp4Vbsm+wLbG47OQZR6pU6neNpE242+3FinPShR2tmbqvhw0P9Hf
PGDtfizItfIMiu7Yv1dCEPkiVcUMK9T5hyBT6s5eenHXOvpqO7Acf3fFzN0RGkAf
bt+SqgdZFXJKP0/wf04qR9Am5TksQAOUKhXa77T/+KJ0i8iNFHw5IVqdrpBglx8k
UE58lKotX2NmuWWOMjDttdoTHeSdDqI18i7VzmukUJu0u1WBxbPzo8QPfcJwjQmB
JkoMy4cqmxY+2xJZHMYjaczeUN5ShNT0tAxcM9tP/UKwRDNsuQkzz1yXtYK4wo6a
FDuHT1ZJOUQNGs1td7+aoedcG+b9UI8sueOH17PS3RgAsvOTuPvBpWe7Y1hkdZqc
2SJ207WxfBY7s8phOU/hkbB1BmAe52X67MQ4U9EDFR3MXHwB5hB+mN98ghjYnxfc
FPDBRqVV9cHV8rS+87NZoTHUzQq7ot0W/LV8ZPr1BUIKzfvhOFeOr8rPrQ7yvQ1t
ZojvorAa0ILPmjJJqlSpwDlJhyCiGpkPiuLsxejtVxGPx70/hTeH/QJwjMVxf2Dt
mIVV3PoJbkyafWTfF8mX5IWVz4f9txaU5aWJ+TyqSPgxXzw/+n/v70G4lUWMne0P
Erfgu/T4daUJvaQg5xZuKijkgmmls8/l/od1Bk/Vkd7HBSVH5I1FW7GQ4NerdX6U
SuFt1vKBSGLD6NrsMfk0of9ZroJkLxNWTUuc0vPqjxQwe+9H2FaRiKcCkwj8pbSH
qKs0f+deNkYtTc1gWx/7rs4lyDzxte3xxNrsCc3iyHb3mdmd2B3kiD2VSdbSWgjA
bKhC8iJOf26MWsezM1RKHNxRK9ZzsC5J8sG+jgERFTN5eGEMvkbB2GGSsYUVLHKs
Uqh2Wl7L2QvJJXyJ9DY+UaA59ROzbivE2u6vlexf9CeH7JVC7ehJBAICpywOXz7B
q6TLn3WY5fQrlp4W9mXYNeGBqyLjZgIM9B7MAA//0BQ4WDoMcswU7Tzcn5MHV8hU
2WkGq/F4v/aSQ4AdqQQ1pILR1lh/HC9Fm7k58gYE0ur/Lnsm4MZilrk457Mt1Qvf
tiu9dAgr1+1L8gX3+/qGHO7VmOq/tCW8MKaincsjkqARMnET9o+DFuwWdKE2yUJg
iXdSGhIeFHOCZD6+xFv0ZyadFSJCSPLXMmBEf1XsBBRL9AjeDXc9IyQtJoKR11tj
9mUtAK6jCfufLzT3GjCe+liv8SWel8Oxykz/VUejZ/TAhMc/XnScbwadYAFJ+Ys6
Il4TczlUuxi+LSQkrJxwpHB/FWO4/VXYvWgs+k+j4ztqIc0O0IzX7DwCa35IM1mV
1CXykDw3zepECQ1qAbtKsmrkMszZwd3s720p+PIWrLN4EeE3ieJBOEWoy/sOKboq
rFNjJpXnDfpCx9dFGav0YRd+3R3O0sl3OjHyOL9pg+rPV6Q8nIoHtkNNNX9T3Tog
tNVJIE+k95gRmLsp7DWfeNwp0ZO2ybNiBO4t3+kpy5foxUiP3SLoIQ8N3WPr90EI
7U0URKlZ48DNuDxIRZiLCcdNqBYesQrlMn91uK9C2UMxTFYsM5JGUS+Dd5Sd/uAZ
5L+ATP39yxIcy6oLmRiC5lRe1VKaS4ClupoBgkdKOwfw1d5RTkf+F/UcKhdRBE2c
tpHdOguicmbRHUNAyRnWiyoopSxZmdUphUXhHS3Z8d3CHd2e5/OH7zNgoHM9eiYu
jkV889zBicL6fcyH18UbHBrSS6oq34p8QltKaeoVXsVD8oTME69Ri3elyYZLSwtO
uqOGYf/+j50IU69XdgoUvOveEKPdu88UBjBxTF8CV73I4KEPVSl/8oixtfAQWqK8
JFwZUYI/lV/MFsFVTonzt2g7y2B87CZiK7xjJAWZ4DQV90VF9MU7nbqC1ljf2D5R
tg/XbnLdWfsQT0tFHp37F4Muv4smEW2yFrJZEzdSB/Lxz+qaEaaKmr3lox+PYFuS
2QhcxgWTeJPFBkIPUC3bZh+E/mUJboW49exRz/ONE7dehziDCpX1Wcm/rJYjEeVr
EhbcrdpSbYkELwpxWZRqM2bBGCKboDw5ZoxMws4kgOwEk0zxnlYtR8y08TqTvWSh
LoZkJPzjP9rwxGskLsdYtvud1kXmAaoN3ouQ53B2C1HEvNsBzbg+HhdC9Rn/fjPC
2jx4J4VF69lp3OAlbZcgrWd8HMaGmRe3TIiJdCtmTixeW2RT6XnjddX/J5akzvMc
g9wg0qoyiKtJF01pMXXVIEcaQFoJbHYPpE/5kTnl2cJJuKgrmv/49Vr60CUZaBaw
X8AthWItVqTUuEH3BypxB1pLYo27XaBhhgFi0n40srq+S2tOHcXET6NzzUdg8I8J
Jx9NImUVChnHHOuE2KanR9qSP9o30ir93qIxsmKHeBcAnjecBFfaL/HGMdqcPtvC
1siA2K25Bb6z4JpavKUHHNXsgQNYCsQbVaVrO6M0Vmp9MweGbD0mBpWofyaH6oHI
BhvWMayRLNOcsk2Qyygxrn3d5kcbsjTbeqY+2wmj/xV5cRV/1CXZt+sexapslPj5
l8dF2sPQORghP5s1mWVNLSK3iAqjr2XK9Nui1oEapwhbOHmsYSfPJ/xkSpTwQZEK
gPLVHtDZ3mwUsz0D27VktKjoEvw9+jJylAmZ4m/mTXGy6EW57OirlqWYTkDzlkD0
iIBc0lGb7s/Q8nFMsP5aUHu23W7wbiezzbZFbsmL2P6KE5t8Sv0uXoRj8x86JFwp
2SbYw2KbSEfcnAB0mjvM8hXHLkpe9eJDJ374YKXaejII2T7u/NrCnmXo9WX46ni0
INZbyD2csVwUqWV9aODQM05C26VS2CFBE1h4SbEeSvtOslL4VLU10fAVG4XOZSvn
9afZrkRaGd/oaypJIvGZGdvT9Fi0VNdDzp5LaARVUyViMHV1eV3o+oHNVIpnnLHr
tVfrEDkpqP58Vn4Mz7gGQFPAPeO0Wd7DH/KIxEyP7ez5iyzEt4+K4TypH0n62rGC
IItAQZ5QmxT2d7zDYOd1naazhtgza2XqgUZtZl3zzRzGK0Xtm/fqd1EGdly1hNop
rkBySnqwG8mz8uty+sRMCmxuF5k1vMnj+VaXZcATxvYULgZwSSNW0WQi7DJ9kS49
a6kMqpfAmy6dOlwgVXGJFQCIyvU7nf42Iksw0QFEe0tsxOCuTQvn/1VhVpf2PBFL
2+gkZM9h3Auj2uF9cqR+5b+PLMu9MGCeoHyzvKMfvye5yv1wu+Ycc6EDW3IU6sa3
8GaT6x8P1f54DAn/i8RwEgfIw5VJxeFNdDUbCYs+rqTb5V7sJoGVdLEbPWu2Nw3n
6KFJqjEUvAlHftB/oP31+iD7qM92/DIKJksdyHtLlGh4Lv3ojbZBSYfxAu/Ll3pX
JPMKpD9u4pKDEH3QsnInHi3kKsQMyP4eArkloft9DcQruaR9yYA2TT8m8cIvjVuD
QFhvd4DdJbL28nS8rkNQ/vOEscimI9Af31OpV+8fTA+LV/b3iI8ORamPz42W/59R
dycEQLo4bCk1PWwUaOjY+y9HRehGvopaqB8eCJcxSih/dzhOIeEe/3UKUUkMPi3y
elC4KbiZ2AeRPNB1MVejHY6PX/45qYSGBZL/87XWmlT+MTFXinoTzIQGe699rKUO
MIdXFnM/2+6xcCvyd8o7hWTAAi1nAE7Il3+NWH8y3PsMLOzoBPMto4zNVRipeHGL
Mvgr+HOY2LnoQOMC6AOteJRZGgbsMCG6FpkTPhsxan4CWiJt1e4NygBjdDTdzQ8x
gMOqg3luZHAkUM0K9T4aJAg4PsVi4H0g3Av6KnPa3gQuoEsT6w+DZ5rS/Va+RQwI
1zCl6uFV0E4Ygv0KkrO07CYuQykn+L0ee7Q8tS2kP1x8BROntW1U+O7nDWdDTNII
2QBjI4k+e5xFUrbq6uDn2cb9mcrVVv0yc9rvRLOCmkyJgGuQ9bC86uB7bmndSOMf
GjLWjqWdF0F2play5s/ph1lOPXDID9mSb9e3gSDl48WW+l6nyy++4Nv5cO/0jAbU
kAJBEUx+4aI7/8AXy5LR15lsNDGziBEFPisSUf7vehW+0u0AV21Jue4R6mFd+yj/
RJgunMt1905Vd+dg5eeHe04IguulHhJb7Kxlg4WAcFDyItO12yW+rMbzC5f1h4oP
R16Q5MUuBNM6xdZFD8leB7bEr4HekyrgDlKjqVFyK5M9eq6uVqs2N2cCQEevd82c
z7wU9qWLbJ5ZRD/dAgzjOv5kel9TVYOfHjQJ2BcYTv83DCrkjaRBa30xUWt1UdYF
Z1eeceY9zURl+FsbHYzbJX2YhKwzOgVAjmlVcguvvg0l8vAzc0aV+QjeLRRi3u2O
GBY75YMZCWCQsfXTF80wqYPQowpDiVQQhBqSmad5eV1yC5m0QvN0Y8cV1g1WSOsq
JagS3SLGApdTRahFUZCy7oPqx3yP98ALYMksoJHjmYYW/3F2gVlByYB8tZgee1SX
6wUYUEbIZ4z0dRRCrjpU3YLExyJ79OsVCCv7LzA0PTBDOxxccZvcvs+n4PtblVvx
WZulSgZKiEoFFNfrTLWkjoeX7RqYsMo5ostX7I4ZbMY7PHpuTY8+TJ50YrzdATcc
hb8iSOxaMC6PQNahxBeW/oYfa8GwL+iTpf3+jMTLy2+Dn8O+Wz11SAB2CvIcHeUL
DTXH/LvAQObVp/1NQydEw2aCcQDVnqrCkFpj5XzalxEvGN/3rMyvAwBBDindx5EI
Ci/MEpgC3VPWxXDU6vVoUN1vAZo9H8vtJFFs/+Cd/fVJQ3b8vcGvTelFBcs+XKsT
SazFV7/Uaxmtdg4Ssb3KcEVTK48a9f5bcpMOjmqWjB7iUPvHtKozEiO9R+X0qf09
pjH/niZ8MyAlsdJB4EKKg2I79EhFZL6RRV+XDfbUKd/F9qWaKzPbJ4lXvbXAXrxd
jh6c+ggDUL9VUE2/8OL/b/Gag2PFeLawNElzX7qKGcanrHeln4rbjGxrHx+MUJOk
Am87viNYAHmvhshBwc5AtBhLxiS1nUvbZ3cNNEig4Ovq73r5kq6BgWxoRE0xeXBJ
Ln13iZf53ijkEBnoDy+BYX7CLBok82OIzZ/lxWO6rtwD4ttKyTbMxSBcYStLarka
Yr5gaBFswxCW66vSB7ZS57ieg9JALSsA3hYyY/u6S2EMlGgAiIkmCmV7dqJcDIUT
RnpoR9bPvWGc1MjEEP2nDGxMJISF6HHkAd3pWp3HnyZ+uPt/ePLFvVn2FfcRw7gJ
g30kRVJs2ZIk66titrAXSHGLZSEUCod2G8flknAQOjLP1u9c7hKhWxzqFEe+elke
ti2DsMcYWyc88e+Y2T3UVslC2RWUx2FMVhI0dPq6Vtl/L052iKbr5nwbai4Zrggu
3dQRfuRNcBFtO0fumPZNf7biVfn9C8X1umojU3uYxBJRp2sizEU05lib1RrkhriF
2GArUBC3nW7YV3oFGg+TnEAB2YSN4OMwrNuosqotxsD7zAyuioiCf1oWtAjkXMxh
vMfvb4asW0++dVs8xUm2aUXxBZOVgSEBL4te6L+8RqM326b8Rm+8/RqoOj07QJ5A
PE1ksSMiH7cyW7rLIR1BImFYa42Okzu/1H3xvAtBFLbcbwhDmG62oagqhP4JE1By
wFd5izfPFKBy2SzclEQEMXwl8Brl5Ldz8O2oWrt+a9R/FfeugpdQKUDVUlej2X85
nFoChKQFAN0JkxDJIvCereyiHbLz83HTMRbvlC0Dw36Y1WzLjGW7f3IYo2I3iKPC
uj82WGLYtkWzxKJAIxC14zVKUZTLEfodPiCrA3IC/28InpmdhRJS/cXJJuKGaA4X
vJSfuXbppzesUHXn3GlsbDVDFfhSQJyrRaV7a29UvtvCZcQVKCRWmysLE0wOdhws
ABbc6AoOJSDuFOrbG/dEQwjLim0jqTSzVMmT4f+TEEUUKkhHtuPDUbZWJaXvEw8q
MHPSMjljFgLzNFkkkf8ZAhxzuQ1aJvzufFubJBQV5rI3IhkKEwDW5mKaPPsSn/94
xvzkMMUmQtXT8OMvlVt7E3BG6DPv7UgrlUM1YM68E2eercQaOKgfZoQN8EmExXTr
ZoqQ2NPPgKFamPV1G+d1mHJGWe3IomZRpQqD992WsPjdjdgfbVcqvGQeS/cbJ7Ls
Zz/p9mAlLj0PnpONnrpiHub1E+TglOzsb7Tsy/G0RV+ztUeKTWe4iKwp5bSlfOX6
biQZkptceJAMlMC1sNPZqChKTg4zXF8xJLV7P8H36S/gjeZ6yq+TKbfd9mBe5h7Z
QnBgQFO/KAsspkg/PewRpfH7PW0f7mNbERR7/O+UkdLbqJRGlHIztusIffCZrQAj
lZYWCvmPFseELse0QOlgI7++0fn29nuB53wXgRrMsVju7XOlaGKm3xHs4nn6i8L/
LH4nKJhuKydUhw+LlFzjhuBB+TSdi2jl4BmmfSjmnhB6v8SM+70sf0L0RVZzV0ij
cVgb5m0sn2zDDuiMJ6y1Z9fQ6YSDvFMLRSrIMvF8VF3HFhFoQM22s3dtJV/aBo4G
8PbPhGGgjK1CiGgNsHvktnnQ/4X1+TNUGEDaCqJyawe+800eOZYvNjzWfkzWBlBL
x3busphc6HOzwxMj+5Qx9AQ1n9rxnpIIkwntek1Uuemviv9jwl3LI8ShodNZQJRm
XGgBdOOtPN+YK1FGtwPuGCeo0rOWoE2fAO1LJqbLLdxd99rBRDSlzgzf6SOwaAra
/PaQbFqeE1Qa83ZnHb8ZZpBxRQALhHmv+gXSTB1jXwgj8gDAn9i59przzUpI8qb0
+q9FKK8O9P0YTfBvv/IlVArqlqIqGuaUK/bVuhEBXSnjE6sHz146tPAcSsPI1BxK
TjedpEJAzuFwQUX9Kb7lP3QDbf3heBPjOZDLbdiWlsZjADGOmXGQM4xK21sbNkhm
Pn3dwNPmUYhhxzFGQ6uzyjDgF9EA1JgO88UrZE/B0vlD3qeT9XK0FNg22HN1/7Tn
O/FTI2pGbfYEO3zqyHyIEQ6Qjg7MTbs1+kYkxZgZceXHpqreQ0371Xbzh4al2jet
LKyFy4AtkseCwRKLiSfwSfQPK2baGIz4zaO+UhADoOuBGIrw12mAouykd03vYu54
Uo00FEUKQ4fbIJWxJy9NosL2GRUjtKSR0GGDgT737abvLudOnDxDjLth1lEs0Mc8
FxVNlEX98yRGuPWT50oU2+1v2pbUiBSvvhjXyDvNBUMlNKmw0CNRs4mgo7FNhL9r
PEMR3jDixo8zWr6PQmlLaV+osVL4Ib9Df6kqSq+DsUql3+Wg6LSXTIKp48kcZ6Xv
BNJZIp+A8dp5v4UNw4DDhT62U32Szqwj65571xqDuXtNTXNxLMhfAlHULa+0suw2
gJQYNO+E3+TZkpGasH/VumGrUDKAcwXEQwmYdMcId1tCdrbv+ekLq79uKKb+2cMu
O0d5DKWxoyvn9hQ+K4ZWmnn4/35Tw0RFpx5xn+T5g48t0/8xlEFD4J1N53QafrAi
DT0yDjgHRx7yS8ED+VEX+5lfWH5miOW2kykDex8br0YqFC9QwgLleOkr94UqO9F2
NPQtqo+7MljNrG7FZkvo82p8GQdlP01sX3CPWy5NEN4ajbbMugpxEFApSBXlGrLH
xpuMteayRYv6v//kBcNCGHlaa9tOLq+1KQR47vIfRXj9jBNNrDwIWhzViQjwZSKG
g1dQ08+EcQIXCJBjuhxHwRojI0vDUBYaO1bhTHzK3+qM+EfV2G30xUmjXOND5H1/
nr/3rBXIidAhKD2YKTgRH0XyKv1xOLzsPRMdUkc/kYD2QZnyKUoXTuSNBLJHSuZV
KKcJDuUlTALTD1UFb0wu9VPcmayOyBfNzosciUFQt9StO1nCCpJDQfCX3YSylfWr
Iono7BG/QMdULmoLn3LT4fmGYJLHNRqt0544Q5xBYupxelDIvefUaxjr9hhUGY88
y11KgMRUiZwlP1GCU8lZtYhaLBffpQ/qqb66EWPj6MHQpP8ZGD1ISlLAOloV3rsB
Wi6LjaWzNHzLajyGzDrRmz37jee1R3JttVM0RCqrOMHPh6UIYYzcAqRcSFkJsjvk
/cols4ob21Fsj80l8GEwVil0bBiG6x8w+pzIyaMOD7r/AarPy8HmCZh2AYA7Jl7E
UK5u2nvkuLJbnqikFHpZmLTiipyj2sktuthqMdMNXuRQJUkIc5og/JPV1BIcmATv
QDPy1CNuLdujUBmgHxDH1E47CjTC/qnxxne8kcPUAWPxwZwOWZHNGsEIntLQo3w3
KaD6gof5blArsmosdsqA755Kie3zS2jF7W2xObCi9FIKzbQM9TceXgw1kfCFrOWx
cu5TH3NyCbKGexlVYaBfpqiuDuwMF+EQyZgvYy5PWxWhYvp4d4DSzcMIxK6cz0bA
/tYerxu/jgyEtG4jlBSBu8fdXxRVjL3KbndgflNJi5B72Spg6p/m0WoCWlB8aNCe
1/WR3CqPRQGPWdMuWU07k2Xrnt3TEKFiKO+o2mQp2uJ7IbcI9CSO/128LmPZg20+
lN8ulRYv2O2yzYwxZH3kuN/gQc0IBBZndJlH33mBKb8m7LmkHrxaeQfvNGcYtarJ
cTx393CHH8Zfx30h228WfHQXVRA7/bF4DaHzndV4ALwH79rg6Jjt4xqSOTwZEWYe
n2dgXp2LuWBAxxmCU0LymVKt1WtvmvRlEr2eWalVQuDsTWOI+vKW6tZ0n+ljs9A2
9ig2hTI2jhkOBS2YBaalLgK1KJLp4oXl8uickK80FiUeflDP4uUTS1i94dc0iZBs
dcZ60UgMacg/nXPFH15q7MC/V4gVpkChCjVMBodPJB2FLcTikjpbYvIAhtV29KNE
MHUobEODGl8Ex80AYO9j1U+/JVOZ3ZDwYNGNxVW/+Fr++dGu5Bbe2s+edCWRnSWl
yUmQXvijfjaZHSZ3me28ENOr6LoVtPM1STkqR2QfaFh+L8JVbiOfoWk/5V96NWoW
qeKjAuEZpATZtGDOjuzbVEAFiw+QmuQ9FrxnXKymFPSp0pLQ6EvnJbgrAhta3JKm
LsOFfE8mvHsGyrQickvKeD8Lq920a1INI03qakDMRJxj4EDG3wBPMseQqAlwUah3
xeIJheiMEcoW4+w/D1S99VUuWsWKcpD4FN769fQCuWk93PSv7q2CCrCWJtgrtAwT
7ZmrZVJ9HaBEdnGJIT/lYOz+bwzhW9+h37hm/mG4e84Wv+NuUCZHkfNI8jG1ldIB
IwdSOc4N5AXRRIbGxGMJGmCJAzXP1O7EhAfG4DYN1OPD69MFj15bV3Xe1RDdyn9B
JBozDtWid5NuJ94pduwE/nDyqKBwIPD5j0RualHlLcxzDbKrVwAk2k5XiuWzh8i7
VtrizbtxdcGgT5woMalHntF2F0AATu69BVPzB76osf2aV64tgWZ/4laWvykQuLbo
aPDdglG8C6sPWpa4j9pcOoywvK6Z2BFDCzFHVJmufHnxq1uhe94Yc7uAgDcQKSdJ
Ekq3A69Q4RoZE9lukaEcQ+a1izFQINvJoNYeqT2+foHBSjf8Pc9JqMznqKrikVfL
YGkJCyf93O3C6G2almNIihUVbuW5zT6HbXn8Ma94IXqc5IjBPEm5U59IY3maAKVP
RY9j2WRhslt6hvOZSmPiP+YA7TeeII+cHmp5EJgtewe2U6yrr+XFpr3tnDIwywKz
AoyG+BHk1szVwEIset1vfdAZB5Ujput2UdSzucXioEg6OCDVkQtzvXmt+rjHkGQn
ztkasw2g4iUhtbskWHYt54rKIDOfovv4uJSJUWjIMfYVVzaF1vwlARL1HZTyQ0k6
3JnSzl9e7IGJU8mCqTU4xGM2Nss1vZUhot408X4CLjb6Ksq0aKX7CF0SU6LQBj9E
jjrlgakpT5UQgI0QqOPdb/aQRyLW7dHqFDhrUPLQLxSxKt0sToRes/Z9EBAoM9Co
EoTgQ3E7JElEOAGX7TeawHOairpClPk3Hs1ES1R8abj++P3CgXaEl7qjtvBvJq1+
//iBk5md+YV5NBE0Gh/bIrZiZWfjaYeMKhZEnOBgg4FSgLDPdkNPqo0hD5G4+fXt
898G/QlJxMNbRb3swzkjX/U5kRZ0zpHgGbblHO8JgCd+Sq6JwIVi/rflZumzIfci
K9y5Z+TKPGj0+eLeMYZc1JPClPfYCUcxD01Bp0exOFxmjA9E09OFk4m9f+tw+YQX
skpdEPu3n1p3p6fqTGQ5WnGlptWI9tDK0BhHHjSWpUjutIovbVjkOs9mucrrNRCU
X9qUJUv8hPMItXG+I/5mLJTq3LHWcpbFw+LMR1JLHfW/bqZYDY99n8NcqnbMQOWj
uGV/9AhumFQmjj3oX6pWUiz3tG/epoPJfDZjKpgJ6UVJqyUkepNW1dhBLN318pbm
JpchwrHZdWyD2KzcWeSOXcOICniAnZytRIVvp2uL5WupvKjjpziYXJAVeQ3JQbMn
RuUbGO/zzUr5334OT1uEbokRJPUb4kjfkMkSZB0FWzOxeXqUMPQUfezoxq4JGl7D
q/YsT1WbiY4c07OG3BDk//vsFq93i2owzC81pUYz/hMCC14BBZRNPQgypGve0me4
WJGrDwv9R/VZBGu4sJdIYbcHVK2W/MGrW5rb8/DM2hyj6+oTsP/mRupobbo2Vc4J
OL7rY/PfVKslZxUrEJiYVRyMce412rJpSuvDfIrDyTYpcqXgnGqNV2vJUXpc0Lo2
+q8c9bqFK+/CVN00Nzad2FDpex0ktC9f+yzTR5t3oLHS/Dufs20Jzh9xlXPRkeEL
NoQbhXaGQy4z3WEacWDKd8G4BLa31IFcyFIeymiWRQr7GHd8h8aPAU7Sz9RSkkdw
S16izsksEajxCVotCfAZ3qmPM4vsIybWb4DCjfkRvm3H0C7RkjGxma+1u8+YKUlT
6w73b0+Te/vKz5MVKGtCUPHpBP4XVUEK5Bb9hZaDV1Tm0JlADHphz/JcWA3KydX+
Aci8vL/1OLkMa0dAdDGMACcXs3KjTpaliGcYZxEgKTMUqZJKlfznuYhMpPlOCqBS
uu3CKupVwSZPw4CcALx0M47rLkAIaIpUjvkYb6CYxzf2n/sFBJnXaTvtG2jEBVUQ
rE02CS81EJrFtp8wssv6gGKYvH3khUkFHp7AxVKuAcdYMt7Q/+dIHFj7h6hxyYGh
Zj0rubby3SBf7vlI1tdTv63Crniqd6Qs59G4oxYxN7I3iqCQ1yLM7IK+n4q9spZe
/2Gstq4W9nzgvqbqnbJV/uIwrzvuYT4Tvi5KbtWfFA0S906cLLjsxrZcn6gUowD5
dOxNqSTyh9Bes2C2TLTlF3OOI/tWk3B3gO4mCR9wPM4Z6E9dzSPHuIkkoUQOhFeK
jyctX+Xo2iWaiygGlXvseTUAXxnd38JR+k4Ftl3V5IczAbZtH6sgTXewVYIafSzB
PhjoJCd5i55pB6w4kAIO05JfiwVeb5w24+zayeSm+xnmh4XrAhLi8mx5EuucC/7i
01G+UDIHJcGo2C1Uixaq9EKanqzIt582gD3FPflqsbvEr3Xb0MkUH/vEvL3oFlC+
6y84Y/nBLeYl1/Fji9KijjAqDBxo8VmGS0ZCqxiaUbRUxSxxC/GJdwlIKH2FC3V3
7LslZ+MDUESZTnWSsfagM424P5CtOY5NHrDD9dBBZmLy1LSt3+0DvOk/piqX9ieS
i/HmVgIxPsAFGAJAgLEAUg7rzToSTVIuyLdj41ov1T9P2YYvIFJsZJb2ZtHQ04+D
fRl2DG4fYSx3zyChKCZt4Dj29/DGp6alUcdBlrBE5x9BwT6AhRUxOEr8J+QlOJGn
diYPw84Rti0/ofnnn7ccDhodQAwgUJVK/iAWwPn9NMjcor+1Q9uulBEKWDfhBnUJ
SYhdKkSo6ITXOZAqr7UDCb3Ndl6Io06GOZRGG6VSsm8t5Ry3bk3uoty/PShvoPPl
YbaWrPy2sObtF86P3B6Lq55CAKMqkhHKWtb0N+0sRWpnlH8/qRqNlm1sLTALZnR0
tzl9v7eS38gT4F3BTRqCxpaMa7TxNMISmjU4P8K63H3FiMN+OMX3bPo1IeBgTqoM
z2yD85HwEwbDLvEdvgcY8IxG1qVYJ5em4MvzO5rHcScgaptRzRL65lHG4aS44FmV
bZSkjfgjI7xISynHzeRuzdKMiRkTn56Aa5tu4AlYkjsdED0Yp8lEfYt5qqnl5PI/
9NjvdBoy1Flxji9pRbkNhtefWatkS3mxXXMwY2tT8lpX9SJ3csm0jbsq8QQR0k4m
lpoQkVyyc0gjpgcWM1lIPzDijg8mh0DF38VXWlT2/6EqSWqXVEjq0swXxX2qMWL3
wLUf1ixJ7qEsRPCzL/vR44x/D/WK7LiKkyYCL4jKiNOOwHmhFp7nFStIQNoAj8Lf
CuAvrrC9u/Ts/AhfBjUgwQAnQQVxTRRnAZ8PXvD8G4nXjIX44521ZDieHcJNGgNq
JI18GdgsSeGwPqzu96jhT3wv1W9mjjNTpePf69WxFrSRywNG3mOxMPogejWhLOkg
oTpjHHTFeWsK47WG3EmwJN3v2D/Fyul6t1tShZYM0VByiPgd2VHgV08v3MbOmmEc
1qAyZL1CBDujlTQ4vGr4Hsp4PIhR1p+fVX2tV3gjZP8QUyDf/NOOuF+N+MYqmPCL
pyYayCD1sCEO/Q6r4DKxezeWLxXWSvK1l8cJlAF6XDouucfoeHE9+DgY5CZYBgQV
yP3CHCLFdVhn56ysmlkRX1iNwIU90naH18THJyXCaiHi88UU3HbQnVLHdtrmEuJa
JwZ/MKYZLRSGkQ9TK4cJgq/XE8GhoPwsvswnlVibSZdFUa/hi0QE+2V8yi9fn2Y6
hRc2C2kSrpuyLiT0rrEVjw4fpXDnQCKcCHmT5cOmz5PEnzrD2kbKwuivti08qYMg
HGXuE+Ui3+K2j6fFxhZaJ95v753tkf7FrDPx0V/7lwHGPOgVNMCyXHG+pXh5dJXQ
xJGOsQsdUA/p3cFhlKVfBBWOJ4IY3upJpYKAnEvep2aHDmS5L0qOEPPflx4ksBFr
rt2Jd7RXedm80oJ6NgYgkgiBDJamRZxWpDa/ydcK6SuHsOupt56kSdjHbD+NLBAZ
y4x5BLvAG4iYuUIdujsD7coH4YRkeOVvB29vQRnlhZG/4gHFjL04VY4P27gDGH5j
aBjpVO6pXvIzkZOCYVf+Z3dNU2nG/huZ89DpLb37ncdk8BvtT+p3TLznMW8xngoz
oE0vjm/L+jek4MtkmstDznUILcuCJkpQVZMcx3qyniEj5au5Nwwk5E1zZYHk45oI
Qdou5TRh3h5xR/ePOChg+JLNJ5jo9C0AfZdU4qMHyai1hXaljAnaOLods/pCXHG3
VIf2EQh3dNTy7oV6kh90I5CccfE/lSYt49TVbpDmdQSFrsR54p8FoHy3li3KgiL+
YasQxNQxcGt8SjupP7lkUFoFclVd1ER+Ds/HyEmEL7GyOLKporJPWBcj4yB1vjMT
eSqe0Nq743qqSMXmoryzUkfRaMxc4NDxlXFnI8iA/pla9lYJCE9Avttfo5rTV1aR
AcP+IMIunnDXU+pFDeJcxjuILSP5M3NupaRVTjaBnkoclCR3lHVWOzNTCsPCFZVF
RTPO/czcEFlNnjD8SUew6RME8IAqZY6Rmrz+TDtASe1WZ6+LAAYDHyAo3bb7dHls
9i4fuUG51sGK4XpSvS8RVkzCRaoLX7xRaTeCSN5EGlVx0bIdWT+3R33M56j6ZD5h
3a9/J1g2003Qev+AoaT8E2Jj92WOyeMpjw3wzPC8VFUzQ/bBZpfj9Y7eZkL9gOAf
3RWvq8kUvpIBAwUN+QCNI7p8WQQ1FZrwiKHfY6eNQqKl+xj/6gT26rDAOm50BENo
NXzZGolhaHW16gWbM4kkFuyrVOhPMFYeasImYArxz6h8QWG2MbWD6DHbu/SbLGMr
ZnR2lTC9a16t6SyaDWMQirgcXjAEMdaEi0fQuC13MMBWOakb8tk8Zf2ni+2jK35L
EAKHzz+DDQkVH3Ur6vVsshoynRN2rAJWODztZIDqpRiv/0/vOwPjszcqhvUtm2yb
grGSSDSCyyshWWMpEcO6gZOVByc9HHlSfiVw+rk5bMl/i+pMRBgntrjr7MfzeVGB
++AMMT907fOIlVhM7dK9JfTu++IEG0XFOXqPuoDuH7bwQzxEa9GqYrah19qEaGeV
TticUzObZcjt/FwWoKqZvJOkF6rV269Yx7O2jC9qct+a1YQOfMAd13lwSgsNqIZM
2LqL0NKsC3LarWOAxEEN0Ekf5W0cA0Q5APqr2Iv7AVdAzl/ykdodup2NnZzw76lK
pLbFu6ghW49zk3iRK7pDpEn0CnLSVa1fc1dfChrJcy1FgaIev5wW7NcLKW9jPtPS
QOAYBI1egh85TuZPp2vtrdCKd9S7/X8/Ksql8YyOh1TkvscqdhMxwPfc8H2IPqQU
G0PBfJOi/HSVof+UBISekzPOxS3orvK0YQ6MltqrGF+jr/9XRS/cQvw+/asUOZtl
8hk9WQh0nJaEFbbGUkGK0rt1if8ANXBc5lu1nR9gO8U/fxhIhb1rRn7R39u8uNu8
10v2NvBSebdPaVvPhBr5XIRxGOtie1b0KVXFSLhC+FP6w0sBJ+TBsEZ0fjb0Zd8n
CyHbPJJVc1lC5R8GuJec+hpvwsQ/vLnvWiTThGVbhWLt2OMlpra5vrIfVVA0Ms1s
JxunrBKDJNn6184UHiNQBEHCB4cxsB5bJYiDWtiJRVezelL/7++wx7nbWPSmbdnS
b/aJHdmoeNF2uSrXvPjlZRx7f4Z2Gr7eIw6TaPXA+fzG2AlhyK2q1IiBmehSO/8c
oVmFNVONlvMeAUBlhaNPTbNpGN+4td8lsiP9a5CD5e3Aei8jdnuICuIKdHVrVjFg
2I7o0aQHB0dMYHk+l6QrCfXQv1DQPJUhv7/7rg0IEMHQ0wxcHUG1IZgyxQiMJ4kh
nrqUN6JNG8i3jHnJlolV0Ad/JdyOp5gUT3ofXxzo+97hwUPSaAc41Vs+e1WH5UVY
uH+0JHa8qeaXCrRY60p4bvFqGjSrFy+VIuvpXojAG2Y5ors3Z+KxYCmUWiRqKUP2
V/wjAqNQrovwgg9Kslde25OMyDKKx2J+p+h+gZ3G4iAbr7BP/ILzSF5o9zRM529P
vEMafMFqE2zTQxbKldxLkwfxxaslWSB6KyCG+0NZ1srRDnfF63pCWv0CCxRdICwc
I9WHAR0jzpBhwLUsOUMdY4LPl+6heGs8IUYRSdxhTEVzv7+tTe/hEXJ6TGdoZRcW
SqPEnYPF1v2SuGN/YEMaDFqj3yUQ/c9ab7xqoTbqgbvXcudvGB36gste3EM99Jbb
9K7e2L2Lik2gQ0M5jlIw2z6h3/DUDSYKnv3afenP9OZtBKhu1IbsZoOnbJYivciC
l3UGQ2bHFKKT039c24Sltednnl5ErN7RYyXIcLULMdU+koPYIRfizUPsRhU6B5Nu
R50BVkg9yxe5UcORISzjnlVMW1elZgiP2i3t8PsmBssY6+zEbFuU0GtQM+ipJXkB
g1ptrevH6O7cTNgcLXsdzgTFPykGdi+gSxWNOPMdcgq4sS1Nkepo/87QvS1sevcB
gV+G9MnBol8dmAAMp4OVwTJX6xXPITeOuwTlaiGbVw9hbs2Sg/ojHGrzsMq+eVaA
0KvrLANo4pvyBsrSq3vmfa07SSjCVra/msPzGp1GLYuix2MeIUVT4CPDaYxEAxys
13V5DJ2rKfhPYjNn5iWO7l3VI/KL5KAs+PtCLXj1XHkO/GW1BzxgVjPTm1xwjf8d
rYFHYmXJYMCdjOMjBDsyomUiQPsgXKG/OsbWCoJCj5Wwndi8EAZJ8ZstGf9EhFyy
3hqmpFlj/e9xVaADs5anfWMTAHsed00vUV8nJg8dZEM8Hs8BIqbtLTLOnRqlWHsV
AftxHWaA1FDVZ9N6pAe1ZwgyjfJDZDYSpvI0TUZ4JDc9Kq8nTs6W7HnzQu0H4feo
kkTx7zTsAjmlTmpW+KxeiUZkD+QhgFwsL6qI2ruFfkOTUuK3fLX8cUH6PP6wYJpc
hxcNIjoXG3EkIITKFfgElFOIEiKg24BFwUiWd8KZFkFbm0LmZtFYyfCYCcGoPZf6
j/CHxDNKyC1o758xBOaDfUnOIoMlrT4sRckDR64EbRknc+/hzcsAJQ8wNxU6diup
/DYCS6oEDwUyWPYq6sol7OQGC8bpKOpJdo3gonWbOQ8WtTDollIjh77XzzSBajsg
528c7rqOdOGOg1Rthe+O5HFCBjozMQ65kn8WX6zVa3F5tXxqmwpUQ/seMh1hUh7x
wcUgrEkbLCd27FEzrNeGYzn2GvoG/2tUiKilxVv6ey4eM795Y5R6EsRq3g7rUvRN
RAM5zddhtu7uODjB2++xLhIur3WFrTRM/+/PS5usiCQIwBErXB+fos/lmjx7yFv0
2VMwiu6SJaJBnpy7dq7nEZIajwuaWKpO2Og0ZnvROL4XT50HDW0EwdbgLikCDNZ+
b6QQ3aYnKsS1I/yRpqBNoAAdS6BP46w6A0d4SR7vwFJ/N5MSvfzAbONwcLCv6vtx
TR9QC0MbVPsNiF29sQymCp97KdvZDwULBsRd6qvAcYBfhsZJBAX7dnQVpjmWQIMe
hJXqTMuOpJLa4SQgg7YwlxpKPNdObgTeXfGUGorBOGoTztE9VQTb/SRwApiIuxVY
5xcNQV384Qelk+lKbOB4We+FTrSPWgCOgyBBCuzsri1njZfY2G5UYWq83Y3gwRBn
GA18WB8V7JwsLb/PsXLU4/CjzYv8wZzJBVivrC1gYBWrrmB9vdxFEk+av8Jl/+/O
Ga8fOLPcwN6QOKpovjZuSFZOKLe5rFnn7evNUw5NVkd+e0xuQXJ1PU0mWg3fh31X
Aq/EJIsry2lDnOVloV4RkJDHZ2aLqDqJ97k3ljQpvQcOZk3OzSTjs5KOwfX33xQm
LECuOLlgX1hSXiMWYWRZadTCSCoZBIn0KHY77FgWIW+wxxrmRU/pAszZU3wEq9bo
wRT98hVMqMfqHnu+z78Bo5wVNYxYI9fEG8e5sarHtHcLa5dboTHfD1YdOldVfqie
so8F1GKNsejpmSDY7kgGrFowPylZNQMURLhucSNN5eTJhVzSGbB/1p5/VTfRijYb
ty5WjioSZbZv0l131nPkMeeD9JwvPyr7+NPufGGpWoQdA2T8aIk43i28PAMkixTJ
QqQAlK5fShzjGgOvrEvrwqV7Tpb1m6zwAMTdhdEUbZJyHlPJa6vOOxQOmcW88yxP
DBbN1PtEBZ8m85Wyn9vXxlBBAlyCooeaUT8gy+yo9hK/EBXR1MYcX4rdIAjxpamC
P1ALKYMAHHz8uBVvmvkgzCkp1pn80R+W1KJ5EqSnrSeRKDosbQrBCTDFffGIo7SR
oK2ni/PWBu2SnrEDv6/3FKBDYC2YVwW5Hxzb4pCKOrCHkpQTVA0EMx6Ffsd/MrVc
A2pj3R5tBbEDypv3wT3cFiIbFvc6Q0IVu+t6z8Vhg/kPMQKN9/khxmP/JnL+d0vi
/sUPZhzAQid5Ch159PXe0pl06wkl/abFqoah9sCfQJkW34NP8SY4Qu3RefwDFhew
baPOqSuL5prB/RbkfErI0S1JYzy9+WwYno0i9JjTQy+W3Z2tNJV445gg4BuMTL4F
zJ34B1Qty76JVJExPJlen1Tm6am1eQzbka+kaFGL+cixfnD7Y7tp2bDT09+MMUWQ
zvdwNLyub62mp+AbMUjtwJT6ADTdWQ1+uAd8ADw/yo8dHTbxSz16FIbZjsBxiOHG
sZ0EVrGDaE5jviWGVyn9JM5uLaa9uzpdznb7Vt4MkNVMcJtpFYbXtuyKuKXrzJgz
EVvmK1+epUV/BnT7eDEN2wlY/hQKzSmqN88g1Or6RT4ayrAlGidkAKfg0rtMF6ay
iY5fGn6fk3dOKmGyV9eBf0p5jJFKg87yUmPSYSPsdA3h3VdmvSRfHaMV2XlWKmz4
8q98AemMd0yYtGFr9bV2PILY7hK+Cfo5oL25yAoiODaH0MMUkxOPgX00ID5sd/Rj
0CsQpuK4luty3qYf9Tq0sgY4jdnDvVEzwoSQ7BGgD2y2vQRXdbN+KjWNin1Xp3Qw
6YkO2qPJrP00jxNeNNUNzulOm+V9BKxawNwCY4IWDyUi/+dVaMjHfWm3Kvsb61Nc
5FBwTcpMj9MVckhx0j2KPvpF5e7yPNt4jYzf8RzjlWaeZjCWtnPGbYnAF5zq0Mv8
k4reE6dWWC4icBz/hEHh+kZriGH305qh+wnj5YsY9RcO7ybaJs/ath6v3xA3OxKK
+Liwv1GamOk8ZtwICzlJSJnwt0hysWTpkDif7kzWoCJKX4+yrDjbQrTw4Hd4Fa/r
OKf9uzIgA3Sm7kKRmCeko/fHEKwD15euxE1DU5GC8Kz3QYSGL75U4giI/iQcHJqH
RM7WQgRPdgBymry082faaHpxcWc2jhNpnW9Igdm4MjAp25BRWIE2EwjqiRUbW0bv
pACpaXE8qvgwEZdhuU427gSVPgS8sfa3l0iXwBmmJzgGWgc35MpitiDtXOgTYX4h
piEaYMMF/fVnZPaNlC3XBQmrq/NeY7AFsK7P4HObP1AtmNtEf7lvxDx1kkJHYquC
orVyKauO0EL98pN2tPOXQXtaqO1Do4TSWNYfEGvVL1xIpc7inHInRrV2s5e7oFrZ
eqxjWZO1byoXbuNseFDaCX9XJxNXC5Mury21vh1VHSMwmybnARZ2I6oVwwNcyYAf
hzXgI/XNxoxkBVSQQq3cQBvqfPNXgMl2htbO0SiGGRpiAUt4nc3Sn/cUc017mX8H
1ie+gfkS71zkPYDWcSgxafEJa7Oyob3qnQCnXREAcyzMlKWDREZv/mNz4XyTaMkz
TprFQ4HpPSLzZTqnfSFe+b45oXMWSzL223RoU2ytQVlqf/ctbAAcos/HeLyWUHD5
BolsBXpoV5TlyOVgo7vZEuQsW0INgIJMjOHifyyg9kYaIGpGdbSnQk79kO7J52W6
vlMZFySyvbQk/10+bLnwcF3phqttavz/YqBCyjh6W9M1T4Iy8tmfuAag60T1Slmz
JFeQv9u9XO8DoYjwgrsZBPHPIbj5FWGvaro0iQk0MK4RLvgaj+oIbUggt3bHKFiu
dvNNwhIZhFRvy7re6R7mmxZbCtOPZCTO6yD82EuN2a1oPRAp46hsBo9/KLOafkmh
9rnJKoyYx6+s6j/oF+5NnXw2eGwIAYYlH6LNUxj0iFVcV0mdgZGudFMGBDw4uIWh
TVIpvhKluoJIspP3grGliLW8XnN8QysQ5l9XR/Lodv8uue4PDh/cvO0JYeBEL+E3
CBGJ7/6F+gh/i/7AHAjOKiUFpyxIOEc8rst2xgQor7SBO6/9OkabEzaajNXnh9hb
/TSHYcRVwm1+C3g/Fkc40466uEb1pSbBCm+v1bxYWFRHahb8GAeCuENQM6R4MjVo
H824XiC0M0T16a6Pe6LIwQpyX/ABrx09zBI/GswB8AIVZLm7zMpf9I3+As5FVbbT
TiRyM3E7IxV4GNs/RuSqSaXvAMYx4qRrCwFJUNrlzITbn5eGFKOBCWUpLyVBM2oc
Svxscip+xgi2nf4/9Ab237wAJVwDDGaIYZFFqP1wKlV9Afa32Vc1TklYband2HpD
3ioDYYFE4wMJO6DUwE99xGrfcgMypEPFsKUEJ3x523Odl1p2W2BJN7C3IoJ3fhkc
UKrTyOdbzXauemanJZnuXkyU47iWkn+TzvPdAdW4qOmWY0W5Y9/WcmNksAgztmOo
/m35gHpeeJE1ZLlq9OmoTOA0rwJ4dtz+3eCH1o6btLuQkNHd+pC6+WNEfTjSqn/x
8orpmI0yRGmZRYuVLWRsOq7b/zg0KyeVNdRizGh2fobGXW73WSqB8iw5pdqX/Gcr
lVhITIaZ27NcMZxzYXMOllpqeVsUnNKq2D7ajULfBY0dOs9WzDz/8EiDmL9IQenm
ncTYuaEVjc1bXemWtGtH72T5spNcYgMUT3Lcyr+K8/2bUoX+f7XewdYL75SGk1sK
iadLzmwrsY0I4TiRJeOXLMnSiL1358XOPrfoTwvVcB9xE7tGfrYyXVuJyresfFTh
IepfQ/IRC2Esf/PhtS7Vp9njudu02ms2vrk+yIQTUNxfB0XcDV9X5wFLZeeuGMOo
NCLJTOtxprQl8ZOmlNiJL447z4eN69L4gv8J5ARKM6FcJTSG+o7L7WfZQxKNscQ4
cfHWiAckY6+Bqjdl3M7ISmrsT7s5tKVz7nQ6nNX7SBKosUA9LRVQLWP3zzNhKPSk
A4Lrc1VH3aaDlWoUTkpxgv9x5lOSgrzSiFuv02F0DuxEShFcQf7kOkFwvChv10QD
Ydoly0rfvs9+N6o6rGa8J+j2MAKMc33jxQl44A9ynIj6w/rwFbe0VcDQs0dTpvYE
G5Mf7x1TEED7OY5BgP6fXeD7mBtdbWZQfSA8yrzUNkuKb9xqHQv8perzoQN7CwR/
eTWqv0+u9pqiJM42M67Y2AN5Y7n23i4vxJWA3dcq2JM5VykDLR+EaqgNworywuap
7+lOcefNsrN4PmqeN3mLEtJvqiAVIp6B2CE1p6MNXw1hu76gZPEg+/LVXXHjptZa
mlBROFI2gAKtr30AdfdLk8vJ3h9hxXTSb8mJZAQpNwFsdJ9UD3qMwzfKm/4KBfzS
OJXLB6TD1TfRCD2yW19dqo6cE0UF0ngGdQ5/4ZcNzW2Ext/UIpyxgcRM9AEjm/cL
VhiusR8EImJLBVJ6Pu9lyHG9kwQSJmU/UIKxX8lHEQgcqHfFahb2FwoChIRSEYCF
KJUbyA3rW/s/OYFbJiIO7Y5f+5SE7cJc15Z6XBhlnOGUXK8Pc0nGYTCVNHGMiuFc
TvWcZjiHl9FZdt7teJD0dB+KwYIz0pyHpHYwjC4DtasdVy18gLArQNkkGxQblz4e
QbjAth5crqNNCpN5FRUSmeP73sK98J5UgAKoDc8vzBPKjo/wHbhH5TFXXaYLIAKg
1coEJoooPanNBSUqPaaYs16d8XSbIs7pO15uoTaKcNQ9jWGyZ0Z3h8mYqmpElvdI
7qfdz3G1P0YYrANtMYYb3yMVRci4roSupMnk5SzXl/0AOnj/yNo6yAtyj/wEYxRk
WF8lIPOHKnnozt/J1aNnpuDh/hv9BfOoTB60VM3unB8rtAWvqeFIENnanfWUJaEC
l5q14+xAFUDT+yCbmC2F79KFU9WRaBvMlcum8DiYNIAob2itTOVtMWVWeVHEaZHF
6t1YSeBzXjgY19pTKvTC9563x00X5I6FA7ICQa8bRkFPRz2TdDfqDnBJR1io6dEM
JVoVJOW2Upwsl2JqNujFVeyIAfFlpRgC0z6VOi4BXSEW4NJKYY25YmvQ/aFIn0ZO
b/uaCF9I8/d+NYBUbck1dXYxzKB9D1HpCWu+zRZVBJcwtM/bkeuoG8LEPwLFiksH
8Y6ggK9I1T1cWRFjzbX7J1C+GD4CA9jBduY4XcbN8gRhek2BKceZP2zCVHyLIUH3
2/sNhHjkgsyT2lCPVfey8Bf1ZrdYo2Dkp+WCZQAD/n/1DVpOdHUt0rqMCJq/Pi5D
5VJsajfCTNa7VjMQC5caJysA/b+4B35aRQEGMKObDkdCPzKctO4r9tHYNjSv2it2
0KUfemC/lCaEaeWS9qG5wW+Mh0Fd9LTdZ/xvTg53dlJVQ5p3i37TTistzoANVzO3
lqvYLb3AELpE5GzhiThYvRBvIDon6/d54iN1rAJG7RU16Qfd9yGA/Y0wsa8sUce1
VszLZhtgAV6BrHDWpLTGZ44XswcrgzypAlMWXjxp532fYCHMeBr+MVnkZSghjfF9
RKrpBFwvA2KzERdzUa7/+A2zgBbWGrlXZFwPI1d53hG5pRAeK+vY0nl+Z4d2snps
H1Qcv4zBnlwmp+wQWMcDOdZ6c8k25l8Cyw0nxgvvYjCArvPAEFvtFrRG3Ybm+MsF
AattKHNRGZjHkjLHOqsJONW0YOOzc5CzPZKUlrcEN2T8eVWVZ7pk1KEx0ht64UM5
PMEh1wrhBmQVGhmBGYmSDPXTu8gdgsGU0mtYnWQ+oIxxDCARCW1q1gf2CtYH+4Mo
ArRTneR1vNGO/qvXcuuBUvvLDucUu6pM/Kyv6DalB+PN73bg2kmrnfRzxlpD08qW
SRJjHzhscfnnuyyYtRbPrWF7ONVKteJEveYovEUVHfy341hTN5M97nuzVjUznhVI
JOdVw4YWSXzOAWh+0eXM3foDCC3NiLrjQD0A47UmipDSFc7jS/OCHmBT6OUkzy3c
EnVnoyuJ/48VgY82KrrBpTFCPUmAiCYsGIYY7fyPg32CLEGT/OlJswIR/Czb9YqQ
ptRiBwwO60zYjNZMJgsBY38Go55DQmhuCZzIXGhXjJAknrRZuSDDLwSMadmizB02
ZL78YJDh50M32V2BSioK+jY19CqCdKCOpB2MMl3wIPAtyEgdmBTSCjF1vLDyRLiJ
97246ls9hJ+tYB84VOMb9xE78Z8HUkqZkqVhtdh0sUNWW+NcwM54eT9RNTq9B6Vc
7PcJiItbZhJH+ih4HM5r7yy4u3Wgv+SndR0jkCpmUg+DjwWdaMbwGcR1zUGgUIBf
kSZNc7m8YmxfE6MziChmAuOaZcDeJDhItecZmoT/uIQmN7AQtqSOtrBBwz7QTt4J
fQ1vsVkNRryjTSmzXtmbtO+Op++csubUfrKJ1zrwOVDunhSjQBgK5kpwjTJKQvM6
BX8ukL9VfZaumkl/A015CSQdl8VE3p/OPyQZU3jOnXbS+GlZ8U/OQV5NKB9uuAeb
i3gdUsNIzxpi+HLMbvZdbfOf0Q757cOG+JROhbvTHFpe0j/SW/2AOK9UMkuQsJgg
jc6b0klVIHAvLMLWMNN9Ep0Jhx4iKFNQAKfp70DeC7BFWskXFw7xMZbbPSLWCbir
6gHeNXp8jatE5cZ9zaCqAXYjYF9JRwWLOk/liXfs2spurUssJE00JIXcwYoIQLzk
FuthiR62J7xeYCLW7TOKz78xNlLqZEtRnjaVLj/ROanWEIG9S8QAKjG2a8uABdxi
dZrGrvZ8fX5xJa8oWzhfioELNZi4ZJjaeXCJAvwlI7PHKGzmkIzEqc7R2J7oj/0V
u5S77Gu+yhBm4EgoJnk82LwRfHZadm/9AP1OswSHzwcsuN/1JrkzAda0n7G+mjNq
1PLSNUKFTqGNFzvQlGObqNrIytK2z+FKB2DWRcGkvX3EppG8t95GRr4YiuOvkPLH
w3BCjU556z4BB9Ymq9YUnvg/SR/ASidHKRHzdf97o++6r2E+3CgkqubNXqtNmuyB
XpL+1c8GgqaPBw9rABX9hVItzxxcNCwQ4voS9XYssZxMky4zBmKgwCm/BfekEKmF
DZppetE6CW6wdLj1mWNA9IvEcOZ6eLVfvYqIvWWLSb87JUWwQpcaaeGPG+XKaVF7
/lt/+0Yy7E/V3KOfi6nfWz5o5ocj3j674i6wBAUTGgqUNwBFSBfOKaIecVHh83Es
PpHL+dfQzXJHWaubAQFM1kSIIN7LOqeDZp6ClaKzAew2Jvtkh/jQekihQLSncXlO
Z16yNyWWgOyc4Ww2D6w2hE15iCavBCPmLh20Yxt+cKH8zW2x2a3CSmfppxYcEAHZ
ffA6apqTwX9ki/ddIkPqjd517pRy9+zqbj1erx4cKXeIdif4UPfCLCpQDXcHC2G8
D1Fu6+lgBfJ05O9Nva1K71R6QmAUXzZQbdkVSGHNZsPiHZeOJi3YR8aoTDbn8pOq
Ta/eTS7Ju3G8nlGEeOVBeIBgVse6Z3yV5AZmhoe520faWbTgs45wIL3jfucRNKAT
AkMLQtlkZDp0PX60geYpES+gP86TZvkATD8Ss666kG4fE9ym0id/4Y8u5l8jfrZq
6bgjocTEJNf4NAu+BgHD6FDf9a5/e7lEMJJylACcKyuHS9/5LQKHvJNQvVhBAt3R
2NWghZhCLmlmzuF7UiIpSONHqazTzVtzlTxecnXXoekWR/zeZXUqrFtdOStC//pI
JKdgyvTo3/ElAV8DrOyn7yaEi7+4yiZElwLVu0IAqXAMlT8xHX9+casAz3cikjND
KMjKD8rHbB18v7BHz87ObF3BDXcXOZG7dnErwmJPgYIlRnaHfs0ubDB7Ao5FD/0/
8fHvQMBrL0E/Mo4hEWymc8ShNnBXkfHJFwU+Yn4MtHQUqEAnjE4Rkt59KZlS5Q5D
K2c95eZeveui2SQL5ATHv8ftglrjTdTEWrCdqeQw1RWcgQDGyUe0tUCm4F+bLAS3
i5n8ZdIV26Ruts0+Dv8qSL4zGQSiKQauuoPwB2lR5sW7HD+TD5WbXehTSuzUFxAa
jNpC/adXysWzuqDWpLP7ePRhy0Zir69Di5SnLwMu7vvQNhq1IsEYFQ03OzBNpk44
eEm9HB46n4CvmsniQ4Dm/g7larqlZvcKG7S92R4Vvzn5p47bQSlaiGH/IiDzaBOT
zjEEw8G5DzKIdCPlF+QY4XnTPHSGRXosXCkiHtsO09jJlHaU5xHFyNuw2zvQmr4n
/BdNY/qEty1QOJnz/I/1AGxE0gAq4U/80fwP3pKhJDLDa2QcXip55a8Wez+A2tzH
LRh55HbyuvNsnomsYTL8E+rVhdAYeUs5f1p1QonMUkSeeZAq3so2IleAhMlDlchS
rfitasHVF+u66uPRRUTtxOuVY+Zu8wi/HNwZ0cavurirZrG6g4oLyxDW82nx+o1Y
EdmouHgEuIz57h3AkMHIDBaw3peIXBQAC71ucvfE0wshMThxxlwEE11s9uuDA6RJ
Lnjcao9oUKibVLQ4QkzAblDPkE683SQTTceDQ66q7B518U1zhpByCJW3k5HQGoLB
RBS57zGelNpzg/aAVHWft6ECSz2Br7jpsZg5LaYcp4CSV02IfFSUYMLOR9kWv2/b
SiA4FSPSdW/DEF8UwKldzOYZpUwY9hBhwo4CcJ9mNHziulcUj7eCjsXIDRzTfEAU
uuY6fjAbxvPnMX9MTbaDTSKwIgt4s6QKrsx0JgvpxeIFfcdz5i7SoDly20d0NABs
qKZdRjszafYXxlFOrl/TgzGOYk6EN7uirFw5wLQn9qHd2QYp+VZ1mcxcgUN+Rk6b
Z7eHmqkeTjyoNuMr/hlJjF5rHKBuz9c9usPWAsaHuzzT+Pc/uoCc/A4ehoc3OfTc
GrGiwQPP5InHuxi+RZ2Q/VxOmUoKwJGpNUbSb+UkH6s8WfHRhRccNNTtHQkk1ft+
/cerY3SOpib5YvH58o5QGvA6ADuDN2X25bSWlW+iEIXqYoENaByeOM+QBKeEAgPs
2DZoKdFBjmP3rCUTa5BdorxDKe9I7+kun6uffdPrGnBHOOCJ8nGjZW/N6mMl5tIz
PE/H8k+RXgZj0syH9oein9fu66Vhc2VLJWTS6lAerbY+QcA846slt4TRWQGVVZOc
DlB39eEPL3XNcKCM7fUk3ODI88ex7E3D4g9XrSsg5C5B2Gxum/dNePRsN3w/YGJw
OeuvyabzXU2DOYjkhNLWTzm+HpD3CLmRFbs1Q7w3fvk4IwZnSKA5OhP0g6/Or4w3
jM1kPrqn3GKByZR1mlkKLoLvaaXLKTD27Qumbiv+SXigkvOGJ4aPW2pPUG0msYoy
TbsOUeKs1oRLmk0QoRe5u7sGmYtqyuXnoUm08xoZ1dgCjH8jFWjnOaIBqy6187GP
PmxVdnIPGtF0nNPsxINA4mzgnoEAubLa1UnnQeu+E5uxDr/8W4pt0hjNokC3RxzS
nEHspGCOXN4gAD4af9AcmA548cFeVTqGRiWL+T0cfjmEInNnVMSi5ShEwqAc90vZ
AwnUzwfqZ2EzTb0fT3caojZzNXzbwlxbYyWEQ8TD1/JSptNRcUJwhDgVLYJ/zgmJ
QNS5HDM/2Kf++Ow0Wh69Nf1y/hlYI6CeWpEHKrvndjH0CBOy6HbhR2Jp/uPCYIOb
ef+XfG5O7H7igMKwKUH67DYraDwGTdhcenHAq8/8O0GUkkWHWBHBKzVmfqBwe/fe
jCrr0dsP3hdfn6x/NRTAx1YIJHQoNaprXWm/NqmMZ2hWF7fMac9YHACkE2FR7dcN
6twELpo0skuPNXZfMbdNEinXov0u33d44jAMU7qUmKwwZ3oCwUJLoR5ZXdXAs23p
e2DL0us2rEzhSCt9yshVqo//T7uBdewoalya160AKS5QhQecAElEVzImCymGT/Zn
UD4nATi5xd5QDZKmgmrJ158/7v47ibGaaezxQYKQLibFusJ1v+mcFSAuYDiDECxY
wny5HGE3lKmrzfdNERCMK4YptU2Rk+zXu9nhRFaigKotmkBGpdzvVjDtDcrl2ieX
inUH1KCll5dSvHa5U1gd9JTP2gM35yyOUFGYm8Llnnto/wgFLJYRgsVURAMNCKEQ
ZNNU+PtFL0RQhhVg0zXqA1lAQneK2+XQNXCFIpdf9fJQncUsYaJEnTp9bEQ9jd2e
w5e0kU1sUqafFGeEcUzKyFD4mxDb7l4ns4b3FXyLHRfD19a5YJWD8vYUftHJQIWF
R5k7V6qjTbN668O58D0lTnnNKtbJTJ7ZxUEH6Ii6bt+VhlyM5Y4kGgSiQCfnIrJ8
I8bgQ/GiwgtVdfvMAm3yWg4zE5XAglNTnAR5TJBwN8hIYS0rkUEGZ86CFTm4XB68
d+EBrw4otJmyDw9iI1HBtM/JyLJN+s+2kNm7DkDG5RTPcRwNxw4syMPBNyyOI9m2
u8BhdUvIiYECKbJwSlMpuKAJa8PYgmCzXmMOI06AwenhCNcay0AQ0Q2VQ2twpiJf
42HJAVv3uNTfzVhWLL1aSDAL1Vxc/pzd2O3k9Cf4FNMhAd3vgBMw6dzxpwjP6mwM
nMh2F17KCOCnDzIoYMYOBQ3P734QlAqqYLwzd46G1CHcHddouj98XrCZA+TNkUAU
N2H6Xt5lPVaj6oJ0CLQWDKgTmIsfdueTLpXH+dRc8WBR6uGKoXTmrw7EUK/oQFV2
STXTbhlneDDi3yXyztahCIewggxVhJUzAmFoIxtglAqiyqfU6CQsr8GzNfiFVfU3
QpIv2YbQP9+F9oh3YAeiVZdE59psSt+jmqk34BkcPHFC9WsgIcVocEdVpMIz1xvq
Xe9k+f5U2ZGVPmsv+qD1xFy2UPstmN/15cA2sstNAAh9mR1QPy7AXyfjFHhhQc05
2Ujt2SHRnOs8oebklQCa4szTM/FkkQ0P7edMV8TJotmhn55oTN9scH6mrFMby4m0
VSAfb6O/DoJQKF0ntajRpC3Az/ifeRNusBxF2HeH5yak1Vlr/7axhgyC56z9t67y
ly9ny4c0WUklrVWJVF+KbL9LRK4fuYORaUJvMp8h3Mu3pj+HwvT9Xfb3oQXSo6Ib
hPKC1TMvHvn94b6rteOBspWro1k9nRzZpMr6NGMMsZ7mdtlaR1TcOpzRapDyIstj
Bm4DnY/aqgfOY+5vphwCvc2Gv2TtNwC8zxFg0+deIqfbLk5J4b+yWWUebA9hXm20
3UMvDPauIcP8kxGFc50WPVf2IE0//zKP+6Jc3K7ZBmVPL9Gg7PWcpYcF44xNLxm5
aQGgtU5Hm5bsG18Iq9eNECF7riwYFmnaSo33GgsTsfj6YI518Z4yqWjw+GxrHLK1
9DxHC3enUkHRWRF996HC6I47/xTFH3WB6zGflA6HtGcUChGsFrnW/nAh9m8+E7kx
i1GHNPL+o8P4wt2bCM0k6QreWBNM42rRwjwDHkfgaKWIsw4jMszajK5+rRNRDcaF
0DWOxveoiFEGDsuQGvAH0PHP6iyLBa8Npp7NwA2fLRN4TDBQcjNu8Xl9D7KEwjHU
DrBJ673Weiz1WyYM1eDR10U5MV3Ojxo+jL43YVEiHdzNGA4KcMafryymBmohUcMl
mioQikR1odjQiyG3YlqAkvn7I0PNz+3nwgWMb1EApdU3/qFKzXpmdOD7zOc+CLNd
alfwez0SStOdEwn083kv2wcNfs2Gf1jvPCwmxtIt9Tzg8fyCj1UiJjALV/ZilIUw
BfeJ3ywXji0DnN90WEBmcIBWn386eIa0OmaqeTwqR2B0kqysNJGpt2v2rd8VIP/C
CXToox0ESu8bEIs7MKcnviovXJjjJn38OmpzNVXom76c7x6JHBowMrqU6NN3Zw3U
Q4rpUU4BLPbUrpjGJVZFzoHSqz//AJIH2DBf6wupGRnCzb2P1yoZ7XbQGykpVqSv
Pgr9aQ05VD+UfQYBQPUfWQz6jBmHUaPbqJdGJG05Ctsqomms/jjqXfxaBYkG2tyX
PpU3rI7G5EAFoIHTdQ+S3zrmXGUBeTfZbWVbNzbQEkovV6QHHK2Nx7GnI28uZiwQ
D6V0DKJb9KpHChj8J4oc2PlH2jqkCcyEGSvPc4z0ODpXGklIKro2jNsBRUOuMZqX
vuycAiPRz8TXl4dTiw4EMRYyTO2X54MiXdj/qL+7T6isZRU9f/7KxaHgxMEm9J5J
qeJ56k77/CrpI0/4AGRwY20WOreGWFmgQWCC54EjfOq6ASQALOjuwTZaSycUpVB+
Qc/T/ZRKFOWAd3GdPpHQ26KmcTTEXcUSylGVGtI5cDFu5Ve7uBvFZH13WilapOfw
au1vTdj44QgtxHjXxb2r8Q6O6gm+hw5WPGomSsCrQK3+L91NDr4ZcAau+xGWAIzt
acGiV/cXa43m8UnvxsubQT8bRuD6gGTRzzU7SaCj4BpKCVSHaiqhjjFlvRfkr9y7
I3CrrKuB16sboDZ+pumaaySh4uYjhVPRyQckad9Wp1ZINYCfq5vdh7tKVr3LrjvG
pe5uLuHL3+pwfU1Pu+cmGwIef/TdDCP8Tzr97Bu4AMk5SZEBcctFGsvFZevOYkWL
tRzbRl5MFl40EzFMxwFIEue+BIPv1KrzBJVAl16l+CEGomMLrdz7NIYhauNqYdZ4
tn0CgFf/UHE1jCMVglUR5f+GucdbTrjtOPVelKkK/0NdFpCJmUgfvx7Kyf77dI/f
BZJQ0kQDV5Tt/wx6ZAF4ViOll1vF6+WTuSQguyFOKQoTtbHKPAse1Gp17OPMj3s1
3ICjosSa8b52T47Gd/4CXmPcPCfaQQYBksuTRXQr7lOTs6qqnbyvShB4p/JGtgMv
FPZlweRIi/ZtFuGFjyLtux+nnLqAOooatbZxgtj7i5plfEu7Z+HaxuWqSJG+DvJ3
F0V67VUM9w2+kkP+mHxfdfy+PdWoJ+lQNOe1Vk0qlgRVWYotA1jb0onFhaLtXYYR
JxOemSnG9ktJRZtSzjzbox4hqijISaFMVuGXjWPd8ZP3qQfyY+EwvL8uj2S8IdHq
VUPTrrgLAlzCcOU4FKUthRKTt2x+xsfc3BG0acwBNmziaSN+ovPRk1mG7KDA87g3
ZvLTaq2anK92u27LhcHoHV0nHmA5m8zJ4wADdJKrSiYCOeYchfguS67Gt7iapZU4
0y8RporVgbhi8AqeO8Pywq6TCkGAqRfXpVBPY6ZAOO9uj/mhwIbHFtTwEYAiA/ln
7tXJ650vRYUbYBC/DxSWGUNFjOlxRMvjjKz+A27ZjQjqr9DQctA/Mk1tZWt9DOIo
Ky4J+A0IZr/Y4iyEiuXf9Ol71AglBY2HKlYnorXlpKZAGbDnP7EENyxPlniaN6D5
haJZa70qe9IYWfiYGBkFPkNLtORiSaogXZYMTrbFde0pzV+0Q8wHyPc1IPMRa3br
oYfnVip54wabdoPfSezKFNw9wEPwZRT3Exwykj+Nsxh5lDpAwu/IeHsyP3YJczVX
YXvR1GfR4OhRTwN/MQPQip/G5CTSadvfHotp+UtmCpNbVsB2EZnEjiOGfTJrqfjq
GF+g0bQ+0lNJ4OTH5Uc+hv66IqwPhZ0DUZx04mHRVNNk4WxQmqu2/R5wG9AqOwXP
xB62I2HZA5XZ/VmXHbIsa+PyjIvXbiO6LDvq90tKwJQmmom12jPhUyU9jbNSsjuZ
/kwDEkwgf25RP7wjzk3+T/vlf09SvA6R/2tjoWc9Wv8sgOFnaKCK44DO3PBqlh3w
PB/3YPQiKguo6OG75YHL/7fPkLv21EP13/qG+6ae3Ws91SQSTL9EbxrURX8ztuUU
FRL4dbGkMBJU+NF3YgnB+Adn+t4lC/sye6+3VA0S3eoI/trlugR0y4N69qYoGK4O
dnHmo6md+LnYrFidln8x0gFgY+fFfcQoUqnh4WpOP7kjDuHpTT4SNx+3/C54buFO
bWDDg2gY8oqpMZ/5ZVz69TFZI9c72ryYB3uhf2eYsdW3S8DsKuv60Q8qwuuDjnCX
lvjSPxbdh5PKZG/RKA57Wg/C4LXTTMjdxOBq21fm/fC9ev4VISyb7w/pjK8HVtGM
JcTbqY/xMwwbEzQHa/eFyYd0vy+LoadxlAhEnZY/wwrTua8EuKovLGVFVa/Y3BTx
p1uddvqXbHvGawXbL9yhREjlmtIP2ge3MvvfyusyFmPhY33OfQACEyRjFispoAx1
hYUMw9QNjTbXx2BeYbLqU3OHNgrwcNl4DvE71yZY2Zw+3ebZnmIv43NwrUqfU1Sj
qeSFlsgwZ4BHH9VOkckFJHHrQ6BwVUsi4VXtvIR1+BIKrnPYWLDu3SWLOX+sd/0c
1z37SmAg7l1xxN93jsD9ya3C1vh/pNsFWtp4nQtnGH9c5NE/GLPCQiU1zjTojzev
ZmYEMwgF0t9u/8sI2VwBqrIXv0ZqagKt2EEHVPdES92otryaidcbnefZUcaQFy45
Okz4qEFv07u9Wu//EePu9qOQZnj1a8leCtyzXiocPefX3f2OyNVr/i/87sI7B7y6
cnrFktKXa3ZD0uNcZ8aP9nEaucMWsuHc1rDhft8UqndsbnLE2W4GoenEtztnWyQh
xPs66//1d0I9Spz5fRHx3y+iasapL0h5BulvbRZOrXMoWzomcBwJRGspyjG4JJiT
g8YT3xw+hbUAj7imv0dlnGVp3hwZPn29lM77Pgbucuo8Rlx5spdQdTG00MH7pswB
idkAssZswO9MkGYC/KHv15pWrfHcXLpZ/jF49c3xCRsphbRd0FvV4MjUxXQIZbj8
XhFavimFsdgDD834LFuDN6AbP9R/2A8cE2AkJIEv7AESTGIB+4bVySUiEroCxhhb
NEQsgapadL45eZSdZCB2998d+WGbgk3uyuKnEYFMfUyt1qgshtJTqzvmiy0eR3e3
v7zAmCgw0VaSP/9+4ie+DQlog58CvjhfvZ+OeGciwKvhPv0gfnkFkLJ8CFd+dxUV
z1A6OkIlTO1hwcU14Fa5Zdz/l2Wl6nzIn4Q5+mBBW5F+Av38ONR7ofRd85KgLln3
sBlmAQMAzhdQuzSAOYUp+yQWgk7q+va7bQ4IQXvsuMBY8ZztInKRmCUahw2ARrWn
17gP4nONN1CPSCMfZoJOlKHrNVwWXtUO+Sjufy8hqmHmWxd8gJP78Y/IvVbX0WMW
s6W1LkLFLVaZ/Y+kT9hYRqN2qXmXl57fTDsxCQK800efOUQXvUf8LwEJwl94RFZK
g7N2Cv91P0F/+vDbJNEeKN4Z778iAa/PBtJaxq6RoHqGHJbryFbkwdoTKY6Ue1k1
Ti75DgHt0cSIWfH1o5hv7PQz5N6leUx6VOpPcnrJeKHni09+GKdIES/IY5POr/Ul
Qkj4/+P1ZUZjF3TV8fAb+nJiwyff4NKXK4ZHgPwYYeLJCCgbetSDL3wfwc9f2w9O
k49X3AYfLn4tOV/Hb8H1kSqFkJVyAClyNxrLkWuSFqTpEPDJdOxaKw252H+/gn9E
lVbbrchrVdz+Ii+NoDSHjmaYhR+EXkqATlvtZQ6nsg5GOh1n/cPecNjwYXBDhS2Q
BPG4tWSnzIEZaCihixsU+roH/BXykrwYMx0+70YPb1DLs5vaNdXYYYSEFfrFvk//
7L06ZK6P5XtX5GCv17ZMacXsAw0HFKBtNhazK9MAD2rDobbCSdtAFlKUpDe2DcxZ
6yCIxWFSDaySriUJFtpUboYJhS4MDQg2g0L8crdMMhXpyUqYpIv0ZVYeaaI3pHlK
Lfjv7J9wMcJm0I0tYeDyN7x98ibE54NzlaBpc4fbnYXJXbUCm2H2fBUtaTwx/cM3
9KzNWTaokLhkZ1dpAUqyuJNnNelk3//e1DIi+hB88J9jUu42UZkxS1RnW9uMvIh6
oQ95F0cVTl/5k7mAfibpSz8ig6K81n35COFpmgEehexrgofCwVh/DSXapJKph8X2
09fL64o0sxsqUDY/tE+epGkj6RAW6uxTBA7JFGTrI0NRbhAjLm9PgsIHMz1ceaRI
ewtRBKjflURpVVsrW4yR3w5R6mILNxybxUpaNPRacCg6nRpkJJILjbZpSS0FMeX4
YSv1Bpuna3uo05K+H1MiAO4axCGyCp1Ns9JkI7aaBcERg5adZLb/UEs8/hTCNP91
CB+MgAJ+l5PFa33+dRsUQxvotG38TS4rFqFG8enDYeylXP6KdVdZyty+oDK/GuHy
apuRFGAPklDcj6XBFRB5ONwjnLsz/OH5cMm68oCHXnG4/d6gvihw9ABuK0x3nccu
JcmGLA0vTAbryXLiIMw30TKM4NRpaKa1kmlMD7+CwfDoIKn211J+2bUyjiH8KNus
FFHrMaPGvBud/nj7eOzBtaVorOrd156Qs0YYfSVrXKEi9RU/8NZQVFXroaw544hT
F2cDX+E9B3UDWAHZ+lSpeyx+2Die/Vo/O50RgJ5mPu85mLsWdGs8xomGZEzQ20x9
1pdBU/1pORkLvAXrnsP9ELU513KhqCMg16lTK/sht0tYB8yWX0/KYAnHLPVFADzb
9A9wFiAuI6Fro73qvfqSUz23LLW6xSy6hZtMLh79yq8cCKwzN1wjVzltm5ynVjua
UBca7J+PhQ5TqP+YNYX9lLTeXssXtg+a9nDtA6X/r3JJ6/QwZiRPIstK/DgSDN2N
oyJEmPeltP1+BPkOqpPUEDAXtYTSGyvHGSN0NsZ/itHCSSdXhNuWs/KY9NkkbliF
qAs8e/WTrr1PhTPaCPZsr7u1jSmn6Lp17hiJCwvy24nevvJUthDZqZWnjL8wZN8L
cJyxjHo1oLQDsliwL86296Je7/x56bbTT/nrz4Q6VO4BXSZmx96S0cNDVtolKWXy
G0m/gq4UT9auBDigfyiwUh45ZufmsnjbfhTpru9ysiVerPvk1BSzLldyCGJDKm01
CGLyzrwxz80XjZscNxoACWwfHKX0Y9Gl9lJhJCcwI1rxeMpNR/azeUqwUivUGoai
yxsUsyZLYs/8gtxHHFO7UOCOHPVtfiMcSO77ltxtn98+txd/qoK3qYBLWQ0E74C+
hAajx48l5zLhuKwPI1iDZq5u3+yzYnYnU1t7FuC5jZvelx/vZCk/k7RMtEJ/IzKA
ynNgaELIHQxiRUr70+HCzAn7ILYNiGgOO5fKofVhRjyZOkQIVyP0WVyDXBDx+D1+
iNJqAEEd+VWCfEilFmgJ8ZKkrFgNS+7U3xAqRb8S3jUMM5kIg0qH0LHNC3zhuXq7
5d9RIjCuG47djnGxNLv2ow+wojbEokVvATOEURHjANd6XOSDi96XvWk36PFgM86y
tzfiU1/29gCgKZsIkG1aKV1XJNgmCWrTpBYB/30XD3xEduHqz9+CsM3IKh1efY/r
Kbdw6tOu86p4TvTsSeCt0sbafs2Jf49aOjPNt0lz0i6XldrbYp7DrXY8Q9f+tkjf
E3yajUDHQ1rt3i8pH3hvO3xrYdSn6YFo8Qc+jvn/Vw983AJNoEK6KDKhaow1B4cm
R1JBqlvJhhOg+CGdm0nGd2x1WKaZtpQuhnYENJF1HyYE3O85XukDUZ2EE/8x5IEz
Vk6nQJ6t2XbX0a/uV/zYoTu1l6i7d7QGAnWC84nJG3i/eKkrS2//gKmWJY5ToyVY
66vR0F00SXKanNKWNt5leXzNKZIWqSDLr+NeLVDCrOhiCVRvqo/II/G2pnm4Q20z
OSm/vMTX3RgoGFHqLmUWk6NWsoQh5HOs8NYk1jXS/hLthXfeO5dkjkfh1hTZfYvf
ikjtIBswkpigxJ5OqWxSOTBymzhPgSX9EQpseJRM2ptagRewQQ4YuY6LnXza+0oX
/mOMmVmoPfscTYXvLO5joy1uTZ5sgq+FqlLGcf/r7z8QzwqcX1Pdj/xjq0rR1EIN
JtByFHnEtkOy/7BLNPx+F1C8TS4bNurX0KuShg78KBN8N4M8yk1vzqvCDu8GF+N9
Nwfh7YcVOvezeIiFXUXGVlPHULKccHCbapx4c6RDnxoytpM/hPGY85dFYNDbnb6N
ed6UkEvLyRLP/RLNRMZUMuRIySEGWY0r7TvSNKA/0j5cgMbepF1WyPVjWxo14RHG
+H3JjwJylw4Wd3xI/Yl4LShGAoDb2pmgi/HAy0LwLYim4ps5o2HZ1hcjegNWCBlv
u/B6VeCCgZJ4SHuQiFOeFT2wILMdHWGkFFYG+OxX3xuIXEk5q8OXokjctEuEN2Rb
oQCta+XtwV3x8Xepq7QEYO9gwGKqYigC7xynW/WJBDianb8v4uZIf7cfHShli0/S
lvfRrOnfVXwvvzeiIAHXyjmKQ2SV9ZZR1UZjw+QKr8nvKKvBVb6lsYgoxkibnBUC
2GDXj6LQpz672bccat6JvB/mE/sgZBiu0wqNBmmbFyoYjtMfk/dvM+L7K1h8ASpO
+qdTfpBTviXz4p1+WghZZBjgRMDoztRqWyjoP0aKIxMjgRLVCEjIAPhC0FjFkTvo
SlS5eAUXEHpqtZQ+36G6JRvwec5B4ttv9JVSsyib/Kb+DViv8KabxkM5YpJEJh9D
NhkEgWzEw028GYHe+a6NYW2Rypi2RfAU7q+ruUGJ7oPXXyiDtxrotq2Z6HoccU3m
4dq3MjNM0y54Y1woba8498AVxuObtgLZRCLAC1q6enpam5L+EMn6i0OacjrRo5T5
zyOWdikTKR5Vezij3LwNUgoYYLqRT3WfeTeygGUXOYnIRzbGL+pxDQUyTBH21Hyr
ks5dPMMBebwZR3l/CiMj9LmTkL1wDqFXIQZvLlK5mDtPsF62JX2AkNnwSu3NAbQQ
H0RL8Vhm7ZEuqyuR+JDEZwNW4kx+A19Khc5OT870cCDF5d1a3FAS+ZC4wA3d1Pjs
EetFGFV1EsKmxiap7DTTT8wdb7gDYfcdPAWqvZ4zdC9melFNoq43Ja+IOpMtemUf
QkaIL3tcrtSj+Ns6QU18h8eNEXVRaGgtrkLGbzoNSlLk7Jow73jLtGx7kSE1iOlU
HpRgkW0NtZUXM5m6wCpQm9v6zFOQVhCY+bIV/+RTdGLM+ZJu5JheNq8f8Ohc+02x
QDGt2du/TjSM90ENwBZFIcaiVZndAoYB15tyXoy72skIJlw/trj1yYWoZ2UhjTf1
UWb7YosluDdwiAuHzPwNTS/VpGRDAhl6/RwG2atDBJBvXgk+QaQZG9Fwm9h5TBRy
BesETlizU7wZQ5r3Zyl5gkT2kbaUjBdSpCZyKwRpYjA+Uga69o6znziQxDtDY11p
dTsmNiw57l6yLp+pFv/IY8CWLYzaRj4uxCs89dmzRqgb9hrAmvS8jG0T0iWf1P+K
5SLQSU4CxUdtriXxuO4SVN+cz7O6J4rbpeKMsUWVJbJlNQ4lnuhzE03NVaf1zoRf
ZqpFGsvf9Sg4aO9+5+jXy+vz2a8xHho/kHbIIGJ+jmstMauyC+J27xcOTQzs6njd
NuGzCWNQY/MlESZIH8sOnHDD3q+vKIhotJDyuAlEyCk9N/vMVzMbhqQ1DxJKSSCl
r8xQkKWmc7EbufAJto+qSG6Iurg0y+0aVw9uLwLaD5fPbeZErN1fc2DC9Pa4ryfr
McWNOLio93cCppF6CbOGF7CB8vIKvtkjs0BkJd5A+2hBF9cHeYN/7Ocrvz5IzPFc
srHJslqfvYYjspRfZQDp+UEnRhmApNM0H3Mn5YPOE+vlOn8Xb45vR5VviZUJzsAj
8zBgq/1/Vsl5Qek5bL0n5yCcP8t8T/f5E4FbCRgc0bnQ2tKgDgL3igAoWIR/3qsk
sS5pkPpA598jSv8KlLoMOcTut5eQ7StCwKuZDsxUC1YgHEy71Lc9OW7MWlF2H46H
q8zgdtXtf3FrLOO/mHLa5R7jcebGcV4IBytziJRt9BU7x3/ITl1m350MkNLte7oG
dRa+0e5p5O0Twvawh0UQNOw7/C8KRDeeYthqZ7xtZRszFc+Q+nLdAQ/dUgJAHC5a
W5f8JUNjvzeYOyLZRgPJaA3WIUwz7Xw1QRG3AtZhsnMgVArgoBZw3pzS/FBVvGWG
X3sD/Os9yvYCJUBZivbAX4YSjL28rmPkP+42m1Qs2ET6j4t0qI+EEJfawd/BADtM
G3XkAy+iU0LC8WLQfDaubTF0zjqLwiZoI8FwnTMKd+oCCdO3cDgEup1in039wPUQ
iFLx1Z37FnpEvpXqLi13hKv/rnCJ46fJNn1XUPEeMp9HPZtsO2LFMuQpBD2EivX5
Hs28K/vfskoep8YVfdZvPqV5+d9bHcbwjmkWf8EUQG2DywepYdxwW2ZXp/gtxykh
VP6F0E+vGZF+68TrVnoelIXHo7AmMCLDZ2YvuN/DrBo+vFcS6GHQOVGEdp/2tVBZ
RO3B8wfoJTImqcN10vUSci6jhA05U1WkwyYAHPC+2tlPVqzEH4XOUG8VNaOCdp6X
tmTdzgIsmHUTi42gf89HOkzBOCr0PUkXMpNNaHm3j9fE9SbUhVhPjd82VMctitPO
wGnS7xS/BIHV/u1wgX49KwVUsIN13zxKxAkoC7VU57oiLxMU7nniW545dkHdaEY5
qW0j+djIOOmm9pZ+PYzXfVAb6aEQ1lTN3T+webt7PLT3BLw9GtvXIcvJdVV+b4PT
cARUqhme+3GyT1iE1HOjf7aLNE0F7fJ/sE6eJVj71+hfFvb0T7mpb22nKM6vb9TB
F1ZZTtcKCynG+XSortAsYIlp5x37FPqinFiPiZill2CZK/2eD/fMaoSkQSbhZ3Yo
h2oZwd508suU7vPBYQr18+9LfFHz7DuWaRxcKsjKsobM1NuDF32mNawIovQdcR5a
UXftdNIN2hQPC5xi7jgKaCHt/B6+XZPFsPu3sDV/3eYnnO76+MlvTwWTfUY2gtD4
fQiz6a5y/TwvUhBP+ozevHOQD0zqDx6EQKh4hjFudUxsN+L5AIJNVq21WMIgR1hx
10hP8pssL2vlhL0ZCohm55fuD2MiX+7nDpuQf/jaxMP0sEPE4z7LRB46THVdYTIJ
HoPfWq4nBV8K6l7aRp2G009coGxoNyP80J8YmSz/LM2BmNy+tn+erBEvv6eFmLXI
piUyeLTNRLlbsycbQxeGeN6L6ii0A2esNUE/BC0OvtrLBDcXaPyqggXmKhoLv07Z
vdcM+VMIVkMnzWSXu1PJHWEaPJyxck1l1fgtly/0Cqm0FCR/gt0+TGEWJsTPlGHQ
i3oeEAfwRc1ZL4NQ0ubNmXsFloPPpwH2NcTjv5vqiXF+9yjKoPHDYbc8mNz/nVir
zUPwfHahycIXBpxW8JynbbBbRroZHkB/Bk5RdwUT4LFKQiEX1hFUQj46Hgi2y0u0
vxsqqs5Y0lZ/idT5n12mS8SIpd1I7HXDVNujStGlbyfCW3cICa1jF/sXHc+Mh8AZ
B83nDbMlzRqfSCBcbRbUdD85RJxVizrE1J62CebkQEAazDcMqwfWHFkoxwcrKJbR
HBHXsH7q+zXAg9nP3RDd4n4PPqB2hWMpNDAMGZIdocq6wnzDiTG/RO8xlIkQVuWL
udE64QYgzl0kgX6/iNEwMWxEQm0GMip7Pzi6QwqkzzRraVt7mYB0fzBM5MZAhGTd
0rjDq70Td0F6CHVxDxRlMbI38myLaOfw8kw+UfMYdSVA2q6C0EVowYVFd+Msw3C3
7Bos8GZ+H0nmf1OtrYIW5omyoMZ9BaUuxotWn1mn3Ts/6bfCvw5x+CWfKyRIvi5O
E1k3yUDNGQidJKYW5bWRNVkBU6HxhPNcC5MYD7qhz+t7HPCy/jKkEviIPJnISMoG
S/WkREqY+3ea7Kj3Rl8LwA12+FQ6MbFQwIN+KtvfQ/H0wbQbRaYPfFTUgzJgggmR
SnXJr1/9TIUvNAkkOyypxAd/iUxiiDZ234rhAwfS5n6SBKFiUYG0HAd9RaSxW2lH
IeQyEpGkFfqfrwE9syIyQUgKnFGp4SXVUUikI+MQUDSYxL+ygVIu1rQavlaQ7IoN
D5b+mZxCJzn8vPJf0uiie3luGfCpIr5quzeggBh1z9QPjuuTaRd5X2QnN4PvmTGP
myTzIs3lCmc7lBDzjVVxLntna/bO7LouqjgIW/tMovZr8SfMrGT8j6UumNkIhBw0
4J1hjWXZRhuPePrLG+ExcWtnUBcwUrkS9FFwaP/8IFo9rUsJSUS6EvI/RkjrgEzr
CuemLo0a7N5oR7jlOx4CVdX9TGAhSCuDyCR8O72fo9ERo1DfHaQ7SO44eEdqgi/Y
fWaZJiBroBJu8F+4mzPOnx5OzwcyBYNnlYZephI7uE3iGNSyb55J2Ei6ffa8CwtF
FPEplhg+qIDGhLSmtiSgVLmbUPJ57MMgS1TX7CaxKahAbZAmIH9uEfXFzIZ6J/Qt
qgr8V8CLjiN7VaI91gVST9qq1HEpWAenS9iL1HEOAq5PDWXlcFGuJ5sgd98EjQo3
XD0I+XaBo9vH8Utr/taW2246DGEuLAkWNmiQPUWHb2Ytrl/HRibN+4T39w9Pkv7b
fV+SSoi4fIcKvKXiUOqCIC4QMtAh+pSvd38prage3X5u2s1Pjb4Zq9rHKKBAZBpQ
9OJNB/+dsJJO8iRqXCYtI1icDAdJIhsbLMcAS98NQONik9tNcGcGR1j+Z9GffO0s
ADOTEW7dVqynJh4hoU39cFRctnedcIDBeahBc0Hl9p2bvoj8xOdKP9eQOveL0i/J
GRvNQpORl3VuaLU383bkBRXdJ628EHSiJqSmniow3mdkbH79J5ygqrWZH5KkRQbk
qGwWfb2BS9pctcj6CEYUcMhxbS3auZ0dLFE0A9YN/4cBBa7dV3AOXVl50AoVQEYT
xYAIjtlTfNRNl5l1lY/XWENe8pS/QRcRxWtCrOOMmlgw4swBf+MlObRe37WR6Kjb
Q9h3MKpzah9C9Gg8wp5dnG9cWrw/Pw28WGl/ufpjWA6yxTcC8UJD2uG8DdPc/pvg
apO0C9Z6jnuMlEO71OrR534IDehBsBbznm90EvD64lAwKZTcT0aVQedSBgISIRF6
L3NWA32dcEHX8mwkeJy5E1KEdTWY7fCIrmlchZpoODgTrfIesjrJ1fz7EKVZA4Pm
jtQbuCQ1xF04Vt8nHUcT1WuBQpwGyab2e5vNVOhLn2BdT4uhlYR77Z58dKtd0Nbh
fm6cCfYb6tHE/XbKp4kS3fHvcWqF9sRWWLme1fQOT+UOIO10rYdjlzQM0Xtue9DO
TsY5u1lb4LIbBpi7l9qTeuayyvrNASYWDGE+49szGzh/b06co5ytkwxvOX32Jb2v
OpNIfc3WTgPo6VuVcvu7tf0SrVnUTY4lSjfLBbSy5lzb8UuVq0sWZFILRYroSjHZ
XCMQtbyjoPksGOysV5tTht4tUTp+OgBNrA9Uvda3Pre0A8zTUrMBrofYFGRzPS1I
2qzky3JMSHj8Psyza2DQi9REM/v8reEnE1r7cdOLXs9KpAc9LQ6xoj7gW0UCZEaw
AcTrGPmubfECClDQxZvCmPfHYs+pQImwUWHfiH27USaLPDnUw1OPF8zc9m510uEE
0067w1IXV6/VKnHNjfX1q/ONavDvuSh14ZACphMVxq5QJYQVGP1iV1W9G8Jq02Br
EADEl46La3E6KyWiUVewR7KYcr27WpYmsBon1zdkxT1fgkwlxS9CD7760k2BLLNk
U2jzkbuYiJO9rNZJCxuA99ZoVIKkeWEygDetMk1E6SNRdVfBnqBKyLoOKjwrUPOl
8OcCeAoTtVMqwHhFFFCB5YmNJ23bo+CkELpRlGKHKnHtGtVkbBzmL78wErbkENSs
kc//eRAaX3v3OekzH9q8L4kO+RwWvRhhWTzrtBZMOSrG9xK9ndH9NDYn+u5DiRaW
fns8m7YXgyVasHruCbhifi3TEjmmqMyOyvW/++/mWBPlaXoQtVjqdZS9Cv6EnZxQ
2gMpvaOPRUx/ApB3Dn2KLiV6JRGETuozl+CkT5+i9AY6F8cfbRja9OVWDrAtNJBu
UUexuFZMywLKAhe/oZAmkFJ+qqAJfxes1OnOqX2E/Jw8bTlkYJNI/7ghbF9E95QX
M1romNWxVLR4xJvWbREUeCvUUPsy72RVywom8JAKt6qn23QUYK6qk3evdML/D/Jh
0ntE7Ocb/Seo3Izu5A6G6zHBldvpDbFBbBJNDtEiuxhEZ+JoEllgqo/PyGG0idds
FSWFG0mwnYcn+Oe1eUiFAx7JeDo0JFSkFIHu9IVjECVp2cnq53zi5jAS8eGiTxOq
Oz3ep9yRquceqTxtVro3IL8yHRNPD+6rDWMqaawWHUb16YicaLFxe/PVqDRISSjQ
IQ/cLI/C1ikgDcEjUDgmmySR5FnQos4W2fAnFohJ5prOXR7M9F91Zypmga/v9QYh
EZf+npSFIwdc31XD0WUBLghI7VK61sH2s6aR3ZeiEchm0s2aUfY52rA6QUlpBZZa
ltvp5o6GsuEPJIgHtZohQQ1WEEAIjU/kJASzIByCQS8C7VHP75Pfqo4YBXjjhS9K
OPEMTXQL8r7WZiWRkZRmycmoB2PaWMt1Sya6qzYLUPON7pxVr+anxzvZe0bXkIHx
haPu+GwLDEpW3vRgRzZH9Htn/LHQ7zvxVcvAh6H4jNa5onkNiVQLnLBcEAKpXVFw
ShZQeWSWt0QnHsLl4y6QuWbcEbS2dgXpU4Yw55e+ovJum/XIhi3Tg/ok/0yrrueX
MDkuRINKtoHVOenQWJAL/sDQXJDVEn3V/RL5DsNB+JhsAuspcLO4UCURurf6SZdq
4oGIlItvsvmzcRai/CxbiIXB/YOtWpu+9/obUSafX0QQ90WYhLPXVkj52vnwsooj
W8LSV9aOgJ4AUMr3sm15rm1+CsiYTBM+DuPGCmQq8KPDG9/o6zDklQoplF6MNN5j
AB0FuFQMYhuRfhsuG+xYBYPVBMseb+BxPcStF7wcQIjWGGN2d8p0sUiRwla5cdzt
90eWtSosqBTnl9xcmj5xz6ZvcwVPoYtgsai9CWCMSoEBtrFMItRmUjCj+3P4+mkZ
BcguXEj03yxQEIE6kJwhrSJP1jt25IZYTQVMEelA9E28a9IKEjtj2kWibfNnmfM0
xPfgQ7N0N8/ssnlhLA40md51WTEmz40FMm993oEHICI7Md/bxZPgI+KxlAYA2hqz
i8m3zmZk562yn/rKbxgtxF9F4VENGaNOyoaBEwm/5r8ZajOvg69dQ7l0ARJlrRQY
zjODOHzeHDZ/KCRbFs27jZwnsGxV1TxppAZpc6gRoe+arTi0PFO2c4DE/P0wCk2m
wmwEE7UbRhXrqeOIzmqEdeDzeR9fcGGH5vt/s83BwOzZv8IJwbSNUf+Crma+lvVT
3lw5xdmwHcE5ja7tm9NK6htDyO7gEPblGKI6zj47FsszzzrumdBGZsRlH98LBf3g
lwaecToeKDNaZdd/rh/7cedt3m0muyCY+J3CR7uW+f06HyYdsmqHO/V30MTZewi3
U/lXlBdWIVQ1mIITUnVP7AZ2A0L7WybBkJDLzTAIHdcSZSKtiR9vTdfmcQ4ucj0T
GeTBJvgVVc48Woc9lcut3AN/J5qXB2sAia9cSwza805hHNc5ucP8COqb/XRGUdT6
SVBBikdoughhZnT44ynA/Cy1dwdmDhd/LDcPWvwF89K9OO8axI3Nt/M263+IVtWv
mQfx3aKyf32yJBVMvvgn0X5S6SquUmGw7OE+XfZd6GXeWWWQm5detC1hU8zlDscF
B+tWdobKnBwxGVaD6cWgD+p1Kzhyi/vZ7Dt/ubS8m2+zYfUYy6OegN6SQCLlxAP2
Nmykx1INHIUFUFp+XRFJ3LjqQPMjRfSNCoo3mSqTXaq5sEOrTRRXEjooVxEwxNHr
hhJdDwnVmNqzvpueIwzPylmUpTxuGnaIgk2eHnJfBAtLh79CWbYTv4QA6Tkj+VoX
AaaqVZLz0Qa8zQ/hIuwkGNKQ8quA90kXIZF2gBTzyQVBQlG2V1iFk4VvDxX7EksS
Ycw9Aicd3/Ef6RIbagTsuQ4TCKywxNYzHE/6ikkQRzUhkTj1ncsj2TC3BhJToZ6z
muhpw6/YAg3efl0ijf8tBKpxEjs/sOZ5w5LZxlrMwlcXi9/ZwfOF4AzEMIVEik/B
sTEoDsTxoPiTQHwDidq5MwEVMunfd83kteNjYsea/4tVSs3bEavfrVkgSv6qHW4d
1x39h6f8n/PjfvAlxGacRWJDpn/OLcDy1tzFAHf+ix6BDBGHJyJ0uRcubxdQI8Lc
jpk2JadLtxLb7so8Hx9F67AMSyDRE+uIiQtSzgl2+Rks4TpKqfesQcw0NN/w5cY8
sz1d7I1woxYUBND4S3DG8GhuWaCfPhx9eWxnnqddoE/UfWdvbt5Dmpi/AfLjZ0Z9
zff1iFEQT1I+wIUoF3wZ2ACGkg8CctVT3JhS8gbV/rNT9smyx9uXmvfmSYLhpOBl
xVLS/g7bDXZIKBb3NZ5YUIqjAqQqThL4vjfv65ynwPm3jFsSq1yF3VdlwFUNpACt
PUez8Eoe66ZfCkb7kmlg21GiTFhN9s7Db0pyhjtrIA5yvs6lZbNM0GBKJCvnMOjP
F3kbmjTupwoSBjlfaKh8+5/8TqyELkOv/jtKgipKTjwi4Ma6HKzYBx5IqOP2ALoW
1zlmEvsGOQfIyZd1icA2kQp9seoawaVryw4NGpvqo3aBTHgx4aHWleD+TATrW8yl
Ar0oOWKokQ8rkbg8U13O+nfX/FZUySrMrYcCKbC8AXaD9DbcJ+YM2d+Flvs5QNMr
7L0JOzM8GApDcSWgxY+1VlMs4aOBpOQIUySQfqIrVuyQldHGV4WqeS+J1ZBHrTOn
K2WQoJUxH/zlbWoAqsI1FG3Rse4k6Vt7I/ucKZX/U8gTerhPjfqh6IfoJCPvSyJS
yyW7t9BmghgYKGE61EU8wn9a5fkjL2MKvB+4x/BcYA2KtsGxz9td41A28d0Lg4vW
D1HswYEwwCKyF/xTGG9SOpndvZaVnVTCrkTCj05sycdN2yPfzot+v5RisphUarZj
MxMz7ue1Tb80sGS2zuY7VKgJZf+qaCVS/IyJvtd321g/xaXA/eY8FTTSwy9UcvFm
lJMTzMk5JD8SS+3Ma9W4tJLChor+jLl/+U+AqEfpqJJFeKahbhOh8AfOwmCiB4Ue
m58wEUwMaR0NTK5owbzGwZS29VLcAiQfrQqkYCPQTxDyOoSOmtPWCfUQJ35h1qW5
8W6nsf/rl8/m/iNutNCUBDTHTvsXXgNCXTgbFBUzYjhoQYciv8Vk7b48Sm3kLLjU
cWSwUXtfLHiZ3mDwbK2EDvq9k7uN1vOVd57pdyE/g/W+1x+sCEKbDHnfRJnC2MNh
gtUvq7CzlHuNV6/TOQg+e72CVFO4plP44fWI2ZfupoG79NyLaQqRW3Wn155D64y4
TcrJfpKiDBtGsEZh/DecqFgctKVRo0aUdBnsX+RVWpGh/1r0Cx8Li+2DKBFv5pQE
Zm8Qvpof5PL2NLif/xC4BY4P67N/eNCU+g6FUgRhqXKmer4cwfqBFyC5XjquwmBP
sTPjDoIyo0wBPhNpPF+tjdjXJ7tIIqkHLiTrkgOYxtpzTaez6F30v7RHycTPRRXx
WWSnw95zntXiA7UkFmmdT2jdQYhie6MDBbOmicpAV7Z0dxw6oY0jxIGTQARUuXs2
Et6FgKlhSQqrdghP7mKoCLaLv/dW7JHwYrBIQtiNkAJ4d2MKwP3XuzNzbtVcDh/G
VT6TaGDi7em/p9MS1hCUspEvOZbPln1DKgQo1YsaeHQDnQ02CfNiv7nRHnkIPrVq
boBHUglvkBC6fNmirh0JKpnKvSxGUW4Zgo7HGMfVjTee9gPcWpXoeG0C3JgfHnS+
KbFnkLhvtZJDRQOD2uKEgRVORsCX64rkUTZcf6jj+n1EuQ3cVc+0O3c2EwvFJEtr
fnh3LDz/3ObTYMKOB/2hEJ0AaSg4+f0v6+gxbmb9OrIPmyjjEDhG/WIw8+JS/CSS
BJljfPcbKaCZndpJ9Tzhbh1vWRJ8grDK9Qo0Zuf+Ay1mtIdVnzm39bm534gvGHQl
rhu1n0phv9LD8vwOzwmLbIY3bggPDbrWy2hnQR7fJQeLekYIlE/u2bXvHfiAB8t5
/FjLVTiUnKsTCUV4qlpAsXlu5uqe3VRP9NJIX128jt7mVWmaELPY5OQ+w6DtNtUO
bs7rM8jEUJtDfjfpLH1l7Gmjz38aLluhGBso9NMOKSuqfmsYD48Klm57R5FXx+b8
YHENbJUk30lX3SW2yhMm71F1q9pPkzg6fM4+zKks+Yb4bykn76z0KCGiOtqjzuCW
xFNxd9mqBZ1K9WN16nPbFljFHOkzjSNgWikywQ9C0TLy/wfvRe3M4Me2kWTqkGDO
d0uwx66hspxJxNq2AG5RY6kUCfWFD8S/JIcm9hjYGvvGTC0LV1dL8LQXvWBaTlRk
PlHsmxkFtpjMwhjg7DFs2r33byY3sIlUi3jnZM3gwKBPdBbBP4KQWZ9GPTlqB6Md
PKyaGTpn/ZvsIIiMAhj64BDMgUhYOY5uLPLYJp0m5Gz6zKjRug0wzaHl/z6/lnA9
lQNzJyqZw+XxfHTYVP8hX3gbkf57TDgRiLITr//gf7/NDq4egKe15123j1tjaAmE
9PHrUB7vX1KTPRgJU+Fz69XucQzS6Rr9ct9sWFAJodRW/uTl1Eh0/1Rc82wOOqTY
W31JynQ9Tnyn9HEuHCBjhYonG62MT1PfaH/HgqlHh+4qs2cHm45GZMEwBau6bDYd
TJlk4UOci/qhtRkbBkjXFFvk06QxUNUO0gGHcmGC8kK3oqsUWSh/AigsTI0Jh2bN
PXG+L41EBaAc69xMkQ6cGJceu+hh6bPA6ahuZEp9/lwz0SF4Dm7d4fkj3pEmw/81
1i3DrnWVxq5FDsdATG1SPDCJh7Z6e5F2EdBNQYLSpk2YhcCKzuD3UoX94PhTExVh
ekKjVXMo7FQgej67bzFPdONc8scxxJu7dnRx9PxV9AuyXG9lgnwrG9LdJj9+Tqcx
M7/Qp/h7i9rXAf1+HHo5hcAiMShFaFighe14o7UzaX5VZOTPpXlQPahryelnAMnZ
E6wPhinFmxahAiBAGXb2SAVYA5YoGPGr6emL9WwY/cNWCFOGCQTodGFl1uYMN/hY
k8caUrj3bTlSQPjh3pkhC0OJkg5CmHRMYoj/CXnNL1DunXfRAa7q4hVf+LqoisxH
tcquVOkD3UulihunMOKaxdrksK2+Lr73X1OyGVD9e7KHIyuSEzzfkBYBXeCsWXuw
zkMSL94X8yiJadJ5NigIuq35okdtn2KQ9UKpxkULFFEb8xk0MQREHdlUiI7m4ZAx
ROI72HXHLWPyUZxDvddzrOVw/W5u1SUCgMp6o5vSWXvlTGB97ALY46yJspGirOkw
nK3ceYle/gnosq9KgfISvneYw65ab6U1ehxNVKu7lkpj/q2oUvHa79QKCVF65ML3
wBlku7L9EK24Pm6cwZCO9dh5081QA2lInhRp521wGAq6C5CspZYWQVQ9SZV0XKmq
8d8qFQuBS10BuAlhUWTm+bj7C10SnErOR65OUPuGeBZGuSRxpTTZbBeSk/ZcGeV5
3nw7tM4lQlOVVOQOp0MHluPFu+WwoLyUnvreT/kVfVmWqVwwPSNayVxfSF1zbAYA
wEnLCW3Q7a5FMHc6R9V4Ca/tG3LfnNRchtB+TlqKvmA8+huKBOzzppuLm/Xo9LjR
EKnzGOEXrBRs6ZRRYZZMEZ0gm6XSN3JBhFLen4dJ8CJYivszbazEOt4HsIgRYmSo
nXows3QeV+yp5v6VOR9p5LC2RD1Hyhw8CSvfFQ8c/2OFYXjiJ1VcT9j7U9DMX5mW
46y5wIacPPLyxxiRkPHn8tjkvllZkfnY1xfsqGB4MBWWgc0LtfGsWuvwXiI9jPdl
APYih2tIMetzaLTh+kscrr7f7PjmO4qZYiGZNQ5UgZz6+nm7YyVpOtSqtTZHvYVL
B37BKStu0jTTuoWCZpHZHEr5yQFlvx8LQmRU2JEFA2bIRqClAW/UK64yO8C5CLx4
dQcVko4CE2ajHlFO6+G/9oMznu5oZiVXSN+dFvQqrMDGzT6Zn27OtsB/UlU7V3fy
sWQzud3dkjxua/iW9azqyZYIOQdHOQ+fkL1NLw/4cxDEzbI7MAzpYpCCQNZllGeo
8a2TffN/j+Mz84GfeMcwrp9wV1djC/PGsr2cdSHgKBze6RYYyRC1VZh1wVBhenhV
RUvBLi4mqZrcvFZMPteD9McVqjfE/Mn7G7FMFmsEHVTGikBkYOgJQ5JD+ZVHfRit
yHywBWSZtWWZnchOrgBTXNjvlod983WH/ilnvpVLvlU4Sa+lq4+APiMxdvQPM/gz
rX4lNZCkD79w525zhgOFGgwfhY47ExgwdEmNN4nCHmL1CKyJ0++yxaw0LisblI69
KFVm7l5QoNxXU7CPqCUcpYlU/nFsrfROIDRS9NabW7ZVS3MzG3AN7ZLitu34J1KQ
HYUx8YJlFtdJjxOclDvsCWEiTyrh6IX4rOsmTCO6AmmCHYkS0tYdmb8memnL5ABp
VWaVJPY2k/vA5ODYKNtVBlOVylsFJTajPNFoEYBVxlt0aEbvdlP70ls+zVH+ujrD
7w+xcWxxWZ5CvFvdI4kfq9d0pHbl3GwC4qIIA0ShzSeBwBdD8X1gg1KR5yhaIyAk
NL1cQLqUKw4Ws215cnMcWeyuknMkb4xNcC1QvAUcnD9+2BMDCFRc+rQemfV25ULH
1HiMjAe8EMmeTT1lCv63axOrSnPiIQiyXgiayBMI1uY7TGHJipHcRInDDWu2osLn
rLOTbO8beCgMbqXNLvTE4IO8aU6rxvkMsFlP6i5I7AIby2O3xTTg1ab/o9q+DeUc
YTgkes8v7bouBFzuO3Zqqs3pEtROyquxkaJ8F/phlrBz3aYV5op8VEtwLmlHJOOW
DPRX9cqw26sRSJcDILUHM1ScU5/Lvy7Aa5uTonUrHTk1EIYcB+zq2Dbs+kjZP8pr
EeJcPgo2yKLc8byY4IeSEbO27Sz5ghnQNCmkdVxkDg3DgO4ZclBA6rd1mAfaNjfG
NbTWwPSrjf1CB/37/pjDhKIFY/BDhckWn61Imnh6Ja9ht74QxaVLZbTfwwj61iCp
o4fxKZRDfEIwOC1HLizcIX9orqHXgl/fKsOH0Sf2bTEwxLz3QgLY28TPW2vaYJu6
dMf8Th5CD1ig8A9m5EB+zjJvTxXu5HX3ixuS073AIhwp2QNVjJFBWc101glNvB3X
CUk1mtunDlMGIYnRXFER/fBN9uIZGadTfq4cukqAAIAO8oeBJJeK0DkD8co7d8r/
PWv/c7MU1jQdaQbIaxuQWGzauioQQUfPGjMDtDBYq8gbp6VSU2w2HYWvfk7pZji5
kh7SSVsgmyc1Oqlr5DtH6HN2d64bz1Asqcu/MC55eJC1btWVCmw2obhUr/XjN+bj
Ti+Kptnbip7Ql//79oZPzOAK9xn52I3xchZNRA6ZSWi0vSrEJnmIHKLgFzGW2VUM
fvgeoFGZfc5Xe17O2osYBG3eWbACFDi1GFZy6Lh9oyIv9hRWaOyaTns3ruwCSh30
432RH1VoWnomszjPlWMgKCLw1h4x3eGwP3AhFGBDiXCLysBnb57XwALiBPyZNUDe
1WTX1GaIjnEO9zwDak9cLAMIug0py3ze2mjz6D+3L3FQeqbimgKvRlFuy+C/bOHJ
5UymgRu24CSyYSL1ZqYOdg/ZNmJ4WyDcX+mMjL90I+HHjwJ5Y+gQqoBc85GMTn8b
30v0tDkC8ljlVga4+/dvfs26SuZYpsp9rW3qeai4gSrxldmz6xMIcIWg1WXgKbGP
v0etsNkr6E7Hau77OSYBYFkLGw0SBpelAiS3noFnKDRfdCVicUgwOFoUi+3W2kBo
rUFRIeYy2km8eofnawYZPe4i76ykkxbEMb41z1CHu0ttZxVU2EFVzzHPivIhH4ou
jVMyeHAZw8ZF3Ax6vTC1EMMP/MhXFG9v6682f70OINSLszfWYTe+mbju4i0a5SJv
vUxO0QpRDJzGQejI1Des8HVYJfM2QkcjYBEoKjiXdfkjfoVmyK4dvS9jZLXfzh78
yZTgiOaxRck9NV8tLNYa394obwvvcDOMyrwe0ab5JK6qf/0grWLRsi1xdjGI58CL
u13R/toMl0hfPl2DmOxGecbusxvzq3eUsrac8ttuYM+z33QNdJhsF78GQBIEDEKp
icUQAKZIy2WTuCYzXQn66ZLhp6i2PcS/4T7TPFgCOK2uDiHKbc2NiFUYkFwXYSKw
t9DnJIyngBtARUujOHU1YHOIRYG5qKT48r8aPA/ybn0eyIOm54XUq+PXIcb0ENK0
EJIcJyLQaZ6rRYHKW88gNrMDX0UCjrhQIw6dEyYvOfbSW+0IRYlqisdClT35y194
L/Y4ThBoGX6OjmqgpbgtpAODv/6/32XYG9uCXgtnk0ihRQwZgpb1AUTj1QFiqS6p
Tt345dc8X2eT6LjwDUIhsAJPOhYSlETYatFt38SjB12iEvyb2Lk4DGjHglC3HCoH
UWROlbjwPTQ4PmCfSD8smi47ke2vDoss6zpXBxxhjewTlm5Z+BZk1xpUtfpg34lG
C/65rXC8VWv1XeBEkSHbu+uI1HQtlW0DcJj+5dnzQazteyIxIvaJU/1BQ4kRO1vQ
Qj4vEfZSfycup+uxSD+yERmwjjJ2MDgnUZqn4riNmbjKwf2MnsjloOifc8ZlbJ3e
nHW/qj3hp+NmHjgT52x82mGSCJgqPlYY290JcIMhV5xkmJctiIzrAVdHwylMSuof
L7siC4j06ItNEdw/+1RVbNLl2bu2328XvR6JM4HIbBDkRaVZ+7NjHEj38HAYd6nC
BjvdMnB2PMcbeqipM2LJO1arLZrCAc4E1lxpSZY6R+geP8APkHEw5OUEUCs6IYxT
SSNPNuigIkKN2JKLnTxXpcDy2aixtLgkXwTfFZoRv7x/rpPnvqHIgY6hykrRtKiw
2G92gP6pb3ZcSYi/yMguW8XkMtccjN1TDZ5dkw1LVZ1XYBW3JIuBvEec+o9JKUjV
uMcGyuhnjYm172jQd5F5F20pZ3IYmnTsZ0MSc8T6/8E+i1QcZj/46oFdB09Zkt+3
wNipil80MXwWbbkhT4ziyQpYjPuoLQIEL37mBS/2QCgO9ql5nnMr8Wg75gbHfgNO
TbFhye+tGynKUW3FYUMHf8EnFaQFMcvzSQYGaR9sTbn4WqEB5hpxhwHDyJfunAWl
zLFPHNejCFcRxqx8NAbLpOy4lus+u07t+9S/tyu5G5XNkDkAKzrxAT0V/qzKK9ZV
Ao4FjIyD1ERCNbB926+T2W71Gj9SecEPlaP0c5loG3Pnsd8D5UlvZXmR9GyDWkko
JXC1iOiuGzV9j9DBGmFmgjoeme61+KymEg4CbPeTKPXOpxAWmu1SKZ0lt9aKNvms
v7tAWLA6CGgSbAnH+RBsuEFlmCQlXq3w81+piwWtDryx7OytSdUX2t51j8zR0WYI
ED3/Gd732hsYz2YhwU+vfp7+GwCokNaY/LnZy7jYKh36lcvF8EveHwua6zu5mwSF
vH5HMpOm5duDswkIQIcrtKIJ0MAnj1n51Wa8xjI9c9/OzAEkwXlny15TSd0pSiyx
sZdv4zrDa/7bEGS7c6+DJ9UNHUnTsKyHp0lx1IzEWbFsLrVyHiy9RvW5+FkW2sQc
BCogBjWXsMuln0XTArWUKBpTjTalGa6obEJHqRh6/2fPOE15QjWC0UDi3d/BexZy
FSdPfMH0IoX4HzHMFkgpDlJ3LUxp6EcnH1fB/K6rloVuBST6pWnHb3fftemh5nhd
evMN6EvvTV8rkDPppEcKTmSZzSAklJWggRXrYiMGN++wEms1WCURsWZmQx/vWVVX
9hqJ1quN0joyCOWKizB1fsbHBeCGLfkX/3gXjsJUDlbOFfj1gL7cPIPcaFT6qHa3
6Dqo6NDK5jD5riPPQRd1kbSV5mWqwYTjUPsJqFWv3djMx7eJbPa05CAj5EDpQKtp
was4whWsaqghyYiDVCFZADe6kQ/bReeCtv2arXeRxRurBz1ssRN9YZj+dUpQrDNy
B7COzkM/j4evJiUZBVGMxvJdxEJw+KtdczZ98Z+jVMdQ/V9yXIYPvCoKkQxOkd4w
LZH09fY7lV9u0crmQ85WCAJw9c1py7H3bKMFzio23kvTMWYBetMN5SofHFTsDA5A
fAc1ty7peXsN7JO4urnCg1aSpP1TGFZvKjjyt5pmQHpW1fD4Xu/RVqni/k2tLLxR
zFpFODBn8h0Wt12BIyez0Nm4ltw/4Zj1iCc7ZHeJSChH2mqbiP9Fk/CcthXbkzig
HLAZu6Z99gZl2MrCoxmJte+W/6fdd4KwRwNAKqnPpCihwtaAnyf7wg/mSCrCzPE5
NZgiYcPWYvC0GbsS2Vq61akbFryU6TtI5vOhVzLE21XK2yRgIG9YdGvwLkXbBFCF
X7zlY7RFRRbQ4J3hepsMw9qJgQLAqQKRvGgWZVTisoXJdppo91TgOiMfYnKnY+1n
HRowNuGFOsOZpHPL+NrpMQXNdkvdU0/zDq7jS2wh6etWCvt/z2DyJ8gIK8RL+BOP
jFBUUiRLBBo6HtV4icwpRQfmdJe4Wqq8EqwjAA9m59WnKjvVblcL8F/G9GWPZ/sn
rEevbAyA8V7Hcws4IE+kzb+Kwi/mN7t/zCKxdm6QDnxhd1YuejbfH18Os3V2JDd5
0E+dHiP/zmk+kYEy+ybkwYoNSCohadj+m80iGhfCZ5rpdCnDO0YSlUYpM2AOvHeb
PtwTUzDfyD6ZefQuzmMLn2LrYB4HJ4/cw+MbnH1vxBnRyUsE9Vov3TgeaNhyBbqb
UnZu5Jfws7TjYmROubWtbJxIMs5A2Ix9kHTuzxRhadjnzfpUUtZuSDaoH9tEhhcX
2Tgx2E8mAfZHvRM9LCrNx8TWzv3+8wSMCMVyDVaIzBQgTxbVLJSSdj+YdNl4e7tE
vqgQTQqOnG1r8fUrmmuwNc0Pq5+QUCo9CNBrhIRKbr1p3Q9y1K1fgFaWtsrl8Ofy
NyRTusotp9YdnC+3+qjaaHxTOPCgvZAbfTrqAqaS9PILf/8OnrU3qqqe0vbKZwI3
aRhuDgQpxMEQmLyu02oCecfTNZ9c4ejtW4CKx871MOTVpHyTdzEPJ9Dior/WCcGZ
kwslYAAlA1pnXUsiiA0yiMQ54SNs37XLBWSOndUm3ZceZ/u/Lg7CuG+onDQxUuyb
We++TTP852KXCyPeX9TBUwF6UXQCacSu8+7Fw5ak/bga0Q6ePBjg5IqXHNCCAi7Y
ImJlOBA9NC9GemSnFTByp612QUq53g3PRYlrn/l0ssCAqMVPXZqn4ZCuAJLO0oRU
ZOu5PYLeg88nihPcdy0fPxbU1jTAjoPvlY6XUT6g3UIFlHDSwudNLf4yl/OJgAQI
sGosrTRTws3s7JpY15HiB7zwzByOb46WWwS6q1sskob5gnwDs3hq3syR6ZZPN1Ma
GqI0QSnxxJX6JLyg4QC+7pNhKbzbb0OcYxmX8rinDnna/MPvQ19Lc7LrlWQfY3jW
vitGUnWsEwQEc2mjsmyCO7YUWbdiZw8j9W1k1ZgUlH0bjWYLoCa9Oxb9CgMXFQsW
QnDY/WnppvypgHAJ+mFlTJIGApfclwsG0v8xR0emuFAnIoD5Qaq0zq7jkS6/49AC
7Ne8wKz34iJ7WxU/hJHhNCGvTk2/LrUqDKH722hcKNeSyVU4EK+npippMvaJJoht
bDXc6A07bwaTFwLCN4seuFAMBlybMA7jEO9jAtieoC4ijOW7LT6ny+L/BakM/4pj
AVjKsBoYLF4uIOI09wL7EjNfCVvBo6WA7eZA7D0by4QUwFLI1QG/UEnRkxKKdbXH
C9plAegCymD+mqNnj/xiqnko0YlB4OWxkv0vUFzdw+D1L0RLu/sCN++qie/zIlVp
sJBikZ7BURUaaJbeoivzbVzxtS04BV7pj8ymC7doftsF86xupuN40/XpDpxVbx1b
ZfoqQ6L63G+UEFd3n5OvhxnioxReS9ByC78NZVuE3OOAiye8uNFOUCPdgzbYgE3Z
zmfmbB4RMzR+F5ds+ZEV9J6vLGuqSY4oW4Mb3hFy/RC99IiVeeOlHvQVUZC1gVRN
d0tePz4SkiJ1cxJZNOIN7dR0DSsGnbBOJn4nlKf93lF2QX0UAdqT4MLGQ5DWlHdk
4KJ6PSeWBDhVWMEQji3DxUIkJpqemvSaq73gRGHrKHmwLRTWVGcwhs8ZijY0jFNv
zsw7g9mdUqHIREm3+ZdxY1KCYApXSrl8sku0jGDyUYCMhEJTYXQHA9ahwGczkibh
HjZPDLRS4xXACIXAIjEnfr2xkWfXT9k7nhcyJz2HjA3J3R+8/dHeAAL+N8vwjBW4
ztKb5fDG/04YXZBKEs28hUECdO2dowYxVwDkBmU2Jbd546z13klLsAZhgRly1Q24
egIdNpIWa66RXRHcHVGmF/NGgl5b5t6zwJYD/7l/o8zrme+A/FhORTw63afo58Mm
/p5JdaK4DQxnZRaWcZJ7wWftSUWyiHmzkXcGDjG5W7nRJjeaW0Zw9vAAHddy3/Uu
CABQ7HrpWHxS4t6EV67giDLazlhA9rizrtVNhZfv+/NO8DuxhrzsVMXLmpywGj7j
v2iGz7uPYgKBC94oWVqSXgGOlO+AAE0+aKRDsMBUluIm2jM9tggnCOH9HmMrOMUG
9t3u1VcXmlT/uJizhEkylUc1nO2YoOSp/zT9phftljaB9YblAqiQrFEIt3moIaGr
WKrzXoOSzYa1tMRGZAb7fnHD/22dMUe0/i2daZhJ7FOYK/efqGpDzD+2m29nYVTg
9Nr9J8RCEYIlQn8lQX+wYcEj5BXKLHg0+Xp6y/xwS1XatCMIqKhn8s19IPPY2NNS
HxZ89se4GBoXs4G7A7wjMvg6PSW4b7mkHbxWMbGTjjAFZWWMsUelUbQwCGnZ5yNI
8sEzNVftvXVM9qGOIyFNkV9F5tCT3K3PeSHnX2K9XoxindHJHrnhvxXNLsNp70GO
RPJXj5Vpt+uNT3gP3B4LdgvYSfbhFaYtwk6gGSq+L6WB2DpNQ31E+tPQbCIvcjSF
J3EdkHXuId8vvQEYcsvl0jJoYDoXmiBrn+USDv9NPtTx1SdkOOGGRb84Pky/Tmgc
x1gEYV3yiDT7y53zzqx+04+4wlgW55EiyE64rrb9VC9lEV08vrRO+dVVmsFBaHGp
TiblokErQ9LxUWefmAx4zbfaRh+QYmyuJG6Dt4vd+55BVU9iPp1JfUHuhBWaRWS4
9IvgDp2I7h2i6iohDv986SkjExJQjgUCoSdFgIMcDNADGCBbJuyEbyof2vxVg+jT
0S5xci3CrMJiLM+V8wvkaPxBcwA8Qr0fwVNc0bLeXKD9NgjUCInDdXuuzuiSVzhZ
hlE7Mtc3UMjfDHWeykwg1htE34yqQlCYu1EfmSyQrPCG/ubtqqMjxBBLKwAVIET9
r5S34pdeoABKECW495AZ2A3WFx64m2tQyqFZobXe/IrVnZB3X3cbFoIW0E0I466Y
F3v44yxrkFaRnis9Or/ro5ECTOcgbD0x9fA8WLFPBG+oL5CzdtYi/GvmNxfl7uyE
uCNJKeH1QaR6N8OVMfJJRco/wNiihUlSs2FsNN99dUc0Qy8GbE0vJsK7eAktbD1Z
jev2Qae3mDMzJ2WS0CzWzbzEQg1I0mFAz0lFUQaifjK0Ginh5QajVCWuEKKoVkFD
lCHsN56T+J31BkgJoyD+sSklWYfQEsZnT2R/QeanY63X15s9ScQY4bSLUUnWBdqC
VFmcpNEX30Qkmec3fgu+CldgccyK6SJ5cn/0PruZgR3p4ze0ZGThGSuWbLULJ4/n
Jwq0ItXoPYW6dAzy+iTRz1W7qUUC3HyuLRY3HVGybmfJRItA0qPWQ7dP/Gn00P0H
qLAbBQL/k0Pgczqt7Ha/VvxyEJ15qWKhDERFOHEpdoayKIbERDNPVtYdDwVri4qC
f/e21YMo7uZ1dbsgSv6VHc+Qu+7ADHsNtAgnYy10WcK9SRxhm1YdpR12p8+c1s49
BHZdY2Aph/S/DC4EBK/3cxFsa204kcsodpG/NdZx+FBL2WKtnhztPR9KcJTcBUsq
GltE78W/+qQulZAma1XU7kbuMVhAoHCTbOOhJ4UuaeWWBlGZlepKenHjjLwANoqq
030ylegBnGHsmppSlTDTYR74opuK4Z2igOY+Bxf30fHKVzpxVsDQsOVXG/7xCn1r
pu779YRMMqfSZ3TOhyd2xiEgnJCy/qIde6BLoJhsIfbWpVVbqgPeGSciVYjtjNaJ
yjDGVzTroYK6rTRy+7QdDHTbcTn9pf1S4vJ5Sm/8+uYrY0iDLk4nmiHjI7UdyfFT
94czy/H8zS8J68swZIDVv6EByt+n0dQoNcDRu1Rf6PqUXTW6jY+YgIHs7sK8c9qk
9klZCuuSJVul9t72GyuzyhMwOsfh50mrndRkXioTM/wfWVrtEgkUsIztlP6tvLhX
hDIYlGYXiV8hQu4zEEn2RgKPiC8Y2DeNDw0pknrxHf/YQjssSiAGskGEcMYH8/oW
1VD5mUMfhquAgStj/HKg6zLSPbRTVL7DoLLH+LF9nqF5G/8oLdsVTwz0gE0CFijc
e2wDHZWNDrHxHwldrq9dCMH/bh9TrT5g2lP76b88hD5F/CKfZHWPvNsHF/hW3A6l
om5Ghgyso5WomHoc5/yzciu344dS9lHIBYWpL+/ILYERgC3QOtBSrW25aLj4SbJc
Ss8ecWsqX3bVUePN8BnWm6FacXQU5s5aevxKG5jbmmWMr0iL0Nh0AazcogWtKS3B
4M9jpc9e3T+RsE5tsUwgeRWnWTfniqN52T63Yo+60l0jCBfE9FTp9vcz4OEVyHD4
/xpUQVJ/G1Qol8HCB7EvBo+o0CFc2pPjsGC1nbna6RONccuA7Xr8sEq4xj9JXNZP
NNv4HPAYG5h3wyq1m9TOoqp8dHu2NlyYF2HldnAOmkxuT3FwFRx3LA+Nf5PsPz3f
YLE6cth5CRWbx+FOJlcZs8K4aEbfPLCHh3cfbhkRqxYRDAmA+3fdijN+j6/4WQir
PHLMmSj7A7e7lnVSDAsgNYUqeQDYytMCYTRDSw+lKfVG+xeIe5fzUDGnVNd2OBeC
xS0OPoh336MEEInK8TkQ6GxhfYlGqbfbfKt1HgAgkaMrO0N+2g01pzCFEdqUZNLi
hpCbShR2NWGOJJulxbUp4sBpqgGoh3GM3U1UrgOm3BqlovwzL77GmGcF2ssz+JGz
goLY0NlCy6inYFmd4lg6f1mldRZvrdFcAWhV4tkJAIR++MfeKLUjAFtxDSpgF8ag
bgNlXFnkOdzxSddzqQBIUuIAbFpKjaMG7dRiRNe+hST27qGjfuv58S/K/QEMmFph
yTC1noYSQcrxrHwRp0hvBbfh3T8YNylybDLsMX0kUf+QOvEc6JfZAqeiYWXpNvFS
X1Ui+uw27MU1f00/hj725Ej45CtCNVvla8X5Ip6PxkECFeHtXrxPji6uYopaKc/h
CR0plExzqdxL3UjUYqkja2KHY6fTh4PqdrdGZZPGv8WmiOp91ANjL0TlWLwMDriX
Ei2SaYBRh61pao752s2MTCOPzFL2GxZ8lVu6mdRbbl6XXcJJsL1fg/UFYXVVK29y
SnLdBriJwzSkEwMh7RmF9uWu0mU57kwzUV1xz3AeVGNyJnG572Mv4/k5SwRzJH+D
3aMGJy/u/SZZTEuIYm5Ti1WpMlMHIxK+enSqd9nfp1ZcUJ/7mUwaZ7gbSvNWqhi6
RdFs6d4DuZ54d1MVdzrNmwmb3SrV0dljXvq+FnahFzOJaEircRLwCdgo8IsrdLlB
ujYWywdn6LeDzD0TSDFvnK/AXx2lvZ34BS2SqBscBLdogMWt2bsSMU9tzPTU5g1J
KmLMHW3UCgCV1EKhXKFCcg4BekTFW/X+S+KyxhumQBdHOA46En07ia0aFxnC3oQQ
bPxgXOHQXyn3Xeiqykrdf9O1u3yaDS/CObyrem5v08P9+e6R8Fsjp3cTPtC+/VzN
nzyMxnKTlKCinoHR91hvcDzov6EK3Qti3L0dB4CBGfJKsOMsxFsCq1xbKOx53BQC
iYBgQYL/L3fyxkiz6+nPM9B581mBEEZ03iHRsynoYYL7kBfEjBssz8pArVFCoiG0
D9Ddy6hIPIicww8GRhHHBBNtbigW7B3zCTg2YSlABZ73cDmPMn1jd/ZlA2mUSUgC
1d6SEXYroc/QkPg0TB3Ty1Do4deZQ4hgDxcJluQqDHmR2yZEjZx/JOWHwAnU9DW/
hhvrSlxk1mixxPLi9o2Wiq/EVr8VsRtzYS3ScbU8BLcHyUliCtJsK+V/wK7/pk1A
Qxt1mdaXEf06ZzlI4jCl8BI3UEzHXYDU62dV2UBsSPLn9Z4N+blxpPXR4267E2UD
LRCJezqMIybwnrhcfJ8s2uvAuMIt6UMiGXQZCrhJJGNVhG2SevuanLk+jU617/ql
KlhVjkDg3izyiM78e8ndKMPI0q7ouNNp7djNWYND8ZxLm02jX+yzo+/KpA32FYdb
ISmyOClQ90YKnnVZ72IyShuQTvx1VOa3vQQXHBU20AREArxvYqQNWqzF2kC9Ksgz
+wVlXNR1g/OdVIVvCnSJwji7uHXYrqEqPQdgdgixkzaZIKDS1g1lHyf+4QPpHWRW
fe20uhneax29uxSaOidER/cmhqMXzNgGNFCOGclXOFo1JDVYgR77ptc25jJV9JCQ
AkJLnqtbCSMJQt2A4S9ahGlOl1921OwDRoRClSulW+qCe/aU1OHDaiYQwZdCOQnX
r81fgwj0UsOkZnWyE0/hLkIQ2Ty9BM2Ico8JgmgPM3No+KP/P2lCY85kccrOoyZQ
kSdjOAVKfA6GZBxFplfz09qvicPiqkTbc8tctw/uE6fnQCPGRys1U5A2ULz4YlCw
Di9OmGle/BCXR/9h9B7mKdaFcPJByo4gvOaI+pv7BfyAr19d0KnvFDTZTpPpBlM+
peP6pxDZkcAUF/WjaTqEgp0zkzR0y23US8CzzbyVGL8oCUCvRq/UKNde3I4r92ZE
5dzC5gGmZL6iYOZfZmAxfc6ILCEv6iTrlz1ryHG510m1/f2YJMRJXK7uCSk1pBvx
AG5oin/g+hYUU+EZaKGaAOy/u4Q6du/bf04MvNnKBIqa9USO0ZOPQZJ1QTdQ1OwB
Ch6VaFCXWlyYstKOUAjhXIgJ+Z0nuyYJ6epEZY4M5dcKckpWfTZKtKs5k0yq3hpU
NtwIvUndyNyIdpz1zVyF+rQZeVd9gQrv3ruc+ZFq3JKT9UztXnFZMg/ukVI6UbIa
TO+7LSsuo+FFeQkLphFkfNF43M+CBadzUblKsGDT3c3i6gWNxuaDYVkEdL2TtKtb
EENMKFB3Z6GDvyHHZHwZNAdxNUthvAkYziEGzZ7BD6divFgenyJcFM/QYTX8nzML
ARNKsjONKC2ZU4zB/TeYFZJ5eWmcouVdoV7EMoTOcusxSbyIbU4zubSH+TDElNUR
xHOnbSeIQ9b94fjFQQY/STa37XY7912p05V/snJuOAtUAw3g0GhGAR1CmTyv7ZeR
kJ0Gb5sEEbsWAAAgc/qvAvV6dI+tT8xHP6BKyuzGPQS8UnDMfrZ4VDzqTYF+GlC7
YeeiqiXc6wkS04EFO3LRpMdjKG0SQgwl+LkiCpiNsULdVjl1MZKZWbYde7/sz7VW
5JwNrxSfwsYjYYGtst4Uh1MjmTmTakxBL1XXEi5sauV/0/KUjwsFAwRmKD567ws+
Z9bdTLerZgXcph8KhVYB0uOW1TkAip2KV3txz6mAAwQyjf7udhfDqQ0MQkSTiZK1
53W12LHwBgahGIgHsdQezOrJYIn8k55VyU2tO+49j/KW5uWEJIG1riBlP82olgAx
K8EGzN9CXFCiW1Nb75RHNmSvn67SO289scJ0nYPY5mCa0IEQc3l1vxYG3jZ4hH8W
NIqG3SAi3KMhUycXwXZIN7z6HW6UhgCCRvdIOgOw8pBHQrXZy3QTjtpx41J9Z9k1
+y7ISvxYWKO7mSaJ2acRAQD5g04CxYiYtUe+sd4dUYF1jePdGBgKbtBIDPmRbNWb
w6OwafnYgTxno1431tTWpRA87Qn+99yaoxuHowxaLFck5npog9Kc+vL6OGccQzjP
Pul6PFQFX00BkY1NNHyVBKicV/hWjDCDfKAKl6vsyhXInc/d9sRb5nvsKpHyi9Qb
JW20E04dpc7l5Ml0fak1OKrwAXkpFudjgLjBgf2hHfJ0p5Ixpbqqo64QKh/FdpfW
w8YWSQv4rVR0jB2aqT8UltTt3zssZr8asDvXbdqcq4HOikh2wgrD+DyIJVbnWxLh
e3WQqn2+3e05cC428dAsRzNYWf1hDfREGeEW96dofSt65wB9EPSNfSNWcivLJO8l
NgF68zUKdiA3bCL1nHexsx0Qe0lKgF1Rr9jD+6QrhLNm3YFgDmwreHHKCbYJCZrD
LDXykqqJ+SzXTse3+kBCUe6uOkXL5IovCY52t/5HLI2dgpFOWKGK1ujyjelzVhNx
TdH+42zzHmIP7ht5Hhnr82cNUksA9STYEgKaOUwZFgNADyYOgeq3IPOTBAKGtGJN
9L6KqMS826ipR7mfUau0QHURU8uElBn4PKdMmTTKn/h+OSbDsZnzlQctYuI64Iwa
gzraaMOl+SRqWAOy76zLvIhFOcyaeZY5pE6i/GvA2HYzXIbkVfzEhOC4L9GzVH/Y
ktgwEfTaDR/sLiRr6+Q5a/ssVD1k11rFoAYrjHJgg3x///uAJK1Zr1Uee2/iO8pW
67BFcZXiIeNhYJVaImyvjvX0BiHARUQc+nkM6PynLob1Dt3gbWErVAOVbunlOu9C
NYbbpOJYCZdxRWJEytcrTndCVsCD8J1fXIfNktQLM9p6TwIKHHs9lK5IPQJ7u/QB
bbaSxZMnU1uCQaYqpy2EGm/A9iK+5D4dWx4W+UWxSa6pWxUJCrePOdkOzLXPzcFr
LWMG1ozQL3dQJTHE80lT8gT8/h+IKLLd43jz+zccf4gFN/6K870c28rRNojQm224
E7KqMMNly4D0LVikRbE1Ag0y3AFuLYLoSJAPGj834HGeqgQKXDDlENQFwgnl1wbZ
SufnDbTsYI3EHi+3jY69vd3XSStBzc65uwRLQ6cf0DmGV7yEZ1MdhOUby+Amvbj9
pRiRvaqYk8VkiMxULYl/nYBMqK9awjSCp9HCNvl1URXfDTMX+2WiyUHoFDuCGJev
zxeqVbN6uPpsh24qQT97vObnMGIKo0fBczK8p+dnE+yNn7wIQsEk3IMQm3WrPHd+
66u1gu+x7Lp02XV/T9/3qbz6h4ubaScwsDjSojPC1S1fmOlP8pVgcGKsA9rvn1+X
IKFrmx8PdsiBhV4QcZ0olokGeMxzP/ZegWuIzAmRdgpz7x2TPcBXkmBn0gObQRQc
i6rfC7ISynWQQAAG4Cvo8npuxxn2lRCFQsFA+kmuhbyp3hpieAsl35AjVfnzpnzp
L/RQHQzWEpxpsvwvD+AbgQptL42/b8LZwHZ63p4yQjagoz3izedhMtXTOqHdLKKV
2YaExTIt5dbQa23twK9YSQX/Bqu7w5QnaNMsE4J3ajIfw3WUT4k4I+kcKK/WUZZo
80vAEKLxfOj5r9t8/eHzFUDRFI5z9T5+0G7whQy+80VXIWYwpriYzn9qVUylAlBh
tNtEzc0oarQ7K6BlNwDXxtjuRUrHgxupPz9TcdBCkxWh+EqPsnxJ1QKYP8VdO3xh
rzDeqdY66Q7K6rK+Wt/uvh9akuEXOOYefOiNhx0TTef/S2jxA9Y8cNVFSHCDdKLl
wLOAoO77/R3s6BnBmgwfPfI1e0nF+b3X86NdK45lh1h4bKNeL3LqP+P4FJE/gUb9
1O5V9nnkKO6ZKV4hD3QunDCWmV0dXoU7m9zEVIP/Jg25sPNfHsp0E5vHQcDfbvvY
0wEG+ki/SCmJJ03WqrKKUExNS0H9vUWoEcx4mCgbsJmEDP6mgh+FzB8X4KCsdGOI
7+BtQ1HRda3NdQIS9brcHxywcREVITgOAwYUC1fxwlPQNTMDShxKc8QN9b+klNH5
rpB2mzUvWGDnFO7pHpYPnRVIJ+diqRsXgV9CIz/b3IEvQULoBdCp5AQtLwOZDEBj
bfnr+SWCcaoV4FcYkEqkajlmTWbLhcVJLLo1eHk++aQRzaQoAEx+8xak0UFPqVrP
OLIq2IekQiX+F0XgD55pXn7/7S/5lVlbP5ntdf/xhGdCXqt17TRpqOtMVX/1I0sh
V+XALgCbuaAXwlwMrtOp/2KU25ZJjAb/Bh7Cqk3tlttD9mL4B+2uUWOE5XoCr0pr
lz8E0MqnkS4ERdN/DpDwlqOaKMZhGGwlvF5dKT8C+k1vrKUQig6zVOMXD3oMSfGg
VFPTWxjTiq+OQtP/P0X/MNQEu6CaEhgkL2cFv9jPrJzjeRBj8qAFw//51IeXQ8CG
2y7EGs98OptmRZbCrRviY5cBcAnygipnlYtusC+Y7XRyDbeGeweBXjiV2pLGmviR
cspkBuDKjXfignYXbekmzlSWRbqqSAcjvXbIbx4M/d1QNWijPxVEqq4orOIiai7U
vc0hjmoO5y6pBjHg/rXmjUkgZpVjpQKNUV79+1HeU4Dd9JMmGSyQtrUthBfd81fs
Li7OucVMCjhMDi+GZ3NWZu7VlLSVyHQAmK/J2+453Jf4ZpMmuAo7oOMMJsZe4gOr
558jvr0ftwDKvLMq86o2xDAGy4XoUJcNBBM4pmD0uVxR2MsIJzYYz6SRtJbjdDqI
skfsnZymLKI9yAcBxCcKUARCoaEF8tEjClGQ8Nr4vhiQFnO44hWY0pYEHIZh4sOM
yPXweYuqvwQxKI3kjR6AJmSs9b5gAIDJ44KEJhwysWZSJ3oENq+ZPUI+y6S8ChC8
64cfzV4IO+LShvIR70tNIDoyhz6sRdbWp62nJjfj922+WrAY6m859DtLzOaMyCmr
D/v61uLElEWOclNcymQGUOU0qAA4ovYqKz3OUtN12rJSV0YNZJiEGZ/hMGSylbGI
BAuzlt2iJF6+JPg09uTmfdgCW9T/nE+CEkAQvigqc9SZs8siKd5U0LJMDbR8Op2C
EEqXwDH7lZT/NPxuEocz0cYWqW2vmTqmI7/qjwmfloaFfqRvNxA5qWZmeUZ4ku40
fi7Qj2WEr1uYdIL/jPTeQ1CgdgXO3z9UGiUY0XfaG5Yht4G3EIpCmkVWwWPTTqjQ
m6f+lsBBXvaCUuO2w4Xr+5aN7BzcXZfYlwXE++r0X+p58sdeHcf3gmvhauHXyW6P
2l4tBKtLD/8or5ZaGSvUI2nySA6JDW7rciEKE+xD/qtBs2zr23sWlKINgd9R3gnb
9jyiPEjGe4Wd4QWGopXogoqtf5Ms1aWWiq93D0FnUS10Bjsdw0Q/0T0MPkpYsYos
a8p0ydN5nNoeGrwNO4ptzr5TjGwxQqqPidH5jMOmJi18G7YvCjdBjJlVnjipEdaF
wyr9G0Z9q+qPl99pi3ac54q+Ga1EkxTmKHEcX0OurV3NTTYGpiW/SOnx/hTWQB96
p8YUa/vW05bfl5PflNin1nSJUExygkPGc0nWHb3HAnPD8BVpbN8WoHrFu7IdFAwj
hVAhmMPDf3+9vPE/AI5sOWy+fKxFbGLbRF53pGfpbGt02r3uFfrmDSr4haDjAnoe
fRYRRpc1hlMNy90xSvaO7haGxJbT9jNrjmVKC3WcMYaY4f8TzVqpYh40ZugrpxSV
XvIGyvTuIm4qtpJeXNxNjOnB0xqdSaTTyFRIiTaTYAKiMuShgQehcIjfk37UO32u
Q++KlzIPa9vyOfaXi6ltFtQUpibsedFUvDeLDL1Op7+8eabZLUlFleWzgPgP8A6X
7zkoMhOGGKC2LHNIgwiqu5EsNsJbJRZGbOzVj8VNz2xd0hW0jN1xEXawfAokN7Cs
sVN1essjOHULrojrQn6Nmb1iesBIFsv8zb+9rKblA3bgchRsGug78ChHkWA0N2Tj
lEDIy6aVN2oiX26rsar3JPjs6f7uQsZUb6QQhgslnqr6yzjUd5sZvoDkRBNLDSsX
5SiaIm3yjTaQtYny3wYdkMUlReHt8vdB66ncKDceKWJ2XaUb5it+9le0v6ie1tww
h7yn1JmqYQvwByXnSZx8sIj6wopq3l5OtoBtEJ94/k47a4YQUqBumjas4Bvei17I
DfUK5K+yL9BIE1VupBlsTlUPbqsfAdH2ImAu/AGiVoJKPfJqdUm4Bwh0IUhXB2zd
Bz32/+6KTud/CbRGNjyCYrm5yKUPhaVvts+7f7OX4XaKI1lB1sismgfU1KGP8UB6
vAHblGVqm68S8kb853LMt4+o651yj8OAfUiwUz/m/F1Y+p5akW39F7Ygdy0xYEXd
pppIcLkQMFVjBwSQ+m/NQrlm4cduaZHdjNh12foKu7j0pRloAD4zlS2EiMxBb2bz
svm4mmxCMVxD3wNGy3Ubs7Jjk2fs9XcBQA9siC+8WXeT1+xZHcZAFYTUKTtM6EbH
xnsQER0vNNypV5vTKij2OOCWW3gzsBv/yi7w/zWIKwhPrUSZC6Cf61d58JsvWCUf
0TUOCbzF5TZUeKW7QFeEM3Il8wem0gt+uNGvgJUJSQulXO79Ao1Tvaa/sdaRj11s
zdRcSb4xXkGrnzfm42BYZ2cOrGhJjykCExIKWEHB0pIyCMTkKlOM4MPbB7xkfBWM
jCH35DTRVcBEh2gtbxlDLhTLfFz9EygKi0JAK/qEiD7zTgBgNEenKBLkArVjC2s0
KLgDNzYEjKEvjj3E3LdAvotetTRUw9Vj6dtHWaLSBgLSJh74ypPZYGtuIHnwpJpc
VWMcNTXUQHTgKZks72eNCxpUUFvpTnhARyxDBynDwhPO2FporH9n/fS9ziDpSATe
qgenfPZAju33mLkdJ/9n7m6L+GCeilWAg5FJkLF1uKBftnfcpD8Mi6e53NvzwNKW
632+mCda95VDsyqEfIDklrZ+pRTknhM/sBMaJCIrARRrQjHYh05p2bsVbb8u/Awg
QioZNTtv+pyYkFvLjN0skyPJJ1gz9hOareoYXAKGz4AEk6UVEsxC1yQxWx9CJxjy
HHQ17Ezy6tHXm9aC1sBtQGuZGkDgxMiZ6g847PcOnzt0nPxf5SfhuwVmJ65/gHtm
IbhwalfwHcIy4o8krFBLYpKjLjGqgKwsOR0Cq+bLix80N3loGMWvE8UFJZCLzON3
t4fmpH3u8toMydkj4sHWa+/22YeSNmn5tSKwykTtKKq4pRR78cKKiowAhzJopNgK
HSlIL+1lLnbptXFBcZpqZmNxoE87lCFBo5kkNTTZH0arHrdWyi3xCL3r+/3zgMX0
HGjzNI1q74GzMGVuA+oeZnqkI03bN3+1MdCdyTapoH1rjbP5l6QJ+KRcr/n84eLx
1VfrUqrifAMB60efHuozqG9XIazz89h/6l35g0DenU6T6RXVKnCEII2Y48SOJDyS
K+a0iPrTw7WThYBeFqI/xZ1e0vt95ceUqMNXUAq6qnFEjen9/d+I8BOxkVNV9N6Q
RYgWInQi4HCOkZaxfpTevMARvLAObJnlfQEVY1h26wvOI1Oj/isgHbqFOby46NeO
nmn1QKAE/cRRz/eqytrpmTzmasGDxBrKppocnJhZR4gIhy6B/Oht0q5X1D4sXtHm
twAW6ZgX2MK3G3jJlUbTdwp778CLIXAV3Z4mA2at1Am2JTdDumVtIAC+REOQk/nV
XQ5zej3RXi6uWIGbOAPRE8q35iY98QQY5DUrzqc+CxYjSIDh3oNUnxF5ZxO35vPn
F9VoMFIqmRHuyPaa62zrNqtr7qoaSpC1PEhOVodbgNtVWi4GLovUiaVVdelWEJH2
nyBxdnNDZQJrIjvAT2GHeZh/cnVUyKhx5SZU7PlwbOXQ5jPNAKzURkiDXlfTggnk
9luDxL5CpJXFNI96Zq0Fv0MFWWWSgfNIhtGujCUj61Ia3UKzmXo88YtmDyU+Esj+
I3hgDDLrwan0n3NVeZDQ8dVvRbhXGT524UgeI2+ihAE6q32Q1ZoVbhJVJ606qm5n
V8Wf2l1ToFWaDI3BrvoQLgsgJcEz2BFO2PvnSAth/NX6f5VTxCvyOaSusILCv+eq
uR74CqLkXz8TSXVznjIbjt5gOBA2BJE6D5aMyaB1efPpyxcyG2VrMPrd1flqyleI
tnqkqP6qkMdV1w5L5smLoZ4dz9ch5mo2n+y6Jz3Jv1Mm1mYyEjksHvzGZ1n2w73a
Wvd8JvVTyQzk6vD0EUKxnKmY8QPGEy8MYZzKLJuhbz6WY/N1n0w+UemD32pYZBxv
hty8Fpg7+lljZzmy+GJ/tnrdn9bhKKVsHQsThS55pYCbrIiwcOrpvVghIxoDBSQL
TuJxBQt0D7eJQcuxoUyopo+In7lfV5tjSSHlk+f59rKcvEiss8ZL+yfToilU3Io2
+enlHV4KrGl/TTszUEG0RjGl67BQBeScmzy04i+Hq4OS/MHTrpkjPeO1uVqMBPjX
pfExMo6DHJ/dPudrhhbkRes/zTcyQgrGx1voIPWzJg40PwaRhk9865+mEvq5vw6j
KfNhvGd7VZ4bmDJAWNEwSNt9WoGyWr6KJv2sfLgzvoe78iXbnLWfNHrTgD1aLfh1
qhCFNtokinEltHePmSibI4tOsHerR2cYF228HwZA0suB9JDUrTFHAp3sEhrLT3Dw
WfbVnVsIFTzdZJcBD9/W7pAZ7leYeJlc+SURdBfPp+363TF34dypuJI+Y76y+jKB
N4V7SIJ4XgbGaHwGBMwKLnYJKi9pivOhK7hOnIAvjo9bEHZNVqHo9gcN987mnX1A
4/p52SXcvZU1UjMqZNpvGW59VBWV9lSroboFfJ/XWbr12X1s5vSqoElxuAFijtoh
FBSV1lM9ecwFLRKyHZF93im/LC/OI0Gp2E58j2zkBx9JhU0Sh2kVUKG+1p2HutYL
y82qZ3+5rWNDgFh8gsdt8TZ3GX5QUk3YPXvK3nXoBPzaxSxCVxMnvle/3yGy9RA/
F3fuwuoHXk/lskMKFx4aWwlCPPAdtVxUw10vP+KQyLCWWbGI6fYSr+yaKaX3QUOm
y+P6yzDdXI9bpncmmfJho5M9mnKARPWekpFsYjk7LOoltGPl804puIiZWW+s5FEe
Q7NlbMYrsC0OWo5upg1uNT4tGo+BltkqGEk99V/AMDEHLDOYTkWoLztOGxMSEIdg
iRNmayHBv429DiuHdPaB3LCI4Jd90IcYSWizlrKPzaQjPaL7CXep/zERz+XjJ5gA
Kyaz6Tt9IHLBC4tgX8vnWnGT9ju2w/a63Xb7RAXIDrVgtj+MngzIkloupjvT2VID
NtEMRJz3KHgkfla6itbx9uJtEmkqbYvfB2Jn5dfa87DXunFcaSoeSPmLj1xUmHNi
rS7O7sqc9Ad5bx7cOBgOTQAtVfZSRmPlLtCuvoVXUmwL9PngUcTmBjSGAtoaltiy
ZpmY0pnM+Sa2FkbMZK7pwiqQG/KxWHis7XlmErMqgzA9OhaKjfcDY2AFpMyon9c+
g88YTVVs7Sy0dEd5BRE8uN0GLn24Ic170xlrpSYm1Z/P018AibN8nSiUw5kMzAsB
pca+Ip99mdKtBHWXDTs0/uB1tQtWxn6G6rqt0wMXwSDHiEGjHFECUQBn1KiZgnXi
urZtFnI13XaFNQ61hHspPyoEPgelqNgVZKLDLd2DJ0LX5eJfvBdagxo4aDwgq1/J
lpFR+U1iHbCtmskzrO5Y1U8te3wAH6szMurbCFNc57D5z0kJjpszBEgjWgOCaQ2C
U5YueEytjFI6qxtUtF30pHEnyykcpCDf2+MqiI9ZW6ivQTPztyuX1ML/Xs1fJwgm
0//pdiEJQOzvM/XjttJb/SUM3qgClzdd+L9JObkhNLnbJKpn71eWku3wMqXKcTpM
qQFFoFXwvu8UTbGxv3N87Mpt7Jg/tIGJAW7YMB94gzpGhkBOfChQYSpQaDdzn/6Z
VxyS9ODosA8QipHhINNwmem6epSIekh5hmsd7Xi2MVm4uw+xZ6ZIoLPpjHh1kxju
+y66zD8lQCsEuAYYF8WkbzdqO14vezVLPVUS7+oelsvzthWsHxQeSVQKp4q5DZGH
eH5txOblJBt5VngM6mN7OBYGKndqmu3qol36G0ioX2pTyd/LnYly8Hrl28b3ZGDa
ewTjDU02TbHFt7as4u8LQhy9Y5aJF7iwt1cLGH6yotwWKDKqs5ZxsJYAx2tp/wAL
PzExQ/+Gu0AAZzn8zfLO9mVFqyJbOqXA3akIJUcrrzt4bU0leGd3368vOWc6Ltb+
9ffwOeiPa0vjdtMBXFVq7wnioCUruwzjnH52kl52fZqAW2ON5wk26bGnBTWyQ83J
JFmYMk/T8O8qRICSDePHE+A01X1XJsbCx3C5eWW1s++Mw1Cr2AmyMsqVPlY2zZMO
kpTrx3ArIGrCs7n+tnrosjvITRHRaXpXLdho1vC0EguxXACm+REr1rAIUDQ8b7Le
plYaKPF2Mip1wltLiVcA8IISBRzBzgTgW5HKXuBxbzhgaCVK8S3rhYEGoyVZ6zGk
51+o7WAdmME4MVMMQ84gTDBH56nlOwyR9q/v8JX4eHOcwZNo8Nn2FV+yzufxICdK
8hFl6/pWwuf+gf9NscVgsd716c90dc20DFxGGRtzrgq5s5Y57PxATPGQd7GfbH07
U57o8IZTLRmjOXq0kBCuR1VNimHDW243nU8J8+IN+Xf7rCTTh+aDTHXG2iUhWDwu
OGF9DK53C1a6SCBvbC86PYAwkkf6w0eSocgoN2yHQFm3+NsX2kvWMcxkBJoKFx+L
p5Bl18/P2lxuxuyVsAkK4BKYB+XxlBCu/f/a5+JAuazV7gxDpsh1eqb8mBpetI8K
WRff9uzGhqDOPoHbLQzNwIHpSYFVsTqrdPmoJEGqykPGjFwhsXxFNCxSqd5IbH8M
bcwin/46MFYAfiMn4XezVmN0EizEc4OG5iQ2TAZ3amZGsWh7W3E8V8TIRPZ7nCDZ
4xto3K0NmJ4HROCo+g3bzNB5CXI9Rqg2f/rOM+gM8U5R+dTW5Kg5EDGUMSxd91qZ
5cXMhqPeSVWuMq8iDlLfY/vfYqrLRvikdliXaBqdQiOnT4A0ylUfqKe28LPTKBh0
6+GWUhXbxSq+cOUreDIvGrqd1+gC+BTpXss7t6dWBMDnJ4UmwSdhqGPGB2bbi33Q
mIGrPi5U4o+F9tVY3JyBxanmzLPEunkDzom0SU0vU8WL4/fIjRWwtYUe9Uefxga5
L8k4BDC8hm+WboNzRqk8J9ZBNKW7cD0zYkFPm6eigM6HDTIjxjeUjWQDq9IhDH6w
Yxsotvloboa97Do6gHrpTDicAr2nH5qB2fWz37W7TkdNqlV/+rlHU+enavwqudtF
JJT1dMhUwBtu9GpBQjnvj/+RoMUHH1F18o2v2adAVDKbaAkIs8jMr+m181+sXrpj
G7P+zJVHJZC++QrzYvxoQoUi+zJrPoBiIGeWuds+ANcKJz6w/lDiVtZT/aVcXIQu
WZohaUXmGTxluRKCvaMZaEzj+D9hsvdzNuhSiG59JOeNaRVKv1pQjS2j3r6rA1PD
Ax7gv52YwRUdkYOZQvWnqFXRNwKuwBRDmSvgzyvnwXcpF3cgzXizkJZEuC+O/e5V
BK0K7REhqjVj9POjkKEGyzM3AwQeiLr1Tr2GnW28Xfdv5SAcUlIzvRQ6zK6H7LUy
6uapmr5hw5rqRYvt8QZe+HM3PzlYJ9Pe9F7+l1mgQq2n4gAYNW4d7A8JbhXWiwrb
0+5LJzKoGoolMabjxwr4QJTB3U5ND464P7Zw3FnLKP8XVt4x1oh1W+t+XFWouv3s
Qw/YRLtr6eAqWYeNiTdixrpDtW+LpwFQLzzu3I3ZJes+fBdhUNcqg4E8vxCGrAFB
cZ7GKp5htPg98w+UenhByEg7e63tjG6/MvDqRpJzH5WxAbutCq0MYXlLODhXsqc4
4B7WAU/g6ncuOZ4lMsCCjsAPrMNbeb3iuNRPd6XQAtJpzKKZ/uWiS8zYztEr+EEp
GQtvrLkozo6VEHPAY4REE9VJHzEnljLwHh6RzErhZGJLajMVSBlcgcSZKKY6/KFR
YeIplff6s8zShTzRP1UH9Rv/oVMIR3zNSefi9zWU8o8GoG7yERnIFAsaRI2LMNnU
cSu++KYyTNwKa40usgKW+aqh900daHDdj0mfYIIrTAKSumxAzeRjpdaCBvJUGz/T
8/58X38zwAMGI3GCbgQBb505uswGbkpQBL03HUQlET7YmoId5lB/RuFndoN5J+0F
eB6XqykXfaR+pLG9lczwji+p/z+5Ibh3zUXi/yGeucK/5w4YKx5Q6+Tm+vgMZSeH
RO5IM9rk4ruodMedubTFVpIgHXfRJU9cOqKsim+1LoMJq9/RV7hTEaz4XA8lOyuj
vrDIuw+H6+5PDOzus/sFSqm/ZzGVr0kf4ATwLuqIDiAQx1rDmHCAWVwgFpmnSSzq
gCCjofnHhDjw29kfjfRBlnXr+WSrRA7TE2DZuFyUgJfydIsdmux4VSpqWXBeh+gU
piyMHCqJXZ8FOAY+apjgaiZW22k/prqfpBOv3sHG+3S0HLl14O+VKmxouMeCVMPi
x4Eh386xqMMUhdHcOjYInFJeQjiihnB+DGEnF71dZl7NfjXG+7lZupXWHOYlzdgv
on+qS+kxB2j6nsDCO7UxUYKuMrvFqYShYZvlG/A5mxSFOdVFaNaI2mih1wt4bwVV
ON1385kQBiF4Wq3csKUNFaRi1PvICBnqOVYI5u5Kev9ACeUTzfnSyANJKhGF34be
RSLM8LEqCoankBARtdPsGOExeOvdxrYSa4A38cXEZUOQZfD77IQxvj5jJfFNdv69
LqJuDfZ7YuWns0w/cPwYiEyj87EgCkhXDJZkXweRkVcL9MZ9OCsYnZ6+sHL4HKO0
oILpTEKx2Yknx1tVOP4YpQPHS38RF2IZqFSEQcJnyq6EIF7Mgwbb1L8r9K95eOmP
AQutWOIVW5Coo1AALIXYjCmjJQzulJkUKBvbo1sIUOSYbyla7kS9fjhUX2SLqnJW
yTlO6cuPHRNqWh64bmBIaz7+CfCCVuCGU8nfPbV3OJBipCvcgmw/jYbA+9P9udaC
PdvGRVjCdcm5uqIOLIgrT9sR6tD/xJK+AgtrtvVTDY1eoBgWTUsaSO6BqsBqBXRG
N2HPkK2uWwBdl6VLF/9Imky9DU3KtmKAiZm7HlPfWymReZ/B37EGboi5IhipanTX
SEUe0LjXa3btFRSLkZRHPPeonYFhmSko24EXEEARlurX+vEbVUMQGuIZ7lmK5QS3
2oMSA9qwwDwJDt19gemhaFRqMEKuEyckXY6TTNMzffgQP0Nw+aRXtxQqO1Kb8xpe
6REhiVy8DmaZkmiM10qABLrrgD7rMqrVMmiWtn+n+d+e2Q8OgfGozYqHaoLXN+++
P2qPv6lyMGFZXmZBaiydZxua7pKeuLkD3AbphH4r7e826u1Z6mvhUiljmUe/ME9M
nHGBIW8xjOqoaokKpqaBaA329mvPf1xEofpKh1oLkyZEICtVDb7LnJiBB51VjYZ/
9mQAJeeAha0PrbEV3HdSSxcTqsBsqKBQxsoDrLVmjrkX9BBMzD8t9JuZfzmMfXCB
gGluoQOE9NPxhBH6OXPE5gFPikqlMs9HjBdV1ZRPs2lHmeOQdnTtkkTZKyW28XYS
kkVP9FWbSeulAD50uw9KSplmzgz4e1+J7bHX9Lvhg2xmWP1y2J2jR7SewfWmwa8h
PAyuJPenoEwnOdwOhNsf1rOogDptWaFXJPzsxY1E3BMEDg+T5+1O0KlA67aCpuBQ
mfC5YiCslnKaGTrTUkqT9K6EcSjzsdV4i6P2JNMeRZPFLCI7YFYOoas7uQ3o3yJp
bM3AFQ75n8kCi1ZrU+mveILamYdtdn6zN3/PcxEwGPTCPbzstDH7rLzDXHrSq/Zz
iamrcSNdNIk1q1Z3ayhN58OE/ZsnyFx8mmxXHrpXglsSOL3IIh71FF54XAG1dEo6
7Pu6y/8pFF2r31RoNXrl/ezoDSiTsaQYav4LHIOTZ6+ZUCqP2XGQZsj1Tm1TxECh
lYsSccHNP77RrGNaRID6NlFEbGNo1UvrSICMYNXfmYXcXU3geORwpMe0IrTGasjM
CpSVcpyywLdZ4M9W8+AQtvh9ghW8DVSPOT9I7nJSiltVOP7WqBljcTWW6Hl1eJZ2
4EX7ulVvmY4xOjRFplRIAj4I50aYxRNtGUrnr5Cpgi5gw0wwFKOXncVhVBSwMg9+
6B05lCe0VqTM7A0+fUcVvSJBmrXhKrSlYwycl54GTFQC2cCR6umzj24HKt5PYLOe
ILnNCCL8n/P/sfS7YZxUTgncl+4XeSaJDba4uglBLC3vpnVvEYbLcAmPX5Q2eXVT
UXXTrCZlg83km0eAflNrLGjoOT6uRVZZIsgPlQH8+tK5l40Fo0+fAyqDCUEbpZoP
6jSsrPoPBqfuoy0ZWDSjzyqsMFqSsev3raiUsOUk2x/ZJGbjvxVRJqEryPosW66X
vgeU2FRKKAXn+fIZXtA3SuwPNrwbQQmB/ONpSNxfP7ABXk5ayKw4D7GFAUc/vL/q
Sy8ABOFex3nD7iB1sN3a/0WWWYLajqxLrYUXfXjnJq+u0pOFBEC9SdyX7pZU/ulm
jl7GNcjQTgA8dwLlf+n+TM9sIAKRVPGHeQ1pAVe9tycEOUizRhUbEwlh85xEnKbX
grWCetMaG8R/lu9pkf53BcNuEnWmwr+wAzNWaApnY8zo4TUnzSHQ7foODdpAd6It
ohihIjpMJHE341Y+7VQGIWOFOYeb34kwxhsrGzHWxEc6c2wDPtJ9lIvsNxepHH9r
JGxMkMK2Y28s2yY4nR5zbpmZTCdLZkeeXhKIi4Kgm9T8TFyV6wZDjO3ns0kSqJRd
NOiL7e329Ny+UTJmxuO9vAlMXQim49i1npeKAxMd/AO5U/XQLdonlMQjOGxM8bn7
geVwuHCpAKZYjYOV4Kdu9nK/awWeoBPY2+DSdgZmeKD1khiA143doQR8oMIotfLq
hmHQ8WttWOq6Tqb3GoPZkb7Tz337lzKGWbRKWzy05WSnsKCWu+ocOP5U1dChSG/4
NetueTpC7ibRm5vPx43xZG+hQk6JDM3tUCwTobekD5xp7H6XxW+k2jslK+aETwAD
H8MUo2FQvYggcMoUoUCQ7tXndRRx8UgMs3VE0wKDcaj9U95SC++PZmtbw1qKucXw
iVtdX2KEOzBTeIFImM8IeioNp7TxRXfBww2kbr8ej6F2rZU/ikJoVrTL8ICHgETm
rzdasz3/f2sqZ/HS4f58uwyTbR+LntbHqMU+oMaCmFUXDcEKCravB95aoNMG/oWc
ykmp+Ca7Dy69X7wfK3mbY0zeSGz7tPCdVM4ruD7SGNdJf8X++PWBnP3ZNi1dGMvC
joAeUPxFaD88P55/LidiyebctExd7LVld4PNTdJuOXFKtLH9Zb/0yK+4k1DTZzNs
6jD1vWx8Or9Uwq+K6vMq9pNjTcfxTPMEZtj4JBZRm8umHpaxSibOq3CfdNllSBvW
jwVJyCjsxrXDKtYT5kz2/hKOpSEIfm3Ks25c3YOk7fiweNulHyykSWuHEHl+aPTb
Vd6awEdvQAfmxSRdRGWM+5UesM/vhWAtHmS5GKJ9DfZx1rBAaroX8ksBZWjTWhom
Pb21NC9TxnyVb/xM0mfbOcvQjDmoX9p59qp4G0coI4M4aoAH3k0u803D8p84MWgr
xmT9AvdU6zJuCTyhI3iPkW5r9aWOC2NaY/9xMoXRYfxVKwY5VLEQqKtFTXAqZ4+D
mJEejG+1HihyVp7/FeN7NqaZefY8oq4GWx2dDtPL4dxxcnnAdjhv5lbaNKQCVqNn
kT8Jky7uETVHDXY8wZpbcb60vWX7a+UijIR+rATDCRDiJsupg0fgKv8z3hRQh5yH
sBo18cxXYKe6atxTX4YVHvpQu/Gy2PH1mDBERJiEEoZDzkPbad++lMusoq3zqVnv
MS3CYTdQ83LMp/lKiRNno9pRzaCKbT7tKWBaKMIJHewKm70CVwcpju0ZN3pPy2fn
+qwqUHnDg7r6rtowC5B98Db11eUyWHYnDtx+oCpaA2OycQrzNTi5XqydpDQyhdfu
R+N9NtJrxhQVuZhMAuVvvnj4LXSNcWztqTWiv2dx3cxl4dFf5t0ubyhypmyJs/3d
0qzO715C5KyDabqDTgkGQ7vmVcGLy02VucfELsRGpYwksRRL2LEjIGc0luGp1jHj
edgw1YTGh/igMm8tFD0NIjcqgS1EBAQmoTUaxYeI7BbY9eNS7HwCFN7cqbMi/F5k
u55JM9m8aenr8BvXDcjhsnufHIax6xMLdckLPBx4WWBwGaZ4ETFx8lzfUp2762UE
aUXioIjEkFyfrn7e/OS7Etw8ZPFVJTrqJk5cMcO3P8BRHq5N29UZTcxFQEUPa7Kf
Zn0t/Rjh9yT8QbQOEp/s6JuOYVPE3s1DrFummDq0Tr7ze1/6aMrirnWfgEXhLrBh
0sIe8d6piYWsg5vJr+HJXAiYz9Oqod/Xy22ZqE8m3fLQOcILdlzCMvQRqTBbTRVs
lR6DAlkbtHeg0rAAzq24CmlHXTTIayWEiefx+qqO8or/iCNKnS1x2h9RKQ9mjbQg
rAPjmeKcscJK0EZIv691Tq34MzL6lXEl2e7WKkyGgh1D7G6f/XCBK5X12OE3XnUC
ldXcvKCSB4l4pxvyY0nUCijAsMzrzldTNpdchDZuDBhIcOr8QVssX1MjCgi+pBHw
1tGStoie3sklvePEmxUwxyzTIQOKomM5ZNct7pXiEPEPy1reNCz9dRttrr2M2MBt
bNXX+MjkxFLCmnUx4qopAPtXz7Pr7+68GDBdApWARQaiWq2eYVS4fKHyJaRACSA8
4pQWG1ir3bpm0K6hR9O7sU0bV7r2kSKTmTJ9rnNYTqFp4NTktGC+4qKXH+oNxhbB
qI8UYp2YOFj1coDTqaKEvFCseiv9s7joHMEhAbEWTFND9ebw6hGStlGyGXyvsPWt
3npseB0/qJmUlbvqpnC6zy6k8j1rrqoqAzfsbrrW+ZKylasu8ozxrJ6gx6onAiyu
0S4Bh43/wrbRJrcwgr9u3jXB7AqGSy3KaTW01nqKHq704Sk7kREdd/Z3HX0J98yI
K3OY51lMzGfY9sUqYkPY2QHjl0PMyr/Rnyu3wG9QrjclwH/AYvVkiII9MMPN/ZSG
ad3+9NAIZzoQ8humY4F+801WXCo/bg9biB+4ifsG3FrEEAvCHTsMgb4r/F1UuhwV
YWPUov/b4KeWNPJaG0ki1b3stusHAowxYwSwD2SAO2F62UWrVHtkK6CaZSXmu1O3
VFV0nxR3y30CGNvO0V8Re1LCgm7ooMwE60yZODl0rOtyQHqcJVu7b333pZfhSicH
5DHBhoO0eSKPQ82e9HxLPWFr5YXzXAHLldaMpD3bcdiSa/TotmFiFV+K3XyIQJV/
b5vo2nOj5dmgNdYOrphxutwZP1aTEh7MdaL98L5zi+mAgEKZ3K6e7TgqQuus77tx
IH9rHIK9txfFlKSuMwSU8ZsQ7+Es+B1Wwrbvt8LmPoNwlzsbSCdy5M6WII344gBg
bXvHKR4ISjc8NdA0jUBDKXsZummPzaEHn70V34MuBpg3mKT5gpi9ZWxnsWnGHoy1
U43+VYcXKf3xgZIq2+USW4+jDdjMKhlGGXOzuIu+zDWrEUwK0o2kfx71OHkdzAOh
iCwZ4+5dzMX11psHfwhSUjUOjRAelM2BuAo0AvahO2qse/gJ3VPTRNhfDtLmNo2t
VkxoHe3+p72OhoUDkG+c4DxbZQlLNWb/g1H/kSKJZFw5dNGaUkm3MZc4y/adXopE
lrEJ0dZ34GqIqA/3DWImTQ/ZRQ0+T/Prk6CPAAeK/EOBYheZuNdY0jJX5FcJ0A7u
akcgBG6XpAAKBKpufhgWxy2NVBOaW2QpZ7+lnv9fzYvPCp08YcsRUnHfukgpf5hb
HUHb+kmhl9IFBLr/rwPaSx58HjxDFu+91TCMk4/6XWcmUhcP+Ft972YOVX/1ehF9
W/mM/HW+wCA64J/2xbCbp7LmRxCQ+tLHqFsU530cWOixTyD862x+uRpHUctcWFpa
m8kJzVeknk6Is1f6V1jCa8frFOZrhjr1MbRsnL+OOe9slpxMhfxYYNgngnDbFEug
WqkQiO7o8TKD2k6SaqU2X7HFaHq/wH4y2JSWgESxax5NEytW8zNRdm389pz5zEOO
yq0oDKkml21jC622+opGI9wW6qGM1ZKna4astP1hy0nT0MWtwhGZtEi0gmZJyWrB
zAqKgXSpvDn4V9dWxzqdUh6rxgG+uvjPnO7nVQNY4L0RPqEtL3Mr481DMk0EkKA3
K37AACO7OWBVRuD0HGyBWEW/DEIxe4DsbYfP2Gx4lHG8rFV8LbEMzmE/CKmzOFzD
ySF++LxfE0hdt8WwRK9yBdFx/rq4ldpGhUe/KkUUCz/ZF1CV/vPhYgi6l00GME8g
LWcZTr0aVxizJJd+B9pH/DeX3FZqVEK4b+RFqkdqJiEc0CxPwFl7/izBJzJstoP3
mgJUTuFg272VoFVbAHsmqiZg1oHbXCmA8chEDN8JoePQ4S/ZXeEijJjRT0+e5c/M
Y0LDIIofTJtVg2LT18mVwGwpdQJUexirsbBSEn2Xigx4ETnVQ1tL2GKXhC+oPEIN
7RIey4+gY4GgHh9Pj13sonVPib+kBRE5CBV+3EwNtzrL67yJNcb1Rz0qdbQ0Bqmu
HhYFWlARfFje2F2RELKFlRb2Zz/M40qWufmLR+Diu6LmcKKQGXFuAENYaH1RzEU7
beciWQKz4XfepCuoLa+nuQHqym88iU1JWEF7giUA6bvEGYhcaYK/11iCDThvnuQL
PDSw0nQJXfcYj4ExKXfIq5YiyG3WalJ1HweYdj0jobetBnohnrF8AryC7Qyna1VQ
DrOwWL1zvJnek62eqEew8BeqF+KtFchleZjUvlHnKf0+1Ux8fUdK5yw+HesEDHZQ
a9Wri1CaZO2M7GoJcnLiv5SdtWZNaXkU2juiivSJaQZNU1COFtA0/u8IHRHOZV37
c1y55Ob1WUJG2YPup/hAoWniwRrVXeK00J0llnT+Cq3QuJ4wFnREJntaUcjWxZMh
WIqaDOg6uv280E5gvjQWAQ5nY6u7gA3H8ZkOnpLtNT14kEN/GwkJS6oyAJAWSEx6
cADi1jaOR/GxKsu2TXWKOfFK3hi/i5Q6nGqUm07EIsqjydaWnmcHAHXJ2Lyc6P8+
7gtyJG39DNOtpWOEpgO782kHJN5BzsW8QwMBtSL1tnO7sCMJ3ou6iO2xii6+N5OP
RXyd6kgbt4h7VXS6vZXlegwYH8/sCli0IfdDP3i6Hv3eBfeLZF8myL8+9n5kluYL
3mNlTU1VOA+C6H6SbQaXXU13dhrrOZ3KQNnlHigFYBCkif/bfwTmTGYKiVDMRSlC
G6lvIYKEMEptM2HbWlgDcxgJyxTELoxeiGPuDDr9DLMZ1yAlLtgvkHmTbK6/UZMj
jaKX6Zr1BoV4LbEIZinvVF07wpjqhYeh21e3kvSBgNrcPr5cbmwjgLOo6vMgNFBj
2sjCw8+hfHShCwr0KWzb/+YS3+jdyi3C8Wf82+mtn5Ftm6bHwsRxc/Q+Pt1uSIMN
oatmMNV0MGkG9h+0trLOnvcCVSm6zcm7Rh1ZEZKj87HkNTpvdn7zp1jWd7K497Dy
UAnfKSH2hRyyGLfAek+gayU0ZHb1hO/zon7wSMPv/WbaXq2IzdXd3BDHBAFXM877
ikqKQLQP4+gMegu5vN4NtLQllJ3xLPy+KriBL71ZL9w1i6uk+vDLyejL0vgtANO1
ZcrbnD2Zt0+XpaitGIHsxA4WSRdPusEU0XcgKDW+ryhBnlpKJnuFTYBbbXLD0okg
ADU2Swl2Ls1GENJqGOnOopqWb5uS4wSdmyb0w8X6Syr/rK6lsBJNMj0OpBXoDAmb
UKLFAavAJ8uJpHSgV/jzU6rf6qL37ak28C9RqkVUwqZRvTm06aEPJEAVyoar0JsZ
lV0kpJODWJZNhK9Iz3/i+yb3gdms+hJQz+W38njKaiABt6KQdtGFjQWpSqp5GEUm
Y8QJTw5WNl2d5peSA/8nKdgIOs2v6d9VwHv+j9z5Zy/g6rO3cUN6uM+FTHFkO5zW
L6vJwZm7N3l2C7lxSPnEQhHsbtKoComWUFKFUwWT5CBUpBeRiReEAsWAYIvgDCtJ
ww6ZF4O4akWtlLVow6sB0KuRzJ+kOSIqSgUmn+085Xd0AjLEDRiLrvEI5TVfKmqh
NANyODRDOomkx2mt+2qeQgTIfS4+meJJjBPofeTZ0aapEeXQXoYhJUDczqriaEgD
Kz79C26kJysN1Ctdx8o9J+a7+Z1GLNoQPd6wQfvueaLkvRgYgvTnr5o0Nqq+eeHP
hK0qSb/B8cz6kwo35qeYCnX9tsm/ju9L8h2A4jQ+1qq/D0RWvepsCetxSnkrQcto
LUBB/zC0IxCqDQfRd1TWgjh0MfGS7GF/Mkq4qJd2sDJM8AIVloxHNRvqiwMikRJc
pqjEkIqmVL8qzzLfPMokOyAQ63VL5j96SSIKHizaI/zrsaGoi5amriC/4KUuqLIN
bj5/mLDHLwQ1cnGE9xRHodCbn6kIT7cPJqtcD2d4hJVvnPKEpgVE/Fmtpg6SSSRy
sVOhaLsAoM79LSn5ae//ELBc7Ws8rmiEkHYxIfrDjRLROZFVhlwd6b6xOlRZwmqx
nwPc7QLpe6m1B0qsaMhc9HnYoPEIkMVwmrRhVWTH6Hu/9bG1fV6Xn22/v7C/Q4ow
BDNn95N/G86GXMRNMw2TWfBlmeUovRqVwUo2QncK6nRcrUubhGh7GnTvziqv4Q3h
YyWDpz/XR3tDCaunN3nJbXyxiG0NunJwWSofbTpdr4mGN+OHdv1o94PmafKbv+cF
Z1HE6A4z0MYEfAWJ2Z6fJI4SD7RuMaA/RO6bLe8YMX5XJgxJZk5ljW+ZS8zOefK2
7FN2gGfNsWM3x4z3PSTlFccdJzTOG+pVPi1/4KC0BfKddIa4Mmeo0j/zL1WOFDIy
IrKyus+3NxC0TxlCjtZ0r8vxzgCE2bPGvYjnrUXEouScCA+KCLwVt5jJfUTjYk16
PhGvdQWYwXVrx2kpywhvrNKnTMy9LGsjcIsBqOxPfLNM8Xl99+m3jJOuJ9xEL2iR
b8NnYrZ2xFhvr9MKHAL4DcTgfDuISmbOPhd1Hl9zTtc3YPXQNbuVwJQNsLXf2WTy
xDTY1xcElCkimcAH6je7R14bGhp1oS3bJjo7FpcpXcj6elAgle/boGlHwQEnnzhA
/Jt1cVth42j74MW9gEsbEAfNCWKfwouGPLnLfR6euZ0prya7nXB68xMJ66j418Wc
4qc+nZktHIZf1Hd1SfpEqJLBsLBxAiXJoHbTwyy3hPIqpXmHY3SCoPZ1sbrTLl34
zYXQWT5qMh0HhSjeCAKsuE8jhEjIsBgIyg4Wc94PyopbjL+CZ5fQGF0sYT94Nwvn
vw0b2qrqA4jlmsJ1+sXVFHk/EQFLoILCK80BVNoH6qJyyJTCKqPIT5N9Z9RKTNsM
8dXAoNM3/sJ70SlF1wQA0VA4ng3XPGgOyh/yotGXdW1MO0AisEIgSEMvPQQ4+wGQ
TpxG7cIzELNuBB1TFBX4mSV3LQ9ZLi8z8p8rdT6VkePWkCngDOIk/9yCaT6+ZWgG
ahtz5E4dz56cLFTP1QZZ+QUISxvbK8qt97cc8lhlyXCd7Gct3slFwb92JVP4Rt3j
B/qdJceRDj3/dKnvobWJXaldhLqmxwp6DN0PhvtpBTV/90QziTG4zk0TpGs5W7tj
9pcM9XbN4nBabUvZHkaLnBkLWkwO0h6dGwQoqwSeyEMWyjHesvpLoT+pLX086KBi
hsCqBxL+9PeM8HeVc+E3Bb16ZGBHltZdxjxpms9MarFh5NJ9ROfRQPDYIkgdBeJh
MZcfMb1oWmrEVDq132M903q00KCCcSr2HMUL1DITjlTZ99DtG1WHG1kZTqs92bXf
zt78v2Rox5KPDofLwqpsAHuVkXbFansYhDCqjh83uzWM+Dn7y/iFiERk/bQu+JMb
XoMCcWUdisNK5+45Cb/zaxU1yVhuQLdjU4+zx8FOei9y50g2aGcaF6O+n7JFQ3YB
gFmz6KYWc1zlC69wU12JdY05SmFtBvGi/HPAvz7c+CY2bLkEzAY/eTTYSzQSftts
+0zYxr2HBY182fBINFf4+trmW4GEexDNIh6+2hwwyvGrwBk3Fma7Ty75BfdPgcB1
R9gXRwvI0jOYMhPIcCV/z8z9cHnLyfW10ElZQQcAeYJGbjln9+IVUxfxmYTmxN07
jdaahN2mamfWbydQXfU/e4/BOa3/9ULrQSlCDqQ/D6BcxmKQG3tHeVXOEIBciCuN
ITRbpS3iOp829uW2sNBH75nggtnM0278Q1+jOwWzzT8Sr5D7ZkGVVUAA3E34jbT0
vHNA2UMPe7QNBK7iMEnLCwxvbNjcUdYbQxPAlOkoG7/4/u6b8mJLRcmYLaTpdtVW
prSSkW+70WSkcICxoezRpimTEns4P/HcB1tHaQYONVG0l4Iwg4wK0F46hfpiKJi7
njiwuX5Yigv4bdft//WdrSpNi3Wllcxr5mNmeGRu8T4L3inSjBZ3E0MnmGXcZT3o
G7ZDbDaOQZXY8Xhm+v9PTq4x4Sycweac6QnGfO5Z4I4lftaAb6qRep103RhPpAve
VQbbT1JhLPSxA4mQDJgCabyRQzRfaXyr+1dFxvrjuthIFiSbbqsN8gF4XbAQIG54
d2caMuMrMp/RIGSim2VipuBJ6iY/TQGGbC+IdTBVa9Aw8W7tgk5VLBeDPDi8IE2g
3bzuPKT/m/93DFlWUiQzAt1B75ZeuCRoHT1DUkHDqF1GA6Jec9tTe7wqMMN5s8yo
ZTNygxo443KSQn9svMk0wcjLGdkOBm1O0vmNRohD770XP2sHrs541LGtJezgMD3M
nzlH4zOORN+OUeQy1Tw72v3s/5vyCaUG9/sbPSosEqkAiIYALlgR1ejIrmbaxqGC
IwQ3Ora2rJMLZdeIaK/nNTIASRV/IQWfybWh9rXStMFo8J/6ynQK+3ctbVdcGW/S
a9cbScWBtBoJiaaKzH1ER06LXnMvaU99Rf1Z/LK4QdQurskPqVRFjXnq9e6/eJbV
Xwkrsusu3MIVS5eVCW8J9JLzGQqXN3XJ55J0hs8d0qrc5IlA3Q6MKgvmM+aCEmxp
js0eXICvrhJGpteaSwIlENvZqdk3HodJ/c48PiFdEPK7Wj8AyopSA0wHF4Mkswpt
Dx5I+zG2x2cGcqspKICiG6ujuIdQem9y+hSntfPOV1N0Xm5KEMTOZoFDqfMrCJSk
zCpkXF9SbzHjqFfHk7mpqV448I6XbZWNAOfqPKpjn85JDMcahb0vb9pvfofgAmFS
URUYT3wdS4XmDQGSIiEuOFWc2jNLMueLrBSS1pVihP++sF28qhaYwkT0Ey9iLqpm
pwdSMp9nNJsbxC+94oEuj/GltSTV0x08lvM/d4ew1Huzkbg+I0B1PD5Rmp+bjQt1
xVReB4FuOggh1wzO4vRvP8PBtyT153O7wVnFEzSaVin6GSeoPsl6NQW5mQWUgCNc
LTuzm7OjDebqMs8965fyhufhUmlUFYktjEDB5HgrLeskEgbsm5dConB0B14PmIGW
wTV7+LkSZWMDELv/3tup0Pffy6oiBfS0hM7s3OTcVaqLE7rFANmSd8Q+zdJh1wuU
nq8ynamWiIPPDSKvDDZ7/Z1HggRfDT/g7kRT3tFBA3ozoln5u0+CGkbjEqdgroGj
clh+xGqUt8STBvbhahRfn/+npEtUOri9PA39B/t2ND7dzqS7/v6aXlmzOMZL0rNV
h28WSFFe+ZbntvSN7zl8wFgsC+2nF1/lY9hLvJRxYEQZOH2hqH2I9SnfxdC6U5Ox
+3C9mnlyd27DqPyHaQ22uiOVCqS9cIV8u94YDWrfFy5DrHyh2Yr4MgHYs4OqiHgi
qtmYLOxkuNLt5OcffbbF0Baun2WOap4QeaGFVR/PdaLBp4+hFc57bM3/oH0o1Ewo
um4UBjTPmV3vXUo41E/DRuGesgod+47tjn73H89oIGn0WbdWfRlmIt+M2fLD5Oyr
Qyg3X0xHPK24EhehOgiLqoJutPghtMVDfYvzho7ha5+CUscGzxtXEz+JFPcTvDY3
/IZ0OFKW+2fdN0wTiweIcqK1kRJ/jk0DUe9oIPqthUaIqXwRTw9EoS4FcKdxZaZ1
NG/s9s67bomgsMlcZL8gw5MQNRuFwzeQBWYHTfCVlVl0SpAB3eLB95M+FxrjhGDk
m9Gzjc2z3mXKQHvFGz0cgC5nh5iHnfaiEZWMx6n/8m1WcNKJd2/YK7tG+Lm3+qp1
hd4vfY0pnwE/xj2/BnpWroWRKImu6nGQRWi1qHp7h5cQSDRLeF/FRXte20peK/Cz
nz2Hfp33Mg7rZU8TpHVhlJUV21Wm69ZTDW1wanjWfTO9JI26wZ1Jotz4eM5mss3c
ltXqo2v17ZMNBrixND0Y8OdsDFcvEAfGuYjrlB8huxR+qrpu/wWUang/mJz4Yj0w
LXW/7c3qe7nw84mlBlhjHxO74q7YoOz+WXywwFS18VtuvtEp7xf6cxNrgY2PvtJ7
R7e69YnUouFVkU0l5hYz7CWpz8eSrSdinPAA7j+Fnl7maw7hq2731oU1FtaLQNNq
VDpWyUw292EWlCX4Vne/ziCqPEpQDPqT2MBK3di+f0Yw3UhBx3Q6vWDAROhUiJxa
/yZdAcvQrvtaIjGUkEu3je8zL4l2jPhQuiQ4lgpD4rx9tDfMYCpuUGRrF9bYvI6F
mPB8g2UrjYwI7Bjy4K008rY/s2Ny18FWSNFN1FdKKOy26dxrOEuxDjwvBHdf77hH
uXTQ89YZPqo/GLU9klli3/68GjysWopugUt6T4vCqaytAqTVTaQL4KS3ZJfFRKBI
lur4ZonxLG9LonZqoPIQVGmLUKtkqxa6lw8Hy1jcGrKkeaAHmgU0gxevTH5Q1vIK
O4i+1UFpHP8RC05EP54AvoxcgUpNIhKCZg58/SyR6fpKU2PJ1vVMUtmnIav7jg03
vn3nMr7IYsp8F/+PkHhlNZiA8+VeH0//pYxkPHwq50tdbcURNLYD7Zx0KOA+JAKJ
w1eExQVu125rzYXvNv0KFuKCmMl+hyJVbfaxG8E8XV0rX+076mTm5GQmh3mbm9u/
NsPrTSQSSZxgW8mgVMvXGloT/NMUlUlHJDCRMnoRCo+BCtbpYFyCKuMauvO1NJzS
pK9Qhzr6tLqe3aHfhuPUAYka5ipVPWeU8HFaFSj2iMeMWVVGPcA6dBlBOpts0w4+
brXfGbabrwrzaiBvoC0u3Zx2EzgXUdOvCYxU1mBBA8fsb09ZCgaAOfeuMjQpl/VJ
adZuihz9WUY8mTIPYosh6x0N9LSq7kPD3V5sT/5cL7C8DifIGNqErbl2uUAhiqnI
1dmP3GFP3I9Vi3MFSoGEgbiLoXoibzG2fPUv2VfUyU675eaA2p2i7Hmg3FRMQc3f
cf9/ErZpzHhgdyZJBjRaxl+Aure75NlMe2+6xPoAWEL7Rp9whwkDjdNU/mtwaAhR
povAhHL2OFbYkQcAMtLJBlWSAO13bzG/deTrakAYYd3gfK9H5devkgltX52GPX88
wNfDec8GNKkbkb5yKCTMS+FEBorSOcdveR4sYH18OTx+XniLcrFPwGlumDcZW9lx
zYM5fnByCw4ELE/b5BcNN5RXG4bV02Je9HaC7/UxLg67oKU4mgm1S7gAyNdjWbHb
S1GMW44HadhVjWi8z/4uZi60V9mjIqhHhMQf7CRWeW2FJ578KD+IIbnGPeUbKq9y
TKbXVmiUBqMwGOwUXRCNabV5P2EAGNlwbZ0zUVCdH8XFfXiDCt/EOQlrbh6w3BYR
MhmXXIgmTsptGvbGI15D8+OMqMGsBRJp5fGOoGj8H8h+Wm6q9zsB2DJ6ZchFnS7q
tLITkJOE/oT1qFSJ05ubm4X+dRV4ksiJO5kUUJ8vllmORdc5xyiOu4u+cJSmuW07
pkqgRq0fNLvz2iontIGM0mt3qoDAkXmDI10Ixxr3c+cEip6cJGYRr2JquuOgR/Uk
e62vAyePJkc83vsE9CnUDg5eVn6R86H0JSlaQVW9Yb8//UBiCqf9N1FsTafyKD2i
fnvoiWyKZwlgqnaIrJgOLiHwQUJPRglBZjfAzJEsw7HZzaSDTKVHRZ3539+FkrCP
LftwEMvpyIlT36QyvJT51MzWpK0cPQDKwvEdTccUy2j1x5CF3lyW78mSnULG9weX
eZGbAbjZwFJSauKYXaqafzQDOerv2DxPiTtTopMiiI7WZYssWS6wxZZIzROtebMl
C4SVQEXSCOW9lZqy5My0MbLX3V8ZyFJIIxYmZk0yQZqiTk4B7kuyjJbOBf21XwHj
Btqoa2We4lqrX3w7SpyepLb2hXtjkR9qdj7+QPjdnUGCp1LWNtBTBCYrdTJicsqu
ag3N3uXP+tCktArr+JCkdj58nupuL0Sm3nsY3Dg9D3JwxfXSJpbrfLPWTmbxlo+x
QKMbLFfBFG+P+Vmd4gszcseoSZ6/mtIHQM0PV8MyUb6+qRmiku1MdskajgkUmavC
wyQ0FJ0yUGgck9iaWM8n5FqrAjski6sYMbvehmg4GkRMj76pMh1ADSEdgzD/aIb4
KA5T3+cwb2rwY37Q5BoYibLAM3qgFHgiKeIHCXtAUHaT6YBjah3Te0Z5u6/YDX7d
1p2rfd612uodjBc39WhslyWegCy1Xl+4NI/lw6VT+F7Di7mY1bbQpCVyRYhU8KsU
/+5k0yd3wu9R3SLsY2i5OPg8qScBwimlsYgW6pPr807qpqnIy9+BpeY4NGagfwRD
udeBf9y0Zek94MoImmXw9XnKCUik/o8szs8MBXvPu1Z3MIvUui6mDzg/dHOCcTkG
LLbztGRSyGmaV8GEZ4znTuuy/llZqUXM4zsmXD30a29rYzHS4T1Y2GMdfVn5M5KN
Oa+wUjHdfuVpmZ195uEXXB8prXSSqs9n1iHOwngpG07gYP3JQ+uOHSStq8WUGyVW
sT8qkS3y540dFBjPlsi2vn2gUixjHTN5EzIJnYUAoBe1/fSu8lQAJ+2W9yf9awe5
5vBYA0si5FwjYBpdwMnqUbhrZrr4XDQyqqLbJ+uqHY5VrOkF69Q2MToWulOmmPtX
HzsFdzYU3TDuqs8TqfvaXqPChDlDPyPFNZUgkkHdEK/8pBXshn1SHym+2N0YPZnG
/OPJpy0iIV/V7454f0kIRNol6942Q1v1a7iIg1aD1F16fvlV0sROmnFvC3HPAyNO
XH77je3GkiuUwH8ivNdCRZ3rWRNu9Rnayt7AyeokPOoetfew1HPlGZgrskgQ+o6Q
oIDvXaCzTLBluzvJrLIj51l9ngq2lQbIFJTcLq1lJHnHWjBcMw27D/dX92lVptHN
KNJ5ObmDd8aWu03LXh3USPAI/7SONbaJU/fsVcHT16W6S5496/NU4iVA2kGT9Qih
whbhFCeO7Ob2ax37Ozd8b7KkBd8F6D4t6MdWrAI6IYejSbvtrRMJs5gQBW15gqyL
eHj81ZEEB5m1wE5PF4tojkdVe8xBJTLZu/u4XnZPXRG6hDdWxTSQn3r4yQSagqjx
+HcWk0yL42k1eI/hYwEwi7n/UvcFYChRwkVqiqr7wcc+QwHlPdUL+VZqRZGpnpsx
BX9q5b5iLJJLbyRLnQzqTAdYC+lejUM7fl8NGKwCYZR4jZSh2MiBLLj/hqTawFJI
GZztjLTsjJmZuinwSvwtG6i3Zncy8+3flFsdlcyePbQSm6bqZ4v8KEBu/BTedpyr
m2GbH00ZrgtP8LprIcgjoNwYaq6MO4SWyhoaR5Fy1iTVk1hb7hy3vT8kYm4yZQ/O
D5ogMKjg2eV5CYSH/zbyCWiEe/FacOUIbMWnbDAR5jtakz5uOK7JXsJbnVo0DluX
Tqno27wBRN1xHw09Yo9XHJk13BlafNvS1bLSrSrU/rUa7eWRbUkNNuxD8jJ1iwjn
W1ihk6nwV+HB4DInxWyVOhg0rIx8rf4qoWf/0tJs1Q9wuXBFigdJOKf7SLdC9YBg
VGgJyBWDdGCgAITjj63LF9k7T0D/mPq3l+JUtjiXX80jgyyX6q5zcBiMkim2PvVp
xZ3h4P3ALrhqaw54MD22jPMrj49uWC+nEtOICVamyfpqc3qcVZyfJAfDdEbUZJGJ
nzyiSyLzTE/dvAvmXgyLH0VBIQCFOXx6kDrprv9ogu3Blj2fIts5jP+v7ZqbrY9O
ZRcLi6MG4+RqufBZy9xpgJtvD+AXia99zsSaV1uDupY1bPv9s9IRxO/+VJ31vgX4
NSmTFeAZU1hJu4J2Ujs6Aum521HncCXSGzTLAh115fAje/xwQMC16oOewgjgCgL8
xBk3qPKtHcEjkqQiJG/zAeaxNeor9RMHBHNWW6yjB5r5ZloNVJ5d3PpM+7KOFuP/
XLQ5Fs7N8PToYwyTWjvUb2gqqXLT9NvGqKuvsmHcl6LTJErGy+7F5X6obuJI2O1+
9kjnTHgoMVGVgHhpfq8KX3CTkolZTzGb/WWal/aHmhnjaTwx/exFNGCOLCNYK62t
7SKS/DWBAnCFU0Uh9XoVdrnZcCjF8ScXJjVoEirJacz7NTfps91ojYgfLaAwrsTD
YBY0O4UM3PLP79af06a1edXt7welGKpGCczXskg0QGwUbYc5Tnv0fNUkpPBYubSS
YXrSQQr/z9wwRj56NFQCIIsEQqS2r4lxRnOYPC+jDxbCkZpeC2QIvd3nVjq9qyg4
dUEuEon9yZcgZb+avYq1kwgg+WMr4VOe0NvVUL8pInE9mwR26XR46xQdxGe1Q5UO
CQL1zsBG3JEd2/OskowjECah8XtJE6V3bcxEhhxMEpZFphBRtb1mgGnsWJbgdDH5
oqFYDQ1Kd7llTcKnqaSPQ692F0hm2PqGXCtAoaqH4iZ0vVBC0IYzUyUne7v+YWVY
NVtjXwBsLSAUx3QwjuxHGQzz6oOi6xleT5v47Ej+NHg0NzRCiWUk3r6cu3Lg2b+a
PvucudS8p/7n3zDZfOcibXgu4rBzrHFrNT+5Vdoh4yCHzXUBPetzJWpdgpd0yVIe
2ukxImDQppXkKszcKa0YY3Ov4OwFNJdUJA/V+wp0gd3ZEpHN4tXwdsXEzZsanq9u
dDM1QttF53M5VdmCRY4JOO8DFomCXyHEKYaOEmQ139ItyaQThy0V2MHjkuNd34fw
71ZNYzasAQx5OZusm1a7HpG2cx7SinH9pYgxM8MgihumKG/v2ry4jJQA8a37/L8w
IuOosiRWY/tpuC9Lyl5cLHB3qvwJsGbQF41C+Y85SOqyNhnfYcsO5Q9DTLorRVaL
ZXw/Wbty/l3PCgLdmmT9vJDUI5cAzddtbYR5O7J8uNNElHlCH93DSMKCyqZhkwsM
D5IPTyX0UhCK17N7hRDZvD+7tnbccV+2u47F9DMnmrNFqnRXohPswF9t0+Rw7yY6
qEC6CcJq0myAxIWN8M/KJbH31Fa9B6AyAsy4TJYYPvUpf59BYN0b/+ijiAb99eqq
pfilmNAa1YWmI/WsJZmHRACgLB3r1MOZGlrpWWrLg9qFM5ladepZ8xBDhHm4u2H5
Eg+Mv801KiZrZl/w3vnNlhNb8TaStVVzzlqwamkokMzUh2W+ppWmiqnrZGWQHWE+
oc+y0OAe8SrNHXtZYFhCpdAuAPhw6y28lkmTmmuHF5KpJWtsKib8vADRk57wV/hB
D0+tg8OpIkF4+CdN46lZjSkVwf6p7fGspoPf7PV/Ay0R071zJjKxlHuYEMYSug+x
wsMLGUNyguvZ7lwIjMGwJW+dfYP426ag7U37NsYNe0APAlRAD0b2Qm+gKHC5DrWu
IX7mIkADkqG0PJUtONSNTzHY+OlFJ1dmJAzp4rm+fiFjkgprTePMdI9iZOsxUNes
11bs9UL5k4P/suHzIVUsJdaOFpMT2SBRFNigm9I9nuSup2yzra2smZMJVbKAyhtC
kZQSKKFoEbKFHfIZIP+6g96kVQ43/MpO/cO6DJAoqoj6G0q5ohibXUuDLC2CSBtY
RAj5fy5YurO8cooguUqfYh6rfM4wiY/gYptDSsSdV7GigRYPBckSILp8gzqj/nh/
VtH38zM2IF/b2ZyW+ISxO0qcTaak0rOMzE4V3magKB0vBkM9mo/JoGsY6PtaQnbP
kx2CevwR3aVQlaEWClYYlkyyUpNaMDm9IOI+BHS5IQJvRrssD9Wksfb7jl98RPUA
aGIZc8GosWKC1FkMZQeDOA7vd7KKPZx1xGGYcyL1YDxWHNTbxPuPjBu3WST3tRz2
mEbRp1tXBlMXNkXmV80LkjjMNmAvN5TG0ULDUsYUSG+ywcrTzsMpzMfBFid8OLdw
Y/s5O7OBl6JqEpj6Y555yfDFAAkn5KvtGvJQUv9PlV3+n3Jbpndi1FOrWR8beZou
sZj77gbacBQl/1HF98R3qdHqCJvBUKap4SvAkX+kyEstvD4WjRBGteAcvYF3TZI+
+sn7aR9FvSUOMM1IXtDPQlDKC6OLVLN8e933ypB7FFtADi5AHXD2B04DLG05p+dX
qed8W/PSZBqKuLIdopK5Ip4igJgGKS2hwjMzbtIkOsiWbiUT1djYbV7zBC2rWpSd
y2V2B8xRorOK4S294zXnNZ1etUk9sz42fhD05sD4Z2bWDc/UdimtTkVjTKRnD6tK
1sPwsBwDsWbvWo9IoVlOi9y6EHm8F7r+k3kDOCguh5VWgcmrNHcRO/byeWn/mViq
nu4F+F003HJHEpC8nx0UAhyJ3xRNNYqWnTVbFf6WTkwinU4wpVKDmssflWP3Lqc/
p2UVbikwc+TlJIpSecnXWyouKP5HFl1LFTyOOgzJhnM2EjnUdEzy2biuzQbxG10f
G0Svui6nZb8uWof1psDny8ph7ZhKTf2SH3bXh0rkZ5aEb1twqf9JdLmMKLPV4hzx
VYXHG1trbnNW6JC6mbItM8jZuVWhTJsDKP2bNwxsoVt/zYql13aAcZ0/4JlmmigM
UDQYtUmlcLO2t/VMmpT2Ns2guXgFqu7FM7om8JfwJg/e1EOmh4pYr9VNZ8mxs9n9
Z5VgWs+qSBp+XGit3emRP5bR4gctMGMP5gJWrYtXQmtghzRrWXkB+mhFajcDawtk
SLd8NDU+ctRgHEQUHUDpVd6HbHo5RZ03cg0AB+txeCptySog9hsgdjWRjTRu6DWi
ZzT9p/P6LTn37M12SWyipu0OTdTJfYiWXL+oyRjC/yg7bcgtzkEJAQzI7FjNNXSO
9SlgpdLMKkg7QdiZTRSDc6uQMt2XbvCjxBzdew3b2E531Y849mx2BL9gUMV6PoSP
m9MozzRN9QiR3YaglIKHH/lE3V8THlfBTul37e51qyp8MCz1ZpLofXP7ltie3bL8
h5TP3Sxga6sVrEje4aZcdL9XHXG3kBjmjtw5V2gtwofuG5grMPs6gc5be2YqayDp
e3xDw5w55Da6zypUdzWgzVEMezUPfadbvGW9/ei+OsteJ9Bw7q1Xm3jnog7Qt1FI
n8/7UJHV4g2JtyPvEz0l41QwhPAFHxA+8tCfOITa6/lqh6e9ROo9Fx7tkyinN4jX
S4V+hxD0cl69ZhLf4FNKpNigwdATUDAHqYE30D2MTXIXWyCigyHfd1txZyBndlAF
41L2U41wxj+2cRUQOQVu0HtySbGQaGqhX/eC5IUyAqVSTJc3TNaRRmrPU7yOL4Gb
S3LwIqcC3Vq+hRJiIC4HHNoca0C6SMJGTbWNaGDzAeWD3iJTJRR3VAm/T8R8nBQn
QRij1FIzO3WU2zhA/1WnYTd/a27KVNgZsOT7mVnNaefoFsqic/LUw0opg5JPfme6
VEjKE050mSMOdnlw7NNVOhdmae21msCodAfWCO4HgWZbF57PpA/fTZxOL0Q11hOQ
ly0zKkKDTMJ4BqAGfaO28ctuRz+ukk0i91LXYBP6wli9uKMmJ/RcMDgoT4g72Tw3
RTTIMUoLNlMfiQIGI6pDUhknGc2BYqMETkAf94fbIOHMFRa52VHkjsHydWbGCdiU
PQC6cGDZDrscrF+sRn4qxy7ar9Mmgnl7vj1CtRJTNjYlBJLsQH4UvyrXV8a0yN15
I34t6Yn/YxNQjyrO6mpBIUHRml1+2E2+CCqFPJeSdw9adjNxb1F6qVyiVMfjRlZm
eJ/yz1ZT4986N6r7a2J2X5i5m4QyYGoNqv9EydVQtEdFp7buvELyrYMohsaWdE23
wDRdZ/IxTgmYNBBlTla3JJSj3YMNbN+lSWD9Jev6GpVz41B7aKPwU1kHydJvntV5
n2BAOR/wf4x6dzBPH+kGiFuBg1FdO0Hp/mC4V5POuVejw8RtkYY8nYVBfhlGtKtW
/HTcWbl+uZJkkZZVwo8BzUDUJTnHegQxq/Y85d9GjctA0PnREikTchnB67/MjG/V
DlEOFi+Kn1jyAnsb3NbPgYNpdSh+gyVwzwActupbtI2KES/DbrJZLsV9d7AMBMoV
pNqpGE5dM3sV40imgCEOVei4LE/z/4Wzv2C4w66QYxkTSHkrIzoDm9hXhETOWbxH
/iIUt3K7oz/2GMGh140p8995OyDB+JVGJwNXG5sJmd0O7lF4afBhECu31GNamh0b
nTllCPoxcQOP0u5CZhAX9O7xV0WgUKkTH8LnRQ+kL+iakINqtpkUaYNEYr80wJi9
45Ix8pmTKuja9PcBFvS5ASXm+sMO+4s83lju9mgcA+M0OENa+G8+hXct6NFGu40E
WqcUiLYcUIxt1y6L+EXfpX0zXlT+MRqNdya22kNkwovfKK5uZTJH/ZsWI65O6u0+
F/+t4JxX6yNggKV1qw6YzRD7BNnzRJ99FydgWZMzTkUVW72+pvMLQ10WQcJfpjJH
pqnmcaSmOyjRs4gxQe/ZVdq5v2kO142xA7y4P48/BrzxaA/BmjUZusIo7bGE8wem
qknQnSGwjSbO6O5SUOdnYJizbIVz3T8cbzugWvm1mq34YU03/wfPrfI+aooIZ2fL
KQ8i67BtMiOSHG8paUH2qJ0eZ6z88emFbW+d/gRDekgvN2yJ+aptRIFw41/cqLty
wGj0E5vR31FjwZcLZYXj1/E79NCq60QtqfpKUrcl9X2mE8AyzOCgEevmu+nxX2HS
78IqHdEeMgGjawXcF0ULLEniVb6J8g98tyFO+FNd/bRRsrZCuGSiQG0cC6X/Slkd
4dTu61MRuAdeo9Fwxmr12/rapY4BRY/szc4H4N9KxRQfbuoVPfvRV4cFdNAaYTAM
zHeejeCs/vlMOP5cmJNePUarBZEwhdYmCnHf8apLpU5S3Bx+Ik1PtOc22XqK2gaK
uuHE/m2Qn1ovUGs1Nk12T8I1cTCmgjREc8xO9e+tz08jzMnzsRXJ5FrCLAv8Tk6u
2i5i1q7u2cITWRUrkXQ0P7he6nnV+OAhyxVUEuQ6GP4zJTUBd6sxkAffWDACCCcF
DgmQ1CESqLpFhq8BHsdO3RLl9gAa1D7yLTPDdlOpsDwNi01ssAfo3Et9HAfJWlv8
tvqyYx2kMWoP/mQpAQCAYHblYqHibu9vTx/Tin3j6e2hxugROzC905xufleEIDOr
b4S/Kt9EyvPZB3h97FCm0+z6t3MapI8zPEwsKLzxWGAvm/spLlm7XLNRuv/kysh1
fQA9Sr7XOWNCT38BTzdCzhTfg1ub7lgVtWzCmCHo/HQ/2N9AGtHBB1jrFImwLrYm
SlolHRrErPcv/ekZMX2gDHuWuHppJmz5h0Fa7rC6o1fYWwYQ54WVP2TRgSutoxJ4
qVhsORk962g54sM+HQvASRz+xdASsiiqTkM1ejyR7F9/3PGZTE9pVrezW/cj8NKL
Tol40ReO8PPKO5ODdTRSrjOztVYQioOyR1Yqw9indmZA7aYzDWoaslTDrjWRJhoN
PHZSdzcyP/63FRH++v7qFTYk9P7dOxfA/GcQDe1H3hCbyM1rKeVk3h2MG4rYGesp
/4xGjkLD1pa3VqTcTCn+fIDc2mfKOmzCasKSmPvSxx4hq0eme/4HaSPHnxBt6aAC
Z4CxC+KE7WBmf6s5XrVz4+6ZB+xuZYl+VUSgO6LQQaZN9TV260QklUAEUHkLIfWS
Zay0LbN5baL30fJi/a557NtNnGlqCdDyEq5dkQg6pLtK9MHRnRJ8IHV5DiLvHtnO
TIwTdk6FiffXieVSlPSCuAIJW3MIH4KnACcjWhOQjWpHjG022EbfNABTjzNt+iwY
9o2ZjL+/omC6Jb3b5oFGDJ3cjPxv3iObiz5otBhVet+aDKw3wuk+0Vv6w/uM29L/
QmyywQZ1vr9dJyHi7DSJV+IDvvY0bVkrpgnIkFLohPkpjA/KAm7S95d9d9vrb+ul
iX3SIYkJK2kabG9bFZIO1VFmy2nxL8S6HRwO+Oe/zJstBvWvFwV3iRQxcY4q1WqZ
gc2QkxNuehs8t4nWjk5F66KuylCSWTaO0NGId60Xrq2WCm6BpBIO5zVveBXiwOsi
bT6kZEQlr7rX75r0jRTW1sahqWhk0e8g1Jo7wGB5JTvN30KpxDsH7GMphysReiZ8
USCda9GFB1por3z1vz+MTgKtzXXktwLZmyU4zrqA7vHI3YqQBIk7/cAkKTk2+9Rs
lslLfqZDSLCR0p/ILWFt5MFtD8zTyH/MMhvI5QjWUrA906Ld63DHur5dz2cBMBvr
XlGR1kqVQoSsbZHvREhDRSeMiX/apIPgGXNYspyCNA1V9SOCH/+5DTiuNkRvSECP
OR7+wSHsc9rDx6Kx1QAlbHs9qPPYtH+HwrbGqD1gTR+zFi2R4yyW4NDeTB2cxW/Q
jMaCV3wMSeQdNXI3d/B3mbIZhQKPMGJQRTa8DEdz0tDJB1fz+yy0c0nuBUaUbTVQ
26hwRxZs8g0oM1azPNhFZDqFYtbVnaWf8dcA+Bs51AB9MWaaryyl5cp6oxJzMkfj
jBcmoSrku1mATGbfPlX+orDkW3papg9Rr9rSLbVgPAbKFKJGc7sONBXrHdJSxTTX
1yqOy5IQdqS+c8MS+Kc/iekR2RWiD0Tr6+3YhOu27taj1LESo19o17HYyzZq9JKJ
NmfEHIXC2hDkD1DJp5UMFHE2L05lo9HRWEflTd/tslyEtGo/lxX8lRdOOLiaVwPf
KxxcYrZM1GMl+jYxzUXPM/ihrk0oNwbTH5vOEkkraHEf/sNnDXQLIqjFWnSbiVaR
LTNiBY7J16BwwS03cXqeXfS73zrrpDAtQSlxyTI2aQV/8/g3prisIE5/QaEBwDIY
NWSDC7HlxsVdN+RssEkd5zCIRPpu893g7qCyrIRI0AUi+MsjVhuS2vPbu0u+VknA
UYiwtvwllaY1/dm+Ed3QMD7em7MeR9Xo1Xz82pKBXDLNqF+VtoYmaz7fQ+2ccrNC
gOh8SLwZC41+4yrozt1MmnYhhRXvYW3N5b3i+OAbFfUSG+arztcjLp55CkFy+7k1
rOM9PcFNLS1nO6QvZJ1dN9WYg5ye1ycJ1QLRliLb+e1DHa1qNWdGBSZ9YEY2B0bm
lnbmwrNZgi4n+AUfCGkC4QFu5vmAduxqRyTxU5tt6GangwPNBWx7hwYFHqBa+zfr
mDCovjtOtF3zNgSY9Hipde7nVEDboCSLTzdiO7x0qr28u18zvBJ2kD1TpHDd7Mzv
ntryMAk1Kc088wwH38K26xio3js6ZY1RpLv0KjFjRxJMIu6RJknwNDPHUeY/DHku
7gO2OW6NKMIsVOakPaxgxpq+C3IVq2byZ/j3TCVrZxUhaHvnYijTxyp/Qj+9LMu0
/k28lyMJJj1cNkL7NtkYuUBfzuT3e2Xy7fXPa3G/eeVdXIHHy/OCzoo+qOCSFBOo
kfYyFCsx4mB12OZHc2olTuhhVbU2wr2G274eQoIaqkQCrYhNit2EYmQOnRub5Tal
uOd0GEv99HBzo1pHF2hTl6IhKoF+qlmEjizSB0Ik7o2YfVFsZEJW0BN60PF29skh
Ab1hIgkSe2upY4WlfDlIDxrnRhnR3RkF5cH2l+gWS4pLVc+ITRP1fdhmLb0L8ab3
1zDRmg+auk871rBFXhVyloTX0YchHbzkVMcRJyYTzY7FjzGALnY5gSohS7kvObmS
kitszZ8vs4UosMjars6XTiwpEvBCq2SXexgHD1r8UILMAncNz1sLFZabQ07oZzBh
gKKLq84dEGmFQ+DqPAM9VyLnVIq+JRJ+RLnKuRFDjMT/cQLizpYTX7zGH2AOr2R7
7B1L4z0p9X0O28hlxd/IJB268WiJx3g3nDsnWyKA0xnxPJ5phfwN2nOdba7JSwTa
GF5EJhBvI1BNZhir0WXog2e1ZIxdVSLnsmLgdg9sLTFSz9YQfGAubW6HSMwNlObj
dQZDx4zMYnuxS2Lv+evCVC3+uuuqqtVPx0OoZb+gBreoLEsewJXmVKPk/5arSmhj
tJpwiD09+PYd24gsgNdODuXo9vN1f0J0HoovbcJu04tQMqpaRPYEdokgrGYn43fq
d4ue4lJESg2IuBHt3IeEQs5eRxgmN6VOpLbCk1e1lp7ZlsaE6WD4jFWvhOHBrjNk
N9glUJIB7cNwQjKaqmLUnyT7jxDg+A0L2rKl8E8GZl0E7A9ecEBTXuNJSwbASCSF
P5MNKYn8vauGN4sDGoeCrVxXOAnQgJ9Kfj03KflXUujZszcvG2KtcKPgouO+2ZrP
3pHAz8OPRzvYyFoo3gPMD7NkscEDSeo42bADGENxtG+Wq1jjyCangpdpVAl/2wg/
BcYK0HrpxAiKsGYR1vt2rZTzL3VrzOJXYwbEeGk7Q8ynwLSTOxXpcyRVjxAmG8sF
bHrdxNfpvggs0vSpU5kp1133Yv1d9hPpt/YIqTihsVo7s1r3zPvuCGvKSHHmEPiG
RjoBiqcjWMDY+WLkN8szTH+G/Uh47xMydHVLa7NlO0f7ZuZ2AbzJ61HJtKzLsIg2
YaeVKCR2I+4oO0HtWLHpclPx3du8fLjTVLh3yQslva8tt0LB07PxzOGe2eQIk4e/
eUxdNUvH9XMi5IWjEasCX0azaBoHjA/DvrItdoUL0zMKeeZRPRWy8+a4vh1sT2sp
Gqb1Xafgp50B5ijKAiaBxpNCY4ybOUQQ8E7APs8jwrzIlpBmVdt4Y5+r32qaUE2f
88bFkC5xsB+xUw8LQh5RhX1qzfgkgqWxNR7dyALTP+rHfquDJ8hY/I7YXbVELGZo
/iGikUIah3kCP2Ief0IAB3A82s3pCKY+WNsbIgDRpkCuOhh39AGg3vPb1+8q8qcC
sTx2G47N/0ppXU2Ja3QwJMRUc/ZF26a6aJAgGXahNYlKcNyvGRy7/vv5wwsFNkPr
5atpONx1P5VrYf0mMKKTeA5rxnkTboJmrfUeqa2MtYxKmAIuy41EcCEyrqfk7soQ
72vBmAJjwPdMukPoza5RPE15dPGmBR+UBz41Xex/lgVXM3Je750S8eCOyYCrD7wi
7TOfCM/bY+EJDumM+AiCHsMv23yXJknHljNqjrZRmdiujS5O3vTfKESYJi0ee7bh
BJL0bOFnv5pKpAFh/6NOKKZJiN7ODTiGY2+0EJ533+DMcdCKr305tQbk6rBBW8Vp
MneL1tRL/CnxtmhZs8WbPTg8wWuKVgA+rpyQhfP62pvJtjdWiAm/8m/Sjr/HCdIh
17gZl23eYUmBlSFkFD4cf6zL1fGWOeL1ixR4/JDSZsoiZePM/QMmat8HSEWqStkO
xo2tjYNnIklXNV6tm7/oLskxX05Jm7/klzf7kHMLa3jKKCx76quEPenOB+gnYjbe
gSmxa4EMTPpKpLt2O4jH+UhEnCjT3h7UH4A5gtoNNoMpCT8Ba8ZV7YazKYcrtYG1
UftPYoCU6QM+yI2z4NCvBHY6QgSzrMzYuMwUJ5A6Ud1rsUsI2JzpxQmetnedm1C6
mwzulGrrmXuiRwmtqtPlIQKtyusjYOQToXEH4zXhwaBQzxhvLYwWS0JfrwOM8BaI
OIkO72vSiZf2KeGFZ3unlmLP/Eh+cJbCYD4XSemKTBrzuRyp4OI/2GjdUhh4wInv
s9wnslR4hqXbV9NK5f2TiK2ShWVQlOczfsUKooVq4uLxiagzWZuL/mpuLqX0+PAn
IQKme0oPqcjPp17m+duKMCmRLgtcg7c4wvuOLEhy7fgcjP1LwGREuqDtZaFgY8P9
AK1v33MqKOZUFrRx57JIqv+/pu3p8xcXEE+pjgptJipI4ETplW7Oimh8iDje7hhT
/XZsQe8LThaheq2VaNC9kFdO9SiQDB/uggF9BnAjGoo7tgE7W1pJ+JFDyAigqVKu
AN2JZL3qovFbjrilnxIoZYR54fEce1dbkQNYhLqDcEYRspxQPp1OXLuS1NrX3Ly3
Vzm6GAVDk8JSJsUKbDldp5zvtpLcZMvgbobj/SdlXZ9ZFwjSi3/PKbPyzyR1m2Xq
nZMoEgVXcPwHJEm/bB5pRm67UOdHlut8sQDGVM5fntTHV+OFPGxK2XDLsAAeSPT6
DhjhpGsbG2+YZtqmDH2iEdjYwoyl2J3nLY61H8ugAvmDNs8jPd9UsEKouD/3Wk3z
AiTohNSEcm4R7MkNP4I01ot/kEcDXLFY/LLrdzAXJZA/s9zTg8tFGQQt0CqerFT6
1edhrMbsV4v32ayS+vr7THLb7kMVldWDsN/vxMRrJ4izPJtqy3ti2kvNP0KNgkJZ
/i7CNhuqYB9pdIFzmNu9EsmFOTer2LUFN4zMCTYlXDAgOj9VCCsQ6LCGnP8vChm8
rMMDmV/zEh/ZCu7Sy71h/YfuNzXOmDSYVRpLKt3CsZeGD18RXskcKrt6O9zqwHce
WZp6FNQRkGKSrLTT3qKNV0BkgjrF74gAgC8W/zqR/n4iotjU+RuLHnegE4H9DrAz
FzlEVrcpLnBHtgx03R2jVbcEHPHK0/6MCIszy1hxT89yGDMcIzh1tpSQl2PUpK0M
9pwuWExZGwicOJ8VZnlZOvLbBW44QABCuXu91RMWijG4QpoR+Z0TUnX5/vGhTWat
UD3mjvjqoG/NI8I/VPopgPxBCAOuUmVOHn9KaObEx9OgoH5gRgSTFeoO8bO+BN2D
3s8zLYOSlSDnr6NGaqPI0F+eheUlhP9aWj8GLp5FCDg+uBgPXMjnHNcMyF542MZ9
ukOAyAqFEFzDLvlWhtMhR+aI3YTOoxqe6DypOz9p1M7BxkEaNwmmUWF4/drXiqi6
9eVN6a2nSeP4tnWn4HBUJ2po9JB5XgOrfxYtaa4zxcvXjDY6DTLbt23KNwJsxhjz
FtyWII3uYJQNhJZ51oS5b4hICqMqsypON1i9duxFVhsESORT0+z2wmgZ8Vg86vfO
0/p8K71nZjHu/MTEA1zGSzURvGlQ78KI5I/QaxdVZrUYeUQDOF8M1tRc2tF9rXCw
ivdXpP25cpzNjC3QcYT3k73h8xaUS8OLJAcMukQy3vSYvaCwP7el7bDM3Fiqu8Ub
sQVOsvyf3ODlRdDzdtMiTBrekpSKsoWBbNm3f2BSf9a2scyhDTD7rXXgfc5ZHBU6
JTSriOx9Obb3lcKhuYC5VGiwn1Vk5npcFLwZFbZQCke4HVkDzEhbwSZPzVgX2dwT
F3loWXEDId71eUqGWxtCjQ3IGv96cezVWSjzujToOVglxI+h6lQaz8ckFcT5e9IF
kbU19QTY9hzlHy+lJFT6e/N9wpospFsYqnomMVFqqD59AzhaEsLJlTYx1t/tnn9d
hsHDtz1JY7cTL1GuqEni4nDwx87629ONE/wSJPP64zVUKzLVwoJ5ZNN/ERyVjLgo
64lklMHT1SGA2XN5xSnwTned0z2fAcqtInjvYhk86Xu9umYEBk+Ha5a9z4tBXWU1
++fFtZeAQnKlx9D3hYgm+VvWB66E+YTMNWN9HFbdFO36NAbo1QMAuSC8tT+X1tL2
xzHFQ1LBXWiH7e9N6VpoE2WDrhAET7eeE7LI8xobjfOJsaMLIcXNurIinXQ19zGI
TbJ6I1YK7NqhthNN31xdXuXEq1yhQY4Vs5oHCFGcS24YsgQ476G4qAei1jBz/XOh
iLQVHVqUyczChYcrIJTf7zDz02sZivqrPlNJ0aP0cYtV0/GXzwVgrP69yZwZpdZe
vpSxycUDWfIjZROzn+ZHaUQ6vPPdkg5WaIKEMV78sBPv73grUU6eJ64MZhco0ZYZ
wmMoT/NBv3iRxuY7ktPL9itjdYFzl2VXdNtZavLpvHOQNc9ckFv/DdDsId9v1gM9
xjybCX5K/iKJ7WFFjp/KgdvrrOxsEI2HxtUr3o2KYnIVw1tX4PDT7JHXFcr4Xe2F
mm1sn5N0ZcYqafuA4PcYMOJkeP5kaGoj51kJx7rb4xyr8T4mfOy85e/5q58hLQ4+
tMkkc4ygUv5hEdzRC92dKAUPeS+Yj1rQLHThBECDHHh06Y/02iyGKNPmmOlfSx3X
ZCLWnFDT/yPLY9GaZ2UaLrLl5B8Ca/4FQC0EVeXu4CB1WwY9YomITQRJAR8iHWav
vFHpfhhMjLZvmT0pFe6gjOCobdsc/nTRhyMykVTqDlDlnaOkA7dDK4b7GzBBYIxw
JvIgpFa1LIxOhGq5E01sP4Tr7lF88zDQKZcxG4SvMi2qq+BzSKJBmW0J2n68vgi3
h7StvvbgilsDvFIOn7agjhKMkxF1aRni9FFE6u+Yx1QrKmPEpV9wyBPrZFt3TbRT
AXHbY08KdEdPn1cdWf7fq9sr6LG/PXeVxcRxlfwbK3HEquJERDWS0DODpbA9lWDQ
ZrcOTmpLr9abOaWSKdZLt4rhetm3pNX1Yiuo4B3w7e6Pu7HDO7WKViOXfIlPsWjq
0nwVFZqoIGJoRlAAn8r8EtjXNLXHv1F33PW029wIz+PilUdXCGve2hUvXQYtkpxv
kwn3B4bh3MjmTVMYX1tyEgwsEoGEyMKG1k5fxeQh3nQbzDpVaIzgu5T+njMgA0eR
8frukNeZYnPq1RuCMT9tt1obuw6sPd7XmK+HzrY0GJZX47PKp55Z4qFOVsHj89CB
/ESGlzHqh1CxG+TAgOJkIKc3KnZYrR1onG+/8iMqohQ1mdKfVpV+2WiA76ra+DaI
vcFmLLF15hmM8Hfozbp/oKPlJBKFeRyllskmK5+X0RDcYgVBBe1oGtD+zGgTDFN6
NgOi+Fk7rvZF4ASkCBW91u1aCJnxiIiWKqFPAmaR0+9UVf6cykdzd4WjHyywumA0
QKy9x+t7H3QquTa4KGh9h0lyt5zpxqMAq49dJeAxuAKL4xiwz9C9i6I9kju2eZz2
/5lT1kKJmkAkFQF3szCPPEYh9OY+tPlEtq2mWMD28AA3Eq5zHVgsg3gdrtWshgwX
1BFkh0lDov+y53rTj588Dasl3FiN6RNh49AjvVDNOzAXTT21aj/bC4ITyLyyNx7e
5G4E9/VhRKpNIzu/pCdWrrsHpbnGSx2G1pDeL8OP4k7nnGRLnNnZEUGR0e4aEBRs
LNXwIHxvqcUFVWt8osXa/DVM1Gj5/8S3Vf+DVTq+I0GaKzV0PjE00lFTNmNIufDb
smZpbhzXk/A2Wf3hd0AuqxD4zFKlbZN+k3TDCvnbBA+VTxgE59/xeJO9lY1G8R46
+EAgfrEoJrcAG50ueIoOhP5vVFrixLkCXEAEry+QCJWLxUlrXnMq34OGENmBvqGn
FArvRUyGvtimZ/1qpF8w0VNaWDguWA1HaDwWr+uDkfs80EA/eT2ZOQeQVJzOrnJ+
rFZtzgUWFWSpwulnCmsZBktbCUtT7rgOB7PIe1pImotRQC/Qef5g1x8jcE67CrwH
hfP+xwZ2UgwJUghKarkZrgnbbXVBzNEL1/Yu3m5xgaXOq1jRHK/R5Qd3LM4GqGHI
uIGr3GBKrQwq6TIdmePnha8wv/2Z+SvUmitBfjAKpb1Mylt/pFPMIbDiO4jjkQ6x
vhJn4lVFcoYWXfproyjHQKlo0GZSjaacYQuOokC1TDPelFIiRQN3pHU9bMsyf+kV
TlgXOmC+mQcj1ZxZ1Fh6JlZbGWy37DnqtiEbJa9J/G8mKNwvR09jGouLcY/MZyXK
CPTVA7S3pyiuQze+MrPvGZtW6ZN098ZWUj9S/jLalVxCTfR2XE+1C9Ovh/XjG3Wn
hBjFqPpGL1gB4iQYKBxnZy7iA1SiYGN2JuaDObHpf9JX8ucqWmMat2suH3HJM2zd
5ULl1T4UiQ3AJJsH9SMK+MRJv4nrRqVY4G3nZvo3+5X6gpFD4k4922iYpPlC193h
9k+5/mEBB4/JqpAwh/K6u/6gwPwbRLAEbYyTANrif/OnzGkXbyaG+A7Ngh+jr/Xo
49bMLh3lBa4hkeM2gcKdUm0qaAAgc2SSA9O4mWutP1oW389b0hQFO9DMQ1+fC80Z
rRMCoQRdTBNuYXS6x6YTN2mlw2vhqMsiccJGRPKrEQnh4mw3DR/vkU5RvosLvztB
+i9zt/sJS9iC5FcAA+3lhZ6btreT5T2kHfEbgKidYLYS0YOqkBX/dbumWEXLaf8m
twl5mYPOh7z66uXZZ0ZlCKMHFiZTgr24MhXCIjRCQV/t3wc5Fnxw9Hb7YtmhD0xd
pUu5TMAO6P9mfmvYcadxWuP2SnGXdaNx0KZ9TSNGjeD0fKDynvYH/j2TNpyOPh/d
eZar/XEyn53R4q7LXoE81Aeasgm9sAO/tNpLPwBZCryALp0G8Ks5kzxrmoenVmq+
1N0YHDqBfpndx78Z9/zB3dhJ+O4yF9ZVVV3EeY9HzT4EP92EG8LL09YFWfuWcNUL
CWlg8o0hwqI7D8kJvb/MtkZYiiA7txwZ5QiIGFbB4fTZYb/v9fvY4/Jhuc7LbQbh
cUZV04xB+qBUiZRIcBb7kvTPxJoytl4hhtUIhD+ahsirdzeuVVCL554TYj8pqtUo
WoAIDYfgEHAXHEGLr6RjTJIyfyWTk07UYu0uNwMarMzwAbR23V2CzWh7asH79NQG
sAPSdqqRPRf154e38W3YDbRRHpn0Y/qzk+aR3w/UbR//0tob3f8eVn3drztEqlEA
joB+t1QdR8aBuIFL1iPbH+Hb7tdXIWBlwrDQ323+lkhetIYfcgOZIbwIhtQHDg/4
jvtXI/Ck9zFpZTHLIVczZ/tzPFNH/GeBhQv67wwrCgHIqdDDmde+mkvxOe8eAG4d
32NEGXglhD8ggMR00ME0BRBmYclRVBQGEo/uLyRxEeuGpdRcB8GkX9Zj9JSJIPf5
KH2SvoFkViemHxDVUeRUM4+r2w3t5EEH3O5VHY/2u+ROjuHH2RNbqrGhLOlvybWM
TT44aXozCnY50bNpdg1nSNCAyMML1m6zKssrnr9PxzFP5QoAurIQ+LNUCRqJvtbt
AmKNgPpFt9TyTRUsuc6iF2zL3mdKaywPWs7odlsyY0DvzX3eLnMvrlGthjDB2UpL
7Wi3zOFDHkrLdERk3/k7ov3zt/qB4VRXwW5F06Rm4POd36ISEY9o/vZZZJS3/IO4
RhZ2n+niw5gEYwHWzK1MlHBPr8cGifhAe+k2FP6Op42Zf346TXbe4ewisK/Voh2k
+m9dkZ/xVw3Bxr9cdKIb6aeIIjyGgunxOKZOYeKCR+zLlEXhV7m1vZV3aa2DkKUK
xlClJnckB6gR1NFHZ8JBSxpisrTo6B3GsA/LL8tVNnxsGREOGqowGzmzz9mooBrA
yba8nyYmWPHPrH/WmXAG9DtxZBTD2gVMM1ty6UAW8bRc5o7bcUFd+OfS2CH9iL7t
bqilHfEp3XNhSm+Oje+rdRY5UvCQTmLOYRTYSz6ZgwVUVMaKaXy8GZLoS35UXYRb
RGsLyIKYMtQOsaGj9O1JvR2dJ5eoZxs5AfUUkZuhoH2HUJUQzmVhh8nwhdYOPLEL
mrfiiWfDXDqlf/6T8Gf5v6XfOfVnXMJRgy4tw6C5mnYD+EvqEJUOY+VqoNNDYh76
JNcRd516BeEGqSmNQNmpKeLxL5c6eB7xXXSoAv9CfO74KjS5dteiNZh24mSZ7rYE
DCJ4n8IgEKf1PuJt7/ZInisnTRvXC5nJSWWYHS2/xvQ6A4HxvcAnjwxEeN0Njbm0
/1zzTwWdYFkHan2wyvzaqXq66ga4JsQPr3c8TgpNzktvqbTSLCtBCtUy2AxxVu40
ZB3kXR2KEipfm4LbyH3JZz2pFHdCI76tZw31GmKVfUg4laHl+Gwm+zsniFpWvT2U
FtNlwinWggCRyweZzn4JbVuCA7sPaYT1ed1CDBOmDQVMUzgETVi5WTtgnmE8wvWd
36hDEMeWQQh2uFJWzBRYeiOiFP641/rdJlbImoNsFB3fxacAS2CH5pdDwHqWPG3c
YhJVlxhtNBqgNS0M74edVVXlEKdIGdMvCo8JM/GlDuHMv2N/9RYMskeyQ7a6oSoA
h4wZDj2IGWEaijqi8p7YWLyr5/If7Y0erKQX2SH214sERnqO91rVTd8F+AEeO/gL
hcWuOdOkGli4nGCFUdpmnsnzJOlwGwRuQWfS2BEIsQCkLIX9yJRP0xLPwWcyxqWS
g7RUpbfw/rRYS9TwOKTH3kl2/w3JW4fbMWyaiaeiAI7mT2Ns4tkrsoPwHHismjIO
I1xelwteTAMu/7+d9D7pPxlIqkr0uEvTBof0CfAOVoErnil7WoUdu8uRBZVCii+1
2wurrLrxeLdvMABo060lf5suGhsb55fBY1YHP24yRbNe2p3sfqWakGSFX9DrR7U1
xurskDlrHGPTDGx0QmnLiE1oYFhh+PmU8RT8nAF2hH95w4faHZTam/1hBhx0euMN
duMMQdfLsQGSxecZpcinUNPfxoHD4jH2PriL37ZSTB5vDyEqbdd4zqUJzCjJrexN
Z11EiyKU5FgCg6f9RKz1N+nje/CPhy3B+xJjbuMSVquCJYXsQCa1fnv3I+JYzRcK
DD7FKVmnntGxPe5D5fCxs5CACgsu+9VdmHOTC6UXHdZAN5c3GcmpF2IKhSbMxB6z
2hHjGvqBQO47OGdrrmAjxgHFGBohxQo8ML0vhulBL9uJgjr0VuN72eILQ906iSTa
u/gOL3h1DgRM7OSMf9HYWOkXQezkxM3nf7UvUtGyh7KoKB6ohyUcwkfAL3Mv706z
HLcDLZXNgm/SKBsBQImxPjtmBNo1ivP+NZVvDQ/nSlER6FkRtlBywwzUwMmAm7sd
A8KHaWKYjj7hJU4wPhC9M+jy2301r7pEGe42aBf8GG7+t+3Gz0FYvq3B7KDLr5ii
M5hjcix+eMTAaXjMZh3a/LnyY48X64ObRCg4FySm9rhQCz9cPWYRmwj8VeZm9bFe
Yp403NZ1kapcpZSixxM8LlC2+tqiRWjiUDEEH2MFucANWS0+stIgaQ4eeSp3BPWJ
7uGNbiernkjrmtdJVRY15GD/50Dq27NiuNsjyAnMx5yr4VUUvQYSBUIZfysbx0tC
+gz0xAK8kmKXfZkXlZjeuY2afPrKxXvb9R56Zupr6OuPRKmuSX/DRxncidjKwZmk
dr+8qkEIiZAp/wyORmXVEhe1SUP9RdT4vHR9kCKjAy6d7nTJ2rZWcecSrpzld4HL
xUMhFfRvXI26ASfPRjgc5dk1WpzWHIWxpyKxrubRtYf+n1EC578AVdKWG0/VmfbT
75bkHjfHPHEfYpU/UZ9SqBzu+wbBmeLClHEYeI90+1KODlr/Mleth+Bzxy0UFxXt
3EWtzWFdrKigoc8mNvjFrLkD7bJNSIN0SDeM+YI3p30HLl/fC9MWS5zPV2lUJNUJ
O6zld80T1sF3IdzrGlPeoxuf5S8sIHxo0yhc8eWQeUUdjDqA6WEsHr2Fj2GHw4se
uTRLPFEQL5liyxc1ezTAj0i/ZkvLqcLWZgWtiDN6Qq2av7GHtfs+VYXoSrCQr1y8
+r9U/oTheOXofzpO1QCAg9SWb49pmwg8ydDKPMTTlod49jXlJkFkcU+cXFYIRnK/
qzpwjqqQWUVAVEn3VleNdcROVGeC0S/Z7iEeCwHfUGupTP4H4gn6tFKLbBrMpAEL
5byDCPM6/6Ro4TeiiO3TSqweh0kBSh3WNraZAws5Kw571gEDln3g/zyV5kdRcu7y
9dk2JhrUKkIXuojkPySSc+osaP/Vvg4zrNCODKyQEzyWp6Uak6wsKdEpjdyvgif+
k+wW1FDtK8zmT7MN1ybieVc1Z4NS0rS0guUGD+x26xMubiV+QMd6Qvy1LjdPgrIf
I+vnhbOm1FqA9I2JIQXZ33zoQbi1JOCIdU4TXaTftTl0uYAAyo5uyM9GxgT9u3Jk
XEkkRBB8aEJT9f6k2o+zULhdXBDu6kzI3U4KYE2/vwmoY5oGWrY3pZaxFwQzrx62
OXDsPwQU2m6i7Zpkdflpotq3ogs7iENRPeX+dc3HHNHRBolAaBSDQOSJVozQ8Yl9
3EQhSzDH5cWFwfFGOkj1n1NLURwIGqdJM2SPrpxvnfnG24MNlCAKugayXVEflbN5
D9obTz0twnrFKt8mdJM2UZZvAnwSA9JrJtDJHe4jMX/qY7ZoBBV4V45TDpEJTu5w
hnL3WxJkTzcua7sMnKb84Tu+CW2PNSu6NDBtad8cHH4nFPLh1JIaanA/WoWMV4qT
Fz0xXH7ttIH0h+NneoHYZxgdnsrDv2A/wovWQc+9ltPpmGPgJzt6VViN4K3KRJzJ
HuVkS89gTu+coTLu9ZfhC73fLHyBoU5ylFt8aE/gQH03jOGeMByGNvJM1AKUJ1iV
LxKnn0HdZOwHvYlVFKLSv2BmnY1HAuvKy4iBD9ZGXFyPJL7fFcRAsTef9P13Tl9B
i/XFL3Eg7ImknPAVOCyw5VVVeU6OXLAsuc5bXkSXv2HXvwEB7yOyM5OhkF1g6/QT
6ovxHrboFBp8bcrHDKy0x9YdiDFNiAsupuufsFLz/XaX6MEXXBi4VQ6t91lS92De
NiigjFJtbLtl49wkJLSKl7d1+ddsAycc+329brUCmymWh/JFXW5eDHFPZqtRKJ+/
X3KFMaLgsQtJ6VQbdIe53Bp1MzW68UbtL93QDev1oyB9Dd5NYdt4Y7qylV4tAjlJ
bZikoirJ84CqCWGyGmK/O0r++qS+VzQ/cEkUxBU9Gulo+g7ebe+D3/Z3gwxYswfJ
BocdS1do9r7x64IIvsuN3JftysCF6rjstQIwk7+c5gzLsPLyOPqeK0iAs30cpWg9
byri81tc7AzzrzWrnKERxzcmcnoatOJIryKxPwoEoDhbcvqCok7Dg8aJZtd9OaHo
eMlDYJQ3OvgZIbaHqIJAnIWfeXuVxn7QJLlEt0HvAfolIpiWRxDNGWDESWvye9qX
eTsN0dISpXUNE/kRveqzTgwMktZNUKmlbfRDzEijIIZgD3b+ouBU3dbav+rhQ7X2
/iWjUH8QrUkqps1mHJr6CgXfuIt76o10GSV67mbSHGriZdR1FZGdgcs4ZDIxkq5b
WSFfg8l/cCoFUZzg7uZo8QPYtootGw9aA0go/6mQoU7e37EaQ3hAcnX7JnNGU7dM
c+Rxcruo9XpsWwB7R7mEJRsP4Ek66rRK1ppUfxfVOCc8wTeHudE3Nuh/uWAMuIZh
1GMt6hRn5NE7jD3xxM1VFc4xU63QTcqfj/r1ZyAaCI7FnhjAzgdgvR5uV4eQwwmJ
ozO3ABTIFoPNG13SCiAM6H27vie9Xp6FimYhs0Y5ZqjBAL92Atks7WQ6ttUCP7KZ
AL7Pjf1fQv6pjVfDiR4M7e1Z9tAdFgKbcQ6FOc6rym+Oge4NwO+J9g2jDFrOA9Gm
kONEH+0/b6hQvEdXn8vwtiA1D/IVq71RCC2MZCidpAwRACnMGUVIaGYRXL7wVb5q
BA2tKphX/FgMqtEV7IV4WpiPeaAhJe9qufWUqjq7JtH5EXoWkdEXO1dQuVnDK/or
s2DqKgp3r+TkPljTz+/kXhI3fwXCdTKMOtbI8W27m1YWIHT981bn3sUdERLGRaKF
rraot/IePtsWI/gRXgFNIbRSUhGj5yGGNP5GD8H7Wpnp9c8VvT6xSSRml+VFlor6
FF6Fuk66/MVktpULY6/mKyb1BL1MAcLABxKmVQst9Wb4Txb4DuDlJZ5XmLdxkoF+
4M4AHID32syNIiMYJS2vrv/pWXqSedsPMT9etorLfjsCse29xNNqK/2qe+6ygCuh
AS8Mj5r/n4rMYfA+lLJkMyEE7ZhZ4OXZxON/n1VRGffGwGlB5mXrH8W3Nu9thhXi
/+EQ/qt6dOxjLRVSGzhAPYfYtOBxuCYwq+I0w/lY0JQmWtmc63PcjzZJOfQi3EVr
MC7KJKylxFdZNEswn+mbY/eCm1aAZ8muTeYuQEkkZRboOsTeSmzyl4wXFSx8LOhk
E8wMhDz10KDlgT9rJ+yMpaN3BVxiH/DfllWi7alyOqmgnGA+iLv04S97RkiTO9VV
qfpRSMM+FrIoKaHz/+zHMUTD6iidT/RNMsYpAJJFIDe7a/uBlN405ZZ99NgRNser
DXyUOexeUqTIqKPXySAZCvvnVUMVCrOT5xD5iB4M/VMjq/0ZdWD4tkVDVHZ8+a+Y
RxX3AU3INVb/EzrKT3dh0+yTi7Iyvc8+a20pnOqC8mI+7Fq8FqHdjgzk5/77hZx/
p8yBD645QrXihWcxSxwdHcOtm0Cag4J26MKT64gmPkNHmODpysEbtgp9YoiaGzKh
/ZtdqZfgFn+ClHHCnRcdcQ+NMviLp0I9anT7vZbYAUTzJwnWlVxcDli/xhq+efVO
j8H7h4TprnrQcrTSu+peX9DQWLbk5UMtSmj2N3ZwT/tnvKnXLYl7F/NDdi2/ua4B
kaDAnERMwGXRFmFJfwOWgd9qc0A8jfRjSS5nrkJAhoseTwBOa1uA8B2nPYx8H0OY
y0WdZ80/ESewUyoFTf1Y0G14o6ktMV+4IAm1BeaPaJw9uOnT37XbAaSJwGMMTPLg
ndSt2TXxaAjkLbbhGXh4lm73F0EsZ0YzMUTbRGJ0vBO5br98A8kjOb+DqG1/x2xQ
mLwjKWYQ+e288XuXE62TMBwdP2/nfnreVmtjhC+hj4dMw17D5ii/0tIOVzabh+4Z
oo2+oA33Elad4bMnfPfH2YfuNkGKxUwhYbfE4HSSl4erdjTcMxtlcHOqiYr28KHU
fIkPG6quIIYTO+Fq+khwrABJ35SWVpBcYNrsWBZ9w8A5sidoKS2iUj8D9HotrN2A
hpxjFlIZJTe3QO56Jq5YVi+hKU0YUl24n4i6FfBrDbLtTU41wAe9FnMTfnHD+SoO
N09T/4nXNRMgFhLlisVHwQbsU17+eTHN+uzJJSuEsLtCElwPieYBGgINpV54B/p9
TYUcjGlEitMiCFZ8zbVJB2TUDBrblA3LSkMsnOVndB/z3rUw7gXUYERX7qWDJORr
3BvNcsQN3Cf37Y9Ctj0CSbVdLxURDhSR6VPBbdyy3Zn6ZX2QsjM92lRauERfcKDG
sPRQtVNvJX2D1P8SOqw/iRkteNaGh4ytzO/6Z4K+FxgpzkXmAoj9jN7T7V9Kbot3
iY07HOZE6XAAvnx5YGRPK7ZISsd76ehxgGOUcPjJdBAX442WufZMdT9HxHqgRZNP
SO2C29HW4XPPZwu7sOs4+pQo3LRNaCsfcSDtx5lJIlHx17qircoZ+7ehkUBqswkF
MN+ULPDO7FrPp7lxmq589+yaqIttbm7DmBXWQqKybFQZpcxCda9y2S9KIY6SJZDn
hPGBrQvw42rayHUVuJ67ia5jgbpa5rbsz1BDS3cZZpG51ZYSYemAWSmGiiLPokjI
lZTtfFsI1r8WiVNKB2D0JhTGS/XA1Js5T/Fgws20okUAZhIMycU2btqLcd1ib8vG
hHXIhOHGXKfKi1ptTj1NxiDOntajLC0hACyyDgH3bE3Z5b+3f3rV8unEEdNZuCEE
lJV+PNpM4O80T1tqV8bXsq/cAVW7vZMo0wUWCzpSjtX1NPpcazPOZ/tuBBhAG6Al
34kgB2syiJ0IF6nsxbW3s6cE9hlYC3TnrCp/SO1HLZ/apRHBOxn9CVhIJ909NGNQ
qdMKYfjgbLAdfq062KwEu+hRDvPUlKX/VZlGNKoJvpqS51+/I7zGhIelCMchMO1o
+60t3XC/N8QNvKmWg3i+YXn3Hcr+B3vYrD/1F7mndcYsgTv3hOKWmzH9yB+DwW0x
oQDXXN8tO3opr87WDFe6A7ajKcJx9evtOHNrxTc+rQqe6ZSJIB90a5cJ3rl4wbHZ
gpbjrPijEwXnJmC5pTNDnC8mctpiFPyeniXiYW5go8UGQCd4YAcj5tzKMhzUKXE+
j6VTSoibm/iRrJsfum8rMigAdk+55oMFOJVLtZO+6EjL0guv9CM9VnvWKaJ0hc9Z
0j557AHK6WGTW6Vw3IUlwPBDL5etot4olpuRqvLEZgqqxbUxR7wcB9Cjo9EA0GvG
wjwwSG2kH4QAFOKY8yW+9su94rN91jNhN5W66VqPrWdk7QUn4n7ZI2bbYIrkXow0
PdQ6kPYQJPf82mlkj2bQ63EFHr/XOEwNjAJxZ2+I7N0/hEptGFYGW/8bXQYW1pDw
CfYs3fg4aLt07hlw/ZclCdNMPX8WqDCGaGSDLZtzuLyyuUdE41tNVtkWkW/5UJGA
nZo5/orlW+KPSmvuS16Wme+Wta5bGg66hkN0FaPWw3pqO2T6x/mU+ij5KfM/Qfwn
o2Lu56Q/RFg5KU0Qzvc38cldbyuoTlwsWZJvZw+LiZ8xtmUjhWl31NbHJsFfzygQ
0mvh44PGTJlX/08xBZWjgwT3UZjJwVQKoIxbSLkI4h+IWmQX83exVkaz2IAUQjxl
CFPneoAdHgrzK+kk2GGjS4GioNoIN3S49LphSm2NdCJ10sN2foBcg3STXd4oPTBl
+J2OrQqp82LCwBC2awoCWNpqf2eErSUACYoQQqZ+n8/4ixRtc4qhewwjGkbLy56a
xjoZeWzV0qHKJ8EHEseib7Y0yzHXXNKyikdRzGBaNDZvwjImtgykX5IsovLItAFy
ail2GhKBqRUn7G4d7sHGKf6iRvWVm/K7g/TbLBtrz3c2xkeIEKzwMrgcLyKsjdD7
9JuFDEXQ9/H5212iPtjzp1L4QkysZX65RwhAg5znMaQdu9kvQVklOFxKx/Rxblzg
7b5jIya7zb3ulbzV808MLpvkZWgvw6KbszHAbQa7deNoMw7ydjGP7HOkmc0rfDMk
u/pCWb+PLW8j/SsqnbDtABl1O00JJhvPFtlrx5fCP37exNi4IhOs6mfDVX4CxRO6
XZ/8Sid018FXLbz+XobtdBvVW132Hl4dmvnk8lYGL7ieUAwEtZAM838pOenTODYH
J2Sd+/P2HGf/+0LfousAyn8qaIxraNejWAHKM9gvl5Q7OUlk6C3JNL/46rFmDmuX
UdJxf22rHmXmOvVk3ctvd+Gy02wspFvAQ6tX+LrAo+e6nmH33zaXzrM+7w0HyyQ0
VIpl6yHpf2gG9cjVDKZaG/XU7LAHFDbSqj7WP9P2dTxU/IdAZJf8JV25t5yC+Xsk
gy+Z/T3JPf0/wzEfcVsWikuG+R4loD0XDO9K85ttN5X7YVHtzLzMF5SQO2zBnYnQ
a64YGj034h2KvMsOfmt1eco02EfEnZj1HV6sU5gXPOn0nF4x8ywtlCtsty372ZlI
ZuIKkQouOd6CEjYq6LWhNgwc+PqBRD4VmBBDRNv4fnEhFLurP8hDfVzejwbNIFSP
AoS/7BkBrD1FdvIeIBogl1e5saUOJKuRdjAm/7J6WdatHG32Iv8Nw9gcrnji32iE
RLxPEgmoCtFIEIKiNclOrbYCgsZVNp4cpvPZjFukzABKqlMJGqwWOtjtBpNmqOZP
o+GtcAfNc6NJjEGz3JzKHV/lPuu9oK5patjZNQnaUrJrkf2bQHvodYr+Jc7lBLHw
RRk2KsbvnUYA8J+TP4y4GDQZWegvq1vveiPjmZsBq3VfeeNOUyYJ4tOpk3PVKC3T
QN50z1Gcd7PNVXh+m07mkJsh1pEPqxsaLXRyYq9MQqf3MkpluNMnVqSO4jta+ogE
/RDjyEBvqXfm6t0HixajD1ZTAgY5xCVJ2wj9Y4oGGu7Qubyeqr4+WCD54Ph3iFBe
/w0mv0y2AiLrIEbQVUwwW3kGMmL5Tc/Cj+KS1btzjtKaco0mOD72eU4D19LvS2XV
6ebc8/Y/eBnIBJsYD3nyE3XZ8P8ACUW30RlnubvlVhPUaKJ5OtQE+4r1vMdWn6cG
N8p1wBRF9K5A18w8ABvavTBdzO8/uR7DhHkMFU5qy/GlsEodqKD6KMW2ZjghHDf6
2sbeEsz0I0DVszjg4Ifj6PdVErbe2aTuENEJ82ciDZVJn0ssKaI2n85d+WZLx/lN
Wippw3P1e0o0KuqajlyMY/AofEdHVjUMn1h6lyAHwzcACkV9A5mp7lcIT+q9y2Z1
kh6bn83OD1Kf+CCpuSyIaaAvM/UFeZZWiOst7hdQ58SjbmRwGw7FqXT0iLW990XB
ywz2ZFh0vd+DrMwG16ccDV+WLLbZb/WD51AYr3frL7JpgAJ1PSydMaL9rjNnYBvz
hp2bpf0/JVcIoWmZhvcWLPTZU/NeGgZFyAUbcIClM/HGVnNcSs/k873bPejBb3ss
HsO+6zMa0jjgMn/6kgSwKOgkh0E+sMoPRJXpgioVwotrb5El40QQUaAlaVSuyYdA
5jQUV7/sBHwp+8NE1U5ykt5aJv8Wg/E62QjuxH6pjy8EIVHU8MRNFJ9m8HnEsfg5
hc8DgDC2CsPkPx+g687pJeWWLUGX75jg2MC3CJn9fN43ARdIPC+wJef9eQO0C8x/
WBLAW1Ubmsl13fNnMjUw9QepDZichVU7WGUfM8b6apb3Dt9hlmHwOPvgE4F2Z6AX
ABQ0k2LQLI4zb5bFw5o1nqdZvwGhoEJFK9ZNl6NWq01ZsE2hfp1N3RV6PQFwa/jb
5JDA5wWgxfD6WLsM/1fRkzEoaz79f45HKhYxIEj0Au+T50mOfYAd0b3/ds1fcGVu
zUpgeHR5jLR0ywPOWcnklIIVrbvEM1Wlzq1igiRTmHzKmXsBlgemA6QSsfvp7adp
fHlaIOWtCGEZimJW2D6vmAP+vMnNyxUCy7XEVLsgH21pgEC13QEj4LZvC8PClFcf
n4Rp5wSL1nL1Cp/6Lvv/dJVQZWmmpHtQD2OKdW5EQhzP64mIpMcC+uCAXnBJmq4e
WlUiRI0UVop04sLqPD6jnbp5w/Vy8CVu8ZCKAMV/HMq908Fo3hlCN62UAF/Sd4x6
z+8PioPNlESx8hltxdLr40omWJcvqWDIu+/jwTWUr0HFzAZ2zQNNRldQPeohGuZ2
Roc+QgASTTaE/zW4Hkf41dAvHJcdU+CVEZP31GfozmGjarQ7J0M6XsOsmgoraD+O
A/QI0pFS7ZlLCUS+0hd+IRM6XTQpHLUfoinv6v5dP6UVaolg1kRKn6DEZGNRnnFb
2b6qzs3i4jiD04b9oXcTf+T8uvkYy3D3qHzcxSppVT2zWWuVQe5XoC92KAio99d2
stow2rarkRsyPfb6ywOMY949R+k4UQ8X3PnANLkf14KOxvrZfpEVhhwTUxoYAX6T
5awAkDeeDS31YAftrtbTJa96XEktAfZSlg8UGcmZh9ZwUCEaM8jyGVQKVxjbw1FT
3EFOHlRv76Ed2fWha3g4s/u7biz0LwWaCDiRX6nDuGRK5SbwLnp9t64pJjqTRaLn
+vyCuZPjApqYF9aqeeWn3tIj3ggh0xR9e81kf9LuR8CHL7nqqCvsK0th1X0+apal
hJuIcbSFPvR1CRP8AaYkPiiAUGhVvbHMbkCDmuHtqyV9Q89Dw2dFQ6iFxw8JehpK
Pf9guRejrv1XWBtTObmCBpEjq5/FXABv6M+jZ6oFUXctihUW55Zo/pp1hWxU8zuW
ncm7i1nhZW6sBxpP2pb0FsI+HR1mt1fE1qyD8d1L7ED7gl19xCMt4S0pkp6eWfhI
XB8bjRQemefP45mFtinZBtGAjJLyEdEwHGFZA5NvaiFHMMw81BP6ZtFZeIssNz0i
eTziK13XCqG3TAlOkHkN1H7otoWx/2bEJv7IEFFif+vDL6Ma/Zs+wVfejWQsVya8
fRmCm+Zn2Otd0J978GhM5CF1Fh/NUX4tu13OaYI0vteg3fT4+Vub2sukaja1aSKx
Ev0MQ6IrQuAfXDqpmrVKK035jxPQ5nBs7D4JwzhEjvyq2/GXJHki6KobXft6zChQ
6w+0ZRJQKn7N7Ox9diC3U/jxo1/zGYhzDRS+VR++Nzo3VrnGl3r3k5KfYPgkM0U+
FXDxQhcW8EkmLEahuArrsTkWdV/H0pBycdERhG5OOaqjlOPIaeZZ1NIJ5Snsbtl0
0VR7ALUNcnjQw2D1l9NaGcZSv9TBpc3nYa/xeLYYNNflkjBYXUunU3moz2l3T7mO
WxAso5TZTRZSDpnCshLfwSos/GCRyWOg0F9XOwgDXVnPCZkdsi6VMIXmApsPhQJc
9+01G7mx/HXdaplNnYAovbXXQw8PJnlaLng4NQNW/Is0qpR3tR2leDapDu/YUB08
zKVOHl15aLqHihNRLTgQ/IOrwXsd6wkNWNYuAPKN74nvyNdOpNZRvTfJp81enWdB
1wRlN9x1m+8wFwmUu2Xd/lPdvKkbMZqFF10/mbHDLLW2X4tKOpstqyg0p4I607ll
ARwhl8gA330vsfgflOg6pFes3R2iMsqyuLoh6LRn9PPSB8aB8qMRzY7odcOBNMmY
psa0otD5djuF+IyhJcK9KiZPFE63x5FN/AcC7rgWKz7oEwyQTUSOW5N9QM91uXbK
yJ+W/Ez7De7i9W+SrBm+SppweJfLK/smzEoC3b9UbLl22bim9444fFc5iCf365gy
txS8WO5YGULCdMJEq/wFwEWdiYKpJxMSE6+Zww8jy/lCfgDg3M7CW6VR1nKM/U2Q
x3McOXLxnPJbyGRCGmQiWlGtGQvccwfBE8+89rli3vv4q2rey8y0b0RcQjDQ3a62
c2nWp61JD0EUrEvq5VBdElKvGbA4j++KLNnKL17XiJ12GBgyYtoL+fjsQO5XN9mS
zrBctdL+m0Z5TpalXKYcY5oTxJ72Zj9TtIP42Wm5DDeMrjjIReNT4Y8f0s71amkW
OAwdN1RL1suT21Ja/d2rhHSr+UozcUEDj+weTzzUXHXEsew2i4cshmsIcrTP8EEk
LK2ykvJp/Eds7RLSZkR124sRXIZzKX3WkRAHgUIPUT50J6B6EMC5aHAZR/DTzwDH
4/kjwWkn+2btOccyffjyysfcZNGYbQx4TXPn2r3Ti4BHYcrYtRf5SasAGci8H7UD
ze0v1Oe0/LjCFLOzSEJ/5OFimxAT5KAZhgkIOybgb5ziyKSFSJ6FylloerpVuUOF
v0UmyVcZMXc0RKQfQ9+2HyPu0ruu6pc0i1BjPddzl5dlqhQpr5PqLozvGJXKdw7B
jC+BkY6EM1op2lK8HGjOPrYIELfR44H4ck4+3dmcZPyNMlivE2L6f5qn2Tdwrufg
3wsvCJm+1i8hQLiY7ndmCIDQisiNltUvxromdH9l0+2Ab081wdUG5zCHFffz6eoj
WIg/dEMphlQwKeg62mAWxgFXiGeXuApX2Xt7EgNhmP0x6NMqA8fNfvjjFbiDTWS+
add7Cs1sA29XSpm8zQrSROLRklWMnT9LFmCe6b/Ujez+LZdl2xuFDtp4GxTIh2cP
N3CljPRf6DFumQXVpCVNC7Z7VAIzii1jPF3FFG7WpXgfpjl9Hq/tjaHrjfdt1EET
wDDFGtciT1QZF48qkMSb0DprSfzr7V0Al80HWOOKNzUGYaHzo0aJc/zw+5ipFkGT
QSb5mChHDwcUTd28ftOXQIYtfP4UyOSm6k+8VeRiZIkxajtb7pu7rGIfYMGNExdX
+qEeDKuAYU6Dk0dSVE9D68eyvMjF1WnofNA2gHvFiwDhN9KBsG4UObdYJZAP47Kj
3Sx60rcPQoRkWrzBOvKp3QNMt0jLYWVVPXSh79qqzg83IcTOjklNzyzW9Jgb2ys7
rGjHp9FGm3bXTJDmDCmINS53mVGt2zbiWa7SUPRFyw1vxNqMm0lA/2vidQwURYFV
rVPNFQw1LtP+nkRKjxLd+Mbp9/PSd5U27cfyAQ7dFDdcwbXVjMA/5moUQbg1eGM6
0eA+sq5cz+MAFXvqUJSTEX/rJkO7UrCwosf/M05wWriXPN/DStPNji4/bMLec6/u
/Jol6/gSYomrPHjK1Zsvd6IoSieMWPPpQleCuKh9vH17cYRfv3yRCII65+c/6MsK
PQsQrSY5SVYKlyh8d8yiPdZREVmznLZSh2t75jfP9NTaAfnZPz6Fv1Cm7RvXp79o
iGQW7DKcJX6G+HWryZ2uAWR/QoHJYWETuJMlOehgl8q8g2SZyKz5p3xqbEvxD3m5
e9/xTP3S4VHPOW38CoQmPogQ6vp7e/7tbkGPX0TsNkAX4eKEOAFO5gJlQKfZx4bx
upU0WeUbnoNrhkAtoYapIEP9NQdHxaJyjtYSi69Poevj+JlH10yk1gkKeNn7BmgL
d495UV1t+dtQnMrdX4GgsPwkz8oUuHNPdYlO9XVETMm4ekwoACDLL2DWUExXImc9
zP4DgjWkOFjloSvACI5kFujxydJwQ6J27XoW8960rzOt5zQ9I4lBXUU3onaEnPKN
F819633eD/JVaxmW5NcZAJoKL1I8H/AgkL9NX1rkdNIRd/NhWpat/7vtVpzXnFyw
/OxD9UnLKjffXT8aP0IJPpQiAOsgaC612Tvs8uodoSb7oKa+YefsBR10v6G4Q6mh
duvitkOMG1PNLltuWMnWNioEvbgC5J1kGtOa6VWnRycBrDF4wj0NMh38JscmAhnP
/Dnp75VX5R7ti4ZAI7Cxgxfmcn1NqVkHrqJ4UtJsRPEldmYTx1A8tEwFDS/o7pVA
kspVU8Vpf/kvwqohMH1cVImXnaSH07MkhbB7wBG6HKXSqZ0v6wg8Erx6n75THx9W
2saseRwH6YwNbki2dlf23ntQMlo3cNMtIvSsmalyBEh9cxkMnHYDndulmOsRX6Jn
XXoooS6n73HAnEfjKhD683bZMUjdSYP7wG6QVVhZ8SU1Yq7lq+J8NOYmEwXoyzOE
JjXvjw2gJ+BiiOIk3WImpf5TFQolrvYHy1S2XpJbjGRtPY4I6IOn622bVRiJ1jZq
9MUij5BaSDEbU6EpLCs4PLcjJIA6HSfMcxacFSdlXflGJXjGOU1B6+eTUDzfiuAb
d1iseWZ+QfOxUZ0eU9HC00l40Tadl/cHHAM7iMxoXw3cZ2D/VpMInMtyBdOA49fK
Uackhy76LRC9Fsn42Nt0ckYrWslKU3WbkpXxhT4hrGQpnmJ6L3kFrRPqJT2TXZSe
ppEzCP8atF69RKkO9TA8GktIl0UF6/U02bQGbrnU4DyTbiabAdqOYkRtlTgm8TuP
831f2UcavsB3nF2u/g2KcHgcpn5HEqZxSFsVbq1RTX0/n2r19ULdwYQwOAqQrqi9
Xd6X/CR1Naj1n/mlFogZFACDoYYdCF1vAWUdgmNSKKOfyfUWIuwTgDLNsn8T4tZ+
P7qfHSQhfv9x7v2pkqN3BBah+l03Xl2IbhcEJ1wCU3WlhXPLegVZh5fpgLYcVXLH
IDtaxuxpoM8PCP1Jp+8tWIyjMq6C5P7z5CGX/rrVxl9qRagum5BduTilwc3390xL
k1Ak4cFKEnV3kSjHY1pJfrujteL6JBDda0v88iyiHr0CmBWwtDxfFQQTLp5AUYfV
O/KXLh8TfjKNAThQDOlX2W4wygzQyL480Xb3uOVU0l4RMze++oKnOWMT/Nk9gw+8
5JjuarqQuNVVxPv8yL8YG8wrlR9mdJwPScRtVXbUW4iZcNXIDYi2oW6K/pxsk99E
hyKZhp1sHbpRkx4VQ3MkHCsGT95h/S6A3bt+PghVuwqj70JIEeSkj0DSfXQBEG7J
Zf+QJOMaprMS3Ej9PV8j4rhxbeMP4I0h1iPWSfv1iU2KkVPOaaQNja6jZL949n/C
CbyHKUrs2yqmdJg5V/6dNu32nVr4eOT+6PdsYq91Bfv2F4TEsj8intslEvVOLccv
6kfYOqhfdWF40b9QclddkA0FrBQuAmXV+9+LKkqxWvT8g6KPaB7rJDwCxXWdP1xg
6NBVAxrVCsmK7YgOu7cZsCuf42h/G3TFsSttaNsjZEv+p2pjbF1etPE5YAcSO9rZ
EoI5syK8t4ELPiqyrO1MBJjvfg1kIiyhPWnNb8+Td66trBfSj9qQpnDW1wnDxSB3
Fs2lzQyhq91pyYOfK160KDxGuy4jOMoiESUMHc8AzADl9Ny1L3dwiQMEdFXhLXi3
a5LAE5S+zgUjjkCAQv6g/XnFdxwjOefcRMoW4LxAuSAhXS80S2kSBNRdCpv2d9sO
TdhPmBCPn7vrc4O9wEb9YXZmA11fKKNP27mWetmaxmBHwT6rzQIhOWUMU4C3csVT
WP3y6eydZeaBMlEDVeIB+Oq25Bw/X96m5IEzle+Tzna1YIwU9jcSQBtiWzVQt9Sf
AEv2ZbSnhQadHUg/NGP7gx54ecjtVB2q+pSVVviVzu1RvYuNqB2A3d7s+O6Xq85s
e5RGCl9HsTJ78yuOTRp5FIfD8q7p+mdbgfBXXiJBZU7//+5erWczMPX9p8SLF1vO
Ktt+xQrM0G1hlvQTyV2qRITENZOBsl7HBt2Sn8Cft7xaW1tXXFiG43GoobeiyRlg
K3+vpS4+jvje0GkGrgzm+1byaphT5BsZsxAEVR1MJlxTPDDRrU4xMKZGuUBQ40JQ
bRIG8JqjtwK9ZulyPhXy3F7HxC6VSnnBPxwZQLy3GQKoX5p+TkwyT3KZiEJPyuKJ
WfAWKzTmXNzhPeWVBMHqiJEkRqiVusAEqGlWMns9YRG7IrgumPMXCLVTuAq0RoiZ
OsVYqUwcZ0aYYk/UB5gKnyGX4X2akU2dFzZKbRLRfLOqLZYbZDNfo3U3CHxc2o54
8ByPvWDepK19UI1tH+4cCkwS7M557jsH55q4QbyVJ82kvOxeumyFJ1O6940MSVxD
RlIGeGWiv3TmvFG2oKWW5tfKvohPvf2bguK69GrUNqBYvYYblLaz3JV4edEi6meA
/eaoK3d4VwpgW+9f63CokFkzX439uL34M7l5FE+VRoFE4naYhjtNars2dcN/CU9m
qQvQL3R8M5mG5bPjhhL9BaT6tUDzvoMy0hr0Q4lNHUFSZwT2QJSJPnovj8q0lWf8
7nRFW7QKe5Kh7KZexddQaUngTeNTT517STvuGTYiZZoZ/bQQjGK1pcudyG1Da0eG
Bq9rSwZPNU957XnDauqgA0kO6VeIE/PPLbcFnKi47+YJ+qQ8b9WPSMknjESWecBr
sVlmJYoggZd9KWpS7V7TQav0ZH9uBxe+FrC0iuM0mVjrNcfJ61h57ymLfocFdCGg
uiSIpUg+phktoVFiUOAcoO0Wg5Cqguv62lTu6A+aSbL8zxs4ZOPAHV7Kuzzxx1NE
zgqi1xnDApCMcIJF6la8Ill43qYqUvh8jR+hVOkyE+P0Rdl/fB/5VMsG5CXo9O5k
mc2DiO0scGWDkzsG0Q154xKZFyXauMD6XYDPf3Wf5XJ2Qnc5XX0zajhjQdTsw0Rq
JPhWAITtFSEgXFcdnySHMQp+J4fVFWgaR0NqR3Bji0Hw7wSnzOrRJxTMiNLKL2cp
lAsvzx2TvGUJ3RO2Rj6mkXSParhlUXcNwVsyZXzfOlTCay58KbN4q/9T879zSfKI
K8/xf+9KWBnxD4mF/hIY9WxPQwj+f7bH1tRJng2BD3FCzFinOfRERRn7UHMA4DO4
XKEb5OKVtF7uKa/i0wCLYtFviNqSzx4Eno1ibzfvM+iGL7kXdvUPBSs1Bkd5CAzO
jh5Q7OEumP9vBYGhe2B2rZXaVOuQBTqkbIOlNKlR7ZNUTmaiocAOCpB8BhpkFl/o
g30Oa/AYh/jqb5/X5B86vxo9wfc7Vo7TjV0sqiTjJ9tbKPGaQTfuK43lC6zY1ERk
AxscyVfOgyKLrndwfua2lkAfahC0CE70Y6lxYPNUrG/1Itv6s0R1TWQ6QMAMukf+
2Y6nSSLlKJgJIgoSb78kTVTzZEDVTybwYdBS/N85IX+tW+OxzEhEp7L9PHA52iAg
sK8QyI3G70njfBoLGlm45zfLT+J5mxvRizILujQVOnlliOlCwSUqIVDTRDheuDTb
+AI7pSzFMTtky0Af5yxogi85VQwGLOP91W5H/IIFZcICQdiuOOpa/PfSBFiw6qBk
NBVnqIKKLZ1lv1Mq0x060wtX8qoJ0WwP5l8perpl2e9DjMQxysltprpBGJ5QF8vC
jw16P5NcjxLe9OVlYytlbsqMcddQg3QlBZb81st/dXoVfvoF0oJIt5YXUW04PQJN
qEyqQ0Eu7n4BLArh3Ez2vCfAjzWu/+uMfQg7mwoEieoYHjSogJ2ouDIvo/DfmGOr
hdZbz2QqerVMiZ35Gokl6MC4Ect/QdxyXYfO6BZQnFZeoLsslPhH5sRZIVvuKDVj
n3kmIfuAwAmWOwQ9BH9+qN/XPQ2VLoB+cw+79C8/ZbeYJRBc4U540Ud/T2XkEnjC
iD1BVR1ENdNdxJd9lkk6pMadrxD4f1ED+tSHPGgGBbFBVepvWvmWp9mwp1NEJqT1
RD/atk+tGhyIq4i+VworQ+MJzrBoHt8CywmrsvJCMMrcto4IThPfdA3EkZ1Owsdw
oRkqT9oI5PcTuvz8+eCco+L8J6s5B3V1ygqMZorhxbjiHCMcXfBkPBIKs9jmuhRM
NBDHEZKwdl+W5ZqsYHe0A7FqKJur9vkQZEGeATtF7RH9GXsmmoF880F52h5vrdh1
HqqdIlVMKH4dX4zgXb5QVyV1LXqm8N0QLLXDbehX8GFf0gRvRiGd0UtwMCc6nN2T
FnoF1yhLDPJxSHSxfGbvIGHpOYa4YkZdRkFkOVX1gstxGRo32w6oEBNdwTag3Ed6
7STY5Eca9ZjLH+Ly2hsybFA9l7LUA402bci4LTm3RfcQaycLcVPpYqHVd8JvADja
2zd4Q4dNfSjoarix24jLSDlsTkqrBKw/uw3qEWVEdLbMhqYOiog5NytrtJpmel54
rxeGRWtgOz9fqIMcSYzxGkfdu5f/GJe+h2tI97di60C5JvZ9rj2dyu5FWOwNLOfI
p0Co57dhl/4Fb9Rtn7WHZw9/PI9UBv+p/2PFG3eco8y0WNZEmxtH93PSs4ctZQP4
UyG0LwoXq7Hf01JRur+vjccZWCFwi+P2xiJtA/PDfX7QBGCMCM95flJAxNpnmcLC
208sZydVBDAp3/56xJZFW7AQHjDrh8o8Qpq+AIeLiD0PnFQvfHkqYOdXq5KzH92j
wLP4yQuv6Bb1IUrHPRdjoY85NjlwgxzO/JqZAFA/B8cHGKk3SgYGw84oOMEAUdcp
jUEi/gRHN4909yVEByiD6J4uSHOoa+MMyytPsij20csfoWsmmZvwmWYDKD7d7HGl
Ezy3HmkTZK6cNORj7hBlPTFjZ0wgeEW5cHueZ+Rnb+VUBr7pqxfWMjjkHF+u+mqK
h+Egj8WaWHOw96gX7RJ9Ml8RxX6a+C/aizD29EXGo1NzXcMcsFE/f7wiWJeok1if
+0w+fXCTvsQpOr5DneaMSjApNkw58oZ91ELckIVC0/A8kRq8GDaQcERosHq/2rHZ
VyizszfqS1cE3Tm12l3B2EQYoZZufEaQvE1LMsoddCI9nUj+qRYXZuiKpV9EjxRo
5ijSte6ZjN/yAxvjZjsvy4PBjZJvw/O48jRlDYZHEQ6bPU7P3P6gyuxo5PdLqtk+
jPBIKXDpe9z5RqU94RBxWFDTyC+CxrYwbThGNj3SaL4Yc1Xjg7i6JPMSm9wBl7AT
J1VCAvsDvtYOXQyrD7emXDlHcG43t6GBuBhbHhUnLYa8eTsDyAx8aSZ1NyAaXJh5
NYNO6hxN2udGZW8gJnPEJtHg99ZXuThhm6YDYTNPXZJQcGfWjtkA89ID7HpOQcTO
oZIALA81cM1dQZm7Xlqh45EtpCo736BsXaE3+lgaunDFS6ZQG6L5LcPy4Up7HLH9
BLF5LsHkeC2GOBos2+2uXyGlddUi2nFIrEhVA+bUhBztfcGgn+BMxz/pkMH3hLmc
Q264QqVQFshU4s6S2azv5T21jqndfODPvRxP4jytLmJA3n43bWpZT/kr/H45qRM1
a9wfHpd7Zv2eyiPwqr3mcVNZCl+NmUutp3sDch9lhLWovfsGYpDvO0woHpyIE+IS
EIQ0BkNHUVU7/CFltPoWhOmSHLYKdKs3uG3OdAtwgNQHDssWv9FNnU1X3USQsXW3
N7RUluxE2++f0N55d6pwqgQ80Wrhyes3khRNjCHRDqQUv5CoKrLBU1/32N0K7kWW
cbHR6qCuFaqstibYS+ecupSBcBKdvwD/sFV9h5zVhXdd4cTJnKY6r7npnpiSw5cs
U4TIgA4nglyGEb/E2KdEeZXqVfIzFNKOmIfPaaTHvDpX37SLwTK99ZMKwvUdBu4M
5jtD9dngARYn7zK9rjWC1+lXNXyg7YI0x5tnuunyDrPAW/A70fL/kX2k+GXDfp8G
yMw/Hmhs9+7KILDZMZvnZ7Pzyncun2EuDNOV45Rt+OkbPm6wLnsop5hAOZ5igI+m
7wDKihJIfSM321asQU3HZODxOAj9hF1qmwu8N/JQjhOKz3f51yxx3nPbxEXnAmWS
h2cYWsG/7gNxQqJ2bJoM9qB5XFJAKtrdZgOcjShFdN3kx/62eeSIvSMpNU8sjktS
Jc0lhf7yulepFvPGgz4U+y3DUgHLXgq1o8wPAVxkaQBm2k65VqKyob3xWfPWIUdJ
yxrdrzoVHSJtAhw+IeC7cChvWTxBJmQZ++WdzB2nMcE7gyFDQnhN4m43BlerT3QW
4A8Eiztg+3ybmUwNvtm+HxO9Si7jcVQ6QHyvIo8ZxWzxza0ZgzjZb5gJNUvY72fI
37NI9FeGVKPhTvldZ1f71db265MobQbRwog1x78nORRt5txYqG4zrbgcyFn2zJH1
YP9TkJPX4Fq3p3L+rVj+oru5bm0dWDfNg/CT0V1Rv+xEfdf9TOfC7nNzx2sLqXHR
esVoZgWlPJO5rjIWV+tKN1nYysuINOxLsNR8pijBtwh+wuxj8L3xXUtZMrzXG0yp
IEK33W816r7UXGZvVcxaOS2X8quXRzlyUAMKCq3NRsGVrwp6aD1a72LNMIsanzab
SP8XVSvHPZU5EYN3404/lqBxTr8gV28Vyvn/xF6DcNn4iZl0jgCo02Y5S81UyvYI
GfZxQ3ayYENNJ53UC4NbV2k0GW2/mB9NAn4URbG9RWJAmQdAzg9wjDvuhG8XWRL0
HOBQKYLGMNm4mpUcGe4++o7AC4uF8EX7WincQA770MX+hZ2kDtI9yiq34ZOkg/RS
4rbihYZcl0OE++SCQjvfD72esmaU+I1PxYuT3G9hJdCq6jXm2+kc+2YX8UwsOA4t
DpP0kB/U5Yi/8y24si5F50FeuOsmfGvwZ0yPpIbGSn4YoeKGNmkZ70jihVW8+CA0
TCf5LiwRufyaF5u4AfrUKk4RC/CEDR84ugbh+Y4nDL9+9ZrbM9d6QVj091PWZEq0
OJ6lJZtj7xnZ4faOvYqMwPF4IsNkcpHV1y2a2C9dHoUUMPydNovNfacF4DL7XFdo
nvnnw/o3riyR2C5sA1TuXJ+/rLP7a2AlJ+s2Is9PCO5cKXu09XgdVGhm0rV2pWqX
CzMdXVAt6OL73X4xzV4t+bVV70qTvNjQm1fCbl/+KMksymj2F0Y2x64uGYfq0yeJ
RjsguK1jVQp3OubMzdk1yxKN9MF7Hqtyfe/OX92KBQkrlqwPWK8Aj8J/RRGpv6I0
Xl8nTpvq5EH82tRCak6qg1IpxWTvi5KDibxdAKr8ZZ6jr0/QcbpRvAVDslxUm1sQ
SWqXUoq8mXLkTLxHKIHtm6FoJxARB18l54SubY3nz3gRlZMYXbjvu5Ty6rxk4z5q
mZpAOiB0zOs26/IvOHQKXaGC5iKBee139JyL4WRp03M+mPo1agcotvZORnaLtOc+
DEBhag3+prJculGHMVtTN13BvSgV/P46Az1nO522c+9jDemRA1XpETN9ubo6boJx
tVr6ej8D22muNYD32DlkExT5sFqugjf14w2HLPs4wOWtQ1V22EH4cIqGWmiestGC
pJv7s9teslrdmMHFaCeKxgQtCMUxxVwDEzoUg2vta61rViLbdPOpc34WibmjwHsI
24WKVMofmXBWJQ1YTzYlVTXMZRCMWbIcgS70bkf8Enh7Z+OWkrkJnNUVfK3VaD5J
/XG5NJzuxk1oYbEejG5BtO9Zt2WOmJmN7CIoGJ3elIeZBGTX0He65Yn/yorFoA9S
pNVTWPo7c79KTeeUUmoZMqsA1wXCtI2gbkzvfnlALPm9LMu8IwLsG5M1UXuLqDTv
ZRgTpbA6Bky2L034F3G2Mmku9pTF5RjqHKZPrEyZrftdfoTuUbidw/JTUdXUawvk
12SdiPOgPq4/AuTXPH0bublVaszMOssc8rnsrtsMX4TUsyejO3QTsQZq1a/axx+6
7INTcC9YWH+H2QouXXdJlcKrLfmLyhzi63b6c2oX0k19TikkI9pHhncoGybyXqUs
15XehSLdBqqe/c7gDRsn6Njv0rFbS8qCSNkDNLPGE8l8yW7ZQyUy8sOsSz+4oaEr
4VavYhIwP28Yg0J1NHkLG8s5AVaVOojtQJZKHsZ/vUPhR15ypSbsWdNcCG44vz2X
Epqsht/4b3xn1toi0wMst9Ufd0LJ2cpE8QMHvysjlR5MpQEiVXqmNXR7I9PzUGtj
7jrqcHWiXeWYhbG2CAG720d0sCoXWHxMI+vea+VsSW9dpwYgevUFgyaNyfB1apWo
calwal9UBbFwgymN8ADE2EzW2WwqVzfuaDTQH0I75rBCXnzpQBHa/ep4a5yM5rIt
XBABfoVcxaXK2Cb5uEvGeCkRiHkN8dRvMWaznOQEI0SDeuog1ZgtBUB9/6vinGkV
3foMFz9PCancBf+LKy44kyfFkfial542fA5bcBmBKIYTIYaBlMx/xaBmkneqi8B9
u/mGFfKhZYNFh+v2YQMHvZUtMmycewv+mIH3xG+GxI4xm9qjcL3emOtzt6k8L2up
2xAE7E81EyleriT54rXywbmfJNG1j/MWR15r/IMPZNBhy0LWa+Z7/zZd29o/CA7A
6SKval4/Rdu6QuusHXClBhpvph2EfthUQn3uDn4YiAO50+vr0Syp/zH/rkkV7dMp
PAbnGr4a6znv9ZpDUu0r3vFrlQtixLHqhd/Tk0qShzwRL9KOB4AV7Jm2R0TICNkO
oaen9u/qCl2IM/88XtakiIUtZDNwN2jXQf42H0p0sVH16HUyC7uqB3gmJb9czw/B
eFFuvHITF2vY2b1cZ72meAvZze9umvi/2Wapwgcsf2zK7PIXQAcgGPRo8/GNFQQf
+dRu5YqLQ3+PwVUjaOE96ShQ2HQ5irMKJ9kF6ky3yis+K8WqT7NHMa+6BcGCRnn7
jD5sdYSYI4iFSuYNkNAAOZ6+52GMRLkwUkTUQaby/PJbLSLlzpjhC58nBptL4Y6S
wlJFZqYVZqkaYkMM761c4A8u7zs/zc1BLGLAem6HAmsEPd/f5inSaEnqwIBZ2za4
TG/M6F088+tEvcQpLAsd61KMd388lX1j4nHI6gFt4LqIXuJQ5uCH5QMJx9L1WW1B
Nmuzye4z94gKryOshJT+KEdQ2vj5P69BKrBW7ox8HO2X4lytC3pEp3gQZRCT9Z1K
N3Myhtzm6Q1f1eDJQC0eAAFa9Nw1gZChVKHVKgAz+alD4r5roCwdqa+UfSHkoFQC
KtRLdAZCzRQvfYz7hy3Gq0D/nhvvC2c9MZKnoNIdZJ9tsoT4txGgRw4jr7RIG8MX
ph935hdKU0yBtyEIB9tPgQMWWkgkcinlAcSsrQLg7k7197AVSdr/usN5ruKrj5L7
sYislP0bZvWQDTt0MkAzf+2qYOyZQCmNl/AslWgckOsH3vD4HI65NByF+8XrLgmd
Xc6SdQK0Rkqxd+cJvmgNEpM3yPY2ccUWJ8gWRpRhMK1h4v+J8WbPtTN01cfTEupF
oGhKyX6ugC35JSY3HyQa8PX94c8cLKh41kEZh5u1XROZy3TfZQzrGEIZUX9CSyr/
PNgGVxYwCt4yDJxD62BAqsVyMhMeM9VUFa/RZ159PxRiDVXCTTaQPY7jkLOLjaaW
CQU/A53i+9fyP4W6jS20d2bDKRcIaZpV/QMofCh0H1uuGAa+lUJkjSkgIPm4Qa4r
B3imIECakkmVf3mbo6Spk9o+TucEHoEr3RxXOGG45c1oIpVnCzUfCqLqZEoORWsA
FTB7PbA02k4f0bHbGm0V4zvX1i1ZlIs/ItPaqSrqrm14M/ucX2xBUQ42Kz5uNY+D
5lKaIJTOAjht4NAt9DFaip3QRP1Y4u5o/kmkAlwMNvzEWRa/8TfbrNDz44Tl5I1c
7xj3taQQMkXlbIg9zNldRgidjQ4wPaP3GajLQESbMFnJeV5t6BI7CVB+imu//Bmz
w5oRkoYhG/CZroHdJeZE68TQxQOMocwbbt0D7xLZxcOrEsxRaYyu6mJMMOazaC6+
Z/PpWXai1Crt4pd5CbuoSGvrG4Txk6HC+QBUZbLuOWThUhxvosZAGPt5rcMU/kej
HJFdD7ciz2SEOC+G+VeaZGjLsiXFL3/xwbbv4h5rARGcGvxkCOycCCjXy6ockgiy
nulICb8mUs1J4wv/Xh+soVmXHoHjnDTEwHre/zP++A9AVI1PshAHb+onHsb6nk3V
fMz624WhHo611iMl8r/W2X7RjqUz9Xud1bdv/mRxKv7HC5blny2DA5ck5PJ/ZZ/w
9qaJGUwl9bCNoNUtcvpBvh1iYtA2eFiwYEyUX4yNnLSupRcs3u0kTMLlWk4mtEIH
8MuASHnDC44lG7SsN5uFq4bhTKOifUKmBHvTAWQ8VrLhO66nQJtm3gM3ivoqJP4N
07grj+qDSSJg05auW30LPrXGVz2RJNcT66tD0pYM4eYVCfs8ZPE+uwAlZ+z3mYKB
P53da7zpxbOs2wUPDzwQEVn2zQFYo4u2YKOBFhIwnMbZ42mWk/Plk3mZGEPXBe99
R2P67s2vYOhq5IdRJQYCzuCwdyqNpG3gWSI6eOqQanlazVCLLcxTk6NqKUrOUhMU
Ig+3+0//2bmpB3rfpEU4bc5bMGhujrVVhytXKZLJC08/CtleKheRtckP5bbRpFul
v6taDD6RNZ/qvyM/hD4gAWoVIHrfLVvA5UBxx1JVmmf2Vf+co9wBaCCfTSUPnWdh
noYEQLlvQvdKRSX+VrVMHqoaY1ABGWsUhioCxSjiEZzpgVDZmXEEHZvH43P137CV
HFCYa1s0nhQBcetESflusTPSca3dSu/jQU4az9w55XxOYsaC4lomvoHgIihBpzu7
EyDA7TJeRAQExtnV82OLX/+WHmRHjih8IccwHsfKgNfJ3L3/GUR3/2LWg7x8wKNl
S4Z742GjACpDNuwVwEfbidf2yvaJb2b1I3DoVkIZViW6CZirVJUQiBl/e/D5aQCx
5OulQNIFBx5k2f3UNwOGOHp2PtkUxVgGG+CphxxqnP6EniSewR0BE4NY4l3Z8ye5
goFx7BjefCMP+BSzw3hba4YXutDDJ/N9luZR65vMbU1un3Kik2+flwRk1YHGQDvn
55dZD8rlVnYAzRAI3eqSt2pK+PxqeNccORJ/yf+QPVfSsPyagwHXLDS7SoLcCzMP
yfltLtRAK8BASTJOou618mPzFpZZORR/Mtf0z9g7uil/ccFYN5s2ifDG9pD/ecKZ
vVUrWUIl8T0DFBK2C788E6+yoX2t4gWU2PeiMBwj3VSjYjXA8m2TDt2EQPwI6rOi
3ZrdEbegKBX29Z4hMeQ3SpDXnjaNiIvX56d6Ld8MjTZw4CHTlsheg3JgOMj06Knb
S2KKl/rrfcGiKdFkS0mQ/P3PGy0sBQuFIxB/Olylu+qVo8uRw9Oo5fw1HoTbl5T9
Gwb94KO/GCLoyoPFFijSM+KItGhhjSQAQPohvKxXCOO9G4qGGDTs54mzGSyunP9G
tEd+t5hiZXHh4e1pzWOh/tF52KOPOoTeoP5pu5CuFgS6rTl7GuDcWHnIaKlsymRj
uHxl3gOJDoplNbnfYpVr7nwngy5osAnvT3iiToXv54ifrT9Pew3zI6bVD+cHUqeP
UFc4F64VPFm0HWoD02b6+YlRZcRuzTsdzC3RF2a/bDdRGnxMN/pascm316fTTS95
fH5YpY7S5b8WEMwPivMcXCPuh3tb1KApkG2SwHSI0LOZGbQOdb6o+DY7s98cCZaI
1ZaKsubXKIMaS1/tclntxIUM7wT943C03FAlLeKc3MSh/SwWohzseD0N6Myw9Dqo
lxViittXAlk7WneZJimM9U7xO4JXIUV+KlnDJj+1O4WmlJWcaYQ5ON3crjRaIWNd
S1HLy739WWVNpbImwVuUvFRGxcy+oaWDhgCoDbFhN0QqFwfn6/25Iwnw/dpa3noA
D4cZ5/reYNxNCLuhgubzDFm+riw+xNGPslU7PKHjgBBN+Z95ohhGKBQ1k1gdO0ES
VMReo8L4AAGAY5u5qyzT1DlMF4H3vz265oLgAvMUaMYZXodLRyCbSVTtyPnmgtWt
yVlaroPlKG4UmR6X8mEkkdBSnY0AEQtggutTRsKSIhh2023IJzz34EAnqqzh46Sr
nwP7GokveKVGVP8sj1XPndrkXFtexX9352s55HzuU6U+unCoLh5lWnkwYPIMP2sQ
ce0gDa0dR4FIoh+LqLcUYUuSxgkBxsgr7QwnLhyK6+vlJp7DaM3nDixv2UKDMlhV
HxTMpvFhSj4Fp2/KTnqS1ZEDGzfPr2SBr0RUYPA8qBL2QnHyG5afwsYo4PAbyOFu
IJp9ETX/7DXcunGdWS5PIG+dLHmN3fMezQOX9VFrWov33Ks7Q659Q8foq827CchM
FYLWQ0wAcZYQGCndamCknGie2G5IuqxgQl0CTLtWUZe/vsHkgInanFM9PM/iBUDK
LJwpq5tJt6AJTes3WlE4Gw1uo5HAvy6YZtRPqBYwHiydY/3P0E/x7mmgXTqlxtFs
BxVHz+bb/ecYE+3xiHoTYmq3jX//SXfbClv3hvSZb0CKIG/m/HBQcZBLAvEzVCiY
XPdIH0OUSSjd1empgz/IhXi88+r81nT+zPCAB/kuKHS/M5gA0Wt2cOihHpGWfXHN
vxRzIw6Colzz9Km8MuBrYSuwsrxY2S/AMdjIN7e/U4sr9+FQtFXGRn5Yt2ysimBG
jsPPfk6/A1bb9daCLHI/nXiuDQVSC0yNjO4/OKPO4ltEMYfR0WwkOk0mdlHfEvkC
c1o95Kd/TVnctrbn3PmWgvhh4Ggzy3veop1YC65kALAjlqxhd4F1PAwMsI58iweK
IeG71QMBp73PayIiqrUUC3N88HjfMhAvJahljNKtpJGah8BfGcMe0W6Bs2qkm8Wv
jii2HyzWMh7UI5dxgN6ydPHGH5XjNM2CapcG6fplc9QcC8EJi9ucJh/Pif+ZaGmE
5Ciijj/AkyvkNQhIdfWmjk4zPDRlEifQpNh3YP6Qx/OhGLzjcAJZ206Edqah/lO/
6DSKMr91ha72xvpMkq+CqxmXP9cKb3L+yLiG47mK+mdk+Y9yu1kLqkBKHxxlFh1w
LwFSsT/0tvfmvEed5eE0zVGDi89jB/PN8WdzTFWRifDWweJfU8joq9hdO9mkqTkY
oHnklrzZDZCaiORN2rhU0h+M+uFrcT5UtSoIOU6B0o682xW1DJhaKndYA/+IqW81
FtWI4Mhac2+V341XYvBYNxFR17JPC3ZFDEXhgvIYJN0xAEjcfMmMZ5kyLS+hpCgU
hptMryotSDSncKJDi3kraxIuTwHKG7TGQ/aXfOlTiiyBKHOVJno+kOBu0yFlMMO/
ET3duDfQtci7NHtp+R6txcjDULtAA1CbWLSP1UMYt2JW7uzHe0AronghgGBwLd0p
x+JMa2PpC/BahknAdoyl7zNFF+/RxCBpHDigJlo04OZpWdkTje9jITSV1VqxU/W+
45swR4e8GzhbzXO+r9x0nkR2G6OFv+7uBBHk7MQhEuSmZH2n4CHYGjdc16faZ0jZ
K8AX4nVHqwXWXS2khGXjNXRjFHaUvY/4e4fFEsbJFgdySC3LS0G5k874/1x1yrRa
cNoFFBCvpW43/fDbZzUP/it4fiEYAuM0gh01jhOJHk5/sXXn2g2Aq61MIND7Ps2c
Cu08GmSaQBFRJcp23C8WaedaLnrhlaFI3efPKw5Gs479b0zrntVqGFmjWqMKuE/R
5FF82GvkqP3PgsOenoxRFfcbiSUz92XQ1SH65wwrYYX0qiwdd6/twnO6wwv3/b3e
jxNASFB1cojeOaOprsWYctG/TNy7Utot/8qbnkSaJ7ydDJL1LkL8CwRcc/8hki9a
7ZsnlU92pNuZkrWG45FQqoSN/QImjpr5DytVBVSHFEVY2yanIflwZ3JgBTcdLxyE
K/Jv0SKIUCgqwdX/APdNhe2N/g2X4LsDlxMXcwZIOHXEMJ/Ft+8TAvXLLRuTgswm
yUQTFzqod9MSFYqTNx39DUnOOUG5vihDFELj3gRrtd2CeDNdZTzit6JkBrQkJ/M+
92HbQTplrdTd/25VOhKloD5N5SHSmlh+qL2qZPSH4MoKs3LwFOlCgxvjRn3Ta8B+
sx0t00wKlJmUSSFfbvqAxiiX2kf3sxwy1ivebQzHhuJ8pU5EEWPgDKB/YcfbKczo
SdMSLRB7NuiX2pWQoZIZZG3m9qqdIUciLUU8acJta9D0nUJPUMEyylQKnbyTQZe6
v1htN+DE0/7FbINO+AoioUCfZD52Q1/bqxcuBsko//4Vh+u1douqOOSc4rVg2CoF
zb2qtkt2sC6O+iBnBmb2p1oRZ97qnhVQ3l48fvSdSddvwvlAjB+iUISQDWZy2EfF
gN10sn4Nb8Qhn8TRIgIj0+scO/2y9H/GmulHgz+yYreiP/2mAlutum2qtGBBsbQ6
FAjml84JiCoEfiR4qr3J0h587WZg9iEEFnQJ8JUqDuWWgKcehonv8zB7g1iwJtDJ
0OKj5IAem5WUDMvgMzsq1c6nu+asuVtxZvqLV9YN8wBXFPqVGyMo/2DtDzYeTp/l
ShjFs1C7A/76vnIh5bcYRFDbhz1ojfFk/ZZLVQF7KdkSZ1gj9mXYHro2p0v2tVTg
buur9v3vxVwz9zLPWhcfsVtGazCjCdl6kpoBRPPG3pQZGYQ5NHtuqTpdmc1fL8Su
VUofFo6c3ksqbUBToyZzSjcDpFx5iHIAo1VRRSzFl/F5ukHO39vOU0vJNBw8ZPO2
+N4nTsIGmlQ12aOYf3ZO0Y4oe4FDofQ4LP9H66/tLPbL07vfClgDg95thYPygwFg
Bq3ep1nEDXn+k1cwUT1QThNNQktnGQ39BCbQPklpDl7Nl4NSoZ7EOsNXfeUsOuaK
entRg7Utiejwhil7aPd7aBkNS1njYFv2TmCmo8wqjBYfIOtZJY61HZzui0VxZ4NP
qAlU70ArWHi4wi6w17bzSy12ScC1U9WbazxOORq2xCpaIZaj70tgCBLknYW8bg/0
l51pfsv8ZW20OKkHQAtnZw1guozfFfISA19TQ3omseu/jnk+lRYzR0Tk9AWS0u0f
27zgjUq/26UZmfQ3SkYvoMi0IQZ3EdbT4y8hoB5ts2IW7q5C0RDLKr+wwvG0Y3NG
AA2CLbVgd1C/5l8nv264QD1ntdg+X+ldc5r1+9CDrFGXAsJoH8N7z09PHRVYmkw4
PgItvlOgVjRh9Fkk4m6v+Fw96Vpra1PC9VXe76R2jBNXwNB/klGLuEnPLWh0U1I8
MLM3gN2sJpK9Iib/Voqi2CBDicgYvsz/VSwDx3Fe+C/QFQPI35cgHCq27rMllfUn
5HW1VhkgjDgoMVmRkbuX5a1ejBh4ljELptvyBbtxoayg3VXAo26Hl5S9Ir1E157z
8O5wBqggwhamaHMzyt3S0FEbObWTFY32FjgYvSEGLU288BQznNAc+qw4yf2ZQKzX
zzUBlg5WmyXGHzwuOesWJ8qCeoJLvztEc7QVCci/4RQ1NJC1Uoe9eFo0OVAcC5/g
vcHZgvp8GCk0fFoCYT34d5KHq/T9MHsuCeHMTf/T58cAgV0npgi0lRfRRq2z1tG3
g7SNk2hLbs36svjvIEmKrXwMkDZbKrxMchMW4SnS/2iGCGfZApOvX2xqi/ZOXw0r
OuulLGkxCX3eW/kSxw2vdb4jiqbFjUwMtErggnf0lkeBfX4WWyVTLoWLX8nO/UU6
NVhxsiuz8gdwxTLj1FFnp0YmfTttPXzLCvC3DKyfN8rqWuVztmSZ52EMAUgZGPxi
EgySfaO7JhKwBd9gaKKt8Aq+/BFoV9srkv1dUrAl6gIx45O3DJCX/A99VSnfL/HU
BKu7BYBuN8WTWnrxSLNjrZ+vCulqh4kx/RbuTV2vE4kmxVe2tIb1Xc0Mh6prgC0x
HxWQKfWLvcNgmTVVw3cHw09vWKH1hzMpQhdgoU10ZZKDtAn/j9ss29ZLRVwslLcN
kjiEox5dY+osijoUw8OWMEZF+aAhW/LaMkoIDyY1KTgw03awXQuWopVvCV7xPxen
UpPHuUu1KKSowXnx+kdmR/G6hqK/wKfGUZgtqsH/wlyXdCzDIvLJ1P56yRBO8J0o
JRUl67Kqg7TZzb6/KGP+WMiG4AUJ9/9sqAbF1MahLJ1yY639SMFG2FZwA7haJ2BM
vzU4WVzfVQZBccLRojMmVl7AnKKXK2RNbJIWr7Ky1tUdwxclFMGKM9O+1c9jYRek
tkj2NAssim7TI+FxDuMKPnZOlDw7anu5nUwocn/lB+rYytUOUJsnZoJkbNnkAsBj
wrxEpXvFvX/I23puBMtYJYQl6nekiCejclF30GzlJGd4MmKnOCktlhE8DNcK1ilL
0vlrn6LrpNMUA3BHUWzs4xH71+6hYEOkG82Xn0jXG32KoT/gBYTChPaFYYFZHWG4
+SxvafGKkElScY2QnA39O+fWEc5w3R+1+KTV6lL8gr4e0pvt84KsC1UbqfEhETWS
fWMT5JPC3e2h/peeeRCCpYLqE6FzcFBSv13iriAvITErpl+IGhKDQlmHFM/nwvvZ
Yq5CPQd/HYU/tFlHtudRXAADOGm85OPu0PywUXxLZsT+ehZlyADtlJ6X7IPrhHWp
zWSFaF4HBr5uugG+7GwQT817DQX7NRoezuM5jhxleVSYsYW3MGeFg0bQXWXAjPsM
3A54tEwvLNI1IbK38jTIx0mrcSpXvYjHI5rYqG0MmwgbXsfA5KJHbxHIE/6SDox/
oLhSsCu2Ja69uI7YtYNpjupvdOdvgrgMz5JzRboEathH7SLB6GWKfUZPPUjIBtXh
NzQVuVzwwrTXCQ9t/Yr9uDAALMgY6bDMdjvs3rc9Bul3WnYdkOJ14BVYRG6aik9a
8c/6TgbZzp2c+oyJEnAZQO0+9K8g66kKrwBwQAII4BkHJgARS2+O0PFvOH9e9aCY
FHY72dr8Wk4VLyg2lgznsn2JehrE3Uxsu8mEtHppVAW0ynGTWQZg3DvWZDAPI4qo
VOSwmGgzXSK2wXxM8X/k6+hZQqJS7/j4LKHtkNlpC9hMU1/nwBUihERQhmAmBifV
zuGrutsE7sztD8Sku1G6CTpzMnG6U0SR81Hq1elkvOzkmVjZnvQxxO3hJu2N5r+R
Z6Nlr402XRjGZXqSoh8esk043cJRffvLlDdkE96R2bsS5rVr6JaPnJcn1hX9Qt+j
JbSRdSL5ZFXQa+aA40t4BJSbFYpvqRVfazwH/90wgyS3tv6UnyC2ExiHnJiC2AkW
UqNMe/XPBYqJpTq782nybU1qAL66NWRnKPSPnYre/kqdBXy0ETL3y6Gel1FnbXrJ
zAJ/1lfhvB2si6XP4gSHUy5cLPEOy59WWEnKlXdHuiru9snYc08FLqUwPqkZKiyL
UOM/NNZelPxD/Ruolnavev58PvSqkf5QtwZHPxobLMCdqiwmuvAQoX0vfnfQ1wcD
vHhi6Iq8oMSjVxeF0VOKJdNTKF+5CbxgohnezlH7WhK6jBIXg0PeSaSTR+d8KB7f
Kd3Gk/E9hpaRxT7/Sj7tfk887pWjqPLc7EvGN6zSlLFju1CIs72V2E/qWrSpgaq8
y1x5AuinYX5/N1wK17oAqoCyPpV2IPKEPWD3OaWg1sOPxh5c4+kCJBfvwwe1bB/x
FfrJjV4HbhEbUL8GrD3xgeUshRgo3eDvFYlMWl9BkaqJwzHeCXb8W6ubIrdt4YFq
7MPBX64B+dPusD4x5HIAaPylcLaZM9mFsio+wXYdnpPb16w2c/gEW9v3+wYJ/9hR
5c0RoZVCF8UJy9HKrDv69EYx8MOIqqz4nLyB2GeSMxHn8LcIRa+QECWu78Di4kpS
kDoIMgi96OLGmLw7OmXHWPhZrDGFyDeWykMliYLC2WLYn3YYmi70Wi+Tnce34ssX
N6DGTId5CC6h4DpgQiBquM/DkCH84uDTlHL5I5vmOLw+DGXBnzn2v9sbfzQ8hqTi
un2436aNI0OCDElWcRy0YE7XdshZ419qXy9ldMcHgk2tt/m3/W9m0JvZeJLy/C4R
g6w2f4SvjBZbdFjQcw3qEH8hRGBd0cZGRZxfz6zofavTbsw34dimiYmRGxBGkYO3
wrM0xXoVo2ukx/nSh55kBFPVZ2Qvo3NsaKMEwoAODvykRrussZEmhy8LzqpCUZ2w
YOaAs6Qlkma7VDNUrCwLSZD52kqTILOhtEcNpD8WzikpxhKeAZd691VTbgK4qNOf
pkcaHXZnipJtRvT1seuN6LDI2Zan9AxJsVfOVnG66oGFD9sGVBK8swSbayS0LYbS
pRDOw0Zq+/DTUTXnPkT3LkNpfIggrb7g5EG4s9/DxN6heDV7RkTO/rV3fonB/MjS
+hvunpHIHAOt2Le7OYHg86CzZx2/cfnSWnrH7sdWcFKy8F/tBXo8t+r/VpzJZ+fj
duUu7lJq4hUQfe+dsdKDiHR/oRd3aM5ZwdM9hwPnWl7NORmFdSeO7LLUhYUMTOH1
97JXEZaUwjkXfsRvenYRHhozbwIh+AgHOWnVO21YZRT9wA9ydx4QmwNoMgHB06uF
0JMoXOw3siljjIaE5VjG0klnu1iwRIqyPPb0di0/fj0nWptVEhdi1XE+coRL3pBM
qgNnMs/lbrwTR4B7O3waL+EvYAP25sWMH8lfqcYl2bp0dgIbjY6F3mQHrA3KvoNT
9tOo7sNfT3NghlBH9bINWVDCWYp+6S1yC+Uvub7xW2Qrfpe7r8WjP6NTxsGQX8/p
4Y4JS4gNEsIgxopG1rgAjwaI9yKkZ9ZdfY6td4VHuWJpifN/ceDxRYgtB00e0vYF
LG9iifaVJxKshzUcpldcnlbeOzu3wC6s2Ra3FqrbeylvfnPeC/walh3hG3rMeHOu
0ODYs/ZA9khSbfnsgQHDPt8+/vgpnxsuBlezCZOo2jcbeyN/t0i5pwydN6s84SLQ
w+pTp2F3nRXlzYe25MuiB6DeYhtWOk/Aj5bvy1AmggjfisHF0LTQNhoS6CFBSzwL
w/P/SFN10mOMyN+L6ayVLMJfQDfbLtKehcnNWJU9/FHA5FUcY3jeTAE8PqZXQ8zZ
w7EwptfbziF4cLvpQ/j/CSKC43zAUk0IRdr0hIoo96F3SL9eaqAw9bNDZEGvyzBr
vQJ5qHvd6dyx1fVmEpU/gvvMWSHgYBoIb3+exhkVusO3M3ktfS8OikZuBdGz/8Qj
gBgOJvNdcgxR+OhrzCZxi6xmSeflGz9zg4V8h53sWWiRsvSgeENoXMtZMCxTAlN6
l3NYmJuS8a6qNbcpxAs9GIKhnaGpuOnXB994wOKU/QPnoFKjFrUJUuTnG34kapN0
H+mHhZ+okv7hG5QBcDbAJfUF8p9fT+pYcdZgesKGKuQowjLnXvmvUo++dlp5B+ei
jQXWSbIJ6ZoHvnAduHulZilAh2yXbLJ8doNrf9rrFlY40wi2PeHR05dB98U4qITT
xTj5XZiCg+I6935Vl7b7vZbSdrGBwmvsrcZYCIzTZiC5AuAzmRx//pn05v5iRowg
o9OopJ094+w2DV1WsyT6b5Cu1YlWypMOyfVs0BIKvukEUQZu3iAs1qhegsvdVuiU
oozL8xYim581tTcAH4PYDn1v1fru0/bmWoeRe0z9FwYyh629N5QmX+IMAlLmD48m
r/huqtBMjkabdO/WIzEXVvFt412opWeIzKOlkVEmLHQGEUTnfRuiQZ7QPvsxM7Pj
6emR9MSxIuSLoIU5ZSnhmDiEgkQ0PyXJV0nZeSzmuPMa1OOpbRgrfWbKuLYA0yVV
Z8WX3at9McmymBY3x2jMNfzl7IaxwoD7DegwgZyxL+TwhQCfQQk9oMMD1BhUziuB
xQAv6FkF6EHrwW4yOEYpe1vg8KDEOb5yRqNd5eiKZ1hidFDApdJ7jddnDT+wBRdk
sYXmlL/2d1f+2ooH2ecX/YFEcJzAWV4r/cEhid8qvqNJHtZ8lxm80vvKZd1C4BGz
ovn8cDDMQx+gophA3QVSrX4MzXrS64t6mx7gGoq+MFvw1ncWX9FkIPH5eu/wbDZE
/nQW61wQwD2TvmNEIR1Kjb3sSb8LErpyQrEdOPD5HazP03wPwY8OgIrjCnBM9My/
WPzPHNK9DpNAmsbw9BTRFcQPS0bKYAms9TI7Fh3gBtJN4rWxQCjK3n49TXWNsdyx
Wn3nUAOY8gDT9uKTs4bcP89SzJYRD0Uq02Inf5JAZ07Uy1cEUxH22/+wlKmZnOHe
Bue4Dn43rie/r+kh1FW0BrF1v1eEB+3dW7RScIbADdi3NdrypLpQVY2TKMejNOh8
OzdTxR99ixLNafSoUqV3V0BARNTprxxsWQbRV1Hi9DFSU9mjB0tSorHX/7qLMvUN
7RW77hcLpAtuCpoChhPGeHy2VKHrK6kP2lPR9a7dQm7T99lsB/pGIsvfugdlRfNX
JsPSxk16cH96CW/eAw8LWbI8ZUZi6PmCrJmxGFo0EgOl+eg6WP8+RZY+VsY7eEt8
4x1SK1LjSaqLb0tVIoZ3HqanqAsdPiNDm/mkdszRZLae884sjXTcVkXI3/Mf4awv
pEwpyOkk8CDHg0kICPpTfCnjg2nf4KRRDE05kzP3s9LP7/Y+yH3WvHTUBzHC7AZi
xG/64SRK4biUSC2+QfqyRJqePQU6Cdr6n8Q2XN3cO6LP8BUovj079PvDpcRJuOAh
THH28pAHUQQd75uuZAQvw9W0CzTOX0EH98gpjdLPRhqdP/Pwc6teGqLSQnbuoykv
6dfgfs6BqT4I02aH3sGBohzhwHXw9BkFOCN6bwEJp0yAz+Jtu6ZQmeH/rBZf698j
slh7oWZfRWIHXcxAy7GkTbE6sqP9zfSpibxkMBq27RzoM56hVAVmX07ZqDmVN5FM
nS2tnzZ/1bSomm4k5Rxt85Hpoomvj7n60wqs19dw470abhm54y8lF2RpAGFQT/Mk
xm+Yw2fSegONKk7A92Bc1Hvs72MXrJS0Jvf1piWqSoq00UIY+ZLl4uSfCeBRGiFK
byxRixoH5N9Oo4MoKd6T2n82sd9F986qnfUZtpebPVE/0WbfEKnaoEb/p1cpxkrL
IPXfG5bYldKZwB+IYBHw1T03ztCaQyGMZAjvh0i/JInJKVzfokUWePwgZNh1L5r+
PKwAhmafl/Xr5emKw+K/g7e/bVZuvVTUoCZqhU436cjC769Z+8lldcbz2AxVsOpK
RkkDHPeCm5R4Imnlwzzpe20zmcKpriSrBrcjdiBfW7Z3gDC8mGg/6Y4FafZkIJ5q
AL/R59GVbQVQ0pcuYnOZX0m4PPrM+f16gPWezJbIJzOkDzlQrWS4p8n0hsjdZHTZ
75c07I8tIAT36TXsZNP5syDUqW8/V4WSe/p9ItAIYmVvyIdDe+whZ1mjbYrcsIvf
Kcauf8k2GuGg2+XDxskuBdv334a23G0GzNNBNRzwV2cUGLVNVrBDnVK3Ze1ACg7M
faspVVhfu1lQ6LeZg7NTQJzDxiV2xTYlNnOBsUPluXukq4HGwK1sQ6YMBjQ/uM37
4eyThmyCd6hP4nHqMUrUL6gKhAe9G7qAhQezJwwcdGq24JCYmdkPSgTMgpjdUO9k
klG6fR2O+7Tio8vJCeO5s25RRqHIT6loKat1YEeE868j75qugC4ESUpusEBK7ZzV
TS0eTd+dQa5eTSxZy+gEWVQlBHg5cuJwDc1EdYu5/CssFXVxgxKtVBaxt59A4OrB
RLSjdX5xFrcTyg+JFOAUn4NCRbn+rM8E5Tw/AayW77tLx9Pro6rvYqfN88lWeVJ6
qv6a85QVWoUaxHAjF0X6LnDJcoeYhZLhQiFSlp9SPOVsInaOV6DclsExmYCX90CD
iAqL68YdhGBFvCMsoyhjt90uONlvnvPu+HNXA37fphBgwE2zs51Ct7zCJSW8ii08
e5AaBbKbNKntxgX6Oh2fnDoaBE6l6QCeqA8t9Acer4mbYrERT6FD50H5ryyyPyJl
cm0wnt6bPLecKB0L/OEyt8oJeKtkFQ0uDV5xYMDaq8v5wv41cibcBPtymcNYv8ke
MF4S1jfZHQjweozUc/ETQVsKgCDIhqIoEk+7hF8hwEZt3wYNAsVbLVE1/tM+LHR+
NHMAVSMsjBBX8fgNx42uhWD6NPw0A8nsJNesgiCuuKwXtihNUpv08GPjR0GYNGYl
VsFvyLqfzEvd33BXtc73oVFNXd0GfPqrVx7h4NFUap0TKC+3mQHbiz/IcCVh5+IZ
xGSWV806VZJLzr25xCxKYgAUd/whlDY6zXYgUtJ62/X6YJDGWS5n9qF9ZP2P559g
rI5Dlc+kdhooTq0okpzVUrTxoS2gIPpFov1wVa48VJ0QSINChd55lzxcyltRrYUs
P+ovLRRobPc19+j1wCZMhmU046aXjoPu72GJ/KUSiCC0+qR8aPjTJPbqTXuvlRxp
Dtz9tOoEhhcsJC/OOB0auzs1Oc22HNzwnChB/eiVeQNa7bKV/3nkP6A3EHGWWiSP
wbHj8piFLUFLxeC0wbVnqEGQHFIyPaW9P+klWKRIZ39Eaqo5D2TzCGA4aku3dYK3
ArOus7vo/B9rRpuWuysaN8s501qBsuWtaAvpXQVX5LGXhuzmBaj87c9ksAZ4P/ep
r4yX25macnPESY/BEQQIfcfy4jAKwQsfOq4Bo0dKZZApig6/QDe6XQmEZKnhpev9
GovLyDnOWtPOQSOrahmAnNUw0joLD/trYeZLq7jM8v9vG05KOsM5xuOjR95Lnf0G
xb9a9Z67vkC6CibP9VaOTRdPbxXN98lbuhTI7cVuYK1qhEJAp1XM8OltVkEjvF3Z
aN5KVSZUCvyv0RSD55BvpPnrOHhRKR7GcLjErWAHEIqeXzEq2WRLS3EiRe0oOQ1h
q8WJNUGpOgOZV2Svvyz9RTTSOmX5hYOwHhha5sB/bekGBdqW/H7rmS5qUFm+/CNs
tqWuY75WZXgBNbB2VzjKLztVpCSDRqbDts/ftarzlkcolhcHsLpdvmCdFmzANN0b
pbc9y5pZGTUopHD4zT9A7BrSKbcz52OS06ryghjDCNB3IlkgH6kwkuMyQn6TMt5V
U6vAx2I3g9Jru6HZa0mX2S74Ne49e065C7Vc9cGOMAwEcpQT9/ZUvZBrMVIl9vh3
mhpV7DoZK11b3XrS4TTJIUCSxqOgivLMzf131wwhB49CGXTHMyGAF+ieeGxFMsj6
Kjx/MJAHHnPak3oSqmLWNOmDcwhkDD2+Hb4fQgoh4VOIXSWTMKPp4L/Cvrx8+bID
8gOgFeKoQsYv5+o/o6rVC8BOH9vseU+d9Bs4W8msRUwRWztWqKaiujAMQDTpVKNq
a8HRFS8BTI/wS2r57ynjMARJDgnQ9Q0sgQR06Ptrh1nzBYBl7jIsufO3keDLVBIT
3ZR3K6ztzny9IeUujRBZ2c29hLuzTAAhCwy3T1UN9e1kwcNBiRYFYshG2wY+AqK4
4FdQnsFWXT+Djo7FKeLlHdtG7Nnaj+9eLZgugqprQmv+wgYTcOWHotGsRZf3YPUu
9sMpbrSnHxEQo7AT49AZ9yfsRTLD+rgIbX/KWELFpknZ6bNLd0uOy2EJWrnZO1ca
OtJTqh34WUP48cr+8rc7wvUZ7mdkm/V8vzRogpQzIE3Lml+rUtf5K8bknicgy6rK
v6NIZeIkfj3gyJVAM9x/OHa2CK8o/zijcVidoDmrWvUJ6pwJT+HhPcl2cgKQl8v2
MG2nBWdp7vjXLRW6vTrZFcQFuNWSgxDUhf0WKqjxyfI+g9g2QBXU/h3KhtTgCfjk
FLVfPMgT9L4pgeIzepHKi8FyfXxo+jaG3bx3NtK77eGfA8GD5+zuVNeIEp59QRPH
cDGsMh6Ykac56dNOYnBoJXtp7zSJ/DmwTtelmckPbZ+FadkK/T+Fv/Sx8Jjk0wRP
mTxuJJ3eNYYlduRFx/jGr9BwimOAsVZyCiVcS47b6L/hQjiO/kd0aQdo5O6wNS7o
GjVyTqKO4WqdjnxW0lwhb5QdBHoPwjz9uB9712HcK3yR6sQpURoe2k60aFNiMLnP
5nHmfLuOyifCQco1YU9bNv4SOUJZQ9ILbE+jj4l0GdUuhJfrR+HR2WKSAWQWRE7X
OGO3uY83mhR5sF5iX1Mcm2P+2QG48B4Hi8M2AqhbA6YFPL4x4C5Rm792MTFPh0vi
CDq5OyO4wm1tWL9vQyYnPYJfcFZ54vSri0zdPIuCv+njWe/R9DbdwMc0YVmiSVTA
OdJTQRd7gGNeb6kP4bW2DZp8+m9rpOyVfZn82GDqyfsJrA+ahH4KAGwA3uspSeMq
N5dmzR40FVUTscgYQ5y4/yj4U+bSioFRk0JPWH+OA0QmWhgn+p39QKDA/i0rZlTl
fhiNgDzFxg7gWCa2NYHHGwReeQaXEkOrrvg3fKv33ldbygHr0Jc23JsBDaJmvRr+
Nplfl5FvE4Zy/aBlhsSo0lvsRehSRQXmP2x76tMwfm+Ro/uCBfGr8uNkeMM1jyIT
u6LRnhs/GntsTOVeH5F8/8Qi9v/anNTDeGwCQlWpBVJ5Acx89MERj772YxNUH3aU
ZIsdAkGf8evBR6LhhlzQmpEWMGphHCsR/HMXp/qXiW2GyliiD1ibJaZGKqdBPlMh
rQvHO7qzHUSdFzVF9B+V8ykokLlGY22JnncOHYrCxGjp7K2tcyHcL8+DQzPrsCvW
ce/dRwTvEz8zF9A82bLTyuHtWSsFkt2rgymzHjt7xUE81KmbIT0CeQOXMZROzvUZ
8aOBngx9ZvL34vtVH2B6zLwraXDkTvk1TCaprcgl0ChE0iDtSYbTdQ8/KVOgUxv3
VNonoKfTd1h/oHyM8mJoq9LuW+tbuG2W4S4niVYFVxyKVBmhuJeVmKJzIpEDxw7U
RMamBT9rYgFZ4RHmfPBRyd4oKSng/DuEQFg7NPIibDyI5AsfJmLWXvYNteZpe+Eg
73m5fWEg9ea82Ivpzbt6KeEsWgJtlV12w0ueg7t6TW2fnZo7nh9+fA0ADsXvjgDJ
ANajOBpbx5df4c7eTP/ldXA3cEgRCy2a+uB7BN5JnN+rH6TAgmJJplxNhRyjWtMh
WQddt88xmAk52ArAyvQc6SNDJR985V79TJDsYw8YL3XNZS1R7Vfh5z+mnoIVhugF
3ikzXH7G0ul0yDPWuipsRHlqeKtzh38zNE0oh3arhJCxIo55b7AOMyB+mpEhaL9i
XSZReldluE9OsyGdv5l5IIEJbQRQKd+Ei5QAIAXby/gQ3JMR/5Mcpe3Ve4VSP1BH
yPzKu/dc0KCz6iUn2KjbaGBqEucgkBIa3JK0cpUYESBG8iB+p+1cTj3NgHE55x7n
2AhIv5c65fTiZkJEvKLP82/k7C4XulxV4EsYEK+KP10tHmWxpp4UuU2FKUb2E1+c
+U9dduvhembu/9NCDE7fFxb028PNsGwcID3Ka64L+zujVZ12VVLqca/uZ1zM+Wyt
O8d2LaRyKLKNNrx1x2ZZJ3AjCrfd3sCj+u1I6BKOHoDhNmtlXsKCSP44C6sI68Rc
/AI0N1WSgcWyXxL63vH/UslR7DttKHsFCS4MNx+aCK5aiGOEI8XwG5LC1SNpfTzz
/6XU6amZ9cAx4X++N2Xn454d7Cy/+9xgZL8CI0i5pN2gks6PQil/W+dyNV0cIxAr
1DlugrLnq4quF1zMDySH7hAm54IlySQrSdqtVRAr2qZVCvGCg+v27efB5me3f80W
2OGLlN5qtB3WDg5KgNy/CSs67YHd8cBHCaKAPr3KKVBGRHpyL58JPx1GdJtqzd1r
EQgfXv2SWJvYBbdDLcwL+/Pf5ZAYVfy3guqiO6srcQiBa8bOF1N62WTzFKEOlJ+s
/xAXsI1tXcucHsADJBPfKJow+nt5KnhLBoDQlzDyHRMzmoJkBGIA6pcpte1o1+Hj
irHKzf/uLjuCrYtOp0iCpF6lsdh3O6gP+OJcvxTI09RDWx1RuFZdm2X/9BWJxS6B
YHtOWv9fqCRDt7a2jRL51o5+ucy4rvCX/9Xf0kSrov9DrD6Lu/oVmIsoboY79B/y
UFeV5aBS39SwfP6FazqSjr2wOAfNbw2ZTVHuZt3ZkDSLoNo2ofFxShhlOha6aYlP
8v9G8aw17ySEfA+r5peKEDZ2w5jmwuupznasM0M7L80G8ALDxQpLO2EeizVSR9XH
1MadNL4j5NgXQTxdjYU2ohAb5AyPLg4JEwLwx0852DKUW+bVL06jkpWtgZYskCgV
mDVC7IFugYb/hg1/SN+/hWtmNvL02dh1uA7D8QeUjScBytkDmb34sNHywRRmlc1O
Sv9xz0LJ0WqTCQRiKkCrgwluVHj6d66zv+0T5R1Vsta6lHfUSHsZgixpdOUuSElS
S3eT0qXrKwWB3n89GKa6K3OGPSEkzycwZxgmVprtOCLlMqMXrKteuY6bzIruHZur
427fGZ6gqhEpSWfhPb9jgNAa6wWru9G1eg4q4kFory7Nm82/cKW4bEOAIq5ZXar6
5LaebZfQjI98Lv7k6pAsBPCbHKkban+87uLWjIUatPzfBDAJAMpC6CtkgJ8B7RxZ
Y+B5GmPtoLkRq0ObnVlzurfhJ7v92ZUJjkMECcVGeU1GCX14Ey0Oik2XSwYDZkeF
EWt9B/dhN+Aul38vczuSyu8aIkqw02kKjiumOKdvfkJNaQF/g5ZF6ax6sEpE29DX
jjJv7CmURUORL7MmHV0AeVun3u0fksMnmfBCy9p5wepZjVQ4+hT0mpEaRo3R45rn
EWQK6EKXnpJLIFm9zD2OIH0UIVwfIcyKovgdfqDFzWvyu/FRTSsdUkUbK3qBkIzq
MXGA6aXiCp8qGKLRFgUQKRCE/nMk2HQhJH7pLFUKnjYVrP4wZzTO+vQa55YO70Sx
XbnC94PzYUjJ+H6vzU0uBLdw3rvBdCcHM8MBlqhgTddy6KDdcL1Bxn0loI7eKbnq
1606NEXWMfPz0Q6XwL5DpiYVHkih6E+IHhuHOOW/j5rOEuVj9PowsViIwPus2FsH
VDlOS2MdhHsogXltpDLQ7nHAWlR9GQAp03/+0kVfSMFEPH1iq4KLeht9DrtfjWtA
aQBKjIsskSH2XDkhww9dI9XXn8aoAn3nKsqjPzMdeS6C5z031t8NbZcpvthylGVo
JtDeSev52PQHuEq7m0xwkr+ztZ+1fsWvFRuo9ExLFai7sLU8tum7bE50bHBrFbuA
5fTJHEzFvllCRcNSDu1v732gcDEsf/RJYgWm4+ByYejD9+Irc1aI6Lt8nVQPNh/i
eOknuC/nNf0Bu4hUzVE74J+zDvwGWf0mASx+6JlOaQzEbw2sBXnxG58D/tVp59DV
MiohMLb4b32M/x9XPD/MFxu1+AAWtdIzF9RKM/wIK2oXl1+X+EKrC20MKGZvgAZm
4zrF5NPK03uh/FWEXVwKr+/Ir2P5KpE8A5XRGzA2Ub58sgSNiNZYfH5MZHECXux1
VJ3YH7AO/rmZnJRMpNrDMF5ESNnG1FOsJH2Ffd9DkNKuDHQr5F2J8LufzwYkeRCS
grS7YWHNWhtYAix1H4VzwINMLqipT9YGDTKE3HNuirAHAcA3p7eab+rI88hnry24
DdKJjXELnzgEMa1MiCFOsuFS3Ck2+VJcetFlIJzl2OVfSl0qsRkl19LuP9X1VKFE
1p6ORWJf5GgG++li2waPzsWqoHBC7wEdSpZThVJPI7gXoHdrBtO246GvcnAHOoUa
tHTL5a4mroPwxNAg2C4UBniENZyan7+cHYJcaGhsoY9DSKYk5yjD+ASpnPzNRpN4
UzHBQb/Ypeu6EF0euuPJNmGFzKBwT8rleqb50K+4JYgUgzGNkGgRSDp0vIBSsi9V
WlwkId+Y4nsAiyMOQEJmkZIDDoQ66O6uAYwsKuSevc0Y43oopE1FjxjO0JU5phXG
SPJtFORWRhM++1mPRS4hntlxvuR6/+dmaXKeJoNmjRHgjoGu6FFbIFYxPIF/faZp
ikf9bnN5TvGF8VfM/+MnlVWMQNl9OgSRcoKDMI/gzJf73OJ4y9aJhRt0lJt8VX+l
qRXJnTTmOycXHlcJXh/Hwajvz/ofXjHE1sxu6MZ0A9TlhruXfcqsjlx+waiMuA85
6wEruJcMP/nEeMyG7hLE3gbwHWKAx/gsaNpzSsRcghI5udw1bKWKv2fCeSdbdQo9
IVGq/iBr06zza0J8Feu0lXcewqbhlZir8J0+pOnvaJhCSNzma3uCsD0YVmH57MQs
jo5h3aB0dnOJlsWimJhjOuXsLMQ7dvFAerRBqyQ0r3CyKsYcN3mRQoEKy3BEEMbH
xoOZS0uhZYaLsccEYEbtLxY1Dh6XNVhNvQMdU6qC4sDFIvLOXjTyCqmHViiKy/wa
z9Y4jWDkq3VKQpWzigy8b9fL+ueoAgaURC48oqBtjxxKquZXAuirdQMe9HjgJcBk
gbPmOdqfH4io5p3m3qIgl721k3msiGQM7Hscg2KbKXCYGM4+8Yjvkaeu/EntpPPi
9nLppgzpAMfVmPFVcZYzzxa4dU8ymTTmCpA7hMX+XBdnZQMRVeD23QJWl5RzOhlU
uGOyMNQATxdDQ2Szh6y9DVd+GRzBaADE9+iX3pBuK4+e6qnl1UhPvZ71mk2aVoLu
4EJl5LeNG/F59sxTxiUE/UbgmA+lzYh5mdItY1uBbpwg8LsMWONyPmHiyGgPVOPK
wz0IkCSpfzp1YYFeh2crf5pJ4HrwggX00mPYZ+oXunnjWihfQhMMmgTNTgCotnMV
d86RQ8I3jta6Y+OuqKFbpJn/W/WoL7iN3o7MudiGufWeMp7Id/8oQTUa1dkHW9N+
rMl6iAJ88xiERJVlsmw8y2YNiiEnQGdsEfRzk50GaZF2MByKVlPPib6kdWpEtuuc
lOQsW6GqsWudpB2cHKTtqMid1EzfiR6IJj+j36/V0vhGNpUkve2Gr/tOV0IJ18Hg
/ay8S9ob2nma6ftiRbJ0E4uiVStIey7D3yNPDkPwaraOrwJaDXQbtu9fVUMxrdl0
Fa1Gx0E1KM7DW0NB+f4Wf7QQ1qckz0f7+Jo2QfOFPGDETJFuEXChGe1Y4Ok/DQH4
KCNRZz2jgX05KegevgO4V7MNevwUeiWcECnmPgAdeBsNMbu7DhM1EegRKz8hyncz
5Ms6lnm/9ELFaXBZnE7jCPzB/sZUXDbo7ma8vhMKNK/5Pq32iQN9R4RcYZIxGgeI
8ckBJorQPk2Gg4lNrpIH9HxdZ/31tZ27PV8KcnRYDpppT8Ltph8TUBxuXRra8HAG
efLDZVONd7TDqB470lCEEZS0zZqLCiqj1tMGvg2g3iXCMpsHbDeOHoq38Rvg71xD
Dv/jE1cbN6A6Cuo6IaZSB5kwx593G+knZY0viwkOfC1DeUXobMQ2G3toUWFzn0Oe
KGmyBOGVcfsg8ylY3YsbQo2r2xCpzWVj9LoN8UlXgtegtHnqdQwwgsTCNtCqviFt
0zT7rs1Ad2CrdWbIO7jKRlC17TCbJJIHwcsGRvLDGG7fU6Kcb+iPx47/kc0/r7gF
pbYVq+/v+liE6nQ46TcyC6IgiOUAKWLAx+wa9IiaAV8i+Mr/1whHRk7JwtLkoWsR
8FWyWJ1BKREN1OEKcX5y+gxLA/wtHS2PpJs0+OGxtErF+UBgJJ9IjNRoHFw2dTf/
t75pVptL1Rolsz7cRfREPIiTU22sy0fz+az2RD5QQ5HVdwS0nlmsasl43ZqWAyJc
pVQTt4uevuoEiNP1DnIy1g/TiiRTFWhfMPyjZGrdXbierf8GPA3Yo5MsPHeD0Q9O
FFMDzBWrMxTx2WHJCEfU9y9f+be7v2rstir5Fg2YnGgY4xaIt61vUZstqYiQGkdp
yTcwvZ0wKmvBQzKPZLtVNfko0QOf5UnkwCG0ax3lcPg0yn5j6mCVM6xM7sSGJVst
vuTnJCFjlwt1WRcAjOnL/DjNblBLkwF3MXVUbDeQjHXRLGC8ZJriH8ZWr6RFqHWJ
9N01cUfmgVo4Q6JG9p2mrD8m2d7IPdmE/pwU1mWX/sOhW5ZiVyS36/P4oB6NRA/P
N9irngXDXucUYwJXAh4boo+ha40FhowgwBwVMatLSwnK6ATdCaLg+PTyXoip4Edx
gUlSCqYM/YCe+cVDm1fgqRA8GTjg0dC+Oz1ecOJE8wDtzRe9iqpyhIdSfRXChIaI
SjRdCV+WEyxWX/PVvegPDb4YaRgnXuKDI8wGjQ7O1EJ9yQql3TvyLc6bZ6T/0z9m
cAUNg0DehCiX2vy3ujk8tfVfEP7CJFO2UKqfYooGz9mntO0RwQ8SKRn4SIB2W7hO
SH9qCCab84L/uZ1sxE4h+lZ+ylcFRONXR0cYXkQy89pxhX0MuL8FRiePH/ZS6wk+
8aWX90gQ7t3MLZgHG2DpSCPGDfWGF40eUsKs/ktJLZL6w6cyc8bOFzpEO+ydsnvc
C+/HKTuTk8FrM+NR8M7klWoZKeW/2J9MW7490/h/DENNSfTLwOndsRWivdexQ4Ca
Ts96u25sXf1tkV5nnjGnXzNdJwSdANoFPgivuQx/3oEUDHzBnRqc+mNTIsDRD1L2
v3xTOp6EkRuIIIcRI0F8ejZCv2JnQhsHA7c6f+y3tVZT/6m7l284ywzgEJqVHiDd
ZGvHgO4CHFurM9gMfEvhnbdiU6/Tz/WzGAGBcU4JwztuAZ52ez/cBaS9iSMnrQaJ
WMuQefg2dDZNVA8U0fEF+60DDT7xdTMCGy9lFg9VxNutS6O+Bpk3oEPdmmK6UnTb
/XO28bGI7MZGBxE+YiD9RvgWYit7XTXMCd0pM74WvuqHh5tUZ9HbvAVMw4c8BZPX
3qjn8PGw/0c9zd4ztMkhKYD5Ykks/TFLcHsj+z1CX0idoDrOrXNO5uQ2G8VdU1Sj
2oRzqP7yXt1VcMHsaM2x8aAldqtB0mHBQxI8MMAyxnHSwktj2GF+vrshw+uMhhdA
qrqfKtmLeAmebsewrV1FZFYMtDXmrMDEedzezWXCYZtIt2jdBR7Wrj9mT2mBBWPc
P8GU4sa0QaoiR0BDlkuonITG3vfV5ItEOYkl+qMG0mLpVNMZqn03nwjExzdtykQE
GxWVnXL3YXhYvOVqQrtK/kKGk0uMEECw2gVtv8b6hdscYP1KEAFv7p9cbdoY2U2P
I3GHfuzOour8vjlnkfmY9t/rX/mk7qp2ZjHLjdYodzYfwoPhxxUndKmdMlBPu3h3
0xhcYtaW4pMI6cDlhDXGyrO/g3aOTF3aPQ+omUCssPpO0UdQObc7Gd/+WLxg6ZqF
ElKujfNiDmHsEYL5xAqj3bZbfDBtVE9yJpDH1jrbXetIRmsQgX/pz4CdGjPW7SZP
hTepxy1PSt6AtjOVWiDQJVq1p5L0fxDBqtVQPop2lyAAqqqxOAkssA1YUQMT9Ia/
FZiuRWf1QDs4s4XPC8nUjf2VtrSyZ9btlly83WME5V0A9i3TDrHSw+CE1JUS23AX
18vBxDwH0XJg183FTOSGMpN13TQhNyNAqpRu233AZblBuc6DhSx/hog9hHj0ycQb
FcRsX7v/8gBzQspha27AS3yNKuab6kLzv796UnOhUXicc/NiY1IJKa74Dif8gIps
e9tI9RXXcWVSdPqAJ38SAe4c41qGJ6goyRRi5gLMmoXxsMT3zNPAjYXg9BsxB9GT
mtnwwEUWO+1Ze2egGy1x7p2Nb5OGxACM8cCU7G2RxlcKSRPPvZgMHjcJW51Y/k22
kvnL0XpxUhHy6DS6qgy2v7NhYCIX+z46rNf6mikC6k5hDbPMG7DhEoaa2YNdXTaO
JZFxrWPvh9KsW6L3t2EFpOBTx56gFNb9V1DCkyG71X41QMXOpbGUfWQuyYT23wEA
Fl9wpG2vKASPn6XLzFA5frSSe8RLfQkLpEIn0SUogvtPXCPp9atieRSZAG4gy9v2
kFWOjS5J2B3rZBom3ntsoiDF+En5OyvIRU2/NAdCrsEkEo2+o4GRCKzdMFW/vUmd
Drr5ogGESGhpykfliwxbPstuJOxBw3phTl/fRtWNqURAsiWhrAUmxHkyAPZKWlWW
7YFBDDz1FidLZ+KlMM1heSMT3cAogpbdGui+vu4wX9XEWKjUefOvJ6GJfRoaPy8A
t4CSTBRzMOpZWPmtjClqInAg+51hCstz7qrV6UDVZzIZhnSyJflX1Wn6GBXPOYKF
X2sp7aC6TJId6e0F79KIqnP/C566sHN7WRK4WqeCaSgo/gF45+/QLcTKhDEgGuW6
I3IMuoGBQ4mfS7TcmqmTanQmYvQ8BjsjT/675N+lBaXn5mpnT4cdW4UhGlzKN888
jWY5pCI7BjLfwRlEKRd0u49ymCRptrh+Fi+950n8pHLr+TOajeQjv/YhtLoaNgXK
sJboDokRsdue1MA4Kfgm+ECaUpfgLQNuAZhvQfD8wzG5hUIZ/yfV7lT7ikyU835S
kK+QEDJ4dabNplnz/0K3F02JDHNMy7vFiWVvwnnRAtRF6aY7Dn18dV+Rd3kDF2Z7
lcMVek3VpVy1GJwoiHaRTQKAKilZm83VJfsAHbl3PN/MzLLE2azxnyUdH6lkdLb4
wurh443TtyrsT/Ayx5cTVSay8AAP0q1DmCusD4C5BgUffRFE+ywwt+/4gV8lcgpy
xbgH11lii/6c04EgISNuCNtuA67PFdX8133ByoZ+XsvLTLeoQfBAIs9KZymrhdW1
MDp611P1d5LYs16bVYTyvymiTKHKQBO5gZRLBeuBOR7qEkf4caEhg4v5WLVu3EWn
Any3J7UjkoLpaOphSuGzw4tdbT/8HM/EBYoNwRn4X87oa1SDfZ/OQFemCZdrhNXV
nCg5VGFX6spGO7UwOdKiFw5o/Ks3GIUQKMgTdYOWzhgM6nIuY+RPIbwNdx/lrbLV
mqJqNPfucYMY+voc/ZvHi5SqqIFDLEEyfu1hI0qT1M45Vtf54SxcBqsSxx1BrLZS
OVS0+YqXgS4Enfwny+bHFV+yMWNcjpyOz6y1YfvrfYsmzjltdirFS7D/spCsmcQC
0x/9jjqBpGFebpU2Ns12O5JY1OO1dAPdyKU3ojG/ERuxCVB//3PGH23VmMoY4t+e
lDV3C7XLeVTbgAiN4xAF7Z2XyYnAiTD6uYtKeuiOjGTm5r9hc6OETvVt2vSN6W3h
A5iKi4D6zhVqMGuECABf9lt78PaLU6hxpJFxVEcpLHeYLWBvviNsAGxiikNKjhx1
oFIJumdxbk/ggT75aaLxpyHqTDS7hNvOJpiAdEFfwNOTJh/zToWvHQG7vIGS9K35
kV2ZQnbB6gpk6kDtmZqVa1MUbaY0vmhc8F0vlRqJT1TAlo8KCBnfQxF5Uc8DJt2s
YKd1ZT11NR0ea5shR0n/sFwea/npGKKjG4m0KFhjcFpBp0HYs5fTlqRUQQsBmRb8
HB7dKWdVwLiIPZzVOpoKtLXKHKohkUNRVa3/5myOpmtnGVgkuqp4sqq861xmt3Oc
7KKiIj/OG8nwBZ/qzuV4+RhLhcWILEA2wbDyfQyzn1bvgt3+RnPxv5Ggn8jglzdk
4W9GEL4GfmAZO3Tx8u9aYnmzcCR9H31w0N2AMRVeWmoc1p8/h3DDO0l8WHMbAGwg
piFGsUbZn43JKDBnP57z2ipwu6AuwCRqSE/pC2g/qoMiGit2zuq204pUaz6xhKho
amMR/VrvgDoonwZNGLu1fJDpeQ2H8ooe/isJWVBEy/IbpP+Ga/TO4Lqy8wtmBitA
Wc2MVYjYmuPHiLbjK30QxHHdeuY4+8MdhvOoRiHv0iNJSHIsh+24kzuf2SbSf6r6
hOaBeKM1SFkJF3z90LTdZ+J7IXjzNoQ5G131QI6lmYMcUKa5tg869tZfsOGY1GZV
NXksnQBE53HE6lrsyw62auKDqSjaBUd7QV1PvciHbK/ETWR+q0YkbbHzdJK81tsY
ppVxYiEB6Toy0TrJpK9DYuA3R9z3cXuXKHwTr9GCimWuDdnfPry2iDue6iaonHJg
ND4WQIEhhYVq4rAXyRS/pDUp27AWFvxFj02DUaqqN5Dfppa9q+Zh4nEs6YllETQ/
T1myq4kdwu4MAL3bMkCBHeqdttpfXuIhuSJaiAg7BLidfm/c/PBhgmKXSpWhR2tl
+cyvx4uovFyU2gQlO+yErXz1SDcu7IjOItfwczjp9XzNTyYbrKbtu+BqOKeLCGe6
aibLZYgnDjmV3yFIlwLF6OvXxIDrc74MRAhTldgZ+wQFgfNvOYXX3INHA0xrmnlW
wOWPXhyPZ7wKPBrjknwncKPGg5kYg83ZoSM9zKOZcd56rPHItkn856lwAuZhe+JT
u2RKsA1ZQ5lUrgOBut0V5oSpMW+KSiY3i8eBr0BMvE8aHiC6VtDv/jnw0B67KSOB
5VSfJphcRkQGu7Lid4YbgUgo055v5wA86zQp/mwuKMVKgDZuMv6yOjzmFamf7iuM
lZboMadELM8b0D2233yVrVvMHmdj+zOaMlNqLJyDj6uevX0mhUIdftCyCUPb5Kn+
gBLIms9ZQ6eCyiIxpwNQZs0NPiFivrDBwI+78fPo+h/aZO3p7rb5RYVZT/ja/21G
FFePW7U97MKkMZ6PZQ0lGT6EF/JWAEV2OgqtkWGpSr+iPEcQJdnFvEvu2qHEzCgr
Z9r+jNx2CPYpNkY2bOyLMO3nHgdv9kXnuqkXWbwx0IOkLaWTVHlhiInqRevvpcRP
yEizGg/9Bzck5UyWm83wjdkjetBPHdywJaMul3MovrU1jaavb4vcw2+Jpz7ObSyA
T2H6rOOgbwQ7bACtbYBVwTnqTiMLn4r3DMBQFhjhQIZ+yJCYA2yQ6jYkMv75z4BX
Bv3/5jpfHMNJIGxOJOBwdJevmrA4N3XkuTY32WE03VRFlMF5uhoKjxAupmzXOF3f
+pe1IyM2N6tPyAvzzR5LFXl4cD6fl4W/dnQlo7tFKMnF08ssl/x0yr0mOV44suwL
hQE3KqeqZXydQjQax8a/O6DWy75lJv+6dioRCByw6mOGrjuaxkl5Tfwv9bn6/HVZ
1MJLZyBdUjc412dv5Cqm9leE6qt2/58WJa7pTdgUp+qIEq8jK9z9b1h7/+syw5eo
pdt5vGl6DZT73zxAsswqFAs9GM74mEfPSLAPAvCHegYAt7QP5UIsIkMt/1EpwKUH
vv53MhK0XG+xeix1Hu8NvdupqOQAng/XInOOCbwj8sHPGBkko2EREjmX0RAhASXW
fYJpDOTitVs35cSMvNjNl2MKNJsJx3KwGjq9mLi9IlzeL4GH6FKqjEpG6oCCrRpu
LBRnARaqfR3lnstCNqH9dmsXwrPTeAjuO67bvZnP+/zPtCQOPTXiXXOjlS3s8rUh
kP5bjbt+e0nbD8xhxVQxEi2VDlfMKCxft75ML2XKpDNHLulO3SlRRdy7LHsoU03a
xzYWoPPFv+A8BNZOfYYWztZcCbi5StMKW/8AnCbB05t8sN+0PJOnYDnvnXnmuj18
mbN20QZpTEUy2MS0VUjSLrBV3xZO12TtqL4g0C38KFp1aZUwaeuY1aahek9SUM8w
aKYfLULGwCM8i0c97yW+3USQpUQ8uMoKDLg2pTyLgAJxvoCa7yyH63MKgP+LAR1Y
rryNVYkUstZapqNcTruqXB5bFziWjB+A1QbMqdGLKM8T3HW8EIypFmzNPsolSW+1
jRJToaGlj3m1lnTvGgH19l70hx6NyWOumIwSjSMO4629E39k5IM2SO3weI97HZs2
ukMx7B39OXwgPhA6JSERUZYlsCb4/d/lZWom7sFiBBJUoPQLcJejwhMNETjhRHTk
/x3EuAwgmus3XtEGBXv4sKDTnje0aHfCuLquWcOOvsKcaV9f+hiyMM05+BFGaGa6
2QNqvqKQqHtJAFAZOHD7niTARSdNfAhI6EygmdSJ1YwLawEYZ9rqwzcHlw/UpWcg
WVQdEciibcMvCFG/mAgz63npzGKVTOgDNbuvn70PCAInzEUHXFBxnwVleoy28LDM
WBhRSRVhgASVHsHKFPi/HS3dRu61weHsL8nnmEbYmeNsRH25pGXpnv1JUqzPNf6u
AecC+oYmdfWXK7FBMMqnHA6pYK8jD2EvFyE8mO+e9QxinwCpOb+m+2gms+Ia2RGW
yo0DQYfDUx2gm6erbhfn+jXASIhi4YN5zQiL1iwMBVJkDrGUTLSygWLKZPoXa67k
7SNin2RQNsGusSoy9cuK+qCtthHvAn6WjwAMkPEmc/6RlxzFw4MpcsmHH/ZE37+F
6wqkw+iGGnUF78z7KX7cWD4qpA4Y8CoMyWqGCEK+jqmWgQiCBFg1mP2rlTTOqs7A
gvA+Zviqk+VSEe11IJ9FcizaakIVeU8i4oiaV8QrwBKdchvdc5v/MwiRARPLLmIP
kYW9BEJewuCA0QCPKYAYp43MZOfSIxbwk7NNvNHedkmYmhv8O4wQwroJ9NBKqKF4
GZbCrpTBIM/L6yhTBRso/tkHMKsEx60xfhZC4bqzSQUaMrQ29Ngyfw7yiAM4oHWJ
asLycdPAwK2rpDm+15046Pj3EhBmIntX9e5/AvkNdTAzofBBXbwPl8n9iePtSwUd
9LS1YvQXmWRy2f2HZSG2peORM0Tvh1AmffP5F1K2Db4IYHM8qecswEyirkzTCUBU
fhpb587MA+bdhzsgri7fqHuH5seGUt+BFKUNu80zgHl34gcxGmOfAXFtqZcr7sCR
ybxozaREGd4E/djv7/vXbXDL1h8bAB5HctnpxaxG0jJJ/+6kz4TkoFA9QS5gx3nZ
K9d0vpkr+4yr0waTj/M8AqZ7f4ymQixsDVI2ddG3arTfEyFEDLCfaKTUa+Zgxpg2
Z2AArl61R5sbef8AQYzQYQTw5+tQPmpuuVzmmCuYxj3cXqRTt8l6q8BCVZgynoZY
wNAvyIZrY3vR0MGLwVAz459rriVOtIFcpFxutbylWyAcvGeIHM8+mYZRaQD+Aw+1
ev+yfRJxZPVSw4ygR7g6TIa8wUMqj2lAMJ8RrMwicfLPIqrC1/zuqUFzYxJiIglI
y/e9TC/dYukxDPyDArsfF3hYeQY8vGIWrgvl0AA5M/EnwoZNl+S92SAYZ6Pkbw3v
eyY6cGJwTOekRJjP5OsMXLYHGdpy0BzFLio7d8BzSFVoDNWcjDaNxKxU4KLScvOF
Oy9sXg1U+G++3tHSdBnKSWgIlWLK9HosLV91QN44ypuO6yK8WHmOwN+puNKzIBPp
YMXCKjZ4gVnQlWkOO9pPJODYi5DGkPtagdJeQTlF7IGKK1bfcRgAD24lkhGxEDCB
yuRN8YEKLONhApRcUOSclDS69ks4/tjaE+ZzI1xer7oHYZtYQ2zOW0AU20BhLEXO
WppveGi+s9kVFGXURglRRVZNe3rSMur31fl9NnmJ7q4nhBJw62XL9bZMtMIqjbab
GN4oeSgoGTzBgMnFWbUJSK7jJ7+LQmbf4xmTOmoDc0yXjpDzc1yAQErT7P/jct0P
mkKFEsKiUuY810BV6xQwP0QZndujyoOzmnvavHk+GTIrmQb0teqS1c2HyShes5XR
CsrF2EwqyPwZHrw0SwIHlr6DUZlLGd46cc+ndZobokoUYdaTGXbq65+jm96UBYNJ
xB74IoJKfJe17IZ7Wmr+nzhOvyzCjXdJi9vUwzsNEZndorct5PTCBb/P8w3Snizj
15IqGDShZlogiAl+ZRWdqxus0NfdcVDcSLDkp1dAokzj2upplYCHBFBFzjn4RdFT
l3zpa/qM3U1pKIF/IpjDy7Ap4pjyviXngWkBjiJLPizuRCkooQNmwgq+weQf0XCg
AOy3SHjRbsuDedYdcn6KzODxcSuwdU6wGqlPt1zNs+Y0OpLV1lPAlOPVx/1pKqFl
tVNVE2p+letLx41hLSOU9ozDCLoHv3NjbzZU6kpZupBHKwHTXo2RT3pCjkJhFJSl
P7S3BQNLwZcURuXuv8Z9M/KUnMcPwF0n0LFyUWhMI3eF35SZaYegvwR7lGHGMfDK
Sh3ZgUOnVHNKjuDueI49dCFsX18qZOr7seUge1h+I9zhjTT/LAmgByeObA/Jdcan
U0EArz/9YTGoahptTMkZnYVoNCQKALDHXeyEfDE3sStbXwNU1A1Y33jkX2Mc+n1o
cvC4zuunxhcHXVJmrAfQywyY8KrDoEYxY79fV9chCxlK1y9aQbwGap6MHd+d3ajf
gBtie1xlPUyt+uh+3gUNc6leJ+1nbfjJdOpFdaBwCBSzvy8GaSv7RNCcw+IFFpAG
Ot/HwgwDlAy7Qz2pLh/co+fBmgJaaJke9U8uP7OCRJ0d+Ih75ktmkEbKtuAJyv4E
5Lbxc2Q2WccmM6uILc9YYkkQvp94TVVc5rx0aEAyYj98zkbi2yH/L2TalfGnD5ym
wjpLloTU3rbIpWEkCaRRHORXr09YR+DZlMpXFNsFM9wOBAilPtEaTxGzmsWR+jnL
HOWceNRXaZr51bL58khSCs1soX74q9xBsmmfQ+wjyv7OVYaLfV/Dvd1j2uYfE/aL
dJEC/QV8kJmSBcKPlhMHC8DTGcI5vZbj+dbyqN1nIEhG3MtjeXtfnirOga37ZBdC
Dl5s7mfGAwG9wEZanco44qoss2kVsjH5yK2ms0wq5d2puozB0RQY7NyBK0LzAJ1U
yKkjfSF+wkeAHQ7rWXzLfvQC9G0ik4t9JZ8cZ72KjCFTTkPJCz6gqGAh1ykbXTmK
cmsRsvUDKQKQU26fys3cYcF0TBOEstWwW1WBrJ8XtnKCxnp89mciLmZ3Zks04oUA
xbHbhjx9T0i8CbShGdz54ZMtaJQMpY4nciy5Q73boZ0fHODVXeeEuhcC4sB2PFUf
2okuv250j1EFGCt3AM6khhP9x0Jf78jHQGZFGFj4zS1YyJobYIqT/keCNIUkDZyx
W4odl7KrL9EXRsBM8ZQ/1KwzmA5F4u6347pY/HAsP6jCXK8VALLAsEp+PpPBkkwh
YacS3C7rFymJftcUqrGtsPFfU14otlqsGigC0L+ZskyCPNhdxGIGawNjIFtxu4JN
IBZq2HZ5h/qI6kVAS32X9Dt2Gf01Dit4wFYDgNmKDr1G+XwLr5nMP1ZjeNc8UQOV
ADuCFyQkz8oS1FTFgNwy/S3dfZfqA8nK/1MJ7hEhZJdgufrLU7HuNlSH++SdnKo+
R3krQhI18w+EqC25JKApBfZ1I03PBFwFF9M+ZXPeijuKBAE+m05kISZV4bFfLXy0
tuLOyGob+fsjpMdz6VZazjO4uO2OxG7BJe1+YDcyeSv8I4wyMeJz0AzX56KOdigN
2i5qldM3trHCGqU4X5eDOYM1oeMpND0S7S3fT8TZ1N+vhlbhAN8KZLzXXBGhaKmH
ltT4jkum8DfT+7zVuAyOermjbIYVIEXoxDPcONgMQMWv+v5z8X85/XPh9ChoVPBD
/UKu66lHpUYfwddN6CT/TCUwFDICaCkqMKI6XwAvxlapjgS8xpY1E/hEnbH8UOQD
cqzCYYkPn4tr9Ev57oThG4wpRSarXbbmvSxCA3tX/UcDwbc7gB+oB95Pm3mbbiRd
UVjpyNJClc+e7hOaj/7sqiqODHi0lpSsUuzDhUwrrv/zxw4XSRNwW0lshiRW9S+q
DOSsR/dK0ew49+vUxeatPa4IQkx5/3cHZiyLvJhHxIvDXG+45KkWVkRvFMvLKVND
7LXUKpfZdgyRjBx/qPRMdAn6Jydjd4W3+LK0pszesfv5io9DrJQVe2EB/AUX4BUb
r4oPzpSoB9dmU+VONVueaS0Lv/4k+/XrQsXBu2xF5O0sJJBc0LDjwZQ5v1riftYH
MJ6xjInq2o+mGFAC26FGY4oEFguJdn7i5zRTM4uDELOnrgyDhRLNrfYs9BAFLvwx
/2rZjH/V9CCQkvrUwE6heP9WDxJHtCN+lSr++j7PhecdHfdId2epGYNVdqOVqDrG
RMYY/lyRmii92boUWDNlCumoboOSs01r4F78cXl6zeXnsd1s2Eu1Jw9eW8oIoIGO
XQ9AKK4s7O04l4BfDHglZ0ybARm2wI/+BPA9E5NWX7IcfJHqMmbDwWt76eogff04
SMERA/3VPTYFvfFdk/23HzgHw6YqfNtH/HgED88c/9cIoOQuAJmu6kBZ8FRlB8vr
Xa4TuC/wLl7rDLSRP6EkNmQW+ASyLwHh7mqZLlIZh+7oA98dAN9gy+6Ckn4J6BUt
JyevsvrsmHgNzHsKMlSwTFyuGugPlm9ZQWLLeKdN54b75ZXjwSmCwlEI2CDBtSN8
qlwBVBLOguc7Hx8+krQIltGKuh7ZzY39eQ9VnogcVFx3VBjuRgWA/WcljTIVQB43
Rt4j35pMeDW6JZZsZElqc0X7G5lvtnVVjwvS99lCWMbpEm9fNQa4KAV4J33mQRDB
sLqJrbbpnBdjWUE515f1AZUj6UQJSHIqnPJYTUMlUjZHTNzFFcqG+ZGB8FAqJWtB
eRe9rSyj+F17JnxAiPKEX9vK3BG8qW3xgNL8mkMyuXOWwQE/wEH26mpO1JvQ0Ckz
3S21mfdaUjtg85fg3DG9RDOlumshsbCXsvYS4Gr7s2P2tj9O7WjwFIslSziv6ttq
vk0fTyoQ0ziGdO77dwOYskUtZtXUbVZmB6MbsrGv/5KWqUPZZIfHox1MtpEV8PWK
7nRqcJG+p7iY2X5eN5ZOCMQ4qbr2n3v/DoLlfFnEDHkuEXwNW7QKl6UFINYzXwAL
9lDlO+7De0/WN54VnU3JkMksxc4pvdNjH/HxEqp0Glm843Kh5qwP2aWJ6wKUGtXe
bYpnNXerZ5TYgILd1vGfkDbBVSKq5jd0I6GV51YFjAYcky/Tyh65F3ezGPIzyrf0
DIGoJ8/bFdRbbXru0rgjFegnBbKTcnOLK3b6XJiT2VSYE8vvJ56YWbT73R29WuAc
oMH9IkHXrOCpfOcE/xTaHBLA/8mqgV6nMA70vHdRwFAHj/dR2CkOMadNdSO1dcSz
E76XEROnBRYVEQgInCXhjLSlZkDtOg65ZTZnoghRJ7+sCSKTu7Wi0n6/BLpR78z8
31WpoUhK3NKDGxeIVwgefA7OGjxYnAIIcS8NE7qitVcXsx8Y4JFaKoZUrLhfZcpN
+rfFW2Je6qJeZlW9rzOpk915pc6W2FclqCNN5eTmevrcYA00AW0eC8ZjIHbP+FvK
mApDj6Va7v835LfwF87ykXyqp/fvjkZWRs7ntpaowOlnWwbbAplesxc/p4V4ixRQ
AChcCePYYUWFWptdJKXfCvJAD5yiFGLbuejoIN/+8HCS2tyUYzmJxgCSapvI882O
tf9WUMTRYk88I43ihOskcCMq6jVPkfqrKrlvAAarTUHjqFG8+QcIL4tdxJdCKpfl
zNYCRrRmbZkTHS8gna0LczF7M3bKkdYlz+Eaj3j0VCrVSfq2357nNzqCojvGhwZL
7TN3ZxKNqsgDiqQmA+2E9A1eoy6GKhBSZZvNBo/XOM2T/4OQau1M5AuwVSlgR95U
Z5wW1U+6Ru/7uNnqTNAqJUXL/2AhMCuwKD4/8ZD7Axa/v5mVpz6QU+3hjliwlzrL
e0cFTrjBSZ4KHSyxoY36ZPcbDG6CtMPMcXHvpOwZUCvQ6hW8GzeDHPcIb2LJha4y
hvvYgNi56miqK3i804r7QX/GVTdkxOUGbncpKb63yPgn30oC1gOZ3chaS+GAZWXk
tbvtlMYBVyIemWYbUhMi8leUbpaBns/FGJ8unA92WR7bnnuiYCiu983/T1DBJyLc
ABr+ZMrgq96w7en4xa1YvvDlVo/a41bRvgknbeQkx94doYOaYMbFUgtkITsfnenD
gmajHD+fhO90tRs0lvzvl8eJjArdw1RDOvescnXPHDdvIzDmAlTbexm4lOhAiFNT
pojwPnV1A8AN1fK1ZBgwom5ObxM6rfKTuqHgwjmeDYeAond7xSfGMnvC5RGjPO3g
OCv1YVndnJUWPsl2Op5KhguhH/eiCnJFja7+JmysiJjKEjUvNLJr4lzekpnzxRwB
+ru31pz9Y4PJSE7v54hmtSMbilAdDIPdqRIBxI9+B7bgWXEzs4f7Ev+bwwjB7qQr
bHJ+9Q10jZtrQWyjpKZ+DlWstu0pZtiNcAIfbBRFoBVFL+LEeZTndsTPNW9EJkeQ
zYTTDRUQLTDBmqlzgbK1SAyJWAPn8n7Vn+612zeEJPtAFRJdkKJOtduulR4j/P4N
5IDjsLDjvUZ3ia+77FZTK/RSshFK+SIXS+AXt4PiuA4uKLtZ8pBSDN2zc299dCGa
zjoOo51tR5QPAjqnBc+sH9E0iEz4e6DnNuUasUTRacpoyImYyb7n6UHieMOEaAcI
wlbbLwrDOCIxIxaaVwus+yicFOHpnoU0hx0cT/bWq/bd6WtUVNfF2QM81uvB+gnG
EXMkHl2ckJkeJFYtQUPSYUuxGuQiGzq8+rcQjaQf5uRCvbEYYVmokpz0X9aOwxcV
XJg7LFnafopA7rrR5uAwKZLV//JEKqQEWXj33FeucT4gXRvoh49SkD7sfkeOA49g
gBhtCnYRonMi4UshKSPmr0tPBFYXcIqSsvQV1vkz2jgOzy/sU+s6yzQ8LPzw9Mr0
KKz96XYCcHcH/hRysxplkG2jg3FBWCu3XeB/1ZyqcI/wdaenNCGVNv/ziTUJt+Tt
v3KWDkPEs2aajWeUhwC9/SwSO4EI8vVCq1JZlWFj6QOvquCZXcn/sUo0FpI2BFhs
Zcu6oH77zhGO9kR0CU8979akjwhFLarwCMS9yAWTOSQ2PqfHTsEdp4tKdnUACBVR
E9OLlGNFdTDOB0gV0C2bbj0q0uOxpvlC+ksjLgjmoPYT066q1Vl7t6lm2CzKvwKw
3NpKvmbNhuGt0UIePvxcysisFGjbs3gvLR8UirfMWQBKvctMXvhbLMjVjCdwiZf+
1EE4YEtt3ZNygPn4uX3LneFeoNkZwXX2PKGS4YePJsJE4P54sgQHdKzV3VCaLsuP
U2jzj/JghbDKfQuiKfvqacmK3ai2yKdRkPkHlxBQc/CH7btIQ8n1cbr/9uCxf14D
OxeQFcGZ+rEZIE2dMm0eEVKf2j8QlfJzA7N8sEierg9BUFKQh7cLf4f5UXbaXzfn
cCoM7OV40wrNO2Q6D0wNq8SBQjxZW3Fhx/I+pmq+PI0aHEYwZ43jFl+NsmATiYae
ruMjs1XTFabiW2Ay88GhPlIMFUgjzgQykeBF61D6mjFbpyuExDNm3+opGhlTco00
HsrKqDTAQJrLAOGQXrlcuWyfPgBFfS8lyR0oHelMg6DGpU6LhHMZwrfcMugmgQlN
Y6/Ffb1q1jM8wtUcfTEIQBt/CMtAMpVJZtggAo1UbAJ8YyMZ8W7fGlHaAsqgLHRk
EYSpJSIlpgskbQskans9dhbvOrYnrevA+G0/HxgiLx7oWDi6WHX1QlX6a5bHtUis
Xh+oo/680ITeJXt7U7a73VT8JiQS5A/94dcRiHERzHgtnVOYHnj1FzPrChCYU1MI
ztLrcO89mnxVjnVMpvAVzR/nyQhYN3MYu2kWeogq9MZhbqUf2e9A5dW7LlkeJTf/
CUcbBZ6FjL/xSG4hfF6Ul5+5oACHQlZAEdpSnzHxifkgnxsVQcfOWePc6GrgKF+I
mc+10Z9WDg0mHY2Fj9RgTJsO/X4Q1ogJlR/cQhOCBeC1vMGMhAIHs8Xo1He8DCvK
7e1v5Etlh+Mmxw6+5atrXFwooCleCeB2TnlLp3P977E4tUyAYhqM/3+1RpDcZdjH
2lOiSzdD4fupQIU2m/JuSVkra1HnXdvVjW70ZryIxUZMHUzXuvw36+zeg+Ve+HmC
/hEeWnkDLEGceFej7yhHpjj+VtrwcP4fZjZKcbfaRTUpJHfhZmFWBZjbNFO5lrvO
v3/sESRZmeGr+UfgffWzuxKhwmjH8+7LN7232jVv/pton2PZN1pcZasbP8V3VBsI
zQWME1NIOV/pQaAD4sdpXfrYi6MMItejQ3GHZBreTKUe061GTHEABlYSx34tP/Xq
YjLdUbZH1nZcHP+KAnMSwbk+RQa7rAqJeWW4IvKOZCSpjDGLh+4A4hwFlPp5lSOX
HOVpDeiNWyyZBR+EWimzo7fwSiW3sR9Inn6AW1kRbk0tpXa0terRYBAtQyqQ6R71
fYTmfMNi+steKiTdiTcTE3LMWnDTpvEZsmqP5T/RxO/T48Emlm0X1lH8LG4KAmCK
Nqwx8c1SNTZ5UyP0Q8n6/PpU+IVNRt/YRtKr887Ti2L8vAlwkc8wwEH7/8OHBSDT
1i5kDVqTPcwe0hxX6yZqwwvUmIHF/Fx4n0yscpFzGDrKzN6yVUn6s65FklqkOXwL
eO4NpoR7HdoXjGAygs4+qQUV0cg6e6HPtofyuBLVoG0HrG7P4o+lTj0xw3+jhuAa
lDc4bO/wQTZVdQ6w9tJPxluIybdNSWuSQLF6tDRrm9Te29o7NmeIRxF0OaNQfPqE
zUZY1qHehJDOaeDJBziR9YDP5vzA6Bb6VnjCZ5AEkXNOrGxiLoSVm8ViN3R2jOIo
HLNLLidx1d6md0LZ7oZoceteVVncjxBepwjMzwnz7bcNe+uOkPQfmRwK045/372P
LxlwiF1nO75GdJavKFBKKxLw5JiqsisBmquK+3vjRfgrZBrfkEDZs78env/Rdu6S
kv17ze18O+6GEoW+O65LTH+BI3yn3wu3Tvlo0RBu1PiLJAsLRioMFkS9Q5Fmp1g/
TRYzmvP4uogfY5FB8KtzJsPIFUgRf7yQ440DXKjwzNW1KrGsxyLDP73kPjhIxglQ
X4Zqrob0RuAmWK2pwk5ncKo0vJE+ZwrFbq7IcAoDxN40TSKo18usz5VRW0SMGEDz
Zodq9b7J5wuxgt2/RA5+kM/ComTCJTO4/d/o7gQizuJBldR5rVSTmim+CdE8680+
CB11D1jrp6J5QOQlyVc0vhDwhumNLNCzrfsjDT9AON3BxNAeKejexW+zX5RMqN5r
nekq55AlkqKVDy5Eh1DujOwjQHyVpETAI/oT+Y9dKLFJ1VS6wEr7jDFGPOV+6xAS
HYZhPEhQHK1Jy6X8J16y9IYi4jkGxYRFzgTVVwGmr5NNe3HtTOLoj1RIvVXKsnzS
uWq5xk/pPwzhghKsP4vzGDuk1FgT0/iRyF9a1jeo/lZgrxsbAxnji0nOjXhHOLhl
U+Ihf4xGOYIkvgNwD0GBavbySYvtiE7wgrmqEsgf4BJtfG+O2HUkxYyK9bXTcs09
RBTu25b/A47ltq5Tbv8U8ph51/6EWtagsBkS21x1083AzE9KWgOtW8FCMdyOO/A7
nhlRUJJYtzuNZ0sm571PxOcFlPEfIGjqCgchcibOIKoqVrI3j0IyBiGTVvS84Jaj
mOpYJYg8tk4ZGdVDEUZdlGBRx3PYSpAca0c7/ZLziJyyEYEXnZSx7J3HTuarWZQ4
dpo7H/f29dIFw25hMyts4JmN5Y+OiXWnm+5rPMadHkS+lZglelmI7pwEpfZFQkAs
S9e35wCi7KPzFC/y13iCHxPzlli/eYGG6dM5CBYkv+2Ll9+zmABMLvyFijltDtKF
PDvx7FjZBcv9GaHXdS6OepfF//2hWWdz5vhCTvu6IkOFJOWkocVZIR2QG2b8al0l
Tuhu/KyrAQ/ltc5XxTiiIMPHizjN247mN1OgimqoRNONEqxJf4Dx7iwkNWaLPHrb
z22oFL2N4PD6VVpp/6b2p2UnP58kLZIROijB/P/0bh9KtSQh2hApoeH99uMgz8/s
t2LERYVs+RsuRsu1YBE/iEVfjkm0enF2QwnxkDBQBzI3Odf+XoXXOeykrQ32iv/0
8EKl0QWdeh6IUMvjJdavISL4kG6vHSUD6viwIG6HYhsv5RbhWiuhWRzoh4XDLTLX
3iIK5qXNrw8AfmEQm+30w14t75jKPwk09WFdV++zNDRU9aYT4N7sb3PGjE3yeiWA
AAktZd4Nq/xGRiWMxxapdRK/zN6LRHK+E64X6HL5XiiQ/+CMma4O2+rZuSNR7bKG
A69q2F4lQHce47hdaA0DwAZlVHB3aO/3fOsH5nMivQt8joAwU2kKTbS220bSqfUO
h8hcZZjqDxPwEv9vUp5X+GxpJrVSXg+jyk8KL8/fAjSXOJbahskjvLSkHXidKY1R
SGiQwA8Vz+iak5HcF6LXputYVlO/VraUJNlPoibrNEJmUxJ0LNOnSlUlIlKWZn34
L0/mc3OhGZ6jTtZhVk41YP4ZcjaeL2zG1GpsAKnwlnvzimi+imvu1zV98/X08z5R
9RUx64ANnSGlAeuymZlevFzpcjky9L8lVees1ea/c8k2h1if9sC4M4AUruZRWslj
bZWAiq8tWAY8+EdiloKHr1LsTKkJkUgi3noHWnP2bkeCuMNN11Dmve5nlGgGiK8v
+N0ic2+FDdyCxgms/FgQv0bII+FjekHbp3GQ7HKwfb2rS5L+FvTmiaq6EGDPQmXW
wZFERR2kX+VI8xuPOfGQVQOrCCRsIAvzPTd1fBDVqAWsAoAf74IE1P8ejk4HFxIF
7QHsx47v8Gy5uBKdlJbtXirHzuyY5nFM4HMYJfMA/fxGJ4yvU5x/xfq02biJUzzI
MvbRIqHmOv1jHLeqoKuQYiOdd7RpKjKj+fGxO8ymFArZGiorICbLWZFPD+3DcIbq
Dr//3dksIBvVkJNPP/HTwmCyEY8sL/JvnUvnCNh5ypyoO+frPwF9qv4+jq8TcAls
ZwsfW5ubklOtsz2TuUebhFYPWdmpPk3cxHJRrn7bRHbM5GgEBqWqCgS9pftgSj7t
dgwJhYs3EYVMdoFiAvJfnpaLX80OosvtUvgDuuXknajht8MVhqy++/mrFqs9+om8
gzv/cAKSRu1fZxBj3W9vex4ngHMUujSHnvvzx1OiL+hnxKEWRdUSmXmLzlDV8u4q
ITX3MT8aLBMZDi6ilgz6o+Iy1Ccq4HnbLe6iiiAUej21I6SgyDm5ulXaYKMkdcil
kdf3lfBttqR9QZ3zBYyaX9oUIg9nhDx9Mjc7GyNH656tuKhLtnOGbkSb1127eWkA
fGED+FT/cJkZO/4z/jzv+q3+BuIASrgKAFTXCOMtHmbFGCU/5NmW+1q/wJTAQca/
RWe00kht7yt9vakaGnEay8FheXxTHXVxYNLfZ2VJ7ke5Vut5vwV/gtJRuPE9yF0v
6zX26THaHRk2IkJyBxd6FXYJzqfCX24UsxPFSF48pPj4tf43VJEgakmgQUJRLQl/
rEPVVdt6gSva7N3QOaeaHl8M/tS6Upt/eYgavIjCHAlurNZQFtIdzxPmv3AIzOMt
jV+c6GR5sfxgxzhWoofSgQrpMG+1xOHQfHYbJSZlvAO9OObKqfr/EwsBxQllMxvn
tQmo0Jl2n0cpIpy1G8hKZejb4tpFzkmacbnVgkwLZOtA/6In1qwfY50FX82gh2sw
Am01bo8/oK9oH9WLDxHs4mvSzqUlKTPwSyY9riTtyTOFTxdcqHebROBojFLgcWcA
LpSWQWZPalojnIZ5dKf7XWyJkl9uvBZTfcLue9qHWQqDnT42+XBt6UipZJRcKQV/
mWib/2rzHttfiu5onB6ea4tkQ9vi26jknwf/gtGLCmgx5HNKJEx/VsBI4ZTzJUC/
7cxsXd9jDl50fdzUpGMQxAahHOFu1V0b1Yy3goJKYFRky59OTaAZlRPzB82qi1VA
O8qAZWY26cn6tfLYbV+tYcqoBnIdwsNH1WAaH1cL3VJ3C/ep8qdQF3FxS4Fxe+mx
o9FdKzbaFIPGdpvYKTD9I9W2W7zLunvA6wmthV6EHIUtvw/XREOxjjgwv0IbKfyM
cfzvlsTqHWgmNqsmEqQL9kLeJeqDAPGftb9vnibNVKtZmXPiCQf0PQ49A5BtLZqe
SFaQgtAE8PAB77Xd46UwibsjpnJsgBWA8qq0J0yanMeheFqhkBT6E2Zx2xLAmV/0
Cofqp3QlIeCeEGvxnCp2XS51MSXekYF4lu6CUMpGni21/+HWcGWIQ4O9qBkGqSro
NduN5v01z2mSROTjmt2lWjyU3/oO1e7X0+mw+L5XynnN/aIx6dQ9gNQ+Ht2FkpRq
BWZCQXOZPMoNBAUvL19uvHunz32dPXT11iw/8cLpdPZo7n+GOVoJ7zFdc9+zrydZ
YcjxxKSo7h5c5uIH+MzjcmtFlEOMq8kmJ90T6BrGmtuN4GDH2nP+Rjt5NHbox7yt
tHfQ96qcg1Swxxxinu5dTJUmQvUw6TdCq2jPAI0pefQU+z+4XB0Pz8Yf1G3shgGF
A8QIfVUDciUqm17YjwJs0i6zMtVIwWj0b303tBMt/fWEmZ3HLQb7ZHd+XvjHeWny
1q3FLvbwILiybNZhIazd/lEaLHxLSESoZ/6E4YxT2l9UC1xRxJaBt5DwpKUmIi+B
kQj1digJ0ICB9XlvE4CZXh361kYIKqudfxCM2MtJsygWUYbC34Qx0kcKD9NtnBG2
2Mi7lZZzZuves5mzzWhC3DsYJ7U6SWjCUrHjRatUnG58dQiGE0COLtNgmorINmVp
SXb0Q2Kz3VtISAv+lbZk2jmANRf3Rn/3rqSS24ibbeidnFkUeApJLwlRh0uNdrYE
4Rf0ED/CmjCQ1yXk5YMiPccQyhFNg/BCSOs/8IVsJe2czXmenM7GUJUcaOLxbU/P
HHJgX0CScv2X0Q/k7m8keEw+5y2vVQohWFrMCC9g+m1nlnydRbjAMY0xc5o3xIPq
Q54tVOjczx8S7oilJaiJDnV15Wr6/44qUDoLwCwJ6qZVXBxXOcfNoCP7BYmot91B
lq78bQ/EFL6/p9D+s9V6potuaaAkKiP857pDIqoqiTlumXc3KLf8G+QRoFYUv7Fq
ko9JLfxnFbePhwL+91fI9n8ZsayAp8q0cfn5B/5igvUfA5MqNlMwguzI/Rz+o+4O
elYHxy/0EuVWbsUZlBosRW4DHT2moreHiGsBRQLGQCM0jKYGVLUELjGK1HCng5N4
wRK5kILvXbDKvEstRewJDKVFUBCPriR+ySJspCx9INCCVp0ToIcdOzbd/SU3Wdgz
X3WKW8FWAtntUeuKqzvZ7AielxKAtssr2AQulctGBkQfZgBVU2JGRfh/Q15IlhGq
IW2/hvKu67WkiZcwdmS5fkfkWIG58NjnN7ch3zPJErWtqwvUMqaQpkWp6/i0Dy6J
PTgg56jOHe9XNnCJZtGjhjYsVa+X+3duzb5IvPFsrYwxcaldAOEvIDWtKC+x2JZs
J1iPPyJP7FwyOmu5JlVtHAdsu6/4bYKDaA13G9jiVWML1VvADPIHuJ6RzdLE5ZDE
q/qOK1ikV0A1Um9OxoTgyD4YhkxRpH+45dF6POGMwAfkaJUTAIqXHecSnndP26Pu
MDqGV7+jXIm6E7PJarumGkBToV2nlMkY0FpMdO7PfFkeTUyCsb7nSHjQg/BZm3Nt
s+mpBZGKhtV+Ll8WJ1lRdfDyJcjom/ug6fEYqsdRlfKUb1n/rQVVyIK7HNYRwSOz
qdzSphhY+YsQ3USaOJLVuSCv1Uyac1k2vvmQkv8Pme4UaxX6Z9gamb9vqR4JE87P
mGfmkJZ+ZM5wLMY9cUNZapsftdEbZlg/dcK7p9/YAhu0ez7PwiIDlJTiwWZTKlNs
WQIXCWGg3Q1RY4xKyAFiduRvCUibwWewlgca6aTIlETK6WMlDSmxJsZXQx1KbSP+
LRBD7/rWCqSRnG20818YLKhgu7BQTnkh6zbgwxG5IGvIKj67ikjLo5PS4RBdEYmj
amUvLN5kB5Z+wcg3Qo87FPyFTAQgRjdw9uVgIHh0aUJn9jqu/gbpgCW9GXsjbqva
w3vetAVPSslu47opv6KeONMtyd147XEn0BHGzHeqCfKJhJVQW29KUvYOi4vxwFiV
KdDPTmcB1q7UXFW2Y2ITA3eevE/dwtHEE2N9mke+UifDLMp3cLM4Cq4Wq4TnMU3L
M5Q9mOmcep25MEY7tu5bSTKxYQn4jaBu3tkm+amyrK0a6gebjW3HZvLiRUG6jCAx
P5zMaCCradntRcSUcqOsWOuFAf+haFiTA2P4n/2scRg+v0DzyA3yAJlkBvCd11CO
ibFQELSaEF66STT51I02Zm/Mnbgowm2aM9j/xvTffBfc089PaEh/wqUMLiy8Wikr
wrBwzbWu9xmP+8kZkRpvafEsdU8k6plpFgBBvwDcT69gGQd1BKEX6VboRFVpMfdq
5/bcSKlH7wO7ZIc3zwxvhtkvsbUYoovsR3OSmykjzow+1rrXV5tonM09wxo7C7AA
Ti+XT45zham+FS9T2sKhlHh2x5T7biNR51eYVf2NaaceKa+Og7ERNeEKQpW6lQGm
WU/zvf8/Ulw1utG4rqNUMiW3jq7ioXyOFF8DnVo90aA4Yt7jJL1ykCwJGp0lZPxJ
iCHFHQuwWXR7MQGrf2Y7F2IfArNfco1WzJeDTuri2xO1dU4I3CwmREiqcxlnITJr
HZohfz3lNwi+kyPcQLXLSHnOWeX3Mcr7tysJpWjjENTP/hzXeToOyDNrNEXxnSOL
sgwRSxY9VEOpxgyJtKJEcg/BtVG457yvXrT/BrKVopGbaua5WiscI8iLTG+ii0ir
UL2soCYu01oViUXYosoi+Dk1Yywme2eE6U5J4MTuEZUoXBBnsF5Upny2MyhKNzHM
UaPmxSe6szGTZPwFYeIkmS5Gy4+doZDKMWHF9AY++2RN0CDCjd+1QNwUvjKRj0ke
Vvgt0myCPi04tgaucMEWBTdFVO+jsy1XEtLF4C9vMI30BUIrn1Z39XaAktuvGisg
ntmRnq9LUAwcyg9a560UKxIPcY2enCrQZhm/r0kv/XCuTOe7g1u855XTiDXONboG
0CY7RhGiy7KxPp0aHk+x2pDfq9vjghHRFKH4BTdAHtGBsTbG+9ED7h7owfh6ioEq
Zwcg22xSq0zJtmhChpDs1K3WJxg25e0Ja4AAfKZvF4Y8//PBQhS7TYJ5uEqBA9Fv
lAAQSK/ZYpBDfhQn2yaRVdOxtR7G1RjDjc4TROqA+hlHPByCG+WuW46SyXrbxHgi
U/LRxDfCnF/BKqUgEoXSgBaAHUR64OjUqQvd6EhJmOMTSLqY7tGZDBi2zphYQ777
LQPblEPcS1f1fgbIW05iDDG409yMylV4MqAKS6VUIdRrCv3eydDL8eQNIp7yYPzZ
dFybaPXySooR9voV7ZxUXm8Y0r/ZP7PF13vkjJGhoXh9aE91nCCPE3zKSkLUaGiV
qNWGAlDyv0P0doaW2ZQ7lI2JExMPH4Fa65OAqHbrEL1+mWGtBp3WolUdhvVK1Txg
so9nI+1I/k+0P08QQFK4Xj79XExD1CeZzRPGk5qZF5tl/FsBlaTc+4FTSNNk1zlQ
6PQzJRzWoAOKFoun3iHBSRRr9kqdqfJI4fggW6o8Jag+boIsjd+yIZ73rtyoBcYL
wJQdCRBYllWi07GoPkUWxOyIeo8lI197vbU6zvy4r0tP2c8ZKzLag7SBMJHENuRU
aZEhldvZaHI5X8hwc9aqQs/Csd2yWMTpls+VJ2BJGO4wLAghLPP/cRGoVD+5LSWe
Ia/RV9Fmp3W2p7+Je/NowCWGbdkzv9LjpGYpthcSQzaPLYm9of+U2tdUT5XUw2S6
cz0yhd4CT+GCFJMdmGGTEXQMvc9FAJmLGuC67zBmZ1EGI2C3ZsWvWCk4hZyCzH8d
TnSjmTRrw4yDDSjVTv9xXWQrgKRnCITKm+DZV/Mx6XNRsKBHoAFwfzWq1XdQ0hYQ
GlMLS3juNHPmwTINmHfCVWsRrRUAcJbfVJYewzp6u6WD3EP176irReEgnIKWaqaD
7dLEj+wAwxR5oERlwuJX/CVGvcm5sIc6/vfIQtQPoV9OnAKcqVPKN54UHbvNGnrb
ilDKkZqYVUu9KSfx0460eHwmm6s7/J60QB08BlANmHIpEWxnCp8mWavt56i1d4UB
6tOGwi8sKWghMhvKCF6RVe4VefaavG4SlJi/W6WBbjEFhECOs4lrDyxKVgQW9pal
B2yvw6G+dyZ456FsUcblMxpkfP5sj20SsLuIcyyVBjxAwQ/bfAWy3K/bhRe3ndWB
1ahjGY1R9h7QRpnHJrL790FdEOMYh96VmifhW6yHUrFIlMF4dAmoVGshtiJiUmv1
piReyKzq5Yohvcv5ywiIBsier+20yjQgaP63QeZM0PyS7nJtpShDWevXRzS4wYkV
rizwDP1DkUBIO67RxIUKC0uHia2W5YNIUyVImMa/cckKgpH5KdtKLxlk4WDPUuUW
pTHjuUweAVNKKwaJrdKarGB4l5CiFfDsCp0/9RpuP2CVEmLHmmMHBNJ2Igz9Eo/P
hwGhe6m86YsL1yCM1a4JlFyIrPYFzoTL1PFPwk6KPyjUAjvcI+b7V7q0n1LggHjg
HBWDfszMezBYRbg66Y7SrZ1MxETY9+DROqPBun+4dsqudeE7gMKvVYOGJWsX+jyZ
P1HWwvvZblg5dvoBmoZAgzcAhqerVajrdq/ebeHKoST7DL3OznMMuKe7xgPfmdnf
ouQWI/VfNlZfNrCJvYc3nZz+LSKSS0jPP0hlTBQf6p+HuncC3U3m/DjBhiIYozIn
3O1m702+lTsX+493HpvkRIMa8EEEf945eaDUcvXqBAJdlsy0hyA+s6vdltZHQP2W
tY4jCIqEZ8jZLbWhkcsFVr+Q0NolAWwfMrhdSU+uu/CSzhQX80POOYkqfnI15vV9
yEAwIiRm3JNKpQOnL66t/I5u5+A0NAVpF2Mil15RsdQN+lnTv1uH75Aq1jOV+Xm6
URlQPLCN0CbdNCOTuJpE0UI0GDZ9D28dgprBbmn5w5WmFEKtdBFdB4jDWKB2PKy2
wdJSSfzLz3RXvB4PaTH2CTXBBT25US4+PoWiEawehAoUwNEHTq1LXr1m/h3Xe4uK
Bicl4mJ7wd0VrXKFHkUI2VuBy6sgq4up4+cSO6w69akNtgcXvFwDonN1fC1iwd1E
z7ZjcrSxvnuDxc7Fl8MFfCabmGx/mkhILGOkCxJS/IgBBRInuwPQCHaw2Lg3QLNt
rmgwV+rKnUQrHLQZBug/rtYlDK696sniOp+/aRTBpVFTCHYMIYSCobTftyyPPq0g
cPabEB9XhxThYIhCPm7mjaDVYqoLqsn/E1I59sQRqkEpOaRHfEmxOpp6dCycnYHk
PxO+5R1HyB1iF71ofmkjEHIehpiHmAqVZ5pYCH1OI/HA79fdv8kkpkgNWYokZV3X
WPtZwB6ImA5Nq52H/7QumfrJSl6CZUupX8iTmTUWJoGL+RewAxCFSd2qMCTL7VBL
0S1sG2jBYQUcLPT5cagEuvWx/6V3lKG20xuJAu/nG6kF1B2DlUj5FijwinCAPJN7
tS0OVrbzwcsQXSA7R3mTO8HpG0J3H+IL3US/JdJCfKCRRAnmg3fZQWx4yQlCbixo
WalPygkaK3ix1ovODHMLiZ/tAcF7Z8tVxeZe0cCovtfKFPJiUdryUijaVj7q0vwa
98nDEaWMuXoEq06mV973gHyqk5MqJqOh9kpY6bRYs3n5qUOmdz1skpkVqcswnrHu
rzkTT9W72ywbbX7YGbA+5Pe9CQ3Bw4jb7UL5DkSi99x5Q89dkiOsyVsedBZLm+0q
5Tg87IFKwPyw7wnVUI/wnUUrW1f7FCZk2zCK/xHxCdo0LdRSPB9MrlATBfKrXgER
uEJnFRobQ+iQJuYsF4GqiAhVmDgf4WOqzGPcMdRNDTIy8X+kSIbp1sKXocHWmwS8
HV6RGwfyWZIGzEhpqJ7MnZJ/6Jm+22luIBIhY1Ql4zGhWQ+BN7946C7DHeJ2kzsR
p0Uit5f2lGFFA9hik0Xn+z6NMc7g5p7ASbhqrAvXu3ZSg+VxhCrY38Ji2H06tNC/
qi85+dcL1AXJo9GTD3uKRt7Z5miPoFQqBi7WOAEHrL962dSs6vV9BzcCLJEO6EEP
xQwpm8vdvtt0mDd4Q01awbO28ab46499LnFFtVr/V3Kujfgdnj5AkwIYR8Lh+xfG
kfxMl+o8Tv6FaqhWbjscQaCIhpqpjvFLYPHHMU2F6CvWujDXriiln5Q16pZ2WReA
CROvMYHHS6X/bfmyxxDnSpD7tW/E/2gs3TA+xrI6ETkU/ZL66VpdrYoLnBo1O2Jd
w33FZBlZDHJ8CII9jmwz7fbRaHk60AL2chwP64jxIWsEMpOK01MQXHFt/MxWNAtC
gatF7kQr2DkK5/dP6ZcIukJdZ695DtNOBumfewdPbBzFNjZkI1q6UKjE9rM9KXL3
0mFXpByvcNlBETko0ePYfuBFagrHD6UB8ttsfmz/HN0jI2jcChqJ16KfHD64E6iu
yql3ClQM83p16xM+yg2dyNFqeGGHw2b99Z/6SN1xjTGPYoySg6KrNT+sXkfVuj1a
6sPHbkR1dbyce3skb+8pjEeBiEkoI7lXjxcHTRmSJ8W+MPomjszI0ma97hnJQ+Hb
KPOGMy9+nraGAYZoi2CoDrS9Oei2MVD2Z5P7CcDjwmBwD6d3QA7e3CejnR982auJ
pAPSUvnIkts1MtznOTFtN/368JMIDAU9x+wdKH+JKBqC332tc2ghZUut7CdqoAWa
d/YvZoicnaQM3o0x4GbBrHnHd0MQSFpnjc0zSo1cAFWCd0FVlKyiDTjprBP6z5+H
WjV2gyewDTyZx45qrJeW+z2i7UVn9H+nA6tPVuXQSSwikZYlO18hu7TcPjqxhMMm
8Ec6qsBDkLTPtg9l90wlgKT32CvkjdWUPqJ9DLErWdoMxXSPMvHIzgwd3VFwmHQn
MfsXZV/NMJb1v/LflH4i/K+tSOJvxkoQ/F4iueUVrYzEdyI6sv62wSxWNG1GHhqA
hu16vad+0vEV3x/8G42843ZCnEgJJrlSJLZvVRZTLIjHSCl01QwqdhqeEEg9lZKY
0gztiqkoYnVfcz6a4AOarIbMZgwzbtXZ6h1esJYV5g2kkqPYoqRQSmcPzLbakLNk
TefIiyLilgvbIdljSkHkt9/En3iY4RUFV4yc8TP+YNTJbPPPWC3UEgE+3QNOGWMh
DZkO61kqZ/bEJHbRfZ9JyfgdPkbOG/VQ1XRlrnL7fqeVqLeiuKYcWjNghow9tn0U
eYzFjo5jAcLt37qznerFUBXgRY63hukAeanBDPS5NIrAbk1we+57jDnrxLad6H+J
pMOaspE6EbvtHw5ZAIZnK6N/FY4Xbu1JwbKmxSpZJCJurlEhcbwR2N2K/usjDgq3
107kzL/cSHzQxIqOgXPpQQcEAlviWdGHJXZkbnyPlG4EZPKix6bRQFCgknXsqFFL
AbfJkX++P0dR5GHZ94JdHopiTzil2PFnf1nIs14ZwX5j78bwKWkdSviuOkBrUR/4
VHZAGsQBwK4qDIzvrwDMJYlD2N/dUDw2hpk68tRdLmA6Iaaduziuo7TYNWqwuYzN
if6TCiTnlk7M5UGGi75TO7WrdiRd9YlswdbAyFjcYNMXsRCNz5e/3d6e3SAvJHnj
tTCxxhWWQ4KXAuorQkgwJUKJu4JDTpg2HIW2By9ia8enhWiVjk1g7596ue98WXo+
TdU3fYFV+ogMOB+WYO0T5po66TraNyx8HxDwqla9ePBytkxJWco1KJ431rGAIwz/
fz2SMLsKN27FQHscDzMowemCWPYKrTzslLBE24DmVCORtrKo8sQIoPkwnLSOPYUF
yEkhDYEMzTA75zjulNR4PX9DBQ7d05x2/YMgx1LygAmXbe23Ydk6+pZLMet7cErh
/3q905F+Jnm54y/1ddWpbI57acsnTKQ5Tr8EVHAJSNfdgu4TVP3h+vAbx0Lj+aLX
DR7tAFC/0QNCpmQ27JKvJnkbLaAU4gUcP9x3rTWLMpaKpCSgkPT+AMf7KkYRnPSY
RohTd4xRxBwXwqIpggHf/UJVnjN1bA1taONWAtI7YcpoeQ7tLUo8EQreSb9oV64r
OI3vPuhyjvMD1Aqk4+0EIv21CUrvfRAUYmSb6UjGM9ELhs7hDUNa4uclebeSVtPf
aHaTe7fiOMCcn6S6SX3eigu/dQcjg1G5jpmdY7zOOncKTgOBTazI0ZtB5JPemHxy
3QSNvi6rDTMyiUIbPeDj1xREND0zullUpjKdklU0k/dY4BDGVeNqRk+Vx5hz9F03
x7O9WfcUNCPhjoVHCT+2sIlyQ0LZA7nNb2nD4HjXJvmbYhpaAXYIpzTgPbwnwxw5
MGaI6dfXFhfuc6MBiEtohimZk0E7kEwFi3cf1EMYqKK0TlwDTWFfYVEgT9jHAmPA
EFRYvzCjCBF9Wf+ABK4RDPWqS6tarUOGFDJCvo6gZv72BA3L2AsLCeyMzOXg61Wk
CWEbpppht84h68xjAUoWhFroDrfiNZlyldjkvy0ZvRRflWl2AbmUygu5dgKXtpjI
YotrdGNjEmgdY1DqPDuaGjIur4QsVUCnCzQIEgu8qNAjWCaq8NGATUVIGr9DlMZE
vHNXGVFwlKfCNlh1IjOI8YDtp9pBhoZI6iLa6e4tSEW4uLVnIeK3Uzh64AHQZuOE
3UtuJC4VTK/T91M8E16Ncce3LYd9Lzy1Ycwcgzp7n6QfOpxt7HBLdnmSjWJ7cnYf
8QhExD15PYhgZ5V5/4YqTOXkmIfVCHyVucJpNKtSEhGxsLCWsU+95IOjvaWdHz5K
oDB2XwpPQAt+JWW/PUhFV7YNeWfQXAy9dRuNT+n9RnEZOwQEhhMbOAdAeNUSUe9M
+i2UoYLmTuSrmWeGdE6o/Nr4bjuIRZsMKErt+occ8zR+IhFnV3uvvJxB2zCUVmiF
T2Ef5Dla+u6AOxT8GqrgnQWVUCo3paRLoyupgxV/GSYg/vdrwVXUFuitOzq0ASbb
pZWPcah3/vKk7nO7coFhcKuneNWOH4xahwD4GhjdNu/0Uz2ICqdStl/QGegLX1EM
BL65Oozxbu5gIBKX3apFeFCPqEi9o/72L7qr9a+TFTCc5qGu8rq/GAtT9s/LpHG0
sXFfpYWyzxiks1WxXjq7zBODX+Kici//TMj8LKleDxiFW2Ej6IBHJJs+zr5s33VE
v09h93WjeQQ/p4wUzUtiiWvBAltpo1NKznVGCP98EQtjLqpLltrx9yFuHwlPQdVE
L+lhmjiM8j3PtQ6gdNwEjYQ/IsuH33F0mWA7tPwES2wVM922LG9Ij72biUFzmkbQ
hMDSLfrYKTMYYYHAuMUp4UCIrs6WX3WJrwCT3mHtJgPEZQ6DhIpKYKeBWXb90DzT
0OeKMpglwIPzAhZHpryQfWJOZB8kbX4UMmjWgzo5JqG8KPFLocpz3V5+rfjH4c3w
Fr86ZEW/gsXjtpefRfFge3KqPwzo+MKfMRR/BYEddUIlTvbdU7/ZdYZC/LIUYRGd
f1naU5N0RpNmwvaT7z3LTid0ODJwOLaTfp1qgttasMEzBfqHthoKRS6kD5TZjxP1
av44ACi4GuCgmAdyAq1qFwNovAv6aOJJ7b7WxTyE8u3vpwt4CU3/k2Egfik1hC3R
qx/ewA3SDsFMS2ZovXu63bT7I+GnPT1m4eCf87SXxD9kxOqrH9fgi4iseb2sEUl4
K++Nnyr4mkwhFh4hyyLUhRj6kF6xxkLoAkvJJq4wjg+h87J6DCDivXp9ozx+Qvpg
rk15ruDI4wbdq4pOJ4A+u7kuuCr5khDIrXxnn8n7ZAutRPtugd9CJGmHH+Dztz7T
Jgpe6BeUV7aZsOSrG8gVHt68fBozMTZp8KpHxonnl/+q3aDY6oOK3wU+G+8m2z1S
jD7/BI4FPLrxlcKdKf+RDfSOJ6XkoMDSQiilhA8HjWUT/a5A1hgpz/cMDOIxN/0s
1EgQVnkJh1RIhLBZ01TbJ4cNzUuBHskoy7dCqH6gl4d+dSavCsmIUGxAqtG6CyLN
y+aSlQUX6GZZQfxaWdz3iKKSGMB8ssVN9WfuX7O+Cbs9cqTSlhZLK2InqAdF758P
wTI9beypPE67dUuJMvMQKSH7NZ1kxRpZUQSqdRquv00p/ICWSE/TeyGZX/kvhRp+
//zt5234TIELGrx2yPDGfbExjE88s3118/Dd9+/YiMsA0iYjSHu7JLP4k4V/Uv0W
DwKFFDUbINUnabC2+i6NbTSkWo6viwON9TMuXWX99LQh/IvHGAgGTuWMVpjUrP8y
17qBJedTYextJVKHhIv5doAkInogAWsApwzZz2/CKPdKl/FWv6WXuzzSMMx0MBMp
n+VEN6QUFhh4S3YAO66DOIBPQGaifZChuw6xuiXqRt+1rk0Ux9L3ZyryOYNP6NBq
sGjt0md5Tp7VQDbUi7vw7ZB7n4BGBJMA9oxHU0427ZUDi8ZEalnbPaphGwZlSJ4q
eomlgb8IIFClgEVfqPqm2jVr5d4OWDSnl/ihZNM2AFHndx/DQO7NtbY/vwC96Rkh
mUW6P8XWCFlcGJDpyu2OBIoblmi1zzTSR3VzdYD26a8XzU3YH2YPgYf/PqBJqLOu
a1Z8FH0qnLABSdDDF59Qs3JM6Hh0s+hgsf61hZwUZ+yOyAQ9oN3lPkfGD5xwK/o7
kHt/V9ks5rT3b3ynBN0eQD/YFYcN7SAZVOTGKThSc2z6k8CGTwQh/fbqs7KWLAUa
x53JojKGk5XSk38gG6BXQ8+AU+gMAgrHFHvmfZK9EAO0/+PZ0rxKvfwusRt2TY6D
A3ZD6RzCBVAAbBgztYvOhV3fndW+hsyrEOVGBU70wDKX7KHUSr7BDp14YhDEl7vL
zXMe9NWAy/huV7DNLi3DKXe1LjIrUf7Btrd+HAZmJBLr/VKmHtX/VUbEI/Ofhey3
B1X2aVd/6+SIqnQDU1hhk6xs5fRTiBU3fpLvI9f1wGZZvtzYGv+CZWoVYSbc3ZHx
fzB3oKn+Bb7/zJUj48GkZzXLvWG8NrnZQbfhrBQvC+/HPaQkshe7NFqVavkbay3c
8+ZqUJnAJE2oxewpBiNT0aKgxMI2TxfoTLiN8/buUkQqO1x2t908zTowghPEsI3R
rCD0MI/qyCRyiWhpea7PHuTvpzqBeXzIv7TvUvjQJl36kZwNP9Xh7qLaI12TP7D3
oKL+jyTJBBXz3trGDXMY/VO19EcQLywD1vs909kSkWH7bXRdVpQQwjyH8DpvBbxV
UufL3X3klo65XYYVYlskkjPiwq7KRO8ygJ3w3cCMYUYQ2rUBI6REK1kIKnOz4wyL
5FVPqimFanuf3cT9wS2a45uBWZHNBmo0alFX55WienDhjeUaPJeUcgEv9iVZaTuX
XgdIMiS5vISTpqv3XuPIXqzRAOPUaf601QVz0EiBerV5BKMOHUpBSe6dHXn9sc1a
fyuovbI1n2NWb1p/jGfpGT6k+sUY0f6mSRUmszlBxUcHHxkLevg6cjCZ8hWWxDLu
FGr/QLBZ9eN58IGMBBNLmRDYviE40sftzBdM4LxlcGzixK3ecekLB7hkMMPtSrq3
7D9BSMGbS71zKlXptR1347L8qjcNMiRw9wcjlViO8zwvI9XZhFc57qUNIu8QR+sJ
D+HTp8WEp0AtV2XbiAfXqBk7czm0gxSDWq0TxCZPb+2XCs9T9lMDCP39TnP26HKM
4GiYs3+ylKXiX8nZ3vsvd8qEKLxP+FBTBdHEK5u1b6zq/dd4WcO133jHcAziMKlJ
ju+YlNw89C+q6Gy+4XWIgWoaf/LKOf1aVitmF8RFFWwneCmrNoUBIs1pdAFaleeP
id+M+lUUh03V19H63+k8oVkeBc06XOFxabUKFubGfYtPWcAx5sJS5ZD309qnln+9
4n/4rFZiZdhaA+5eTVeQhVgA/b3bKElZ1p6fAEgzRcbxUZqE2Ka2xWLoq6wO8VDI
63L21lKycqLjLlb2uwKY0zwigXrcaIHfiVV9eM6+Hxvmh75kGIrK94izAOXhIVrb
tl/gVN70+Phk9qFaG/K++4jPsI3V9cd6ab08FZoJH8xUTUXPaaBtSqahvjfejJGh
NY8MtYvXRgna8knTRN+TvVepDA/jKHCADUEObiG1J4Ny/gysrAQcrlql70bWio+n
ErSRG/bi/ifduxp5i1hP3Bqq1i1N4f547KZgdwNwhdkpCODlI9jHR+psSbW2jA6C
ZROCJbNS+5frwOMWWAC4HpDe54a2OtD5oyWCWNytIHvGGnzSHJ/139wBwghhoynF
onSwbArgzEtpmAbA5yJgPwqYe69r3v4wxBchMKCYKvHuUKsD7QZ8JuaFNeqUTKbb
j3tXgw3oLbY1Ik3q4mjqfeV3goq+v1Fz5nufKk6t2n7rfxFfelKSxwvCOeINosTu
Qik+MfFcYcoRdDNrwxk9+oymEWxCxes0Kw+cMPC0Hn0rRZfk1bbjUSpO7uNzrwsl
EeYy0XxitUyWBc6BuKv9FvXf/CaMFP/WHSPbPGfIF71lRWDWKU3gcrBQ7XOQsn21
zOGeC92GDt8c2E5n8smneQhzG/+SZ6ByXHGpBqpPd3lgQqd3nGPazFgdMckWeA8f
YTkCSC3oV09pzQQGQrOHP+JIV66eCE8tYhtoi8qP4rPTM/6eIL6HS8ooTlsJOSVe
N6F+ynfnJ/bnil9K7wTB6KQvGBRLNA33k9rEOyDhwBtTwVC+h8EMFdEjJK0t0STv
6bbGk8peT1H/XDxazNlevhSi0QMXVFleBsi19EU77EpY4yzfx2M228vaesrsAfg6
WI1TaU/igYqHSdynyqnkPYoa8AfxXW9xFOU11gajetZrhnWjRJeQvrlfyQ8piHSy
kfrb7AU5Y5bLXytcQVWwjBWMIrz9jV10KeQ4kIGPYIPMJDQSgX/JH4uglL1qCTKI
LEQrVF8/NCnIjPNjf1Xohyu/ToqALWt0z4sKY2NCzNhDbj4coRKUC0/7cTVDbhvO
AtyYv8fgCvHbxqZwWoL+kwfVm0i6Hnxt2clDSyukYDnJXFZUcJ5/YZGvPBsFDe4J
hXcImz6Op1KgqZ/NJAZNPPSdyO1TLMJiJBpgvTiFb19k8pb6id1XI4ESPzP1fZip
pT2CJAbnGOLV5yvr5DHC8fUm6yPn24Hg07USJDAcsgOE3EEv+/VTNR0z7vzMsRm/
RF87NIigxNytb5SSzvpHl5mQj0Ml4uWGWCqFiuBSdaWZtRoQzy5icS3wLPHbaUdd
PeSv0g3Rs3/KqYLoV/MePaWqksO18+M7OcpOQ/xCGNuzBzBaAfXD9mjPQFLswSY7
DP/sUNim3nr4F8xuFf13jmAKGtxNbZyJ3UO5MpdS7+urT3pUCTAqo2wT2WdlpS/s
pfs08DeAVRNPb2X0aqWTMC8hpgQVmL53IJejZk8pSwPeQP+O+dF2KcU67FL/oY12
20Fi/MY2qU7UxsExK6YTnqXVvgl1x8t4aId1lhF1QumUAwpM1LXGgfleqMnCOawE
VqRFZrfpJ4T6AMpL/tFI7E5XsAr1tcKSBmlxUJIWFrvY4dCjljZuA81UvwmqFJAx
T0fh3BbyH1+71RHoA1t9+KZ8cDCNXLtVmG42Fp6/gARPpWTUphd/2MQ5Nv9Ap/q3
0RxJYcMnSNUqtPxVr4fc/bNKJ5ALeVnMiatJeW9ECUjcLBgNVTS9NXjAia1fJ56V
wAyFQN+5QjSK35uZWadOG7+PeXmQG6qVKvr2xQrJN///9H0pp6sMWFf9ugPbVEXg
OxfZHjC4sua7I70Y7a+8hwGCUEpMXNh+UHFzmD7QDcLRYkkzlFENkWGbAJPmBNVc
KG+27QjUW+Jb8W6ASTdtQOLiwFcEy/+uMHw6Un8WfmR89OU2barWUDQV9OwlagNN
hdQ5QzMreUd6UoUEBwIKbU/nlMUwvjHT7mTwfpaI2MCWOcKUyRuY0ovuql3Zjq+0
1+/eZqjbdNITVNXA/JfwMTMAkkNu9I4MYNAGH+U1Ml2nLcvHkhCqXLCnLr1puNhu
oP4Y7wfAt2Ql1USn9bGhrI+EqGqK3ryzUhlNbPGqEVa9qN7aFuFL/aWnBg8LMZ6D
Q8mDVKwiUdVY31IU3hqg6REi3Pv5p9p+zcahQNOcyTC3S5dqelYmSOIpl2qJQKJl
BBgHsa//qrooUw8eXwhFMfl5SQyOJoji3luzpX/zjkAiyLCug/K6M403ksaUU9BU
TxTYOgq+k9bXv7bbaj2mWYpBV1EL9LUXMuoJuObfF7kCw8DF09DhLdxq9cF2BpjQ
5QE0uplkYuXRyI0Io+LGTQNtSTZNuXJuWzs+Tc6mt/ilvVm7aCSmx5aosmozbyBL
rzxPf+/0o7SwZtC3Mqe8vl/HPv8Kw1a6LosGezK2mKU2dCLzvsxW9cIYxQvhnuMT
/m/hKmGCdiaweoSuWVOjb0aU8Q6v3naok1AcLJyENwpwkBYYO073oba5g/f8iEaZ
ScV+MvYq89e551iiGul4Q2EM07Uz4Fm63nH8Ic6YS/2PDCI+sMd+jtYLNbyt2qVG
fm+yGrCPEyAp/tzi1mNW4FGxxT9TiWYTtSJ/90RiTi5CDZEJ8jrWqvykEEWggo6M
pNfRGW8MbhC+a5y0RFlo4xoDZI9DUvM0l66Ys1GDAzuM6BYkrasJ5gRROYHP62OB
EdxJ2+0jE1IS5Al4GWMWxHUfl24i7IaawP/nE5Yb5yPm8mAVUx98S+TqRwMYrrph
luY0QakT5YGddp3nNaoZt6DaWHLd/0w58/5CuE8d9CUoZ2UXHgrWs1hEwTuTaR62
HrtcFGC5N+dR5uOHvhB02CV8hyRy4TgAcHMmq7bMiLWoOoZMYGLMnSBHforswpVo
xqEIQ2Jou3/PHSv28DBttsqL0RfDXDe2oEdh9dL4AwFsGk3RusuO19pyfnP111Rz
sTq4Ikgjqzov2Z/tjCuTAO5+Yi/ByoqAgRblSjD83bKiCbv6VLjBWYaI8WQCL26g
al3SbUe2JAL7k5hYcz5HRGgVxbUmJTqBdbtfVGT6oe54gCNQlahzfwTvyFbo3KuQ
WHlOrO6FPfiHwKZ7FYl7evkn0mpdKwb8KTUDonROz5unKJR56jzeQFp7Je7anaXR
ldZXgKjGBqgUxOeZTZdcCVqXNNRJrvigBUQNmJGNtfK2LpGWuZdkrx5iG+i0GVf5
5NZEX0lu7+Vl5MAU6o1Pd535jdyyWzikoyZDZEfCgMNjycTAjmsAJmcOkkndz7ww
I2fYvNSA2LSJwfO5Wi1BtxAP84XKGBQ4a4SYrSV1FlXe3JtGSxovTJ3idgnKNMC2
OoUQwTrUCjEEsi6VMS+Hi4GPtDWewoTAY5opjesghUmaYVLuR5olRfWM7WCIlvJh
vZjnH8PvaIBOxi2UOHhaRsuBYYRWJV8OvcF8RDrrPWO9eeCZYQsPlmr6lP6ABCEI
oGZ7uqk21Y3oTv0XyFYud7S/gXkAj3LY9RjdfOn3MqnBgErXExdmkr3UifGVn1a+
LboMgIyGAiwFhF8370/0zzMh5mmRHekNQKLKYf2NPSljrCctmqfAeHdUhwHlllgU
9ubYCPWoVxCgAdjPJpv7ro8+Y0im66Q7scTyEpALWymLYpL9Noe2gmUUn/lrW3JF
tMrgxu65nUNJZMkTzwdn5YHJ/YBFe6wiSDZwDjh+50aLEV0uoWD+WNNVSeaNQsKr
Y/M5yuSKvOiUjWp3VqoSf2ylvaY9VDaL87sOTeVY/dhTgDlZyb+0kQqANfNorGXG
Ft6hD5SwN+3ElS5+N0/s+QXIjBzNJG2G6K/tp8//ZIDnVvPH5eyHoZC0Q5Wa+4p3
ZQnZ/+Dem2kQS1cCSaMSEQPtVdQlAc2CM/8hJH1ieuquKCn8VYIX1W1IMhowLoan
f3yvNNXdX1XXKRAOMymO0nDvT97VGo7BhSdI2eItqq2A1i70y2NB969ocegO5v/E
6nZnTMLDsKrQlJ9Miqn1ANUIwH/901dmzgfQErBwaaoKZ0hmEkq7yBvrlcynTcFm
heHRmQLLd2XszSFssMSN7ti1reCTRsXWbpMYGsv1FtNDB+xDbCp3KY3T0f2Z1lmp
lJaW8cnby/1H5aOvx1uGlhvWUbjOtwwsQZMapse5Z07iT9xZo5l82r1ODsEPYdGj
rWBcuR+AYDcPGJypPOXtRMh6quQ+O5o3GyUJstgfvGy9huKIdAGmqjIf5Y4sou8m
UTPyOLMkCYaS+Uwrm/acCKnj6/prkuDIMmM2LYEcsWLk8WUwMkvI4DOTuPkbf/ID
jgF7H6GchLnI5ZomJXnvLGoL7bUitchtGrXCV9VLB2dXVfQRg5vtemWxUvR+Tppa
TW5ULunXwyfhoFLhHKmlZ4ssD86ydck3B1abx+riKdmxLamFc3jg/DSO1zHZ3QUR
8dZXGyidCjpcqmGCgl6NpbTxvsiQ63GYTyTwcvzKKf4Wv8K7ycsXUOCWqXePstIz
RzepYxl+XK1NYQz8s7f1qoYWeQ2T/xorMGPAC+MuMvGJZ1GtGOClix7ZkMdEMQyH
FCr6shwhW/hmIQYCvoK1hwvdgGZDgneu4PFEsOD1P3yMcBi3KHywEKo/KNqCZICK
q6rnVVB4iDjTkrFDbflE8bMxqgR2N0qwZqP3oBvlXox15jSIaMG+kMoR5lOaS7Vg
5BAIq1CqNqNAWnYuDSyboRLXO9PMBupbPITJm2RLVI57Ln83dQqzEnLCl3TdrH+e
TkH8g80MThk3t9KqzRIipSU85n3nLjCJUVcg5xRLIMjJgsZb1XcGMc7/S32RlRnu
HBiiCcBze/8C7kNYvnkqnvTMzTZfGGla+k9hsX9xyfECFH/f8pzwTcfjutXCdXwm
coJfajt7tz/q1/F3wW26YTQldsKHlT5IGidTbqX44lJ2GdIvKPbMG2YsLUL461Kq
yebZM9dyWE2JiyTwbcMDicdgZoQDOJ2KX6xq3VbLIj229xmLDMLiaNHFrOORgGc/
7Rhtd8ZxICR6JH0vBPE/c+7WSDy54737b9MEervzB88jDLQxnCjCaFw5/0yLPYQj
Uus+y/inGnPYrwE7S+LqwBtYi4bOSbukEDA/D6JsIan5SoGNEC9S+cFH/h/CRkKo
qlfRVOmqJiEPnY71GIixhX4iHrYAbpZmKeEKQm5w+AwEWjlm+9UHlx2Y8Ml9lhid
O7tOwlbbeziGyWwIADoy+dnoT+TPUFqi7OPFleGIFHn1OfH8HIEiu1fQq4RVq0WJ
5dkN15z8VRwqmrXcoMmnD9YeCZm19k/F7Bs1lBH4CfjZxmZJNgyR7NKKIU5aYDhA
X1IasGMGiMpy04d2iHX4Rn+FOtg5RMHbOi6hOBCrTRYPxv+PObWrTisZheAhQTIq
CIck+NXWhD/0tgukLoBOF/DwTMSOlewy+ODq3R6vlhuCnLO6QqTpXT4iQL51S/jl
uaJIsnvqExEinCHqFUdG6HqJ2JKr2xGvPBpyAhV0gVHxuJxUQoZGhVHgcbQaZHgF
WNWZX35DcyLOEv31xwVeJrPuLrNpvuByrTEAE6ufiIxN486SUFh8IY1FIK3gcjWU
cHpKssyZUaELKROldTXHQ56UpwjmCWXbZaKAo8brymYqwMerm0Z9Avtf2S1mCJSO
pHbHwYHiqMcgBAW9TS2RE9Amx5EpT6rVbYC/KZVcwCB66YsrLne5cBjq6VZjIDuD
fbfGK9SlcDdTvqOZ3AIZzQdsPoyZLuJjxWAm/Ei2GIztilqmUkyuNAVFNPuBEL9A
2+FwtrgUb+Bfj8uh4va7BFR6ekIEx95f0aa18z0ydrz5C3m2gLQT0P1jHS7osgBn
zysGos33eNSXS29GB3iqm/kpe/KqNU9VmRwXBZUjs9XwzAqReWTkuoCyH1FlVMRu
zVv89aM3RmLjgk63ro1dwjSfldTIj2VDRKBqpKq3N7e+yM+jp6L1wXUVanCJjQZC
tGpkjxZoDrHS7VO8sQfPVKNdX3SlYLBpgmJ6dtPZPFz1OkemEJ8sHJubCJA3UtNW
2aarwaVVoQjRH5M58XzjgkxBqEdeJu8xsLomoGtXasDA6m2OeCJUhRapGOCuq19Q
EYSsfR8sjKbTCR3X5IR3CTCpP0Hl//iY+n/lfkogpPvbO38JOnrSiOiGQOckoiN0
eO5wO3YFwK/rjR/ChY6luAgC9KwvNIHbCGAAgV13igwpkt1J8WNUqGgZa/eXnwsO
zG6O7ONB47C4hPcJ21kKGlricGm6EAQQEKuTw/MKfRSX2SR4SCjzV6NvXsqFbPHu
0lk1cotW0nKChEo3lA/1q98RtIE1vnpUs45Q03LdX0HowZC1WNkc0ucRJB8Lp12F
OmJjwQnhuSTfsf1rMCY8nnTBMIaL4DGJGmMWmouvrFPY4iChQL57ilRrgv3ebpA4
M0jEj1ep+hi9irw0VnhOk2e2JIfCfAv4iqK9G4GNiihIDBjJHyY8KW2NKbUCKukI
YsdtySCDWY9JuLz6QdXj3jIG0c0tXV4uu4lUQGwmWU1r9udPY6t30CfHWgJGoRU1
rPjwEcjwF/1zXV1MIqx3Pj0ifKyNMD99tYSiE1hMtpIbjhQB+3f8frDz/FPxhzE7
Tc8MgCWr0xY7kilEdIkeOdK7KULSUPhdp1iHFy04oFKToISdoCMfoMoD5iQe0Vre
As/CTHeva9hVUunhn+e3k7ZU0C+8Ja7fzgkbpkUXmgaU6kQyeHfioy3kaqL0186Z
ihx/EEX7Ta9kUr3jRrWD+Ff4JTfDSfolX1ZkXn9krGaaydHPB1X4EClW8T7OcmbI
E/jTixMCyGGt7ovIy/WQbCyXJqv9Mm7YhRNsMcmz53YnDo4rdfC1qIuf2VUSHwgN
zX4R7xgfaTKRFu89B2rLSkn1Csy5ok9gEEXnQ00956CdSBsp62U7PU8CgGPyvJgV
Joya9988h2egi0jSK/1XyIJcrLHDIhGpisdpi3t+wMBj04rHXmsBWa7gLl4owlpK
ZjTuPRRVfpPm0rhG35drTLK+BN5ZPmcj5wcfQBoltXKuFpjmYnZyXQbE6PS+ekha
Dh8t/n+kBBp8+H03V8YpdkX4VYP3XiGXKfJ+W42vLe5jZDOHQEhJHiY01fzVUJYf
xyA92VBFpNAEZBQLiEaPI5Mgxiad2hz416aDdCwKJCMhJXDH/eDUJfTWjP/OnPqR
Nksw1zqRCEZuoAM029nXLoGw3LxiX7ihXQu9JIK9CA6EYL8Go38a5L13DojhL9Bc
Lf44OnSEP8tp1UwUaGaiFeZpI1fI4S9NcKCFcSBmc7k4kccpZqa9dumx895fp349
elBIhI6gYskbbZ1BWsa9tsLgmCeFxybYo65IaHXBmxQNlvD5o9+DXMN839qjxdQM
q2iOVDKQSvbGsDQHZNlYSbEXwm9Z8l4bqolXpLad15AKlFD0A7ePzTfV7RN9O7iW
amWDMpjnW4UDHdRKy8NWcklb/AAPgfY/tIwHxHMW1ykfttrs22m7S4HfyEcAqubD
Wb0ZomFfUDTMYqBv4ysMsm2TWYT28NZgk7TksQcHbjowgxBX8A88VpsQBuIx02lU
Tnj1+6PuDRB+OkPRziO2axb12iGWQAFkHRU4I4Iey1tjsqjWLTMxzO51VkJuRadp
OsnCRQv3xvGtdqyu+txC1wZo8uxxYCKyp6XmioIY54+aSOCF5vYR6k2QZ2UH+fQf
Rh5YSJilRHAmWcNLHEJkhNlhvwRi56k7ie1s6dSZB0efTJt+GSHupkxVdE122nqI
+9UqEqJ58ITq82GhWOe9y9nsehIehJ9c+ruih87JEFGc5WTKthL0nPfPAhZ84XJL
r9j+2jwEMNeCkpPOMVz6kOavUIejG5aWzqNjWo9RVPtFWXaXCgbcClh0I8QyMrj5
QQfBPk6pE62d4HknQv1CwdrhaoSil7rDJopv1kHw3glnJFJ2sQP775SJ6tJ9JnVn
q0QdInmNTjCNQC70wys7lqN/CUuii5tsw1WPXCE3sPvVl40BFmlzmXV9kev5asxT
z5Cx7unfPsaQiBG7qGC0hqPBEYz9P0x1VYpoxWcyAC13moeq3BnVA4DnUIAZioBr
ZtflaL7g9MA3CVNY5B6s6oxQFXjKCFaJPeJHSNLaXHt2hJdhALM3xhcqEG8ng9N5
TjU/TIHPYycGesb1G2wnww3an0bL3tAj/Gab4+iv9HTpMzoVjFopzVysdEsXHasy
K/0AN7xW0Opbi1NntduORguT3nEszNOFPrjpMc2xHBwrxJJnIewjuLCW8JYvLvxO
pJwUXTbkA/9TeZE7cAiB4xH6CCKYk/y++scMC4FiDU9yxfyqMN8gbGbATuTJ6Ghc
oCNs84+M/cM2sikWWyKH/pz3UTbTokQDEh91ZRz+0oRGJPlpzNw9W48p20dwnPBg
S1bCOq5AGfS9fWxUNYVhdA75sbIqK5WEBN/WJlYqWu1nmnOmM5v7YPjrMbKwRRjG
ESHHcq1BZ//ppGaXiy31IzLm3on7QZap8yBvzZxaLzqG6Fgii9dg4Phe5lZXWOMC
4MIIyj+qfrpOLO/UnMwVe0T2LdlAckYdmoPb0s18uLb7gOrSQXr+nDY24nU88AUx
OekcO3hUeya6tZK1pc4oNaA9xRIXiDSQqAsKff9iEVZPG8svtf1mg6DOUUAcxALF
ab7GbNvLnCHYUPOQZAPqBwJ3UXtq99ajm2SfI359+BdVbdD2bGDBYPcp4IOIfWrf
tu334k2hxbvVyNpBdLI2jRVEUKs5Bffvc6AImKmpqj7X10spFNp/p91LQ1YTgSUD
E/fvMVZhzYADFJYBUeQdsclpfk89VtlHR7BDvO1tEFkei7ML0tXJOd57/4zckvIc
9fnKn6E3eoi5dJoFt/GbT07d1v9AFbPHJCmU5dW/yv+z8SmUrrtuxtWKYeLr8dkf
88u+7Nz3PNm/IkPmgT5MnfkTbThjzIfvAHxjwujqfG0oyGkRmjB7Lsv3BeTk0Gpa
d2tXoPC53tYgZTT00wvNN1x0jQCw/ygVtNj9M4fYkIVJuSDgY9XIk2rio+UrHQIy
vbqZvN+nZjZNq7MiDnJ82xZ+hsIg4etUPK21G9Cz3SLYV0eQkyeEASiLCeIvera3
IBfCW3E3bJvQDwHU5MbkwSfuzOXDA7CDSq1uGTAsUbULew6clRcyL9+0RwF36aS3
oM6//XvyOWEyVMJYNQvRVo6I9zUmr8//4cJldz6rQxdN01QAoTIDJhm1yPoLsRbV
1dpmeXwI6CSFy8TaeIqHsAzKp50AP0LUmyHmLfe83N5iaL4BamEtHsBGxhiTN2qN
wCszQMiDAomHgfA3h6IQ9mgfv0p+EJ7gMIeQuCKRHn2NtHmK+v1B1Bh4QX85RR3T
NJvMnikvbeEt/G9NGrqruTk36aW77BblrSlveQvq84T883d+In2ElCHpmg6dksjC
VaWWjlVBvPHHjikg/deE+vAJ+Kx7v3TM2wh+lewX6nLMH1P95ncv3GXpLGfGq2F7
B9AW1EPOEDUzgy2VeKOOP88oKiAoiFkix6drcWoVUv/+g/MqVL7+O4q+OvtZ9fta
qtY3nAY96QHs+fIuxwX0zAcLkuW61qLVhIE/a+owp2UhtCluHDu+9ICM8B7w76cK
p9oJR4C1mbp3iDCmxKMg7mSrAUZ6vXhVqtUUjcW6zpbs91gTNxoFQECTsUkVjM3P
SDmc8cozUCetRvW2emDyb6BnBEF9F9EWLmUHMYBdAoRrHyx8uBi9rwQ9jnEQfHr5
sMf9jg1LoKu8zFm7eSb+mDSVvRfyppsAm9ulIa52zRagKezRUDA0c7bkGKeTWm15
Im5IuY0ggrfv9fB+MzidnnxOThFoBxBzugx/1azPJibD02qlzR3FEk78VgaPFz3w
2Axyj9mcVvgCzPjpscNOQGT4ZDuc/BTCQLu/YMvXLKAKZv+4xYE4oZPG2x1mp3nb
8dYxvf1xMKfwM1lEd+D4WRYRFHZYY03T4R+1JDnBVEQ6WRkE49sX4KSNZkd5M7Qq
BNlRPsV+2OHqC9tFN+kkGIGb5j/CH4lDgPYWFMDouNC4CytDre+yCSRTEf2/Fz3V
341bsRpjMcUgMhIOfFSKKDGLvCNNY7wHRWOtCc5Io2gfGiGpSlnn1vQ8cnWJvDX3
AzNlzrivGqxaEYgqM62eyu6RdWj64jQO6M+i0r5NzFmt8WfFqtJb9rbJ5EgDJO0V
k+gD3RW+OjJCn7C1wYoKlm4Y6itXVDnDZYhcdC//NvoT+xr8x2699GPkKizOkKVM
6nEeIPxbhihMv5GzJ5u1VFH8GuBietOGaDv9kMf0/wsHeTiY+ifSBoD5myqUcy4Q
/xemw4QrT8smQNNzOxcsxZQ1yEC42YmCVxUA6P5S1/mE51N3QIHP6rIkBCURWbqn
VPznkzREJ9vAHP3W2kphGplgD76a7b/fZc37WyEy5OFECPySzAyATcF+ckDP3cGj
sD7iF/anisNPNNeN0CPHFbXdEwfOS6hlVD191ZPT2Kp5VV3v+89TMTKwq7Yh4yan
VSyLPFz40dHBTLj/4kZsSKRO22tXsteWEyAkVD2tL3AEPLaiiWLBhsf7Kef1KCsx
myCd16Xlxs4hxQes/OiyVgsrrx0lDWRORoIGb79lNTx4iBg1sHEeJ1YysfaVlnyL
e96JM9AbQxjmAcQwToKPDicn87PMZ0N/iIcoOWomCVJQ4ypss/HH64y6tEN7+Mld
E4HO3k8jRN675e7He3FP7L01WCD4kEnOUlF2m3U3lQiOxjAAxFquJkS0kdqmWAPG
LTpIMuZDVCRcSgNW6l/zsRxlkttg7snXfUdHUcjB9tJLj04e7eTyp5DHV1rWVUkN
yCIHTI8pbBfoHsHWETr48ZXIKtIlIYLu01x/uhHe3u0OydRE87MgMDgbWpl51yqn
N/HHOmkRa4uVN7gB5M+X5vUlwOYJ5WZzEbdzLuMBH/ZTfgN2t2Ld0d0LFZyDuhsH
1r/HALeCTaXK+FQbdy11wqKJPc4RpO+ljG1yGRbCi4ZFcG04uLeRJsbAjREaa9pA
39QVnAPJ+xAeHh1L1557EzSXe0fcbjAwSCuoWFL5llYbD/Eoon0L2eLLgffYgww9
t1OQeuEsYP9+5sY9Zk4vgKEXR2V9yhRuR5gAgPZCnnMP+UQWTPByJYxmqlLyT760
j8wDn92LRegpF0retn9eWo3/La6O1fV5I59cMtc2Oh0iJvynRIdYM/YKmcyO2qOF
swsKsmgKFNyPKBI8rwO1WO66+9QDfLQloFYG0zqmDN/oFCXfI9Y8HzNGNl72WGvV
LYlbh8dfShySFoe3uDonzH8DrdZGOpguE6svzOgvccY4MZ+/vxHtVbLqeXQAmX1b
iqnLg2ZYT1Ujnyf42I5hm2cteGB7qgppwJ3orcxYbH7zRJITFgyifb+aJ+Xd4vSZ
gABsBe8V/vp5PRFsG9IYLeGJyYqcIdKfp5BBIsi4piqXvEpVX7Pv1P19oWCeb4/A
QCgYr4ALBLyVHdc2TSFoXJq7O5aGDfpXBJoRvgML+JFn/bGq6pzWa8wdlE2ckLN3
ODBGVlxAc1bzBoeOC5G0DPs0+ZLjmWwdJssQrkEIzZGlEplj06s9u7Klxh8D1VoF
vL9+Gc+hT9feYTKSLX73zL3DYMDtz71rpWZXZbrtq5hQj9e7eW1bs89hYHz59x/O
OcsxtzUTRScBNxYN1Gp/4myFQYNepOyUQVx8gUYjRRychr3LRBtrOIVdgH807Rhf
V9kgKxRl9tlkyI0WdDcfGhYEAwLuWWN+ITiI4/z+aRwznJCgLn4ZcquBcsTrHqfm
qEQBzb5tbH5n5csegAkC+VKPbxmT7a16/kuJTh8ilJwbdiRoQiFBlg2Lc71sU1N8
GqOU9iWHhTzd3uzOlmlAF7YwXOXtraTLfNx0OQm0+wT1Byg1HLwyZK6MQqXJOksZ
j+32NaIaRf1YNkZjWK4p3sf2UQ8kJl6nbm7efaxxxbKk8B4z6VjiFuVCAorupgg6
dCv2jDI/S0B8i5hlv/Dxlp2mSDmqRCpELi9MVkwa9q5yao3RCNaWOWWM1DwCV1M2
3imrCMMraBf1nA/Qi0nBtvHCCeweltdSHsWBs9YG+geW74kEmM7xxUZh1nRdN/vl
GbvGE2aLcjVuhYpX6ESgNI/fS0rUNyM4z1sKs9d9urfabwziRZqhDGjsRgeSo7vt
z6zzI0RF9LUp34dVoxy1ijyoGt7/P8rnT1FIIGnfkMUX3l4U9Pq47e0jmx/0qxg7
A+6VLe+AAB/0LnKbvfKJsJeSENASEhAe6+F4fcQhfvzXk7mRl70vg1lrdnZwWXT4
X3YkuJ73eQpSFeHnrbipf5WeKbzEQDX3bzG2/G+W+dCVsGNzqVtvqSY6e9fjyEUn
TNqz3ouHBSYMJX/EaM3o0EZVLp+5+wRjcqrn0wjAAvmBd4I43hdjN5WaxvFKsGzk
6XC9s7/GD6r+GuOxo0QJLomnxrj1iJa2Z6NUW3HLw4JU8M2CyDtYBhun4cCSZktt
WVMpk5ZBL95QT35eJQpQkJen9f6+ARbcxHlH49khHVR0EM4u2U+cMfLnlAVTXkTG
yL6CkJygMF+4qouvju+8Oi4Ll4NTspmsQofL5oNyrjbk645M6GgHUSlS3DmIJTsV
xfkzVPVF75uxXxPcKv2ucL51w8h9P3qtmf9Qz47sCNScYjiBNBNuwDxw8UFHxQja
cdGzPw8WodYv6IATtHioFXEMNxAAHO1piInVnx3QDeEH4R7G0C14N1K9KJmk7APR
l2vY6wZmJtFFSS9j0MLxqcY/W9lelG9KF3E55v7yckB64VnNiPB5vgRRY0imShSv
jsODG9Hq3neXxaq+cwnrD2GEas+IJIRna8NpQAj29GwuDFK8m/gk4lO47nY+Tme9
W1rzDPA5wRTJQT/NJRs3TGGJ2RcLhVm1x7drtDmD/2/a6Ft3aPJzpWbKzvxzqSe3
Fi+a05eZ99QD9ulPni9FWVmuHkjxjgLcL1gOSlJb7u9mmNHgCvMzzjE+hzqNWL9r
zpoUnl5jOM+DGo0b123mjQKS0YI7pjtKp49Sy6L6b6vYMShIIfsG/9e4phSvUntq
9pqlz+CdFPm8R8J9+SLBNPLcZruLm4sy0BbJHy7p291ej53EmlAUX3Tko+B9Tkc6
m2x0IWo0mpJnIwQZ4TJWeP9b38GhLepZlbrJa4iKyvk2SIY1eKZgsA8rdDaTBe7z
jGnTzO9vFZiub7zZ/KBvKLYZQVO81aV/RwzlyVX/mKS0ONDK9FoPXpDa0m3vO8n+
0C3JJO2eJmOBMbOeIZOoTQ7zCzO9i79dymcwK0veM+ymOHNeTOB7cDwkGLUSuMFj
l1gTJJdM34o/7af2Vq4Ae0AGNUA22n8+9ZA6DfKdNaNXcEdRJyBcSLxEpzme43DB
2/pHYJRHekfLbKdyopqy5GyS4tPN8zyRDjVT8IGXlrOXtYkhqahJdDt1AS1TQ/nw
kmKmDK5fnQN/0n9DxmC7wkeTSMGc13kpATwSgQTsG6n3zr6Mk/2N5mZSFG5rFAVV
R7KHksTdECDHzOu69PsqOhi4U8xaDv5YTFXsbkEijSrK01In+wguCiePRqbd52iB
hGGbcCZ/aJOzQSlUGVFwpvvZsaXTVUIRw1yr6Gc15bVyLrkaDOVij21CuuZCZs7h
Tw/t9VU4f3r29hJtsrz6vHL2RPc4L4a7CV/RoUYZNzlcYJKW3Sav5Vp9aGA/Xxph
I1nSPWfsurcZELIGUkrOcla18do2izjEOkaWh2U3/qyf9t9nfUXQrp2p6dXGn7OI
sDDow8RisudTFazjV6+AnCaAhfOKFutPg8d9Rh8cxn9sBkO9zkX+pE5HzZarEois
gpakA+/V4oPVNwRJjuEROWY81bohBGV9E3u8Gcv6v7EhR+TwqfNEaKfonHN1Gtdb
l7o82UKyErT7l/giOAZb/kf5VyIyxE5O2VPXHzc7gNmdcfhRP6DBkFW8scsjfo7Y
Ha1tV4RUQ9NTNYKX3ECX9uPthmRtZ/RU7DCdej1GMHF+TAC5uRoZlzpnjkl6ZL0K
ErDU9XkZG9eflgEWYNEg4MBVPjtMMl3QmaLz7AP24NxC+GkCWXtg3k8ll03dfOFW
xQMRseIwTQf5yNsHvxFWQamyAb0YUIzDvgfxNs0g7Lqi5B6jPtvuXvNEEw+abGYu
vpW3awcIGmu2Nso/tvfuIK4mD3Ln98Zul+/KHUPr/JalcnU/g9KtIG2rCYtJLpU1
WH0OcD7ST52TvmYH0ZaKmK+WfFu3vifCdioR0gVxtms+u/atOStRe17bPjGhI+Zv
fsWcsx1qsaWCZGDJGGLd1X6wjkUT9oTyOMRFLJ0eZYh+sp7+QrOI1EkCrMNASZzG
UYaEPizuawkWQlQW5fh1T+DRA/Tejvi/V1E2LAE+K8BkAr1XxdFvnm6kyDZcYRNx
PEXP5R8fmcI9ajuW3GP/o9HaoELH++l9oukgaDKBWVF2Ggz29rj8//LerRWB3XM9
mxZDMcCqmk6/yGJo/geempeLx0bkyIkKNR1VgpRHe6msBK/JxwwFFD95E9cCgbBK
KWdc0Z0ldI9/85K4R08JNCEjb5zsutYb2b6yvHVVQu+SiuPTJ+/3IDBCfg8By0Zo
4jq09QQJqYQBh+jT9eUfkW+eDp6EYeUrmGiFYigN3PJDK/3gkd4CaP2cxkJT/iCE
tF2oeT1UdOgtEzj46/YvFI3d+EofNw2vzY2BG7MpTsKLFIzA9CxrMwffAHAUAoEH
eVeOYQsTF/LFlry/bCBTzL24dZbcKi6F6CotEgXA3ecTJ0g6w+QJ4K1i2TqsneiU
gzTaRh5WlxUyrUOz1O+OLxLNNuKGMbz3H+fbc97oQhXBngET34gvaryGMlqRHe1b
+xHXxMZOcatydS7fDyRQPSi2nf3UpVr7161AcNtaBeORd92upLRFKDw+00s4iZFF
8nl4TokOAo6xcNR7DcFB+sDYiwxSaTFX7BhgPoRVA9jea+j1a9xl9ZSkKJNBJAPs
zujRcau+hA5mEJO79yqy5Uvcc9myQxfGiCNAYFb2Kje2PT779i3vtevAzoZQOfmf
evSOtzzdZNWA2iCJD0lsTsekbQpaojWw0ByAZmI6rbWIngWvSzOThlkw+KdZidTz
PrMxch7YEErJs37TWMh4Mi691q8O2JDgcdCI7DYDfFP4DSdGdK+oNSDunfQQJdn3
WH3MWMNXAOlPI0PSS35MNHWnf/F7JrS3+qJbQXvix4SQimCP3FTZeSIvcI6K0fhe
CLD2o249IoqcZ6zUCa+satf2IFbe8RLhqlkb9mg74CFHB5IfwR3sL3HXZe5rH+IB
K1vhmHzwpDSD+/u0DfvLg/yThbEXhtCn0FfR/7DtQutEoBHv/a2Au3UZDx5a4qWE
Sg+K+8SsU/Ruglwc/zAyOpDI8/z0JuoUbdAsPV/ohL7PkVjhyGJNnG83DaW8qCSb
qUMb7RGRDlt9AiVFOQI2BnDumTNWtxkINm/xSB7gNSL5olUUIJKeSmxGK/DDxXai
UnXDcU4dYE3ox95I0jqfPiLCdg1h6I0lHixNXBtszq9/GwNtrNqiQcA1A3dVQBeX
a7JtF43mgCMgUvDtuNKoQAtMGVH5gYRwSq7bNI7oVO0jkku5EtvlwwLycjMCDoiZ
al4Z893zS0ACKHAkYsqb1hluXxs75rsW7O+aDehg50X5S086Vfu8Zdhl4gzjHC2L
8/pJyltX53kNa0GId5X55CZb5DrdNB2n1p/Q5gADnbtERhK8rBW9AZXFXwZX5Xst
gn3XXtCrJggj1UBpJOE886MTfw21cgai5yFIVobJNGAupYiEiIttgTxOpksDL9Rm
mG/Js9eTQGK0GoaKw/G2qyr3nUFTcR1LOLtftiXE6qzmAodsU9mkUOJrYrroh3qV
ffVb1AjZ+zzcMMvsXIdqXMsMRvuQCuemSgYogYwsFFmaRIQp6CvWrTakHynAOHYC
sTsoYoE7ZBv4r4whst2yfc2seWwqz6Xm0GHDUX3mVwHhXKRTVg2hWbOwApo6cxLO
A8dvx/qxICwkg7dv/y69nOPUq9/XlILcZ5BRYlYmXuTmw3Vy3EnH9WgvheGBGXme
w5RIQX1KdvniZH4L8ttWzkJbZvzxs53KPpV/TRDRB/tk/UnaQs0aBnMH7LwFN/RK
Xc4Cm1SDdJ6i8ubNPymotl+yhk3cJm/T2tmNur/sxFfctQpCKsqP0lQUKnDqrXjy
K/BcK99Z8wPOUFq2sIofhq1NBnOvYaToHoJBPx+KpLhVKx8Qivx0DEKkjzb5ZcQ/
FJiGgtJrksLOKt8ed4AcQKX13K66wwq9za+8TyzyC1l5Mhtsz7jWT/dlQNUD0T17
GED2g6JTUrs0HNIJFEH6pcMd9KQ/oREsiTg+9rvuLx5R3aXS+JWSzA7mdjbi5ZkK
sGRdXi/jZzqFlSqq/2CX1S7yjz1Rp4ArvzF0JPccFoOQXnbNk3J/30KUKl1pQaLk
HV7X+CPeYXURW9w3tm59W1d/IXtoqhNH5aIbTDPOY2vzeM/gRq8cA7Fa7l5qj+Zo
IJdIvtMxzJcqfepftkvndI0V5XPXVTD5bP2ESgMdtwC5gPlKy8AQs6kOGDCksnrd
49DWls5Lfw/85jGf2GTTTbt+3tY9BcBca/5On7BXLrXyNZy4kf6exqyGSTNat5cy
4mTTSYTL9VlLIrHPMMOHGhxaPte0mucxyF7CDQgHtJEl8kDPIMG8UeicWj0bKBrl
8pi5pp56Y/Kwu93DBLPOYLbHTRqwL3YWyD5X8O5pjSEVUYpnZSHT3pHGnwOLVigM
HFB5Ay7CAdO4YQgT6gTwFo+DihMX6uNyxvLTPgbttIr0iG11cqYBqmo4tQ9OiBIy
Z8+zIxZ5tKsqb5OjsulAg7K29ixnqh7m3+JY9xOq4C0SNZrIKUfhZXOE279fB7bM
MizPpZ6qEvK8hDmIr8kmfpc3XS1IVw++0atBtGdJzfJ80aoeschy+BA0mAdmUAEc
aPN9SvGbM6KQZMZQznvQoJ+LWGTLQqa6Z9v+deWK3AC56Gx+t3RJnTwwS1Ze+PAm
MjwMJWHgYv1aXbmmCn7RlmfRn1rkIU7pYB+342lypjETBVLd2A0ax14ytqPZrZ1f
d7kdREEHFXkA6Ewc83GeRJ4gwjMUCns1vwnkNXZlC6jFHd9o8hTNn5KQ0KFNSKqa
/NgoRet3BG5ryrcPo363TPK7S/cPtaptTzMsl9aSBZgDTI5RKlNwVSNpHSW0ni7t
Og71vNFyg6oD2930dGaURENxajiXpZg9ZsJ4goy56W5cLX1sKpjgIPRPUWdlLivp
OrcyvnCixlmgjRgmfnrvL62NLfPuirKrT3RSVUf0GUYj69N/tMq+mtxc8johReXp
SJpKY5eB193fs/poYOYGKfiYxFXN0fml0OgsnhzpDzDin2qIbJBbiHUZq1H9nY8I
F6SdLHqweP9KxC2WZGIiv4MnVzDykUxQiW9aNbb/rhbCtSJVLaT4V2C6XQ9fq+X7
AFo75MEpwBnel6LeP5hQ0WXBSOcwPDcKijs7HpQcXQs0rFGeDiSGUfQNCzDLOAov
LHuu3OGxncanFBRqmluYslNguXpLPzhstk9sxTnVLajTLou3BRqMuRXfdLepK6n5
JeKvm7EAE/h38Vu6dUQ0m0j4aTEwcdZT1t5xokBjgN4yFOZBgkbmS8FkLnPtZOaD
YRB2j1LhatCVxA0ckzZIoJEONj+ayrcArekYoYZTiYmEHVmf2StylvYx+2ub3nZy
jCwB5Ia6WXrdREowcp0ZrgjIFujsv9WdH4v/6DE1BpnMNXzdieBeC71UxV613gkj
MDw/K+nOeGlk7SnsnAy8ZmZRH9gCq4DvPdmXpa0USZZ1ayY9xxzMDO68lXreg/XO
XZYHpeb9pm1UZ7l7A/6J0JVpfBqwtaR2meAWCSdNKb0Gacd8Qg5q/0w1bm5pMS5z
hkP3GaE6XkbHlh3aqw1W7o7bvTQyYxSlCsVwTdOnMuDVdiLAQ0koHSUgfPsibyRG
7qVo2rlvWhL+DQCipVDXXUFwBCINbJJasJJHXKErT1kW87wXWVqxFwiJBLI7357h
NnUpf6dD1t8/ohP/0zl4F3vwjnyNptv11P1zkYkW08HaKI5kJqDjqV0pgDBVuRxh
1PWIecXsP3qHG2WtDEEkmNhFDjzsmednOvgKmVNvQfXwm99I+o2yMAJD1FDoiuVJ
yPdTdqiwmI++sx1+46Dor5sNRwy3tTIiq0o40EwHxjyL/1Z30zgAeDvNqYSJv5WQ
JCThgmnQQswuLZJK8h3xfSxf+K9IZs/uQOR5Wz6nNUdF5FVvWt6iYVGgpy/O5/vy
sQirkHdM8sA5eyz9DVFGbkNC4BGeT5ekmVoIyojWh0cgiLXy91ZlFmuQMurYwUTm
GyGv4rFc/7u3XmMj37iznij3w5THIrVZgqgqE6D8OYP7hQ4iQAmopXB5lSgRM2Ra
DfsYfeNrAUNMbLZUA20KRfzeRSoZZtrTdF3rrM3Lu6RFzh8vba8ppL9I4RBlnn21
MTN/8sFyh9dm1OlHGNni+0+i8BuQttqxey6y7Q5toBweXNu0AA+R61sEna3Ir/mh
qrskAL+LzUVWnp8wpt1eS/vnuSsu9k6Y6RYUy91Vy3H3lTrEkexBB1keKOGkxx02
O6Cpm2nnZD458R3NOC6inWAKblkWQcjFQkbQHeyT9Mhof061as5Qzz6vxlgIE1HP
OsX1uIHB2aLz2CYO6A0u3aP77iY6Yf5yF/eCMD666BWpq7aWb/Yi0tBZIEp+zMtg
nMWYcktwdGqkMe9I6xFD+rhWJjdwenRdHfCjBz8p0jXZ10j1SiK1B2bkoqmUCRvH
cCezJ+405gX/I6iPe41IMFrJNf/zP+xSnGaAtrJWCny39nywPfGSg1l1KTXLi0Xy
q6LN+KCmUwJBATfsAX6wHe6viXF0XaqjM6s91ccp4An4ymVn0zKhG2EWtyQs9Epm
gSeJr0HJZFy0YpBF1Js84TPZxQUcQjzDuaIWkg/f/+mStmMSPq4uS0U4Rge6/hnX
6xb1WZ+V8FSPNY4ZbFDD7k9Xcx3Mv49fb0JJMh/LewhNdNyZW9yoyNV8I6ZrOAX5
B8PqAWBiwuQJodqccirvGlfh6zrDdINEQOGGcVGnfnDysWE1rLUMIMXh781xswD4
wHsZrG70p4rZL5gpcIs696vsonK/RvKros1gg+hxGuaU5CmMoqTz7m+He8AHkg1j
o/tHvmhI+moZhnoj+AMN0UjCuUXHRvh3QkRv/XZMb2iA/q/Y4ULFOEi68KsJeFLD
qWBtAcWW3go+INmzt2rBidbd6g0sGs7pOXrz1BLtI+nw9o7qOEnf1vgbDCvfgrhN
iunBlE94q0YWl6R++zLV3bHSaBdkNR+fS5WVnsUhfBGqWa6nLE4KDpOex49iioTa
wQ3YUMUXQCjIc1QoHwpMm3Z+d4i9Eea5/wtvaVMgajdOx6zTDiJJlaeGLOSrBN9y
JvMURNxrLEKGtnsQlvE1+CPGz1tEo5JeCodPMjDs01VxBaGVmEgZD2t6zXGvxLrE
qhXzG47jR03ozVTPooxuZsLBp/+N4FKvkl++kgbQKryQ/TrKuN9zY/D6IFtngPNZ
PslA+ptqzluA0O2ScOI2tAzBPLbXrCOGN8wqKgaovmjI0xUPn245pmBJQgbsApS/
ZogMx8hAmIP9cPduORWdGcMAg67BPEdd+WgBM4PG19evEG5mmy+YFeUQYxOosPeK
n/cL1Qrk8EWQGw+Y10JmV7xmABVijtMOX2BiMUcaGqhClyyKJz6gWej+1EGR0IJq
oSpfI5oRid24UBoFtH58uxhyez1HX480JC2OwlWLbk1Um1kgQk9mkSZTY63eVgLP
Nv519ogcrAbOjCMcn9fubBfcmlQVm8jB8fwMPldR05U04fcLRLsjk/NVAqXOfk1T
onzt+WvVq5ps2CUKwudDr8y7luvw0uZBYoQOAB1ybxSVQmyqG6P7x6r02FYl6JxB
dmvNqDURiIaktKZ7uqMoH46R7XDo1bhSIJGVzrVdQ9A60bDnDJUTgqz5x16Bha6O
iTc4OYF9Es9m6+yCR+BWSBJVNiXt61+7B75WGdY9YH0FCGGY7Cu6HoSVVWQvYzet
VMG5a5H6OfisCAvLup+AufgZswmZmHfaVMhK4gQfwu/7KqNHBANvp0JoNsPSQnBp
ZlL/yJsM4grjTUdXb1AlZU3kdt+VhsaNIGEML2jJV+k17DZaLzPoxFlWUxmU5WSj
ogbyGmPfu9vnuwjNwzjJh2tn8xzUe8UlcrNue46s6wmMJ88FwoUpCOC8XCAO7c5J
2lC3QqfAIU76FfbT6pecIPosKOpOedpUYQy3jpFKHr1RsUQnxUo9W5O/WNxgzDc0
Jx9ItcOGK/tml0QEuI/kztDbjCrL7rLE7Xs9z11ATlxFu9nIQXb5jHAlaaLo0rBD
5G/fQ8jpdye8sa2iXGdN4zkhYNI97GxGwJL3fd12s23uyerpUxAajuWOmHkgQGOp
HBIlmuZcLXziTM1nsg+KduXEeU0x/eFTXTj5ZR4KFCQshjntbI7xy82A3n89XfAP
6tHMf3QOKqCtdS/J6YGd5nqut/XgJzEJ0KB8bVBZ+KAxntyCQmTJmVT6EU4xKFL5
9IXFWjR1N6ke0BkqA7KEpZTWFKqq3Tf34e9le6jic4Mep6CHpJfu/h8E0qjG1brY
lE3xeWqjgdjbIquthRao+qpF8YS07mXoDl4cjBhmF0DP7S+rsxwvKWZ7A5tVwRw7
3+svvVcaolnqAbgxLoHzmL1OPh9DitQzyF7xnzqJP7y4U1Jkc/P5LY+8TdzryU3z
vZgyh+jTb06122qovJIZD0m3Nq0maQWx4NVkwAQcLglznyLg4egW3NihZfevvpMD
IlZ5BCjawKuEnDzJihWKRLd3I+57HW+dg5ihNf7tNVXYtTUR8PaB0wjG4nEuPh+5
tYWhjp3VMOmvO3RXHaL39fLXqRLXYQ69PyptBGk/SJSpFE+AjTiD+i0Rdfg/vZ9b
zaB9k4wPwI9oVNpdSDr5hn1P0iGR917D/zabaJGF5UMkgMqawpyNOx7zOVIAfExH
7rrXTvfNx/C9GythprZPHLYcPVzfbAaLtE4uEAOExhMV4RwxofFDfF85Qn+Qx3LP
B6RQ84pUuzq4og9cvoQibDJOyDnqQZi8PUKwSJKtRcBhsXo7C20TbG6tzQpgxjqT
+8CRL+J6/Gp8PfIxWVxCNGoc2FO0L/0LF5OOI0JRDfaRUq1OpI6clnTZn1eGRMFF
W8kReXsu1LWYdoAqQcJRkC13RuTMiokh1VfOcmChFffuJrjYZM4y9+EvcCcOYD+0
aiAnPk30sOWPVlSpfQks3UzhJJx4ubHX1ZCbU1/JSaIVeaGRLMbGgABqzENgXe3N
GGecdP9OG0wI30hFKXqotFzzeZgpSQSybNAh1xH+2mCJYBS8lCctux418lxWcM80
Dse9T21e25H8Jxr2lcqFrdvZg7zz4yJmH5KobOE/Z5BSzEFzAo4cZ7mChBTCC4Eh
L+QJWaDSkS2UFhOYYKtHuYIczltvzYkTK2b741sWwUsPv5Yo3rDuPdW946Siars6
TO0GQva3MTaXA/UyR8CEqW9yPQ1DHqvoIbDPlRuvJ7r6Jq8Xte8CWaoxtA7SmLSw
UKL8EAfX9kvxPmuNNRPXs+4RVjtq0HHSuNyo5pA/6VvlKIMZEX8nkhZ4MKj+o7Kl
d3UO0H8HwLUmsK7gBpgBeyZeYDykceJbTnfCc3cCD0DxG1S+5s9Do0tsLwfG0Vrj
WEIHNshcBDQMd9V4wB6suUrecZizMDaXvdPZ8DDfTxVmy1uPh3yOv8JixUbEaHh/
nb7uEBCh5kYcfh+3hjhfh2VRaX8Ar5UR2Tkqh9cNbAE6kiSS0E5uOUtkIPKkg6sv
YSq70nCvg6MLMErOKFl4cYN2EVVbhIGDBHJU5u1dZTjz8KHTV9NSg8rl2rwhRWOR
8oIzxIboiJ63QkIrXOya06Mtb5JnNqcMYijIMbXJ27EnPew2oeIG5ZFXTlV6wHEz
/zez7/kokSdOC14BafM656EV0wj+hr1W526MdN4/Dd3kyLE2ytNhALpPRL982O5k
G2YvoqhieSlmg2+NNg0tvtX1r7UBCXje7sFWizx0xBuWZk0/tP4AsXSVIZV94xxZ
z1ZXD+ZZ0l1F6VbcB96Cchr21d4nVHvF2uRxgDGwI0rdM+qS/031Ji+6IwF+pfu5
1dF5pKTuoDrsE0wHbYCEw/3jCpCJtow41Ptmn4Z4KgVcXz4cO9WbD6VS1sWWIiQR
wHTaPvryU2OY3yMYMGsRUJU49MceUxn9u432Bzj6SBEEsjF0q5hcU8kWRbSdQrJN
HPuB7VgrC1TTDJawBs8QLvAw8o1jYJWyzkiDHZH6kB6eCgH/wYF0AEdF3tGib7Xi
tFTGrBlkIqfgeThimMPTXvB5TpvFfjyZ9RywNvavZcbYlC5Q2GoAhGGkmdF7uXB2
oOclj5fthRw2v5nV79rtoM0OrI7xtbbgnmCDnnprtivsDXY2fWZSwVqGu+Ug9gD+
MbcUzF4DlaOnX9eK7DEi7jqtH8imkN9V/tYHkyr6qDTdYumroRvKlWvbHnChzAXa
6D+VNFBkuXNQcJDP790znaftcH8eivmOgaDwakScLGJWcFG+LPojllRmygmavov3
eT/MN+BXi4HaumZuzsq8nh89BkE0ZnvDlbTgA78R8U8149Ha0lLPZDZ8shp34YXg
hM49jXtCTIgYhxbHADbyEYI1F8camDLJvOa4o5lPbcYE2NRAO+2R4+tjEryLaN1+
eKk3Y5r4T/IAuMKldbr/l5CF1Q2sGfdVYnKJQfJlZJfm0/AUenuyxPTgOd2mM74Y
6PH/Dd1C19WmlL9bPZ6n919Y6IXnMLuUI5B29aZMh0ivxWVl/7bAaEwG5PD9WmXK
S97A0JT29yI2HH6mcMivpKYNQH0nqcUEDcBe6O5x1Ma/dYdkmkppK5S59VfG29K9
gi5CwDdkw/DAjjDuRcwserBAUrkblqsyJ9aHrTcadced5iRX9Ra2cHs3jBn27Oid
18Wy+hUaUY3vcco87eA1rap/WauoAujpcSv8mIeAFwGgz097a0AUzDsr8hSkx08A
PqfleAftMbuI+dF59SOaCakX9Ajl+moGN7EY3tzzS+iaREe8NYa6HEKeLBGRPcsa
KlBUlXBvPCO9rO99LBjBh2BlvQThXu5KT1bYHww+jyW4tjtDKpn/ZWKBflpiLLK0
1PCrXnl7xXEzLH0yPYIvUehJHlcyKWULFcdjVv67YBonU/VbkdeviLBV3Ya+6A5T
T3qNPlKkseGlj+VUOTYkfCaQyIr/nfPhecA7xiAxzDTzF6dSe1Fq9TeL1vRYIF31
H1GZqVIWem8YgjvmgD3g4CJLW5KuFM+JNCPP4QvkPRI/tZEIFCZ8USRALkQZM2iQ
RKz/LiIif+8LBQTZTmOy8I+DIIHkGACNxVxZNSrJBNwABn4q8M/eRtNLPm4rkZ8x
xWfjDiqT7D+A6iSEiKbVGY1lGFVAqIgn8VYEJWajf+rXXqkvs3btir+O8aOZ5loX
Vgy+wbzmWSnY6XZETKLsjYQQgLanhPxT5Qr68K+gyhGnqGYQF+yoG4fJCaWAFCHy
sdCIc+7XCTU3QyiTajxXfr8xzUi0wk37ZqKhCZDtZTz6uilB8nMDoEm4MMgMhNgJ
BQSMoLXo/pGNeipxiOUnQZ3qGDSUEVTo0XjHtliuC8K99qVRxkW0DMjr52H9Y7CT
IIF3NgkUFPYiA5alc75mQkLUhGDEO+RU28SFsWcdbbr1oI11gZDsiuEtGsNmb7/v
GO2I43PYAr+RbJ0xZFXtmOoQ8GPzWWdp4AOx4fR5xjQSm6VkdkRufrOgRflwVrc/
HVNJ74LE6hihIQQJmlJxsiFX3C0y13RBaWY3gzR3wZ3z4FUz+DkXD4tkKOW5OnUI
Ond0P5j3pUpQ77j/w2MRJxu5W1mEYfAn5nooj5dU85eRGPcZ2enH+cbrKB1dkD+C
N4KFXrw1eQzhdgpVyvfRtCs0YUEPljcIax25YRMdHLzmsBRB+JPIF536FclVETiG
3DO5XUR6EG3dBwSaKT7uxddyoMJ3S7trXTrXzV4uCTpM/7zGoynpW0CuSzba8CtJ
WhpDezARYgIbqKWCUjN3Tacyz8TzRDfDYW3Nn64lAczPyqaPH3+Lg+hURH7m+Uz0
pdWQSfA7dkkvtTYVr2csx8XTlIixR0Sm95RaqdiTpYctxnYG3T4PvyubkDLSsWJ1
h/x01E+0FJUGICPaYoqAt3Gtu2EMH3hfKyb9bvIBk718zAx7Pvj2ylQe/tucYG8H
2OymM/T5ovyclHXo0QodjJndKmLfaTsdeN2FMq/U3WrhtbPhk4SpBDX6gIpJ5Sr8
usiW9Iv3jSdFwWANn+X8VR2vknEzJIurRg9XdWr/6MEmVBR2GCaRbKw7yBqU8BF0
pqkrUV6VvEjkHRz3WXLuxvn3gCcWIPCV764pq7/XefgmAnASFTpzyMx/MHKXbYyo
DYQWgahMVW+7mf9konG42LFFaFcmVrGvEukFfUX14nsapaWDBk1lz0oS7Uhx8EEK
1Ja5x9A4vAi8BdA40atlbDnueOSbkoleCdW4tsMSU70rpW6T8mQnAtdBRpZpFo5U
JHgAbQqpVMXNBx/KGjnGMi5QluWwPV526TNxerzWRZiI750DcsnkhjrEQaRV7dSb
HHoBjPcMgLuKA4TpgHYEv7C0B1GcRJbOD2WU3bA8GMl0YX8H0sMEsTgNasqyB0VC
oJ8TCSZF0DKDnBz1lO1WVcDNBtx/uyArB4rUclgNW85fDC+ChC4OG2zeD3McA3h/
pvPdVWyK7Vq6aWaYt6gONolOG33QYBCF3hZdiDJ7BnYkV8iKZTOp5Wad884lLf6k
lGgdeVkR72AAkeEtV7T5N/cHF3fUC2v+akJMYjWeE5Ogc0bL8bMDCt+N9/C1d1P5
RCv/o9utFLrVwxMVNSSvVT7rCqMq9CcMlbglPYCASCyHyAsbcEhKy6C1LknL+RwB
j8xslUYgbC7LbAXGE513xUWwGGIwEyhKQdVut6AICOeAiRvjBK3jxt6KvyQ1m0ZB
428xG7QbP1rrOujygbQo6Ce/62Fs+SNqx87zz7vufpJQ3i6BGt5rEVUPyBn0QUJr
rVmRkM56oytiJWM0Zn4Nii7ZIkN4POnmHozvVDoJMH2kIRH0Ts/8NyMo0PV1Ol6k
wXiwJfjXCMRVOIs4bFHMcGFSdkltGzAxElcyewcJKXAR3zAhWVrIR9F4lEO2KRWi
8Zxtpl1GJjEAsMqXMbn+xDyujYQ98bRlULxuO1+fe5ZXQs6ellpl/0p5MPu1ZsDb
Gmnv4iRv3svDfIQW5DtIFlQbBH7pJ3haWAnWJVTcFVzB2c+9JtfWrqYcff2OPlDF
Sj3kR5y5HC7bcjTiRvTg9l4fFLzPlV7LuGb93DEltfeTYOxGOfnsvzlcfGV65YH+
RvRGnghEG8mFkVVvuW6SvaE0FhmA5c3v6Y6IMTfLQ0osAn31v1n1BkOLf6v1Pr4V
R6OX18w88uLgLxqzS9bWwsIBS/p3YVzCkR1TCX9zK0OoT5uANYUNwaij5Aq5BQ5w
46reZaXqb3QIQ7hJxTdlkmsmr6P9vev9l/AtQ6lDpsUJT3nvb0Jl4hXEre10YEyw
eoZmXrB4qTBybsZ5uCAbe6Kc/BmlVMg5JMntW/9yoWZ1thdAos+NuqrNRvsIZy4N
5TWARYuvEHCdDT55ffm4A0Tekj+fYdSgfPVL3fFOVGWfNdJG6j8EnLDhbaHotH4U
7aPzYWNHPB9cxDgTd/Qtx22cTthNa2DJO4zV9H7EAN1Fi9ImuBUGyJV5JvO08sOV
21i6++a4EmvO2OknvLaocMiDvSSal+Y0bOkozqMI4aosxLnWg3k5Zn7NdDdzxuWc
ypTtoTshYne17xwga/h1ARw2RF3F072rKwH5QXbMHGxBwgZj6/DpeFrphgULajYa
QYqkSPxjui27uIi82CigW0F7113/TbFhtI/T2gOIgtFv+hM4tbx9nGbGjQLexyOM
HzSjVJuq+CjUyYyhVkpEW3kOCXlHQ16eIXtAlbw9iPgPWrTo1bG/0uhqKhfe9HRX
RGbOexJW+F9vZyf7gS3xxlAvrCP0s8eCKCR72RRh9+y3UOv6FKcaGWlxKfrPSCiv
q006pfeBsa2w+VaGnk9+arIwCPvm4III04CQhhDlUxNx3Zpua7wXhuiV1WzsaQpT
fkWimL/e9sAGJsQTZqmhCPNqboE2jDC0aqGPbJYR/VVoyOlZkfB7VJRU4UkgTbMt
l3LrCG9KMHcrA2JGXsQePZvtjpSjRLu0Eg4KYUlz8Zq0O7x8JOlDI5IlBmPv5ycT
w3Wkv+FBjBdKpddqxrIOYJxtNWm6Rb2Z0Rpxytkv9sphReVjxLv2X22fxJ7lpEWT
lWVG+LS1qqwTZ+up67Knq8MhdgGYOI+axZ9w70tO+bKnvqhefv5LpzLoXLfVDx+M
YOXGQj99XiEGcmCSucTnZoUxAi1CEFDPhZrLCN4aa3wRAtGU+EzZFEUGyd1CQW7E
WF/04sC0jCi4aeu5mD/scRe8cuCxmDAg62GinWCZaG5nbgd9FyJGVahwErIM1EYV
S+dmjGbKzkGgVYrtUez+esIGAYkZBJlC/9rUmH9pifhAQM7b1n1S/vW7+vEK390y
nC8dZPrg/8FUpknmC6YaJwp3u8yETKIagt7IKIgrOgrPKovFnJTK61jhT8Of6Ihs
DeNoH1RiXEzeTUStTn08l/bJTJynxLybZhHSJAnT7WTP6eTR/LdOCcJqBIkFyl6Q
ef4kIEHr5/2xrZc6kmT7MjM7Hu0HxYx8nVddiQM3qpfWQYxbF/yoNARahGq7JH9w
8QWCm0JcKywgQ3HQ6/lsWFb6O6XblyWkV8Dx95svXkQ3+6PLlF3w/dvLtLHR6qgV
wEnEhMh3aXBLbiA1kKLYED3oq1HmQ9d0S6viIdb4MYcaEhMrjANshKkZ34VzvA87
STTUsgC9mfNZxLAchFvKdlx6gQGBt/8RfYgpLu0UAMuo8ykrGzmyh0drWtShJ0rn
wk7baebao49AnkQa18eev/M1TqbZr9bK23OiIcsZXGFpw++VJlBJ+lLrh2iF04dq
oGvNEBXgl1CaajD0EfLTFamA+kKGTI0Vt/Tc4D+KglWrA1RhqCxecpdI6xKkU45/
XMfjT7JlMXO+wUMU7sPzLSw5toqIXk812UwQmTFJSPmjgnOI00vN+D6ZgUCwd4xG
GAgxFk/VZdcq87RtKFdzAOko2IvWByNnMyaRSQ16/HHF/iHgjwd7NbA0yYfO/79D
GGOjrPX/fL5qNQqJZnMIf+oOCSUKdieRTYzjxsJTpliDpf4W/EJfjompVJN69SXd
wjietX6Po+C2qkfyn86bJuPQ78VFhXCu5XYmh3zjBmnYzxEMyj7voDl94vuoxbfT
QLS7F//Isl94ClE7ynSwUFqfadO8i5GDPbiHD2JsofjFGYxUWeGXmkxGWjKZpiIs
q83CaFGAVVhRYSfcJAmRgXLXDXru6LDSteH9PA353qxUnuyAc6oyhQ4vZGTw9GdP
rFU3xDUsXem7Y1qufI3agZPuk08RKQgmI0/Yc5xSj6NA8Djeti/yE93diQksWnm5
PRrSU7crR1yEqBFakg6os/EfsnSQzbSlgRONZl9KweveDDw23IMwG8K6UPQHu1eE
Yy9Q1B9KBCFi1kfiQATJCjvjjT9Q4n5fUzIiVIB5wLLwRl/IewyAsFM8vUMXIl1J
8iuClKkcwasN3sEB0kgqZ90FAjW/Y9xJIMc0vOXNC6nvEafvE2nPCG6aVihQzYHg
7d6VX7oqGyB1yywc9xVSS7G2pLfF02I+24bnT5cAk0CBvdIOZeL1HiZ99b2ki9Zr
G1SjOIKb+Gofcsc67N+V7uIzlksaabrPq5n73t/Dxl4IUpbNC5FRs/DKTbftADBK
77RXfwm/PzlBN4O9XPSkUgr3Keoh++ltT2oNthgaG7yhnQM44o+mYeeldY1hV1T3
tJqQnZuhNfaxvxPeDUxfnzpCeWRC5EJroKD8q7tJvtOZtAPDKkzFSU4+3W/x+O4b
cRl3nJ84XThLE24u+1UxZN41tyJgvHcWNVVFVtt0SrZ3ZSzKDtjBRf+B4/NX3cri
p1FTU2FBDzg7ZQvTxGVeJ6HvSuqf2o9LJy0Pj/6Xjm37eFHwMyOBFDGRUb969Qcz
dYi6T8N7Ukv7+5l62o3+HNuEzInSi2WkZJ3UL97hPzj/jLQp33bwWpPXH3sdtBqY
SCdL2e6IVKDCNOX49AP/5qyjOWONlXZ/sM1IAmYyO/TqGAIyudn7RlTHoIDcFORi
qVz54rzRXH+156ZouacCbJgJenIOIckiRKWwDPXVn5kGCgfQTCiwzYG2E5eCkw5B
+Xv70gKEq5HqaiEN017Q7KEa5a9PLrKnlM4fBEKXUYZW0/HrLcVf043LEG39BI9U
CdLMnwOj8NAY7Tby8yDpJOKOk+jGjHfTpNI30gQSNt8v/4GIxOsjCZuv5e7FKFaF
4K5hHSnqzmGbr16GNCCC1VjzgbFsg/c0YlXxN03i7EwMXFTzQXFHpBbp1d7Ow5Zr
8F4SFGAQxQ4weninCkFHBOSgWrHUAOjZxCXsAOG6g0ecGIBspVNFVQyycefSij4C
cGgFE3hN94NPCqUt4FkGSbmfhCnvdt26OnhJNPyloH+N28jfxCONqX3wUCuOSVtJ
yVLFxPv48xWEpMAvQ4hSGF8p3G4tCuXFzhOCNisYawJHr7Uo4mT6Apzo/1GAqhwK
nu6WyvNdKCD9AtGdSPYvKtyWqzBLO2DJcVtn6OyqphwI4mYDuroGf/ZiBsotm6gg
Q55soAoOJXYgsuAH9OEMEdh+3V5MgHSBNWejyQCoMufuo3i7mibk7Ee+uSru6Qxz
aJWtD9TUWHRQph0G/ZsIUfI7GtuUC7EOBFV0+LKIIsOPi6oC1q2PRIMSAakzYWSe
LcsnreXinPzW9mmFmQuE3GsRfeCoVDfhYqI1dP0SjB9K2drTXSy6fvW2wHUm+yU8
geyWtkLaTOlm3BFkiiNkIzBkcwoGUvbfF2gPTl2NOqh0GFYvHlZ+N9kL2iev++X9
fLx3tqnFCcYlojN5Wjs+stvmw6yXF5e4STyOsJyUzoOXdZbZs21GncF8XdySD2KC
M0Vuok6U2A/6zqViqV9NJhEtvLHl+y9W1XIUHlgYtofLl+MBqjO9gT/3pxQ1S46V
R8XbZ286PC8jtKy0C8kDZhISZ2XnXzfxtVTwLBYFilvs3zJ3q3d54aFaTED1e25O
owbUaoNKCvrgF6aJBou1yAEpeB/xpcI9dj5p7PvUgaAijQEKgT2EpfvwO//ns0Xi
HzC4l9rSvHyC9wnlR/vWeIc94TA035suWontHkyGKodPVeIJV9bivAjIjm20Nh+u
/pViZfhsZCKN1+qScCjUvs27nx3hbrv8FprEbcOaJN/TaOUQsio1i6M2ihE8+0Yk
+LtlCPZQnG7WeTRRKWRerOAUIS6kWfZyPKBQRInm99SbSWlfxsFH6V5gyFJl05im
0G98UAV10iFXiZ4eFZGTKL9GTkWZd8tssyJBXb5+9ctFQV+q0QfpSHxvoiJJSj+A
GFgoR/k9sY63CXoLWsmnMTASUrI6sSWGDaRf+7A/AsGbCLx3trUuIElMVAI5JRmG
W36U/DzXb3PZn8ujNdGn+PlP2Gv5DYT9QiP2Sy2qoFrkxbsZ3yaMb2ejIeqeQkrH
bfxWIgsJoa6xVsKWbYpCNo8nIeGhZfixhv1PH4QiMCbJbwfw1Vws32RBxcDRC8pv
mWtK/Gvclwy19o/m82GdCP39gc8EM5xJalxDXRjhZq5UCgDRnpQg4W7v4xgUasRs
GFvBgkPsdar1Wq99UynDYrgQHoeZzU1DjNZCsMKr3ng/kBe4G1zz0SpE9U+ss1po
z7Lk3+Jrw9hoKWcOwtYK0f3QyGGsKO+dlvVJcEo8YY455nubZOynSkCqnVCjK1TJ
B10Tnaq3eRSJXiYGZncLnzLEe/R68A/nfoVDAi1k039U3xo4Iaar/931PuC/NkHa
5ocfH/sqT0c6k5MJFeRMSpH5KsPrUKj2KOWojoe0ruyYxbJWO3RJT4zddHuF6c7+
+Va8uJuXIWVKPov5v8YGSfbROdeB0Mhj6wKutC5KO4vav4dNhrDxrQvubEIXu1g/
GdCEUBWAMNzwk7RnEsWGHFiUcpC8BwTUBV56RKbEpgQwzgvf5JFExjztrL8OgZcH
hHxRkA2YUMMtwwfTIDKXyfw0x1Zw2ZR9siybUVsGCC7j8H+k919KbVaeAdsZoDXr
keqxAvJfkqNjc/uyds3Zx3AT3n3M4Pqa+H7lwt4q03BCOVIkuyTU0HIwc3ybhw1+
9jVwZPp+sH+iFdl3WrCSm5c9iyTB7lSQw+2+8xJaHR77eLIcZq/DmjKdVoNhS531
zhFkHnmXupe0gjgsNmurru3NwKtiI1V3WHkKqXFMX/Kd6WwMMspvpyw6ognZSma2
mD919zXymq/tF4dMahMrwXRDIwPpWV0aQihsMJTFc2dSsT41/WenEMHBrb8qRRUr
vfstwpnjgMFkjULD3lFUR5dXLaVWpAVhbyzPvQe0hmKBXa/R6G8WZZmPZfQ/jW7f
72OvqTx/IzmU3ihPPAblUHzl5swA78qkTmpVKWnAUMjzy9j8cL+lqrd+7p8/7K1W
+zlggQQkhzr4s7dOUMuYFHMu4HU0H1fWWL8hNzzqAJcu8fazbS2zArDcMK+x5NXP
bpRedSK/NZkS5axDU0dE75AXWEVKiLIbVxnn4k0sms+9kuhwIyXPEC1kuZodycyp
JGbR27DjgSKeRO7byEYbTEzFRE/Vrj/D1e/daTl/ApR4xRTS9GiackLxH9QdGSPf
thEZ2/s+zMWbmUaom1LeHdUgpcSRefksJRX10aswT/1UpMf+g9DJRNT/irzl5SeQ
LOdKvuPE1w7nX0h2SRUGY0b+0F0LyaLAQhNp4FqK5Ygg3uXuDVrwdJfxzPU5UB+F
il3qxYFanLwDMuuQ2UwnThI9SUHs8o8s3seJopsi25bXv2ljacPwToe5osy9gzeF
TbBCAMnLqtOtHtEpWnjqZd/n3FmZltPUFYwVuSDM8GsTHGtIslGVNmA+8550SZs/
+7oSSntTnqmGmbn0yDNzHymnhs3VGdWn3nKruwsfWxdyoTgdZ/Z6QSCwMSvZwoBs
LAslu6jWU+iu3lFOKB3VRPLso/neugdk9Qci1ANLf5bxlg1uafPcaKI3mt+pSNYj
k15TlLDQtQfG8sbg4n9AqJgldsGbNW9CD2uzZDRqDCFYvbZsYprndikrD+5iHOH1
bfjlAFB6ztxIKbsLSCQMLG2tdWdTsMCGHMTdWyU9bFnDcF3u/QUrH9RdM/2Lm8IL
dW6zVFDpKsH/e+UMqKd/oKAWe5IGPuAycmkV2+CXOJHKl/fSDxVGx+hpTvZHvQRl
MSiBBa9hNelk+eoh9I8eAvTDKYMgiUTlZezPfmohECi1Fupr+j8wmT45rMVqKqBy
airx8Xfh2xVYyPZ5EAo8E5oOwsvGs+h4ifmJ5iMfsV3ZE0CJ5fIrkzww9qBWV/Sp
njCJYsD08chi8vuOo9+E36uSQy3AMiA8/U648euOPT/IKzcERaLBnnBxpQoxJrpp
ivGSBTPbYFCXUjjCrrpzuqQK6fL6fy7OwK0iiUwicIOODs41GCRMFiuq4wKz9INu
SsX0jFC1rNnY7JYdXJv+U9yspbYlaW230X/CadDR2nAJdVlL1yN9Fz15kMvSMITU
1nDokfqlz1CFPuJn7QZAH/h41kaWfAc5JEvMi0q72DLHWYBtE0qe+6tHZdXh7QVE
8nDhllEFi4O77ZsoJrxQhVUccxrTM1vV6Ztr3TZssBWiYEaDRE0Tup0CJZFu71JL
BkEmuk+8p5EmA/FkXMCwf3I+ZyDHofTOoUlVnJoUss5o9D9DhXEZqjgSAqw1Sfma
KM+MmHXIlcGYG/G1XBPzM8opFVxQby7EbxxCmkYbiN9tJWP9Kz1FpUA31Xn4kFBs
hBYfUGvYcISa3pu4lH7B/tEtA1+ziIFkc54SjD7C7Fr7vDELwajB495PVRYxyQr8
EzJVtZblLgqRG1B+/PX9vz73LU3ksNsh4GSDsu69l7gUs9dhPSaRnBMRbBX7ql7M
0/PpCZ6WuD/hruyioBVprBhAbNnx1CJeIkDwTvL6Ix5Q1F9Lf2DQmu682v613+Rx
/Sfk9I4wdXRYyZJXVQ/3eavyfXRVtDek1WEptg2XwDFKJJ/zuTqOKevDNCQIOA/t
iPktDKU+nMDRv1ge2kKYznzxUAxJ79hbX2Q8R5n75eDqs2vRW04LOnVL1zvUav7G
c41e785yq9jvahAfBypThuEwtaxNmu7ivomu+WkPeuXi2UtCqysJItnhvU678lfx
YCoDGONGtDKB0kClokNlkgiyNeUPjJYVws/T9tQZIJJOgC0tbP+Qs9wUUB4fKvZ4
kmRZb2uQ3OmgEmfNsg+nFIOCikVj/XRMvC3VZGJTRHFS5TSaBn4TdmKwc0Y4XGPm
u3n++Ke9SxF7bbsU7a+RS/2Oc6A0i41HLgen2ho0toOkp6Ng7HqAGQKypu1b+sef
olrckGqltAFv1pWriWnUadJRaKkv7Lq5QI1vUAFc2OLM6644/i7JmVLvZfiAt9/h
FDvjNJOkaW411TG4lpqoFNBeau5XsVD3IWsNSev7yc8jgrq9Dhw/e0AoVKjaf2pU
Txa3x1mgfZUjgtPNCYebRw2LUpJoaVpv0Mg+3gmG6Yaz1zIQPYxTvdXNGO079CSj
UC/WFHjn2pixUk2UOYWoHdXXAz9GzbSD7k/cn/2DPSYY6Sq+xGUmpAwXKDcPAGet
aoCRob3SV9i9UfK4F7LBzjJKqCJboGtgHbaqJ/sFVYKJ7bE1Bf9DRuGFYfs41RoS
Wl+4pxTV2Ou0s6p62WyzslBjQjfpM9Ts730KDlLud+YNOS4+IvtwbIWnPkcsb5jD
2ZjPBv66mVoPZBUJciZaoKVVzA9CuCAj8t3rcPuKlHeWDe1VvXfIWoPh9MDzmJ47
SU/ABOOraFNpUWEYVOUiYVdy9OgH5zvhIGNkr7SMWP2b6MF4pUQoOnsHJ3DP03UV
BgyBP4L/I5+tntZS1w4qp4Qe4U/M6fjJwN22xmLtBTSapxT+MYB/awpN9gJo9+bp
/4REKbODwyVuM6e55qIKdlbDPufA7uSpnwVZ2rNy0zXUGkv8CgcRJ24gtLhDKP2+
gNcB/q8GbuHsvy9vAAV9Sv8yMp1ctGSuAhyY3YMd0mYw4Ijhjh1h5QavdRw5UXzh
eCP2POqDhHjhxILNXcrUqtxLeyHNUk0/E8dMN6k+z3C87Z1JskGJn+ovMcHfr7zX
wy6L/GlD3Jl9XVSQsNTHgm957cLIuY4MVHBvqIQaZHPCtRmj9qUBWyNlvb+Oba5j
H5diQwTXfnUqwSgIz0/X3wrM0Z9TWzTvvk+7N5wX4S97dv6qgwSrsB2Ru6f+GMU5
VuOLoZkAaH1N/y/u6kZr93iG33ooqqXN0hB2MWxbyrdEsaPgvCQ0raNzoryiT55X
zVpFQZdIRJBpbngCzzPWdvAVJf2SZB+VWbG4ryMPu6hoMYwkahKegEsG4Z0MO2RC
JZpRE4zb42dm5EvoUt/N5pg38hILdf0/rRa7EGxxorwDL5t7+f8pxggA2xk8hfNE
0/DMqrCLmhnT8p7FZBmc8Enf1pvkgDvayWm05Lw6h0gYIdU0iJ30R9HgQlPW9Kat
OH/rMO5QJSyYRSUFqVPLnP/QhqvC2KawdNbSICXKq69UzCSVwhpSVSslRdxednuD
8ZUK0CZQYUpdwBpyuXvlSqaA5IvGdlY/qaY/Q55NZqAkHgiWeEIOA+3slSU2B4LT
M4WkiwZZnkvtDbj2G1HmuUJCQVkcKTifP5+fKyCkS6zsHMYTlj7Aavbp2Tcuwa35
KLeeslhLqmSKTSDUs1OCj9bXzZcNB+Juwko1zuBZlkXmlcibxZSVsiK0Je48ugDm
COA+RmTWoGm6x7VtF+BEmxq8DUgpuOrS0BlNgOJfZNQO5QZAk5marvJk5ewb9oRH
m6j+j+JAOE+oIZ2uw7os5F6nmKmcYfbFV/2I4RBb+3XPV3zy1qvG02jdapTwMAPK
u8ANEiWICoatAyRzDA0BOtfS4nKfZtEl3wf2xcW5DScmbPLPAGPRbT/axpt2AauQ
zrDiCNUNmBKeUdudCjYelfltNLUW2iM6DC/jonwT6Wp823CSM2BbAQC/LKBzdkNE
oQNMx9JQ6KltWe8LbeUN8SiqgfbdHY98AVP4+RlDAGkKpu9tk2aKslm3G2xqZ6Oa
YOCHkpH24mfp6Fjhgw/1H4RkjRp7eZ6zYZRQy6OzmWF/KbUh9/Na1vb0GQWnwc7h
tGjbTiodrhjgpQu7oV/O+s9NpDIz5EKZK4LJFwKpHj5oIUjSxaccTEODN/sS5z8Q
ozDy7W7OIwxHCkF/RnC9wcYPkdHbTiTU519+vP7WoveZ6zPqCLYUOu5m/alLLmsb
QScXjbCqAY7fd8xz8CKBRyrsbLqv3wWLKmYo828osvGLFI5PYeMF0zY5kNFBvuOE
9O9RoHa4PIPjJGCcfUX2oAVjgCGCDp66aA6yQJca/tlNHHZbIfOJwtboofp4BHhR
P3duhZDyGH/m+3CwxzuS04/bVBm2E+V3/itEwRFw80yK85i9i1/h6dPhZk9yRiBj
jnsQ7Fe9wM3ceN1SjwsbyU6KlFPN/x/mpK/HG7Slj+nDZwdoTWwMuoDHsOCyYVkY
oBfYNKSXB9AgAvAg1N7ZE+jQmG1zZG365o6vLgkQTpgXWz70fFpQy8wxAt60k5Zg
LZvQEiL5h1t9c/hV7AHKMHG77LshsLAwgR72PbielS3PhIDFqOr8RcNIafMKLqmw
YUGyDTwWg8dnNPpKXcKdZZhaWMzyZmhIEObCoti9NkchmAwfUGqgdy7Z24/CNT2w
FZ2VwBnygDpWmQWYPXK4owCK5501U8BkiOEtzjGaVSgRrHQ8/UP2G/O9ShyJxgKF
13rOXNpVjY+on7TbeAXpmjB2Q9fQhgAvZxsxy25JUqyINLBQ7aafRvjpCvfm+RDf
uff9aICaYRGYIKetcxiQWxB7+U6MGMadEOOMdl7WFypkwugnGcGhpzuhR4B/K0g/
iaEPqdAV/B5r6iY1aw4UwhkNa8dM4XBX+t/8utN9b8qZpTMDv8mxOoI6Fc/wtiUj
hePs4PlV/XhSpgJJFPUZu1vj8NJ9TNC1q/3ZsCiZuQGzsLda6l2/sOa/7aaMvuTB
qeywYmY41dWIixAI1SLYOhknOTnnxZGyVN+WFz7o3Yu+H+TF9+QFiOOhJ3+JAVoI
qsaCEa/ffYGJnhRv+xjFWjOmLrdIXWaQwkNbg9hQde4PXiouRX720eGM6PsG+Gos
8oInAH9KpSqDhwfUItJoRmeLnTLCEGfhdtsLHbL9IyHpFmQxiFxW5xMoZ0ahTjaD
yn5cqERYn4Q1FDqUWMUxti6D6Gp9z2TDB2Z9osSAQN5DmkvyFXKcZeTTx+jgHmiF
hV7L0kO+HWrRcDzFl7H6luy3oAWFwwuIE4aGAzAUEsaUBKxh36bOu+K3nseX8vxC
fQHerChhW2Wn0kivjH6rgbZ8vXkclSIfOst16F/5wGDhrua2ezFwhFYqMw6B1a3n
kY3OQI8LY+yaeBU+ue8oUOi8IF9H2l6xCorGb9mqOcblvMv9eGfNxA21d5e8qf8g
kLjGoLxWsvDR3ch1NiM4m2SJVApiSoJBIrhGTRr+hDINCTofOcEBHL4Y8oORKnjk
co8ja5oBewLGXJK+AR8FBfyP9wNSau75Emzl4b1W4MCg1sWkL/p0fc85184lS1GC
0uZK+OwnQXzoXhquP7arhtuT2+3okD2Ul8LKywCpdpUiNP1+yH9IRCBMC37TCZZY
ve6i0lktO6pNOEFKklIjpwAH6i/IvLnjfsBxvFj83vXttMP/SIc9FsugJFU1o0hz
eVwbVo14LtF/y/1LJo4gy5VPu1mtH+p86hMSybqx6UgAECNC/kIg5UkWmVbRxqYr
JwCg/55Kaf3XUtnV4wd/ARwsg8Qi+PqQX2P5h20tGSieC/J0AVckVd3UEKWmLQLx
DOj2+Eyw0IBdHn1+F9Gcgr/7Ber4Df/hd5LLkbg19mvrV6N9DoVNzyrlJ2LsUYHK
UylZDGqU9oE+T6xlVSCKAblIjNzniBWBGu058jGsuq8dqL4ZQAazswYgLwBzyauh
yx2KGL9UNwgTKkjFFKdXBfecFX0J9A4F+mA4cVKarO6exG+XxBXRB9GZDZ3JnojQ
9Im+DDqdD/y2WgOyZ/0zqgzI3U8PrpX/GqlzB+j/dZtD6EzvqaCm9IGt4laZ2eAY
c/TrGs4Yl9CQIOOe0aNhxejZQmOxhDaaawzE+OCVa25eQ5ZLVEysVAz0oY8msMfU
K7v0J4q7AEYJtyxmR+RJI8CcDAyXHtcIGx+sv47wpcGAxAtCcQZS5Xv4jioW6/zM
od+nTh1mbXak2+sJxoSrkh8l3hEpUDQqMrcUIZ/A+i7vWnkwXHUJp8ponuW6TvhB
axNC36RMnMG/YPxoP2hahnnhPMHeWsdf8D9UMuQSY0vY9E+7e0JmPESZWmYtmUlv
p1AI+TzHfa6aVw9PjmrZm8U124y4Js+tOWnvPTVvx60P9tqd4P/zIZxEXxtLB0zd
6NmfmRF1Z3GQjq9XVjIjlEUMKvDaWQRcejrDiot1xbA7ngR29/nyegh9UPk0e249
o0Ip2+6THse7IwjsRVpYaNVws4VbvEhn9tJKjb4TRJvmsuAhGt1uR9LxzqKcLaln
+rS45HnZARfFYs2mKuwcJCAuU8C3JDqBMCb/Mbkp7BCcAjSb1tvHyfGzr/3ybKqt
iUgYOb/fEkTxgyk+hmklIi+X0ibDFBOxWxtJZEDictI1EoF/y44rXBZZ0LZw/IU8
IrXzoPc/G+619T6xMBh3FfqXqHWWjV/EFyfyM74bQo2wipMT5R1iamB1XCyMl+CX
ciUAUGja1THKPQP+eqRPByRrUzODdFkUICOn0qqImPB6u6W+XwIfigQ5EN/5sh0k
9NBDP0tRujQOGEzSFxphkaaCkEGTpFpYdpxjrVTTnSTkpS6BIPNZ2XqhkVdFgeA5
3yH3d2pIxqHWZuteQ+kDcoEZzh81izhkc9I01OIpBnbf/LUTfmRkmMJ9VPAI6WUl
4Xp7d9KV3hAMCTd7eRVQqrIyUu6gIe3jdok3jDyZmmmYh07S49AaPP5Ph2MRRJCx
oBC9mR3HzniXsWWvu9TKk28yynOotBfpUUExUe8sdY09zWmSzBDUB7TSnzzSZDxh
3wyBm4HpMC3kRSEOi9RuXEi+2jSpauQe+Xpf7HxskfmxfcGi1qwLIEePlo8Z40hJ
Fg83bUTxzWno9zsqGtzx6uGQoHXaqYDE/Y7t5brLKEyC2tP7Exn8fVQbsDh77Jky
bMA7jDUfolwrbC2SVucURznZumOb+BxHzecedfj9Zs0jI0ONZ6a2GuBP3Vfv/swT
DfgHjTRN0Fr6qxJA4lSVfpuf2ZUVwDZy1N7Ooi0tknbK598URM/ERK4I5pvma6/w
pOlcSOcIbgk7nbVczZ/Dsiqmx3+K4GBKfp7Mc8VjBgUkDf2cUAU4nktoekbT6CLL
giTrVJmtNc3mBC5/F3CznX2bIZOmAVP02zmjTIxAfHWKTORxIdzXJVM+/EzlUDaB
p3APmz3zYTp2jSpN6+sbXfmOzWGAyiXh/jVnfm8cW+gu50X23QkLLuE56+x0qwTJ
29JD1gFWzdnehmizkXvo17mhU7IW5pXzD0ly2s03KT2iLUn9+2W2oKVw0Rippeeh
uKiu0HuP8cNYi6TF0yhkWdzKlkWdar9tYP37GiV3bftPNKpk5You2G74f144Hc7t
T/AG/ObsbRJyQf0AJ4v12UE+XyC938Oi6MWLkEuPnMNyU2mMWojDl40JXOpmUsiK
Iulob3nM5XjGRMHLNUjNzekCz0zH959BzR00/qma1FmiikeRpvK0W2kmEWfda8OU
nhj9Req2m6hdnwGyvjua8W4V2EzGqRxv/Kjl2JUPdCAsd+hzzBn3TZI0MTDlw+oy
zJVL+GKgOpvgd8r9I0YcfiK4N807+Ez739PWLSff+bTaiUZ0Fad8Z/S9pFWa2lon
M7UQPgmm4hqkWAcNB1pYm658tMs18fOyW93tO6MGo8ibddljomvWhrxTvBdyTHHT
8ds9D+0gWYj+AGDMf0n+271G4hg4t4cZ57ID/k/8Ezbf0YDYatDHtrcvP+1073E+
jIsMT48HmCLYbvT9n7x3SBpjwHjSOI+/sr+F9Uk0xwyKL7BCWqMsbTf/2kpCcRLF
a/7ThHwPkdimXvjiPyTLrng58J9t5Y0ynlfH3sLYGs9uBbBn9km9+AtsdjWCpQz+
1hwfzFbWjItK97jnzc1G2/SIQdnAySyWIWX+RRH2616cj53PFfO80jKmFvXL2Dzk
3qMIxgtsju3b8Q3G9M6ll08UXytPCmT2l2Wx8BVAR6XSJaGQSenc6GxNCvQeU5he
J/zFcs3r5cKjnkDrf0b1oR1M2QnQAtoy5liDY7gyWI0jPVUUKYtzBUdwyQzwhSWd
yGIlBpi8EYi+76dqua5SpMFQ/zgS62bxLBV0q75nItTEwvbTFlkSmmJzuw9kLdoS
QG3WNzY0uvuImfRW98R+fzLsT8HHp2MXpYfSe9/2x/mkdUcDd0j+B/oUXV70QEdQ
PYELC19Nu0Ihzq5YFxnamiLAdYYq3sFHqiNR2ScexigVAJbtQOzvMxF8Op3fIDS9
SY+Gr2d8+nwuQtPLHRM0s0LOmWR3OKHRLJt9+5HN53zyNkQcMJ5qpGCmnl+bv8/P
I8oV5u9ff0Ab0ImmhxZCglQ222nbR0l2CknPG+0wMERkjx0NcVNd66X1QnPWfeJd
tRvljEguHRYZmc6CtCkocaSYD5kMiLXFv+hvwlV3rDaj6oV5yEi2sI8B3cCLp8e4
UpQGFdQUNsKdNiHutIKee25SLPzfqy0wRu5slaUFDPvIVAbBObgvV7kAj8Milbp4
6FAZd1uLo7JNezsETwdEj8Hjl3e8lXE0SXj3vQ1UCErDHD6+kwdJha93tSwJ7yPT
+UYLYnZiUocJ2NT0MJumx9gXSO08g2+8Or00IxYEE4gkVykUr28gcXjGgXn39pRg
qbLND38qSvXlBMXVTrsEZ8xDC8Prt0l45Z6Om6Ah3JduWi5dRDkz4FEk0qJnIwjS
ppM/FqOyw183plbqxIc7MNHSa2OZTjkLJbHOeydiYQOUCaX6FIdMwuBlsLAAbMpn
ktFK15dM+WP5g6VSux6qqc7VYFwsoQfwnMw6p/GGSyxaT9JaKgEBLX9W/8q9LxfS
FwP0lbjq5xq2iedG9MDyJe6cdYSzbGcxQ/kSSoQpIoD01NE3ZqeNLr2a7e4vzu9N
mLcbeW7XtciMbnTVzU92G2JPar20OHKJwM4Ybtb7yOZsmru8xB2PZZVjs/uNczd1
bwMScogglULGQ6ewYoKqRpAMXq37SUNjVHZEBa8wuL7uQmePcwQbCYaqthKU4/F/
IEnsId5Luy2zBw5gTqEpnhjGTj4WhP0lZe7gvRIkXkD0mKdZiqqO1ySFHQChf/GT
xSzslT1SgNXDp6PKTt0eDEez1w769nXaq6SQgPkEzLm3HpYm6lmyFtJ8B3RDLN9x
o8BzV+3NjffcnTeVD3/cGHnFYfkpFJjzLhzW8AqD5gZOBzb0I/jzHrv7BukkEQ0f
i2dpRY1FytfkUZ1PBBYpcKPQFoijsS5bA0vmFQ52pFhRuZvLnLdLpa1mep0JxLy8
O8GJkm8X+DEmoq6o1deAK3pt0fKaHgC5I3uqc0R0r2uSKlMyGoju25qLUNzNpnLL
N17AYwhOre/Pt+bF34kkBgRyPRmIKQzKP2iemHwT5suP4+ldrWLatHkI8G6sR4XC
p5RKUjhsfKV/u+sr2QQOzwUicv2zKGVxb6MKPFaaWgkN8xx1+eq0yO2y/+S6jkoO
J8n/mY5tbZlkfsr1WMCusFaLn3Ur3/+diAt/rmsAWVp3T3BS5zVOBZ806pS4A5z8
z4+P8lIrOFppcqVTBXsk0aNvQ7ulugbE4a3qtp+FIPi0qp2dn6pcalAEHiniK9u0
5uqfTN6WLXY2HYs5xuDSgDtLfPzupdoYMen8VC0OhqPd2Cwncs/mIJuJ7PF5mYXy
Wu03vMYw+DBQkXqfdq/kd7qoK8Odhu/3WUUycThAlD1JfjRvDoSah9bwvaaGr7AK
uFhAiE8WUQI4TGrxe4JpznWjnm9A1r3nLXeRRKyPG46KtEFs/YzAXH+qGjAkLcEg
/I2/v3S+s5lCkWENWJ608TLebwU9r9/kjQYu3IISzTbQW81bKgr4eOVMf9JmuMaQ
hUObRO5v3dKHGC5I2uxhIQuvNRRz0hDsMlvLiryip4QCNq2uxOmz18FGrKHqA7iR
XwXUCprlHs4qcmhsInv27W4tISXn6hDng2qfVjieC/UvGWBJIse1jkcP/T6nuheg
90UuqDXIN+u4T2EXB+tM81oPaAq8Jf2cMKBeVpsmfzT1AYTBoucyBVcan07y3eCy
J6l+A9p0Y1jL88VyLjS4TwHnIsSts3efjAai3dv9j3ZFsyKd2xV0VRP1oxkFu51Y
vd+ffkOLF3eOQ4Q26IZykmHq+Gm+5UUoBUQmld5HMGbbEwZ7NYg3T0L946aV4AAx
y+mDk3A0AxClU1Yx26mx0pJh27QLFI9Ke4vBBVjE6LhC8peb7uhhp5zc/Le0/Uzi
JhBsceHKBZrjIGgEmKEaLefIpb1aO9mOolXA2xU07H4aIgMupCnogRpnAQ+k/Xm2
0wyygfhYyvpuwE5YbXyosOwk3Ghqf3fLcVlnXY4EYUmBbqZELnXrCdpB1Ekei3vi
XveGgo8OOMUyA+fog380Wn6f9mM/l5sP54sxXv6qQJoT2TFnS38nz0+stln4fHtT
meMRdsjMQJl3eUi6clqYTL8aYO+sBI2eNl/oK+Q75PsS8uPcSaXomm/lo8m4z1bY
jxlw5ZdSbkST2DlvcIM8j6tR9g97dzEeSA8ZWXcpHR4nUDmO8PNz1SElvye8YbIi
fcUl4rFpj3uVjKlqx/pF84DuPO3tOlPxbcYNcbq5I0vDAT2uFsr/GuDmYlwAgkp9
F4qcMYkhY0lsfW0FQimpgBTmdpWs8mffxxldBtnn9x3ZWHPQBKrNhOfM3t+Q9KJS
jAD1Lq2GpqBc7ezigWMUMKcACoByKMItSgHhFt37cXZjQipDb7itVigMKIBBx5ou
2sWUP2ldFB05iyX9mlAavoRMpBXZyhJ/3Ndmz36jlqiHRx949B2TvS8tG8UKvWd5
WZ8MNkoMWHphqiSb1Cg8wQsKjeE9CvxkiEoDeMzPVR3W7F7oq8kaS4BW9WinbYxm
uiuHspPME+M8L4dH2RTnhmv4vSv8T6aiebRJvoZFtCJAhbzNW8ggun4Jt3fhx+xh
I1RElPgcVJwaRrFtujZ5zOOIXzVG3H/7U4PwAv9OeKnBlqK0EEVlfIa2V0wXMyoD
9ERAWojiaMegma7nsa8nSsbUzenQV2Zh1CN6tKOd79TPJ5t3yaVmq5Lrva7NNZ+4
OzuyktZk5MZ3VaFXQ+6jKGznhvLc0ecDtckik7XvlIe3LYn4eSeD5jQDnemVe63e
8zBV/Me0FWm8mtens/3UbVx+3ufFgllDFx+rK3sY6xooSdu6O+0Q8fbMMIo9Ti0m
XAHiHra68Z9kho8SYJ5zGpUqikodvi88C+KAgxi4iP2OrTeGBOw9UJR9YCGdjifU
qfoPvWWcqm9GmD/1M1dbMyr+qwBWEULYjtR3MUcXKsaY9nJnDCvjDop9PEF+A9xe
6XeigAoEij0jmPHq7JhfuKk4NKL/03DT1ShEBjjhtHI6y6OeZuMWqtxYGmIM1Xgm
zk6mSK4gtIUmW17UuqASiUde+ZG2cZlZ3XAtcVLOfGsePzqZPmxMNlTarKxbpwXg
jjNZKnO2sR60vd38vHr3dqlt+MrJNR2IBh4/wxx+uDH0jS+Okihoi4pj/N9UrArT
LW0+K+D8AOHhwoDC5xEa9mA4TnVnjLzFXPORMYLYa4RG1AbO2/6yVYf40PTAg9oc
h2EobFqp8zPIdnP/JoJcuu1H5hahXzPIkT5es5TB8+wB+xHZtu/g6WDaz0lsBfmB
/3oTSdT+sVX6rG586yG1dlexcQ+UQPWWpgwMjDsYHisEQoFJbUJKgrID03nr3zdJ
2Dl6PWMB+PCcBUJp89096UM5gg0kuIIrk61AJq8hPXkjAqi3UzClWqSolMQVne7v
3LMl+/m/tsoPtRenWffKask279m4gNc2fw07TYhS7wJJHtbVwqgfmmZyTI8GhpUb
MtSsxgG2yhEAUF17OGPvy2M/qWIqjD+CgPRgW73c6N36I/ykWa0NVcWtrCoLmzsw
7IpH7r1rw6BlpgDou9xl2dgYPXuU49oONCW67oybC/jEham8yWurNKCqQJN0+8ar
PdRdaVXjuBXMhmxX4NtZ+/zP4WHjRU1vnnLFto25YYkRg25pKrvTe3ayTaSLLlki
ccAbTyWl6jsW7NUFmrb5mpt7nAmK72oWW1lxTEfwkBZg6t9722Q/hmklYi2QuMbL
pxKemZ0JOFs0RfHTOmTrptxNzoPxgh5e7MgNJftTKcSuNFF0StD6sWzrfEAp68or
ao00S31nVO7MVY3KQBm8jYU4zKCK8uQKhpsnU4uo8cgFLXPaB+YWrRXNi/G5juUC
GlGDV4RFgEKjCiYTJ5nq+gf3yUmOdgrB5Q9xz7tT8qc0//vGtNi5a87aGYAGuLgv
ngS1sRj5CJS9CJaKtH3TPVi2iBj8MJvxvLhJ957431ed8CNVEgRW2oI/Q62Dfxoh
boYvshqsLwZfZVABOJ/TjCaI3bh2Z87cH2uLXxxRqwQXKLqWjKdwb/Rf2nN6N92g
n9uJjac3LMuTnh7GqtSCyr27oxsx75TXTeOQYObNGmb7qUMcvAsctE6+xev9ZJjE
BgAHfTQAFcGp/RqZ6fwUrppjqvhW6pxbc+xFhg7stXkecFbvDtcCb9Uj1yL1BJzD
VsM2kzaWhdjxM7DLCX3F7y8hMvS8audysJAH2aWuMtXfnw1YYeCrrAi4r2f0tgJg
JGkXHlvGguFENCzRvGq6paUUVqHhf7BMEEULToOhD/f+hT65J6TJOwlO3FmOMSY6
MADtyxNGVv6Tq9f2C80A42ofYJS4xmzDNYFZYURP2yeOkl2QyH2wkBbufAOIBEh1
uVJYp0pt6i4fQMqZkmh6ruchZXkFDPjYSxK0gL2/rT8c4TpQrkUFIUozV/C/lCja
S1EUUAHIyGR3VBbU9NkOwW33qH6CFkhec3w7BoTeBa0lMOzt8HYMrNDy2hFGweMg
SaJUCVUgi5M6flrbOznasJrvU7bEsHjvkCt1B5FK0rGDM1mqJM9k4FJoQ0L0rA+/
aVBF8SK9pLWx2qKC7wJqmYvzpxEJXpERZlg7mKbKRqydCRP4NaDrOo/MBn9Sqwqo
RA4lMBdX5D6mlLSI/x5KNDk0DoGZJV2P/XTfTKpjxP9GtZiJ0JCYz5n0TxSWZP5k
OXf9gs9SqPtc2aWWynTQEFQNbmX1dFNqz0bOuy8OH6cUrVRoxGoQVaJ7F3XvAheh
TVSSNCEdK+zqCPlJuDhLvLP8EdHNHR3XA1crWKDUuutBKF6LXFFGtWEJox1XW4ix
tKvdQq5vPkxuAfko2O0Wyte0s56TDv21Glkpo63t88IL5DuSb/IqLvm50j6hkTtT
LXrimSmuTVQjJX6s0UJYNp1QhwKbRdchZRyscP5vqZR1VIs8WNak6q+wmpM2psqa
Hv68rg7dWrf31maEEsZR0qsM7wIOwWVv5vNuwrf7MDTcxChoztSPnHsDAAuKBqS+
4Iz8DxS3I61DZyh67P7QXSYc+a6OK7tLdb+lK/oLpzSoV+x2YTOCruTeheJa8H8v
ucIPS9KloRVvZMgEpZpFGDAT6ccBPtLePHNGu4HIHLMeJ9AjsDb6FpkeQ2mY8B+z
C4tIsEfQkYnlyP7o5+8KjyUPLw1bRll7Ln3RJzbFg+ikViiEg05DEzLuNHAheJmN
JAOf5OhrZylYRf3lUpF2MzwlWIyK/pBV5ibH1yrT5pLc8qyIVGF5gSJCcy8+sqPu
0D+AEAQSksUJHtEkNg3zvsxVSOlw6oOtXfPtPnsfjNRE+BARVCKxVBetCBJGQ05k
kxXgG9oxmccT/vjWMmTchFoIlyisstFzqTBRILlpd8Vhm8SQDqUX+8Z1HpbcwJ9X
rcGDy5BAt2VbPD/yTvJF3Gd5PmSZPh6S41rQ+0K2ke+LBpxmZ5jtIjjUu7dnfW+k
IGqsoSAMF7jXhKYl0h+Fi/dAzq8aJrUI/fYFq/Qv9LxMUowvJ8qtRDPvYTzABEyM
QRSgaGylhOmrJCz82XUSPVS1cBvhX8NtXggQFrg1POS9B2Tk3wyL1IAgLj76qsVz
ArvC6WGBj7qOxPVd+FUxuDoUYF4tLAitrWXCBAJK9UHSzF8AfdMTVWpbkzQTYyna
EEzifs6Zbn65Jf2eKCrb6pGDRBloSvoVJ4ldN0rKg1RJMV0IDOhJ051lx+EX44SR
51+oJw9Gmp9AhOaObhPnayKagxNl6hXsWN+t+gXZvn5nVzsB2Gd5cqe6vZbK5t5z
HzoO/IZrTAo/3FS6dLZEhxeEeRS9PKCEz/NPwxvW/7nQlF+xyn9oMLLw9srfSwZE
gpyGEy6hDkka62/1C+5rB5PK1jRJG4E0xTa23SmTzYxM4D3cWyroVGzAu9tr+AAY
Ek74ErRM4mOxKDE3WQmpNDc55olsBUjoySAtQEgtmzrNmExUNm7S1bp0/bnvOVBW
QKAqz9R241Jw+dvYOv67lpRfK3xbObvH4jXZdMFAPQWruNdhm7Xoe9X8OiB3WQa9
vW36YrPUM8NjJdQv5UmlyaGQ7u6SJTkShf4xLe56nOlCgxE9EaLu4DmOWRyAaN9r
HS+rG1Bd+88kvnxj6UbW8xWZr/5Mlc7JBpauALnMPzN3P+Em3xYnLwkovOYVvPIm
3B5hnAjliff4+Q1DWEHlUqVFWnA0WkIihEZf/vqV7PqT28mx96sy4vDwE/DB593G
hj9LnZk5M5Cut0EbjPUUFeWKscipnC/VNRJYb/z9WiQPIyUNq9z3BBfnKFyHehvK
GsyHD0LJzei8L+pOPg7ozC84z2LgIHCVZdN8kMMpr9GEHQLSqDKuN0oo2XpuUmNE
tabKaZU6xekkroOWSy6d9Gd/QevbXrXvZbZZWSPgSn1wsPWY3dgtRNmzf9o3u3KX
NFxUaDRAClS+DV4l6/KYt2/p8V41KSZjoR0moKG0Nm6aqIkORChIwkPpUUai2cDu
P9zeybUSCMu7ToFSZLnU+NAec2tcJAyYrYrH0OdG/G1yY0fLHPrpgdJoClmQG0kA
L3344mlONzViM5Ye8ederPW2MFAyb7jPul4wxHamQof7ZYZBAfqJn15gR/yPbog+
eXnPxFdO4r73ddp3ctPBsi6syIlYA2Tybpy5UBr1xIVx0RE1oLM21NdKKHUVxcR0
FneG29Kq0Tks7BuKX9vFs8ya34GxLyGF0ewTF98HL0P2qt7HhRls17IRJjjk6yf9
jHgTYHFRd3TAEQ/4jAwlx4PWlxRlmVyAq6HdpoJk0klA4xBlI0kvbGlDPLZQaJYD
cEQTQKFwfg9+B9xUXsbLg48wQFlrM91ygk3qtwibG68qp7jJp+znkUBI/JdFkAV8
OWwpvTgw38/nbkLWfwtK03Zh0KRbWGZC2DjHIGs7w14pw6Hif6fKbpmpJaVpnatr
CgBLX0TnVRVhJ6qr0dW6rdK5xz44ydKQHtipgb/hYl7FL8+3hq98hEEvTkd7VBm2
0j/iT6cxju3aTQaFm+HqRhkTn5SAq+yo1GZIkvkTRFXiAn3XeUs2kQ82zXdUpTyB
GTAf76W/fOxv06MSulj/tNQv9TbxHDvv+iYhAyYaU3qt7bLHyXd1It+rGzLPU7Ms
cGBieOBLVmAy//Sw0/H3s9xvfI8Qykbrv2ev27TGOXWSTwk5lWNWULLhg6ebUvEP
UF62/kxNOv7eJN5pT0L0pJEAW0jbKRjzmwLoCRaU8Wjly7MHjWO7tcNFcOlBsr8T
mpIx+R6Mr0Xvuo+kgPKb6SM40UYZWPvRIFCEIfk0Msc+AR5hbQG1Z1W1qP9RO3Zs
uF6shawqWmFdiPvygsvE1sM6blEtM+HIbp9VFYXb0W62TLUEQiMJ7yd4ipKcHheN
ve3s42N6HKbEOpTGc7oYLlTp9+ZnC9ekLZDVfhq9+x02Mebd7SoSQMDlPWCTgtH5
j9ocKykK7jOVNcAlAS/KfcaCYjPOdC6p3qegN0s4wzoq161rE2G/Nes3E8lL36cr
Z2yV75/ZhxCrNv8PIfRSiMCVffbkb/WUyVcnWZsMdRXJRLVsZmfI5qL8aCxousVL
lT9Bnc8p4bzn965sLp8rBMzJ9xGw84r0Yv69379DT3A3Tl8n0FnLINW8uJGgXe1j
zmRCcdr6xKm3T6lqtarMTV7Z0u2za7RFSoYp2TrDAcJN1iWSr4LNCycNCCNTw9QZ
SRD0OzZ/rM2xDiRu6jvx/d/bNnhZwyF6cpFv+1IHxJwyls7glH0lw74Tvbq6WBT+
grnJm2g+hg6Wa4+8tiqP40fCcTuy4G8qRqk6/s173mMnTl92hkjwoW/Bl68hfgv2
LqUpI2s3CjaS8yVyvB0sZ5a4YNB5YO6I/df5jYzqgBWOd1g70OjsiQIZMZGdPJuk
14ub+hW1X645QbtH/4mcEVcIppv8xjMZ0dBPXh14rLCj/u8m8rAz+xmBd1RdqgBe
gHZ23i28Agl1KLQaVS9f1tHy/N7u5jUSZclPVaU2XbDQzJQMEkGbSYbPL3hmCiuC
5WDtRkPjQ/0eCvvXw8u0WuQblClkC30LYDYihjI+R4X+Pb/L1SkQMYTmJLUcivE5
szy/vt9slmQ3sAJmBp2bRafFdZvbQyw1k4RCyVAh8MZ6SD7uHiRXDu5S7t73f8o3
DoqXbaTW0k+7Q1TPuhmU00dr82g17+5mdeYZJcHpVXWQ6ENtMqitn34QqZPiOZZj
D73e3gqliXvTch9rLSpVtZmvgdxXjqwG6rXVh1FEXj8fGj2yCRpDBu/zdJ/cGMrM
1WzG0OA5RXkEg19mQk4amIjsW/jepLHuXud4nq0QWiL6AiXhBIUwleEpebbhB7aw
MFEiklaGlZW/BsPM9SgQnIonznYhMHZHfLXGMrErNB39hz5ypSFwDa7NUK2ulvbD
oa/9x64Evcxyz0pvxE3ABU7Wa4ozl756jxQd14v3N01Dvd9XN4x3B01aUglqjz7U
gDx7sFzyKfKmfFmFOAR1oOufU/mmzjeNyCZqdrrE6Vjp2gxw3ktZmj+a+R9yE+tP
UIe/r0ZbpIxM38UrqCAmI8jC1xg+gYqNYjbnQ44GAyj7IoLdDzWMGpSGgxihqCRL
F6gFQnE6pwSaOVRRh+Dvzf5SSFltNdFZ9pgy6WEfhpZkIcuZSFd/kHgFuqoZAU00
gVrqmzjcPG+NWEn1SEoyYCZMQdQO38DzAYXNWMyQjFNmb/A2ay31HeYE+yA9WTZ/
NWiKLXfrlKj6iccRkqcxXiteQvLuTNKXrn3dSLJjQoDp/azWJkxGRZBFBUAsku6m
EOfU7VmvRfNGAp53fvkjga2TvkHWPmXAwwl8m/aC3MbvOF2lgZ4ThR15/7OUlET7
GPeQVXCHZ9hosEAeY9/NlZJ/zNsNa6Rw4ObBI6OtFK0xgDTbhMuW6zOWW0P/VP+h
7NjOQKJdz0v4yC/x8Zb3WLGVLZ/kWg3dujEeoStvcsRt+dLwNeiuJk/YnMis/Gw8
WxZCd2VipeA9lbQX77gQo6RlpZdFKZlJVBHia7eCh3byi5zzmUeJPfhuVJWLmAae
FGgj3Lu8EmG03O0PZ3N3YPgB6t2uxs5oYGEswZm4mutPWaMOvFlNtwd2hTq168yS
Ltgrojgu3mRubyt9AgN6omyCbE0Z1ci7CAA/0oG2A2PIbBIsNF76OnMiGSuvgwzc
npdqjFP30AQ65eepq3XOIMBOIaXyvxbFWhp0rwdCcAOYJxfzziBG+4UJL6+gYKA8
VSd/s+6M6swY7+bhLR97kWeJQ4rRRZFnxHC+V3/z2SCNtbDhOcZdkl9MgCWU6eW4
20CsFjy8Bvyzkwoa40g4cFoY1Ep1Ruoy1ifHUR71Eo4jv8rAp4g/P7eRarlV/kjd
pGHqWLmXZlBRpb7JM49fVkNNkneohcsEu3a1xMqvc39SarhsJB5imD0CHUS2HWYG
dZHTrn06dQR9hRwHKVVPcWRV2yQ6k7tq7waJW4B84BdU7512gHmMPFdFRUQ4UZAL
YTf845sI8uOwSA8scKbLYTulObi3/SBAYo7QxC7Nxv+jR8mwpWUi0vDpkLPKkpZi
oiLBOiTqefXxDJuaDbFVoQ41mAHahM04RsuZXMcAwhHwWCYsMG1e6f5zUVI5t+qj
ummDkeDsLp+r9foMDSi0YzhRIDFRiUOFxb/D/J0QYgNiklDKUm1UblDq28h+ntNc
0Pz7r2tntwjcSV587LOjj0hmuROv8oWfnUq0VkmNVMtWU7cidYq4As9gWbBcyBKz
BZcJ4xTtH7CRxY/nbBrAOYdFz+IErt7ca3o6nxf1dwcbfeiPNr+KrtC5HmQWRnml
0GAP2o6qLFhQvhxZ0gW5mxu1TZyCcpxf4c8vruFTEa0YTn2zBI6Mm7x8HgTc/vfL
bdA+FxrDCfWgtOB7xqtKJTYDaH4kiZPKe7uuir1rOhtcrKdGyXvoxpkscxDly1E8
G6bELwuqezBk+Dtg1YSkqK4MWg2Ix0HKcU7OdyN5gk+epec1zBmeoGhgOl7O6o29
1weIIX0mtKVPqrunyzdhgZxrl2FFhjUs4DmLPSbSgccGhcYcs7bJVcu3qulYo/fb
J1lhzsTttjnpxFhBuWJmOtbNQSEGK9lJ4uWS8qP9E4lNBQ9gPitWR7Pgm9j+qVEg
aWs+AxhoFJuLudgPeyfaCYAxUJdYHPtWEXHQ0SrQYGPh/fgmPleu7io1Gnxu5Dui
4YJR8GaB2CdpUX2XB1Rxv5OFpYxoyqHeWBho9JGdOZHbsGLbWruwORKu231/Ka0f
B2sBzQumy7gDSxFPAWW7cwz3fyW1YppgbK9HpYXHLUX/OYHCpBQc4gUTJGFhJiG/
yStNyBSCRFnzctsO7ry/GZ+IfIkORReZVlbClRd4E35EeYTCkNSvMGyg0NMQGjTs
fO14Hv423ORORo5OJFBNV4jynfhggRONUxuENcuat2/aDJr0t/KLdWfHHhv4bvrt
LXd3OrRZHynp157fXjbqKgpzcdnZkiq0vE2UJs1EaFk52Zis5b0/oClbnVe15/cK
cbtlrCvf9rK/lJCH6oTwndHtra3yzccj3YCPYPskhioz0cBd1BdtgfxbFdqztlYE
Quc8Ghp3PDCyemBSn0EbA5kfK42FvqFZK1foS/ayTFIAc1v/pquOZ7YOHRfIIDhl
KR5Xpt7l75BN8eox5q/QcNevTsxspmnpcCDWkY9J75c5PCC6a9yV1Q6E/Bk8nnCX
mBVUPZuUViXvvZ48jGrZWbwpGcCTCUyaqhv/zvlSOul8PMpYK+EPQ1vTT2gxZXea
y7ZJicofi0uibE+c5z0L+OP5NzwKxWefJE6K3ZNq/fkhUNKSOLBSDe9W2LK3Cn6x
l2KclJSxreMRtVgFMc4bglYmP3kFQP3kUJg+EJkT1kknWufKOFX2RZyQ8d126ef4
gNqiUjBUIWuvi967rjrielO3yZ9bDu4i10bZoQq/6raC3MZrLoZ235lOfChs8o1w
8oC2Ab/Q1FCYNeF+TU0b6GMk0MM/dIf9JXoDTm6mJhFPtHgeLXK8LE5UEOwYRAqo
9yGD3HoSeeFmE8YaEi2Uki5SbW6djTXmDcYLd8Hqvk1htqhAMwNyBeBWVr5/IxsT
w9lfB7a48tKbn6lvYRq7kNisaHXTIWUeEGHPR7h9NVG7G2GnamWw3NV2hJ1FAfL9
/2w+gNfD9RaPxd3w27/S/IXzQq7gUS87ezRCV3By7kJ4LgFlhNyU8TAteySepepl
aTL3QRE7nHzF5YBtcs6AImPTWWBdhZ9wcUFeDkuKjGFTme6aosbmVjLQZj5JSmdn
pAgMHxnyHXH7spklVkMKimKRuj9OqNXhj394STtVpmLZxbbVGktEWi0ipcJBKDlx
Qfuw4ArIAYqY8CoMn6/eC4zZasPCCHFv0qPVX5koPAK4tLf+2txz/2U9zsbV/BsQ
WmcFqdZgffUaXY6tqODcXJ8F7dLZ2TndmdUD1NxNbVeUgMcL992d8DCdzNdYLZEZ
KVTxbsQ5WQoFa54c0XqBvwudZcLrrSb2acxPjq76tBV7V8FSI7U3uvjAv9H/Aeda
3WSxC2O2TH1KsL6Gu+yoQe9ChG3sE4Ftj+cMNCnzDj4Ww5hwudKy4mnk81No8IA/
+h5EIdk8sCS90JLfZyr0sjU4KMYj4KqwX8bwz8Qo+0GWOhHqFwI8Cof7RKDLEw16
FjZjtjXzakoiEPtdkGnIEA3giWC7vWIYwBESh9hfFrjDlSZmaNPvGi6RWGsymVGS
RsoRBcIrNHpyiXJFporx6PWuSe8H0BdIQj2IBx54Py3ilGr/SsYYTON8Gjwd2NZI
S9w558iZwItxMYFMbqyydfAV3BFUQZEZ61oFuzQkpQ4wb1io0WNhwUI2HuZCtb5O
2IiWTBeMetAReglyJwpLW74324gPfkX0XGM5bQ9pxScl7YQaDuvVbF/eGXMrclK4
FjFtkye0sdoZO+1NV+Lp+okwtMZor/lUyn4OI+jP5OoF9XCvGh3hvM4bCectePoX
6AXbmJaHHcc4LHE1mBlwshEEFVA/8wz8qL6TNEXFHlFutpPWoVd1BCszkkE2rSN/
xVEU98RYUgLmEa8XPJiGTmoXaTxDPnFuRjtbpjfc+CDTZB7vq1UqcURygjCjt6B8
xvutqioiDp2lTGagiB71By53WcjACe4sqmsjKzTMlgk9+QhDzeaybH3P4ugrs7aP
7oyRi6hkQPSio6jOJTN1tSfbN1jA1+y1CdgjRXY4qZ41VqemXSE5FzXa2Q7pD8MO
ujzxSICIjUmMeFGhImNNX53KmYuZ98H+ruqcGUNQG4NLquGE9gwwDyAIVzq8yCFy
pRRu5D5DY415fpCLhZGluFDjqm0jDz5cbwZtlbT1zEKhz6Df61QWmV+FwoCv6Fnb
D6Bvi8zaZAu/cickxzg+ZTgYs8gEt++CQSAb7TZB2A8s7BCUz83l11VgelRrxt4r
Vz8gzI2KWyZT1PsvLGhGLJtJr6cQhE60jteElP+F2Rg/wXOYdhG7Iu/846LXGLdg
LAyKx1ik9T5nF079+QG23PYA5z+v+LbKwB5AE3x0GCdbN6lMA5RGDSS6HjIybwxw
LOGfn17IeZ+tu8LLK9qapaE4w+kNQLG29o39pQlwgDscAahqg96VBl1hPzBzBiHA
R/VGMr9g22+G2lQvzaIIWKbDVSiAFIsU+7yRFtptQKeIaiLMZDlTj3Ye8m1Ima4o
BCalyViMmIHR42ueqkGxV0wggk7C006AO5ZD2OZ+H6PqXq8dGMXnOc7a/ujsQ9+I
RFTuovu+wGZEsuqFp5uTSPIDyyr5Ws0EJ0b6Q4/7hvapBKeXY07ZdKlAgU/07/mJ
ienvuJizpuSaNuPEZrJhzGMx/+iIv2RpzOiwSAdCaC/ObXUIZyj4iT6qJxhqRlYq
ZR7qjjtAXaSfOc5q96Ov24pVDpohtiqXaFPfGMgiqamhagdLEIxBKsbZVcmTqPau
kBm97r1XjHWzEOX9lIihwZmcMjzyMVVIQOtOj979NFU3ZwLC6RH1A8iaGQQ502KJ
p09X0QK6FTYUFTlpH0je87JdWTreKGUUghJQESbpxnJ9+ZCQ+n27SKwR/5e+Smlx
HzWF/oYuhz+l9BgUpI8B8wsp+UMdKLj5rJb2XLY9bchTvMG7+T5e+pQ5TE11/bbV
yvkrTqPmJ8dl9zbVZYchJvilYzGBoJgwXuC6uK9ds+tc1BsDyp5Cv57zaID7w6CO
5d8jUSgXBDXdts3VM0IWgW77hsUzHBojbJ63MCvT8nCtProLRih5ZtK8aHkt7B1m
VVnp7x0A6VC6ZMo9oO23kaTsw/KD0u4Vm6TQIapZHbMVy8OQrTEQo4EGAcjmJ0be
/jU3OChVaIIOksUT/RwKbgAni7wW9Zajy3DTyQmWouqLO3DcjC0XkRyRdpJAJ6Gv
KoveN4mcy4z4Q5nG13/K77Tqa+bKLPeyneNC9IpDDeuBVOGLMqkl+ixtd54Akf3A
jqGTo583JCJ8tL7UfohyjUszKdkM9lRejZ2gHOSlP2u1Yvomgi37wj4yNq29QN1s
vbODcYN4PHYaRocB3y+jhZSPdaq5b/Gcj349BrDkNrW/uD6w78tsygT/7ooDYuNE
k4kvvVj+TIbTuFVG4NFvZTN9DiLl0XqppdOpKq/Y9wLWZ1fRT+bTiLMUYSHJaBhM
kiVRp6scPW8ogkAyQxoGtJocvVyl5sKjBlyUj+BNI+/ZoosYzVofpDr0e6Trodmq
9vcd7n7GrI2QCcsVDta/900nRO3wnE3cPSPP8fGFeJTBY6ytZOepS9zpFhQhko91
g/+JXBK9s4PjMhArQX2aerT6bJUg1tA+zyUgYyrCEG/WAjx8pUH7t+8nA7lZxmfd
y1FnVMweasr3osUe+7nGaOiRW3epdbUSKA0u/LnmSBDVu7qgahk1z+fSLYcxJLat
J7mbSkpgSL1xHIBTzqrzi94g3WYfpKBIAT+4X8eqMfMMINrgEnTUNqh8dWg5EAVU
FGcPBmAFWC3FU5uGmWgjsSfcjJ0VvjpU35zB13yqOXGE6nblNGu/X30sE6mHwUTK
19ORDNOILpPoEhHGzlwaYEKpe8s/6VO7mlFXHQswbncC0fyn6fBLxXHUYiYyqkVl
8fnbcGS1MBeq8tqxwzj5i6UfmANmCAaVM5zvZkRI7xk8sSZhYbyS4z43vDT5k8lk
zCxOrAjsx9a1xbhaSd8pZ9Aota25uO1ZY3f4Pyv+JaRt82bu5HXLvTulvbkHX1Sh
XecArohsDwesOEdI8xz7dPovSJOTYTNfELcklnmLpNu805DlY34QecovRLj+U29h
i3GR2iaFBKNTUcEJ8CJYCWjQSlMDD87o767FGW8n1lqnFMt/IbcWg08w+lt4+oYi
jk8aDB7koF3l6uI1EzB9NfWcE54Ow9KG6UvT9tOKqFJ5r9O/oTo1sdO0cmNZzLyf
92NAumllgp7wzWr7YwF0C5FRZoJbJ+cT+CR1HoCRQ4n4bGPz/8Ct31Q2UvKX//Qh
DNHnIDyVRYPHnzsoAfVcjH4pKjtcDmzEgrlyFZg8+rOo5ZNXodH5eUmElJlBVQoe
z3bhbBBR9qdV3ZJHNbKMZ2Wn97eDddxPH7o/6qUDqAqFSAARXs8+tOcGN4CCjBdd
vAzFgepPdRIdXmtr1qK4Mlr4Gpc0K183tppxLE7klZQ9JkC+rABk+Yy6SR5hJtAw
Ha3iiT5M9g+nw0lmSGH5c7vxyxUvOzzLKlyfIbsOeBsmzN2LJQoXLyDg+ayzlTdy
i2UiaSX+OMN8byn563pWwig7asxxLpTuApTcUMGToxn469evLQzYdbhyepQaCPwC
8Jla5BlpkXMf5L2UKecQprfvmu/ty4O2bHY4URm84PUU+REJk27W4PEwalZlFuVt
gC1DDHKW/nPmvei0S4G21+z3021m72tb3OA/RxWk8yY6+px2vPdlUCy5LT53H+tk
SoGKfazjUJbmF7PVqJNhuVVe3kyZoUSvclwFn94arX270FscsVAUJ9TolH8yGZLh
yo+OuH2Jw/5+HBbb8pWHCtArMpqxcNZ8g9t1EKS1Zn9kQmEtpeTjLaD+vts2mx/O
j8Pcf7uHuXUwlqe4QUKxnYUOPYQ30qaSoPqq74L0aeDl3VqT/Z1ij16JrK3Tp0cY
Uf50YNJhsr3KtaB+/uQe9yy5udM4o2veq7RbvbZQPi9IOn+ud1Jn2CCI2hyR15Pw
RDxsQ8Qxho5J4MUX91aSeyQbIPWfcaofXFDfAZzFlq6faD3aroRV71gqVMRsHNC6
25XeYAb2iITO10WIXRIvR+rpFqiHbDDuBbG5qWDpfAkyvjE9rvgCNl2vlpr0hxjV
rjeTv6mdVEo1YvwrPqOCjC4/WD/Eygz6M6HcRh50F7h3/yMrq/jRw9DNUdadt40D
NIlSfgwH2oi/8nQtgHCpLmyXeEbUnSotmdhaU0R7OMJUblncG3wEHmVK9XcCMRsK
oxpu5A3HIWOks4Mg3yjpQCERuDKvQDVNcFZPfarPoExh7gdqwDX4a7Uj5P+r08IR
WypgWa095GykWMXT5+mROdPhSSxcfFickFsgiIQjlJmy/Myt06yLLBoy5LppnG3u
KMZYiyLl5c0i3Inmwz6HoOgymaiF8bB71AbPdEs+w3W2aNIsbDl8TBsAazbUzzSW
Hn+1q5PxF5j7IGwz3mpYjM78RweQXbphWpJfYbPOPNHAKqZzAXkW7wtYZ9DAsV7M
wBN6I4Hl/Lax/LixRSvobjFTRQ5C675+gV39/bFRepxFg2o0mQqW2bN9KTVpZiEM
ytu74QXIqfgbdgRgHtPnWIKexrD2D0LC8Scywwcgw+2TrTpI6ZZbIW6db1pE1d3M
ZJ3ZGdImz05cAuflddBjTXAxZnZi4LI71vz9T6xT4Z72wSSjO/DnZ+KIJWN+ilt5
53m4dOmHPYOKFvj1WlzyD+FkBZtzpe+Hlf011g+eHe4h06MZwl3vFzAgbodDKz4p
MVrLzXVFG9PSv2on7HdE164aDpiRx0U9CBD8pcG0PX7hB/fc+1V3DXvkv6uSNiHn
3RyHtxy+o2JxlN4URG/nT9+0vwfLOvdSUI3BJeGvj9Jz9h5NrI/or/TKCXgVFnjD
r5H2FxaCBsf1t7iV9vOLEwfPtjFY4AaXTGaEjO3gNBMmbkfdQsb2kFTotnS/z9MR
UYRSDFSc6HxrVyW7Qhj7vl8OaFUCXJwV6Aniyp93v+KdOnRbP83UsKr+hrDl/WT5
Fy9zgIseG6LQMjBuGTAQQRgV09JvewvtFt/4vc0w+tT+UbXQ987qxZsH1ejD0MLj
dq8Bn1d6MGRbQt8j+QJ5Wt8LKU89axA3dQV3jnzryVLXNlXKyFd4iqVpPY40qEhD
aOQ6vWx1WGh5mVQzQqEyB6wvTjV47WHJ1ue9jxx+wvqujnQ+OCkn9aOAppFkz+Qh
XIbIPpGZ+QR6aI9v4Qc2zauDmbhmD6p7MasUDAWbLlytkgU81xtcD0OFCdLetk+E
clGEqjR6xksKIA5wmbz7kgN9CSBHFmQ9AecM514NPfX4v9u7H16JGuS4niIb9FqH
mtMS/2tz98RTzzdJbL03Z26PIGpUrADJrSo89hlMSk9BWHwZHcX8WZhGeyGrDFio
HbDpVQZ6HajkebhvrogzbeYY68JMJvSaG4kogeLoZsvCNPLVRDubcy6j5POApyrq
jr/rD1T/co7DSav6/iBFbmEFWXwOZp+arB2t2G/GGjY2R/ABz5mnRbynH24T1PUA
2+5/VRhlcJjX0CO0c601CQjWbh7+Rw+Lcu8pzKcP4/ThwWPdbNSYFpKWJxHaacUx
kLqLrb7GpxmQC+FvzmgQQneoAziaEWIjZevovo6xcJxW3He7liBGhfcGyn83EGb3
HeK4H+YDsheXuHY6HKhPRggemgNZBcSwfw8f51xeKOfsO7GfDMRv+ykox3fr859Q
nVtpHIj9UuvEZwKFtQh9DA7wWQiL73N7BgturY6MFNhXyw9Kd4Gwiryv1QwSKsyw
30E5wawNtbmo7eYrpvc/0qeWulc0BCroI1Q+/fyU5aFzEnILat/z/1FStLkrQghe
oPc8UGXYwFL8b71Q2l+67aaMVh3SjYSsc/ln+g0LA8cbwjIk8JJPs3xsmanB8b2g
2ypCgEWPLNbH0xQ0A4NDQrwpE7/UPD/cmDJPPf/0N6wThxAkYeJeFGXIB169aIaf
+iL9Dexjre6TYcx/Mq+sj/i1dsEC0PI6F/r5ys87ESlK4xi4/6gewdkMpzobD1rR
UPvlHnzCFH+ZAQPhxiHvcXgiM8EmmOmeHppP89UtYgowaHApFg1NsBIvO+F1IJl5
IuJNhhp9LpgJnA09MPDuZyQv1OoLYHPh1vak3iMcHyMjdOksmxPx/naABa/zXioa
I+y5jKiVmuLfrzAFTsKkTEqqoajNsAAfUzrfm3fe1jgSRYDjTmlIacIA+CPnTSWm
DTn8i29/cTm1+5GCbAD5KvXJAeuOG3yIGvT599SopyeLcGzdPVHDgl947joSn55c
sZu9nJVsOFEK5ejl3rq+Ie5ByAOzUFFd3JiL4nDpt/uQmYDMYZa74P8MMoI/w/Kz
mqJz97oKqeOvyjCvzDuoRdu3W1xMecGue/BOu/fmZNQrpt6wzRwy6rqRqy9kCybO
P2xo9tBjUfB9gvE+Yc4V+XcyqoCqR1skiplzlS/7mkpWNYsSIlIoqzwln24iOLFx
9tLrUIt+AKEtkwpoBOKOJesTZfepkqGjU1VFD2YFSOaLe+LM3EuIqOGYP4MOFLAe
AAR3H/c/fPV8xiTnv/bZhgUcPtZmyhsVxglTDndMhRtJX9WBZJur89VW1vbSM2QB
c5JyLVNzBbgL/RjwHVd72r7gnA6d5SXAgRFhiYfiScTAQT+0E9pwB2RuQzC9h47f
jRVhVHBS+6MgTV+p0b5rsDMi7MtnJdIoud5MWu2rR4TcIkTTA2kRiRoEy3bF8rA/
Y9Lz/EGfqK/p2D97fvsHflCcWJLklFyNrxxQ3mzSeToryqs92gLOXLr682G205M+
AzJHUS8pa0656+iRbWMasvZFtbYtG40hkDJ220JhPPzusZ1Z/Mzo3MWjwS5ShpZA
ul/nzZqs4mumrsrUMejowdVz/kFsKFxfkpqeh1ls8Te0Z/uq7bfgE9DMAOcCw7lw
3WJKUHf7faOauQpP5/nOZcTqKUIn3KmgiloLIIb9OU58De7SnnpCw1kpWqvhiVew
rkWC3UM5YJkO/Pia9tUrydmm1UrXHT/Rr1qokuCbuq/iNyTSl3B1sBcU/MsWixy0
dHXmQgjucqkxYE8UoQ2UBWsOVIaKopit4IgCSdkfcjkfYe18uhL5CvctMgQdkzer
DCj9dd7UI8ph0myBUMKnt5j0m591kJTeRIE5L5nFpEcQNQdwUgjPDMsWeao7lVpV
DH+m520xAh3ynsUT1EB9NTKSBIZaJjzkUtHhXidLNDK1EwyTGMhWzmNSIVSesmAd
5LsiIzZniFS0jsYlVbD+h5jb+ZVVYx8/2QB6Hyrcsu4Z4e7ZGxpaykwZwv4+ioqw
NM1IRg1HfDz0HXzIVFM0x4u/sah3thc1xjch5Y5SxDP7aqaBLDMJGkEUbyYHVoFq
aHjp6agu1sVmsGyR8087/B5MGNvnPJq9ckQZW3c7Zu/T6WxPexeyqSZ2QBZNyKP+
jVlTFJBXHkPw1vzMh1XrvcsnRAV9c9hbsYbZaliVPFCQTaMu8EGdKI+Qz0EUcSvf
gFkq0CC9G5Uz0MNn8m9AwmYXrQFLO2O54mtcuygP37FgcXJoXvAI9wANSlHMqKQ9
uujRJnb7UDlFiZLDLohlNx/isN4ZZinDv13SH7E4g4F+HRhCmjRqkNEYvrobPX+x
CPvjUz54yZP7qUzP5skviXMhEWqN+PydPvUFseWmIxYHlCCFEc09s20A0toinI8k
llBGP19Yvfn9MMcftR8t+SHsaX8WXCUPOj8WeCA8Hm7ilXzlk3FE45Tfu38vMiC3
QJfiCvcmwo1fbiiHxNnzsizpcBAhvT8N1ANY1zoMWT2SpvsFQlNfWUi7qh/YcbuL
Kfo3NkrOZ0A1FJlSSWN2EU1ZPR51GrbY07edIfAKVm5rcnRLQttGbzXkyKjVoH7z
WUL9T4whRj58foGWuqS91jZjTqxOrRn8WIbNNzimyGCJ5d3X2aanB9L9IqRB9HKE
BBCYEcEgiyFdciZRsAuk81EwRyT3TMGc0TH8LJZj76hDec02ek46h/niyjjvktQK
9XMML5AcddjYnH8peIfZaowex9EJEq55jmimEm+WIZ0RBB2a0dlXlQypJ2hQIDfO
8O6HROq9hEGZg+mZlC0cs72OvGIneWJI6p4UGTBMvw/tLKKPtx4WIJ8Vcle19o6w
+LmTVschey88kJZYCQ6mwQNbgxJrxJxqnA+WoJ8rWn7OumFD/X4e5n7tzyAfHZwi
NShTI6diz6s1XW/NDwF3I7FojRFW5vPBiO0WSJLt+goWeDYxWBKglzVCOO4BSXXc
iOLdGPFvnEoTcCBIVTF8QyqE3WbheO84ZcbkmTaIncSkUXe529Fmlb9yI16Efukr
ShlC2A976r8OWP3DpL0+OI1OtsyYmtTPo2AOPVgFnBfIb8i97IWAfdkP8uB6dWYw
sT3wwNZVRALILxtUjqgkD5Or+5o7Ghkv0GWpKrSYgXAOdOJz3T1gOrVva0yxn2FN
3DMUVT0XfwVdyY0z915/KfgI1gFJAdMVKwbedyFtnmvAr4JqfzhpY0q3aMJnNp1v
xyYeFl/FBEfCQBQdi2GXN0e3got0Mf5ECoTArwHBljFOLCmDdTNIx/+KSVlCh/a5
tzgrWktrT4wim/EQHqVi4BU22nmWTREUY708sNu2knSq3F2fTYTzrTEtpRTM1MRw
HoSoLCHKEOvbbH8CewbT/wRiqMU1/yzOpJN2Jvv88qJAcw183Jj6/Kw4TNost2+b
oyLtvDQtTiVQk8g1ldW1p3aYQcO28oUYiybTh+Z0l1fls9mdas8RUOVM8gep3whl
918bekzfC545AkE/OWyfz0jOHP5cL5Sm28KH4ruCX1qUnU810H4JUtgymBO0Ja6b
pYj831MQDZUPoGZI/b+nonrjCMkzDxGomai0mUMH+J7n32WoDYYoTU5xqRW6KYnI
oaP9xF1ZciQHOvBiw76QrPByjWDUA528ud4iDDH+DL+yDTsPM1v1POJ+tdQIixeO
OzyWNUBJPCWWhat8njk/++Ivt6LIm8/CIjJA72ntLEuCQcShfHasOqsr5hQceh7W
WP5/LQyUsynCns8c/jRShsAsfpG+isqn0bdhUw4ExDMuwSq7oa2bdBdbxtYR/NWf
xuFjqABdtd43e7hFM5uHAYz5TpszbzbFHcyiTi+u1K20Jp6qa8K/LFTKMhZBHUb7
6XMLq400fC4Rif9NR14y2N87E9AOO5xYgk+3cEQuHUQ9vHtL39zQ7lEntBcBSLUS
yMT+hE0R3mTS/+Z0ouGpIFTDctvrFzRfX6VRq93lDAeWWNIY2PWSElj+Q7xmahH3
6OZisulGjfNk6EUcoMHJ5ZNLaprtGbG802Dw/wmo2amactRJxB+zp89fohu7aedl
mqXFH6CpSdX4Xm8r/JIyi5QSIjxmCbsm5jhvVZIHZ4ZkO75o7U5+6yHW+bZK59hh
5pWIdgBR8lxF74oydBjm5scSo6xis0rQ2gE30aJsWCfU7PMjCyFMbNGQMZcvo9eA
5Zx+G/9T/vb0Tg+pSn2IMx44GOEgV8cV5FdI9Em+K2jjxBajMpcDawS+lcGnFKtx
htSbgiftbo4ITtDCJLY2BfDGbH8xQbDlhaqdIgDkU2Xc0a607VrZk0/e0KeK6nVn
w2mDULcYs0NpabP40ssiTwixCvwQ3IKfGQDI8wEfVzu9Byzoa7gQJKHDSd/+PqE2
WzKssBOafdoY66C4iwv7d0GINLrv3s/P1m6900c3bEq3Ovk8+8UNCdYsj/35NEqb
aaUZrk0e8I1JX26uf3slc7feXxfWSAiozkwPQAqB+rpLu0nb5I/j53I4SXJd8IUL
rvbGXMhcZiSRJpPULcHyA5J8fpUwhtMbQSVF9cW1HDLvj8BdjF1VkrVpbVwFQyvS
pvNCPZYBahYL3iBmRs55zJARSxbUeYIdIjgJSo0MfXOgbhc6AFD3x3W2Ztw3CRWV
QfQrKDdHXb1CLulA3DZ8291+shWj4jhT5fF9tD8Hm0lbsvIe4W0+AyzVNXxF9Zwc
z6Bf3ufSVHIrooatRn7zmHZp4iilboK/Focb4FodHCt0d4MS6i7mel6w4o4RPIIU
NPF8FDIUv6KiZixYZ8VV70MvQEi/sWTD6EsF5JGIZ0gnouwH9EoBS2qD73bNkeJh
4Dq5ZonAc4cMWQ/+WmoLo89NHUwrJjkGGbI+2F1jvOMXRoALR48kAdbPSxtpUC+N
N8k9ZkxD2B0OPmiHDzVZ0rij3FP24tW4Rh+2MI2Y4ky+IYAvC4e3cN7mZIrEQieJ
OimC/LOnCN7uCPdSlQTJ24nRopjzJRUfeydr9EjO63yUTzDqNqStuIIEcfZJTzbU
kE+KcSCl+oGdCtWWLYO+RgNf2mCUFJEVt6WleCSp6f2UHr/dVhvuiB4lhDIPmo5A
un1vX1LDvIMpx+2lUyjErli/oZUisP6U3CSEOwY9DKN5A2u+sHuEb6TP2tGSvbVt
wEkeliU6NA1KjXfxcyVXoaDOqHIBCZFzVR9GrfGr7ZEhBbx0MjbhK7SAXeH5xlnN
o8XjJIV+fPYBYoLTMawqhnokK1ezJkZajPMc7e7XceuWhG/guY6D+OAEPD1+PB4p
L0Y+AZIhnSpueYY3U2SquF4gy/qHEmKpggeZEVblhUknVSuA+efmk8MspAipbXhW
2QPJ2F4f2Zf0SDgrHlD0BUad4RbkxHGXCs46r5rrAuUZAzg75/x1q/VPyl/n9F6R
KxgTVwUXRK8oVQbd8vxyGu3sG+QcJNk8avMrW1TCYpJKDOvVU0DTIoWB0TYYuSYN
fpIlaNXQJiRa7E6Of8qSfW+D+2KQzfXT+8R3kRrmkc/5Isi2nPfB2ztH5xFA3OYV
uAbgsO6Q24xv1+LRESwMYpyKJ2adEPJ7EOJmbSYLTUAIB/ZX7M/tj5fRb5OLZB/8
QcFQktjhvKYhraUhTLIjLQ+23J0ckd3OrHS97M8m4BOBgiPiUR17hYLLy0IrIia6
EXCTJbkzoFK3BPE+e9+9dqxExcMU7QvZQyp8YwnTQk13+3AbkcMV96vu9wKPKS3H
cNykBbMqR3F+XzOlE5syU1TBKOIaH+Jsj923trttuDw6eKdkA8QBaxwFfYZxM9f4
JQ2qJBNWrsCJQYEqc73Fc8vEzu4kCsnzOybeu1ilWo6qP8xCXJPZ/4zDGiMtpeBd
qYl1Y1omzSXITUZFlziv/piJ2ZXXzRGEocQrcwEIgHBtxOeTqCXcTdZzSr77MUy1
Ebz+RlbnyerE2mvxg/susicm8do7qmN1P32phxr9UUwa5vw+RWfr1x6k8gBLghTN
9EPPIoyNvb5wU2IR5aaijsWAtN+t1alY8LYQTqPlAb+h4Ph3Q8Oa7GfvofR13GVX
wPK1EeDNR6OiYXQSMO0bUI/sDUWM+Vo8A5o1eGaoizXrDNU+LJ0lpSXoIgnZyO0d
mVCJYTKpE4fGLZzesQ6ToZHRm673JFlUAdmQkHd1SwnnPjfLMfaZGVqmoVwYr775
moXnleSMuv+x2vwNhbbgfoIBAFazn6a20jRoWCWfQY2LxPkZqXdBiiTWB1ujYhnl
vu26ttJJHfSTcis4HraMNH28CSkHp+neQ4Rl5VZ3bG3bsPmuDrN34tPnjmhYYfTU
UHP6GXCmqTzQm3fLKkRRvgs1UfBSTX+XfSi5Hg41jQlbUjXYTPnM1PzFJliYxp4/
60st0SwmVcx2itOBd/+1QwTxgpNFSu9vjemnb568XhOqpyK7OwDEeDQJXuk2zaKq
A13hd0evWR4VwhyQcS24KiqX1B8ev2QIia6zYO6B0X+6ihHny0PXqNX8YpFbMu8/
21YaiIspo7B1crRGAniAIfb1CV9vELdzX4uEYp/4fPxHjFFGUmvHPA0Cqiauo2vS
n+7300tUWg6FO3lSc0G7HLJjsIY6nbqEgphJY3Zka5EqMoVzULwMwh+Wo7l02dcj
5NSW5LTX8iYv1pT1KfrDBRICLQsD8CVpO0m0a42YJv/jb6YKNTeMYRF1itia0DK3
/x+6X0GG1krlCTTF2p/37+8saUjOUkMh9HDru11+Jx9sP/gkxwkoMDvKVwpqsFcx
1MFyPAUTeeJo+aS4YKhACypUuQ8yj7CsmO15eJTZYOKLxXtYhthy8sqt+Zx7EImZ
oZodUPDPlKUoIMhv6AZE9Z+CJDfdF0Dpa7NlPOdJgzb6P4F2hxnvKUXkXqTV1B1U
vkXnop9vsWJsT2+/m5iDn/PSAfk+v8nafVo/T3G0g3txOSsacTt4faWmvbWH/k8r
5PTLDshqlQKJqbL6Sfn46LYLzLPNiO3INqcAIducUtD4lJtZ798jG2EhhkiUjgaH
KkrXENa8vH1L+cbmM7L0TrmeBikEOd/wq2nIdx9F979c3uTt0o9VxPtZC748hOlT
2JaI+kvl++a8eooYxhi/897dh+6GBdSAnInxDMXmsLUeXtt1NDrkcM0oHKCNDENZ
gfiTIWjKuoBiiZHfaE/eLmoEoErbUGYRIGRfS1jlUFMWJvIXr/oumnf/LIjvwZTL
kI4+kj6at4Y+JafXA8nTCfkG6A9Kq4cZ2Hl/7fcWSDcOpnWeEn1ejEOYKU0qo4Fp
sGu1KN6/YYJDUknQGD8eN9nxSfmrti78t2r1xl5zbC4cIRmcKwLCBiCFMuadfBld
FrwqBkGG8V5XyDEuPs0cBEzaQyD/aMsA8C3N/Ucn8JyG/cajwE136H0TI6msxxrG
9EjD6uJPEdJv/Y6QFSyaAyBUY8IzwbpgnwJiFodpz7eMV2co6X9VFB6PZztOxVI3
Gc1V96Sb6Tguf608Lwb+dQsl84F/X3xtivEf8iaWIW58rhnPaAf39MA005W+fnVO
HkgDesv+sYkvQP8eHIpWIPJME+IFAsL6RZbK2KMXWrupHRb1HzN54WFlUkERyMUG
nRYtFDhbF2eIrwAfleZZyPI3DGuAHj+VpRWL/AJlj+Mko9nDunkiDJ9TZVSeZjH9
lYxc7jPmKhwrKrd5vN45wnCRy+s7ecpVzdUchhPgt2h5ZkR+SIqo49qhDhVWiluO
+JDrXZs+r5qTeqHIqiweDRoSxZz3PNiKkb4GW3P7tE40KxqFnztUEKGJQ/ZLy8mB
IyV43rLzcAkRNjeAle3qhqEWmk0gOH7EgkuBedRz2k//qhPJrHyn1HOMbnHlG/Hy
GmgP8AX4+TmnHUyf35mPTiM7Fy55BJFopsGhAw+GDjgWxt1jjI3++36dpY83MhnV
zKjKA2TqoZ9pPQ3VtDGjzCfvFbJsSSiSq7xp3QGpvZ9TB+FWnqHc+n0KLwG3bhvq
k12W5nnCQ6i7Tr3cwEr+5b+pjeyKlNF0A+XLD121z6TKgAenzTZWCIhEzPpjfHut
e76vYLPfQgUgEokhLzb0GTCjDBRgj4wKRzUYnXkouJEBy8tsDgQz8fqGvIQq/OXx
ilAjsIrXqcbmGTSebZyT7wBTAj7buEijqg0ezGehBm8qVmyS1QST2/Lpvds5oa2p
uHknxkyvfv96yv2A2tz2DhOOAjLWKhRfXIucRPCfUc3czzTcJ1LoYCWNo6z78voI
KO3E5o7prKWq46MTgmmlwoemqmhhaHB/OTZrMMaGjA5fycpgr8/DCXIZ+5f1u2KL
FOP9++PW2IY6zQH4ZJLea66VezMzBQQSR7R23lnIsEJWTiiMQThyVI8DaLeo56fd
BuMdvfUoJfjabX8KWXnkX/nEmLL4/3WoqJG70lcoB5w3Mv0yiw7b+t0KV6U/dZW9
OI7G1P+dDWIP6/OgaRwLe3yGmBdbzrVltM3/embO+faMeIiP8Doi2oLGznpWAgFg
cQe9zWwzWsKdqoHLb4cu5Aw394BLSf0PYAQh6eLnc0jd49TeEtaFUSJ2HqnyJeWx
lC3XFQLrTSbVkNVoedFvkq3lFQCRm4XxRUxsw+hR4F5KJLZzbOWWQ3b7xE+wJ2cJ
Jag7AuK4XItKlngpb921hURb4Jt6kmOs64dFzm28YAl8XBgWxovQKEnxOh87MM6g
Vq2xJR0ghScHOW0soOPPUMRMQWT8KytCGRkyMvj8QvYyckg56Nx0v+Jr6azi/cOM
8RL0WZpRRK8+pvF4GX3UCda3HAQw5oLOw+DeC5BXXHogMVl3GHacpjnXeQ5rg7+6
VH3X9LLF06TPjfKwPguQoi6SUMxUrV0i2mzhv/R7z3LN7f/NEiETJkbw+VIuhohx
h+J0xrXrqQUToCuSF7TQTJomrH1YJXypcf2/F8q0hoCgr/10Vc8rC7kMm4mzwbmQ
3iEjGBXGkvZ2KpSNQ7P0U7O0kvhMAmgJTnQ0MaD948UhwPZn7NasY6YD1Ebb73cr
VDxIA+6bPEb15DUsJmTeK6Cv6pNDnqoGKtGIX97HEK3Vuje0KHmnLApF5iZvFq5a
ymtYENLb+acGhUjY4GMNGPVST8wq7Wt/Eg3YY6e08cLVITx4R8nw9DnmVgCkDJSg
77dUCRd+cKLG0zXO1OTtwCuGUYDrnlAWTDDPLC62wLkEFCgW1KIFWC6DUq2lD6dD
yZu3hD3LHLya/0AHiE+8nixKDG7bpDU9HY3ylSXuq1LljYCbaYB4Wcxqb13AWDpF
LxpZe/5BmrtChobDguYT+UHhpIL4GI0+4AD7qV9T37FT/N74mX/P6O6wMjhNjT83
qBOT8He2gRnMyDCwZlF8w8Gb8k/mMVdbRX+duP6J4mLAcya5MBX8+7vK0LHIqBIU
224AMbMR6DrQKqwh3VrU+5Zqx+FGcnCd323XFNYiiZWUcZzpvW0lprL88womJOKT
AmHjcrAqKgnK9x0iuXEeWqkUyeaEr7jiOR6YgUSqItbfXPpLbqeoFzcHGZ24SOYa
zvb0RlCm4JwTo4Vtp99LEEq3BgOYUO9eannk2Tr1266ugD9tNUtTEoBHa93biTlE
xy/Aw5TMWIYdI/Euj1pm+Mczub21KmqFKaMr91x1IL572kHK5pAW9fBz5nWQGZlk
6Oq/32g9pPGS5Iih7LkvvWwz8FLEmWPbcT60kHWUXf1EYYbdgeEaXH+1+adlOSff
M2A0PTjPW9I3tPko2Kh7tBOnAIOmdZiU1qfr7qxzyS0hSZ5NXxJPR/If/E6sH5dQ
sIy2Ig5X1HK9q21Z0knZlZdvWJoUI39X63KYOeyXmWWoGVCgM/2TN2wrl8S4Yzom
roScF4n0fc7KXTZ1hmSv98dkgBqDotu6dqaqKdzjouCPqw4Zw/7iJWmsiwyX1VHX
fUO47ETOAwfNR6nIBWCncnB79+AjJgEScrVlgP97QuMjpfXrPNEco3iVJmmtROnr
cdFrSW5F3KrzXBymYdirAa43ZN/1zTy0I7PhmBP0ikNJdEefyvYhrGduHAngUpIY
2oIQlF7Vh83d31tC5pyHL+gjI8/fCYEaJTrqYAMfoUoYlBXz8GfosW+tqu8oD4jD
MWFHLff3cC5TsHH0otcnW2NTBih3LgJ0ANwoab510NjXSvabct6+Cd1CQGxGxIw2
VlQl/7J91olYJGikl49/J10QT3s0iGSDLmVhXYP57IZJsJXlQsOITMw9b8MM1GCJ
EJyopjhmHjGdDed+wyW+qbonIf9CvZ3/MMUdWEc13CcM6Kyf0xpyuKD6CLj/hRkP
kIxoLQVDRfkiN1x12gkRmTBbBouHHyIsAbwbdzrM7KXnI0PWh3LfZ65DfnUKHI3K
unhbcrqYhyj1PumBvIoNnuIf5oDSNvsSpfM2/SVNmT27FMjfAtGrXvbMNEFNaYBV
dtOLFKCbeKBEyOonlx9kf0+MUrDVd84ZaGmMkeHFBZDgbNOfLwKrGJTuP5GFHSEW
Td2I6uyhS6fhtTVg2RSAo87/sBDcjGJ4JJJTfXCiLgGXx3b0qCFBR15QGxQSHCRg
zgNxXYMUOwPQQWKs/b9VcPSv/B+HUtrscNLUm5BHNnMABXdZvm9C2FCCQFxAKkrl
LiK4GMKufmeJwvA7k/rEGrdU4NeYG3Ii3fA33i4dT8zRIdUb7oslenX1qG+aBGsU
dh57lCRBwQ8puF1TxT0AZnLUMTt1k3dGzOFPybjX8vwszaTFSeXKde4TubLjU/aj
qjmlWNvUIVWFoiGjQeWg20Q+uluExhRzQGik2MN2dcPIumDh6n/BwSoxWjlC3AqE
p7XyP36GY9ptnOmG0oQ0tiv/cODDm6S6ocOcEEoJRWQzoC6u3pEaz7WfTTs8uCB1
w3NHBKE7G7B7Pf+p4G4Q8vLYdQW5bXcIuue/u7n2tOGtEOXESl1squa42AW4aFPa
keD9adjEy+RQsBOIt+5TVytgRlCn8x/SnGcB5iw+3y2KoqEHh3FvhMSm4JcU9y2C
+1HY877g+OOYeWbivz9VwgXhrzskagfCQTWRfRMV7BgVCZ9fXNOuxMPlwLdXiqz2
Ioz3Jn3+ZXnQgfyVNxH5bOOVGq4h4pEH/UeSJc2wERkxlnfIXkPrwGFIWbSCQ8jn
YQMbpKGvi/5PY80tRTbjr6dZxpQlNwg0jLYynjuGrNFR+ya9wyCDMa1qtn8srgZu
MXIfle57tW+o4vdJax61emafp+uQW/a/HMPpgt8x55joxOXwnOESEkOSBGfwkhcR
YDhJ8anDziAIvzwmXkHRuhe6t8RMo8VB6ruwHCA1xNqMmaXfR/iEBjA10LkuG7RG
RgLOuMbWpFB5+JjfsOqg0cCasEkkX6W2TKVI/669dgY7JNSKs8WF6DO4djdESgTD
2PENt44Xv4GvDEjpI7UqY8gsJi/f7dbT4T1Vg7MOEsEAptWlAR2RaK+uDjdPqWfX
9/vVmy7K8jLOfb2/sD4csMeWcpfbUrMROoFuMEcFEfjoW3OI17numuzxI/7YI/mZ
r5x3hfS6zPZxB2XFVBFc6qmZWlgp4XTf2U+G8dKZ7XBL+O90UHcwF/gwbTAHOMq7
xIyWSLDg1eFh/yEAbcPpBrFxSHQAeWgXVrC+Bvu3cqSOLdhspzv3i9OQDuKd71Gy
11iEhb0BLR6vggXKQkjZH1kz2j26RZmFf5TLLFzO/204KuUV4mL9q0w+8XHhje9p
wpaezWWrA/CogBvuX2TBkRwXcfKixtqWlS1UZaX7nEbpFz7VZcjLQVHn6fx3ZiAV
2/EmeSKrqLzdmgQT0gUohNuFEOXul/IwxfLLU2GbfEzrTNiOuP/ECAupZuEN36HG
hzsQuALVA8OgK433EXx9/7HgA07mdRvIO3vNiRS6PBIgrmxTRszQPdowU+DdTRui
qo7Naah2ofXEbgkLy1XbE2XaFjYqkgvMyrPtkI9lxgiyjO+p5Ki/qmmE63fH8SNJ
ExIsiyLEszNp02ZfjY+4fQfOJ/WGWjwurlcaxTmW+KxsBqov8PFEhIGVcezKArNJ
J6Ms0zaC7JLfyqO/FXX2wI+H72OKFa53G0ny4ZqGE9ZdOvgVMG0Rbr57F7DZ02IG
EwB8XX4XBPc01ulsPEe3ZXIul7BjShE0srSUqEPBm+jv8NFTvhSLWIljpHHleT8Z
n/yAaRzkxb0enu53zJSJG8wP3ub+isiYTQvNOhRhA+uJp9F9Lx9T8EqhfbVn6bjI
KpTpbi7gUJUDIDvI78xIy4twHT0/PcCVii147YCVykDUkTBQuSbpi7HDK0wrZ0D3
Q82EW0vbhlk/nSCByuCAybVIGh0E4aHL7KAbZbMtflCexfCSbQOlb9v7gVeg4FDS
R1APSLeb9Fe0gIfsGfanPNmSs82TZY6rhJTGCeefTG4cagz1zTKHElfbWiZ2Id4M
flvx8sRfdpKBWvjfwKcposJBRuJVndXw+f52FdYPXJxk1ulZI5zMKFURhJdgN1tx
FxdU8MQpCi30TZk5xwD1Bal9OMANXPar8x4zEIdn842Aaktbd1mvFMXwK6iaq99k
ORKj8Als1l9poIs8XVKAs4GiBDUHcQucsoX9kogo8I1xn+hHwmYbQZPt0Aehw4KT
SvtWNF0O7qPMLUyh/fSHoYajp05OgTh4E2nD5n4il9w/kwXZtDAgb9kEWu53b10L
1RNKoBEHIPnTaOJWVNZsEngmMlMKrRDzXYe+olwWZLfR7ru59g4NkiNwlaDG8Ymy
wNWvvAcg2KyC021wfj48Q/ghH+ujytERlM91SNOwT5X+k8Fukf90/wbOb2AObpAc
B5aYN0hHWqMA6k6v56JZGgeUJ5/dqZYvwrZWDFX/jDq1O0brRswNAdATh2oe85hI
HnpsdyrYaemNEwa2YYqTljxDWO7vuhMnlsQphXHWNoNYD95UkdUpCFStT7a/DMRc
YY8p0FQlWIdP87ocNMXiRxCcIRNOm8V3QA8XMDxTNoMPuZNqh0V+XpVv5SjcP+8O
qpejXmMSGB4VmSkPIZVHOtq86iO5PGqnpDT9o5dzvGfmN3scnQ534KxSgyhqSPMP
jgkarct9Zx+PnseVQg/OjVYAOOj9HWQSKDMPyTKg2cuPfGZwcvj6Zv21kBug8GCh
5obMnMhGTKUaSMhq2Ejkk8CsV7u85lepM8g0FF8AycYyiMub3Z7q4IfqKN3lp00j
UZp3FzjYMsNO7iYMqBtYW351TkGYd77NMFWxfu9u6b+bN7OT7SYOYwpEFiOcb7g6
2IvDHH2cIjE+5X/f6HjB90OYyK5CB5WGC7p0bmSfI90ZXQXZQhBf0VjUxQ2w8fhE
t2YdpltoWv9Bp1bEHwasr3dbRn89+KD9ARJ3YsdBdtey8A8fRg+HQCrCMvNXYIjD
cdxZw4FMM38TufbgPFbS0OapM9S/afpxnQEiFTJwq/yi/mP5ShaHMYgB9VATB1Fw
iCnyqQo+ci/cJrzG0Poj37Rzxzy7xl3SZj6RC7VMFmpFV/qBQ6DWFJD0eejRq1PT
uAeWgAYnz0Nl+OVZdZ1qjzHY3x2TtppXcXgXwyiYEI0GYayEDei+rCMBJYiNoXJn
CiX9q7vWnlqcbj6bpAEYKo/bE/u9d1M/dO5iCts0xWl4YXLwtDu7aNp0odv3e0Lx
8bLhjoLEeAqu0TMEGQqNoIp4HL9a/jhmnVYuvLWVIfDlf3qHVlnske9og4ZzPWZ4
FOjx1+ICI1JyWY9a/w1Yl+3f7tDZrOMA4H1hHaYYe2flRHflCEh3pNwA/UJMefLJ
47fnuJMmCYf/yiv9Yho4yFMcAykHSByO1Plv8uvzFRaBV4jfOsViM5FjLBptVVPu
Ol14g3gzkuy67AndGeuuQfWDa0mci1MdbUI6X2vbMA+Z+SFdmc3rGWi79itbEo4j
bT3OZrGVVOsOYRxR1cYWllAonGm4teyxgLFCVKBFguZPMXVESeRR79Sm0/DxzgD0
/Hq4OggnMlegk5qE2GbmqUDXZf3elVIzwnY8oaNt7JEeQNtj7UuaUQNcp5s2d1E5
rZM/S2o3IG/XVZQoo/bXF6Tt1voe9HdDfHSVf6LpKM9pr5eof3YsV2uNF09M8mPO
bMp5ANIlmThOK+w03jscDFO+lrggo5uMUCeIZcgOK2zNIx3r2soFfMorKP8L1Gw+
Bei42I5Tp0laxbKXJMA2fXTeSaA4nb8zamjecG51oDlVDMPdon68H5EtIzS4fbcv
l5wswgHOvNZ73J0aJmMlhA57bNKZq3FXkOgF5RhzZw2I0ZBGp9f9qFCEQ8GPGa9B
jlqPyAtzzX0yktlhoXzw5FlpKNpsJc9D5w/uwf15kp4vWWXlGDoGsDY+TUVWKwex
E4mTQsbkzmGHSZ6e7h2PmpP/C9c89ZhLHvccX/tmGaLLUQKN/dHJa10Z8BmivjVi
bSfNSKzwx2l4Bi6iSlU85pUwmBlMfS9B2jmXoNez8ZWqyDm+CHBB8Y//IyywtbrV
dsCiFHNo6TDy+ABNdxi05DrDLcbN57tLVSW4wn9VW/UHlnfWNVqTlbpMjVqspxXc
QyVZ+hk+N1aAN+MgIMbzz+BeAD3WKxz4cSW+FqehPqetn0WZPpJ4LuM4mZ7bslC5
RT29d+sHiz79iYAA/UKxWDRhAOq0K89tQeR7M7ypH8fcUol7OqKg26Oncp5PQbdI
uMLJdK3BzsouuE9pE44/IrROWLTTmg1YUPFfuIhqdjhv3i/vaTMO65wWM2ReY1+x
tVE/t+ivja8+DUXIsMVbhNbihYiZMkvIbW6NZsdzmnA+HKsF3+gikfTSL+H4gKZK
nI1XVJg98mEwvngSCQHQOqzloIIywjtCxekyiOq70R1PChgen27maNIrqyDM6y3z
2AlA+VcSnGmtjG0PAlgSYl7l4rt2dAIE2IE6vXA9eGRB51oC49qmS6W2ooR27n3x
gu/h3bo1JVDyfBBmVjFeWd0zPYXD1vJV1QioDAIgJXiDNUyk6RCyIQghIpF1eT9/
NhAqn2ed899RasDKu21HUHpou5oYfRzk4TYBVr3p6Tyy2jr3/9AjkP6/IHGcqpQc
o6TPuxQ9hspLuHsLa1TpZLGjGGk+0+AlIxaxshPzHiLWHTcHy8jO4DqvYTlwSsXi
vYVnQvPk7V2m+lVWc/z51jSnaF67/0uAlwY6eAzfAFDGITMmkhEa1fdSO5DMW5aR
deOtGXL3ZbJbVtBXK0/nkFEI53gU6lbs2cWhA98i/Y9txSs2ZSsvFrWxyokrbDmA
7BiqImVcHnJpvPG/P6ii8F2YWvtAFcwqLH6RXJAEo58S+LH9kaka/qArF+z3s4FW
L2xCmz6bXDdeRugH4BJ60WPAQMDmKAHnTs74JyauKmt4qrqU2uQsEayBT6GGagUZ
czF9WbkW9HDMybvrEPUZhN3pB20KUL3xstC5WjW0vpevYonx6VGCCxaySnFL5edi
eLKSm8Z6rSc2AFl1XjmOf/BcntGtYK77C7Yun5W6Yy7yOU/IwZOXmuAhnxhT9L54
g5AFGe9zuAuel+++Mnw7GlM9Hzli0VAK4JmdcxS7W/wKllhhX9LJGYaIRgWK+0KS
2SKAyQYSbTvc0W9exJ1mRrW4hLwvDxPw1LMmNiDQSAPtzLU49bNcvRGP9FBjycoT
Yyqg1pVFiw+w1DCbXEu1GQ3YZEzeCpnQexwdCZgtk/TglGSWew/aRBOUxR6HpXoI
Apth5dAXwpSCFBzvvaSMmkLB7l2IlP1k6BPdTrBgNdDfE4jQ9/VDZK5Lb7fRNJVQ
Ypwr/71h1e7s79x0rWau6v7O0pBt7Mtd/BxRxlA6QRmi3Bxgy9DxQjTgE2VFfsFH
tJfXVO2dWB5xhlUwO8v504OgdKcaiVb/Ge6g7Ua2Ryl2VWhCVMNyBtD8LSaQdfT8
tGmXQU4jqQDgK/GFQgaVpur8p620UBXW6FQmTx8ZqKwODt1+0gMEKWirFtUek2RF
Ks8MTBrkYoMl1apScwoG7GgmqpeSUZUBM4lrJIY+0Ba1xUx6g3B++/yB68zmGAub
OvHwOTrjXRPxi9bFA5+RmXQLC6gV3MJpc1ZTutdtsGsHkZVqoyq2li10XgZG2QII
Z64XCop1+WTcCX5PpunMGRrn5oeh4CjxBUdj4DBbhKYOL5KxdOIltfeBIvjcRMMK
3phiJNfic0UfXjsXPlwI63zLrEQIJSMWDIberB1omIfWcLRgfsBtBEo0AzvlFVtR
bEoknf3Foq4aEKmacI3TvoKBheBafOIfZ8sExHuFOSSQDxAhAAJ327JWdg2T+Fz2
H45l/rl8C08NTOXuWR0aylEH99vh/744tb7ocEkwV8HP7bnaxl2vUa21Ed34Ss5g
lx7O8H1avJAst5s9gCPM5Gz8ww64bpkbXYDInstUCbIYGxemrIMaGqw0h3o2ywXk
wqGTs7HKTZKIfIZ9qBhBrGxstE56QGcKkkiXQ6VPvmCPgvmNUIUghtprvkqVSuv9
JaxBXb5Wyjhe4YnxUfl+wSBpT7gt2+N3UOdX5/q9e67Evtb7ze+O5YlYkIrFxZ36
j34INAEKX78MmVDPmSo78w7WTsjo+dga6oCVdzcanQbvGfRqlBYY0MKRJxWS48Kj
b7wd7+5IQsJREOmvXsXeuYLGfVl1vG4CKSINus/BjW5e/Pn2Y2ZV3JL/1+T8XcIO
QC3djM46gh11XamRph6hXSFybwiM+ksG37Wrl2d4LK4IP3NYeEll5uSz0DWgLLeo
RwP1K0W1EyQDqYLRF2ZpX8kr5OLWfc+AoBmui6whYAgtuEhPq0V+zXLewEtR/3Ea
yrNUC4/PP+8hfoTz3WlF3cGJXoKZfCaXlEK4idPCR2syLe3UNMxTlz2h8rzvT+ph
QpU6m+tQE3LS3qckgwuIQhNbR3PkmjLN+URNmVC5n3btac7QCN6U1hOS22dBAa5Y
k8L6locafrIpOOA9dC0J1F6ouOkHXWk/zZM3g79Kkv4TGcVtao1rIw22HbHWBGjh
9OehfIq4VkSSXDtndrm/f9Ah3q7XOBrjh6m5HNwZdb+Ix5ZKBb5tW7AiNAsejliL
SQ/sXNDVJhNccW5RUrw+i3KZf2zlTQrLiJUMHYotFPpg8M07heVWZh61IcdQIPv2
BZINGhwQg6m8XKaYYRWP8WYDtyGqh4Tf6mUyONO35l9pVGTcv7CQWoiy8ykPeUhU
rqt/QDzHnjW5WPWMJgjqArUtIiMaOI/1SQwH+fix0IuLnmq0FzcLGjhRH+Pkz8Nt
YicH6bkmyaBFAoNZk8bLNdSIxey6tpAJedPY/m+aN50ocYRoOAOqvsfqmrjbOucr
vntVnS0gBW+P9/hW6ephNDtEK51xYHFdNxlRKvLI3rTjG30jxkJj26Y0cALnPOMS
AbdsmZTt++nUcbdby+AYFrG0hRVZyXHseXgNN37VJJRbp1mMvZU74l29uHnDcEi0
GLG1K4sQp00XuDDpE6VcEA/wmOu4ObcVryBLrPTzecwOJGZv7RqqXkRuO9N2vXrJ
Nagb/d3jJZTFz8vNyFjf5SicBwjSJpbkcoFZBFUXuFgaQ6c7hVfUudJm/gBYRboL
mtlVlMIcDdesef1Hd8MfiwvHtF0nvqRGWGnQyNs9ex8/JXz3as1uuG+e4yWgki6y
eDnLr02bP/Izp3pCcjyvHq4atrbCh/y9ozPO0Rb7p+C6E98iO2ftystlbWMQS7eI
FysYbCvmx3dYSxkXNFOvDcd02N4hfHTSAyARxaIJTOdULrM94BtPW7h/lWLSSpNf
hmjtyY+Hjn+RGcVGVY9AWBVKG4Kp0H8i1NoUMDVUNbigkRR2TkSm1qnnUlITjrAt
e4O9twxr/XY5PdkerB11KVmzkDVmvc0p3OF6nV1qKd+5j0O/cRhgminZBRqpvMLg
nhnYCsLmaX198gZjenVrqh2EX6Zfbqqd25Ix71/5LArSRxocLOpnjXdXh8hmb/z5
KhKGG3AQoRiBaZKJFp8O1RqSIqftYxb+N0Sl/v3VKvDdd2KdvKVTcqE5MfiTQokC
O3zGTqlWr7uFXq+LtBc2TaQNgsPkdCE5ev59leR8SJvWMlLGLH9GPO6mRNZmhCP+
We1XcXXSAh9G7XtMpazy6eAaQTKjo42zboWdAN+apJz//yvBVJjbfQlrhhCgznCq
VJ1MzMKHBeMTlQ7OQOE024lH1jWeAv8J1xdIww4CCvKkHtvK01pPIDQbotYUN/lr
VoNT7lBgvzo3inqlTArP71Nh6u1Ee/CLfOt/NNkZbb/0baCbYX55P8hd4vm0eoCe
4nJuGH23X/yjkWOupZYtfe3V0LzBO4EWXGEmUQmOVO3ULmG6TqMVBLn4zMh4+Fij
hBXOZR7OMc14YM/CbvpnkZQZwwObpkxbMf0aNUXZDEkLfIjXkjrhKJNPNVSpqrRd
OrXPpfdhjOhZqHidMoeDfGQ1OC7LyFueySbHIfbZb1WgS7C10QTvCqxqSilXVj8o
fXQIeNYd5VAAjvJBo1z7TeMKUWYyaj7DO09IgA3F8kOFJV8cg6KxaDpu8aDVXIKi
otmvMF8uD0Q/UgYgeK4uOMlhh57GGvuqcqItx0P+5MEP/3YHwKvuGHOlCptOr3GO
KfHNvMca/EQ994/LuA/E4ZYnJwsIZFRJSXmgbRvjnRLFSDwb1cvs+muSGycjRv2P
3okO4bfdW1np6gYgFG40c71WewtoBGvepPFsRoxONNGvlYMCj2xYoM0FnjRMQHnz
BY0vcPcf+bFJZzJM3B0nm1DajygIzJRAT58XRaIk/7h3+00Ftdb6QeDVmc/ZMl0v
3rzcO7PUdzv+SbHoEMkpwJmgrKPVi04CtOySLIP/8nXFNMCcwZ9E0Pync+bBZ1xl
UHPlgOb75XpXN7XwiImZape8woEhtyuojSJAcYdo1OVu1VodLnmAawv4HUn+uP7O
Ggn5Xu2A2dZLYRnZRUuMl4jwVJxDuzDHZRdS+E30xfuMyoHaf8gNSKzxcQiXadqg
/o8RlO1yWMFzfoeCNdO4/a+phvKTPV6FAnoUXVIyp0FNE2jQLE1AqYGY74LL/Pq0
dXQz7io4CnVmhNaVUSBmLUMH3FGmzdCVxzwSLiuBi0wt8StP6DPl4wZnF4/OEvRE
dpmINiKZ/yB1eIlDDNhrsY+bud5Cz/C/gx8O4ETqJJ7vKOJN6mxjFVvfkTHopq2l
CJHtenFoAEGnkTUC8EllSGs9mjzgLMA7tSqqSBlaUvAZaZ66QQNvMcdtdAdmj0L4
laRiNL9XSCDNdyf52joc7KPaYavGdxS1qY+fhfR4tDBDKInvem6ZCrve/Djg5oPq
t6DTA93mZFVRganBLvX+gGxFOdTuWJpv0ihwVIqyiqIlW1eTDYutS8Sc2NAF4oKa
08KKQhE75ydaZLvENQqrmXDA5oJRaHITswNVw3CEm300m4q4+DRVYUcUSkHziWfh
nbjC3fXFe3tUARpH6TtpG5saxqMIu6FcpkBb+H4maElazIuC1k8Deg6Cu/mfOAqN
1+IigRMsr7/uuAaIF27UKH4Z1DUbUko03kNnSqjRuf9jVEwJOhjiDhxWJWf9LyMC
gzQJTlyKv8Wb1mOButhWOD1g7FdB1SdcueeeZKnOSULVxBYUtgLCn4d5OphnBk4l
3hJnhKPu2Pzxsn/K39Tdg/GgjbX9X0FcQrC/UONmzANSepTVoPMgjxZUBCrOaWrG
fe6Jq3QUrAk9niihDdrn0tEqR9hZCTCOS13yW7RgVtW1KfBY3uoJnBWlcg8m0VyQ
vYTzhphK5/XQoRH0Svhu+FVWODqBnOy4d7MG2sRW+Kuh4e7YAjxJbRu7e1db/y2A
3a/1LVidpyRNFzSglqizUE5yseo+kCuv+Fc0s7V2D42+wcPE7ayvAx4z7trYV5Mj
HoFaZXNyTvJc1PBmI5SIiSw4NdKIcLP77DuJHc0oEK+65aAuC/eCsordaZOoILUD
VZGlwAmlbLOHhfOK9pottTOYfXP2/QTPtzhkMvg+hEkOIlVpcSQ7yH7jD3uKxCYu
0FpxJH+4uqbafr66DOmR3pgI6gp7kame0SYWCFB1eDywH5y3D21UNVYBU9lACVR2
I7tkNWUiQIVp4FDVXHxOyG740PoDSUsnhQQMKkBfQiKcMjowZNJ3gZKjYGc9WbzD
Z7gI6d2g7BJL4wOkHU3YLR2TxEf9AU2DWN1muHffvM1uBqMut2C1SA6Bf3EK8Ozf
ZY/Tb7Ezyzce5kgCJBLtvH+IY5MCs00q5aHgCQMmIUVlbn3euHF0sYIugDhaYUWi
Ba9zEXLZjxs9aG1L7MkO1O/QBxdbYqbUokML29/bVJE2IQB4MRGigvgRFjQAXOtl
II0ZMcD0aisLO9VFX43IEDSMTt6/B1zIagWXvhK9pX1D4UzxuMlONBAM2cnaNBRV
eSxNP4NpnUIHNvzReGWip3Sb+zVc6rXHwJL32uItkxsfWVr8NrduxAfz2xswLxKF
mg0Qy6trplpKqCVsfOyyKjX6eWB8P0CrAnC/Bp4jS9t8nmk3UvTnPNcwQHT17lof
FrDU97c4j6GHkXPDpFz8UIX0titUiwYJQHyLxQCfDGMxgAXSdO2/HhK51bfeRsxR
ibe+bfPUy3h+PH8QBpOdnoBpY8qL1rJEK3kGCRj7o1R6FEZEyP76iO2iCkSu5Mry
sFqsYdaF7aouWEIDhhr94gLz8pI1nT/8rA+zmocJmI3Zgs+VH0mrJuMXg4dgqwBc
JqybuR2meJffQR85jckmlP4jLLUPmb8kTC3/P35U3aE6/N+nHwfYEZqjaTlyMWQZ
T7yyBFpJKxoHIzcORvz0+3qMGpBI74LqJccVqa3FgFuGuXkyLdNDkG8+pa2RTt5Q
KmieplOYwYLiD+NF7FPXpN59GhOTur9gcsMUSZxglvq6Tv3U2/NfhyThVsAaxI4M
9jG3KnVktbBtos9Dy6PJe2sqWiFYkBardowGM3fgZtM9bleXPILAxFM39oG5+n9a
wWXvyai72Ze0rEEHer86o4XPonJVcUP7hubiF6nhy+z9xXSHphDqcPLwsMlGhWlP
Duk6WKVkFAUwxN1YyZrfMPo207o4BpxXkIe7BI4V4WScikOKO5wlqXBb4GaaERLo
7ETJvyVuOQEJRJ1N+f/vTpQ455g0k/dNacArNExRfBIZCnwCW0jzQdzJW3exKTaB
VtXNWhMGLM/Yo2XbGOOlOSLjCdtwpbuIWoWckFLYy0mnFWFjJVKQpVN8pSTb3ocU
P++HxIehslAUwp1X/sz6mRwI6rxcfBN679yNUrCi38g122f5kdqFI1Qs2lSpOb8f
+pla4AgpnGw9eatgP9RydKy7JOubryQCiAoEyIzus+/NZdWDkHzg3kXkm6mBdd1L
VOh3R7zxsQj7DoGiaaqUIfuuqUKFaoEFXYx75EZRj6L+fk/5SlkKT/72QwzCdkAU
Nc8wEctkkpOWYiq4Pt+eowG+SKjFEpzBLfoYW7oJW3/PsAk7+XEFi7/aoei2UiB7
ul3zXopyMUlZMtcKcAAJohKmUVbotsRV25MG9l/P0D9AovZwndyh4200TAFfT914
XzwySbsrzoJSCZlkr8g/Cxi9Ovsd5MfkGG36bgJ1/SDyuv5vWhTjmp732itVZbIg
CrLXf4w6+rkwgi0dmLyrCCpmbpNZMwAoyoHlxrAucydvsqbC4/AL/cjapGMnxDF7
DWUVZX5w9+pS5F9giPeAlgO6bB30r59xxV9zBxBOb6mNyjUm6Eds73J3RH4H0jCM
uQPEt26Yy79+rrd4yaimrTGp+X6eXKTZ9b8QPhmVDn00vOeATryNzQ/KQYJqQ3nn
WyAysy9WleSP2xwSknICJksdK8D3H8MpwKgOxXvcPBV77C61j8k1TltMDLZYbnuJ
0IkuEQpd7iTKQYbGR3Ig6qPu4HoRHWGt167h3SYqJ1jfLY/+O00xmqUO94/itIvC
jUObXtyjyAIuglGCeScBf3EdVw4yqkUobf29VtcMdy8eeNteh3qe57ZoqYveazxi
N8F3WG4S0HMnnub3dliwea996pnqbCSd3l85kUu9T9gAxsiYwK9ay188bGiaRpKU
dynYRyMk6/GWQdciRN+kkes1svsDkjO75T688IFF214lYZqwAlilm+Sgo0J2bb98
kwVE7cJpH1h1RL7F1IarZF8kPAmVNzMfD/DA259eIin8zG4roQBLqDvvZRdAtcKd
UHi43HrlfCHfm+Db7IAAn1n5tvuQK+f+vzJdFacScUGdVErVaq/mtYJqjCpDPbjF
FZDLeqPAwsXyjCDQ9kGA0EULJTxI4yvToFWne4DOnBVThrQwqzigorfTcYJ60TnQ
ymgr8ay3QZIebUIKH1j7Xmhx6tjvyWi83Bw9UHCGfFEPgvXJjZGqRH7mVO9ZCuPY
E7/O+UruuHyTW5qYRf/CDkwH1r9k1+3QvPHOdROihzt+mAxMcY5VrqTseKJsONvm
iJZvavmXbfvtI5QasUD247Uy/LCDFAPeu7jAKMnMK1hypHQvTa7rGDCFXAV0jROP
NxcULa/YWrrgyUbUaK5BHtO0e9CsgFgsJBvVPHrfVSw57zOsrULXf+VO2qXeJX6k
4rV5d3B5ioNFnIt4Gzp6izVfinF4X+wycsCEZSvoiBV5nNz/sdV39eHQRRDMoOkJ
K9isQ/zqBWJd1ur4glrbO67uafezV8fb4c91NxrjMv3hGWNzn5oY35QL+3gFYh9a
UMBoDfnjWfrKA6QotMgq0L6g2QJf8OddrnNYlb56373lhkEMBLqJ8kWYKOs87QW6
z9q2aqiiee7wtvLc8TH7snFNyJiDPet8uiwtYu5mrTlYWYdDVBIqcxkSb5J7hEv2
SSUmK4DqFxMO6LRrS4XerIBbhH7o1l7scsg45bPB5JYFD06QfpU0zQP9HbV39Q8Z
dguE9LCawg3/bCNOFAXNXuHybWOZHK8N0DXARJmyPcznZJxCqw2ZSPZbmld4YKXz
iPlSlSCstNl/1dshTwwgIXZDxWlgg8kXQN1qMje0qykhDYZm1K2bk86Jb5nvHbT4
TqCOt3eL9iSmRoXLOR8ptYZGySotzsV7fz5WkH9TlBOQB3q8nO8dQTjDO1cqgezL
4vZu7C5kEskQIv5pJ6jvmdnM1oYYZCTx9vU4KtEcgiRLcM7FAkEthjT8sCPaL8uy
RqxMTaQvoZx3qCE0xKltw5Pxwedu7AKFA+pp6/NCZDGIEb8qf+KZL0gN2bm36XWK
exoW7d4wc6GX964oARcTZ0F6PZhtUl0EN1cFnMLieFAw5a8lQd0AHfJ37tAveBUo
XHAhQ9tLUbHhMB45CQprfxtpAp9nGHqTZtCJ0O5MUPSa1TPvJWcvYom9kbIO6a6k
raYp1QdIAXYYYHulGbNb0vaGmtMhT4VKPjvP91RVXX8Olr12RYRq2Zw9eTf5r0W+
0jSbnf6z7iYHn+n1lfy31YsRBmZVpKoWiJRklUiooZX2NX0XtWr06onWMBuSorNo
xZozbgG2BaVVped1FXOSrFlvv9OHLQZbFwtxQz9YpvEfhlfBIszpC3bN6jAa/Kua
+ZFdOPD3k2Wz8NRO7d+bl0UEi8M7/Emvpp5uqg2pKfBK6p7c46khx9keiWuvKQ+P
kDo8CJsVtjzn2s1dVYhDuIk1YzZQNqbskbqZd/wpCHNPEe5co3y6Ev5QtROcnVFh
Iz+K+9J33z1GMkXfc8ebtS51EmhB6zIHoGv0xJZIvK3ot1MnxoCQgngvZHtXrPRp
8zkfihtf7gwHEmvAVezeXUL2E1fDV7uySNMH4MR9WL0FCeo+/Wg2c2xslDxpq6tl
QM/Wsznuq18psTlOxodLflZBNDlhfmwKn2GpZKIOoZ3LE2xGNzejTG7rsMnWlrn0
66qC7GvQC86RH+aLSLeoCyrGvazo7IVJTiuMwmGRZ6m2UzO2GpLysQC2E7TxmcMM
5xvPpAa+VJakN13rzv8fJS1jio8og+5UiaNWRw3b1m9Ky31raY4SvrBXYwDKljKy
zt7vC09O5cKarITAF3/z3Wp1tdVx+C4nRrvNUGgLQAaMLE66GwhigrKBm2tZKgxq
xYWbDe5dNjJriMGsZRLCViT73AUzsSHVCm9ILxFAd4iZuaICew7TJvUrXleJ2Qf6
zuC4sl/wUIFFckeyXfTuCr3Vmf6b/X0u/pC6PPoqrFfcNIk99sJxL4y8gYTL/g1d
9Vu66D7fTPzA6zrz3aK2LqkmBOLenQdgmdbQvnXi/js5DYc9e1OIgHYCGtn23jd1
JStWGrOvlEoli1S8DXk40kqNz2EnSpS6z724KrOZD2g2FqfyE6SJPY3zC/ClB/+Y
fglj6Eqidc/tAnHj/LNZKXE8SVrL4ExvebEjTL8aXyg7bI9BT8WNLUpLITleKF+y
JNoeDAZtyy61eFSDFWfNpKltwjVKZCXNsR6nhZXzOr9NjsRhF8EjbefrSHG5KkaZ
x+jB/1dBKob7QP36raq6vVAHtQCrn1+DGMc9v/7z3rGRpbDuzTJoZir0/qK7HPid
uY/syMDk7NWG7qdMTQ1xieF43b3fXqYTeN5GWV1xsHMKlWsi80hueoYDgldgDx8G
bHBcWFhp3IECm5IQjYoYyS4kOjjz1FDw0YfuksUgFhLRDVFC8ddFG4PTSU0nPHfg
zn8KZI/64P18aW2B2p/h1Q3gEAnAQjC3oKH1A2EH9eM1a4Pxd0ObFlxDpmaONgS7
lWk5RmnyiyEGTkaEs0R/IcVol7j0dKKn1x2yE4qcF7XJWF35EbF726gm+gwWgD5r
hfbChPqglHdlb//CYl0oBBCWe6cS0MAyrd8ED8Xf8CWvTbiWlg4PV/ivhXLO9jwX
ur+48K3DzBMYFrGSzNaNYZyNa9/5rJJT+4nzxaJlmNyqkqPFha6ok91gcVVoAwdX
WX9p5RhQQv4Gq7rCTK0RlCjTV5KNk02CURzeWBSUPOu8xsezm68+DLHWw9cfpiV4
eR1OpHg6vGQTaPonCbnSGilgqXBqbAOwbRF61jEBIOoSOKP34dGmAxxg2wn5puyY
ONitveepPpYxg48/XCvnbbQ2BNzbrCefVBmftmo986pTT/XKUrJRxni97M2xodWm
mk/Zl4uQJyvTVsb8tCIbG9lzfGY9tT1tSDZwHllddtow1ribAOEDN5M24VEjXUK+
EQGqxRHlSJRouNcW1ILZV/P2Hhbqp+9TE+GKUycWpZVW/WdaD9On4IA+On5Xv36I
yDkWqBZwxZcOeOfx/33GZwIKQaPPAW/B8s7h4nppmB7PEqlsgw6vC7oPi1XVoHAL
8NJCz+V3O3tEOzJl/GRRUE/TYEL7N3zBfiYxrd7cQf35eiCUpAN8H6nX4wQEkf7H
ZhzVQUxxQ4QJT5Vs9BUu0LMeXJezlSSjZEDCjqRWYDW6lrxuFQr2aq+LP1F7Plh/
u+Z2Wv0M17i+CwzTGQdtUj4LgUqnhTH7G++1u2tsgRvfwXBS5Z6bAKDoCe5bKRYE
UEeBzSMSaCOHEon8C53T0J6Z2RPt6hS+wBNlAXE/dQavKvWDffPK77tu4VAiQYds
Q7Dl4PnhAWdDlpJHVM2/YEuepsqO2derG7A8Rs+10DH8IRlU7KqVR47i+ds1CtB2
VE2f8Hnl8kjgDGHuwKrH/5n6GKs44dHoMI8yD8z/PDiI8V9ccyrNwC9HBATRcU96
Y3yv42XtrdYHavNGhxXEz0kaLrcifB8tBJjPRYveaGfancs4q/5qGSc3clRbbf0u
KDyEBH/ketzFjXDGbTuCX2+r1dNFl5Deqw1rncoy+sefTKVU5/lsO5pOaE9wKwwa
nqZj2A1ZKNCc27qf0QXOMrse6Zk++DW+mw1bjG1oGrnwCj7DTvx5I5RdGYsQEj47
yNafkQCs1npdHWcx3ghRYks7/P6UJ0Dh8KNaMmTs/5T/e4S3WdtAU3YBFeQV7fY9
JBURUIPPCuUaX11tW5bRxi4N59KrCApBb5jP5l/swIHazK8FxGGL8Rwe1UVUkcXB
LoWnVqlykKIzI43Y0ngZ/h2vrzGWNhIz5q2NZMFCR3d9boAeOPLj4pNhUhmQUzrU
WczkWs/4O+UmnHG1D0gwz3tjeN8rpIVfJAiqMbYkAifYuxPz19au0+IpiXRqdOtR
5xWDYHvK/5ctPnUD+HRG2Zm0mAY3J9YqOH+Z4E4rCkUqqMw9JI0lCcf6ljfrW7UA
RiRCWg3RDgC/OyHjb505fQo4YCGGleNzL0swA2B/sMOSYM0LZ5iCBSsygyf8jTBV
xQa84IgO9z+sH0HEN2ClC4Oa4agJN57wmLAklSTiXFRc35Uv/5a4szilxKnjEqFH
x0F5cyhEiF7WKYUqUeGUFqvUmXPoVbpBpJ/mK/doWx5qxAA+xq/D1W0WOJVaDi0q
MAi+0WzWym8W8KsXERVNSUyOCGb9fhkZ1UGX0PkEF06S/S/H3SPt0qeJhAplkauK
wYUTvU6+2oj4EdEzW3L7JEXItdmjcqr/ieyTwTCoNUThlsl8o+6/dkgJc6Y/AMqM
VjM+nOlgx7Kl1h1pvIPnzSTyJhnPq/Nvl/LbskG9eWz+IM9Hw0BJWdmcRrtIeb4u
H7Dwj+3jj7SYzZA4HUYD1crQxHtInRkGN0otZL292lEozHjfi6vLtz8PEYMmCsQs
xxxOl7YaKa1I96tjhXu0kOQsVQR4ZCQ2laacyjqJDJNE8jquvNMPNTVf6qkvND+H
13LAndOG91LA4TxXLbAs5Lmh17e2L0U29fOoiUiwrn8QMWZGdFK7RwCgWyxib/IP
CthlKdymeHblm5AYl9kHpUIL1kX91BF+ZjxA900cFaHUovfuG584xisKvW0wYIaZ
X84xjoj7C80DnikHdL40s3yAeSOOl6PNUwssElxCKMBCWcG5LwX6Y82K3Td2abT+
g2bnHjWuUZ/TWilxvRU9dKk8tCc0itaYsSCveBYvhttLeU+Ydhs/5Y9OtPxHaSuh
P9NY1N0txi6qIZJUMKaQKtEmxyIx6WvyE1Srocz64/f2ncC7JC9PbJGt4kzzbK5X
bN9lkdxxu+lEQCD+JGlsyiUXk3Zj59JOqj1fB+hC5pG1jTpNjro1lFvuaPY7Rrvm
mEb6RDxZcJnvxnFXJ6wcONo/L5JbR7rh/6urU/EFlWa1HL5VL8+aAT/8WktfOvwn
hFOpdl/Gp3WVpBZuOzziTkFpdoen1IVfzuy7RSnW/WLTXK5A3Y+5EhAUgolBzF++
RgF+jXDKJWr869UTbHAAlRqqy+mNCUcw/hIYaM492ukRwUuTJFFrv+NAv52bRyxU
3QrhU72wZ9tD70CQ0hw685PrWUUTe8vJ49W6TbmkzCoeVyNC8rfbuBFjcSrL4FZn
jigZOkmJQEwsqOeTYv3tRhVPyS9Rvscl3p/lEmI/8P9q05j3dFajKb45rH+F1Qoz
3HG55O+Xh+26ekjHEkqGlZ4p4qdqPczk/tT+ONzHbQL7+jJn83N6yaTPf/R5E6cu
a+6LEModRbS+umdVIqBTCFy2QFfdckgzcjT5MfDyuAgxjK+3tc8Nxh7lP3BUc9C0
iP4ynlLfZWLiWT6Or0FxHIyWT2aR8XtWRm+d1X+lzSXuYdkLxP26r0Z/qyUvXRbx
8JyvTiSiBXeQO45vueMGv0d/6weffXCd6PA4IBmLj0qQZE/7dSRIP+C55JTdT8xx
x5lqKnZxvaKDYbI59XM4jjeGX3/H36txehk/8ZbeAaw3TEprCrVjdcQDslqFsl4p
8nYK7atXppGt9+pXY3gi0bZAj/hMAIieMf3XUZG+hyvu/zZnw7gowIxR+vrkXZD3
jIgjoi4rYzGOnpTObOJlUIUgWvY6sJg3+xCr33utyIXEhMX/22nf8zBDjmY+/X+i
hw6WGFYFn3jvSYCdLLJjOvWN9Qxnp5QH839DxuFXerKOEkPxwqTdtxixhgZUTzcf
rs64TSUGxFSLrl1jKjs9lHWcSCtxT3P5C2XH2EAHzMRTUqo1nIDGiRdWpQ4BUma4
RCJP+bLV+gOK4ZNaqXPcL3NUos3s83vZgCq6VDAhwLtYsD72O16FPvUlQaG6IJbK
dohiVaHXnbyIN2mNHt9JgdS5qPBzapLgnj0AGVtShfEf0Wx2/gROGs609nGoUZNF
JUFOc6aWmfUcXaGaEHsqnnUv9tF3OE8ThlukKmYYy2UXQgJ6vwkC711xHh4znEZs
7FEtFEAogkV7QC5tVG2ZzBzpdbmnDhym69soFaa9LEt68i6cCQUEyH4BZdDuyCth
WhqkKSqOitWiWGextv83RURLEFO29VAFpqMUv0p74k5P22n7Bt8fOSf7txwF/tYU
s4uzi8VwGt98pK6pSl3jcK+T6kMRW8pCSOywK4jDKPBUxAlNNXVZz+x5O4gaWiA8
ohAvCcw+Ilng/LpQv5gK9V6XC706pjSgl7PigdWv061i2n8xYknL32hWPFCuyELk
/36LSIrUHbKFiROHb5bPqA08GsT+LmjGP306T+ehURA6ZGW7nBX+nOCLXebymEHS
DRnSc9oHlz7T79aefnNwIDdXQj2dKy+Oln1LnnN1wodIa7IhBEb1gfnCFDryG20H
QuoY8cgoqnswbZnGymnb4wfo/6kbUJE9OF5eHnitwS5jKISOz0DrEUO9EzsIRKyX
DQeKKsmVsUSx6VHhYuwcVhT6jeSTvvD/5lIaiznFXvjOL63YKaIVI7a7zvfG3NWW
A/DUud1zmf5baGXxamVH6TGK/3yQ+LoKJalb7MtgwZ4cWWt4o3wtjmbr/zzSJcNA
/lhrwmG7lVdhiwFdvbOum6GIntCNi9XHJQ4j9KceLA7h+xB+HWweWj0S4tWP+TcR
8kepSMvt5E64D8ctzWtO/6qLcnS1ulH7yw4wFJ4iy/nxGfNq8bjEGeoA+DF5ZCiH
dCkFmePa4NjYGhNycfKrtXVFdEr4MmWqOCVsbya3ykPPzggxQtOEuE07juVpW+3Z
4/qh4ttkchcEizFmnx6BTQlXdPFzHB49+DQsIvTGqa66qYoR8I/Seq4XEQX+5njn
UypLYgWGJ7VLN6rWeBUctQkR09RXYQDwqX1gcmhphL5JutEGkJLznzTYf0lbBN11
UEecmQI1jZy/rFRbhhJVujsbS8INNAY6jRhw9iA4bXBvigasC/xPWOUD7xpLMyui
YTdZsyweNKIROvhtvBI8jYJ22I+l2W/wIG9kPLupTlrgAgerMkghNLi6CJeMEIiv
NR1ywaS26BgZAPQo2MDcZwwgZl/BTextCwLumAKfyYxjS/9Mdw04HYOSzEU4K7la
RxqQ3vXKRtsr9ACRs9fjyUs/1qhXGZ277tXJevv4oU+lejVYeuaZPwmKfwwFKIsy
Zprn3Uru/HtEg9o79F889gk2cLyeKfDyT7uZiukcoBS5ohWTMzYev02qWuyHfXs/
cMEWJ5UQeGw4XK2pz8ozS1rZC7LrcV7DtDL1KYdI34/MBp8Dza86HY26rclP7wf9
1GbL9ep47m6HtKrqV688TGuMBQJgv5RWzP8vU73Kh6NK1TI7kjAtCDywVsY3SgFC
GusP9qgUS0YvqZYTQMBTJuNKxOesKsrs1hQmibqGBh4EmRrzWdo50nZ4KFSekBbt
PGIaevkPrpNW2dXE3pBwrQz62XZsdQp8+hl1TTxUNYB128k2IHCKLGPNvGftA/UA
xGqk3Xmuiwx3+75lKoGuPYH1O5jAFOxO1Us9x+zMuYDv/E0T0qbrwF636/NBgIOq
dy7QIlvNM197uYIplPdWHv2bA9p2w8jkZqbbnym2JskUNYsayWjFU+yklaaue8de
jy2ivWBUPw+pLPcCmhIePLBVqSWgFTEVdtGi7ZM7CoUSL6fnbuhe0PPYHuvLjDMD
eP12+31ajtHLM66Tw3rWrnqXhFcEyh0+lpjBGyJ8yHibtjaY9GvyoZr/hBnN9tZC
fNvXYSV6o7m8EgYR0HXE+VjR8XPdF1UdvawLVxWlZaazEXKQ23628B6pNh7fUsPi
yYGstAzj5Oaj2Fc8W1GQbGqY0OJMVJDMNs7yXh1R2nyNiA6x3EDrdA65sRzSleco
PA3Ki9+I6TG3dCr2cXlwhgfdq0Ly4LnV2ta3BUJl3VAhUHlmFEGqvke38YrQ2wFU
qdf7HbGdoF/7NmbTRNZn4fe1VpvHFftj9McISunELZXdrs6ZSiCpysV8Nx+EhMt2
OvBpVPqGzIADXqIf1+GwKwVGA7+SstPWv4/HskSwrlJdC0uYuqnOtbymUFPTp7TT
HIaSfqXqm4/XvvrB7ZmSKcagvUTq/KaxzduMelRbYF1wnmV1rb1rZ3LG+xkgvon6
eSbqLZGy3vJzoitaDuOwgJV9du5vbGPe2B1LJIJTMaxiyPgWqMOHVyAYVyYE2ro5
XZtchxkpTB9KhSK0HftU6HRoztR7bV7bgPDU7hLPpR5kiY6bzUGTh8y98JvBYxE1
E23vHgLySXaA5V8OpxcSaGamUXC2Fw895xvpoN7pw9I9/3Ku3wrK6XtWaZdpnweV
uSs8BuFkQ1ZBv95jAmIOqFPjW1Ret/kuwfZ+SDK6lg/UPK5GdV2zSzbvsmddxQIZ
GGB0V3qdzhnBzUjyBEva/Em/DvUJU9YY77Z2eBXi0e5whE7q7FMSVlK+gn+niyni
UHHDwp4a9KPLw44sL3Oq5/pOoYzZCFQ6ZbhoUtC1OfRFDuF/WGwVpYPpOYGemMKh
O+0o7IPEU+cUOUSWEXSXvsXRH1QNUcX6kc6xcyn+ci/uGTodOuh0IEU9ATp/HO0W
qKXx1ubezqn442kXxwQ2P9scW7pbQ36QGharS5zOqOmoSbYBWvog15iJif0JxffY
XVjyn7tDD3r+r4pV6nd9CPtjzAjYEDlFhM3ZiuCNDEEQ2w9FfoLVRRbpNFIDmouZ
na6I+ISIViaa9G0cDhiUiSeMjpc8AIz9TW7tjrz3E6tnvpDc8Owrkw0D78P60TN4
g69rafRppGHibk27dSwji1mEf1QMKJSghauPJnuZnfVnDYUBWwBh+UvugEtnZt+Z
/Dw4e6AU1KdYK/StD8/VHAivCXSvORFx6yGcPJ/Byd5o6u1DU8ekwqcxCrDgoWnb
jYQPKcRF8rp+KGayWknYgH0g5z1CHOYugu0y/r14olgWHezqv2dZvo36G3hJRfE9
nbhnMiUIW8+EDwzPTBEvZ9zec+uCrGLwxdHxm58qnJnUrVX8KBL/DsHRPN6c0cZ4
J0OPNvqUVVts0fbL5uN9BdcPj4exOuVcd7uUDgbBPfEs2SnNExjQO7X+2ip9WVOM
Hjoeizein08uLFqMDegZZ5DD9PdVhuS2QmGxsQrpZzrEYstxjg7Wm7eomgU9k9Hn
1qUSRwCqQfxXWX3kuj8irl6fL2ZKEtSSw3s1KCqylNskZOinqlf57hkfMNjJRwn8
VX7Z1Qm/7Jp2lIdr3Yg7Om/i1o8rvdmexXcbOvRgt4xPuqvtkod5kHxRhzgpU+lF
NIcAUAPiVx2D5XqXxyCx3NwOWkpZLirTXm745Nmx1e2ozLi/QfrNzM0D/DdnSFh+
3OXa9/khl9m6aBLqpd4SnVZosgNPOCjTl2qpAlqeJ+If5ThqmjLMGj6ApdLljhYQ
p1mWsiZzpnstLjdhPylJSZlgECxbW9CHrbir5dGmQVg7zudbMIIPAvcxBIkRxI1y
JP8BA0ZnVewwwljUZYMjVeIkvEM6R/YoRxwtcPBuvOhj1Lslf6fszGz0yRrfX+dJ
kVlA1yU/TKP4PUEAeuj2Y/7j67MrPxxon41D7lFILl03AdSX4ng04seWGo/3833A
egyIs0GgqCS37bF0PSC6rSMYEfYmNFcx8D3ENImH1v9hjiMBl4G9AE9/Xpk+DIfA
HNbFZriWchO97NSB85YZIWHn6jXTy2wExxIiWw7KsUJqFVzypwhPPVJnvlPfNO+u
vhiTH6uCoEahMdRL2ReJKvEXqmzqTHmJgg1o0n34FwC/kxML61rjwfjFx343x8sU
dmeSqEDmNnPX5fj1uXURzqLdaB3AloAbKjJNk7P3LbvqVMDwpFuu+Gc2puRsf3nj
YfRhjND6wtoNUG0CFLK67CluQxljSscPGHDE9fyUk58k8zK8TgV8JrfrL0NH2S3B
4vd00lv1fsuyD9oYzvFAOL4Dvj/nK3+JXgfzGUIYyZ1+dJ9H+L/TcE1K8ytAzSZF
jnCOLc702kmlCKRIhBa6Jg2BOe99h1W4BPbqNWMlv5qrQOk81W78B2qn81m+VWVc
01B0lY14L9bnw+ThCq4RzTegpTKxxtmKfY65QgaAaMujJh9BsQU7UZFgm6YAHOJh
O7RcWg+V96ny1adT7rre7KgxyrCDf2CJFQ4ERz5EIgwJ0VOc7IrpCgbJtR0XnRmL
/14Y2HvZ+SF95sdFP28qx8UImNR7hrLBukVordsx5kVzqcexr/nj8RWGA6bHLj/L
5SgixbapOdjhLXS/8a24aLXu8dYAQWXIvn6Cb36zEm4WgBhbRSUtSBNvvEeTv1xf
vey6qQGwKpZUAqPxH/6mWG42Tr8BtVKuKmBFdxs/PeQZycNoraC0bxPLcdXKNmmG
xeZLsUzwREu7Wi4sfmNBm6VmYGP8NUYr9AjWjY/8xJ0a4ubawRZmHa26ZM8chAPl
ijDV7QUggI8TQJXf0HhSXUdhU7w9K0iTwLQRLea1xjpZUepB/akrzHA5V3ZdYwVB
4bGWLOyAPv9bFbpJ6hO9utCI00TO1bmknNDAhJouyX7jZyFXaX+EZ0XLtUpSHFrb
1hbq5pyFZpNz61YcurgAublrteSEOkA75zv0IDeCX0lmObVI22CkiGMM4Ju7B9zy
M5Ezzj6Fai3iS5yZuD4kcihy8uRfiGIn3MLlo8ROu54nl6x78TKIP1CvrfjLx0gB
4WQp5omIZufvoh+GBf99tUysWWcO5PiNlKUtHGvR3/eCT3gEcbxHIh20xJNikePH
hcATD0zdMaHSe8/XaIfq5wGX1ltAcrkbIIdfYJ+c2tb7pumJFHWeJeTKMmShDnaP
Z7qvz9Ctl9eRN3hBULZQDQLomz4Jmyu+l3Exs9Z5LstfMYMThIpRqU5GPwwtHe27
6u1ZOuV4uQYzOig2f6fCRwsL4Ze+4FXeJWuXGXIGjBkvf1vDiXz1qmYQp+GXLbyY
8skJPUrs/S1YwfpQgO1/xVd5I2ELokfOlimKy7r+gnAQRVy03SfeBmX+j9wB4oag
ggqS8lkzv8TLxaw0ZeMUs2XpPYg9TOemn+w/B39PbirOgQ4ZSRg6Uc16lH3YA/mN
HUAhYJEjN7i6JCT55DuHDKBM4niguCgIKWSBFNYVq7q38HaISSDwa9APN0nWp04N
1EzW37Bfh9SUXIDYRHSKuvgf7MpMviTZ1SiDFn98b05EN9V0PQL7IW9KF/2JXQp0
Dyl8bCnxWbEXxJysHaTzqfrx51kRqDUwt4WmIZEdiWrsXYrCBzAuYx/2n9mGXv6n
QsM+l+gr2dhYaw9XYgUUIN0wllLztglXQonIZsgN/xkNT2y/10n6P1qk6UJKzMwd
HYCZQpgtRmQ9QP+y1y2nilfk3be1C71uJWsKKjd3ysGw8kA3mZuqRZHIwmJ1tfgx
gsopOxmTxtKt81i4Od4n+hW2gi5xOiYB3fcvz2oVNoqRYEMp3FVmTHRVz/YRLYwd
Q7QEQxYfUcpGVf8O63T/FijwtaL7+LGli3tT6BJKTcmD2grQfkffchwXJ2pumeH4
zXXrlKsc9v/4ewoEB3AbOQGsV3exfmSgbE/kvup1wwJy3PuUc67huuaVqYn7kwrB
0YvloarIhfXqhYgxHndDeWp20U9puuSGgcmrUpeKcam998wWfLExntKnKOIVeld2
BIP9En4Y2+n750mnpZ8Gj4ejFmVMztB5FqJ5mkTqavuZb773Q3/JtG4uvn9GunHC
YgNayNvjBY2oqM7Yiy2RlPxbynq5UENPna8FQ+ZeLK231whTbOOpzbJbcarU/fvs
qQ1dUevPusFAm/CSn5+9ryIPK0x6Cklpf+1Cp84VmczE0CnBbTNmZOwHzI+nxGK3
lNVXn3OnW4xekyteIMAzVAjzJD1x8EQkDFi2VKN02aHxLsT0uY53t1vVwq/m/ya5
xOV0xwr0Eqsbl3mZRxMoxEM4KF0yXSsctAzXO8/ZyDN1QIMuNOq+EADPxSgveCR5
bYNgci3nLPvR7UBaGIX0YROtk1htgphGPBxHVVZdPVS4uUVC38bq3juo7lWOeKNl
DVNFSiPRf5Aq5phSihRbFsjAYqGEDzQujCSCDvXEtgTG41MhJs1LEnkzrxxlcSPC
oaeSNtkneVwFFHqabdF9wohUJj9rc0as4HLMP5s8gmwhAoQryc8y7yS6xG768wrr
Rm4XF3sSXixYBECjnoYCO3khbFVjUgKTgKkzJJ4G2ADDNa6aVpylKoKfvL4wBVr8
GKZJDQ2jbS3NIXjfTYo+xm8SSw5a3BNNN3Tsr3/s97PpQE59Ma6G5G10BqNkIXo7
C9rm5Ai2CvwkBklU3EyESlzg0zV0et3pZes4gV9TrX3paC3FBc+BAIf7IiSaDONX
oqAlO0j7xU8qwYnPNB7odejvvN8a46ZFiN/5wxNhAOx2XsBX6JTV1y72aqVcTqp6
ZvKdbp1BOxkUeiZF3C7dai8sXu+1YB4YfdBaI8wOEWtfC1PudHajSWxvgbGCH1e7
6wUXq7Vtmm0125865bCJl0S04s+R2vN3QUgbQgwNlyPZIZVMGQ+SJu5vo+EXjBrT
G4O42V61v9cSI29JV2czaB59Cz1LPZ8IUOg/4BO/G4DTxoq+HUvONw1g+i3PLzy5
P/IHoG/hJp2ai2HcGCM4BHa7oh+chXpcS9vIVfGmF6yMPJu5895oseC0TVsiJX27
gSIG2hacsDmGzW2HRTvRxRsqTyyTvnVnp36SPKcp5xBNwcfav+kOXh2fFXauQNMt
dyCoIxoNQkH8szStdNvsjXSGL59MikAHhS/KEWL7eDYAuJc6FyOaIPqr6OqQGo8X
50AEOJ7/4Z6cYz3PPlvJF5AWiC45GwWi64bjlpFpgWrFLleXDJwjwBw05s74Jjz/
5MT1Rte8Ncyt7NUNkTHo/+K2O02AM6Rj4pCiJpqDFTI53XpBRISgJX6L4YpFbTv3
zTnjiDcY5aUWApr5UHETiBXQIJ/3hkI4ZDO8My9/mgtH7QwKBhDtWDOm18E4yg2g
fZqm/OhZROwrcZuTBU/yayz6lLtvmqM4ne6a5qfBxE5pnzhrjl3XUYeWHkssNumw
f8aM310WCpyazEiV+Wjke0llPhiAWlrt/vYbqXE9Zfwe66LWyMTQZzXG+/x5incL
f764u91WEU2p01ssacCxmpEGNPzF1WhvZSZXR61YxnuacJ6xHcQMntQY2T9Ft0DO
SezWWy8NsCqg/SfsPxCkhEr4refKzxHDj7jWOXSkoW/J1Ghk7YHmFT78RpIZH+kW
Y8Z2dU3v1bOHXG7jdJNki5Uday3D7nEvkkmdP1/X2MZVJiPGlx5f/SmTTk7Ecwuq
gfbHys+ePEYF7L4BOwMJfeGTKvyyv4IPbWzrknk/SVmoFDn9ErJ2b36f2R1od6Ne
MFEycBMtxQBARknpyXrPa82mbHcNHrD0mrt8XGUb53UPMZYGzGN3HRK3AwRz6wve
p4RSyeVLgres7JtVNhUkZNQGtsO2W4OQsZEGl6K7kSt6NsdzQ64M8jiSDen6wSzS
ZaY5XVoDr/oNMcdUgcq3kiuRLEkQk7/FMi/48PDnX9e3EsynTi4gow3knxO14Mp3
RGrTWtxfOvFtb8W8SEUnxHvTnTQiMwxigaiuNlqOYQb0nl41sQpFGZWzK2jLEvs7
CaZN1zY5IsAvpeE0uXMrQYelFvwndUAQzzw4yAXkSL8y8LA1nAN3oJzKV6XxrRi/
uOd1zMecdimy/9qxDafNWtU9yS62c0/S5Q3Xczo73ecM5inkLaMJw92WVCaPdvTf
598NYIUvpHfGNJUYcQRr9Too9G1FTxdjWRlkN/VRdqYNXtwz7I4gyvdT11tasTVj
9MNQYGRWbyeuj2+AZuM3/plIr+p56wa2uTgRIcDXg95g5IYApprfD51Sk++1eJuf
3vECmTDzEnBskZJCo9qfCyy8ScMCAeJX0D7/0pZa94xSJSZ2saUGRYX4XNhvfThe
T2YRLlfYPU3CmTEIk1nCN7WF0EeLLnv7ke0my85Eto3F0LTeBUCqoGujPkhZPrNK
UhqwQBsa7dMP5Xf9ROWTROd6UAIptXrFOD2yh2vq/mRAdEre1G6xuL+3NR8jGldY
CUgm3NbOFsqX76Q7fF+QglrV+u4k0gpEbwo5y/5oS6KZp8RHQD4T9CeIsbzbNK6G
7LQVp+bF2uQun5rzGfPJaE6F0SeLnzKM72uc0ApwuL5ZoHVmD4ENp+NNGHsVwNdp
wFCuYVv4qtrpccVgwaIQKoRmKordh/llG3TMv537gG0eh41ATrsZ2CJhVrAVfjvD
ex3JJaoFoHgwPJ+QGEz1sBuTzIPyNYH5B1xV0nsUALDvkDTE616wAXose5tM6sUp
btAf8h1pav7WcF2Mkug0oqUa9DqYzVN8/jsc23p2FoMULDPPZG0LuTx5yIe6kSq4
TfE81FCNOAY/UjcNXOmHIMvlykcqhHyvrxnU4QoD6nWd42tLe7xmw9rDNvdFbLMM
QmLi7SeGPMUoe6lWgowNUFImRs3tsuuXFsnCVhXYxlXhDVgHggrJeElPT9Yh6P0B
+e2RqMcsw4BInfGsXF3rkoIDt0U9l0u+Ih2JoIuVoZs9BIjtEVfr206HGUDnbVME
LVWnAFg9/wGlUzxqbvCQNIj9N7TjAE9op+D6ppaDvciOi14orzM/GvuRjmcR46cg
ntEcYcEg3F4ZAJibGNbl8PRmtCNoP4qQk7bsp+QEJ8QFF1F2Fbk7Jg/C4PfDsK+1
nFnCx4SMwJo7j5M3bY1fGqSIGQFW64E3P1hswUkZ1tB79N/pULNjwxNCqdRobRqU
be75OSkelSpYZWUMVfBlsPEklOF2z8KfxiUkWiCItEpIJGUyQ+ltDvbTO9tAbsqn
HHqm6ZdfX3CxVbPaQaTX71crSa/sr1PNz7Z8UMkLmPoYBS5lMzdPD5WxogBJuPXR
kqmaqL5okS7sUQDl384E7NrbanZny7Fm+Sm1ZirKS3hAw5ke2JxYVg6ptmfmdqNj
NrTyD2PbG7EYuHB6PMNoP3oi/wysqqCi+hyCsgTZZWkjaysE+7xjZKe6Tis9eokV
VHE01YmI13eeyHs3Q3Xxd2oP996wDeINWJJ23CilT1bMixCZu5U/mKIprZATHqeD
8hGyPsEiCbo8rFxw+5Djm8JYuATRIwFEwsuPdg+mQnDQ5H5Aao/aDVYCJ5vcZSrc
sG1CfgQt9D1tDuwrwhOcHFjEu+3kq2hBcgxIYSJCoFTf6kFUs3Lcqa8INKfgy8MP
jm7aCqkTLSOKYAYNESJkIGyiqYgaVx1taLl+U8B3RFMHNO895j1qXYdD5iZIs7B2
B3oyXgVqMgP/595K6JYqyP5OzNOESmnYdoSiaE5uSgS285UgHOkjmy8/83ryeMcI
oajuFyKb0/6Klhx+ySQ0IMx70FP+cbreh+aueaGxSX5aJgtTp2Hm6t4UYzbJyowc
IrxoIdW35sAUPXVDXMXWevHdCYde9Hn2M+LJwFNaIMb2dgqeg41nSWXmvuiLlry4
xCnmyr5TTTu5SJZLVJoz3RVxy6xVFCC/Oz1WnK58zqoDW7VqZO56m3R25CAD7D1l
mcgiHc+XETw8ryvd/TExmbGGE/ePTWSCVebwVRt8ahg3y+BYlA1L0oKikw+x6+ie
P9RHvtDHLLuVJ6I3aon6LFnBor58Zj0CdS0c41M143z+RMeVTqXJxsSTsX/pSQlM
G0KI0m/dbvG6rNHtFvvL29AXC7vekK21igmyhWo1GLmVRCVPSlFfxr4dFXbuRAUP
so2AK5uifa9OrErk3xcebCpTCPiuObUeNSzQ6/wCSy0Q9fo7FDA9Q8yO2MCozwb5
gpAXErTOqcEimzN8IheZHmI4qoZzMW6eekBNPoVQjTKIvKLPhqBIuoMwJulDY85P
bNd5h5zhyeKYVDCneg+9HZscv2n+kTgSQJt2HXald8t6Zs7c5frt5WnWO2mQAZXh
3qvlIG67IR6tl6UwgXi4DQhIaEABw9KiM0YgUKjsS7+WeZABGfxQR6N0LHp1Y5wq
YAPS3PdVogTmJf4PEw2ske5kpl8bwM83nCEl04TpjBZ1OPez3M3Pr2KsMb3c+Msv
E/br9kB3jxbhN9G9VJTdnzSIz5BfVUxVz9iXuaQ5FXZVZ4MwTBWSJiXsdWFUIhmT
Xs7bPhf8qVu6WfZ1/3G7Z4vRO9HL/f9+vKlGIGB+eu54Me8Jl/oiC1iB4gdd8drM
DDBtC8qMibe7g8lykf4OSX5jx6RCGjItAzNgD0g7PEGJ3KCnfZA4cIfCk/G+vg1u
KjAT+fNNFZ4qzmcmNAUlXoSN3BtpCIN1lnTuA4TZckSArtISjz9skPXHYy5Xru+h
Fet8UYf1pcJnqgxLpdYnCjVivYNuaPu+Shc0XI7ImxdT8onWtJabxHnRzi4lgKdj
eRkTmnrD9gM8fcwskkulb6PMRPNhwimQBkTf5l4qUjHRGMKY9nbEFKn70zvnNiQ4
a0KfUUPyzXQo2PjOxm7+V64anCyandGoB28sErzKJbGeg4PSCstesHzdVNeHRbnm
5QafYuzPdECob4DvWKS0s0Ikj1hFMB0Yuk/Bg9wBM9CQVrBohSjl0+jtqzbmKO1o
uzgLE2o7ntTbA5Gxefupk9MXzzeD04E4ZCcobk/CSrWFCx7Fk+YiPrhD43KXMvbY
BDG+H9iZGEZzbeNp7SAiwcGC/UEO5yty30di9WvDNWrsCkqUdB9COjH1yhSCi/SW
GBqf4HU4lc3VEMnLTP42eavu6c3N2ManTuNIoKgYQ7SbV67rwa1/lYx1JjYwBHZQ
iWuUw0Kq/aKtDnruditXUpd6Ezv9pXBHVP4vZKP/To+12k6i7MkMXNQVX9c2sh0P
BPpUSXpIBG6EoaDss1ZXHhoJb0X1COcpxaQ3t0D06sRTrvSxf7kRdk0dZ+biFilo
tmCpbS6sLXmiiSB/UklW1Y4AxnoQYL1zdfAn4SKSKCXWyg61h/Hpwe0nZgzxQt0m
cldMMU8bh2UeWS0dJ/LvLCvO8XbJphXzNV2P1+gS2WYDArJbKaSxnQPEC+++A963
MC7+kkLJZAlR3AHFxblv68EqwuYTAPeXGNapiHDszJnU0A6trUaWkJePwwpJZ27j
fyumGbOMfbsTPQlr3DpOwdqrpOVMJULEOBtZ6CQ5Fz2G0x17A7c58gn9rmd4bixl
O+Jx1vJ7kOE+cpLFj/SGCrT6fhW/RahtY/i3AnH+rHwhNmEMQwZ1dt7GEcdLDCni
/4Is8SarLgEsnZ1ZerxR0nLkPr93R3ciQLWPjNDe30oLrjVyxo5HOJn4HkYxzmya
tWvVaTSEb8PgcjjNervNeMXb//Idi36mMdxYyI1I+pIPLVhf3I0HkaoA7LcJvD8G
w/b+HHMUoLI5sEajMAM2AlX4zM7JL0yQu2EZ1ZDQMYqxGDb6Brgb1CBf37FJvKm+
YdqHjwj+9XrEzgGZWGJhBPgat0DujIowYmcKS7c57yTX3FxHcMLWbj4nWTRmz8et
DuCqZJ2zu6CHdmyGJF6R2KDX56KFrwOzcb28q9TWvd/py1aqvd7n3v3keODZQtjT
IfGSf5NpxUOWdmso7NJ52D/0+qWibUSBc9itnYq0xEKyXTPw5UgPWO8i8avEIEZ7
zETNucKtXD56025lG4XoABZErtucmA2pbk2csxnq7bT2ectOvBsqMhYdyhmDYjTr
oUMObHWrbxIDoALjOUqblbL8G/2+QRoa+tKidrO5/nU5D136DygBiov790ex44Fn
whMFotSPn7oMCGR4ZiY1bUQA7OxMU6jj1WkB4Efzc8Hvl0ImQ1zX4WTqL8fkBKbD
rQgkiKZyi/xlfm1Cb3hfWOJO7FXPJJpz1gwfnkOOlqQxy1LBbYuisU3JyyFERe87
Ek5k/VItdKMAg/1NoFs6kB35E6Z2ZDpA/6eZ6XhcrxX4Hrw4yZKQWrpHw+ZJ+Jtr
31hCLAgNIeE1isE1tguOSLuDl5vq9fOITN3+a9uDkrIyQ1kSsxttT4eGf5HSA2D0
y9s1N9sabM2vbPw6wxPbX0zIUHdFl5Puo6Kk4rRbEkraERr3/2P8WGQl4S7xZqPE
ESs9Ht9OEk/Hxhe/8xjV/WImYOqO3yA2NfWsTzV0SFEsAUGw2WPHx7Dyne7LSqXh
iSpk92DPmkuutSeOig+SCjTMRUhXrW71vzqpyP8dnd+a2Yn3MvaqCtJz2JeQ9uO2
2OsDvUeD8dSzxEBSe3Flv6NTNXRNrhGIBn8YcNvmzXAPPUQNveYAowkHyzzP/fNs
DyVjs01dT3Ea0Q+66QD+4+MaXzDRvdXTAalzfhLv90f9gukDEwNphN7bx/kfEAUU
jcNKtp1P9K5k9uDGs9jTSeCQEzmlFaBOv/Qfb85qZxUBE9ift3O6H6a0zOj72/SP
zRMSLdmnjGeZvF4jvhjENrYtT/n3yWRkejrqWQm+6INHa8xd1hqqhpuPTd65+0fA
NSE5RhR3vhUvttsMLwwVx8y4lABWtET5XPuNJoHmvvpsSq3Q1Lwxe2HUXKTZnhk5
yWEU3AccE8bx+ngx6Nnk7J6986VArL7Ahp6KoXLtbkSkzTZQNoLF1jYIemVEq568
QLLYlP1WXbfO79ZZOR3OJ0EuHb89rFedgImhDMedQYHJIm6oU1JCXD2LgN+jTqfg
Je8CoEuw3bu/fgPAywxrZkAKGX+FKIeVZaZdETm15uXpxYixlFcanq/DciE4Ypv+
AYOAuCLhcCsKQdoQzG0Dk8T9IgewVA9of07g7M1SoC6vZbsxe8xplMxlOMibVrxv
HPceHZYeOVXv6YzvAiJcZ50SXpW4zAdmMXF2Ec4uY30RqExQkxaGdU9r1hQ4iwAf
QujiLLWWyh56kUqebXLN2VuJnlYsdkoMxXiRBWB8/G4fe4mRk2dzIyB9Ko9DmUBM
pghmQuVo/MRZDoYT481YfQ3nvhl22QGkoPmNF8SH5nQ8MasOXoRzWgOdKqjp2+JS
Cp7pGVqA7G7rXUB4SBV1ewKCE6G/S0RQjr+kerf+4s+gSpbaLjK873CzjJG+L93a
zJfP35NXk+GSyfL5bLor+MvwYDJ9xUNnpYhar1m0gF/6mOvuz0KsRSgXNyDMOSZ5
IMfWngL96/cfutSw3M1T0CpZu64CJzeKfYgaE0vJyevHbCq/Y0kUOiTpKtPxDv0e
yLKzBm2AavdDK5DauWvNgFoZmZjyEFWvXe+qSnAMu7LFzsESXDmTl0+SB0y5MI4+
9g1Pm45cY5+bxqHeGiIP8AcPWHUY1k8KDmtmo0CZSR3g+nGfUT1JLeO9T6Rdrgn1
iLz45yotKmWdKScQ+WQ+GnjN132xAr917k4J7ufa8jVVKLnZx+AHV+GyFjDiqGzB
DPctNKTFZ12NFKujwSMqn7tlZH/WD5XfP1diBiGC4Tbuzm3xL8Ox/MUK9X96cDU5
JA+JuGbHW3ijFIZkQT+SbsnQZ8hL2cRyNxGDI0ey4xImFXIazB+L6APGH9GtPXbJ
xQYRbRRg/GQsuCqjgbpow6VMiTJHto52hl3cjs5fQe6R/leGZukmnwJvmuHz98AG
lU2SK2XWFT9YxFx0gB0udm7YGgmQuDWS2TeLF2ov2k+Q4mVoF1ZBn9qIjXpFe1nz
jabIacaZQACmKDlltfgDV8gd3IKQcHBfr0W+KEPDUWybFFyYUD6TbcsWV6OBgYYS
7mDjTJiaMxUfrsbpcfy98qfRp10ERetA8JgndHCndrPM/SllkkZbz5vuA2fOGL10
7tADPftkcGIXxPgGJ4ROhBCz7Y8rSTZAsdTFQ308zqHI79qZ5MoqzY2fZraeUcvs
WUkLonJj/3fcRrDZKFsMWE/hMzmRaflmWj6N5kqJmCZMaqIn2GKqIvWukrKslCUH
GMpMksYD6Z2wFwxTYsf8nfl4YQ4DcEwYjUreTs/aw+Zd1axwq9P18c5RnoKOy0uq
5RbskeIixrCPGRBlqGvyZnXVTui73/dq3yfZeY/lKxRYXGnYNst4se25ZVUQHgyE
QhNR/Edyvo/GF67evVXYM0b5Qc3Qn65NInLHO335jn1sfKXYafCzn5GfEDwu6UsK
ZDrxr742El/vFQlLV0HCMx53xrEYSXY3VH6rYkukUDOc3FNhHRYPeW8kJajRhNS2
0SrfQ/chXv/AW/MM4nnabYzM7C9GoDF9S+NA2ilMEVBFu/SQX9fcO1gnxNmA4UyD
PT3cNR8I37OojhS9vX+563A/k8nDxb1NBqDiAiBmuDeMWhUF1MHMGkkL1TPcXnrQ
lL22eiW9MYgNXekzbZDMf2d5THqr8Hw2hiLs9kU4RV1EpH3vYTeDpGNGp3rErffa
T8xUH3eSTFS5U2LK9PQspDmuE6FBl6f9KaRQdmDTMPCrzG6e9KzEQyWLxdloBjLv
pRhd/+28s7L9cwbAhQnt4qL3W0bd0W2CeSxz1B7ppk7CGJ2l7AsllNPwAcmJfpjF
rHLVFadFh9cQ2sYQ+2krWtj3hgJ+ldgpBcZc5zz8lg2ee1LYFw62btgO7yu9sqWH
LURiDSV3a8Ye9iCWlFS8IV+VjHzp44kiScAyXz2wxuL4clWzfI+SKxqBiXip+ciI
SG8+kVvUiQVtp989toOfGI5PipdPrLJflMdR6N+PMg9mAGzBP9FvJIGk3ylIPC+5
T4T95LGYFcavfSl86w+t+3yLRVbnpTYL8e9fdwPE9iqSOHTvufqIJolITkxDHCvu
vltYVFhDBu5SiBB307BtWpRv+1h7vJro9c5Y4wExUZvG76TzOWzmJuxouWfPxYFk
tykduvuuPJx1WZid0jOa0V7xTtLBBaHj75uv2NaMPsWg4u/0feFwkvmTbJ+oobl+
jFQ3E7rNoOBUPY7tJ4fDcKxuEkj6xXk+FvqkiWqGiP5D2MMNpY3UrT0HJmynQNet
hAyvHBqovsvSIlhi2ypWfYCBYp/pva5FwDvSWQqCMAur87SwVBAjceRoHa2Ltqbb
EMABySkNhuhXEGJKmOzT9g4+OgYASJk0vAJuVip0tIXpL4vGEBKVrmFr+zTIVpX/
WZkUVnoqWLUKNqjT1IG6d9Xt8VuEPNb4BsdW53cdiOz1F8RtBldHaL6TYBXXym9j
lj9mDbUNf0MdPpyIFohsgJXNFw11fH3gaw3kZY7qzi+FQiFm2+RCDB8n79+V+zvN
jx9VN/R3QpTcW12PtewgNlh7yUcGRbMSRc2Z/cpLuhNrostzN5WV7TTkRECaZdzc
dGiUBDfGGEuOmB3zIZPC+MHO7HBai8k71h956crYD42TGKCnt7nryLjRMOOzc5OF
8hkrUx5cp7Zaa0vkXXlds8Rk98NaF8f2PVw2lB5gsaZyNEGk3BRebcyoGE8sLuwm
CyXDUynkQj+pV8yyqD64t8hfwJ7Xwwx7xJVfCxWwdRIGtBuJGT+TVAGEAh0W7YHY
PzZyyeqr/sSNBJLypYqDw4FOxz6Ty6VYWihLEAI+NwmgnDPw4SJ88Npysp8abnZb
fHN1mEek3VgRj14VrPbvmGyj/qm+GGPU+CnIwRsvMlCTnzCc8yB+pXTp2v22oN6w
bujF5zbbpq4hylf7/DgEFo9n8RkGhJAtvy4Nk16YCi0wM69JLb/z7pvllBCtbB+R
PZPNmIcPGUlUFP66aEAK3UctglYDunyZoQZSq/vJa2g9xwowx5LgWcUj8l3J4b8l
mQdzhaAXpBRaMx0WU8plTtej8o6RMVfiq0GGDgRNDBQY2E69IDotvp9Z+8GGcWk4
jh46G64bPMZLR7sJd+fxlCwy4L1Fhqby+qA3NOaePIXhqvEX+EAYSxpsTNhaS02w
M2kQi/dKNenTEx/XaVV3ioGWtht37LYvpLqGYtNVfPsqaneGwwkj2cyL5rSoGqdh
ukuNZyXC9YXNlF1wzjh8rrph1zbAcnebnqj3abFep9U+KVF3SGkPUZ52Ut2TLlxa
mjFw1O4hlVc4QCo7qK5UHiTQ1Wi80rEDMzhpP+jboa+O7vJTa0DSMxsaH3xSxwPX
08xgNPzUewbHYs7l66Dut/YCDcT7wThmoPuI+eMzqpI9h0IZ2qrk+U8F/QFXPXXa
/fO1vTYj0qQdYXbpxMz/OjE0WX3F0XF08x7lRCzxEX7HB9GhaTJBoo0T3qIznRL/
UcPs+rWwOSl0hAWiBkBtrEBY4a/J/iP1WRE31hZGm3BSgSi1TODoGh98LZdQm7p6
qdRQQ9ud7701ed5VfSox0v59a5l6uIDACpNkfxRnj75TLMhRwr617Dy0nRqb4/5C
VFzjpIbcEUcVkaRq1hzhhccmzxcH7V8rIYAoWkQIRtWWPXa+STzrjbk4X9SZI6A8
O+0S1ZgZU15FhVslHxWzmG2oORJItdm+lXI5weN1H+CDMyOC3CLtWKx0uX0Bule1
k7d3YgTyb3F49UNQFncq4mIzRuMhfoHIMTuu5v6xF/qT5QYMMl/ia7Bz+6LIGBHs
TBw5NUpD29On+/j5BCqFVWIzoRvtBUPsu6vS71j+2K3iNWDanBngQ9YmMTB0rcwT
yHX62784GGksIAySBPivpSTYDXytl4p/+VTrTYYcP6MWOKK54+TlrzNqp5dxJMag
yYvw6UIMvDEl06SVVRFGhe6+Y91MgXvcy2EEm8xF5CBp/qyf/XKNoFIWrwsYYuDl
oVVpBmfn4Vb6dQlOkX4k2sRdWAX5O3L1YixHCrLMeruTIYHut1k/VxzJTqsXzu49
KpsQLkvLM3R382NfWi2MXopTZGQiLcs5yMt8EQf2aKZOOkf89JzPgxZH38F/dT8u
UxTFOBw+BtY28C4i/3bRH3S7moXktrDqYgfGxQnNvtbyQ3P36adrdt4Efyx+2QuY
leh1xt9niq18t1NE06n3ReAgW9q0NCTPpPE4RO5t+owLeX+EIlx0h6dAYVxcCR4U
HPJnD0N8egOLjJKj/MKFO6kvNLfxaVo9hEKbMp2I6adKw1zjB+bRDbypAX9kXVTf
RqATl9731I6dWhGDJfCXN0ZZ3CVI3lhVnDyAuF+ZNARrOxDXGviUPScfKYynq7Uy
k0lctG3ZLuYUS++zjt2Vv9NEP18M6FHn38EuSBA2iCTatmKQ5FvImWzjqJG6NsRO
8Dk9xpA0ae4BgxGx2TN6Zhhf4ojBNXOna9fXts5e8XGP7RknxNq+FytVUNyad28b
uxN6KjA12Is3klnJi0BqIinhG8cYlEeSq8A2DdPPTuv6m93EXvmdlEfMhKgaQs0y
8zpBcl/dwkdZOC25XuDscBq0xFKfc1qz2C3y/no1/fYzWCFH85MWJb4NpVC5Lk0v
sC0w0G/Ax4DCjpfXzmgpIXdHp5aMX0bEN5e9+1U+TF/C95XfQvuwea2hQsY1lz2v
ixlpPIjYX3G6xnelp3bu9gLmtPfVw2HDC2nrIvdEbtgtb6Qw0BU5lbRKswDmfxiS
2OS/rI9UwZ8CddEieb9sT3pFZ8JwWhHfOKpGpXeTFS1KXpYSVsugwsMhCfotAJOY
mKLCoyyhdUlrh0t9fTZe4WqNIsT4IMEVcvbta9FNjC7FjvJ4oViG1FRZCZ6xaeia
pF+G3i6cbHA7tgM3oG2WtsnpW97lLJxaawiqq+FnnwYOK/3ToDngrVifBm1JNXS/
IbZ3Lt5967q3LdElTS8D5uh54DjWW2swL0LPnoORZcMxikzMeH9W4KEx8ZBKUQPn
L+8wJ5XQgz4Nah9skWDWI9rSrGnj+NjoZ5UjbgUsevkIXfYYLKJeVZWma2DSBbF9
mY5KZggkZfdZdxPaRUO3nHrS0I/2GrDVscE4lPYLEHSgK9o1vTzqewq5SVAfpbLx
soQg1lCgRMGZNmHW0hfZ98djkObPsQyv3hZR4kwrfGPU5Dg3LZNe93OBbvQN+M83
8o+b0T26PkQ9FhkVJz2hgkObGn1t8RtuiMCua6slTm3BHEW5sKMlGZhjiFpLr3HF
gAOgV1jdvLmIUX8i9zOc4d/RgCmSZ7KWo8l2CIEpGcQui5HEG/ETgNzZkOpWfjLn
46CPzDEDT4K1+MNpqAp0H1SyxomvIwGtde2oNisb4Y8E/hf3EvWibhyIjocQp32R
PzArBNkQmrzmyFI4t/H0CbnM/EZJA3L5VtnhSmhWV3nj+zE3p1bTDRgb08zcY0hT
1hmY18CvYPL6euRcK4eUWEQQu46Fl0V/D34yKI3P28xiyYAGW+N6kdKGOhAq68bJ
tBcRa+rIyLX5QrSiY6umqSXSfYxO+cTigIMwVkrREMLC9kPOlvDEyjZfYZCOcphP
Mb5IJ/j2a04pdZOBeiuqnTPrQEU9r6atjMiqPCff9r5FulMAvsjp3SR+0vZU2dhp
/+4cyLv3HcQg2mntIXFmy7tmakfbs6F9+DzZHii4DaeRg4ubiQriqxugnOyDYUCP
0c+dGfGW0jNd2jsgp1am6zCbQm6PJN6jdui4yPl/wdkJtDcV/uKYM+gOzwOidudD
rxf6WWcKzKq/V750r830hyuDwh/yDXMVLBFVRDVtnmw6Mb4MYi2MGpkMM1TcZOn7
FtdG/YDUwg2nsEo3QEMp/V0iLO8jQ85KghZ/4x2L3MVmmWemytVRXermCoAE1U2W
N2yg1p2WzPG1PGYCTfeM0pzW4YHelXIlSPTfD76VGRmtrogvxghRGNaygZCFnUcK
JhEfoGsZB4CD/EFgiODlyaDC3Xi5ZjsLo4R9fj6+NwzBIwQgSDWGtjlP2djo7mpk
/qAsdSh2JWaSKNM3t+hqW2Zw5GEoh2RafRspaBBG0yF6OUi0q2Z0gPRb7pou6V7X
mw1J2N4EFtSxbNF5YH69qedCIWT4Ss0nTe25eF3aw8mLFvcJaC4P4Ii/4rk8u5Mn
/IWjwn7oCuIn5A03PUyumD/KGHp4FvIhCPo+E4ko3eyOCSFqCLN8ZlNyGuLO7JMY
a1LCIJ9i2XHYPhkVKt6k6uhf68Qf47Lj1YUKdeeU0zI5iPG30pQaNOU71YdhLpIb
mG+jdBkOgRoQQYviPxmc6Ks5ctsuqrAkwIkPYv/I0dFvYJT8FLf97AgNuYZ1gbGZ
3ItvlIFqyAtNRdjclFzg5eCyCasFqXBU5TV9dqMXt2qwsLBb3/7Zli+Ug0c4jg9J
LXHoa5QyFPk8pJL+heX8kKWrznUOZ4JWtCZCzq/XBZkatPU8WDfPwvb+3pEd6IFd
sU6/sqLuygmr8nrlREZRwRB4ueoW6NcO2DuxiNn/1he/END/vQX5bolHsUtrpXhK
OHE/UaQDiHBhaWB7ACw39yDEmy9cpZszXXJ/Q9ZLo/WWf14Q53ujSVOQI4RfBnKg
DZ6Zb6/o+7Rvak5zVabEx/TMEkCQnPdHlCNSdeBaBCk9HFh3mhKRctqNFuPMJluv
GDeRAa4yFzEGupqD1Xw36iiuks1P4dYJBHNM9jYmLDwnPJ6Xr9/hp3VSkbzaTIxv
aQ23m5POg9r5EstGHU+aOFC+BQsPQ6GadZYTpcgAXFSowRbsO9MfGNgasTSGoJoM
m6oZtV8t6B6K8YyxhVjtp9e4X4cn58c1zvjLckrDGqKEpaiqV2cpjmEUy1ke7DaT
lvu3SzzMKPjzQHsWtp+SzeKDZ6bthaRrdylt65NMnQwfr+Qdy95ngWZnMh9Kfk2k
rNJZpu9c1/xrhERRusyYnlcZL8suGYBA+OjhQt6zTJKRiTTLbpPWIEFy2nqzCJPx
00fsTievAsiQjjZVY4UDTBcczjxo+quMvSCpPkozs36k0beg1FVhLcuTDOYTb272
0rsZJg1VafDIJv/mwv4bHfbVVwEYNcY6oC8b9WFJ/UxqT/tqgteDYB8jPyoVa9k1
QF5rcxSp2Wnjks2KJaROc1+negXeymrA+BTM7prBnEs8hkw6UkhkIEYcCSoPLcvR
Cbz8lHlHGWRx//bnByoPHKpj3Hd7MNO5zMm5vSmGOkzNvLYKxymGyh0P+neEgqbw
Eiw0nyva3cb5WNKRtgN1flUfd51bdCjAzbV6/14kL/LATKAyav6+RxkfYhTkHwar
ymtSqW4bhFUdjTob/2tT/ZJo3aEBO062DgiVHBBXz1fGDnYYNdI2K62SASwanhkm
Tw1E6jm20LQkHj6q036m8cx8nfv0aSwvd5eSZak4jSoxN22NQD901doh+qY5i6bu
3xMrXlM3s2WnB6QH+IWGxkpv14yVuw7Pq6FdkaqjU1h6Lcfm3i2OCoFCXi5Y0493
AgTZRoqyNcrD6KBSjAu5hP5D1ZL3Sa2p58ojSzQpZt0TbbiWW48xFPS1URmttx76
OP5GNhya8OPZofj5jXfiRjTG7lBWGr0FcVfQY+705ecl06wBbt1z3k8wEyzAbiyy
o/yQXAPZ34T+c+UXowmxyXnMnfJ0S9TDAvae+b5cN4uwS2vDEcjKMs41M/tuOrHU
sI/ZGzKQ3EACmvibgwZ1URbP/m2NXhl+DgWnzOy6KYoBquIGpEMM8khS/kFY+dJM
kX0xs80TXZh1j02EFQA5x/is3ySU2PLOSBAIoTEYHfPJtBP5Cj21ZaC8XozMFcJz
jGWiu9iqiCrOV5v7sx8faayegX1f25Ds9d5JfgYCndsIepP0nGxAuy/9edHUEMZe
3VAhS+MMQouN3NI8cXREVw2NvaEu8heWcGQd79nILOz+7Svlrm2wWETvVigjNKS/
gzqcEUX62lb0aWXQOG7GOik4tirKA4bO6q5hNYFUvYE6pbf5jYhwTtmsIymu9oZJ
q9jCDh2Y3TXe75LlQxIatg52v8fDZx5cL2jXsItwdY2PYzGHTErAeK0ox/HeaZ/c
iElPPU/6arXTwYaHLizEBiACCdzpSjT72Mjis3j76MYaGnnNO1FJf+22yZBYS9wD
XKJmVzvL6zJZT7yKFFsDu1oaXUqVvP+G1sucws+bs86ZjFAVLs1KFiMckpGvlKOY
/wWv7hRTi3oA2EPEH2lD2sNslLpJ6TXAF3bYZgJzjigWNFXvmKkeCJdjr3mrxKgD
V0aG+VrKTzQdusb2oCXptimg+ndJ6+j6nbW220ov9ufHYsAW9twpErIHYHvtPtaJ
bCJnsePVQHVyC4401RPqYV5w0h9GD4BtX2Trq5fyI1FoAiFWJNh4N/N13YIhRFKu
pASa3e1nT62zxmtkrE5YvDuqkC0+TIsz4DRT9BJYWmXXt07nkQiFuHBiDM7FvYxp
XmfAM/Zq4U89MhJepEUdhLOQlWElaIPXq5j6P2sm3bep+o2M9X4m3ce2CMC+6Uqh
XBWnTkm2ehbaQ8xqbtxMxexPIYvNi3CmIid0VXPbg0Qg7YPunhGZ8rGqaIT4KOGk
ucfQsVD3qdEZS5YE3UdDizDy1f0bQ62aeviONh1exh+tuX22SI2X5nkfu4hk5UsZ
tJBcQE7TCRzuNIjVPUW8Ru8fMU7ls7Bii1CVvNV3syDnQisWZOac5Z/fj4aLF0/d
JlUJzZXdC4dryEvFRQu2uxkTPSLyITJyJLRQcTy0xNiSqbKSabpxmVToMX+gUvHv
rnYacvtqToELyAalHtZmCdPGesaM4P8JWUg9DOKlBhvMuUxAPoOvMdxR689FrUA1
BtfFLbYuJqGASzmkU0xloivd4AuqIKFVE9SWQUjM3nz/lytwOIlS7htJbZlVHlNv
QYgAJczS5zQVUEEqVH0u4lHZ6Vc//tJeNtW1G5cVZwd5ymOEYC/Lig+rbZRtwV62
ConHyfb7ADF7ZHkceju05cZiNjD1zfpzLCeimALCbkJWs7gIe7AalWBWpMfUPIEf
jA2R0bTPEr9/0a+9quj9nwyJ73B9Oh+3YC7JOUQjZSO2perUIgS2kIC8ofUwclhc
4kUZaVE/dY3aZ8ZI8RwmuhylkutZElrnS3yFcFBdc5Xlg7d/HTWZ73GOvs0fZxCL
ATC3eEESCRQLLBnFYQATBFVGtOlhGutMQKY7ya/DVsfNAZoWa1sf3kUqPFCKbRAX
5cQzN2ipV4bX19lSydYAtvzwRoibabxcyBP/+F9EnwisgYBzXvT0oRuLOEb6aMuh
booEgaaPaFBkWZalEjwlvhDgElGN7kToDEvM/RxQk5ugvw/mAptVJvz7wQWsVqVd
3yNT4ENe0C3iBeJ6Y2AQefaBQHZTQ4CzgDDLci8AMqtUYnfWsLe/SEk/uHRGhEKB
dgAtOSb5ucmQcUq+CHqNoNVxNfisvKqzsAZURNQ1hTVdzuH4jJ21SttLfhwXINgD
opW/fwf2eKlJfq8wrcCO2tmPkzRqJc37wNaDUnwE2jD2rn1p0yLgi0GgBMXaR0Zi
2p/czHLFhfLx+o05554Ma7cYhPIHFUwDoeXdvaVfVzs0qxVMhuv1dr494JfpstBu
imfGr29ISPoV6GsBdEgSQ0RuVyJ1D0nefOKqIhTDNnRHUQIq3SgPBQ9IsbaeIlWp
hQWH8cvePVVdyDqnMkIX1fJtIVLuQ7DT7QOODSs0zctMtfuYU00Ow7DRZ62W/mXI
daCN0Lz6gi0K/N5acwMllcRYUKEiwHVAoqDhXzf70CJFYliN93Ozz8MOinA79MuO
OLwVtxWU+EgHqc7J59V0rDDc9HS5vmERXtsyGda/OF0/VkMCCRJLRunUGj1PcwpJ
2F4lQU8eUZKgQX+bYjVsKi4zSp/qG1Ipe7AHBRVx6laJ4ZLCXydh5iU+iIeHk7fh
bKgfetE0VASaVH0JnGpmQqPiJKg40Tk/0LrqvWxJ3bGJhVGARrqYR5DHIq1Z2CxB
S6Jsd2NtD/mN33dT0mYTX07QUrKXqkZ0wLwNzFuoQC3uGc+X0gf3aEaAy9CtOVQY
QvMcqWQtDoVrFbnGSK0DOQhnb+Zhj3EnCudHxEDA1PeYM7OSo1LE6Lp7IVAwH48F
wMxdCi998nQTynbHGrWTPamGM8IpeAMBfmfELJxoquQRNEWGieZrKQuTpmorZuGX
1M0z+cf/uSwZcFNsokG+rxaE2S4CIQY/NLYQYUw/pvo5G3reQC4z3KJiAonx0WBM
pTy3gQzk3dHbBsDEpp3YFig0UCPvAUsrZnMiadu59kJBSlLC/bRq3gdQ5vY8ZRkI
fYYubQZuiKySnVaN2i2uvvXWWj0U93izZucD0QJvknW2gowQDXBtRbbewU5EJdFO
0Jrts4datHaumK68HQdD/bs9/+bipGqUf9S+cOwXPS7D62GkibtUILQQORlbWKsg
Vdu/YBvFcVxa9FIveF6N4jqPfBcu6OamaqutsXFJusxafF0rBH5sZDzO593e/ObO
R+7p/4Cd1A/B8jygdwA/3fU0okP+6iFxw1UQ4txPUSxERo9qDlIg0Yg5xtb7oqm6
ElDQKmxG1elFfyG6wA1MgGYbDjK3gQcMkFtY8gjL5gx9jVhOyC0BrawTHvmtZMId
tIwSFoSrOLCKKMOi3YqfjLXt0CVbp/hW3iN1tVm8D9SIxGI3mjKYeEtyMz9sxYC2
ik/wf8P5uc6BS2zJHEPPPhdaocrjrwNxMgRvriAfB8/I2Oc0WIZsQewiwm187Wk3
vpXue/QwhFmUDKwJpmMESOJHlhM1bMR15Lynova7zvYvo9Dwy9Nxgsp1G7wsgd2V
mDCgO6gpnZK+VG86XJnzjliMqo9/ryPVp4YxTTGHB3HR3Sp4jF0YjeHblazMfT6P
+8O05SlAuFRgosfG5Cskpegjfs4ZcqoR8V2c2zqELGolLZbTcbDJeh5pCG3SXU5g
cLEwSDN6WxLsp8fB801JXTVGXFxTsw7etYbyO+4cGSySuluizdg+Nh0NBlkqQXw8
Yr989mmZszsoKlwdhehRWS6U8mRVHHIfIG4xn6VSt9z6MIL+r9IFja0j22EyI25R
dwgPNg6inZN5721L3j+vLWjD3YzKbsF9xmebwytP0LjXR4/JXlK6XiHowfRU9Oea
cDjUiabd7I7C8fDptcIp9qcJJOr1hh+AxrR6z0trfDsAZgLp6xEkYhB+eIka95S5
5TgO+4oo7JlrhyPMnp9Nzv6KGTwWi1pwkcj+NQDPJN/QK7f01rTk+rYfF0VbCiHc
g6Z3nGIjmy5ynC7O5FSO+ulr0DBj1KiYzn0phKDdSiff3FCJ7es7039Eein60aM9
e3fis8ySrdFZGZaFPEQiZGnlU3pKzmtjxxfZvnF8txgM8tUtTnH8OtNkuSPMKGhh
YwCHOGwmgjyXATA4a/kYctaR1a1UHsdm7Z7/cFiJauza8TEArxuizrWbrT4OA1Oo
BqmA+750+OaAnl9CN0SmdYRM51xtY2moCInoyr3jmYFjStMMRC1rnyYPeBeiKb67
LRM6Ab0M95MZXWUfYNMEEHUjGlITzVVZA1hcglsLA6MIlnN/d+jK/kDmFrLP97QG
8c/9F9FSB3Y57UfgWmd8a9e8hA+R8BrXSwzIaDGb9DQbtkQ/6PgijSLfvi/4D3i/
6Dfj6z+cLkHj4dz7kVPnrwVFxgh+3CAONC6YgVop/XNsFenc939DpdVCCZaV3Zqw
v7rx0n0aK4ZJWoOotRIA9HpbfVFPpCwK+2tv3Hk/TIHL/e7PyxNjjat76T0ITxf+
KaYTtUc1aRjrQ4dG+BfbYh4Zdza+a/StU+LDt8bWm2iV7G7I/wqJ0fYi52sqwYe9
Qi1n0KT8X45WBcEX7zTMGLMsXYx/JkIiD9XkVx5x58qTifZG85bgd02VHSpJbw2J
vS7fjCezgBphoQDipAX78Lp1i6tWML1eEZrFwiqXTdVd6mOMyO8JTHX7GMVuS0Jc
95NIiYlJ62gmvarO5ZhN4h5Dv20WUbq/5IXu0gSmXGsYS7qKQQLyQ9qIb2j8LqrI
/Ve3mKS1Sc4i/DChxmXaL1jbAbmCH9g5eiGqhm5W7p1KusiHTECRRqAbJoqbhmrt
ilz0kYzWBnkuCnKUCJbVSRzcqnD0KJml5qPYBzfFC0bA55ARE5mXIYlWNTmE7U3Q
cCyED3q35HLxBdeNQYvrS5jPXfKI0glHiw+/odyg7GAOE/iiG3mU/BRtzW5m4qwG
yuow0f0GmJvJZ1zvgHnssnVO1YApaD2OOmmzDoWnolc1fhO/4zPQQ1kwxGJvoPLw
I41o4r6PVG1Dm+XrYYknPqkSoayVW1kKOm21nFT1X4WgkZF7a53uCl4sUaYKZjFA
9fKGQoXFjUvcjAGWZd7pS+AtCUQ/yl0+dwTPf1wvatHIodhUrgPj8MYfBrt6DLOC
YEeq4M8IS6b6F/xV5BIDfvmeDz+kiNsMMYjtpVAJF32SVBrZ77VRBM2Ua4eYDm/k
rrPvlBfi+oDLaKdRVbpKEaozaJlYof6SCkQzdQWQn1O6EfSFQXQn7ksQZE7tY0UE
Q9TK/syj/k4rbgGo+iM8hAFcv+DtoDO5xKOCm+5CM1UDB61RLQ9kNWtl9suSZM5D
SgOGsyZEItVJmv1u+3D8WuvJ7/r7y2dxTqDutE1lFzKw043x9eQq9MCv+gytsjPs
ku0JbtxfMfaXg3+a30Gc0FfV85z9gTQLTmhr88XcrYdDYNBbhNLmAXMRw9Ef2Hrc
fTYmCV8+r1xSBTkfY9reBwgr5c3HRQWbSbPYPvoH/HhUKbTLhbgTEbONed3Ji/h4
p056MXE25fwhaGM5/nST4XOpBcVsWQ31vhuU7+b/5tUrftfxsDEs7xEvsMKpP2Lz
RdB5MRta+GGsysv/xgL9eIHJ+K//uQO44whFW0czLnJ06Sfe/pJNKTHkLqCb5Idh
IIeMpXRpZ1FhX9Z6CQtcAq63438mXDs6XQHkzbhpKBld9grCWf6G/6INUaPLIS/Z
D5sRfGNqJEGq6A2XMm9xxvRN2x/cfGJz/74X/bSnj4IjKTQmWOUawOh3HXF8dgHX
nSHMnwwrx/0oTJ87sqorR6UHB29A1gEDWRuhJfi4bp7rbT7YUbEk0ueKbHYEVD0u
z1FfXiSH5c/y7+JLESsjRlvr4PFA0DtsXmXFvXWpE/3YXkdQIlf/8HVpfO2F32U+
gGxq8p9ubfk0uhlhITWyNBJL2yi3HH4u1O0eWsw8KAuADhaDb+jI3HQ+EzogTE0N
nhGVYwmE9p6aykUV57elOfp+5ZAsO8DgltiVK/+WPVWJog4BZwJ5BiNNit1ExiIw
8GUXmI2+KjKHAnPj0pqCl5sFeLwLtXZBCVS+2ozfpOABXeBFA/b8gjF4aOSanyJG
dXeAfEaKJGahQyu9Aa60zty6j1oaz16g4+EXuGduaB1prdR3WXNnuJwBxhVOhXLL
ZGS6NtR3DQfAzF9S0VC2ZQ12tvku9Cb+Zwtq+P3fnMZJzHMTSA0LKwRlt1d97VYC
mbXrwDlB0X4Zg9pLtC5ehFVYMphicTqYMa4izWh1EJpsouB5Nqup/2LXraaz9LYf
fdYJA3WBAsFMHID5sTC+/sjPjnof7K+93hwQEdfLZNrO8WMAy24grQnSm5ctq+eq
denV1trYleAbp/6kk/5i1ojBjM1HmWQZr0F4jEsdmVX37onBvHv1Mc/4Bqz0cO3q
5yEJj+WFV7TrDK+kRWEmGhATQyew9pcPoY3rXArPI1BIYyyU0pmrcZz5y2QaPq8Q
/C1CDAdtvCog+8QGTIJYynDTDc8Tb2e26qn3qlPZ1xEhv8KEUnq7wwJIubTy6IUk
3nBBgprWB0UgkJliM7uK1p1vdtmMgTpRvec7NPiFlTW7DwM5di0Rjv0qKElq7TbA
ZLm6qeEQiannI/6x1wT/liy+8qvxPBDy7j7ncO4psgz5h+HtY3A0TmZE8W00DXze
eb43xiVNzSHJxBrE80ZmWCtRBgIfNKHZDoj4OjI6XwXu46ue12to//2vvpc5yPjG
Ef1iiN3svrPw/LCN5IhbKzsfocjChq9WthT+zaD3w6PjND5CXXPe7Tm6VDloBrEL
xUFbBLFC9sHJH4IFiNn3QtntvVjy7UUcpew3xLdS9VznjxqDDjR84+VV5HXwkkHK
mRGYhvcmebivIL84KphoKAieITg5Q+A6fhIGL9zakpnOROs2pomFCFGPaDt54s17
zcEhZKcobMIssgN2ZAh6ZLbcC0hFC8oL2OBSTmDKIUgA2SWl1mB9SpHOtRCisms7
owJCW4h0qF5U/zoZavtl5vkQdfimwTt5JIKVap1CCCQa3RETCWi2Oi/xHajlU9WH
LmcjL2moA5cU/UkkMn03l+oqv5FtYPbGsuYnlKM9RdYbFQks3a6CJGiO6Or2q18P
Q/VKDoZ6W6/YF1V1OpMBO1BFnAyXSl2k0w4Jl3zNV5lCbTkoCSto4QGGL573aUMs
2ODsHGss5EJfKAXfNLcRZ2BT+r4IAWrMEjyhz7niKZACpyed+OCN3P7l/BbthoNj
HCBZ7Kz6czsqJGC/HspSM2fSjU0XeT6vTgvdRTR9VfRCo3gFGIU9Lsy1gzh8/Bj+
qiHBSeQSiUZWDReFHeUhvI4NyonVQVNyzSkqLRsGkO2Z5zpBUYsReEoGJ5LLMjFE
lC0OnCVRZOt8gJEq8jqVFmWJMNMBT3aEzeI5ShQyQzxmTN46XN8gtttStgF0upsj
DC3dqhFoWIlPiWe/Z4mA3pNgW52XW4AkrSWMAuXY4sLtsbbepLWPKbfETRSxIdJ+
V4IGtw7JzuppiKnx2pw+1dxt/xtWWHfUL2wYK7vuB63pH7ZDP3G3cEMlilFXnY0w
qdgQbtnCPXAf6OV8dl5KnwULKN5m+U/oXTNEV1UssaYqTGcDxwWzmD7o2tbh1Dt1
Rtt264b+OjN2xCO4+cpmhVUoty6Me6XaA+Le4jQ8UWzjEdDIGn2WhPNQdwkt00tJ
n9H8SkovnylTMbEa/MaoKg6r2qv+0V/Y0d6WOQu2OIbRilegBBK1HLCHU0zG/eRZ
s/dpNzQVVDPXL/BmRaApVAKi1teoD1aa0WNe0m+q+jt1vz6nmc1y8dN14fxYeFPj
OmSGgJBuySaKeY78yQbHfF9ZbJyxz/jt50755lo8R3SX1zsU1Ci/pZm6X+4md/jn
o4jN7+751nifufO3NyHkoHHYcuO16LRw8kf6FdnGmQfVJDWifytqPn1aiZ1vE6RZ
wkNZ71rMJy32cLjnsR/oKNSHeBDHBQLGrbcgNBN2ILicDb86Wd5ZUglbkN1f5HTR
qsELQmFUzJqJPGQvq1lHMVU/4/JFTLJBTRRDkqGgHoQ5rVQQJznd2RqYzRSyb7Zo
Yn4O9kAtUDmr+vL5QwtyUECTbLkRsrYru8tgj8O0eWTSJWl/xnGnY1oJ36LQ7QE2
ypm49kWP/g23EJdxGjFy+k7XnKA4nndT6AYQAmAw+WjOYIjcwpinpb8Waa/FUdNM
dUW1yU7u+TZ46cedC4NTQSX5HRKumpjiwn2FBeZd2ht2It5NqDhE5ICYP6Zlvzgn
NCDlqHF3lhJNPyGRnQrUcwHt9SAI/RXiBBMZWDstiGg1yCj6Rk5Us4865HKEuInR
3TteMTsDo//cZ7DuJx8KsMSskgqiJGPkS9luV1845WV7f1HkJWMd+6OE1BXoT0eA
6eUr15Yy94DZVLFKqPnfzB3h2EkR3tlLlT8GQWiZxWEUMw91zNk+g90+tfjUAVAL
7+xfdGOKft711aafai2C/aeqhqQM37vqS62gg3oRiH1ZFi3lLKXyo/nxEi+n05kq
iiyW+u8S/qjHoJ5b0yc8gOB/Js8uYQnoGyZD1KxoU/p3fm0hEbzwP29sDdxa07Jn
FbmMEhtHa55y5sJoZAngIsOSjrkZOSrnt0IIAVBFMsQFJs8If9q2U2TzbxsizbEj
QiP8zFnqPbr1vaR950Xov76v6/Swi4MsVuCuUu133FYQ3YAR8h/igMPhHToDZlc0
9GzmINhgHLG9VeuDITns04u8x1GcNNYm31Mx8oWg5aQkuKDTHcpTLqYMQ0CjPw2b
dBLm3jghlJ/1ijx4lTr5wqZmCpA2aHd3cajuRd7zLorzdWzLl22G0I4TglVAGz53
A3XUS78lxoqXvOK/Ab9aAUs8P7aCDtuAz7tliQJw1Jud2osLQmmKcumW5u7MjsT8
aAcmwYc38MX9NW8bE2XoDbA3VZo0vrzyAa7PDd4Bq4bz7PjodX0CPIu+SVQJTG32
sFGDBt0XytEaV5fqaeIpZ2xYwm6/QKDs1ERuEjs3CgIvU5pA0/zKnQxHsOoFDU92
s1p0/BmSaszLXoGNyHaT4Zehm2irUj69ym12A8eiQDerqsqxf7tzEquqm8ax4mTZ
t/DoAYCwkrwC/IyHApyBEvBpf337Ndx8oBXiqcZ+SFumz5t42UYD/PfutbZXeSZW
l5J0lEbEO2zxz/iEdWHxiZ/0pNBd1LS2E/8IuVfRzd7p8AA/uScAPWlWFNHGuRIE
9ZiSvmHiKHg7yWjguWOIn+MkZTMX7UOzLA0TKgKkYd2TJmeDu0pY6J4ogWDflcAi
IWjTjffJQ0XoOdyKPf7on+QZ2g6HBuq2m7wPaVQhAHoADFYHngU2Gtv7XU0cSMuV
0cHJRwA/x8SkrL2W9n676VB0sIuZVrvcPTVGk6md7njEt1UpP0iBeRYBIwmeebSH
EzoT3kwyaKdn2LVcHusJWVpu4Y6MwhAsvyQn/Xsw3EtlcLwrReylgZo1pjy8C9FW
Y9XJoOFspas0+BywLaK25QD7QT44tCedsOqVv0DFuy4yDeI4/WckVbVYLVDB2w0n
vgRFoIRzuIUJ29eo5BNd5ETSYna6/1JhFpC3BLGOcjbCqbTsFOqsG43oDqi296yV
Qf+M0XvYi1/AmQukrqHXfhvuZh6n0fWLr4Vti4HwS8DwXagNzNZ0hDAymKm5oX7x
LWz0Lhbcl3wzOzAEzbVNZsErQjBwgPaUDmHmRCXdtvEGslHFXYM/B70CgFC3wsrC
QP7/0N3sw8BMDmD3PaOQgu5r0Xk6LfUo2V4zLHEKOwnlmuLcRHINnwQx3CePsx/d
crzep2PxtGEHoHlHjhkVKXFt7XBiOpJ50oKuBurm0mIUZgLJDWsZsHmGCUCQd8tb
dLOkrTuiEeztVqWwKvtBNhpDBqM2MZutfMYtN6x+DMGm5j2astF4hBJEpS7sX2xb
bMIGyjayxpeYcAm+HwnbtKDmi9nexp6iguhtrrFL5qkfyxwv8WB6lZNccBxUhZny
l0Gxj5gDN92k8JxY6aOc675vibNslMYpQj80P2qry4jYbMUBW1aMQ5cD+uxiYuc3
LxUyDBWjvEKzipIxAkWiVXfY675Q7zZYt02BEVwPczp6uDGYAnRoZE5tQ5CthOON
7HHNXdk+wYN+uFs999WDHaJEXTCAN+IDdTRPHauoLGt2eMYhs7t/Nr2g3UM0MPqL
+Jd5GPtb0R7Awr7nYyNLm4JKA+69ADEMkl7NYkHjgFwU62JptM3uJTIY6G3coYiX
0p2jE6XQlT6IFfpbb5C1RSHMFeHYbjj4uBaMRq4LgnIyTzb9HcN/gml+qh2j71jI
odw/o6DjgUrHuslUcvYgO6qtj10jJ7EHSZFj5m5i2Vu7uFF1eUpILvSXYFFU1uiG
pw06wmXU0GBf87M0BVR+K0fyrFdIqJYcPZbrccs6kF0YKcLCzDXAcUNMdZTIdPeL
dvM6Y8hhjpCdTrkJxSlAdIGUp8XBBU6jNxmXbg1z1Yni4gBBTGyFjBCYaDWD3QrQ
7aduA8mjay9Ci0DOBlNDFE8uEPWvOvHVAk345wBTrupJ1YJcLUMSKj2FD1cqWhnG
pEOmQRyHul91uuCnk/pk0j2fmG4T5ogQod8OYaeS06q7sKAASgSvOKHGygRwGnCM
w66ONnqRNt5uSUrM9hxW/oeEiCB33al8RUkzbMyaRQLfev1iK5GUpK7rpdobcFLg
9ZSe65Y3vQ+UfiJK+8+OG+zsm0muRCxstJpPX+7mxiA6nb6mOna4lw3TJQGcnzrm
fwFNfATuJd9tnbMxR+kCNUv4kQuRjVjuFau+RNRrbrEuWhYtVoSILjIdl+RxS+95
JGWcpAwjpIr2qK6UJyj0M/AsIapzF41+b0+8tshCpfpA4KM1h/o0xcFTn0qGAcAK
pp3G5ZCnGyHBbciNHMSAF2iqNcvcruYqYyxA0OKFUeJxPHEkVVz+mN3jS+nbIkd+
Jp/AbA7t+J9pV56etbtYwAQMhvIYtJ4qdrWbfQXNRBeLdPqa4hIvGrJD6rcCMNwL
FcLUxLfVceSeDUJ7ZynBjmw+WEe/A+y+r8C8CK5RkxX8o7nR5ax2onWIIrwRs3Hi
Kb4n+UaHQ5kWlawilJbXwEBNWVBYAe7W5hP2PU5/JQszOnLhO61f1fEKELN8wo3H
tIpgiHV3mFXUG8yteiMV6WZkKmH3ErhK5dfxOofilQGds8BNRHaC2Z78QUhlZDCc
ZqHWlDrDdJvDl62B4m2EalJLcKUaVQBi2tYyy969WdFLF/OR3sZQoRFQWNGSscCX
o7dvAQIXuEV5HeHOxIl3lFGNr61F9dPNH71MjvDZs/r3eCUUKyXqeQH9DdeHO/7p
ELJ1DJKq6/Jw/80/x4LeJ/30hmUZE0orbg+steUOOPFAjIniAPmMZoCday+4toSK
RQGjPaTm7IPlIQ+oYqu3qgbziM3SMIhVcZmrJibJdQOoB8GO+wuhS5wgL5XIG93X
kdHeEhSjEyrUjGfW9+MJrbc0najkSJgJrFWApR4vpmng/c+q8nFoL7s63DKCqkq+
A0rLLBZteAZwtbDiyo5PjyrXbf7O0EZkKijj3V6jDsTMDd81uUfa/2aUwDo/uNbZ
9O88rQl2uIuPB0H4d9dLO2rF0mkAzrEIsA0lWvvvCcV/1IQOVXcWLiiHdQNyDCHg
ZVKy4mukzjESQvhrzzQLjbk/HdkwvXZgEQ1fedEKaqpPsTo1RxR9C5F6KePR93Kx
F6TS1wJlb5rXFw1SnAz1NmXzp6gtWP/+2dBO84jiwqsWQ62Rl/xk616NmgD2MwZ9
fB4uv5SHDM2uX73CuSK1ISIBySsW/PTHZs4CAT1h1fJz3R/7S702+OZKerjoyVHN
6diPMJ6hmytWAqeplq1cWhgDWbBrtdOb6Z3Zs8qfF4/6u3k5QMlVNClQtQ4QmM1c
XFrr4ju9qyuTsPp17ekctUfVyWxjy2WqlIY5AUnscdXQKSaxXNgK17Ty6CMZiZSm
nub5Em/QNT8O2c3Ar3dbjHN473Lg5pQFIXkrvVUSsk10BNIAdwNmtMZGEbVlZ65t
xXm0sDq9h4+TGGv9RnTJhbOYRsHaltDA4+rReSBM67vhEQEKKUEHhrE39hPnBlAY
RYjtTiTrRj7nMgYdbQJy4++Phw6gJ/EGVteQaLY6gv/06Y+QqEK/0EfwnBILl8nh
BWN7ZvAc/ZPv/FbCJ81oCS9ve/LZBGn9h1ch0WcMceDlPkhM+kmFoOPbuEz/fHje
CvObAO0cBywkxOFMeFx5XQkHMncEZ0Y/SLXOpklSMjDGG4B4PSi6cPzERdUd8Edd
y3EQY2MejWI8M7IOBavy66iAPhiOAS5iak4TjV+gjyYOAWwaDbA57zLBvAa2diSt
GVuH7brzYsxCr1nx1J3mI8u+X23C4LZwZQRU7HpVFDnJ2Jb61jVCJuuOy3xwrpcb
jAUF9xAdDaIPwzNwGf2MPN8Ech8BfA8/apGEcAY1xIwWDyndBIpgGIcp8sbPbFo+
kugK6Z8ajnozXS8zs+LpfLCtwjra6L7YfNX+pF6Pkk1jFRi8G0GbAGMXebqxQ64Q
MBu6WMljb9g121RY8f/CqVJz0ay1zMgjp+xlwifRbIZW2t/fPxnP3dIL3Hr8u527
Gq2O5M+vqhZwM664S0WCDOfekWCjoeODLZ2EQagIRA2zl2sXVMSqc3Pa2i21AmpY
eWHExHK8kT+EhbtsCrQa0eDeT8bOWR54WlLv4pRGXd6zW2hhxd4yYX8Wo4iD5wEI
eupFt2m0ZfBzeFWkV1XR3Wcw8gQCulZra2ukwQx4aPYrDHLcsel88XXV/DR2Jm6C
ndZ/x81uTOUYBJdlnYkAjMmuaTq2iAfnB4LeKUWEPABEpkYxHYzxI2TVan85OhSD
Mqoz2acZNSQCYThx5gyfqGn32P76f8yK3/ivqSBIJrkF7N6L8MhOeEZMYqoaFCkY
lDk4ZxRk53YQaCMWKi77JoBJNVBPY7gbc1a6eRaDdBgkKx6+MLkTi9zIcuswVSCb
OvIZuOOLRrEjmbC+cqw6Wvf/9csF2QEyCxgF1089qqB25HXr17tbtlIhuC7IBxZx
lg0d9oyPx6F/2v0afwlzKChwgEQaZcA/8t1EZIBscrrlCT9hasABI979/PJSRa8P
1atfbvu48Ih7Hngq/2iqpoUd6m65APRI+xJ3igMthlZbuLMTGBTgSuJ+cYLvqxnt
Q5gmt6k4Tgy/s2zeasscLIA1YufPVbWCtERPDiUUiowBHXoB4GOlzknQG+QJ++dL
lWIKgHtYRQ/XO8l6oMRFqujv6s7pLgCULN0c0hDvxUfi3F4U60fCDPsMxfcSl9zR
njND78ifU5Hkxdp3hipUyTfAHC1rPlEbLyyNYReSNeJbsQVxWvFdamX7DLMvxPiL
38OJsJADmh4k6QTA0X7AaI6X9ghs4a0SzY42YtwHodA0ANlLVKL7s2HWrhUew8oC
tykgEFZUrlXZE9by0Gn53WCnnqKpxHiHl0SqcaWbAzuK4gjD8A+1tpc63D+NHQAa
GowNaxhKMV05cWOP0SHYI129ymhh2eQ9u5SEOaoz2jJHMudpG6nlGvtE25VTz8LB
wTyU7DvcPOkjh0WFsl/pwLINt56rV5G37XHVNPVJLfOzHNM9yBz2TMuN+Q9+/wcp
uJAIk6XeUHLL8JbNToxAGETZgKqNvcP4SSpyEYZCY1ekoqI0jqNqOvdLURA+GmqI
OeZBJkvBr2FAyXwnAV1nQ27bQgBHBVbQFIKaJawy+J/4KrxrDTlw9hx9HwejfM9n
e/2KvmgAzVHwZA3eK3nipEhMiAuZ5GUl4vcGZxwFGzrhrCZlWl4dgNU9vN8imV3/
VRz/DnC1EtxYrnBIKyoLE6R0oz35TiPCeNyqT9AdIpyV2Ifd6EB/Uu5V9TlKKSMx
WcdrL7fxWWBaVv0auLegaOt+7NBgVgg/deYjnyjn8L/qcj07CcV+9vHMkC9Hdeth
UwYl27WC77MPEQx2p/RVxItayDudUy1j28f2omQ1HWk3sac+dX1/5WArwNunVtZl
TC7oX9q9DTZxZTzgZP25SPEf/6U9mYYAJ1q1N6MJ4M5n32XMB0qxz8ERAz7UpGuF
wb6NlTjz+yQYPF2Lqp+rQkeVvToyECwkR5xpx5DKmlp+nSOwqSdCUy3kDiMNexFq
nt4vZAUmL9qxQeDgIOClwcts5G4ND6t3IWzixpstaksJkiSpQ9YPda5AxWzYATJ/
gKnAaJbkZGIrdajPjgYxQzGNO6RXWjaQY03BReaRVhJjHRE2C/vkOMX/CFqxm1y6
OOyYgcjV8jvs+kO6QZQxc7kXrAoFAxHjus/rR6Oe3Roawk2TCHnAtXBYClL4SJ9K
A3JpOOtn3kf5XliQzETEJBxH2CuBW1wabc8yzXh00TuzzrGst+EL7AONYV0it1xV
bQ/tL2PjpfdpUv0LI3cxt5TZ3D424Kbt1tRIuB2JPsw2CW6ZvyuCB+CbrUvucGEh
1v0jnVzeJhE1UKA0BfozFlXX4jRH9TUBKxNGrV+YtXbMCUJbrL7GuzX/mlLbQolR
vNTs8Fm3+vbZDG28J75sQBgwjpM0tg9XDY8GJP/ZmQwRb74eY30OBKORFsyiBJ1O
w8EQHuJ3uVpSZq++8zm2javfzbKHBRRF+2gPprTf02XYwVls0FbbACPseafjlbAx
bE/OHDUc04selzy0T+IBDJi3SuKi2enEl14hay+kE0w04KLgHLKQNC4Qma2bYV7S
8JNvYxshMdi/2WK9zF8KUC68p7z82TViGXk+vhx00dcuGb/y9S5JX0/VeW9Sig19
7eySXQxWcKK543/zm6SXvM+Tf/pF8TiZ9ctODcT+iTqTG5fgINP8o6EKExnY2REs
0vpybiCsnaZadeygqcTzdDN538U60Y/jHeSfh98WuDRXLzGV5C8Zbd0ZVE4XWtYF
vpNooF9rsH+oKQdvbyxIOwBV8jO6VgFG+B8xPyuAdxkQI7jGfi0CH6OiPAZoEZyg
S8X1y+fIYwvSQtphtTz6sxLNvH/GAVGIkvfl0sIVPRmmnf9ikqHx3eMuN786+PJa
GZuUU9EF8Tx4HBRyQmq6tzHt2NjCsji72QVpTAsyqF7+mdiZRWonJoXHI7dsHSsw
Wtkw+LvXfHH5Y1gMGeD2loAUb6egXE8TPbjkeQ6jQkYQFTNR8CBaVDaT83gh+jj+
sNW986wGWsgbLRAATWvyn2KKHPe8M1RB027qOB8H8IzQHl62hrSiv0TsEYrVcM3e
weRkjaJtboyCMQDt9DDIVKJ1fmLQND31P27xd9kH84D8gjtYuCjVVp+IWrTjfnWG
nSKx9P0vYcjolN6JFdf1yP/vYtCYpop7kEOlBzvNbcqeu8BwyCqpgDzkQpmjO5zz
l7NMepPwrnvNizHfPGRp2ISzGkc0DGCGO5A869G/1xbAxMA023zbstQB6V8G8X/z
NFuKqN+GDaNRoJln0/4VBqk8TupSAfoe0muS6zBA0qd/OSvybhRcpcyOn9vEzRoi
bS9oo+6JXzhOLUmfSE5n2Wv63/xkS8/9f1OZCVkyzFZqJZT1wM/jnirr4134xLwt
RK7GPDZxW5w3Io5itMcfExi56B3Xj3mOIt87hxV0L+h54WQsmKy1oadHG+QLqoET
mUmSzsL/VXPbHYjqEXNP3mXs5YtfBUPKs5a1JLOyp0n3viWRSRAf65xnEmX6V+pK
/DdhBv4ZgQ/oC579sLVNhzZwqAt99/qwNbf0WYkNFkO6b1+ZiWI1NDRTVaYKtssB
A7faHCevdxdIZ90ViJe+t35pgg92xAGCPb+fn2gZ1hE2ytr9NtfsyHzf2T+m5/PK
qIaZgm1UoO6du1RjjwUyFdib0/TKhLNG5HAMQxx+2cYvR5dredMtqUxawSdOaLx5
mYi5kaPCyBXLUQUeEFadVwFX6ZMd53tHLepSGRSbJ48TMcKn7cuTq+HHT7LcLlm4
w7tn8sUTwRGgR9e85/nkPKClZTwYYIzrv5KVQp0IQ5RVh1A9N7ScXfWXE+Uvye9G
i/vWqJIHJj6SgILwIKYlWKA2G4vObVoLd1U4v832Lk7jhH8jJ26yvVySowIAxh81
onb4UpQZj2r25S9jzQ3jlHGc/fYkDmdakKDQvoRKEsdfz5tuRdd+mhW3sUpdEesg
WYCDUZMVSsWRisOBmE2M7UbMCrf1Q4B522cxfl5xXeHKoPWSizbKmJfGHQLQkvt1
kEsI/4A9FsPzWEyfvl5f7Io7U5fsd6tRegO1ykoXEugo8DySigHtYOZnPVGZGN0p
//PW51niBwaKbUh/rfwJo+ca/bUYH1i2Dts1NZDtbtRaJsHLtUhWmomgf5Q1rzbp
jqPiaOZeL3raWUwBHefNM0dyILHt57+wPMPyz/5j6Gm0vuSHs03RJ5rwohDtToZr
jBJt8COUuo3RKro8uVY1H93JO41QbM2Qs6INRmrmD8i+kE64BmNbwMPHSF4CT37x
g3+2jFoziQZHwOM5KEkDbssfwf6bkiiCakY+mUXJeiCnfHa+2Mhqb3aThzNvTte/
ssGZveOU5h8RVEe1HFSpwtsLlLFIGeIYkC7qVp0+ibrS0amMcyZhC+CNe5+jJKVM
fuaaCVAplzTVNAy7zDRXUDBo9QG/pX83eO8nDpNk6ZdC3zT5HliNVLjhR4ODQIrw
rzXDA0WVeSUCkuSZtxX6OI3NZ66D0sqi9X+sPWKPiX4WGCAFdmYuWBi7DEEDw5jk
kG5mHWX42bktmnyI2doaKhHLpEmxULW0mov+nFTmCfi3jD/F6Es/kMeO4tBuGszp
2JG8Vo2hwochgYB4BxxJZdVrwY6tQjF56BrmWdk/jP/4ttAG0sy35amt3eCiEvQh
2IvrRvPm9ZnGQL+vaR/1PemgJOYzf5NqRFyN1FV8LGnaTnk9u00gVmdNZyqH3ZRC
fuu6Zp9jP476wvsHkCE00RW6ttCLnEejYkf9gca17aW8yAtz9+gnkxjSA9UlXMHW
Bokz+tXovJr/1jmBA5aCexh1te1l6qC2nSeuWwovpoa2SB6lpvZN1//wqH1H6Fdo
ZYcQ/ZmTqGu7lRPKHXF+76g8tr6ceEF98Hdh66b0O3EsbrKXoZeD8pr099rEHNsP
B/yfuNMl5tshQ2ah5TSyqGm2nLRduihiZf+EzxwRvXHZS8GrrwyqbEM1uXeIcoIZ
dHV+fkfZgvwH77dsceC/XI8eTYkDWAZkrEEpAQzfvtpAVzWAfcky4mbM2yZZN4dv
yL/HEjw+al/AHAx7ZfvcAvcy28YloqBqv1HduDG7/opqEzpEsiuqwOb+wg3EJODD
apVderZra75TDNnleCehWdsNh3z4cxeIaBrZfFcuwqeD3B+jZTNpsVbaqVrI66bv
Uu20JvwlIacOwqfSCUWJGDt1FW5Y2BbM0YNg/TG0yMI28vQgvDsZzoCan+4X4Gdh
6aMDviJqynkdt9sE5Y/sVPrzfEgFpmx23Zlu58lrxa9tXv70l3AlSKu7/1vlM+SF
Qee6pUa0nc5HYjqb8t+iZY0Enx/lgjxJOTpMNH4eB0aabcUtRG28u3GpGEykDz8q
uxieERmIlt9t2w7ooc3BPK6Nb+erH/Xb2zee20vTn/O7VDKRbiSN8VuLy7xG7erD
u9FyL5kI7jSCIZ66KREYut1b3MjCTLfxY6IzZ5hVoyT0R6PpcdkSoVKTptFPOkbb
EoIqCO9WkBnKCOBsilUhXlAco0tx6uKNzFTs5VTqt8jXTCKVBdxugD40h8dWdfZi
ffbI9/S4pVm8rxhEFB4oKYNBpTHvvqCtY2pMyhE655V3iJ48Y3UGwI7hjH/YkwG9
dbgAw8fdLvSK0jAAubHpV7tofFryQr/w1YgTqQ07TOcFwUdRMVIu0OC+pPgduQu+
5qiMDSKsHN9Vn62e+kzdkfdc2q+lFv/Cn7PGjt0U+xxVunNMc4e28btn4c2fD4lY
cuxYmg5FqFllOprZsoGBd0Rw1KzNPvDR0EDlnDirFaUgFLmDvxzCrIrjJ0roc34p
HEmB0n1/TfOSHcskXh/9LHWoO3rG96PLuZSCyWF39RpePNvPlMTyJJ8tAF9DdQ+j
VuSaVP77chc4Dy+kH9G7KGE3cV1DBNFCQp5DfGjpML5IdQwCppgFXjFvKdSdbbRH
BkPxNbrZjmaDafGPgmLGkCZ1ioc1tdngx7ye/Uwghj/XAIk4l5bBTvCTaHUHjYqv
uISsxzTUP9eKIrL0vq+/sZOy2dkL/ADqCJD3RjnKcrG29KGU3xuwCw0r2vR0EA+/
wu9EFbQ6gwiHELqB5pwGkOj/3oPDqavM1gC5rmXLGJZENlmoZodMGfV+CXcSBbfX
kiZGVgr+UMgJ9o50db6k57ut3zqr5cBn/77hWCAYBWnXEJ8vnuL83yN1xtZTpnFf
tcWcm2DCt9j3DoEwqS1ZxOKw4p3FSuECVrH5yvfbpanjawj776q9Hq8iEPoXFGUQ
qN4UlLH5x8foaAGFkbRdgo/tQzH1NgeSMW2F6n5amhvLirQ6dDpMHzoHSzpEmQcx
7sTN3B5ZZ8IHuUiFVswTwS2V/FcOFy74DzpB4q3VeECLBvPoJ8hKUJZgCuWlMj8u
q7ik4W2p8cLLkeWSYLa2USUIPKzv7TO9sa1MUfhGOcZmgPO+BaszcgfftpWR5vkN
2uyy719Oi1JfI7UC8DS0EMv/dl9Aj5QpjxSzGx/OVC7CMRXZZz1vqEV1IiPQbAAX
1lKsLZVbaqr/AvncGx9/DtLUnidcqHKxVdCZ+EuqEhIBbT/HS2h67jE45rn+Z0iV
b+/u/ptukCphM+5YjTFCxUM3Lf/513qjnot1eHEUDceWD8lbkWopdSwgyxbMC3FA
uNl1xpugBGRLMxv8f/SD2g4loIYWdBv5PM29Ju+EAaHGaiFuIRjnePQQq5G4+zA3
2CfrzHHzML+UituMkvuJfq68hM7m5MeHbcf5DtjnTyuWxOBlLUdoB4R7/0BdEhp8
KSRXAX2EX4z1jcs01RuIDONELCXuZmXcwxJjEXjE5/jxAj7yZQtHP/fmXTjOwN1x
e8aJI+Qogzqz2KPcRRX69gtAAQ+kb49U82bgPOmY7OqbxLNszcEWoarwPbdsSBCp
0m+b5dRuX4Ca6GuShmZHYj30Jdj+liNx5CSFKEibO6hPUWxS/Rssv2D1lMMWphUE
OWj3Jpi69JGGwOfbnaPvVfbs97JueCC4z5KPbKrTyos3S478920EIVLoP4KwJA8B
JUnaCdQ+noByJLZivvIbJ75c73IG56UfYke5lFK59PtTzsiecTVIDLRt3NKKhPdb
yZzkB7rzn90p5GzaFONcgZAQeSFYw7fdasN2h9W9nr554yMZVM5RvgTMLcCvKnNV
qLAlJV8rdGBIjVm7jYVcQAxIgmjnpDC4UJ7oAsqJiDZ338KXtoWpR2MHKPHNzWh0
ftgyuhHcrp+oeVo9oGJA7J+6rR9nv6atjiACr+j4kqutvQGgzZKmArObYNH+94Xr
FxQL6F+QWGp3itMtkaaBdkwJ70q4RteUMQzkkh2ejH87bruxII8TY8s/GsTtd9yh
N29BW/y6ZxC8UV7tzvxGkpwZSgis6/lMIcmr0xynkIu4N/X/Pttd/1o6o7eIPA7C
zPiihcH9MieI1ipEtLzMZ1U3AZQJjxD4RAAJf//FoyvuBn3crn3UQU8uZ198veuv
mtkuESanU4znBJsCEOGmUCwTdOuJOHlejqDgurY+9vGDjSKSs52agVKvLAxlyRlJ
GUM1TQQToWeCOMrUqpTAxD2Iptka0KCRQFjAts89C7XetdC1D9U0bpQj5WYrD5l4
51Fi4xa6vb9i0B2kltyc28H7IhjD+RdtzoLzs2O8OA1evYzINpWr3r8ZrzLkS0EI
KkxRPUnIitxD0PEggOZVVSskmuifI6d3urEuFFO9EvJyWZXlUVJaUQLVDkg1YN3T
ednOMeg8q3bloZGvwEry+S+0JrdRv1qS381pVht/unkHUmDvBXg6PHzdeci3B+ZJ
iLxWS7pyGwavwgIRuHnTmBKB/Ii51geBJXaFiUI+GmBGXGOhddb3AmcaKmwv7jpJ
phharqE8ay455FjKPKhca883CssTr7GL6KuAaalxTnujh9RAMzzVnwltu/CZwF3Y
pByLmGfN3I3NiSJyqiwPMD3D2chzqcoicUq2QjqD+daPB5ZrkpMcWDunQcc4Qb1Y
1vLqCTbTueV9AsPSW3e4urapd4WqBsnxVmi3XSJXloh5HXVWPwZ6msjyKIGK2u/b
h/zh4mfE/XBy9e/0UG8Crt7T22h9GBu+yszIF8voI0IooKrfIlRJgqe87F0g3yE1
vUm6160XCU2qoKz8kAN5tearW/bq+H8JYYjRR8jczRDf8l4ZOOkgEsonQACNZMsA
4FEiDJ0TKs+jnaQUXb1YROMKD/pH1tQ/MtRtxzTOFqPLq7vV9w+j/yC6aUdRZa8x
d0NNoUbfm+O/oC1SR6Vwoh5tHstTyl3zJVRCBYDfssSpsXy3aThdU849SxDUF0Ai
6so4DXp7ZpKpplXRjNSgKXi8ERnFABM6zkpS2UdRiKgRv0wAk5om9Wa72gFw6jmU
DYRLvFvUQyqrxnpwdEkym7lyWMNelC/yZrnn9HmybAKilIRqsj+ssD8ASOkMtlnH
YPlcHZFkGZtcat1ACI9T3vRH7Dt62EAamzjfi00pknRoA6rk1Yr6G5xx3eyz+GSR
yH4orJRKgvsORoIFpFw6nP7O9bbVzoXcI9TNIFGwLacrzXpLfyI/2YTyzKorQxQW
MOS7tHItVAZbnbP32XXMV4zfwP10CVrMTC4Rxf1dHx2kOPAjqzCeeeqNviVZ0l2N
JMEmMOOlyY/BZSY9pj+e2+qDyiSajj7aTez1upAbsesu2yhvfhCdFSdiXfTXXI8Y
J+atYeYXysj1QQlqGvlMgIjGR0yVSzE97XKj1cuYqrlqRDDYP/vaww7bUeeW85Oe
ukAsqUlGTuAR7OawdzxwxnPz65QOhnNwkwHKjNym8b1qRFlHO7Y8zi+d92m7XHkl
3m5yhlXS3+8u4sT2Y0F93Y7s0Bp5OyhnbBycDNp1DoUyBh/4oBlsFVdjo3xjsRV2
Pw63A25OImGX3dbIZkkTuHwx2Mlb9+hQZfIANRdyEeKQNeNKzl+DNmeB0amHhS5l
iR/8ldwzRROS+SpnRevyQzaWjJt+XDUUbqqgvhmJn10DwS5FiH/H79PZIErWAVEr
vGfsuchrcKq3GcdS4AZx4RBjLH53dl8mrmKXwaKyiFbIPmWTMjBK6kI9hmWuMNEB
05HQBK6y86jd3zOk9LPYvRuL+V3kX3hrkbCKxWEIyYzgUCKB9zKiNUOtSk1JA58D
mWJHWcD4GGKeIB3bARN8/rwCDkKnb/Fy2DsOEtabsYaa/TjCpUOeOmVU8bR41bH4
cfk95ogsFug12PPbTTBqszuV5AwTdYqAgPqEtGjUGPZW63emUj+q4FxAsR2/8mxH
hRlIKL+VUDDKvLsfRM00mHB/7YY2tU3D2Gq2FMkavU0BwV3+4IMrknqynMNwRCng
IEZNKnNgG9DpYDjiLosAyfutjd0eHUgkdiyYNv+eaa1KuYCXDqcyp62QjH6cHVy3
FYyt3pkBnsUZJbbQz2T1XRaaCiBUcKjjjaBZQsofx+nU+WP3J6M8wKetW8z8XUZs
opm71Pwn1NMxih8y6BcKYyG+Tc7PVgC1WOThdAbTVkMhyqofGtedMbL9AHpvZm9E
YTvVQsUgpAIMa/ov3QgUA5CjZQUhme0J+K7AamMp8cOYkt9LE99CI+63VHkB7mC7
ynfdVlLLl4qvg7mcM/NOcHKVJjE1OiM7kvCPi3yNyTFmNHGI2mEsPaYe+gIWT6aI
kWBy9GJLSYtpZPKTwfb/omSV9oRh4PchXfCOxx+dYYHBwc5bplwspRS1lNIqWkz8
JwTi9BfIxrgzY6OZOLDrF5vYnluNo+AZV0iHYyJGHv+o5ekShYtPa0A3/pxHoo8H
fjhSEJ5A41/DErBI2HmOLDnSA3a/29gr6SPB69swB/YXKN0d65gru+aGdSY0Otr7
wfuCq4Juv7kB+f6dAUgX/zJcDt30Fqa/yapUXLMuNU+cnCzT3Xiz361qp1iCPKWq
Rff3nmMPOOIdRFrWff/ncFBZ410h8s/jJum1VqdVkMyG6gSGsB9guUP5r5ufrp0+
R5Xao3qKA4sb+a5Jgfm4/L53ufjpP8+7+55fadCtV87Kv4ZKG5ToGXg2jj/eCuJ4
kxQlHGa10BDyLTlnvR17pOQiUN0IcSR2W9fOoSqvBfptn9CXHyySAriK8lv0Kd/s
PYHlj0Npq/t0KKbHfK21nduab3TNWRwludt1iexWnZ2OEnQTvCgAARf/xEXIPAwJ
rvMrRFsWdE6sjJY9Hu40CwnYTqKEI07jqI9iJNNpOf6hqRBgHd6oBi40js/lFXD8
nny5NmqzbUbeuOF1MIDfDjCKmwmw1r1mJ6moxyM/AP93R0O20SpyWsmuS8R0Mc2P
Z5rC4ujiDVv87v21fRChKhH6Vus1LkYlluSatWYiq1GWy15aQpUeOFd6W3DHNKHt
5HYCsPx+P/g9WU8wdvdgBod8hWtgUJH9KF7+k6oqCIeivXMBpYfaE1EfntQRc15v
FCjacysQo42MbmABtFhdyDp0NmskIpjL8Slnebi3Rmxe3V6IwweEfr8jwQjI3gWt
gKpGsnugXwNUF1QFEpUuRSS8ssZUX7E9Keh5doXYtxSMCLwatfE7rfvOvi4ER33J
aRmhTH/Vwve6ywv9zklDyr/XmjMKFUckMQu2Qw+ktbsU9eYFneGPedBzmtR9Ohow
2lg+ueY9MCF5axKxMRSSyiokGB9cPCG3PN6KOTjFEtmuar1Sv9VcMGAJSDlysuuQ
c5DDhj+ta7liX+CzduasCqOPBXofdJyyCl7a9vN319kAZ+Vw4ta5eODHDZflFU1T
ruT/MLE3sfIsk6OP8c31PIOG2mWF6LwkfqatZ2eO81Jb6su2xvntIq72LM9bev3Z
LkyYrC4jb64XHvSTDh478jI6D5oo2xNUnS7zQ0n/Bix9cEEPvp43ooIvgFrpe60Z
YFNNVydFaZuinN3z9tRm9JUMoj758ewk2FiSc6Wl0O5Ux/Cwa2c8EUBt+wLAs5h2
q50XrcrsCnKgxLuWV1wMrX18xeI5uQvZwWXz7cIyI0WsumsjYvLp4NkKpGiv2UOn
8hP0wnZNNR5NKZUeVHHSgN8lFL0s0tkaQKMFTTuIYu24wu4cW+jYHfr+NyudX/8V
3P+Tgn540IcPCurhnfy7qKpq1sL91iWBAOpgWun6utTcI6cVObtKBAgOueTcmuwa
VRU2Lj5bjzjuLqw7YKS8EibH6JT+LKGNxmRzvrDxZ6ysTMvq7BXWdrenOPX6NtBS
JYdPtN3djpZBJtuQO0I1/+JbH8CO8mWFwqxPUulRPvtS7kdwqMSPtaVhFmp+rpeC
dwTPBS8z+qTQ9pj/0R42m4zYRwmR7KDwXf0iXf2KzYBc3mTL6C7u5jHBQFaC4kpG
Umh0cLQymZqFj10jCaGKG28jruBFXr4fjo0NcJq9Ljrlk8omNmLDZWFzVWjnWldi
T3NnsKq0HdLshDFLLruln05xNSfiuAxQVe8ZN0EDqeGtmYwYJRtts+83jR0WZtsZ
CSTMXOrpYFKlvRFrRqiRjV6Y/q2F5bHral+ibkJGWjHWaajr4+Aye+/eiqonIXwD
y//IP/jdOFysBN3838u4SsDOgkyFu0zzzhCpFg5vf7PTJtxi6GExqtNGvjfFN4P1
Pd0xXntZgY/TA9X+bRh0G8bZJrwtRJERSy0kekV+LSM9G7GCu1JdFYdz6IqpGjM1
J7oT3NL8gesS0FhpqZ/NUcOn+hpGjVDPjgdhkCsOZ69V4AlCTWPIWJNR3FsUkDSB
/vTn81hPsK8M+grvfocdwtemFjE0a0NNoHr+XrimSFWGL84TysoCGHPueBzyd9vS
Q2dXQxf/1fholvONbUSeXUY0AlvOeT/tS5AZFuU60p7du+nroGfkHF7ldVP4qObQ
ie1oND70SlWhZ267XNVTmbNYf+b98PwvA1CM4T2rMbEwZMUptaNvBDzO8rYVBV4E
z3BtVA3ZNJ4tPSHTNnetGdIik8n3bWtQb90hLUmdDRkv3CuAcPqBUCgBd3OCnbO1
mVGH0Lo77UDZsotct9BjWMCa8oVkox89GP/m56NWBfrtHc7ROe/gtsYE2vuDO7yV
bR3OT2D5vNjXGgqVBc9JMfkq1qNVDKbnGq58a0w+9owXsH9MHMJaVRAQacP4w4mH
TZ1I2OjTS8/yKcIaVpCBZMp4RP5SG4he2v+Gi5m97zHMnSgFCI8ItA5vjr0u4vlH
kGwEcXzqYWvq/xU36cUFOfMNVE2gTDeR25nQSqXCJ+55qemb01Uajs/kVjg6OwnF
2mXdlTQwEu4XhcreP4iqcIatNrhRCgBN7yD/SBPWrnyGGB1NBJc8yj0bfy0YDIQ4
6YTauXB7uNbR4ldhZKelKrkHXs6mQktZEFdz8EwCJQbju/APPH24f756vMsQVyPC
JvhMcyNNy5ryL1/N0k/eKPlvvYK8st4lpIc31CjzJSjLHhw/u62UKSYaKHsEV3cW
PEKpJ1NVr9Hux3borxoDWMQhN0azWI0XQrwIDYtlNAuHRbFKh2FnR4OIInJVjxOu
fmNPkjMu7ty3xd1bFuSYsN2WT/tNZA2NkvNYzm21PS3QEJUzhX/kG1aLBEof64j7
HYZPiNA9ydkS6EWdHofylF91BOweJcBkRoLeqgaKg8D91lNv/nRm/v69h30FYJZE
QO1aeUn3BiRWLuP/52AeFPL+AlcCPZza/YOMiZ9QYbrUjwlEXiryTPQW5C6dlrf8
JAZxIdGb2k7bpqLkhAF9mbfNnNl1suNNFjyrkoWv4CK1r/vUVE2A/ICObeoz1BMI
6TBuvm0b2fDqoQ1Ijs4BM2jTtwmmr/jwYmauEzT4AP8q274pwXeBnfCfD7XiKSkD
c8lyooSlNHyYufM+XNIfAgimyfAXSD+yti7nMnogNTAaS8DbR+VMSbDOFgH/YiJP
LrBslJcO2NS/8bOqsnzFYIQAjdrV/JpMgcnV2CxfwLZuEe6R4EYkBcOITieXj4k5
RkKFMqcoA3RcQ/tsAoq9M8i2rnAE18H2SfGxxNiMDy5GgS6Pp0rD51Jt+DQq4/GE
UJ1VEELVRlr2mwHOcpKaPs5QbWT8aFwqRJ8M4Fh5q2xX/s7C8+iJbfu7NpXu/f8/
ImHnRDIytOUndegh8PikNKp7+c+WTuvN7kHAATb6tVOe+/FA4yNyJHbRUazXX9xc
mmQTMV5fRzK249E6DavYrxzZGbkXw3JyupJwsrZTHoqnNt57EsSimlN59nkPaK2N
d+5n6DDDLNHsFEzrbQWEWwrJoxKziq/9gdy8N2psHQdzD+SjQdgPohjvfR54ah0x
UHL3NYIZiPz6chlMJeAc07gqJe38mhnDnAdfPLWaFELQIgVhR4vpTnuQcne0aFJt
zlAJe5fbXZau4/mAQ8bmy6BMaZ2GjFfZPwuYrePfzpnimcPNcVQFmhWW2Mc9W+Zr
L+h3AcLPGSlIqzQ2Go0u6maygbpGyfeq3JfBISXJ9tb3GEaAvsjLRcjisni2NjXO
r3gvqPOMUGs7XadvMs170eGFwWM6mD4xoe6uYjIOs5MK1IMZsQaUq0sZbq44NuXr
xVhgHFKDxKP/f88Le6oHg88V4eQRe+2+izt9LOIdCvGvzIbXrQ9QEzl6Q1H8MBMy
CZJTrvLUz+dju7Hi65Jf3OHn7kxgsvb+wBN+a5U9AAySXzo39ijZykYY/2P1F2t+
uo2SGi68Tk7B8h4U+amfhiuHY/P5q/V674rYSN0uPA9ywHLDmdS/UhqlBf4GfChl
a8UzdBL0cYiiSogmIvexTai+3UZQ36WPBsf5G6iGRrq13rvPKj6VCBYR3cMHmoMw
Vz9P80UrbRO7c3ldgwnd8BM+VWNuLPYDuNLwJ1tLRGEacSInsXvPuDdgnuWOGTcm
kZvu8HJTpQLeFyopZCFzsG/nOdUcRWDLAjh4o8dUoqdu82ZkfuxcuUXnzPXTsalw
37NMNJJ7vVM981bV7w7HplMvgWFltExJUU2+RIUQ8la34Xv9Mkujq8QPSgB7s74R
I9vKoUcCKCq/4+Cp2V1UKXEjhi6/s+uSVy1zaAfUTdL5ROilP6RO4u2aaFQ/Uc1Z
Pv+Yp5jz3H3a2LzgDpU+TBUCDuTYQvHUs4EjBu9I0rrMTwNBWmF6Lbp0/UCZ1T6C
lfZlx6YDCDkzxAC2YavkgNAHqKj7odzTCbntbJuwPeFNpWF/r2TJLawtwMtYchwJ
PsozMpA5weukQq/WJiELj9p0fCwhmqAG6E5ziP13gNnYrtbQhS7N7eVESgVFgNrM
CVEdUXJkfP2HvjQCeFV2dXwJLGUekCVSh6vivGRAnByxmbSbepAoO9am91IAJeIB
+bh95rRcRK0Y1ybIYVosUemq3SVa8QRj33W12zf2hgBqS+XmlL+xc2ANRsE9A3Kb
re9HosXk3XGrtEUFwVOQ0DHs7XIJv1yLiFxHEEUuKKWdHEF6AIdwUhv0y3/IzLPK
fe4d9YsMVkNk2vdYAS2e/9bdixB1L/6SZws5dHetr2SfsIs6F9BU+U1Buc0FzvLF
fwDAnF4MqizQ2PXj3T9ksz6dQiGXmbyWnfBgWbnX0iamkJvlCfOdFcLRgyUIP/r2
2tPCX8WQEW5fpEDvszDOnBicr9ozdgTsDKXUeQi4rriJQSb9eo81lm2wRUAAms2o
aN2x6lD1oGuMvfYOGHjlXEVGVhwRKutGeWT/ExJ08kAC6my8dHB1+o6XQpjLxcq5
M0ZDL2VQDyDk2xUoVNxv3X4Ue1MNk582/Xc5q/nmIIXwC5kNzHygmdO8C3dxlMZM
c5r3oCwLlpkDqdYCjE2R7mTbUQA+/Y5c9kLwN2xe7tFmciIIP8og4ADezcqpwWm0
l7yXZl1UnVbgk9TDo3vza/YqUAac2YYHANDjvXNxKxEw9O+iGpOafSgSAUz09SRr
ueQyDQCN7MPh9vUEev3gAnO2nSNE28WYIEJJ9kckkb/RsMd7GuwFlRijZG2fhMJn
7eGaFOhprUqxAUw6LoZhhtAoBb6RPRM+h0TAmf6YUolXVF4qtPYqDHaoErK6YKfe
poaJSEZZF37+iPdkjo4LYu3u9SlUhREunFReKRYu2dxdXvsjYoOdZn5amLtO6VNR
A854J3K9Njj69MAu/kkWmgZCjWkfnjN+BTTFUVGzJ7pzpLe/56k/u4qPCX+GcnPA
Pk4BBfaCO9cb37RN80GhN9f69XK9/mG8MdmZ6UwO1QFGCPobhjxbcSwxVZ1wlGkQ
7KYnN2nQorSuyD0rRyTwrsd7yMS6mq3KUlet5OYcMSjD38a70bBZXKLlLE29u9vg
21Nzr/iGnZLMUKv3nN883NaSFykn7M1EU7UznInA99P5Th8bUW7eJJeBF7uBW/rA
6OXGdbuuTjneeHb7bzhdUaQAmrJq61iEIYFrm/hVzGyZX2IrW3WuOmfjoih9tPVt
TzLEBNzykvF7CPYyNiiZjQxlcyKfwFIZB69GuNV+KostGqRDefAcuo1VcpkGowKb
LYfQJtQlCaJzoiCPCT+64f8R+wDnWKQss2P8G9LP/7jHTaCQ74ES3IsOL/sZ7WwV
Ew2HVtwpGjNmKMh2ExjmHpZnubFrgWtB9onUo/49uf9X+WNtKy8xF28Xca84Z9jU
Go4YC91lzMfo0LkiE87hAKQMZRTgdqbpa8rqsSMOrhUnEskYhI7oOtZUeMwCqhDx
7Y441qyZa+feQiFxRX0NPU36p5pO5IdJEOJ+6neaPMBC4aqXkatU3W1LmC0wDkOL
ui5oFZV7/WyCfdieBOZwA7XqcGvQZ8Co73REl9zxvYO79E+fh/1OjV2pvzDnghIb
VlAX0TPlXmEsB0v3Nga+8qu8yb6trJyEVx8H9W4dtY/H7FeqUbUy5f8ohoXOfv19
GjoNOIOP32khiFS4ASFkJnHNYO5YsskEtH/qp/pcAewhctcfAFxN/JfchYffhL/8
DdI+/8hzZwKEv9fBRcV7b3owq/KzKXVYJVR29RfmWPDf6cLVp4b4on5puC9+77Ud
PLAMZH3k6ixZv1Qo32NUAVfj81x0b63Rt/DYUFpSmxZHmgXm4jw0Y0h0otHX0Vzh
22cyN12Pk1NRqrwhO1IsOHd+ESPN/WtLjfRsypi/q+45af+l5lsmoZcbz4CJC3cm
Yht9kq6oMenTvNEXhX9IKuF+OaanEyTeWRi9QBe5K92NrL0uVae2TtYhHLS6QH9o
zHxRj/DQh/iJ/L8P4qfq/6/YQfCs1vBrW4pS6MOxkwEkQZs51axDMwxrukGgwybr
Pbq5/QYm8jMMCImGhphv1T5EM9fVZl6wxEwOb7yXi3ttXLJk6SWKuDHPmoVfgABS
PLr62VdyJoezuidnS4zbcTEppkbP8W+zfL8tvRZkcS+1JfUJ7+sq9BTNaq+O3PUk
fEEsMrXaoqwJ4/FaorD7SdKv0sZNIxHVg/hrrAQioMpMyukcEshILzdjpswUivY0
asLTbY2CIG7WMRbUyyq6G60Tpp/Q7CmLqlepugKMXNs4c+iEZiAy1r0y0j3RVnaP
Mnoj32U3zgfM72s1ClQXwVs2EX7gwcb+g/UPgaA1FUwuXIt0gzh2WeoiYXoyAkmw
9qvnybN7HgVHc8HgkcxBmzUb1y0PpHyw63svXllScsnadXjcqio7/D2MPEYmaigC
FOJqnRBUEWKd4kiHkC1u0ZxmYGEWMN5FYqLLMr0HRAL5y/Rvo00An+j52uNqLsXF
4Qof81X5KDzmodSwTn8J2kj0tLzOAxou09KcQSf8QbQwGDLNe49SS0JfWPpd0ugs
wBFAoRMxu7+Qs+mhGGb5dWhBT5gXWxCAr+B+MaBKlkIV7vgPFFSncqjOqEPJu0In
jLjP7HfBOldfg1iRB1qIae+eSEePayv/iDPrJ/ohLcWTNP+tVJ2+KpkbHDBHlv0T
vEyQ+DmVA+R6RwUhHdVbp5VBJ+lxf5MGqqfCq6YmP2z4T6mn1QW9hwtLU9QSHKSB
o9gfORZ/oUQNppMXG/hAMm8kI/ItXKrT2z+WHTlHKWuyBc/rrDdtnpP5abm4n1Hn
VzNNyugvu79yrW0eVq0F3CT8Qss3G38CJvjbnj6HoYz1rxgMbRq2nur7EbbI5/sy
O9N2MItzrS1tK1nuyOUgVj+IvJCPGxxodYKEajsLhPI8cQwVlnJJzPV9khJOPxIk
f/w1CdgiqIe73/piL/TOmV/4gO6p1+O2yZp7lb+BB0LRydBR8EQvZ25UApNhEr8F
6MYI8wknPIlhjVCkjldZ6MERCBl22lXB33K3zq8odgOt91/WNsRnAKjCiNzmUPi5
MWz+Qh88nebUuLRAzMNbwOMnd6EBWpNXxnXuUN7Wrs9FWrCtsdGz+vwN2ksZXOOX
CIK5sIVGxSgo54z0cMf8Xd2aXQojTsYF93e9mF1zAkl6lYGn9Jot0q8O/YNPP+21
teusQ/s8QFgL1QWpzQHnIJj4rDvzq7nQC4a322HvgJLbsQcLhzEj6b1i2lwlb5WA
5LD/7o127+qajKS7h9XVR894Vimfqk9he3Khu6eQrIK96JDJzLYgdxVEB9Jqwd4E
piV/bz1dt6hKcYazKDFDBiwgMhwxy4VS9hMHjEK2K4IgKj3hIuFBgwCif6Hj+9Td
3PoC/eRQa3J5RUBOx6U1bfS0b7ELgsRTXO5cWr0gpyKv8fV8mcSMUvnFLwR1I3UU
JamAT/ZPUfTU/ObbCv2kUoFxMj8jtJGl0KKP0LJSJz0ZW1uffs+VEvSRkClpzyLz
PCbeYnIyQNzUQbo28msIpiyRiCKBTOiY3mw49RzXiJM08Fi3oQUZgsnRJaTz+3KP
kR7NO+gibKCks51qYhpPAKYwmTuehVY+L+PAW2ICK4iHdEKZQw/1/CUijhGcP5ER
o/Hlv6YEdKEMd6ToFBWTaq6QOd2hHOSdhpV40mqXG3xF3aKHV2eqRzXITfqVmaFk
A1DWRd1FlW9soVqwuXc1blJm6k+47nf0C8Dszg7anMH60BGdD9/c7/ZXJWkVeTyr
K7Y+rDtJYifFsHvjKnjuNxTRSffxZraGHztEsZZyDMzvqbMpk+81L6DlDUraPM/P
Ls1/aqrzT4nnhx67M/UtnQIhzpKX1VrfcrT5Yw8/dw6IMEz/i3hWsHsZVHtnAurX
vXcFtJe6fphgvvnvGt5Yhpc2LKog7FryAP3iGSt2Q8+WeNI1KjfWlMsmOc7rM7oi
M9xwJb0PLIDyc6ONzLS/vbGkGamK5ZJ7OWPf8g6O+yokWX3gzYNgO6Viv/4uViT0
qo++uVfEkAYjXq2Rk3vxZYuRujeyD+IzPHjrlVYS2J7nZlWBAnTW2TQqcKSoXkRk
ZuofL4uoMFkUWxfTlPjAszhRgBab2RDlr3tvJCgMoWV0dCZvoX6a8NnJZJ1MWP0u
gF88DJwME3flb2C9Xz+3YZC44CRktW/gRvEDdKulWxA0Dag/xrfZPqGpHnFG5aYG
gO6OtPyJcjjQPl+26JmcPMtJpsonSS4C9vWnQIqoqNBQUjQ9o4P5BCfWmTGsmj88
aY23yQ92Xu6Gdf6VElk1CikgTF/XrZyFB8e6zxWYVqjyPLzueSdknVtAAYle+RKX
4fwj11t2ZJBYhHIlSG5iPBgue9xdqndM12K+WX52cqJcBrN1kz9YJaVuAQii0p3h
6+i5KgrGI99Gv2E9FqmlpVUGObN7geP6sQWy8whY1+SHUFb7X58Jq/yewU0k4VhS
6YHFfYMN6bP2o4BtaXYJaOPbR6RY8D7iSwYfBqTI7L5bPrvqvcvkBzlFeXDiAcJQ
jkn99S37PTTn40CSN4D9pWBnyj7cTIgVoFTn+RHuciLb9CYxL/m3ZZVyqVEhVN/p
rQ4cjr0RTzug5TNyKW8fQyIDfUiMVbH9TjyZhMzA8nEWoEYNNFuzBBgxnMssiaix
0cdONaQODlppWhERS3aBLVvMxyi/3i3MYlfzXuM815hd7KjQQHwVS7HRHFEao4l8
BgHb1AXCDxkmZIGwo+hsxYjRNYrLGrbf7xdiJ6EE4yQ+mrd6gNhl4IMYS3wuqQA9
F7Aarvx/e/EECNv9rWW0CnYHQ8ja/a7T5TXusdP/tiIBaVGXyqqanie1DWWRQyQN
hpvIEBbuj6Z71hdYGRCYftFUm/41VJktzoO2ezlpOjhJiK81md30QOdTaI3C/3Kp
E6lzs6+VE0GHoGw+g6fPvHbsopaOPRSDPkVUxIjL5Ax1vfAKsK/bW1mBjAtxdgcY
8kFcrSxzCpb0B6L4dDerocGdBfSfZI1XoNnk28LpXllJ0x9bvmlHsZrc8iCgg1Z5
R98L74nTWiXhCWsM0yPedp3zWQJDZMB+jIKv8UUC0Snhl/RjDNt4gZ576i1Slpif
2F4VR8hUQdAj/mcw7gD2fie2IryxyGV9PEu1Tk6ZFQmCNmDNfX/gS7bKhOMWh+gy
qY4pNhpTkBgwkDxtw4VeTe1etDxYYq8rzhjiRUsyr+pMScfHNEEoMv+CqdWGqtea
Oh3tuFReQkvS1epNlVgqHDAR5G+vvLD4NIpEEplAtJUcj0w/mNgvT9bDIluShrz3
uHs+CKtNEx8MArhjWsYywrq+IpuzzdwRP4H5K0vfP8rXvwXIidKQjwHTmuqCALmX
oz+fes5Siw/RJ9qHDi4LLPiOYY9vg/hyE/0Cx2gMbVqypIOnGdaneV/h38DLFt8G
PqWb000zSC8uum83cN08PLYEf+HLWJL+DVEzkU9JMtwA5vjY4mTSz9UPD2/7tzdU
luQCAAN1qeXUrQf6XtlG1HujBBPFkWrQ80Ge5NnIqd7G2MwcGNyQeuiMcSax3rlQ
CL4YJ3eVscfEB0w3Ck6gU4fmI4nTqHxbceyYzF125zMeWVCW5m0y7xmeCEtVEHrn
YbujMxYVaa2Qpa6zhEgGYy+Y1MsBbx3UYUmBnHuUl0cWsa/ArwO5QqSTlaAcLhOw
sYK0hPaMy75sIrrCKgpFu6+ndfGaOJwLhYy2ASCNibiyDhQkDxPiiauh/iIFcSgb
Qk8KYs2SvbzJFxqo0Up8MmbtEK/h4x1S9QMMdnEHK03ll35Rw08VmHexpaZ1yDbH
xUuhJGsQSIfyHN+BhoJkn8udnooWiYEBdaWJ2qiJatfrPvu/p0fBVdKx/2nTHtc0
fy9RsqfP2rG2Qk5Y0zbPDAtm/Si15T4gPzt8Ch8cYiS7NGfwEyrOac4AX9U7Hcrr
IaoDNCr7E0WIhYCDGIGnuhI5s58hhDBoz7UGSZ3LHxlI1KXYmEm+FK4uZCznTl4Q
AAb/IXZnqt2oYYLhq4kw/noI/dtZe9HxVzBp1ak3utV7pT7mmOTD/5u8W13djtI/
KzX9yv/fyT6MhoXQXKlXHofLNWjC8rfJUFdNBDP3vEe28Mb/j0DAaSaXi3qpQ6vZ
iXajLl+31IBAQ2R34hOhf35Ci2LxTRrh3Q878sXcsL0rzo+qZzCgv9Q7UMMGmnLF
csXG9csi5gPUum9jD1u6dQGlJXiS0VJ667J4GF//u7DARM1seb4PY/J02Ob9kCF3
4WYOrIRdn1Ura2impxDHk2a7Z0ITfiXLVVLB2Sa7oyLdEgAXPeeAxQ/+IckCjfRp
yoN3zzazBpa4TZjND8KfGenLT2RkBEBUkBZHfJbfmLG2Dznkil+y3jxicsM4x6Wp
I86Y+Rs5w7N7Nv7f5HH5mv0BSZFDO1SBUJhp4ervJQsZLT9Pq/DE5u3uG8KqYB0u
WUvIvq7ld+zSUVV3WyIYk7GPdmBcIfNAI4obVDn25Svj606JHpvQGfAJm07s0HmS
wtdcnPOuuKKxqt1l4m2ineWLPE4IHU5w1NudPqvDWPkXVhBemzr7QhnhKByq8/JA
/p7lc4itaTmRWXk3Mi6ElKZe+yLYJjsDCGRlKOUsavXa6Drszo6Xe5WsFm1UU5r1
39OO6RnKcOFVybxKxm1po+9KB02X8K0ShBMJIS1ptoVxc3Fb4707nKnLSnV2x1lC
of5B9M0Jpjps0Pghmzk2nuPjqA4Gj/YNhPkLwS0uRPYzuYnxhVHhxQKyh0qJx1Rg
MCdF+SweWDPrg8nGKVXTcnTtOAjgnapSr5tQsnUKftlDmE+/x5ukXqh4yxwi1HNr
NPbH5+yQEo4ZhYEHUM96xIis8MCETX4GI3nbPliKd/aX2asVsO5aPTNi4L0KdI8X
rfoGxFZwxY5InaUoQVMFUoeC+QPl8erUUGPM5rjUpy5BIbMx3aLS+7WqAjWkIqUm
bkdI+C/gxsw2741FWlZ3xRFJKMgVB8wXKwYPrWeM1w59bDJ3vgJM5ukWk0OhUoBx
aDRAWcg9jeNlDCh19reML/SMHUw0K4FKHwE+acYg7jeP9FcQTAUY7yEsuIeR7hmu
LP4DhgIhGMo075VNX/dYxOUP9NwFqWvxM8aAtA4e/1xZiI/A5lGGPtbs66UPqXh+
AymoCXH2bEqwmKtJsEfxHpnLtBsZNLlP5DaEq+RCPrYGq0uT7JbUcAj/Mm/vIzSy
XYrw/LYXVaWd3m7+UoTdsbAPZbaNXkno3UrpSe9r9PAjsG69zgtrv5ecdZNOpq9Y
eEI7Oq/4BHn6BCsHydkqs76RwOKm4soi8gwAq4C9ffvYSzCbC5paM2iOuKiBAP2E
hcB5hCIDyvPyZGD2tpkzazbfrubx+9pKq2s/+E1nVVFmO8WBvWR+4bWiwfLBO8aP
34rrojhqqy11+S4dK60m95P4K+OcIMqxI3Z2E5kMv8OkyTW+8kPX8ie7D7l4gs+F
JgLx4W4PXDsLbAxKMz+lv+gR03FmgIwWn8MnJ5xfcJ81FWKMeSTfaahNu/0u5xcp
9YVoMS01ddrPvjgZuBEbFr3VzgQrzMTGDds0fxfF+kQmt5QWtf3vPUt4zIg1Tx/g
bxk/3OlveXVkS3iKdUVRChLpjOfa12rTZtXFH8vdnNRBG5pJSstwmyPf4Z7GIBiR
T2sqzDLbqqriPcF/w4RXcpflbGjyDnZtGAY3jZAUc6Nmc/yBEz8lkmCQ1J5oZ9vZ
IxmqeUKDUYXE7BqTPC/UfecmeVinidBCHNrlQ5SNkwi4P+g5dsY5lw7ypVkBz79J
J3WnJ/+03xivd+m/NiflXCxuQNwF6guGGK5T5mge9Bt5JZIPed/37f8MSrypAqr5
P2XMSsjA8bvpG8r4Zt8V5nsufC2AMCdcB56XSx3riAQIx8kY/KGBWgNa1SPgZbmc
f9WdJ56WdryNN0O4pygsQ3FPLRyrr9l3Z9yfSdRIHWzSQE/1zlP8M88NWVj0XWeg
N46d5UajcSSqGfY27eHj/XmLgXVxeoRliqm3DgQBsSKPHe+gvaF7OF2sseayRR8H
t35wFtCd78uWW0ZnCLAzRM3uVWkCsFsMNPcaJSws6WPyQlz2Ia28LUj847elgmeL
Q92GJO0xaCe5/ErcMWWqiJJDzojMAjOiqA2599MsE/Eq/em9E+kU0U9I5OoxOPJW
pEIJMcy08T539oAo5PQ0U9cZ38eiP3xZ/+R2XpB8I+5etJlgV5BzU9+dzXFecP/j
hBQ90NUjbVTFcHQJ3egq1SWF3rllZToZvBycLl8Ujxe95nU+zWbeP8bM456LAAtw
0R784D5RSU2zhmUwTaKA1WurC9Z6GN/venZCLNgn1dU77qf86zN5FoiCJBu7O3rl
I1MrTlli1htZIi4xyhGlXsgAc0teHF12c7MYs7jLk1HmW+Dgs68SmwtuydV631qO
I5su+Fky6Lazx1E8ydigwwA6QqaZpX9KdR5B2iwr7BJ5NjCFFMPjF4OrN1vUBRex
g1FVKkzaJ1UtwrDqH/JooY4kYjPRXKLpoJcOIhRHnjD47ZFPFuFq8LJWK9S8356y
kKQG5rHpgZQD+W5YuNR1hnKf4QdJk8WeXqyMteZnvkHKLexNkyqVnEZTxw2mbHK7
isFNBkLl17KKrKp8PPiXVdulvddVo1sRcny+nmKQvnZhrm5lYtOToXH1ciHrUHul
Lq6Dk08J+y189T5+zMZRSzYuOvC/tYV3K/NNNllN3BKlmNbv6lMELYI1G6tzdzjR
XPF0lsnq9h42umYJiiXzZ4zjYNjvRzQ8317GqmBaqtwuXK2808/W7xJCJi/NVg7x
mgWqQ9HnLFKZLd5M2zQLfm4lICYLCk9Yz/kfESQchLz02AdehF9Dw6eLVDQ6odV1
LDZFb9CpUcYbMfLlb4HxPVz2MguJwKGOXM69RJsRNKePKpidIlBwN0/5KMhw6K64
hQgw9YuXIj9S85Udjjx0/ds29y5aVRBpuWOjCQZSjpJUrcbAhL2NXw5Pr50ZPtun
s/VDrJm6B0ynZWB5PX5VXVC2ghm5zs/PUkUjt2yzIiCLOAv7A1jGh3ru7Xoz8PCM
LARd+ttVbTAkY7mWdgYCyXg8jPXHcnRMDlNUIJVNoxN9oZ7/zg2mEpte4tuosoZ+
ZwHvDR8gFnsOrMbpXNDjO8Js1cxzbCA6R2AMufzRzxUWV2s7Fd+I+wRdikMZcXr/
oQj90MUGTgtm06XWqhCkWQ/Dzp8WFKZ5fCaXP13VtlUMQgwOXSgsWrAxA2/AD04O
/jrL6Il+SexxDK7mL0cD1NbUyIZwP04Ph31Y0fffQTqgAr8r2xeXKQeW8OmqiKwl
OapdQWFOn5cccR7ue3CINNs/GeburZ0jt9zISstFY1L75X7Cm2AHpEDlzCewBvhZ
Dy9hEQ5u/U1zB2t/EeItiZ1KarBiQA07GRzKsSRUPNrmEsIACyXYcdCyjlBDmeCA
ZLSG+oaI56kNoomDTT1nEPYjK8Xa/qyL6RLOpsZnsJ8Re0hVWU/dtjH65q5AfvkE
b/PV82gD0l5BQAWQzf1Kkd6cqMo7QqCXwLiWnemar/Qi2EzuSbrgZgd4xNgs46+o
haodAXfjMLJtHW+KCZT5s+B63zIEIEV2vvl1IZfoAdiMVRyGoAtaHBFZL83MwMez
0LkeQLmvTPmwcX8+XGqvwlqOLTWdxlkMLqtOylm4pNwA2+VqPPEzND3TfFvMFFwZ
/24ZBxLyxJSe2RaZAM1cCut7ehEBQ+DdSNBMn4a5AzM6BAl4LfI46Fa74km4u1Dn
jW+F19DLOkHAqJUHutka38XT4Fc/DoSAlaW5gu2Fu+66Nl3qNk3slyHA8vtBndvM
pXnFNrKrXme5uzPrZxL79UhB8Pj+Jpr32xNMxElKicnQ1WqIW9hwd0dx+jgVuIRc
jDe7DtWMIpSIzvFZYbFQir9EaEQ+UkNl3eqzg03Dy4hOAfCso3qzKD0qVDDhPEQ4
h+XiwN5zFaiHqi5j6Xd5AhyIofJxgx2qzhs1QukziLGHDX8bQSfr9JR5oYollRWI
UXdCH+oXIHpWppwSFe1h61C1k46/A5Z6jRkG0v8wuuxkooGp8OSiZc15vbmbHzXQ
VXE6YMQWRj33UM6HV/LIj/kskQCOO2wJQsGFC8uN5AaRx8l9KkEX6VVu/JqJKh0t
NUf/L3kTkgRufWBHGZzerdQgnxPxBgFFxg7MG6Nk1tPIBK1JoPi6me2FdrXfuxuf
PV7BFOA56DD/DhS7CV2fcyPimTHLD1a4imEsYeX5IisrNp8PNvb/9CtqvuCMYpsl
NUj5qCYkqNYn7RjsOnzOEtqDwkdrrx2e5en2BNjumkX2Du8NxaXG88n7+s0O0ac+
4o0z8YSUPqtosJMkUTbkWQbGuTPobIOUwBnNqqX35arMn/XVVeQxLLw+r3zYx0mE
5Y2PO3zyVVMDxyGlsioL9+NjSAJjH+O6psIyJATe72PntazrCHnCUtY/qozsgRQG
oots4Lrxmpx24MUqXiC0ik32/qyl2jNoNuFXH6eQCNDFFmxIhTPoYY5taQURfNOf
cLs4qYr1W3/UbgEZnAnPskEtFk6ypnhiXt+NwjLxy+YXCD1teNqyc7YJ1hVaDGAU
3LwoqB5gKmqFUVD02GsQdpIG4WQmO8J+khfes5jSveM5j89iruIRV4Aj8GEJsczO
dK+zWz0zqOELvw2/KrDZo/xKLhrr4w0I2uazX2rwx/b2w2CzS1T/Jw9yu+4IGD1f
ocBEsoNEYkAfqaLRbn9h1xKeMxcS5yIud7pwZOqrlRfsG6jU7x33N6hbp79EYFRw
AuWCS5oFSt5dOQP1pAK6vr+ZTdQQcPjaGzFpFiiupgQ2jY1GLrzAJanlQ2RFPUYO
9YvL7oJ22uJKHEITMiFKyUYdgvBZP99TlS9JC+UqAAxcZiR67smmUFizvcD5+3A2
NTyRR4kuyADDcwD6XBMz/OLhJeoMUpPLo8/qJK+kxTJUqYQaS5ka3b9hbhaoLOE5
03IflrjcneOTBAC1r5nzboXes2/TA4a/HUAoji0pQixOf1aslJbpAuVuqteFukNY
hlLDUQKCm4euQNm7e7AmcdgaxC2gKS6yhmyrKveQArMrtO4vxItOScPtwt3KJBNO
Ojh9IjDBS/NgN8BhtkMK2hpifJ164jyY5Xf9cb2Ol+oaP7AftXxAvs+VpBnuuv1I
4HvEb+zC/AoDwIYfL2haezuPhyZsrhZimywjdhQjIX1NU7w4omKX/f7Lr7uDDtFi
RCI2YmFrPryJVOcYAKIG5lJ26vqXPzgAJgYMggY6OXmGlx7z7KT6496bBh2+2tcf
IB2LnFYyv7A+Axu9HenmIpkNFY/v7pKIXeq3sXEsMpDxOmUjAgt6MHlX6+nnz5Jj
Q0gn0BXN1+LUXWjtbUirSWUWH3OZEnj7RVjQy4+5Ebtm5dot6AxuTRo5i3oRIMTD
fTWkvSro3WrAsOgBFLVWz5AhlOSxykhkbp3zIjj3UhW/XlN++uoVZb6DVjR5caqE
WCeFLriZZNJQu2EkGvFhjGgN6wbu9fhdZyRQWIdP5ed5vfheANQerjQPSmao3v+W
0jotm02golsKznHMlfPLh9RZAm7L/fxJ9KONj7vmOf+WyqH6hU/AxXkhSJd74PJC
uUbpHmfLKtAYy9szi0hnwDj0WPdLVepy/101H5+rjRy+CZIonpA3pao41uBgPBuL
bKw0cbKKengRgkzy/OOtXsseW1mr/GqQSHnQ9PIahJNcpbpGbo0njimbZENOmQxj
zfmKxNd2gy4izZcBvXNbXxj8VHUovuLaALNftk8iqL2NTZ7ZwnCjCKQkOX3fFA88
WNIqR6DwY4jRlG97YNPMSeQdESilXBIF8rCiDvIXDGcgQSNoMGKQGEqdHpMvjaID
V0cb+dYbyRKh5BivZGZ2A/gZsSe/NGu+O3sg86ZWuYbuACiTCbvK4kDeYRgHz0r2
B9KxfwILwpOvylGIgHCDErkOoo2OMV0fpgJFAwEYHvlzZzclCXjYiIJBkMNaXntF
Z9qOdeH/+IcVtrvNyjAVBaDM/ko0F1qpsh4LV1xX0P2PDAV6Ftk/ytmqKEbxj0uj
MSe4cwHt303dpxConplqDhgs2X+5nMfiJiBc/7813A9WkaBPMgHevC40f6ge9Y27
iMYDeQX5gFzt9kHtC9eArsEqOW8hJdOVt1rDgkNMbqoIMmOO2zvAtE89EnAinrip
W6fByMmXlucbX96umJU3iadsLeEbsCHecpsus4GSIrjfZCkGoO11567qbWNCWRRi
PGDVhnQq7JBijzePRpPRwASURZYO5Al0qaQ8N7ULk7oOg38fGDI9sU7hgGpE0r4I
fey43GDHVLcpJCL9HBVr5OxupU2tMKTAbDw3hhO2lA1i4PLscQFaqLi206oCzmdy
pAuvDRbT2cxYy1PNy+11i90n6qdS42JtTnLy6UwTk9L4qiYd58flzyKol0bby7sQ
QqBMyXr3l41qTKSNWrx0breXqQRGZcmnq+QNJ+N7Rt8/yKTuf2a1hYUUotOBIf7q
/vhzpAWcCKUYZ4Szxyo3ksGDNDN56a3t0+dOH4jcJzQ+1BMK9uwPeycon9/7cknF
Q1XzvRMTrqrO+rxaASB5uJzhWXp1qpk3V4bJ887r9rx1B5W8AelR7mERDXUmoiGL
TfW+kKNDmYsocrFl2A6LHsDRKhL3kbDEmRvouVvz/vpQOBlsyl4OrqGNFP2J3f8q
SDsidclBx+bO+cXAgzJWUuLbkhQuMbG4Viy93X+idizY/y0Q3Jtp8fLIMW0kMGSP
1frt3FG06k7wxiwWwKTeF82h0qI7uQF8Tf/6oPl0b7AelS8LssXGGiHGNvESyB7s
cL4WOkqg0wxl+4S6odsz/CO/a+VPD8zOqf/2AFLuU3Cu5XVfIhTr8eGEwQKUKvqQ
XWM4YpilHWZoqQvZYOR1/FVPEOuzCLPRxGtA9CZkaHJfsWShSLOY25RCODKqzPO/
XNv+42kk43Am+98aMw2UuS9SQxS0gaJp5jQk3CzJQYu79o0401RAoZVXz/4gyGL0
KN7dQe7lgOORKNh14hYAONyWdDJBRgdqTh2TYWRwoi0iZy3Pw7XtMfpPx8ubJyk3
2zBjeNXBh6LDS2e24aMpEQAXJvMtTFfyfDS/cvqQJ13b76m30lnIdENHOlBUNyAF
3TvKVX/wJ/ouzSMZZiCDRxtspAKNg0+5eCmCMRMHoQXt7nrpWmM7tiVRT6YZ42WF
5dcs7VL6+D35NyHnr1SetfOXi2gTB5CLHQXWsxe4ccLdGLv80EdcbmZxXVrJ/GXI
ETfWEgPiflQBem/55ispJJw44tT3E+UTQU1BI1xdyd2/HPgRr3SUrE5yCNlsomGJ
f/2ASR/Ftez+dWJH5g3PZcA+x7ldTOX8ZS5cDyvAdcfwrMVknqmgSKpmGl/v6hvw
0LP9Volw58HETUf4zJr/ipGqgV5bb7LMPmGjVHu8nu4QZ04u/pa59MGXtP167H0+
lBhyIsdSX7S2L2sFgYMA3W6YIeQeavVpzlTMwbDSXK9gdNVfA5oZj/VVq3A5QiED
10tyAKyxIKSAtwKKulTmjx9ZQ8oigJXUeg1qi0Lo0L/CvyctJAU3aG+Ra1w1rXfJ
nrcbOWch8waRj8O3Riyspu6Z+MXdr4G07gSh53gob94UNIGzXHCsOadExDnORbne
cl6SwGD3k6IBHrV1G5AMmGLxlrM1YVAYw5ermnNGhrp3phn+a4/pPn9OksuwAbgz
aCMCCJbXgzTWJ3bKzOjeSs14B56u6SGZhZDaUbeAr6+hcS4wNLE2q/YW+RjrDe5e
gOBSpSnd2SGiUgk9flitmwEpW2hl9Ba2eC4XayPcjAk0MUOMJ3Mqml923CJ1XPU0
GzIJpCsyCklBXB3ChZeotFOrh1AW5rd7MnQuEgBe6rqY+EmFxpfeOGOi0uNnnoPC
a4Y2WpW3RrAX40FuNetH4miO8/rGDNIOqjcTVZDHgfTMELShCZ9+qdzwZzg/ZVb5
uv70p3Pe453BB+smBHXNMTPYvvRX1gV46ZealNzwGLubrBr5gvNERT6JI3yoqq1v
WP6CXExbCgXcIrDi1UJ9MRCAcmGjdMqlhH7LftPYwM2XZPOveLFC1cLwolY40g8I
WA4OFmlv3N+xyuaR2oAQPCYFINGCJiY+uiXkOoBNy0k9gMmyh6YONRTZGdylRbaS
gCS5OEOnpQct1rWTlxC6gl01K3PsHMv/7Qg5tcclR4V2fsUfQDDZQkT+XRSaUwMa
YkQmTLB1z/SZvi78GYIFHWR7LWMM2Flu5uG9DmGOeYrU6VQMxUVwM7ferWZusuo8
0PDCKFNVHPPNNUhsATYWFjHT98QkHMQGW2ObtdFmBhUuS/CNRlC61Ivyz+AfYUfK
qrLsrKLdmFdqJJtSpJErS+xM98JxT17MQ3ZfZHaOe8xJqpg+k3BoXU6yhqNJmNxC
ON/+S++Jr+/gS4daC+Kcqc1P5REC1hs0QJpF3yx0x0vKCRmmz9vJeVLTpyRpoDg2
1/2hS8sxK3bflVWFPhNt2usQfGZ6lIbDLyZ8Y41o5nyuQiERE+1Ya2tv1LvgJPQn
bb2x3tY0yx20/4nAdh2eMXEKOXSPlXhMpGBvu7+DvWskBLF8o5tIIBlvT/c1O8pw
PvHs4YGEvfi0/tMxsFEkhm3ydSTCs7q4lSBMG42mRG6fqqurooQmJ35q1f4Ln8ug
jmDWonvE6vyWICWhsSowongFWClO2xGDRNgZIUR2TKnzAR+vIx6lj5kdr/4ca85g
ptIJyLkp47TjwbFKO6aSc5jueNhrQ78MmK+GYK1Mkulr2RMonX6UShjLhPqRgwOO
tDUKti1ANqtF5LJV8tnGaOySsgzbk2jVz/GCcxSUvbPKGj13kIICvldW4oWtU5IW
CZNMdKpA/tRSrC+4MhEcvyYwGZCdjBRo3yyIH31XUxg6QSfJ+hYGg3mD3fgFDtfz
5bQ5n6633xQVtGOVnGmj+ouGyHrlJggPTyDj+AucR0z1MZZNAApArEd0+ph/03SA
tH2e0Oi+lig2EWL9yAuNq6l+AyOO1RDDMoVwEfGc3kc01QQOBp3lPRaQmqvbhvRU
jRAZyF67A67I3gHH4rRWb4zGvuyqv9wrOKZgc52rF0Zgrwzd/BMHi/hEbWjqFUt4
AQI6PvGLuPcB0TzghLD6Rg5pDP6xGS6VA9Ig47QfsEBx1+WygImyFEwPGm/vZ8sr
cqJaPoHO+hgV0QEttPwY9QdOf59etOKaxDXvtRqVBy0SyeTCjyLfCqAtHIEyyxhu
KMcmfLft2ee5++QT26ENnECIebSFvBzQhfq21uDgZjacehMWFMZnubnn86r0h/a8
vdWOB4oXxo02gNAMIuZH9Io7QpwE6Kv4dk1uHy+RQv+F9Xbq31740HL7mq6JbG+b
EqDczmuKXC1pPwWaMaIOlbN/PvRDL6bbEyhR/zNgIxciplM95HLwROq3tJsacdBe
fDflOKLZdf6FCGVW+xVMON+XzLccWg4snmaQQKvM4oqRtVo53BZJ/o/A0yCEBTeM
g036ufAqKEE68cqXL+nXJlS0lYkMl6CZh6ZD5InCUxiFJLflKblOh8S+kKAdpbnv
V9PGbKREpPX8uTDawvyAS4apmhmhizet0JuSRcKrZu2a29kBZuhT5UiYEaedQ8k5
Wf+bgoCnX0bEqL4LAnAP+ylUlp0psZERBcBzGIK1XVUBRmFDMRtsLPUOngD2XiL1
qzBGHkUkxHw5nQZJD5zWKaqLVrjToJ0Nz5jzZfeksacfsyntkGUHL23ZOJigvDYh
sA2mmguI/uZWN0TTejZSe1leN8xcHF3/blbz7NmuH0roFabPic98HKuydgx0vCNv
qW/PZw2u3fUYEFXyKiuwezMc5ftcPQ8TPFFesfSL2cJkZQvotdqpOpTJDVA+480x
7UMa9M8wYROdFeCzI0kllV0L4nspQrWPiMZN+fSThgdZ848jMiINkZkTDyoO81Ba
EwoZXdEgMybCy6KLT0+Wlvyrchy5Sk66JVsAKkbqtq21VwfA8898bw19XFeGncP7
BfGcU6qHpKpf61TlVwhyjyPS7dCu9o/NY4wZ8O5B5YoRvpz7fS6ZyZvY+otk5cLl
Sc5/OZuSZwx1GO8a35virRPhd81eyaMnh1HYotdalbymgQVqz5/QihD/1/H0mbzQ
1Hq6AIX00mh6h/1CVwy33O2JsCd7c97KjXMr0N+++zGpm3k15Y2knb5pR66eiflV
eQYjx/RQ+LycFmOtKLTL6jNb949y2D7lQXorHR2xGEUMw9NXxPAhuTL5WhHIemL+
OHCi3JkcZJmO8LHhcO6HztHaE1l1X9CtoA2Y91E+OxOW3nC7wKeAbvQTamsBqEQi
stPdKUNEQ10wAN9jZHKXkk1op1VuKB4yuQC71W1NJw+dNaN9VMafAjd/dhABO9Nh
5bMJkZbSVVQqGwWQXZfgJxhmPKtozmfz83Cc8gAlk719U25zX3Tn3Eo7wm/X1j04
UvgA+3CRoQSUCrFPfsv9ByEXzFvuuICcnQQ0FYIIpn+r1kWhEcEUjHtW/oklAAsm
AV4MKSm7kzUbJjIvAum/NutbuGn5G671sJSWtmSNYlCxbJWiFUBDiLB8cVDbbQwm
6p0C5uHxBprTGmLVT+aHCF8ySMRa3L8JXlJf3dLVCuNaqcVFJqMZy+ymRS2V+MBw
jeMGwP7JnUFc4jUoW1/HvAyK832LixRevz3kP9nfJ/ukMQ5VrnJ5ghZw5t3ETCsi
eQAojhCaPPeMddPeFNm6CJAANd5QmHNHtIgB47Fmaf2sB13UvANyWBd+k0rUZcn9
GtEpTvCiRIaWnQHOVK3psx7ctOUBYVpblDltaoDnojlqPK5lsqZ918QexlnZUm/t
vf9Q4wCOcyx3aAjmXBKahVHjU+mMidP4TuduvNV7DFvc3cF5lN1SAiVYWPyOW9m6
FU/4fwkGHdvXKXBAU4DiMUEYeNWzELgDALke4jE3WDeYb69vx+UtefQ81aa2T3YN
By3JOw1A7h2Z7dq28eiOJyZac0hywsGNp8HeqUhheNsW6jEC0UpxNp/x1B4+S8Gh
RONfqHHsKsFs5unaXVRielAgG8UlyG0U9QwddaAVwUhZ6nrFTND0T29HDFLbMptW
XeTTft2a3iaKdfei3ZTOZdFhvLaWtXrNfESK1YLU05vjLI7W2OhnDjSqQq4XJKdt
fwOfEDNIfdAwqjIR37yeOQ2VCTuwfHaEQsBQr2dH6+6a3RV7Fai4gh/AJgDpxVij
KHOMmQNS9Q1XcUfSBapewywoHWLl38O8c6SK1dv/iK3mgfmO68xrS6vndrT+7Ju0
e3+OlgeMZE/GeZNkCh/iVGfR0fKx5PkJnRuV7k2bimKPXfCH2rcU3GU6B3dhQCCS
ThyN09l/YKbdyJMPGMB+0ZSm+2S8BZM65/l69lx7fAuqvch7QxmS6mK7FdH8dDlW
gvnHflpGlPIvIbgjq+VwnoN++ySeFNKLH4ZMi+U5yl0VoaLEGVUnUbkv3oZJcsUh
Br3/BL53xemCTq15uDTJk6lUapfKsr4HaQkKSBpjT2kzXcMaqZNOLOmbTATQ1vgl
vPidvHuNdgMyuEJ25O+cmOMDvnOWcWrukyzoEIQ6Ans5h6S0RRjIRIma3b1PBLep
2zTbyARDtJlCh77RJ6SyKKg3yoakTk4ZPi0vbJWssiGpDOL8l3x0c8qpyPemgpUH
2tijQO87IfxNbm8neWZdCv9/wRfTUnn3xm27pfTbRcBrCNC7EEsN9Lih2EwRIZB4
9Z8D0QfXZiol+g3eBdF0Sa2JiIMVXJj0n9CRX3wHG7O3lvurFrbsCb0KhmnEM3Xk
SzHmebeGmcVdH+OZL7OxWBYaQM7EgaDeIEkRvDC/mJ3BFHFq0kOvwSHvgCd82xS9
Rn2r6g/bYQYoxeDe3CDe03ULoOxWC8P5i46/ptTl8lUNvjZ16cG1pgmtYdZsxuMM
vNmbtpKtJ3dqsCGcmdk1bJO1n1AFYmcgxonhqsfNGgooXg4we0/MI3JRQV8IoUiT
VRwAVPAQ6/kpnKQOcVbPDdMldah5/V8jrBdFmtIHqoulucBabxk+Wvg3qODi/w+e
GODUbs6lMkT0aFQlz3dC3mp69QdXHx1RmyFopgle0fjGxAt6eahziofOtRWjqjob
QbU2ym8CToLVBWa2H3g9Ee/yeD5eaOkg5le8Fvm1oK3plx0nojOP3m7DtsNf24iR
1zPxMiOPTXVx62RsTTM1DIif6T1yiUatwL74jXM2JgPHhhvuEde7/IM7rrsbjrwS
AUjfWHWcUCrDjoSThKKNECnRhrveEoDL/0omme+GMZZJsmF5gfe8Q/SA9Mfia5xd
sHwcUCpVg39w9MCThdohFzlgE7rlFAv8i90iKdDwiHBw8Ada6IdYU6BsJY68XCig
RLTVzKlhTD15FgncB16GF2J36EgTQ6Y2q0QZCfvhH1YJzSfyAG4fKflqJ8Jsr38X
BgMeGz+fpvByD55T3UFCcGOBjZB4BZ2LMpjwUqDB+C6psyCJgvxahXnwZqWcxCDE
vt/eaaqhVYc7UHZRJ3l3AjVW8PfdBqEvcQ3Ui2VRe8rcTgamCh9uRlIUd8VCKabP
apCmi20F0T5n1hXOpK2R7uo2GPiRK7fvCazThnYYgcH1ow/1pUYw4cQ8V7qzR/yb
PmdIPbo0+Bkj8W6Fz8WeOcFn79ef1lh2wSIpkjiox+DbG6OKMr9jCr0qvTxnNoCl
4IuJ4bt33fS924SIVBLX2Sm4U6oKIWnS+jlMaoamF6tjvvim54FxYPv55r97YUjg
OB8SZ/36dP8k2gYhgxkUpTieCX1qXywNVvRtD+ITZiPoT0MwE9+numppZpeh9QT0
P8s/NVAoP+Mjj1kg8aJifMI38Epb+bGW+H77FDigsXn66RAxPcz9o9ZJ2z8f422C
9UA3Njwy49tZmGtVoUWxz4kpQiE2qI7eQStCrfqWyC4GviiA1myGEVDSkPOMkbVN
8xz2PF1lehqZ3TXw/nAwggVljVnPtIiBtPO4lIRmyz6XnrrMvwsUdOkSqJwFxGQp
a+2AuNUBsDWkP0Ia8CtNHx6fuNeGqPYh8rJIiQiB0BD9FbZU7JLoFWPjqA7m4aVB
20o1x7PZnTBX9tOWI2huQBSDw1kKADf9Obwx+9fdymDYU8/QVo6hP88XsRpWjrpq
VVcYo+VAiuHGTlI8dCCQnBCDbTArt/eq9P7KA3ZMQPK/B39LbzI6FN0O0Zkra4mc
8UZWFnPvoO1Tac5hD9oOwQOAGWbUMBKH6XE4zdK+g8Srhsu1a2iUD5QkWsaFCLpX
DzpglnxVPAfSYkvWUf0aYBG2OjVDvUmaUCq0PNMW7d712GVjWiZpdkxULqqIJEP0
uu5KSawSlixV4JyIHukApDoVqnzuQThkAUksRHbai78xB7SptdDIS8CC7cGgQuSC
moDelBAaRrfJ/nguXj0GTYYCnlVGXKvI1rJ1LCq1nMkZkMRWCIhntHxhseFAh1xA
+yXTgzu2VlXoBSd1az9pbjg6PmfX6bVIpylF58JNjc9JJSP3AXRx8/v4zbfpWy+p
kGspO0Ds4P4RYS/5ed5zb0EWGVNDeq6/ZtMjZcXm7epb3ajA9wIB/bsSWVG74F0i
FiR2Fl7/V0+4HXRmxBL2K+3yU9mxqL8+8eMuqX2plF+xIvicriLbHvi3ppI1jKBp
wZt/n2P5CM1kEp6+nazdvIQx5aPSCZP91y/h53Q9I9nBr+kD3BKv6H3BYM9mSiEn
EGYEPFMeropnLQxlIYPzbu0AdV0laC9/uChK4LfO+TgB9FXR+gllOXCFuUO3D3Ye
PBA/YRd46nNW3iBl5Dzfu+M2BmZK3ox8bNcVdxixcLDwZlqTvApDzNH+LTbifscW
zMoKNR3daA3WRZ0sGMVsJsymNHAQEH5cmKyEw3XVA+YQAsPPbQ6E8H7un2N8XsXF
ybR8M3Uahcb/EyY0+kkBU5GmMpniHe0nS5HhSctm11mq0vx6UQ6c1K6z/AsvJYGF
NrOTJiDdvHn6v7oJ0gtJRfBPCy6k/XqzwX94opZgjaZJdy6guvl64f00xHYVOSR3
IxGgtJp1F5nOna9msui7HQyNjyr8zWHNkk5V3FcMRkJKKimmqNYfE4lHs3emgtEv
1m33BxgmOOBSF+7hjLTVwW52qNXnCqTt30VzlmE9RT1aEUSzix/GAfIP2xv9AKA2
JQhY60ueK6OGn2S5CfyH46MKSH9JBGxkHUoflafr6RuZBQ+Ly+I/Y5labWoZ8aVQ
bf8QHOJ3Lgw9gzkxkZYNaDf5mcY0pAZYNu++dVRY0LXazC1E5wZ02pR94xxVNgNX
Km5mAeDV8LBERlTDjyLLolQSg2zA+SlJfuET50epYnlh1Y7sCF6jkmGrdPbbA2wt
olnk/z+K0p8hQLjZGaupX4QnQI4frGO0n0wCahcJou3c+O4FCfL3J0TAwKVfwavu
AQsOHMDKEMCENN6rIgN4PFaAc5Z+AdB8gT73uBh/zuySX/ZNofQ4VlUlVyQZzPmP
RNqs7diMe2BeRKH+LDT8SFrPktYRHO9RS41DR4kFIlRbhclKC68nmzmBFxUeoz3/
A0fxmSvkuLI0rIG4NOgGn+5NmRva3J2aQybRQM6NiagcicB5Q0Npmlr3NsNMKhFc
ckI8aUbnRN/ANvEDqxi/ZL3cFL1EL1rPUf99kblBY8d8Q0E10N8eD9Zv+9b9NhXD
jw/WoBr+L66B8YxX+mHEjzFIewS7Zh+o8NPwlVcj/VVyN3+MuLlOI/LPPYXly/Ja
J0rAiBc5WsRTsiAflRpvFN939TVMbGHUKpShPajSQsrvzjZ8grY+56zIAujL1Nn7
mPCqFJT71RFTIVE2wAjJJy4jRm3YQld4OCW82L68IRSde4rRV4GtzTk4qVaAQwmL
nsstjRTxi5jdUaaGu1i6m/uSlY9WDkTqTrb568TundtizE9RMVMHBDJ5ZJwy3PxM
yrXJ1zuMmD+ck2RQqVsVpmt1W7Ak1O+9N9W+KlMua+D5z1xg00wOL7zu2DLN8vmv
ll2GfZVs7Jg5JfHxQL9+D3PABvv8o2KJBjE/B8358gpLiyeRBiM7el/tIu933Mvf
3Bsf/uf2ZubOP7DP8K2UtSmxYGMNtESb3ZbnWmU5pJen3LqSIoCIdktPKhc2bIKt
MHi6TXN2IrcrYqlCBLCeH/ffI5WuaUJQmBvPEfewznNRxtMQrAohIg7knfAgm84G
uKwI6I/ymA84sntbR+RaIT+EuugMomFRr3CH56GM46C7s1D4qy09w0i9vOypy0TC
mUgh1emCCkEvbMcOvtOCq/hzHFJEOH5RH4f/77kWIbg/jyvZetHu45dWEfgCrVjw
aseOlLZxR7Eaj/SRebB4GZTHD8ZM/UK1wazRjeKCSLqvld9z303XjyikVpX1lgVl
H9uurgtvhYeeusUwZrWFRGHvFovMgVWLFb81mC7PVnVhTt54wc6M1bAkNDdXRiMF
RKP0hMf7hYHoezvfHrKZ1f/QQIp3/RIg+F5tDhTvq5dVfqCpUHpbrTakPYuwOcnS
j3U8FPNrobJ0N6LleuJ3Vx+USzelZQGpzeaKZE3DjJPWtOpOe6OyJas2sUhTu+4q
FgWVqP53PeCzyY3ypPbhQB/pxcshCdMvI1gzzK4EminX4vSgtK7MwRz1cldeSNUu
8RY6HXYpsoo5P97QZxGcf6UllmNZiaoL1ei6DAEOWqM8l7FsCjNwCJYVLWVI6PwS
RvnMvrLmFeEDHq5efuaFTX+n77JBT9XT3ox2X6kX+2AitFXZAeZwsBIXZ7W8qhB+
m65XiRliYYbnqp3+R7dzM0mQ+W0vEFcMCpUBN1aBSazr7GShSPaHyVgxGxe/pgZ8
7K7T6TSTq+8hQGH0ZAngXzDz/KERLCXzEw+lxt2eUvPTf8Q65lfj+sQuT3ziivW6
Tt5rFViTcgi5NIhgARd8WrYtjx2uiVeJ2r6ORex8A3zHheqmJOpLSt/6cbZlOI5M
Vabwnyu8JcXTPxggN75UYh8kmS4iYFoF7ibHvDtNSD465LYu29QlwLgkKyFAYj3T
Q32Y3ABRnjApH1+/S8vr/w9c5D2IRdXHnV7axdcIozkBdI1FmLpGtEprWL1J8izu
l6qvgYe3v7YWMXOnk0pISV2fXtXrOue7JIVBvB+BTJyas6AVw4eMrzraZh8Bbvq8
rrmfoGYvaEoW60qwIKMZBbZxU4nbomIT5UMRB09aNrlcartBur8zmnpTbboG1cNT
42UiVg2CZNhHiieM7TvXBwCfG/dCS+xxq5owcCY/ijhu3vT+a7vhiKqk98v8Ui5I
VL2gST+ewOX6+oU0CUSOJ0Ar4Le5XHALt40C45Xl5TCcFFfNCvBeesy6ZU2UZqMZ
irwKSHgPaYeL02EbvphAufSGOerEWDoGLewS7Ac45SCkVRBPmUbXtQEssCOW0Hxm
dNg5TtMH1t5R2RRjJko54V2PhKa0GCmFLZc/Ws6GHYLQar5hHXmxWuYTtCjDNj1o
6MH3YeCkNXR6tI7ZKhw5OMuHEflUIvW3vanhe0p8LJgFWlk1T+IQvnG3wndMU1os
6yvYkrEulY/D4axBQ8oeQhx6/3anFVdOwvwy16BovcVH8sIUsA1IKgQdOUFUkLt3
TeXKsGb8h3SG8pBId4NZycWhIR9EfhngRRuMYEpD44TS2nH5gKa2GU94N4uxO+6p
I8cu7BC3pUF127MU5fuWudfxcoi+moKQCtmxDrciNwHQftxUHK037f6RbBYc6fuk
84I+pVkaCeyt564INklYawcpJX5YZfwYmy/2D3Puj8L3CZNZBj6LK8q8QBwkmCtZ
jU+NjL/jqt6IIv9pyOVAgZZevW7X0Jm00qhjSpnjRgqh3R061xgs4PF5MP6nU2sB
BQDHbIBs3kUZkLrC4ns4fwoZQHmD2tdvKB1PEIl1peoq8CDtcxLpmd4r9NLrCVtW
b0Wi4tt2fqoxgKBFY9z51aIWS4/7yoyaWo28yumYyBXJ0UpcPfAbzdnGs6hTR0tJ
kx5S2bopM8AN2ieqhqdS72ujQ85RUqvom2eLcsAxjFyKxIppQ08mxEvzuud6E0s2
oWSBj33kfmq1qMKeaiVIZJsPxSPSbklsSvPU51WZ3kLR2ap4+g+URt+wjjnfPP7G
8nWSLLls8tw06E7aJbkscu5dCqueXrtHAVpXKGdG+5oJuFMMh/tD0REOvL1mjTT1
XgGYdMOjj+pTxEfMM/z1LcunHteAlKJcJYPS6eTJZ0Bx5Cq9+jfZfglW3gDfu9tc
m1WJpMCKXodbwyclLdL8veVzNmy1pEmnEFXWcxv1Tv9LKvvzxAkKnU23c2QGKxlU
I+dYnmEg4FPOYb08A5d8gf+h4nQDp3saqMo7BpBd+K214IBWLMge0pZiLgeZqe2b
/LMTR9vpKgztau7OxtSyDAHO5r9EN20z+GZDYIyAkWtcRB7TPp62KPZE3O5el/KX
7kmi3Y8iREVdri1lxthu+WyB41s1QhyD+EnfwdmCnHI7OY57URV5r9kQFwKo4/Ap
sLWh2GKz0ltdzQPz+dQDuNorFkglJQB5zSNC3IMVhCe54HUj1Zh5i324MWRVG8FX
0bH5iHY8TgsPPsuVpxJ2kh8Z6/6dKJ11JyvJVhMVeVfDJ5DjwbHn0qLVVWm1iBsF
54vxNYrdjtgI3nwfvQMdUvb75o2EtsEXjKNBafOnpZI9eKfRP6zCFtLBRbQj3lYJ
ulCFmX6FouLiaPeGwsmZcjk91L9EL7DdSi3MGoVi/HGKGn3mOKvvQeUYzJRYvs+j
/ulclTNVOeff1r3XW0UIOuZOImY6bzlo/SWWc+x0St/Jnpwcjk7yWLZIM7NPug82
D6uGo11m6l3k8/3OEcSLVExEJClxfTim1q0bXigjxD1V2p3LYUx8LHUutTBF+cO5
5VjjgPat54ZBhmoD5XaLBElXlHdJDOOlEfLQRwamIFnl9Q3cUnc9nDdrxl4v1VlN
g9g9fDGixe5VmdcH1yWLqTSsjC2kzuq2+37RP33X2TY+O6eJPY1q3M/t+kfjZvmh
M118RABYEV4w+V6uB6DyNQT1u706koS9Um5k1QQC8S4MUsxPby6ryLX8OcxDtvmm
ODs+HPolbbM+5k8N0z0dCFc7TISjKhOMKQfykGFD4x/SZYvkg8nihpKjU304i6Mf
WwHnqmALMWJde/uFSKEv2yOPjp1KxPU0qZks6G5f0ngX35EASmHkpSBCy9iGGhm9
YJNMk+H0vQvJVkvQc/FjaLBv6oJ4gwHig4xk/mAdhjRbzYgXPhV0+iqRSNVN11nF
4QtpP5OiuQ4eshV4aUgB88uRruVHUkf4xl5u4tHmahX//yLLz5PYyC8CW5lw7nc3
ewFS7gjFaso6wjmvrU+T6nzcIW/Ugx4E/Mb0Q+U9N91d6n0Eg3hy2v60GTJv1Oj3
LIsLAJntjulE2cY0PlLssv7wjo2ZZN78OHcCsojNnrlnf13h9eHv8JrjYcZU+ZoF
3Z1R6s3GYByPU9QZWd/veTJ1+czZUsC4r+hsF3Y/kQxeg6tF43iwsolNy+xA7yWY
fc/F5dbAqBxbziPfLc97hBF0MId9ADmXO+0yn1fg2RGUuiofNR2+wD1B1Gw33gc5
RZyM3OYsUhcf161o7U9gu+DVJuz8F9HrigO8e6Wqwv+QWK/kjzxDipSGNgWMHXug
XUGuFG6mFjwiqy4R7OO0vsOQVUwB4lgXVblRVAtPQUL1G8HDi79SRXI8CfxULPtQ
rIyaacPjizR/fA/Z+PTfAB8qd8Ve9KDib58WrgH9IX1IKZIH/50/YWYwe52+RRNY
adU3xkIaZVleCjPXJ1/C0qlRw9uwyTr3zK21SDkxr6pFAR0WuzZ1YhfBOGjLrb/4
IImUmb7nVJ3d39B9KWEbxGvyb1QCX7BQVFccih3VzGholv7ZzroUkudEwvaE++we
wPbJJrZphau4s1dQjgBvjIH2pFyk6WsBeiP1dO0cjhVpwBkrHoFGTI61fvbbNPH1
swsPALVoSIwfa/PtF7QVCUYpTOOeQM/k/AYmQ2oJj38mU7LF0u6Zrx5KCOEYFr/4
ntEDhQ7r0byk3NzkGajiRMuaoASXBBqqDMbS/3O2ZJ0MfU8/IbuXnV+1mOzODxq8
mFkUOYeWI7+N1DHhzFLtGIFtN3mDwmwgrKmJ/iD8O91Rt+tAot6q43LCP3cMX3pw
/d63Se1mfpppz9WXoccZDXRyLKNjkSQXahGdSxkuRWNX27tP0OdWoJk0210MQtGu
5rLNmyFIhG4I4FaGkksfxpXCGjrKahkrnwL7vNai8xIju0BgvDNXwv1nnN4KQXRn
AwpDSqsEFpWi3ARQCTsm/lx6zM+F7IQlyQ+qVp39mWybt+uwPF2G50T36WEurnFL
yFZyyF+65+tg0Xy75Ii59H5+cfkmkFYw2x5yncZ+weIDB9AEpP4pHvPYKUbAjuEK
ybx6Lgvg8dMOZwINxDkNxS7tqwZ0SU7p+JsH2J0uc6WfR3/0goTAhcNczISx0bLf
dlq+pd43nQZ6cEr3khivvPDuPw9a7D8BL2Elpa9AuFbjHTo7wf4AD6eKJ53nVD2o
bxXpmddg6/oUBNSAPWTztbuPr1RxQSy4BAReaUGuhvSIwEJ/1j3zfCEJLwT3HITv
mnjZ6f7SzPeAt3cVfqcpCdnU3P91Xuk0o7OW6WK5RAq20DLCi1dQbeXy6OOZccKY
c08ph9X/wuDLxACTrMq801l4GJqE7ttpOW+elwXa3i66HpEXNWPODCIi/OIbzsD5
1vdmuBokwerhjJnpy6HMCW96Loyebu0a7oLzihWc2djDqJCJVaRrV8OEbr8dfUVd
H2gz7ykQw01caMZggNhAZ+gxRIiJmVW8JTcVkfPoq+pS4Lz5zBPvFHqpL7ENawgI
Exs+Ml+lCCySa3/buOwQb/Eh5czk//rJbZ/RTE5+oRVXOaP0F5B7vbwIea+8xn0M
41PHWXXNr4leGlKW0gtsECme5VaKhwF2/YdPl5882EZEMLu1CdSuEV++3UjouPko
V+YqLF7iENlcdIgrZpk23L65cR8vpjAXehLl4Kax/njX8tjV6rRElh2WXWq1eETg
zEOZxOIYIY1Tz930xDmLFPQWdevA9d+krUyoXFnXnfkkHUQ/qorstsBa/XqEScfr
rwOQFGg36+uuq1CZZuQat7eCAxE+EJXOJSusjXI8D5VfEF+aTpKFGyGiuhClQyij
xCNyqa8bUg9Klkb+Pj/JafuCDw/GCPKdPmiuo08Qnu/qHPxRBR7ugJLDapoel6IB
p+uZYb7PVLobuLcaGrm9FN6SSgEdCGeCys5tWeLIA5ppe0KJdPAinSS/VM5e2W2Z
PoGiqMoGTe02/O0BtoZDI37cAdmca/MccFrJCHEmsf96di+HtI2n5wIDCHjC2l7H
sRt+xzpa2ZbbbNea4Mu8nI6GPZ3oNLtOIO6xxIUzzzHkG6bJfFVne0nfkXDF9JAw
R2MjFKL1CTTqx5jwahZ+o3Q/IVLaRJtlx2IfrauhN6vZn5/PAnymJHLFoqSVs/Fa
Hkz7B10hTsgqSwY7oGGqz/Ndfmotx3KdpbFTnP+xw9ERArb/WIHXhLlEo7XzYGuE
sKuQ9XEzLUWtdOkvou34hft4yrmCBebCA/g7nB0TzwVYcDKwpIrXIwy3/uLdPEOo
x7FjcrpfrKeXRv5GT0B73PVfqOLRgiIiZqSd2ZJ6/eznDpzEfP5cTQtvqOjQf8zp
8HTA2ihW+PmglJ0OX0XPltk6IeVs7wXlMSA6jtLClzA2WLQX+krahGNLH0T4gMGq
qIRdlH/KnQsT/ZNCW3M6TPZHQlVF1KdQQhiwhOh/KvR2AiCEpnRyU19rRC23AT6c
PyRiv5gcvNmhI4BoklntZtvYzLYzbOaHnzDhZqmcWf9nJv45hkOUaunNTU4lCiAA
cNug++VaGkwkinWol7uX+6QJN3THjZx0PfsLnDhDEIHP2IMW2rMC86olelyA4RDX
/QTez/yzmFcsGwkhyGt0jEhWOjahmvxnMjYf3DP01ht9/cn/aucqhcJuTRIkHzC/
Zc2k4xbsTPQR6VQ307PtpQMYQZchuinZnavpEBI4tFUNBZNz+eUipP/zp0yciTLT
p6CqCNy8+u4DXVTTZI9NlJPs4f5F3DmvuMNQrOk8YPFnRZwGJ7+/AO43yUq56zK+
L5o7NvHFPD7xCLiDr+y8TbLdr8NTPy63Uia7dZahYVdSgR3IAXaSf0WMIOFfWOwV
pkoZPXYuhhFBNgrtbh6hrI6SZKrjARA23keIrc3d1Mnwsvo4j2Dk3VtO+vStxGuK
JslZ9t4zWv7MStRKD7DSzlnPzaodZVWbd3Nx8ayQxEXRzgIlEbjoAT7XaTEibsWF
6i5ltC/P2W4DwSOrj16V5ywYQbdwiSgD2513JyDUjgovQKk3Evy4xN+rp59qrxYf
LirX/48kd76u1EOb56QPUNLUpZ86330kblJQIUD/Fz6S1cBv7m2Tw2K5pH/0eCi9
yiRuiaK2kKDGF3eQeZIXoWYvv4kTqKTrrF6F4Krt5zV7gKAtwIYykq7bJbPwhaCZ
iEAIhDTFaevv0uGZ3aLmGWRJKoMa+ZIbVKqH9vqg76aiXNvNvPLAE7kNWRokDYeL
Gji1vBWDTw0p9OrwP2qHOQSC5zeapPiVbkP96oHtzwNuxvKJ5i09oLKgTM+6OgGv
wA0I+iOh//qnDGr33dq/qo1cdZy4v3akr2ASWtU4+CzCxeLc1A3pPJWtFB2iwwmq
G1CuupincHG1hYN9mE9oX6PlIJlarKZpCt+exulpqf4/Zlkr67gv8lcXJVn1UVJH
k5L0rwEXPO+I9FQXLXrP7jjkN5TTOhkKZ/INRtcTGCKqG1JC8yJkHMDTss0Kbh7M
F1rp8JH9ht4QBqEK7jZ+FQAPEBdXA8r9tOybusBBc5lfkRbYE8kXSI/qIR7Csz1S
PR+gxKiwjqsYXx4eem8Ws+SG4qckpkJHAdk4nn6FnHOEXKmBYdyV737Kxa3NTEMS
TYuBpl+rMSwB6e5nYmF1K5XNXPLstNGx5b3O5M5pAgaczxEgVC41bIJGDw+GtY3J
YUM4+Vovz0or0wJkSYRBtS6CC0VLOLMWI5TriIX8sV4OHxIfK8a4kmfs7x/+roSh
fQ+5iP809v0a2/whSTQbp+asCbo31Co/lVujeqpvbna6MbYtItQsrJuNrD/fHdS/
oj7QMApQQAou12Hfp0yjobSC4FGV5pimE6VquccLpITePRT0KtDyPCIvJ6mBw7ZC
w31/PK4vmyxPMrtS2zrNhihELNIcGMBfkA2aHwcxfeN5GZ6IoTGb9+t0HxWUfDV6
r/5BJHhmvys0ZP4Lderr0REXYqhLJ6munAzSd1v2hajyvNQgwgGkCWbIR357q3iC
WPLfAfxI+fmE8FvJmsfpZT7jWUL5ueXOccSJEQGdZslVKYIYheJ9CsCZhPvvjolg
M6eyxrWYJxsWtYWq/I/v9vWFo8ShxfPCuKcc5k/2KsjmTFC3egXrAfsE/NSpdc1p
sN4DZsXwmAYktfNopCmFCExXGDrL2YQWLyNOqfIryMMNhsoSy5rTe1BNYY5Q43jF
235U/fQnSnQPy52gZyXfqoDgBVXSIlzdLXGGbDu6TPy4MQTrRif5SXDJiqGICzpq
NFheybr5JsRIs5L+MUs+kEqzdYB45svlaedAu54sTKhI50jmlSVR8xK++y88IFLI
e+Tmzm5LhkX/lSuyAuobNMfH1yVDAGoiZn2cgkEQ2X01K7wsRnUZSVvDqL20/wHn
BYGroIkfmvg/hhsPPxPTjdiON4+dUdR4YCTPEfnCS3IJ0MQmIFDqQdm4Gw8Ep3Qc
RlBM4y1utX6c3qtyqcLLpZeHhDl40vW29zm8PxMz7jecjfByjc31LrYdh1He+QZs
wRbo6JNP23R7QQd2f7zEAK1gHOL0vBxhXwwEmCsoE1Nfkb9G6UnSXtH1jOdLd1B7
dcYE8o4pzJQTF9bNhXk6jU6Lkrg+9dCedw7y25XK6ywrnbKQu4tmcSgsxBPhOwww
pKGM54HR+2XMVwkenN2Hs3ZEwUX19HyaIJPaw973pFWKgT8V0kRccCiz2nxo4aek
X7+rSCQGFSlFKSZRi6BN7Xtj3p5LWBWDsnwm0xkMUUQ9DXNuptgfgi576y2gOx7j
kZJggzKPrPtJv45mn25DhnhXcVe0icgGZjoFiyViGJXJj2L2qeBHzn3bO0HmAD02
Yyc0G4iv1l05kr34sUWX4IkcHWyU30VKnnvp1OtIROdLT5em85VOWKDHQ/mmhgV5
aWGMSA4Q7U3XoxOCy9eEk50QdP3ibFEBhYJNVkMeolj+7YKJYZhmbcGFhEB2BuCY
8rIXUyU52yFJ6xoldCr/0/erf57TDytXnZph9fztzks2JO3NqLU38niBSdU1LfOz
ZpDIEfehYXrFFzl2ZMpaFN2arviildcFBlhkMukOr8uN6EcaCb9XcDryfr0PghYJ
iRHlwOc4RMTuRIrG7rQyAtQ5EI37dbLkyHUhk23GH333k1HphMzX16Bbv3JpUexQ
BkqHaQemLsB8RO3kwlqLSRbYPybh6iGrBhd401DcMUdwhv5WDCK/e9ZO6Tdme44d
K46CG17N3DEX3gMa6w6+LXRbZ2ke7X097k3CLuEHlAIyXtrK0zgzJktBk+iqqLQf
26AbkAsnrNQPBTR4aV7gJfUU+4Mu6ug4gQrXr1q9G3VzqrJApn2+Wod3EcsV+AmN
DeAYA0jG2TNRmyIw/AV2c4OUvATpTLQAl4bFI8QDyuXq5Jo96Tgc+APm6MhWLyTS
4GWuh/qEfw2+3ZPRvw24FDLgv3g43rNIfApe084y2CAMP8e8UGn+36FUXI6FLug5
mR2C7omyrA3v5JSsVlwuGBm2mLFZ+E/bRMMKkS+A5q+VrHhpZ9iM+fTepoPR8avW
WyFzMdTyHePWjHVu+4f/I2A0URmXgHkcGyPmAni4IcwBiD4NnSlxqTFM++2PFq42
byM+n2FtL/dZdYJRRuVdB2IM28ODYRSozGjZgRn49GZtZwXeeV3Usp1rGULYf9yo
aEcBJw3NejEnoZ5UqFWzu5taqBuulfXWeMDc8lUIAb1Xg5FbvOAvDMpq/au1Mu9I
2nCSsY2Cwwpn6VpwwPjaAGX29p7GkIn3AiPi9CkfXyBT4I0ynDLPM8N+1m8l6wgf
1uVzIvgcSo9RlfYHViXAkTBZvneUcIw9mLFzsQCCZWp9m1eUJ59jJEyVeHyzRilu
Pp9UuBgk+ICBS8JZGCw7E9ao50NmNO7XWPB/dBPotvqmEM8QRrKlyiLH9SGk0k3B
yGriVmjAxEY5XjQKJEoh7ViKOdtzCrk6MpjKhEhOIFYb/AffPrQgdyEf93MOE6OR
H8v2a3c49TE/wMFvxSuXhCVv/Kj6dkr1K7FQ24GYiSMISoY+PJohWkV4DQGXyO8s
sNCQ14qj6bUCp/vmKkRiwa3wgSaPxZ6S+RbWzdXJNnPDeDKt9zNRuFEZcClOncGv
eNwjXJv+eV0I9PQj6lSAKzIdbBFj7ow/9dpEI9fG7eQkUoZkpoV+Ive0FpsYTnwM
Ytq3hWFPlu/6n0amSazCmHBsXvkvHg0ZLjAoezwtDdGgHjVhhtmF3+heAhTAoFTa
lE9bLvJCdM0kY+GAwUh+jpMqaEHKJhefvQAIyphdVVXtXND863dhniqDKgXu59Es
hsuEgRyCxB90vtnX+x/c9l3EzefwvLpx2C/rxy+tVBbJ2B1iN2cIJSeuszu/rMLs
9rBt+nzpALM1hOE+0qujcgsfKROJBnO7gLWSSYkJe/qz8eEw7KORoRDXJai5YLe9
qsHvHgTdmbAA9OaBfLZGgox/KKAA7iw84d3SXGiBE3ltu5y2i10yb5ztdiMhdlRo
XNDL+ocDAsBfiZwxKu1/N+ytu3sQZ0NpXPc8KOrREetMKYBtjdrzITDJj+Ne/yLI
FO2zWpafyX5CAva+7ZKgSjC1eQgigzPmSFWym4tw8cA29apfTxZG7jijjBcELTYG
G0V5ZRZCAyI1KAkG+aSU/N8mndQUwlcimz7kG/tBGk/g115ij51oG3k7NM6Smos8
A8xPyJWkyZ9layH3IpGuMFlKvUPQi5gvwzMZhZynOySEO0U9/P3u4WRqqfYTNWXA
yEabJnUaNPKciYzRAEl6L8MGrJC2+vRvO4Dk/felellhrN2EJIHyNuVM+ASAy3gY
dhE/nTsj0RiAGtGu2ASlqD7vyLP2yNc49aLNleuo4pUcwESpTWPdK/CUbez/MRiP
fD1O2Qh2LL3h5ytiXIOoevuFhqyFx7PARsMEw5V/COGoHBqKXKAdhC2Xqt+rAtyh
jUqCNAGQHdiOaionR/1hy8A8q1ioQdsgqvEw5UqyQGngXXUm4Bb3zYPDzwGIWADm
XuGj9IXr3GOvMbFsHCOTyV7tkGkKWzxHB/MXFXXOj+SuSs8OV2AP9SIOCD3oeKdy
dkW2Mwp0j+brN9FXemRrNSf8IP8RTY5NZat0uo/oSmktCyYlPteCMvzILdRD3WWM
LWClHIYJE2Dy+dpsf3+Uw/0H5CKl7JFlrFZrA21bIWScNZI3Enr8jG/GCMCOjtYA
wnXYmjvq8YCC9J4eF5wHKnfHaWI71RveU81pjyDHpnDLBe7vVEKNp+mZ1G9YObQM
rk1aoGuOLBkTkTpWm3iWQR87IFZRl9AN40yJGasC2Voe2cPmNMd+qA0grWljYI/H
ZGez2nC50PnGHAdCyvMisYvfSZhzxLuAb6LTNIbz6q2T4aLl0IajTW6rezeO46Kj
qSbnTk9SQCQtTTaOe0jU6H1BQNUVhOXmprN/OhipDXS8tRPIp2d9S/c5vFUm8CCH
/a79vdOtLFspZgJ4grtSy/myVdEg1PTShfn5ptP86G7rIWMG8XDatcA+gOBxTvda
Fjcq0iGMpjZlpt1gdMJNOY/FDT0Iy/EZwVM8QR1t8y4EbGAIfNcHxSBydJiVX+IQ
etF8U6QbZqaa02qfdL70+mRFHeH3naS3Dd9Qhn2my1AKxCRHe4xCxNNKIK7npOMA
ct8l6t5SV9gfprPKrGqjp8U2MwESOCvmnOFQYMGQDRgewKc2IfXJzloo2iHQmvML
a5A3+6xMyfOlE8Gr8m4LNiU3lz2ANpuTTdBxEpwiwd6po07ssEmJWy8MSLEqih/i
9q9TGUaAwNfeFw4ExQFPKq9VXnZWBEXDrUQGXMKnunWuvVNeuzCy9ZM/KNHef4y1
zEKD3Vrx5YucqDQ1Xs4Qc31Jet+xlcEWUx5snFHIgnbLu92jWelv7+8qgmWilWgc
xM7pIkzmh9Rs+XITLwNKJet/BVYF0KvDWr4Q47241NvZZBsEFEmg5Vc4gvle38+3
LcnZQUrEaPBoFyZoqkaY6LD8qyhBuNkAUwB3oWbNQ+Mo9OZaSZrZB8A6d9SBn09k
YWj014+qHW5dzYXNoHRtjWS9OwnYs35jO9eds+ImNjM+t+QMWlV89TZm2lgUf/3z
xHgjRGyu7Zd8oObDNnd7kIuae04D40RBkKC7B47B+xngGjb6yLan9AyFzMIZqnfZ
E6KxITj2B+hXxgkxbBOLsrrMyVOHnOnGV8IYik3D41qeJ/YCnZVA8BRX0u4sZPjV
KGtY9bOWcMjuLSuNThP4ttdZJPQQPfp+I8tIZfGIxVKZtGk/kyOXpfe6Xl1hyB6F
VOGpAuNUZAziLN2zREboSSkr/+OtTYZNH8UXy9Yfv/zb9V60qiUVkYzolpuNHZdg
wJImOV8QKqcATrpFmaI9Dnd69XAMfBsoDCu0n5xrYJRMTPfpZy49xdcTcblI/tlN
D7ZU7igCCZNP3K4TWRpd67x8w7/iPXuY47Zxy0zYh07SYBQf7JZYy3E6z8QAKzyv
B/rcxXLdUDK5GvZ9dCLnvZmJ6pkPKcBTYTUrbu5+9JGNtx9xu11C/pqgce6/uIO5
n3a/0Jk1w3y/8JPYwuex1XlKaoMlwLPCshOkk6MqX+VUzgbl+2U07rDaCWldjKpn
UgQ4bv2bHyv2gM/KCOR6wICbFkNPzHIPKwo6/AsDesapWm9HEGxb64SxWQ0feDOT
MLdhw8d7MZBIUvq2HTD4t5zP+bmODG/M8ni/bD+2eXdYJjtVxdh9zWw5XYB6eaiM
DIaCPaR9WZM0gvFuFZikC6K5XYN5JlivRI+tgxIuq+PECe2RWrzRdhWBmvI07sGW
fjACO+LC6QTFz3nkF9tbkE9qQIRX5mmumF6AQKsDMD7nop3fkmE1424Pddeo/lu2
ZXtE6yeGX64pFnJkLkEI5UdvqIYHCyesPqhHtkfurufk5938Ki7rJ+3Ooihn6x9+
1fk3tXKvRDRLPFwW0xlizwG3yzWstIvxA4ddjoew1z2wYFvvwOWliyk3wVc2ZPP8
5ul6wGoYIzYT9nacGO5+MWUsQk8FxITTszsemgL2JXz2KwwU6u+h50vafLq4S6TN
8aUXD/dSv8WDqTVC10YXFFRtcnq9J4oy1mmfCm3Dmqz/5zm4tA8z4UEPwrSKEvWM
COwV5MhttHOYfxw6Y0zqzn5pKlqUcsw79z98Tgm0g23Y6K/HVxRrWlKSjjphy2NI
JdOqubnUCCWDHrHdwVdII9b1SCl5UQnqetRJbKtd20B5fUVSOz3yta5s69wAtNPK
U0I5H1kDNIj/n5NFmCPDi3U0HRH2t4/XpzyPg4+vnfGu0xNwV5TTRAJDKmhZnV6F
yOQ5N221PalQkZclxXjAE1kyYbVi3Fa69AjZezuef/+2dbgehhQl9V4hd5BKua26
QFbk1H14gOuNJHQAToR7I0kl1eZo6+rbEMxmxkgdhhf3AxCL3gCuiAErCUy7OjCa
W0WQSK7TO7HVQnH5OvdQOwFBa2pV3rTMALMn8o0fT2AkWroPnN2OOi8SzAHPaWfC
g52OiUa0Wy/X2R7mFnXJbTb67zw6Hx6BCzAi708fA08dNWTuYhwNyPqFwM+a4/cV
3ojTKTRWBKJQ8TO2QZESsUWBa8J2T2XOj4VPQiCNxTayUSnS7bdic1c6l3ZVMkIx
mTJMrUgNmjbFzvapGQ4rhfiXaP7jtSUmW5Sjf+gP6aueEPJlGqYwXZlP5Wffn3bU
auP29rvwbFMrYgDLcnZ5w/1TCzUdCy9t7IUgdlGWandB3vXNVSK17lKZzu6lJngm
XKcKO2d1clW/dVtBNwW2RLT4HQOc3jeDe8X3WcF6QjNsvHJNkFk21tbvKgowjmKK
xw4QUIvQHzbn+cOjysP9BYJgRABl15+5vRb4GOXcZYHg5QhOaTpfxTLYu2XQ7KGU
5PNiPMbA0z3cXsuq8dDJ41iwjNaGL84fLMWrsg7meB80aNuUWrupVKe+tqW2HVp7
MmnL/hum2wPh42T3Wfr01BoKt9ius/sgLg3olfAzuFBj0XdkDNReoFXw20D2jTIc
E3vg8EPDQaONnnvZBR8xI1RMOHvf9mkqUT9e2kvlHdCD5+eU7ElMrmZHvN8heVeX
99DbN6rYdyfhvzLkrCqUs8L5V6vA2Q0r+gcm3vq4IdvMbnAL9MdJ7V6Np/n7Walk
rwEry3w5whmU+2RwYN3+jIlOpxZ2zybhL8ITmxjKJGhkJlpPJIN+sRUqjNXVSdUU
HBlhsbAKDXtVxtVGUczGxGI5dhRKdWaMljdY52iAEUt7XeUSk8m69Qay2XhQrkBI
5tGrXYUfMaEgVTn6Ado+GbqWPYCskKPuf/LhbPLIttgLlc5+Ep3VjRJIa6A1vGvN
93cBmdF2ZZvs5irtSwcmYnek0EkSzoajs+c8zBRlzmQufJkCZA9+9Yia7aj1Zr0N
yCooHL3lEtRviBszYNfpS/QX8+1pTsRhQNi6qvK/YHN6T4mbrq47p+Xtx/AUuMKb
6AWPSlSPak3EZ7ewm2SWjuJEBkZeOzUZloOLMw+FQo0aj77RMq5he8ClsL2sFGZQ
C/C0QBAivQ0khjZXFz47b7k080xGKIOxQLFMKQoUX4e9yQaF5H4c/gua0rZKbPJw
2O3kqeLmRYGIl1uLV49cP+7/elZr+WNEnE1pLl1Y0UTM4eKtuBCOMDsL5U91DMN2
ATuRmnTFGWi3Ejvu+0kTUfPNAxybNt+1kANJH/8E3lvME3dYuf6tS6q5rm/pVXfQ
D/GY2/EdCXBGGKp/MtM5iWkrd+etlrSyT2eZiYlWd2I1zReCPq1gsiGRHsxOyl5A
Go1b4tGvd+r1jElKjZ+Dh/6BFOVwwHv/zj6RIugvIdmyjkDZOGjIc4ykL47HJUlO
nXLJYp18JrqBAdCQUAxMbsbZd8vgUKvjNdKo2XkeVxaKwiwPLXNinECdrAZu2HGN
oeuqeC9HMbF9TECFFvCND/O5XHl71qOxWRV/i3/7ngp7P6FsP9CSZKkG50tAyMyP
4gnvo08T7qEzY89AtNFlQuDXvtu/GgyJt0Z67lWkL+Io5mXgICIZ+g3ol4GzF/to
YcLmg/jcHlFXOSj4crM626kEyZ28YA37F4iRVwbTS924ZF60JA4ZYNSBOjanmVKP
mrXsKfbd34GlDuaihCxz4QBU4Q4E+PIoYGBqEbOWeKYQtXlbMc80q12QT3pEda5O
963rYPPUFVAG8m/yf3a4pkYbl2pmqXojOxBKheT1HZjXiXLJhYM84kqoWB84fZm3
KO7uy9H4nbE6MA1y0ShOb7RYudqAxsU6zagkAwhPbbIYj5u8BkyfqV2R9+oW+e2L
ll/m9RyN2l0wG1AA4kAO2Ocy5ioLQlBvXPOrCEFb8sI1e04RPb3egN6mlDOM2FrA
CGbdAhJ05HR9CX5MSXnp+uR29PJ1uX6UowahKUFNxGsr3UUPpfutB+Y2e+2WXd2X
81n79cWvoh/dDdGmwYCLwtYenvBfuTEzC6ue85g9uJHrx9h9PkL5YPSfltcRyq/B
bvy2WrXInfvxQ3FdqoMVnMEscgUxq+Xyy2IEOWGl4dw3mfVhXZLP55wY+wdYWZV2
ssm1bRoa+QQheNIqHmSMLHiMbqjY/drBhsFW/MvV3Y3u4A2UBE1gwdQi7iqorLbJ
HJ87ZmQKXP5IoKG/b7RvOLdiCEcdG3b2EXYoqqjyjRvCsSZtvIRvTGtGm9eeKhNt
KEyVhFn8Wp+AEDnzswXFNt/HcaxmhR70k3Mz1001eqz5sirP/oQAcx2SPm+cCBca
7uhtT8FiGaFpmmkOLeBzzp11eWvyw7OUGwL3OMsDavnoJK4qH6Wz9HCwAVjbwQjF
s99hlTHOUghvlnHp5AheONn/3a4PCwYxhVsI131D6GmPti5XiZwOdq8WKPP4aAP3
Wisb9T8ESijOvAVHwqtV+REN0R4xwXngCiC5B9XYCoaFzNiSKmZUH8lzCyZIIq3L
HYzqW2L2e4PkI6lg51seAwX/KfnFeW9Y3L3TbhTjiLB/7JaoJzJdB1BSPHuavfNC
wos6lpcpJAUDGBkJ71aauQFgPnQgVR46hIJ7Hp8B8brXDyXkJKiV5LwHlrFqdTxl
2VeI8zN/2MMHJDMyWGEi3SJ8jdZRfcn2CJC2s4I/kdg5W6jjV5XOeMQ4w1dhq75T
8xkx5moARaRkjkU/OiQgEozHyuyIKMHGoZjX5UQbuzA4Cf5tuYoByKwuUMB8q4Pj
yUDnDtK6+qBiCG99QbVa6kv/iogzKh3mp3ItcxX5PfixiXQcPTU5ID48symyexm5
maYz/qYuUlWV4R1DE5tiVRwXQCAhPFiVOocPthYDyOE/YQTiIfm+k8dHKmCWADHB
L2tCsOyei+ZaBN+Xbgfa/ySF8dOJghVBxkfKjmaKAR6jiHXpMc8+XEoERBP4+E6B
6geJ98c+bGQy/zOuKJh61HJwGdyqQmra6udqQo+DORiw1J/RsRkWwrSoSaOgG4ld
ayrYL/4OUc4l5ycObB5vTi8vBIj5Opo6/eFpKBAZ4SZ/applMi7oRE+YnNoM/z/N
dfTA9tZKCkrXoGS8oYMuDKIfkIsTHZQ4hBHZKb6RgM6RtWJywl4oCpXHNgdYqYRR
4RrdDOyiz56CcHOXZQSLrPf6aLsoXv6CeIZEfOm40Dh782gTJDgtG6z9/fvIAsbP
xm3V7njWnlDqNsZFkRLC6Zjc7zoUhQPLW6kJ4tEjl0hjs+6cjGlQ6WFGvONYgfqP
cY/N9SAOAaEXknRCyMt2Oj3tTJPvT7q/eYMQSYNI6jqKJLOToiGdZUICf+DsjcJZ
yGpXlaStnlYr4jDuYYTpQ1LIhvA6YIpU0dpTxZGYvNcuQL8rha9m735yl8K9N0dq
spjfvMJJjJ4rnR0NF6UUkTLrz0alPhg9a2DUiExEa9b1RVUdTaNSpnS2HwIH6Zzd
IX9jVyJyUsndl09GPxPOcWiomHjS2OTvWbP0+YXXw4ikvn+oKtabKNS6O5LUBDx3
WR23FCpf6PcPjJDpc1XtBVujYWuEO8u1GSPUpH3WfKIxpGKCDAsjRgb9Txtds7my
grV01kuO8aULAYCvolDyBaKxJ90EJSNjfSCNnkbYxzZ0Sxy9CNDGoyhktrDK0QHH
SypHFG7ZSmrVMwk13P+Wi47SKditDh5Ae92hi2mkQv4zYBoWmf9C02WT6Czt9/yb
QYQR5/xqHUod4JbMDI3tkI7Wc7P4vJG96EevdWVeTS6hFNJkuUypY1Gh9LrUJScc
jQZ03vPJAtyrDR+xUXi/bdbhdGwt22D28iCoV3abRFCZm372yMuCJA0M6rSatqc+
N8pp1DgbTyncSf04xKZUAPb4kywqIUK0Yy63twC+/qa4rQzPJ1Y7mFQ4vFQ5GfrP
ebZmm6HCYAG/h0hABoCm/rCU4F8qi0XSWa37EJU5KxtnfhLOgcQ676WHErNPq/QE
d+LUcGxYdFHYymv1K1hobQ/4czfOaGulHi32ylTRk9QN9/k+TuauM6ak5xRJcYiD
Bt2cHm5HHR1BENzQJ9mSMiHm5KGIgldn68OEaxXfnZht6cvxWUMe/npXb7WVVgsJ
TbvH9P6/OJvqxzfxDpbxTPjmuXziyCrhmo5e+1n6BMkiaQ1Z2JSMGtUEk44glfRy
pdummVg45bXXN1VEAnKPJM/LwleKFLnNOluK4c+7d2Przex7VDO3TzSr3WjxhwRw
ue6ahcQy/Q8wx8gccc0EUWHuq10w3hmJ2D7PfH5zrfoQ9J1JM8Gatn8x0suzZX9E
ZJ7KlasmfS+YuVi64rz9G2uMxyr693jmnoNp7E838z3zKdwbkeah+CbESMPN8p5D
f/WofpCZm+tSgsqcPt9umi52QJjZTo7wd9/a5wrRCeSv1KXl7nH7sDHx4DFjXpFz
IxEOq0pE5V8L4tkL3FDpFqcufUP+FZHoO4lrL7Zl/V2SSxz8PcsTwp2JVFca4u6G
9IwjeHWwEMPVjLPGjhY3GCL58wNjMoNkPJKnVE3EDOo5FQnKrflrhOYCgjwi+IBY
O2VEsiWY7GZT7MeyqelNyEI+Xfov0t6lNsNWglU8DFX2KbO9MAinTPOhCUpUvG4n
ybC8VEweS6t18FkpkPP0hnVsp6UZcxy4oRXZAF1tDtuKERFFAFj7n4YIoybNesqQ
tUI1bqC6iqMpMjLIgMfxbP15gbso+2PoB2tD5vdwfnG7MGDZ0eGSAEYPcPLkh+Hy
WBvPEgtYlTozl88MTpcG1N6DvazbtZE/Xv5RohvBDtqEGIzQ2A/dOyu/ILsHjRda
HwKSudor7tL4GH17MSBR2QU37i8Mm+oqxv491J813GHvMc9HfR8uBJ/Z0rQmE+3G
aVTJ5fQq6bN8siZe9k1dODR9or0zYytuhwBQcs39NKsGKOwxX961cYyw+8nUXPoQ
b8mC7U0MwidlrmIzQg/Vy0/nwDwB7ErRzOHpVoTy5i8zGnsisCIcWl/6l5+9E4LO
TATVYFy/BWeKodTSYCdAcyNm72wbX5aSnMoH8Akx/U/rjJd2YyToI/Wk2SB8plQO
FUpaF5TbwRAw7YDjx9c+4McyLPZh7PHmV2pjlGAwVFXLmEx8UkwHioqD0FqaNk4g
jpBM2k+y+YWLDs2jGzQ4N+0hrJbBvq0zhV9x5R/yYhetREHrITMVhQCPQgTX6pbA
fwlBMXjQ1WjM8Z7wfJkoMqIsFZ2qbQaAR2aIYMZnQYoglX5JdstHiOHXLJDsQQlb
FyIdQAs7FussM2jkoIH836koLDKUAx1Jze8rUzthle0ZGdeq4JclTgOLPD9JsCoo
gy8KYKiQNZXUe8OYlKrtmaEmc64zEC+7zNBo6/UX74ZSFIKxUDZtMZaJ8XFaBbXd
GwQfkuIYIzh7iqQaqqoLpB/PL8lb4bFc2lvK6jYXgIqCrwiwIlm3a6MIPOmUHf/y
sqpW61oZqxHpO0lrs+Fbv4uAYkgbN0ND+MxAbINgSteK5TgORqnsYzA/ImcYs6iR
4wtW5Q+7A/TStI03/K33ObjEVQzNzEljWVV0sVlRyCUreNB60tnQNO34K86SiQjw
Ce2hccA0Ir+5ITlXQugJe8HlW0XrMa10Mn3Gab9/FOya2n1PbAlLYH41LH85+mjg
riXo4XLP6BeFpkxhxRG40aqITYJUT1AOtle5lsYlyJh4uzNkF5bAsdpNWPnsile9
IKzw1dkyjU0mEqLek32lnqPZcT95rrCKitXw/R10bZLoejgvWwT6qy++O0v8zXyc
1Xw6Cbx6iKQQUCOgy375RlgSFvFfuney04vbNI+m9ZMArim8VADwCgWFsIVs1ysZ
ihj1bxevZAVQv71dEMGCICvZjiPkzMO474LHY+Y0/3ioPXBZeP0nGMz3zWMHSfVy
3ItB7oa/E6uiklhuhrMZ35eTGND5jOJ82GvEV6l4FgCnBRv7LD5u2H1dEct2WKa/
VqN/EziQInAjNxDBEuzsgsHF5uJpvLaBOY/FH4gQfw9KEuahE7fKOTLbKp606AKH
nXJjuoeGc9vPX2UtDksjjOhbkMWITQ4kj/ldlPz8xAFkSq8c2ugrjMObZtYgpuuX
hhy7YLdk5fJu0YF9Aa2GhW41mjokvuAfOreSVmoWp0UsgkL9QtiJ/Pj3HDwZEqje
sCAzudJbTy9Vi8NLJM8RPKDWLNPTLcEfxiBETbUJD8lGmy87HXR8js9xbphgd5sG
Zv1XU+okzTrFRNUSmnyW520wH+YZAE9mV+pkazwRgz5Yb03hZ0yKJmoECd0iZ9Jg
9B5G3e9QMoThdgq7voHFWG8cLMEoYtlNjUmyW7VKt4Y+NXev7Bv2WFrDnveHtuZH
JraS44ZDb7PPQNnGDC/U9DwGkAXxvlFvV4qFGQFJeHb3QfY2XFl+b33GPO8gjcgO
58gSUfFa/3fH6xQP1BjgOAqL+OTJse78H35FY/scIz/wshxFArFn6jlaIRELjTU8
b8KfYIRqqCpd1z2R3rOX38gz+6BPk9axCsNJ16itpTKm0J6Hm899qhR1r6fCFi4w
gBSrHlhKDHJNBi2UNuxOXAnBcB4hbanKlaaGYstbjeoOLkPPlZCGvCtM0KRsWde4
JOzgedy96U4HAyUtXXfkvYCixkXXug00V1xxLLaVGE15f33f/yxHKHrzNmH9etI8
URryB5m06VU3xzYz/rZ6wjPVckMXzRoleL7swHEoeBkxg227MWaDkpvMenjKfQU8
xFr7IP7+lgM3Bh6njlGYpRtb8QI6IXSP3J8o/4ioOpHwLd0oIJqwbrCtM1SXNRm/
6AkR60htoZhi0gT4tHGgFglaqH76SRoAoWRx9ptRmvBo2O83vRWh5MgFG7iVT0kK
Kqm3m7d4L6U2+2sqBz8rcTi3EzR/h/IDqVYxEUE3x7fg+BbESt3f5AYeVzMd0Dl2
HpF/sp62NBnb2CPlqJte1Fi7p2Bg3LTb0axBJKgZtRjJJ2PyiSKCdvjrwoPtcpLB
0WlyESlaQNXn5w8/e0UQYnB7PAoacygroq6T/j+q/xVtgaDK+HAIV8h1fMfFN29H
IGZ2vEPQmxEoeAbq00ymaXeJr3clK1JfJbpwEZpxiQKGgrVAiyHUg8OVu/nFvGii
nhs4YLnfOmCztRweZpwF/7iYNEQw35jzuFsEjgpkYxP899YvTGHDwEq8bXHcNG1t
S6XdVrSmUeP4y7odv1AA3gEVFWftk0lRSqGn17FgEZxFZ5M66epibAQUqT3rB5Zk
M/U49wTKlh3H1rD0Trd4jsahOghD1lRg/NENT9eKZZSEULH2xVAu2+bxC6dht15D
3rr+egGAyKGT9ZA7llv6ocQzN2Xd4ZOrd0eCL5HV40AIj7OHLVYJQ5tNzugRQG3n
oJhs2MNbraG8wXLI7gPTyD5/kZhmTSExuLAsiFoPj3Psoat8rmiMuwDfaAzDjiWq
K4vvy4GM3lJKBQjjypknJsqPwlOnjHrRpmLCq67LktFPqtK0YTuRmqyfQ77cDdvP
GXbrK8dQz0+meNVAj+npCrfmhJNlHbnWiIeMHaeszX+wEHznzCkfZ2xo57VROnbs
T236qBWnlGNGcN7B35wLSPPoK62n8ZcVCmGW70TzKGLPSgoNG+ijo549KdWdwuYg
7KiFw4SQQZC3eJps4Jx+zNLb4o4qbNNibS3nPFqGqGGJRHEW+6SkN84N7eL729kv
teekoWHDkcu+xuqsK2aHI+TM0A3JVVPfRnBVQ/ANjzWHYOk7nmKX0ygwHQFP9CL2
evb4pdbnMo9DzLXpFwVdF0gy+oFR5OqC8li1RkGknnnmtjJBvXzu1INwOTJhdXA2
Js3uV30mc+mNNDEKxZTeH5szPd5wy0YTLf6aboqJHPHrcbIKJvHh085zmpIwnIay
fK62bz77d/4bybNfY314EhaYYdE+Gn26gaOb/RGAN7Nx6cNOvO1o87KDDAHTNsUP
9Sjw3beOkaqVgG9ixWwOtBeGIfToYIIl1QkbcKoIazRF9yKGzDWPymo221+AgEV6
hFhaFpP69wxYOFbHO6yt3MoJNOKwDGoS+vmdN+O1x347s9flOjy+c2211sR3PgyI
k5z8B9ZdZWyhKUIOIICcgfxwsPcAh7Yq36Lp2MTpbo2MaQPRcuFdnlxMO22aP7hf
y9/4i3eW5cxYDmVVNz5MRoL2H05cGxCSkmdwThP7rM1lJEf1oJl6U+kL2uSN0B3f
8nNdQC5lScyY8Ct5JtPmhtLlUwsvXq5XITDu+BM+/9B/OgfL1zW7ZuZSM7/NIOZA
k30DLT8G6yMhpJSm4iE5y2+MHAz7nGOZZp2V00W2j/Db4oFz9l+AM2xq6IxZoOSU
k8K+pBh0r7dpNukCAsWOqrwZ+UAokPFjiVPaAC2v7pHlLNRtPc7hph54n8BqtQhH
BPocxsuWAZ0q/mItjhxtk0hNY6JdNubMWOx6zgO3AFEoQPVN1+esQf4H/HW9y+vW
Oz1nLI6SFL63epRbDeWBvL5JtzJaTOXJylWkDzICV8GqhESTdWUBra1nSJfH6aIu
pL6jP40GYPiOqRc70VETNUlGgUEEaCF8fY5hSfSFAgM3FL/whDC7leizMTth4CCI
zWHS/2LI6/Z5P5WRpZdzdPISpo9zmlm+MoBvgtWGnIBB3R0nzGH7QNzmo84eAOGy
OIO27GSYp9yJEMD8voQGksmDYH6mdEB92YF3u43jqlpJHq3Tk/XHNgTZFVeQLl2f
D8tK6hnuYOb+J4MIpygM0ko9/LQD+NUgsYEHQdJYK5RCGqf7l4SeiD9hQDb2B0N4
BQnSdV7rYV/caAK1fXTiXTxq69TmWRJJbyNjmIjFcIupPzOWBNORxjRoSLeaFQjY
lsyTwmqXlTRZ4FvSZXXBRPdU6TA+Bs1MRVzeEdHpXkSRcvudjLGkligbOMHQq2wn
YkMDyGolhdO1rP94Bos08nlfuL6AYhhodVPV5s0V78WNARGRIDV7lxcjc9Hwf3DP
MF2w2Pqifz1LVlFgI7x0K5NOxiVylMvbf7I75UDM8i6GfI/ow5pGPpAefkEmTjr7
TxxTul7QevMEA7Xh7i6JYH3YN9gM10Yzqv6VshYlfwvuMk8WcFpeME17E/TLRtJI
uny27zqr7mUdJyzoi6E5jWR1jd4PK2hzHcYP3jaLE1O5DrdJ1BBOMsIOnVdl8JuP
Ybi9KhRvUbOVFhWy0/ikvhO/WSqcZTo1qq/h8pqA8AGQ1hXgkNEZ8VrSJpLwA8Mu
hnTyueKOOTUBYQfydxuJuTrzZRTLQUQIoBYzUSd5+0YCOTtWi0NkrPVqfxIsvbEm
RC2XpJ6iLBco1ppgCt4agFEeexoqdvYx8y32CkmBkkrlQK4b9LwzynLzOZsSpmtl
b8nBrIndnsi7MMdp+piWqNTXrlFPk9qQk5nuhqe3iSLWyi3mVxBMIdwp2yDy7ulK
DSfWmQdNL6Btb5Z670b7Oi+eE/SqNtG8Sn2fyaG24qC1RUjdcZkoo8Nzgg0BtvHB
xQKSQ3ds1v6EhWoHsO8+vp1KOJ4Um7rX0XTFz/+fKp1NvKGotjYYYrKUEkTY/ntv
wZbVycMQ97NdzuCV2+DlBgc7Uu1j8iUqjwBNfI/Htspp8ASRmcJtN7WFyroeKlom
NxYgz/HUxd+h2IdSajKcW54Ta6pjK/Lq155NjnHWuFzvBcUsmSyU1UWYFQfASTFU
weANYuOTKLM7AjqnXdCnDxob7WJGghOLiBx5ShjfBOZZupIZhBbiyEO5zFFBYEQy
0r6vnAzlvZ2Lx7TKX7pj0I+nTR6XzJC9P44JsxLb1tvUhRzbQCobo4cAq1gtfC57
HRV22iyYtAM0PdSFfqaS6JnNRKlAmgzhgDLiZj4RN4/765Pm2sqck+5RTvd53fL4
cysH8pyZIdqaRJZfpdv10DHZNV7e6rYKJeGIpcUfUPBT/Z7XDX8B9mDUlfBaIiuQ
TkPPq+sP9NGA+4XLwa/MlALPDo089ReyJeQVTZxUa/l9izsdmo/SydhbsJGACBVx
/OmWEMgg87lAuXgPj0Hsrg159gb+nlaXXMqv3ICzPSYZMKPllR7N57fkYzdqFLtv
zMDmUzmYzNnKbe/dbMRpptRZWXK7q6AdGIDdADFgkfoctOHq5IQOLClzQV5+Y5v1
BPRZXkoyBVTmV3A3cwYmtCtTSXVIczxJTyT2PSVPS4HwSdx4Yu9RgsA5uTuKFCVH
gMkqYb3H/SO/OMftbzN2uRsYk95wBL37pv4pY1DheSx2JS1KdDtLf9jpp3+Q+ViN
ecNI++zVtV3dI27B0fJbGyKS0woujcn3WEo4rZDkHCP2ERJiY+Z2h9piUJO99Mp6
4DH/B7LTKFxjaoHGjekCz4L/wcqyUaK+SqXCrVj9QeUbj/9g48TSrbYg/grML6TO
07h7Dedr6B++FKVT9LuJMkrqHRYpu3WkXhdrzcxvIvOqnUsXZe5QBYPo5qa4XPVr
NURPyT4tmghrSZBzeDbdh5ZQbMr1j+7a2nv+fP0SE5p6/8D9W3xJ10unXeBiLpfx
gLga7AoIWPbF9lUytJfbL3lj6ifyykmdXd8++QrZqrN8CUEavPitIQcXs3QRciKK
Su9H7ymG2ZhSdPnIxhw3c0X50qw0A53PgpE/o6/3RQ6wQUxbtUzqh3brtl7pK4j3
Jj8dFm0dj31yX16Nn0FIM3aaxVgUknO8OWBEfWb1zT3nkwU41zBEZ1BnMyrRcAyf
xUOwHwHrJ0AeAqdf9odvB6l/BZh1CweRxubLbFhGznQjrmfEcxFlQ2jeeoe85N62
xu3IgfAEN0+30ulg+VC/OmJo20ITWbZu6gYQcsyDJHXOFzFXcNJ3jqdXHxsdbcrB
kEWQVQlEHpTuGKKhvNSeyOXAVUGuqoDXFrDWcsVEg/9RiFNo+gtQ7EDg2q2E74i6
5BFQAipcXTrG6sZ6EpwN5nh279GAbDwY9XAg3ySg95q7O29rjrHN4T/+Ey6FYGgX
NTkLUHTQETXecsxKeSpLHN+uy2cN0q4QaQ0r2mx7hQo9efYgnePRv610aIcxcNNK
jhbm36XlxVWpgV94DK40lcIPhWFEGmknGMXdssIVOqABSINO0AWdkahUHg9LT6py
+KmAk6VbV239ipVpjytT1tN1ye8bho8Uk4CY6LZ8DhzbuysxUxLCQZEC/2+m4uqm
DODlfAdSSorpOJolmqLpomtvlEMLLKWClCSRMYrGcO2UuwE/w4hGoRf2DtYRns1d
M8Z/Whyj1s3ljB6GDBZLyxqUNrxKHm/YSS1vdL2lytHoom+ow4DtoUcwf5M9lIuL
wX9q204cfOchOzdJjpPdzyG7FvSicYmb0Q6suwyAUIhqYqXE13CQMJBnLTQYSZT+
1/P4jyY84u1hoc3PvgvqCGUXsThfzBXT0q4/yMxp0FiU7Xbn2UDbHldnWQC82Ig9
xgSaMicOm9jpw7e+oAD0LU6QJJT5aedz7bRj7hHeAZkme9hyxmIZhl7rRPTg0zRa
jXn/uEBxLnAaYjC3g6pEIlf5wJGofYgoKJbOfWrmCMLhbCSZQFVXPWiZZrGOcINa
MiGCP/1X032gL4cp6FdZbaGVB9fTr4z/LoI1sAsWHNcZUahD3iRM5gKJGw0ufbnE
ngFj0SRBpR5jdcr1Kc5xkCqZW4SgNv26PpRVXFvp2G+1h0d3j8z1y3rIruWhLq9m
J9ejdOTSk7GMJML26PCfz8mRFwZ58nmlTe/hb0Ao9X/0W09qXzvJ8+x0WWfnmJwp
WEmiyiQ+9iKxRhSZabANWkyVmA+NkDULODYM+50Q8ZuX369hHNUlKsxjBW9A2KJK
zE8YBpl8U5m5PyFl3iwhCRUQrsw6iTYE/8dBpRtXZ8RXBm9i0HWm0dDj5Tr6XK1u
jWfw8y7nX1/sQX5wkx/cPWTd9ja6+4iJfxxYQV6EP4gd5XJi2P3LbluukTChUNx/
pQofbXnItKJpQnnChZBtRhW+9oD5nONIzqkLueg1bkqhQHXO5X+QxO9hTrNcZcwc
u7fhvx51h8677T2UmO9vFEXsFhLCl/W0BNAJafhTNxhZYqs3dN0Qj+5KPwmeGvmB
EghJs0B/YBfotfEqzBJ4CNYEefuAlQPKSf89oF3pHI1V80IajbY+0ZVE+AR+LaUF
hGu8rXz4vHJ7WPJ4ybY1oC8z+SJK6cKGIXjuBa+ExCdrNETMAdkx9z/Niv9S4VUd
XCS3ezioqhksnKuDf08/S/IDqigGy2812LC3kiQdfsfVon3hAgLxRswF+n0bEkZC
RZCBm34bAlxJxtw09nuQVy+dC3/vpqzzAaae7xkbeJhnTY8sXoidTUvvnqpSaeAJ
aJT+0BV9nyuTT0YgPCuDzQ8Q5wHuXOF/SG4hqxvkzUM/2UlLWtLCkcSez0p61RhX
uAvxEvowTdFvXbZFbbGA3U3vS4KMzv7uK3wCSbEeEP8lRePjU+83cZmeJsRYAliP
CSyxspvOWmV45UZ0uKTuwJhhglEo4ZrcmTx3J9a7gGL+9Bv2jBS11BUlM+ORlCPV
8B4ZuW98DYp43tbIaxH081EZ9drWRlpHeupJ/0tjASQTEBysDF6tLiHDlIZec12H
+EW+dcfWaViCDQdBop2b3vZtYc7WSGX0pBWQU8BW5J5JuK/mX2Fb22S4vm4RJRSg
n6pnAkInyBVr3IcALuEqmuxGo+0msWgO4lTLSlmIcWE2Q3iLwweYvwFq1gIabHOc
2QKPC34KJNGsVawkZcLgNXK5KMPB3x6NfuecrZfK7paUim82+geuJheT3OXgfGBo
I7dlHLmlNuiZ5dMEHxZx8ky+NMIKOT38ZCAw7tvjKur3GbNSbdove6dPiiP7ovYW
c0BYJR0gjoRUNhCvHn7kOVFwsHMh0Hv6sZegm/Opuz9KLXCh/9nFVCXSLVPXzbME
1Hy46BC95khVwVUINYFTpjhqQOYzomihFZIK4uDe74l7YGt/bI3QKHa3ZpZNQnB/
r+h7RJc1qWGqrIBpyvcHx3jVaI4IEKbbW4MIvddWX8J1YYzssR+R8c7kzLrIiGco
vH7mYNyz9HpG7d+GncI6UrWaR3vhFu+MKkAjPqFixObjUsJ6wkKyOabPO8gUWSGo
bdwbMDhNxr231nMPMcv8x+FUQ9ONAlHFIdKb5gu17T7GYIF1BcPgTmiy+iZN43DF
8rSf08MAvpYDmgdJ6k5J5v1EPNcV+7HqjZQbh13Al+vEVrWiO31fij8I2xJT9oRc
ibYmSnaxm+u9iQ4dqhjYS5GKE0OYg22/O8YprojmxkCjJ7f1Lr0W7l0/rWWbbF5B
43N5jbFRk3CvLn7k7H1O6+MXeKZ7Cb7taMiy2MNWhL115g4H97Yx53cyJ93E1iUf
IclbHCtJWJ4U6LsAgJB4X95El0Aclo9XbgSLiERC23f6PNF1AHP9c3lPioHh1Gxm
ghaZPGzAXijlZuFtRVe9caLG8AhBaOtvEBbYnHuSpw8HuxXX7DRKZHXG12iBYAwi
DupoQRdMfE2fNIpn1UX+soFLdmpuYFHm7e8/Hc/TbPU0YUmpixZ2IvHj6/PyyBro
s2eyVx/pxAftKAr4wNoMmG0gOLVcEUz2KDkVeg59Ye/LfzWziUJ4np6jLwgv+GqP
IrgRY0Fb5c2eU5dHKt1+wXauhqcOus1Y2jsAg6yqDtgies4p9/8KH+E8EtjWPXYT
SCil+QBkTVG7CD7qhh8BgdzojoxMrq6X00JLKD7tauwyx9YSOGW19eY1eYzp2sf+
gE01VfGqqEiosZoA6csOZFYbcsfjpQvloQJVbdUJ6jdptfHrQyuBOL67qVh0gvuo
vYFZ5YEKCZcAKD89+uenz6GkM2uVNDFGU2uLQeQq4daU5XGJqKp83Ac1V+4HmAZP
/D3/MLPAi3S0InsSgjvws3ZmXiQ6SqXg4gJ5aAd9OKubJxhDLk2saQgJ4O4T5HYE
DQXsIhNSGehce1q1APcTVLS2znzzAg7b1RO/P3KPOzlwLzVvEDi+k1fP4qUiS6ae
KhaqCEVvDVVo1yLLXOa0z/+edHAzhbbfmiRKA8wPddf4JCSoD+PJOTQdB+7sYMX9
ZTRpcigE/HYmCH1wGA34n29Q07Srv/AshjJWqz2PGfU1jZTFxKaewHKupN/kSW5i
Xw0EEdi9Ojzmhtv1rmpnAjgYJ3Odb6OqzwsU0OL/hzmcZNnQDVJHl9Xwu/JZkjUo
T11op5O0N4PQQhh9TyN2PCbdA+xnbiABlWwd42TzwdYazeko1+ZondnuGhNY4zyb
gtylRRWfgXLGWN0pbd7Dzelk4BeM3tNTQEQnUlOobQEKL45vQ/oLR/513jHm3fPk
Q6qcJV8ojOv7eue7ZIptW6TuKI5uB6L9NTB6hOUbJyR78Js/SXf6dWfux3fxkNjL
a0QEZfmTtQAgexNDY3wpiZ5Acl708BLBS+fMictJBjPUmKFXjOTya0pO/mClrL+n
VWiggApyfoMNTim5pm4l34CB46SZCwWuhL01X+J7/+rH3BqP1vgTpNFayzs9AGjx
hzt1AUrBGylYvRPxK7OiEb/OlfuT56D1i1960ME6rS68Kw6ev5R/D4yANpscOBKu
jWEwBpzmjwBKHXRLAdB62JHobW1Bh1g4E8IZ3ivY3ThufeeOlzgWIh1m7s/BUtN6
3/empPoIZVUT0c54916ttmv+oIji8qXMopTH9Zo2NPFEbJLpYTkSLG6sFxAOSYYG
4gtLCN/JLc+YpVcFpUiDNEkgBUxomniv33siBGtf7vdJ2QnDA/3gFq31F8hSbuFv
qbPY80nY8bnX1pN4Xmb2nEI/7kgz4ponNBg/HaEeSNs1byUVWRZ/wJLS9qFnid0C
8PPktA+R1MQgO7JzopDNLhOE7oqnzb8D6LqKKjPHEbZK5jnST+WzggzOZvgYpgkD
voZvM7W7Ntw1wCsGbxMroC/8qjkktEuOB4/obpSfE7VdJqyUuTL9no3SIIkOrFP4
TYpCRI2oIJETTUp80xGu8Wf0EawkI67Ro6pdDEqH7K+bb2Ukc56cwR3W2xIW/wtI
NMdTLJemKGidE2pTUkL5FDsYQu4NcaCh3VrcWYxhaGh++j221EdNThbCuGkQ0O7U
+VkbOhwot88IBGlk9CoFz/0JkCXHQ4C+e32EdXtAiArgqabAcCB9pKym8l08Hikf
uRhAf2dXkYRdzQmL9znASpcGimHYCsicA8D+V/55IQNpKbsBSKqqkFvOILNIwHIj
UTYn1XcnnifVvkZWTCHI6OpntA1eFaxkMkBIQ+hHRzzn9AwGOYUW35YUYM8vKJhP
txLDN3Bekbr+wpspTXBW7EIPzBWPVWbcl+6TOieUrNe+JQ1TQdBdMSDi/v1lsqPy
RM55Blf6l5EzuDAjkYF+LfDcvDHG8tSfjJwgW5QcE/UkFPAiqhByMW5tmyQR//D9
ARw+MEoH5qYFnCim9w2sJ0tdQ0XFGP3zO8xMNAERE71lN3Wv3z73luAREc34ymDh
6RRDrNJofE3i4y7S1pOUNR5vIOUK7lSLkXt7D5gorPrMX56LrKfB911qrBEsSTSj
dosLnaXh4ra9qoyGFoiRaC/jTbgKCNcSU0FCYGGQVy/vCaZKXVxilrlbxnaHij2q
kPCs7F1RaIOiFYUbk2ncOynZ2yT645a6TEojmZiuKXGDRZqHB05EWwFElzgnE1oC
qf5HEbCa2WepLL6XFrqCsqI/rYMJFmPqnFGi8819Ge7gt1lXRJBxsrHIBJBcx4Hc
6kv8rsQm+CyKxOMxXwTH+HIZOuqsTumZAVe5MgqPbM67UrQ+Gl2u8al2UXbVrSLk
gq9yFFWCRbIQdh+GB58sG5C5jUB5vyrowTjAgS+uZPhFJT1FzQdpdVDOZvYgLNnu
zLbgpYxgBxd0WxVN62Kr7Zy5mUL6x2Qs9b+zHPspsu+wZYu1OMMv4J2L3JLoL5wO
iZA/fmbHPEx40ATZPnICe+yyGX/cdhPH43M7b4Va9SGYqR2AIu5q061UsLGzVL3Y
xNfzJZf9q1jN3ADy4lzfN6JSJr4eoGlL7tZ/XkDrP/EV4VYzaNPHUqmtks09SS6l
YrTtEzpu65mpJBwTj9DJJ2VzoXbEPI5QiPKVnvMvyFoL7jhxuKjBI9Wx6weh6XcL
+UjhAGP+jH3PNF154LFfsy5RU/gYd99wqDbqeNWEA7ODpeaAcymeiivBsaCs+X1n
brH8EggdcE1XlI0vE7vghKIe8W5yMH6PWZPMqLydi7tvV4/YqWONRM9gOWnp+LpO
8yL1/SIO/mh9gcLAMFVSuAksiQAWjbqZCpSQ1JBWSTL7uqu0LalntGCJ1V5IeU41
njB//w1F41brvyNv1Bpcq27JLpYTkVnmpU+8Xdk9UQtuJeHo4HhYSuMwgtFdNDtv
rd3TibgJeZvBAbuHebOj9qEoKVMRZgrI1Ju6Yy1c3IjOlAJUawPytzLpcb8c5A4t
Sewucr0ecH9jah2aD1izO/w5LoEwyjySYxjMFYq05o0nA/P7yXlJVGEJSloNE8ag
3Wk3O1pxWckqt8MjQvKd/opf9qVj4Lyw2A+MxEqz3lqOUH9N7Ggz+qG3P6So50IJ
ErW9oMwPyhRNvAVvkXlY1ZnKC39GJqkaRQdJZgZFkVKxTTAuOtL21B+t/cvJ9zCA
rd9mbEl3ntPs3Q7rDZpbp6W5neKsEqcnIPMLaJiilllVz1tUxzSs7RkzDMj7zJao
Gn3rQglr4XCahD+LN+jvxiScWX62P5KkHyAdpi9F70j2gRkMZGWUn5nwKGtQtVTm
l3c2Ad6zd5GRYHl77we/lEHc0z8A/EliJHFmwfKQu9A3y2GzPNTsamvf2SrIoldA
XUuI2NkC/hdISb/uPqHjV+68l2JiXDF1rLrh5tIXrHLhuEC4BYvbD3AowLlGABzx
vNbFGlDyETbxvGG0GmdLFfQOIs7xxujy1VC76v8Fb1zdkMpegZLxyXYateyuvY9J
BE1p5ouhrx+wo5+rpwyeSDUv4i5rJXnulL33aTb1/TM/fL/xL4UCcriX+1pacjcA
V7x5PezJ6QG2qujlCVAJOgNh4XwuUglEjpg/2x/UJjH7wGlNy1X1vN26+wcThg8V
nepmyYXrxzAB2vFHbfyhsghewtDC+oTxFZzNS67z9Wa0Pqs9lg6pU4jQOFOHR0LQ
zj5bhUObwIB9fWRv8NIegIfomY6bu9IOYObyfigJGcfHUmnvh8fkm7LXOSXFOaP5
C8nCpGzVUfu1+yCbhffxurSP4V4+/oEU3lhCKLfbYJHczV2IjlRy2Kqvf65pmmb2
MhfviKqX6f9c8RtT9z8KRZFSJVLY2ZsTEYFiS5anJnyTv4SAD/Aiqi3LSKwDvWip
OR/iqzYk+bqvDFMlqwlTtYc0ych5BUY38Lede0zEW0brg8H9p0p6m9dExp3SCTNS
iH/VEVgWfxdWMmJlrIHxY9ijaisvNtSTtQhBZ2pfPEhXHicR+uvs0+2xtAtumzND
z0pzFbzbJaQxvNYCFEHyDLDzciRz1QGwqVa401LEz1ROCnxz/PmBslu3RMJqIizz
hJIW6tt72IDdAN9m+e5jyAdV8wWIqe/R1qQUpfRHekqrcbcpoG03toACNDjLMqJP
nWMomBEL+CfYm1DXnyQxYj79xFWoSmMiu8kvIp/p6XqvfIjw1d4CTPbE2RdDv3P4
nT43FrNPJJjiSt8+CENvGJsCj4M5E9e6vfncErgAE9whzZlFbo9ugVtLZPw4pQEK
P5V3KGYdQLe7GcuEa0pX+aJ6EsYSFe1hi2vi0Xa2egKeBOGIAQurztCuaUjM7EF5
wF9cVOUYEx52CawmnovezgRJDYqXF6dB42gSDNWGl+QwIe0HBUu8YSdSUAGInutq
SWH5QrkuWo91e60/Ex/llC4hF0OWHs7Ci5mkl3h5FrkPK1MsvaeHDvogwx0tar7z
6dCKFPbxL5kMmOvYBtM9XXo2UWk1onZIzUjIgcdzhI93cwhgpDRw0nGknDtBZyvo
wPc0eFPzv/qEDii3ESLksep4eYfE1udPoztocheFqvbnks+j3EKyP7LanYXMjqCG
uWbGrox63cFDopqD05oJ/hkutCTWPec3KLaUif/gnKMicvu1qWbaC12qCoz+k3A2
Iix7eiYg8suzcLvX1Q4pAIrj+82tnVvM2/dq+g2skDa4CYA3UjBUbuoY3yT2ei2n
U4KF34gnduazACWy2kaxVkAK7Kp03zFy9Gr7SSj6RPN3NCRcS/l9buFBuSPtpcY0
VR+6hEfecm8eifEpYmfh8fs3suy8a89MVQv4O5ligIb8HhHBeQbCk1GYM50uvhH9
sI5ai2S7pChnHaTJIQyiwlcjWe+iiwMreTsuRPxt0ZDeWDopVqiYgMWv1VHdK32a
8ytcL/01/G8sW6yQBKlkegwMFvCkiye4R4O5o19CslJwahQ33R3GNBEFf+P7B1RO
QRq3LJ0x+wJxS9keccrT/clhk03oaDllNddG+XXybb8aLAhIqyKOLhvu5I+3kKBB
LS9KkeIP0PFDVTHQjIXQ/rgSBBP8Nx15D6CAdeEXyHfy+PuD8O8joUFM7IQIboYX
6SvHkTQvxGGQsuEY0wZFDzqqOL3iqGc/yC+iQiUlpDO9vWGElhfmNj8nOipQSdGP
1XY+9PSyFtmVKTZc2N3PKv2GNw3q7ZjvE9tE0FU4AwQjDsrdi1brZ1FlH095wtQ9
BC2pKelzUAhHPi5wjxiZsyNzOTp9roDhHxZAckjjOs4jEj49A4Cg1720EcQ3lgQP
+AE4DgmptfH+/8eXzp6RC0K9fQznC8TpXs6A+zq3GgRt1lZZSjpAYaFmuea/YcOt
AIxgATA86EIc5gKP0kQ6Lu4B7aw/GU+taCG10PvL/mfTRgVYLloOGlZ6jD8egB7i
kN1SX03O9zTl84G+tjeGb5m/rnjend/2L3fgaBD3Tcaynybcqyf9Rbl6lc6Xcv5R
h0HWqNw9zx6CS9sYyyrHWoF5fJy0PgB6AbPe5nOoC4eFhRZJpcn1x8HVZbM8U83Z
WjL6zAxCGHzflf6YySCSDRvdynDrHJwXEen5uRFOUQTJNey8UhfFJSh4yT5+SGmy
I3qJD7B6G857VOvJFbHmLGk9F9YaGugCVO/saPUBnIHgNp7jJPgAXNVSDdZhHsH5
mTcC6BjP47Xx3Ez/klbLscYxfwE/nweW1mM6JBfVqSXjAl7gceuoeuoasFgBd1G5
kwl+28A6ARLzSMDkDTDU9Ah0BZs3pw7mk1DM1oaUym9UYwLkmHojHp+CQzQoDvQQ
BQH73aymEx8YOqpUSfEo61LQoN1oIRLWYZKhSaZ0juWu1Pxu+hJKgKcHBSFsYS4e
bKirotDRtaSyKXzQffigGG27yzlziFYAV8fN9RyBzcX987OEVsHOhLxH3o6CLumI
tDH0yQIhCFM0cWU/NMI45w1S/OHai65Mzp9dla39m4WT2S5HbAUHIi+gKVuKKal2
D2XFYYRqOljBFzFybUSOveUjOSaN4wP8P0YMx1w8kd9Q57cCM9FJTOOamlkjuc+D
I+xRpvh3ymKHlfMkUM+L4UEtAcCvI7b1gWdLwR4sd5PPCIIn+V+SlkUHunNh3PRf
ZNOf72Jjvcd93gjeXbF9ALu8EVDy/eXRLG8RoQusQw6w23V5Sx8yOUnHTRxEMMq4
I2tHXcBehhPs6LGdnyWzcg6btMHPWMsA+FhlmxGb0nmJ0X38PevbzAlV8I/mGoXA
+qX2vLSmxwVieXOT6Qo4SbGUwgwd7X4ehKYY67vt8b0ltN/vmca8II6ALu8RTIVS
5jqojMas9LFkDejtCcA/u3aBGx57k9jeKxWFg3l+F+5mmSmjhv5IMzEsGZFEMLz8
KobQBGrtmU3/yh5z+gqdNPkyBaiaZKUKtMiOiOarb+9xmOzNofH/TbdBTmfHZAJl
h4k/Bv/P5hh+ATMR22wvde0Fsrs6HwXfp79T1C7Y71hu6pA5Ze5QX9JbXiCoAjki
jstAwyfIXzfD79myzF8ACbPPUtkxeBhkrnGThNSDF0RoG+8Z8B20UakDcOOlGASY
YMbZo6fmx8MOwqMXSKpK9H39/itdC230d2TN4d5ClOHSHkyel6kdm6PDYQyNxi2I
sJMq8oAYdJES0kuYwY+tM23M9zDAktocb7iryNVLLNb7oYDRgumE1cg4h0DJO+oF
1/CkcTCZNNjr2OMcykfjFkj8hwFwJZzMxe3467bjRT8JQpFrm+9vdJW4LNe05zhA
mwJd72H/f1RpeM37vmYoJF3Am3pHeIAvK1/yROky+YLJQH2v4fAJU14xm59u5N53
o6O6LdAcA9t8EdhTCJbtF0mCMiFvaPwTCV+Ol4YwGl8nF2oAe5427DNw6pIuj4d3
kCzU7aq11W89jpYByqRwFasYnFqNczxd4UNYVTP0g4YZYt55akn6OiMIbSfv+8ME
6pF5UO9EgmmL6IP8JY5/8OtjiBnUQNcgPTfDb+cUOySXIVb4frVE2UhkC9B7p18z
PBq/rIWQifXLudWtbcVKufzgG0lJOTUFiSnK+Lf9yZUSSIkBYIlXs+bCV+Ofiy7y
8AorqdhCQ7jAiMBeEI6BMFtFunaxwQombp0FhJUzvGf/RvngybTYJlGkee+Ot8gd
1sCLjCEy0efyc5Cw6X6suVfCQo6oIDvk+VC02K4I2bICA51uKz/PwPxWVSjYJqps
pkBG5bBuFKLcKCKdYQ3ODxfy7VycFCK+M1FGmDHyotbw6BeYdEEJb+wyCkyQ5Kwy
YJyjUrczlb6FN7LZCnhy55xj9LQJHlj30NrrmO+aJiKSi8DLoXAO1dtbDh5+RMGJ
JfdklgGlxoflR2fZg3aVpDYwlGkwjbdXc0zNa6TYEC2ntIHYN+OEDw6gdWzQrmvy
QhRgfc3YGnIZ/Bp2XsoOjHsotQyh3ph9FDpXnR6ARs73z+Jb/e0h05kMPM8PiyhW
srIKHDlzMHne0zY+bqzVEwD24lRf5jdfjTfzFIw4fjFR7EKcMTaCkY7d/7seuKev
h1DLhVkkMgHJTAwueU8wVuZQO9r911JCg/joUlnRJc3Hiak4NIAZR0PeXv4MsICI
eKaLgR7td4qjyyVLTiOgfeCOvWUvRHLh3cmTC2fBbO3TB3Cz/bpsoQuSEJSm+TOb
L/69aCh6eIbUOx0T9kIjV8sRV7dySQkp35UF1IZHdPTs4B6f0rMW3kM7ZQVTqSwY
XgpzMoJpa+ncn8lVKHqL8Mfqx+cJMC18K+4EWUY9XXETofpiv5nhZxd8eVLrFyYP
1rb4zGCS9inUalcoMywZ9Kp5QCGOMZrD3DW3Uy26q4cVZHZ3F7VkuAonv3kjGQE/
LKg/oOJRL2oOeHU0VWsjMzvSnZVOOTQOHrXMmJUjNdynuKYy8G7cOBpnPeJor6n8
txMvSbk+IsANBsBCn2hrcGSb+/32GbRnj98OReqDdDBQPIzxQgIdpKZP+fzLIqBN
jekODb7msRmKINYQ4w6d3mNA1QaPQAJqdzZ9cYfVaLJgkvzX9jZ9dYvZzFms30SI
y6pz/UCzBdIczSBWMUN7OFoDJGyINWmFN/7vXLDjYH9Z1/CI4l+7QJR/o136hJBl
lXCeB2a9X0QTcHXEFu+33pjvj1OH3LMwz727JRpc88tmLEcmBuWGJIN2Cjnb0d5e
dyaGHkkQAksrQrh5dUYoT/frGrj8aGJAXzr50rN1kWT8e96hg2EE4pQDs7gFP3/T
SKGhvSQiqum6GpFljmeH8tYCuBk8LbV0v1KkLOHqqOWXYbnuFWNQh4/9T+uCI5Xp
xXBDbnCYb9xgEUXKnPRlcGYyd/fp+nOgSkUTeDn6ptxXp3vMq0tlgQkY0P7+qCar
F7PP6hPqqq+lleuea29GVJKsaQTpJJ5n3YvK0tuUG6cCRc1mDSR2llpUbFZNgl6P
JO1PKvb5teU2B9ullY1SUXRxf7bo8hLV7t4XbwfmMjTQ8HTtrgnMxVTApGI/6OBo
nwGhnP6yUzGKorYR8dG05IJmKpHIYXbpgD2QiSxfXFhQjzgvnGw5BV5dzeMUJ455
1lr0J5DLbvh/XbiMP5VfGqK9a6RH4fvjrKqFVxlTpibScMCt5cmzH5LiIYCtNTZ8
hwUAvVMm+dn2LLWuP+sGuS9MFLEHYfyIdIwyMy14yxXPCFBwmFFVnc30jUuvk3/U
raB1SDMEE4W+KqSmT3fUBJ2Dgsmc8XtVobujIFaH7tgBwy1gcZoYzwtU9w4BWWFq
RyThV7Zc9+9sPPHzpjqbCKELsgzw6TyC27dqM8i5GQQpSYQ3iHsv8Vjz3IRmvd6t
rjU23MAe9e90yfOT74qHQGLcPYTUwGVIoYJ3LycZd6KHNTJLi+97FJ//Hr05W6kp
WQZyADx8qTY0iMWO7NDDRe/o8Co8hIVeYVuTsnRAmOs/ndWw5syJLDbws3BLtM5p
qkWYZ6kDFijAXTr77T9IzPQmVCXLJxuotgMd5HGI3yJct2EtyCAVaAubNfToRjfJ
Z4nDkNOfImOUZpr6/YEsMKIEDdfw4PhcvNLuGhj79nKbhd/5ib/MuUpwkN59Q734
1cG+12z221lmNCFMCGoWHdBf7EE5+UuZgvVHgLp8Df7MEVvs90FT1qtAQVEhCC8r
lCSyUxzW3QYkUBoIq91Bt46CKrNoVAjG541hEGoYIzkUjF/4eTxTkmT2EeTwB1Vm
L9zXyAZXB/vsQyDrnOqfmvnM63PVrz192qHaTI2cxLr1H60bQ+HRalkG4ku34XR0
Tm2HrQB3OghH54sdjU7aKgQkmZX5iD9FGDtaFTM6jiQXxdfordCX+aS8yISflGr8
Pz0skGh1PhcYd61eh0Uk0niu7SZFk0rJcRcjxyJbL7GNeCHUP6WCMpV1OleA2TAr
MgOs6dyyRA1zRRFb7nizF/szrugAC+Ljo071vkb6bleG+OU53TSE9oABhCMR0kSf
jyyK0CBKl/vEXPvaqyBSoiw18Sw3t5e1CyOzPrtcIU5kiCPzd8x/b8wR/jjDbPVY
RbFNhQHo1bV6tx2qKosaK6+ooxQ9MK9fk0vvpXG3Jsm9tJJbeCwDNAqJtQj6zzPR
4SYsX1sChEGlTlZGgqBHDxAItwKdzwqp11fUsFNWY5A2nhSIqNh9gmN9qkBmMk3I
Fs2hVpT6cj5roVgavCCB0OTHRXZv6T5vBm2udNfsKbkYvE+yBzWYS+iK6Kfn0+qR
IyOeX1NGIvasewIjq8O2w+0CcHxsNR9lPsbEk/omRWBq8+ahjZ348BSCDnIh/I+J
0C9BlXoDs5WFJUyYDDz4bSTB0mzUxuQ67ZTtYwlbPxLwYEj8VG5IxsF0zJ9SJe/I
iSySFPw+RC2lZiHsXpqKYb8fVr8c0pjh7yAwyOj7kuASSQr5MF6T3IHY1XkYCVbX
TzrUPCpApIpeZxN1OI7wauZNPWjyObVoZ3C7leseMsEy0VbsBfuBLQgo5F06qE2g
ALDXz4D254xB1bsdbzSNNUre2O2dF5FisStPHR7SBI+OFOEBCI4zozaDFupDAOLj
3D6gPSGeYz4WGBDhi3ke8g/ppImcO7V7PZ49viyxn/wGDK+JS3XfEEUo8UMKNz/h
3cpboI1QK++b4D5C1EU2zkVYK4/umul6T4zjKzed3mOYBGl9YvpnNPJeYxZlmwln
swWRpdBD1BeZcTjqfT6JoSO40XiRVSkmzVeQjcOnwH0ysipFr+dzTy3LHEvgEsq4
kohY0n322MPhHycpYVwh4IJWN4uwYRVVDEbTNvUJBZtNaNVsmrgCK1MlBHXvsvAR
vGHIqEVSZOhj/fEB6MgXlMIUihEp4Pjxg8LFEEcyeMvjS4+Rmi8AIJLrYkM/+yb5
dgkBpx7ocFWIDqM1o0rKWR5gZZQ7cDG2uCffgUkr7/4+ZjTtrza1DB9qDvpHi/VB
NX/lLutyI3TGA/kojfHsTWBV048o+6pZFbMVv3A+x8u7r2Icmw2QQ8ec5g/NNPsS
BW0ZsNyQwP6IA8SNzFohDeIakdRPZZkxcnaJe6Hi8L4FqCyOZt61RaN93eh01dT2
d7t/qWi/+K4eFjXGvUKF9uxA1qXdfRHMYvwJwznYDycIC2Uf2qMei+WeD0bXZ18G
4nEyxLDNt9FwfNdjsTmkzbGWQLrfdMa470LvxaMUkrpHDpNm0mhQ8kmHblauXNna
z18uFEuUF5Hrx+IOCXcyHONi8z3lT2+2sBPTo1DKn7VuiZMhK7C5RlzvTJ9TgDMB
gTfiXj49Sbg2DXRrnKbw4z1LQnnYh2UqBmd3rCpUDiEJ07asMSJkkXDjEvq12lfR
RXNDth2NJsPpovXjOVSXZU971dYqWhrb7DeY2I6iFi4NoMuFwV3Zcc1Bspli1WaP
8nmYoGcqqlapoI9wJA3RwZ9bpQZR/Z8X0l+lrlHzV9Hemm0gRMnaHYxHVnXLkCyv
Cf36M3iv4TvKRGaKd3CyxyfwBGc9A2VrBtWN2LN7PVh6tkroaht+0HYx0VybRJUr
qAIdMDuUOqYo5jfzu9xdm7IwivXKzVVdny47XPjb0seIBMNiYdbC9jIyADnoq3Mt
f9eia5rOcYqj66LUu3CvJl4ixXhfOvt1bNeeZQmo6m6kCoFJh8vD8LveCXl9KRY1
C+aLO2tD6LGbF+N75i6H8qne9lhS0pcYgWv/ynJ+EzP+VspmobfKtCMQm7EfOU1o
rnVVPiYRorqkyAnUZbtvGAEHSpPdQc2yCDg/o/B1KaUsxHgG2v6hap7TQKvxo7aY
XL3BvJ0WCtHig8BRZDtgiGthKPovPsv3p0NqqI8GlkIdF/IKc8vNmQtyeQYUnF7G
qc4/epKyFAOjnV80D8sJ56HjRHexjPvpQjmnYdA/uCnQ5ZGkXyZ3nvcZQvDb8Tmh
EvcNRUVCc7dchpYDtq5tn3WjCuP/D2a9Ur3C/uF1iagFLgyQieiQSz1gQ38DC61P
veCPODSxeh35ItDRZZpts5fq9/m07TnngaGDLMTv1gkcFertgqsIQiL45dSNsvw4
pNNMqgnUI9/gvDRc5gGv2W2+W9mKPqcDmS0M0IZMb/8/E78afl7IxWh4WLWAzvOI
lByYTeXQnvH7uqrBufnSqLHEnzh2SHsuoPRXIVne6o4fW0SYox2NaV20VWuSJ1xm
gqBbMyakvR/VbLlLFT0rTKtfGOOH0hdjSHUUuxOUDwYUa+C85rW0D+zkK/wn8ySn
ly01eYjpXY1efAoxjGoYPubqBIekeB1V7G75lJJO6ZQsAn7g89BjjHRU635dCLey
0059v/Llly2qeWRF3s23bgdoE+YBp7n+s+wuZ0xRhT8uX5b6WEvK52O2Pqrfn3nI
RR1f6CnQmrAkGu5cbtzAWQSkeMFwpArkHEptKSw27hc7m+LmCkjJ3+KfAcJXrmda
9ED2qFHkc103cBnxuFqA7+8Mc4/JLmqJAt/f8yAoEJzcUqXOGhHVxCwJFN0npjG1
9AjMtP/a5JvVFPEjL/Cg7TvKu9UP0hsjsQQY3gcow7Q4JpgJ1JThp7aTBsOtOMUp
scQAsAiZ0sYM+8fWTS64L+RRqEt2CNhUQyEfMWAfwugE/vbye3q3h5xhGESzdy+j
Wnx457LBLhyYqyCadxfC4mPfxS70wwp9Nm9Q+rya9wf51cV4q6WRsK8nkoMNeYR0
ePzx2ic0mErKc3ibW0nyja+6mWhJE3YezeEbxymBf40aGxhpRbWFrTJOmz6oberr
262z7gEXDMrkmBqDeF4boNomoU0rBAooXKaozflpOklf7czO+YGUg9YKIXBTMxAQ
nXz4xBRSHPPgeCh4aED4VwU4SqskRaWSab45BRC/g3PTvSi2lUbqFUdtl+BOM3ZX
+HFdMzbfkD23wLN60m3vBDBXXoxcFC/x8yLHhDQr5EvbAQzWUki995eP7pfrG84q
AkD16u+jDkHqYHpffxKFcPBmSH/m+/wBO2yrxmSi54m0IKXdRO7Fbla+DIHCHpDF
pJUAnFLnhx7KV7jHeFAvYvVA6ulHb+s/R84t7OpnGLdvbSWelDpLVQHNsf5K8qJ7
CBREPL4ti5Py34pLM/CUJqDQ7/fIzbjLWmbsjtHPtKKEGZiU8cwrKovv/8a6mJsT
tYIFc8PQb0rny41AQw+t2WweHllTjsoQZTPibZv+/t+QmH/ubqzaR6zxOsvMMVXt
BjDbk0GCW9iCx8b8RLQiFo8YpexjK4rADUJudMG6nkMxYNZJMLWNvqboZK+U77Kb
EV4pKr8LPZ067u75KlfAE1xtJUjBeqw6chrnphpu77/YEtuZiE3aA6P5SjRZ0VzD
KRWyWmbwmqakMnoZoCEKLMwsP2cb+kDc7GQZ3PMCwVSdYBTezajRHoLBDcsQ66ZM
3i/R08zG/eB9naUfb6opNLj/cu4jO1vzG+xyjM/jwqhVh58/eHV6QdjG5BMfUEKn
ETmjZwR/8IKgClCBbLYk3pf/qybhNHuUkuc/TVjxQDv6VC18Jj7H57JoofGcugUO
zsJzF+ao/4ZYh8ZQK9SCl9d4mSTLDtFAIlnijcXCsoRBZvXmmhpHFtEnM6iQbD4J
u1lhU0jQAj5jtheQm2Ll56XEF570F4uY9urRK8IcsHJJTA4DEUGdAI1o5ZP0VIZO
gy4NyZNz/Is6SPRh0QeQUcAPzVI2onXpF7vHl92r7cTgANaP1kOxUyDxTR7fEawp
ODmxAWH3M7SOWQjz8umcTSZwpq//IYRNiEQaeH0Shtcf/Zf8E//uuFD5LJ56kUbc
QArx+YuEdETS4OHdsDRf8qm4ACcQ1HLMu0PXNseVxqTphnZ33mLDCE7caJhhW5Lc
3B3adWpY1E+qPYkRxCxZ4BBx5HOj+gN/tu2q6oKIzoqNVjaK8grK2se2q/lXvuQJ
3PpaG35ouEvhJJEJyesiEiPE+FIO8p3zlPOfELZwkfgHl6b5nqD0Qc+m7IpsQmx7
/qo/KTpzeM3IkaROesLL4LgkG7Q7Jb4bgsKgWjU4hEheWFhBPJclpRRyZbx+CmGB
+OD8evm6UqsN38CXM7FLvMUbAumzRYDiFqsaHokchGMu86fdJjUnqLJZzkhukfws
dFLoBex0YvWRDUpU5YJocK5lztjClf1akNxrUhr09sdHpz4zkDGQ1awN9LvwOiGz
+sQ9nD7Xm8rQeZFy6M3pYlTekVody1GSXbjICjFKrns9z3hD3D8rkBHyDRaXrgKL
uwW60SzlJNyuEBfIpiulIlKY5GUCHlsYSFEffcL16k56vm3sRnYQCq0NGwQB/eom
bB9ofjrRg/Lw+L7ZW1U050vPko9+NNV8gc2upHwRzVI2I101Vyoo3GfIVhtbCFPk
0HRj0I37OqAwMGtk7L1+SNlrxNkUQRivKkoVRJ0aUdfRe+B5aniYhmT/M9OF1H3r
pA6PfUccXEs4JKdWmwX2XBMkdUJrEjctPsXyPMeQLUAHjIBnDaHPBPJCwnodR7g2
0IHRf+iVSDMBCep2t7J8c0zuxvuwltau6mEPGUQScL1i/21qnjHnAhgdcjVB9SyX
/JvawmxieEenicxZfd1c/X35pjc8+kZKmuDb2zpDBAC4D0/hnfEjyuvp6yQ6WAva
7nmLEJWUd4VZo1X3iFuBGGZnc2xbGFoCG7XaA+/nhYju4KRkYi/UkGEo0SsWTJgK
i6yCl7055u+2mQ17Ag7UuA7o7U9OgjzTvEpbm9xDG9J3O9MRjEJ3B3R3TgnRYOg7
cYH1Aj542+g0mNRxOVlbSCBe4mrAZlRI1Hwf916VDuaTP9aR1zTHbtkyN0xD1+h5
fABGhd7JhPzwnFtXtYCMpyA4APQyqWT/3zYknkxCJeeudjbT1CbywGxQeYXiETFD
HuJyaY7DW5QrCFSAn0xrU2B0ElVbaI9ojRZaRGieYgYiG4Dd9QzFJB2mtlO/4SuS
TJmy4wYQcMhy0DzorIoCQesHbdFXtjydBEgFxTLKQhLksmBfMkAlve0e54k0A+W9
Yud6DhUKIIUI2EhJuex4rdsjNi0zGt+uwu4zRe7nJHjr8JpIyGOxd6PndAnQgPJe
hfQZHkFeh5i2d5VpwiLBRSEp+Izc7ZKwJL4W+k63I6oPPxqjmVNOwQylGVsR91xq
P4UyQ0x3ZyT1m65mS9FTYwoc6JVvm8w8z5qaMiKSX8zV6BD5+wiasJlteNasUQJz
kAVfXyYPgeRTShsLUBs7Phxnbnwbw1Rwlt7OKkGMqVO5c58yz78bh8ZPGN0iIEV4
0pm1+J+7YP194C+0ksWKzeIVablg5OrqVf5lSrW+ApcBKa1rPitVpnSJ01dcUdpL
q/V1HsYYmLY/M1NGJwEZrhhdp8msdYJnE0PqmSrM2dqOde52aiG/0uLIDoM47+6A
bxHREv/SBf9mHpSWffcN0xDMp7XhXgeGsl5MCq+JNNUqtOSuswMxJDa4li//AFxq
WfygxEa1idrOeP2M18tt5kTPOpkayhxyEZMxzT1q4UeBkhKYu9Q7dPIou4m3Y/qH
qzuR2S+gDfXjfNr+HeXPw5DRRLEOWyR+lUT40tn/ws3pg8u91xlKVu4gJJk4zxrB
VIkzezxJ8dnOkOpzURLpLYdX87FMcxfZqVEtJeWFAC+w6WbxUK/suAagrUq+MvNJ
K4OZFLD5K2yNnXsucM4j9Pw4x5MXhsiVf+9CWw6XumbV7h14FIeHrYT09goX9R5O
Q0o6tFmfVJakX2V2qMWV4TVrlitu8Uu5drwXBeHPsA5xCgqrM2TJzrLI1nV0YNnx
jNBD6IKXxTGtJ7xFRmKQBz7kriTJau8KZay/lF3MXkdvz0ldq2KgZ7wtBga9o31E
OcVjxPqFueqfRdzR4+A3rIXJFoqm58sdzLhi4fzV405OsA1ToRTbkygKzWBTefbR
DFnnajOUBd2mbncNOjbP7cjstI+U2sCs8+IVCvItYvANQjlFdTsacqTY3jx/dVrC
j8D2HGmqFXm0ozDOYyFfnXfLWYzJN/ukvegN19b89+iJZYbYfuiV8rL2edT9AAbb
vYrl1PO7W0+hnLKg+omgMe9I3st4GCdQ2Q34Mk8RgEo/Cht/R61L4gSRPowhtHVE
cmdxtoE118R4e9ferEh9PshR+KAjSMWwgTQUpTNXu8FQ5KAinHe4SVskAKYlmWIw
KhEVMaCvXGBD5AMGmDNaPgK1GdvOpIZp8otvfB4jPntHYi6UlhCsVZD59aivyos8
ySgXLtM/7Fza66ZEI5cSJX7Khdc00I5wpOfTmj9YF0Q7ICEj93S1wyFEigluzlLf
MVYN+4OIrQz5JcHTVB+WNcFp530QKx/h8Iz+l1guHTsFJC9Hw2JSiP65W+lveOoO
Io7OzyjNWUGAb+KPvVPhw2VStoRKTw39gHEusMRij7WfC5zv2vFHJRsF4DMlKRTd
IvFJyW3zV9ME4bTzvfiZCW8Cq6q9IoDsvPKr7p4BrNdN79pcK6H8Nng6yZjWZk7X
yhlo/BmFKrI0kwAAPUo7mgy4FUc0kBH4I/Qt1Dl5KjxjszYLyG+KBjBnVZ44Q55z
wIdnFdP1wcLOMDrpi/00Nc+n1+1miVLGMCWuAxNr+QzUx6PaaoGj7pat9KBdHFwR
up9bj+llF3mJIOXg+IJsIkweXQ4UM9wtIS+SaJ+RnO7Hk2+MU5pQuO0czol6nzPA
Ht425OQS2LYL0c/Id1jTlwKj+U+I+ikLjzL36FZVcAThnVjDU8uRm0n8I8cfcqaH
eFR2p5G343802DhBYjBWj7jhCg7FwsNt/7ikezyN0bXlVomhCZe8mva1OVNap3rv
KTXiMPxgN37uVdUZAu8fLUD533YxLucyifDnVEN5WeEaGHJxa6viFu/acolfly91
E/b0gJ3BsAtoGaN1Y8AR7sfXevmtzk6K59zYYpvx9jN0gS2FX2fNN8XjhlRUYx0B
lzlADVeIa6x4OgnrEzyRul0jBvohws6L8SsNqBPnTzN7znR9ENHMnYQkuVmDwlkx
weAO7t2ByS5jyOIZmRsgLZ/ieZ60OGxC9ZypbDPHyomzyL4zhjBmkzVE/mNxjB9y
NAMJd/Va3nBHW6ypff5cif6sc3449BnLKGFLKTn/cvRDmOMUHia1RCxJApMk9zX8
XcnzFFKu1TTNNjUml9gP3rZhGWBGg3uQbBk2P85KV6dV7SQdYGLvbDHXg7wRD6ke
qgXEIfjaXuRG4zWeYv/HzLWEoZq9uXH1V1b8XkYXzayCzCdaUgcAfwIST+kx9qP8
DUchiv7TSsWsWy20MlbD7j9KD/aGo9RhX7t25wJDr09D3EttepZh2c6f2ltlwTNQ
5RziDzi7wjaTyU9zUXsSWJijIEFZRWSv+FsDZD6LoUiGaOTXvn1QLQ8ADC33oTwf
JRziXIkDhY/NitcohQ915+Y1otdAUzwh0zDPU/SovORgQR4G7qO1iA9AR/5aNph+
kCCWC1JxKJh/xgAZvCEcbhmg9MvKmFO2l59kIhQQBRmpcLL7Smc/yW/4YTvJ1cKB
uI5lhakDfrNADxKr60vnVT9YDgcL3s7v3zsA52Y9KKtowbf9RaZ0ygcxcupFc3PD
SYWpW3h8ogvBcsRF/RoIdEBufJLcBOknB16Wjj/9eDQtDUwUIZodKXySq3Y99V5n
laf1uK0oD5hBqkuy8SxRhw3diDBabAtnIxS3RxSism9iF05W03ks6xp+nhjgzJlU
/zmdVidp31Muv+Tw8ydy3OHDrOtv50yRW2d9GEfhEMc3H19FP52dYt7bkJexUiYa
EiSA755KU/fVttQEja/hxcplD7FjvH0q6WTU5shpRGbQHniQ6iCaSaen4sI+/hyQ
7GPDjNWbuZzhFnelEXq2XsjIXTMUmef3Vcfya23KdZeo4Gp2cbb5ESKXpP0Jp9mm
SYjLatHNPvXGS9y8IcLrG/bm1gzl6NE67imFZAEundm/9T/WyCvMDrnczPPAzIEp
eSWQVA4NALARgoJv58FYXYEBwSKJPWJP9nJ9ecnC8XRKxbPm5/NBoeY1nUTqToMF
a4g4UAdPtmFwgxeHqfJFv3h7B7DkaaylDArm0pDJ9gn9wXjtkmmR450Afem/jA5B
TGcn/Ms8w5A8umYZ3O4geQm09SRxRU87bri5SAjZJXa9fAiKlFohifIwbZZJkJ1J
spu/+wSuIDsu8R7p4TfHYZ9TrUXOQWW6v0j+Pw2Pgv/sFHG1/7ZZ2VFUnEPGC0Qg
fRcRZPTM1Wohbb5VVVYK/Qt5FtCWdsT6hnaVlmYNaPcAcyQrh46BZIKHaUvWWpHR
12sOICBz4GCJoeU0Z9bjv+2dtO/82J2aONv7YGS3J4x51egAUHR8e7edF8PZ3jAh
2SGa5VXBFPJWlKTlWMp09iT32NLuUf7Gt5eapnsGgUV/2Nyej53nxEIPYOZN52mo
4HMC2ZCfc9Qp25q/GhOsY2Q3lGflq/sY1uO7KelkhrnJtmRSiKh6XkdOLBMynxBv
9wOLAyJc7t6jBujDNVIxskV/PYMcX0Zxg07exq/gzWxJbCigjGtYUKOTWChiGfZP
vxLVPuAbcDoi8bD1rL53Wxqg7I9ESCo2HH26LpuOYFJRlodNRTHNr4dmKmMGvJZz
rK4etE81Rcp6+f2sE5gBgkLicfezSE4TTxkyOgXYdxAKS50X3g/j9YyhOEw61zLY
XwzBoRpcPmbc5/xRrIwN3yUV28DN/U3+WglKYVSaDcWvYveXwCqBuT18CCA7fDXC
OlO6LHZspsZKtxpBCfSnNdOVD1bOvLaQdo2CgcvMklyblpWj+Mi5R0LELKL8rZky
EFuXiOaAs7RUAmlk066HZMQ0ndJO0JEWeIV4N6yPpnxBer6MZfU3jaVB2DNUkqJc
39OftZqLcPGhO6rUHVBs4H5AZb9i4mS449l8X5ZYrYVIE9mowCelU8A04eRoecjQ
Mn0M6Q389akLoe1FXiOXXZDz0C8Azg+4TFtnNzsXA2JDt2w2p+dBzmzzixTSyOcz
PuVh8dXIrPALBNRk0Blj4DO4Nkzc4kpQCgYQctgPwsF6IHRVRqztIIg87mVuLmKm
sJMCevxGaz3sRoLWBDwH7oOGley621dD4zVLSIYc0PnF5qrO3tCqkIjr1PVWJ4Zs
iTp3RCEGqlsOX126e7StoOaaDzDFvpQL23Se6j3oQPAgB6H0W9F4KNUMHLjmRCJG
LB9EzD6p6nz+1ylUpAWJrUeebqR0kzuUKmjbqpycTP+F1mSusIBV34q7pGSiFv3R
g4uEHC81z3Sd27vqL1R9GzOB8Ia6cfl5WUhdyeuyTGw6R28eIcyOwgkYYNBKgy4J
6s9pfN3u12dkBWwOzlPwnffg9f+9PFpUz8Yb7RUBLbZeMQZW6lWxNERuCEDyvU0i
xL9ICjrK6DlE+kM+GHqireKTFMZZaWl3/XHvzWUvt3/NVGcdTYTzEIexPzN7ylm6
v2ejQVTjlgUDgZlQ0px8K7BIa0bO89VHN7meRShlFs2biwMfNzXOm8iW3eWftBOs
qoU8OnTrFsh5HJ9hMt/CtjLxtl3vUWsD26n8F4rzolgBKaoPB7nlTyus9B5DvIzR
1FWyFuuUokq4dnvHcDOCL3VGfvxetWiyp7mZ+Gv9EmLhtxByMm3DleaPWEATjV3G
6qg/XG9JzNAArb7Qreqdx1qLzIr/sBKirbhSv1iV8g/+F2Lh2V4AtYrh7d/az/b5
FsNi34ox+4+HOlXbn5k4+GUKWYWhVaQ4kv9XrzxurQJOL+KVzCbfES+rEMj1V0fC
B7lzJ4GOET06UPfEDkiMPNJHuUGwWzF1HlioenqGEzhPJv5eHT5kENUqHl7vpdEj
poZQeVzTjxtgwSLFu3vW2LKGch90CgglV3KrLP0hvzI7Y87FJPuoWu0qDNF9yhzz
/jm1qjriy0vkMrZYsQoF9UdqILywoTG4aOXXaPFE8tp/dy9R9tyO7hx3ogefL4zh
jJdJxdfYeyA5oAzEkdwFY7o5KM+U47yALIZYdVd4izokS9++LBBZ4YBGd8f9zVmN
zHrTvZIfFcudPukdx0qNDQyZn0bf/h8rHHjeyilK3nGyy32ZXciyIcgUb5oM2gS2
vjakItmDLH/Z6+rfadvsZcwabj8h1xRiEuCgrW9DYgEnqtIwjMISBCjrVeaQwB2S
XwNnj0z7U3xjQXNT99LmjOp3/PJmfgQRagy4v8QsCetiYAGXVy09inWs56rAcx2B
9U7INtZI56mu05oJoVwdEJjQQGkud+2R2mNA0CbcGK0hq3XUj+XZunzyZNexzkc7
s9GSq8yu2zEZroNKRe3IzySB1RUgMtqVb1V9NXglMWgE55Qemqs6T+EuGT4RuGgF
h08l/QespWqJltgqKNYCS6Lxd9DP7fOxAETgDZuv/QVHklsXSMXwWVgKZCRx/di8
70JQUQCYCkDbz6WL9QTagyDmJJX+QH1jyMIMmEcuZDRdLmzUPBzEYhYnN+RVAl2T
q+z+IJgqhnWbh9RAjpCtK4bPEMKQsTTZBv5YTlyzVcRfw5vqGwx2Bid6R4QHU9uZ
hx0ISHQbkful+SB8L3lUVBvJgluFZb7wOrdK4mOjeal5To6l5byjAjXi9tc0+Xaa
iF5tLApa7lHgGY6/yJsHga9uAXR9faiu9o/ykRAfXaleUisfeF1w3wgE2CungZsn
O/u1dlbC+LedCpXsElw9F09M7V34Fd5jpqr1t1zTU7af3QLpVJLWqSNNo2BIy7NZ
O/r8lUOo/66+EZq+6DZVQK9M9OtAXiFbnMWwFRgbvx4Fgn2nRMwYP6n2EkbjIzzs
nQG7CLIG95tlPFgC1FLfaILN9W981WcZpb4foE7ky73NMLehGiGACP4ozdM53qXx
f07Zy5O2dFBhNxAS3WN02p2zKlth0vh7jqm7Ut+FcOJhtEVQXNmzKlOPp0u3VMw0
wCZoCDNAza/0NhP8wsRL4pVVBR/bh7b3V8BVeo537UQbveZ6dOqxr4vEgReHXNqg
jXo+7S3/UsDOZbh/ER9ZyUqNC52JBTl47jH5uFWwaUTfhmKyjKfhsqY8lPBJVg3z
EaM0dyRD39tHzz7bCiO5QdrmOBMH0k1m9TQk9ZYMp6N1+PGn8v3kNwqeXLeWYXj1
KbSaj+ZJk+oMdJ1SfLLvWjs/IkKSmXfcnxnbeyJZGE7zXut4EdMlTyrIbWuSo+qu
0PbsMNQ7lg0SGOhVkZCLsA0ZVXcyIkvIOegA7YrSwKOYvaM8HRezvSBnZwM/8Rjz
4kzNuKvKOSAXaSZ5nWDnNclo0+4MyM39nA+CE0WLnuME4mqpv9eAmLYuy1KUpi0p
Ruc5/nIvYfAB+ZmdY02kb8dW+/Wb1bUKhfHOLkoU+Eu+PcTWqPiDMxKj+QFDpc/k
y0uKwlXP202HT0BRt+hMyVnLO1EQWktj6jdGG83HG38HRlDQs1O73vepneLjntQZ
dVbaTJ3PjXbveVown6AesXB7M3oJ0HfoL5+WqVL/fJrVq487bL80m/Wy9DTC0Y5o
tyuD3OHNjhfLVVn3wKUlbUYIdrY4B2M0nOTwbaMSWVGuO4bM8wLqgkzPRaFumckm
K8spEHLAVC6M1oQOSyr0ZTvjXGRp+gn1AGxYlLB7TIeQo/WkES85z9wXV5YOCxZ+
bEw0rte4Qv1eOG5bjjV5rKORSUVlkrCECrIRc2KQLYjefPP6gimTHGNu45ZUZual
CNU+MCeM7aSvfNzgZ9xugFyHSWhpKLuLHz6UQGdKaQ2W4DLmECsHEShsH+aIVe6a
Fdc9lRqWl40jWuqZmpilNJhAfPyYmQ2weoJCXhqwBzxOn9IGMZq4G9ve1TiPe6y2
489Jlz8bioWH1EZzF+Ypk6dESVy9voDI2n06Jtoa/CtN7MsbeSKwRJY72rIEmA/g
I9UI5TPyxdIvnBlg40+H9zxO4j0+Z0DEyQeGWSYe+s+Ko4TGynbd3QgZtXsUSIAL
Oe9NE3KPtYVsy33p7zJX4nfR9+tzjLSdCwdiMcYuyXQaWYKi6H3PPG8rSytBnJox
cLQkZt6wsgcVqFC5VsTe0Jl+6cYzzQdpD6a0XN95XGabSN6F2Bph7RQLEmccR/nA
wYF41O+zLqFyGxbSsV+NhijKa4WCRQiU/yoqbh76/ypz7gMTW1/LgQIVDrvOcAzQ
p0nNO86EZhF0r0DtdrEQ+TWNkzOW3UQLjZNv9JTEDGrLqFULXPt2cPkoJg4V8/x+
FzgttWJgTpCrR6Yvd75nfuPGj/59sBV57BiqZ1aqUajR1fErOs+LfDEn5uH2x7JM
ZVhSh8wm2ktXHHtP2xqS2gmfNvWo5w9Xk+CmQEg3VOiDm1R/m0oB6SiyO8Sv53Iv
eukxmb3qllRADgiTBYVLnfEHxK9khvq+Qq/gfcx9spf0l702S3q1nISBBTtVx42O
Ajv8SkWxwmY2ZsAdmjMpsPrKX1lVNs/vSvzs67drAwEqCduKKJ5DBBcUB4Dr/QWP
mKanWnJ22aAs/dqknb9/i/HMm9QMaLKCun+dD945jHMzG3n7i7q7o1v9pGIuAWsd
pNNtYDZuUzSDRSGzmalPK36URPNkkVjBpMRW+xlg1kAWqeMtq80mH/1dFCIsUqSo
fyfE1pTtAza1cnxoqsvvAUVUgZVGile/kXt8ojDmywkOysQ8rZ9YmEilP9GGDXBq
sy+4AmpcW6ytzDKrF3CzjKlgk36GsHtrF4Dxd28aIKvOlGiUkzvE4TRq3cRjfDGy
GFhGGMSbjzOfM09EaWhUsjtaPBNMTssO1DleEqNlkEBe3LcnwPK46ZNysEa6pVjG
KHXgyeLxMjYcOCAjjX3lx6U8xPj0kr19TuYyhg3gH6ImTUClhPSOt2ZcPjFkV8wP
SA9gbF3D5J4ozWMqf66kvh9k8PW4MZwaBevjk4wEC38fkzKmxulihqrceZi0xS4W
93Z410GJoUg4bMcrty9jQd7sUj/jIaY7wTtjFYoGjEdAT9oGwGxZhosStI/Moe2M
q83wwD8UvYeSZtI9ksWCUjR1DmO6WHobA2xIg0/Is0eyg0aXlgm1RsnfU4g5Uz3M
TWryDAjUtXmmffQ2t1VHrZdokZBp2nNkGTB5xL38GHGyV0JSBzWIm+Yym/xjtgjo
zjxfOl33qIaRThmvHFk9Q2l4ooz+Kv+pYoyjxP5z21AD2uj8CspFzfSagbG6YVwZ
Lwf+wDRxGS48isF03W03FHU0Jm7xxnBlz3kRQB5hUyD11HU/lOIetSPc4bw9VzB3
2pB4Luu1fMYWlhWyQyHqjWKX3szl5Ca4yw1lFL1ITgABjiebOTqyRdE7kLPk5mG6
lr0XvB40Cm1EyJyXaUgV0bwqpGO1IBVjJBh8sBUC/nsEw4KJy7XrpRn1fPvjYoxs
ru9WV0i5aarWAJyhWsJAiMWZmsZeNz4/bOajBY/UbEozQMC5Id1MusOgch3PHw2H
KireTBtmaXmbI/3Oq89iA61lMBqj+x2udVfx98xCziHDR3rGi2w1jjFHnDKqdKkQ
UQuA6BqO8cL4z3Yiy+3utfJ9+sSj7meSlT5UYQJj1ta/39Ts79gEeV5+CkPnkiiU
45z03DABx9cm82Jl3UmbM8DeGSdgU+wYCmjNLfuc3B6X/fpdvQpAGAN2NyqSil6H
tvB69FcnBEy+SwztLZcYEuD0j/wV4avVWw0Ama6Qa0oX6KjUrV68KdKXJFMPXLLQ
vGl4e+Iz6/lEnJO2ukGv3Xe5wB1HOI1CTmqibNDqvaxPy4Ks1CuYYy+g4ToIWnDe
mz68fUKvxgNYFy0v255sQod2JBVQo6pMbw3DIQDLRD5+eFTkhTf3/kdS2DsOFF9s
0aByoVnSwFTcoMu4Q98I1Zw7bX12jqzrQu5b4DiJFfMM3eKHMt2ZGTqZIf/lsd5q
/0rm0zLTpYVChmkQjO54pEUEJH6dKED3YmvM/HnC/QHP249xGc17FezoA9natsuI
jrf48/Y28i6zkiGQdKOKdlERsmsvc5PHy2brB8Qo4NbMsFeJHy6/FgtNpCjvDf/Z
ZX08P3N9ok02d29JQ2DbxrQDXfzQ2AyyFMo9sdRy774LSMXUWky/EM+tLbtQiWNo
F6LFBCYCW9JPkgHykMXpDZnE8yiVn2DYWoBHsk/seAJRWW8c+7dkKk/fxVyDYVMB
vAQ2ZGN8hXAjEFRW1ZfXz6QgWOGew605kBGZGijds9rE5ZCjqv5nPkmo3J5gVPXx
dUmbgP+L+iQqyKBNCZWrbiBbV+rt9r5TDBgkMz/Df1EWpWVlI8IJ9zxewitDo4RS
fgzzKfMv/3um3wGef4OSOH0FUV0gFfcDxqg4XKfbhTo38DAq2Cq94T625lcwbl4u
hbpHJwJuPxzg5YbLfChpcP0SAkD9ieUJuPOQfdVeLuarSkCl/jUb0gWETv9LPpQg
xFYO2hLcLLReMKj2zyAeuxtsuHfE7IrR8vp4ebgbU7WPzVuQaJRmNxP4Tb1+GDz6
DS59RQmgqLHk+SA7DVq5bGJb1ICLeyzcW3E6OQyHa8KUBae79ROop83ZLT0LXIkQ
Cl2vMn8Xv3je6huTOG/RJtl2RHdmdK36m9pzWbJH1BmFQv2VTSF2x+usgGzpZBkH
MQ4PlKk0h9TdHWFsqQYZP3iOvbyjjaJbyV8xLkfwNcjRkLePeibyQ8euATC+dziC
0dvn7g3uWVsRuQfWOzmZCYpaXsQDR/J5+ZcvVdYRMgJqdqCRgHIHWuOvQbvqHQy0
z52V5flDbhXZ4PZTWGFhyPfvcXpLxVDQy+Rf+mAICvaKj8gNV1WtmqcLDN2i9b/K
FDnQRtBvFG+kCDbA6m6d5CEeRkZFsqPk1AIXi/jRMujP7r9Z0zXP58ST3ikDunrd
6LWzcM3QB6p7n/FY/AwFP/weGG+aK28oLlOI3MUdsmAI9Og2Dlx+cyNkQa4cv4TG
p1VivYMnWa6bAMk97gQKwDOcIaSsPfbcbjddBcBiy5OarMMIsiNYBLtG5zJDP9Ok
ZQ1GbP1hIugpqkrsT5NyBR67Gsz2F3+axZLGUsynNpPLLmaJY1Ulg1jSdFVJgu3+
BNjBRuSYDMKstcXsc6Tb2Hsp/UJeYZeoftJcq9zaMlKLB00QzukDPrgref6ut7XD
K1mHylQsVXsKREqSnDoch4lyqb6FzjhQwREppDYCvKNSZcS79lQlYp6buaSHOZFV
qiIwz4I0x0SuG/B3pZz9a9WmG+CPGFHP+PSK0ItCv14oWTt4DyFQvhKYhj3s5KMk
ZFan35zAyoDVbyCkOrhBD+/8w+rUxx8+Z9YlBycyQhSHTLqwiJz70CMLZVgM39o0
LQItkzWT+GNIkwd7O5ilIU1iRudjjnCrvzApV8PnPsvFQ1vwNaPugYuGBOyoC6qO
s3PHeu25f4KLQ++G1JMne6Okb7bz8Mcr26RTe1kwoJDDsU/Hw6wOSEa5Sakd3JDD
5R10xeSD9aUSB39ObnyXt+T9qiMXrlK+pir7m/fmw8hm40179tFfwoXoB1XptGmn
i2k/Q4uNCt2jxnljZ4dLeSFWQ4RwXp/qfjeP1+11cpcG5JhXlFk9H+BxCppyh/4i
OaYzEuIYgMKld7uga0Nx9tcn6fJyCSluxPYOeHxMZm7HMS7cAcqF1gbJzvt/jWvY
BcC0fDzUYi2foOX4LhKh17BGCyGWHzyxA3HcN+KJIMJBwRN6pxZmY++cFx2gj7L1
GbHyIG2wRSr8IWwdoyth2KVlEBVxeqQTaA5akufaRsW6I3is+GvBSRVCYJNY38XE
YCUInpWqxiMn1oWU9tonK50ES80xfQmJdue0/mUd+RuQKV9HsZOPOeYrPeZInIMX
GFySRhA/nNzoRm3CpkQBs6Ph2abtJ+32VP8hHnTNq153YMu/yHvMB6NQvOw2iAWk
YLZntVMqhMroJYL4SFJRStKHYiTJ96jNyIf4wPREcSs016plY8h5yHa/UaW19IOA
tU8rtaHO+zOJa3+BYaIhCfG51w93Xrmr8YKtGXNKXtRI+XFRU+DCNszBPGdJp68R
h5EAGvehMBSPC23QazpyzErDibo26g+brxwOM2dNjZ7w84qYYi4YKEJWd0mzmM19
IxaqKQJjQR2BoURfHd6t4RQtwHgkkY5bsKQiURzOVsJ6VX7ULwe7f/4MGxkAiGBp
FpSio55H9gGW2Svs6gPyuPhU/N4CFmBYAdpZUUnTsdEn/HPDIrWOsJwK/N6cxP1J
INBWtMvL8EjWaMSwKkDEw7yhIV/ef3pu2wCE5dxa6AfTJH2sA3qNh6j8OXpH4Kzn
GV4BY+Y6HyL1XD0pS7azo3j+36fU82bJYSC+dZnwDcjElOhZDqSXkqlaF9vNRaY2
WpMNmB9rdCDn2B/c80I0H/cbZcBdEb/pIyWmtOYt9q8813oFsE8PQBq6m4J+qx+a
IfE+gsE0YkqUAss/hyyOo8jkoV6pRi/EHIqDJ8kNZ3C4+bbsv9CPhXNGxMy7Cd1A
mJ6SBLk/OhSLEN897Bv5S1ZR47YnAhG+W6vdN7slnDJ5gTaOq7r25GH6J7UNPOgU
nmlHpo/M304Ek7DiLYBdS34Hin8PyHk1PeHZRtVkyL/NgV3SPgylbXYByBGr4Zkj
A+xXUbxWFq7rv/soGWYkLeh8hwCCaO6O6WRiF88VAbqm+I6RhwbBO4OnSUvl2lDs
wO/8DRtM0y4P0EfO5MOYKNwaOQaYUtc4ROkFwDPbBCzOyJmfPkzweOz7s46nv8nC
JsA/XG7YvsCHRNGc/KxxOC27ddtxNZ8N7Q+YxU/DnwVhV9uBY1uAMFkLjUKVgJ8S
BU2XM8aXVgz8U/a8cvFz2OKYMkoF4m81ck0gdECTx+8WP1+1Jq64e2WoN9purI2e
2WxXxKrczmrsAd6JQs0ZavxiuSux3x1PIJd4BIzpVIahenhMB4KJ3n8/24sK89Nv
BdekdFup19xcTTEqOpgsG5UbHqcTENA8rHSli2ry6Q+guSkT0IXUXNJXj/NjjztK
R7VfrXeznm6J3r1MPM9dg8usQeqvdbi+6SknjeL9UjEnbx75W46IHtXUNXJw8avT
HBonJPDijwsBh9+yPOw7FTaOiL7Ez4NjraX95gjg0LaG3vGHelo5/PEbrX1a7ZEU
6mwXCjRu43ZaMXdAS2dz90zmvPh3vn4dS+LzDJ74GxaAQPTjjwKA1LLoNoO+2m4W
wtjR7ny+rJa5u0OXUZlf70DTYCZVygMCvNEjYlepnn9lBpIEKqQJ4oWZH3tqUyMd
hytD4GCvGJdKJoxHJExAv9XcGb/jI9rgV3AQUlXCnbRUUBYFhyGZYRGKKyBHfGCl
dSS7B2I6lvNysT0Q/7VMs+nG3NAbRGhshCFFw8I8cId/kXKFErjgqS29/VulA9bM
alR+xnhTVY40zeZ6/QRhTtXbwpwvG5fFVY+QRE1+5J/5wV4+RSw2sWYK5ATPAeQ+
69CtGSQ6vEW+cALwJmt5/xwlsS/uiWXhIlQUyiu6kDUAxSqqaAot8glZ0IbYgHAR
EkFcqC6tUsxc29LV+908eag4pVSjAt14oxfgEZUrcrwIYRGQVT/7UtafWgH5gw8D
W8o55bWbckNwJs3luSt+pREuoZFYZQY7JBb7DuVaPAPJTC7TRTSdLgyNPAgeHqY3
mSEB/+c6vPkujv/plaoUiBdXhwGKaB4zdWnZskJlMcS30oObda7hZFU2kM5fWMul
QN8ZiQYQ7lSHP0pqyWpmebbB9cZq71VXjRLAtg3pRLc1ltyFCdICCgD15maMby3v
aNYGGuc7guty4j7ipFFMtgln8KqZ3O1LBfFLVF9c7SDl8POPSCcY3WpV9Wnjd30y
XLzSlXnjlu3EvBWkmzaM4ghnngQLUZzMG9wR63MuoyHiPpkrRMy5Ec2/A3vCwyS+
KGmWhzJPbk0cHk0V1bcMd7Si+3sVyai9DouGbSp2BIZPwsBBlguMO4njIlvkNUGM
3/Vcb2aBZm2bH0a1HCpMcCCvexCeeN2JluCRj6e7GCOki+kQ0EtDU5tr+RNH0r0j
+O1cPzxmwSlFoyJydCmS3Kkn2eZFomb5R/UcNqpFoJ+CExhn41gfVGDKce7n+PTI
2pxGHXdIq86P8FIswjgvj/j8qoAH0fhJP1y1TldZsx/KJHk9ziJBbrzhlfIlrNha
33m3s0shssoEhhBTW+7cyq2N0BI0esG/65jhWW59ozsoqFqjujsvoeAoY+kQa68P
+p8CiPJSUe7FGWJYg3zrNVr8LH1S/Y8W2+K9aZWeGZEsIJb/Goj/PF1pmmDQC0oq
v8WnPt11rrktK+XPWN2pexDPD4kfQrpig/08Ulz9/5WiwVYRjNs0Fk5gR2ZJVRI4
VdkO89T6k0jK5NwWhoy8d+6MwAfCMlh2QjdFCDpk1uheZkMegeOhmLcX7hEE5EFD
hEgJx6WSGq7uItCZS0GpQHtIJnst8TgddPxIYS6HI6cR4RDfZuMO0DVc5fDlK0MI
xRawnP/nQ855OLn2djAQ3gsXwKqncFvblluK0OHb4O9TWuLKF9HUNYmTVO5HbAIk
3pEKT7hRuLDw2Ex32Hcy0ZCiYO9VdqdPSRCpdeBaD9KIzd+4tTNbLIqEubi5gGz/
4L33Hx3Vj0634xKTlliA8pSUfcfjGRjRr5svk1g1lBszlyrbOx8W0saABZEzSMb1
ol5NuuRPmuap56Chki92A3M+/LLH1onyeFQkRQA9+otb8M0poX87oiQQROdpsWgh
ZojqorAuCfJtLP9A0ICAs7RoB06cq4A7SWH7osv/YQ+DSqRvnA7e6ysfSKOiqnLh
+dmpQWZYcqxZvnyg5aVhgHnS2XoLdrm5gh53Yw9DA2Uf2CR/7JxP/6geumIYOqqx
1pGRB0zWugGMQayoNU4eW+MeWamI+t9TkaKzlREGgfzcaTjT5cWKDlYscciPbQ0H
k3XnFBXn7okWezBRkFlQwfDgDeiZsEvO4Y+/TGpT/eyYTAgaOPjCWmV7XjF7iiij
f4OUtVyXzf7e/9xX+tS1a7i39ILbnUqhtDG5CJ8/p3ZYUy8PGsrv0czDr8vzav4Y
LXx2dEpqLM5YScIiTZ2a0SK5KPO3tqpAZ3fWAeZxn02L9Q3ENLyywY2b9RL/3s1v
J7TmwzNY2GwBR8ONHjkC0dGX+W/d8Fa3u4N8+2FIi8zF2dUysf8DQ7fVVgoxDkrv
Yaht7XFAmLXV4NpDTqd+kMVnejDCMv0AA2kt6gWPvFX8c6G2IlsXo6PSkRv4g6YD
1bfB0r3yH2Vfgem0MAjGOtu7/ejtyeRFjksC8Fkjg9azEvvc0qEcKwLlZqzQ9dQs
g6K+wwCYU/1Wo5uY7dwW4JfvF6PLMwMibhqC3MuEdGJTjnl01Dm0lX260Pe5cXkf
GeEQlXiXTAcSv0eQQeqwkkMWUqPMFnh/98i5/0EZrWf1Ia1C3KtFp939pfgn5IBX
PL6fuOWqUaabZxo8mviepKfRg2kFiTEzeD4fDVmqVawviA+zAdwiCbiWX8StjLBz
sSpSjPtwgjAXIs6Ryzaj22umBcy3eoVvlQ5Y41fx0BpwDat39KyKTwQEl41D7ABK
HqSRybX2w09UQaoBpEyjf1qj/wGF3dF92wykNcA4JcZH5bBSjnjwCWJRpN3y8gMu
t3hlbXK2SvaP614L9WMd17WUUp1eXMFL64UwwdqdYNu+mJF9w/dHCMBPFEittmPc
DYnv+vwAIPq8TqTtFFgGGFmrU9mTigOdqgEkRiPOLmtFhH3DdMQt7R1bO0DuJA3b
TKEOH8YbXhn3B56tr79i/69iGDT6GaChtz2eqF0fArBDqoQXjxiUsZXgxZtnaDyw
M8uw6MBAWI9SqpOIuAKuF1hMvn8Y/I8vlOygCunIlD5b0p7h0TEIEKKGLgvAlXZE
MVCn0mJO7MiYwZ0vsxWj9op1cWltH5m3X9qnuUcTFbqPp1PWx02e66qA6TfjjtR/
/ejzJmGnk4BzGUkKDQGX5kSOEtgEYGDMO585K5SPlo+TJ9V0n/1EsaDr9nuyqMP2
CNMeXhmmQrPydO7v4AmS1TAObZcPe0g83ckof93Egqk5uGijgCmXk5+xqOdC24cr
TlDKqSXH5PD02ufy5iHHCGsJh723XBnDV/pZZIn8CeznTFcG6s0qb/bbF/Odfvff
P5sOhVtIAvIRGdrIOGNyhskCfvub4BFpZGWN6GRuvPGyq+TSFPkUy5hXgRdNBets
3QndqGdW1Ucpiizqzn9sHfu5s9qFOHTcoF5fVCGFCqbU/cO9mH0xZpn6fGk7Ni5D
E25ANXue8UB4yGKzjSjIbIus2t3EjCK7CLP3UeKJfgoLqfLv48EwSrYw2QB4wKDc
LkuXIBtBVpRUJ9ufrARe6ivnQqDFH8uu1I2v0/9oYRbhrmsL5zAgVWZxPI/iuoGG
5X+r/d9lTCrZWPi/mMYJbfcE8cExs/kGHP6f4+en3iuXh6rSuCrDYKhdfg8lZI3v
XljGK1wagA9xR885ncABYBS//8li/Fgy+wPLogDJq8y+oBU/Dhy4YobNkBZ2V59s
9HLDoZk/KVGXZ2InwZ1IHDED/wJqWIX3upNhKqnY7m1fjEkzCjvVerwu2Loc0RWz
/v4jZ9q8I6tfLsJJ/4koLneNVnVHUHeQWdEGcD+1dbpUNU0C0J1h9OyIMmJuoorq
AHfw6TSxiHJ5ywCHkK+DJAe5GKQnajZoLLUknqwVwKkxE3aPx9TbV+Br2FWlAHb7
MXcUn6t58Uqc4Lgm5obQENiZX3t9qqs1fHXmiA9HKvf5vLsGaGfyNLOtKQCdV5my
Bey8mAV1bLbQr8H/zZZdGO0GF2Rjkl2Zbnbit189nO7KKddx9RbqYrHy3Ip6IPhy
ZWEMchS1G1FcKYthJ26edg6DJ20D2xkDkYPBc3fWtDdl3O6N0863MNYuf8PzxDl5
H+RbgLvDngk7qUbycNQAEqSxS/UY4SBqo2yDehPeMar9E7mDbKq4h32QujEbZVfB
09aVPXA9AzQU1iqfzrOT426BBh5AWJ3V1DQJZY0c9ZiYnakkdb/B9eGMkTJqie2j
3WxDwDnNNoh6iUshykflRWF/eb6JXBXItGEOtTjmhnUapGNxuKBzPwN2elTHe/Aa
D8Wtm/BuwEKcxoBQAmywZAaqZGJE4LtyjUXJheCyED/x5duMrTNwRH/g+l5JIn2F
uKwqA8QCppz+uCsrXcKD1FWFfLHUOL86KIAehLNixWRJl1gjXKIZhHQfomhuUqlk
PenT+xaARrTppZXchoMB3O6fRDsJ2CWPvUNEv9qjkkUKeC/Yka7yhMhQfCt7uuCE
VWdOe8FFOP6C8tGwte6Sc1NZbepxww+iE8Et5VN5UkJ3LDMr9HGNzEqSdZNaxFpy
FEDusPWpQAw+GZNmXH57xFIu4H8rPwpwxVmGjbYFb3WIlVxoPjOXj3T7P4jiwU9+
1gDgR0cXFpa1Rqf+M2WVuZTWV7G56I5jLuoCFD37ktZbuK8or5JOI/xuQVRA6dGg
JVWs9vyV20IWCYuQFyjwWneqju6NLowGe5pF8SvM58EHu9bgkf77eN8hwLnkNBww
Io9cZQjNO/Cgg3A7UuvsROhBAzat2dJVKe0/QhrBUxY+CD1AMkk/Y3HpALx5z1hl
A7T3vFL6Q04lymzZ2ke/Ab0r8fCR+ds9jUG6p/0nSssc91EcYjZTHxzveMvjTHxz
YuNG3jn/G1X7fCa6kWwz6543SMGFA/vT7aB9FFZrmYpvL5vFrNfzhK8qsgfiT9MD
LJjlNnCFHYNGw3merRXZoTuMO5roG49TdwILP+vprYe9Cmzta+oNRSFuEqI3pUBJ
Q7bRUB3WVJ92fFQ/IRJy0S86W0dBRrUIIVzca0MwwvjSXvy/oh8aDsx/Baycg74Q
6inAEdeNlN0vBy8fS/MnNbvAqHN5Y7VxCydMJKVok2D2rAgzUBw9SyHUkk5mbKrS
bvBZKA3Bomd/3FWJmh0a4rJFswqyR7V9iJxeGBGOQoPkvAmNyB2AcLNarZ8HT+9R
mwzI8lInntRwnPXaZrbqaHSlwmdR32nJwBqG0F52U9Y2fJ8XKpoCpy9WXHBv4tAD
8Isyix0jdCnuq+uoSZUQ7+e0CIy28mQeSFOxBjlLRP1kxW8gyThj4elhhKcMzj9t
A3EDTq4WrpZ1gszN+bmRzKFy6oW/Sh8L+pqQTOGvSbO5eArR1JwNfhaBctnbTM1Y
ZD8qW1htdRPJvmBOudcYgGsclkpcdWtg03/VRtAeRNpDEz15PQ3kpPeRemJ8Cpkk
uuyJnMd5kCOUCbsSZaCvwBXYSo/sIKh3vLeZM8WGoU5Rna1oPvbPk36yv3psfMym
dHksDCWOGDA65EMikN9deHfpH6u1ihVUJu8Aqrg0u86JMlCKsoXVpvUUhv8ycIau
AfKHZYEYNov1KcStgA80EHWT9RhQSKdhHV3Mw+eN02oLnpxRxDPjd71YzRptgUYI
hxuo3WsVnqBHgmYjoQs6Qrs7RMn0ggapBRwdDxZts7Jz+v9mDXsp6ak6iNNGHia2
hbmDR4Ki1AiNNWVvOG9mmj1zGmLUROM40QwMGZrBN85U/dEtbKkELmwTT+nJ7e08
P/KI4nSL3tukBY8cyjq9B2auFUS4ghm403kBs1k1Tz1z/m1uKyDAHQ9tSeXRKMq0
Z91XU66I5MvKArrEb+ViHNuJB3+np0nMrE1+X2ggq6R7qveTfnyGEaMEzrKt2dg9
Gkdw8GpgBMmBY0MMh4e0NsIlkUYOUZTD//nwxupPNuTXrKXtewH+VTt4F7Q+rdqW
g8cb4FP0sW3m8otMW6PH/TGO84lWVOLpJrIyA5yzt1eavM3BClbf0OcplGyYU0nH
3FwHyO3Rdmf/e/vHDdUpoTp3C8xX7bpNjcLNikKutPWgZssP4D22XUNHChvXlJll
pRHd0+iK4W8s7PHXEGrKpUv09PShV+N0dY/TSNDSBYIzh3eptb8fQwfeZaMiA7IG
/mIAudImZsungO4NogrGnuLbvCfu8mSBHdsadFm/6fRRZoDtWX0fDOds6IXRlgHM
W3e60nVB6l/b2gT7y4xkp+2GC4AJ8k/lGyzbWkBeyvXRiAHbY98xXJsiJsdyBHvP
hjp0oeLGL76qk9AFJAP6xsda8LR07kgQTyj3m17IoKdPzdHsiV+MTbwMwRNoIryd
BtA9NHh4mCt4T1ZPs+eHSI6KfoQAW9lgqBLBMCKr58SbAumz/EeZAjGzilWCsz85
mrbO4GBpqkP6o7KnLnlo3q9OtDDs+uUap5RmPILg/vb85jggcIIegCxrllO2XNxn
q6leOmgfZbQiA1om424A/U9qywNeCfENCF/I4cafwaj9yQCTXkf0kaeQ3ylGSdqS
96PqAZeBO+3pSJBSc1eqYEch1H4XmIjKOsc9m5eKlCGZ+iAebgRSBgYIIvle5U3Y
061oxhi94ntLBQtRX9sVemwAbINyVbtKREOy9UQ1h4ozR+Fap/c4i+rMT2e4r+lr
8248TmcO+gAlbjjnzLy/+jHE46UNT+tuq1yFi8Pe2gVS+VwDJCkLmyWa4YlKpdEG
RIYDlF1yaiArGcVdBJsLAXoD/YQTtrUhL333atzha9JybSesQDnLVbbJnuUtdsrD
iwyXMChoXrEyI3jQfFURioUK4tNmsUWIypKsBZPMQO1JfokLMwVN0SGqhhFlvjm8
juQY3BiX2opTCMBgD9Yxrc9EJCk0yscgX6oFlpUGCYqWRmEBV+Fm2wS2JAMlNURp
WEJ2DyJimNb97ElXRMGcxohuNkr4i/I740k/xT6EAnBh9qmA+25bx4OzcoXZ4wwD
eyOAyvTd2+bikTdjLRxhd686+VuOEjBk9BXj6xz9VA4yEQPZ11WM91+8t1aKDDcU
y9r94n+hX45wJsFTuINWdsgQiwNeaGlYnsjX/RG04MrjLe/rcGyjH63vU/iPRKVk
W+9usZgzh8fi+8mmPuZLgAXYqtiXlsiK0m2KV46Qb1dIxrIvixXn+qecFgfbomA1
zE81jC24A1NbnYc2xF8ARmfHvmyBO1V/xQJz4Q9XCU15Fs3JnHtnhXMuMQZbIHIc
Xn/0bhnjJSrbsHXFYLhdnoEeb90mNj5glXRsi0doQRuG6vDJ6UwBLKnlVGhV7T/D
zvuq963j+KAxEyPHguvj5XeBfEzc/LoCp0sPWDsu8eh9sbpgBM4vZRIB0BXa5nx0
KdXXRyey14arijBVZGJH7c1XgZQ3I1zarfJchyEjq5dreVLUOJhLqhkfJeHIBqgj
Ejny5u/E42TTnN1T11EFCmyAsc+PKoxYjp+rocMY7JPMu6+OQ5VWfudb03fodEt7
+sJbYm09A0qjqjIV0N9vg7kmpoj1c9l2WMvSg9wfJsZEoosktoo+AdC5NtPf96RZ
XRvnG0JqxsoxW68PzCT5NfFZJdsgewdYoQgLoDxtlgTJJF7kjez1UMX9GIIP41fk
SyM1ys/4A0Q++2He5a66pA5OYjY4N4A77XjXPoDEC2Lk0iCO37O0bjSWHqoKbvJd
PzlIqBBPxGpidvmItnqh0uIbWczBeAcZ2zjXCSI3f0PpoBajEdrQ5TzVA3vRTd5A
vWeO3TjT0ES/1Ie1m/vtNlLhKS04DLYAUE6BZ+sp9VyAg5kjiHTr8LGN6XY+vFeQ
rF3qcSaKDY4R19yDm5SZ4m4aFPeI/OMQsj7n8U+19JEElJ2Eglo3jXSzWnHbKV3F
EAGA3qssFxs47HDBkHfl6dxRwn/7lBPkHRFFwBl8v+IDTiLhBiVepw9yMJpgRZet
UtVfb5OSyTZftoGMMQmMitCRKcJpQDbIfEtVB8lt8US1kMN3JBhFXj+13h25wx+/
UhSNPfAIgFpgKqgqPephgTp/n3gQ3paxXn0+1jhrvbRVhxH/bsUwqkPJ9A59FtlW
BIMbAD+tUjGttYB8YZDOOeCVWqqFzPfydCjCqL58ncOz9B2Mp0CpbAQWX09/kJSn
CZ6uNQQw5EuOEWbWrMyd3MTbIt7yEIxbdXqvdGnD+nftYUfLjbeFTcFjjrGveZt1
X/i8Evxz3hU3ehdtRrxvo272ORR6FVv83oNO4IcaINYsfVhWkdJBoCfdLUXfBicc
9qJaWpYmKb5hMpD1mv/WMA55NSsjNXJ2PIzFahJT5hou+xBhUzU6LKPjcvk73Cfa
zD2gN0NsQ4RCvk+HLEGGx0HXFhAI2v+z6D4sZDma2tqDyi7GepBaA1avRuUOFQQ5
KPWx8nmZrQQsaqKQI0icLfvGbWFdUJOHusbepemkft6t0p2W1XC1F9X+0Pc7W/hw
c+3u5AZ2zIAYlwyOPHCyvMq4g4x/HT5A/+M3AK44Bdm4tghrRVvwZ1RsXqfpnRYC
pSIKvmKiZvzVK4SlpagKAR/ApgE4nNDgojIYhi+PCGckMCCxl/TQGW4U2aGDn2Ut
hBV6kA1Vj3xLzx/cYCom/se3E3gDIDJXYowM9DsNOAAsAujiSMqorzb1PoUSChl+
EQ52YJOjubEuD+0+9jYOjxO8VuKLhYLqPy/+z2tgjZBlr7T/In7qsb8wsDQ10/z0
JZi9OL2Uw9LUJhBzBgUl/6FvAKJBQjNqnXl0tQzijNVytDkysNadgYZJ+PAgyj/Q
8ABoS9BOOnqoUxZsivQSCav1U4N8qozj/9EMNFwHbgAGAIOEtxA5UFp/sqyI/Nod
XBTtZQIbgybv/5Q6GWDVRYpI5TZ5Mh3J83NBdKRGpMYm2oJN6Uynej4Ix1xpMp0t
FXz5H2bV813GdZWUDZnl+PVJYy1SE1bwyCwKmQiN1V+sXoO4C5UTbE1FC3WGN49K
NfMgWANhZ+Nk0EqLb7q5sXicWQT/D1/7zuBAXLNZ5k4cNi72VB0KvXNgBhA0klKL
vlT8vGahZOWOXo/V0jgUlw5cpib2cMXh5T0ljXdbgt9kOi2pLbETo/B5wSFZXH4j
VgQCUWOicJZx4lTLZYIUej9y5E0lNwap8GGhigtFaD/eAja6qp3Fy5HOuLx6qWOO
1wgQrmhIPpWe6Icn8qnwy7faTSYKXMPD/b+6r0YtwHnlJgwmdA8yK4bv8KUlNNWE
3KyQxar0aaQoeUGp6iN/MCODNRz/9xvBfBQ2I6NrtDC8gywEWypd0CT4LlcIeuUz
W+pLjjVuC/1dWEPWQooA94O8e1dKqjWmcD2A1XG5UfzEHp3tFnMx9pVqzbgL7crl
5u9ikXIBnPpJPuHc92Xu7wTyGhlLoPvW6FwE3Tpsr35Ud9brB5hlfupbm+yB5eX/
fBIXLMy/QkEE4IOukkT1rJJ0sob8tTF74YbgJZACBHN1KUsQOFIQ8QYBaIlZiKWv
gF6ekoE41YqpWLNkWy7GTSam59RXfxq7N6kyrhg2AsaN9RNyzzKfbFujfUHgDFvj
ojbbl3vEmQvmidVzE0Ct4lq7uBPsO9bqlM+WbQ3qfE+2dxp13imBqhEoOq3bVLuf
gwqgXQeGtAB3WjmUEl/0DIhGbYa2A3LeyymaZe/Wgb1AYkXHyFUWqfDW/nHHB+g+
Nzg2Kk5+vKzTmblSttd9otOD6BmfUi0n4f1NvcGCLB2rfanJlIJqocrieMuNFAlz
x9/+uR+BFi5shTQ0DE1VFXsvvbHvSed093pOuX3ajjn1FaYtBTdbfTThg/JpWBg9
FHqQNtSx5vnXlQpJC8nj04KhCgm4RL2sgN3wKf4yO6no+r7iElAs/AMwI/hjydvd
3CvXxbNaUt0jxEO5MTLgm7qBmekSf56Vowd2LnaWTqs6JMyCyFvNZhGjTPc6x1Ja
AnzbnR7x303T9FaCIJNhmuEsrZrZYMkdKxpRPjtorZnXGS7T4VexWAwXyrRUl4fJ
/XsHAzLXI9Z0Kh+aQ7wsBGYXQqP9Loz0/S45E7Qjnq3Bo5Hx6exDqv5eJxmTBK5v
ujplmWeZcNzySY1qg7YPNwtsPdHdtoaaHVaclpFvWLZRgrIjaXOTqDeR7aDDuuVy
TG4+kRO2/j+OrXAUkw/A0PjiTMaIq3/m2KwX7KgshIG06oVM75jC0Jfem7WOhDCe
fgK/R8MpchFj3FwTl04wCCrJxy+uPpT3bB4ElKTrEcLcK7ACfyc4cSbbLR46vxOE
8/fFMQIY0ReFWejH15HRmWqrUvoZfl/z6tPgeRZUQ9eIdAy8qf9vmTu8bAai28lc
HMxIIGbiUkvUZnUTWtV2Zug3OS5Q2DOlTPScCxUCEP8o/txK6R5Godkd6OYVXdSH
v1CR73+GxEpPtPXpwWeTtcvkNTtN+kfEmgm1/5x3GECuD4Mgtj9L2nqG4IGJ4Yot
cGpWWgyyZ4IDr5pkTcy4A8YnYckU6i1Pn6xhrhgET1FIaSCX/gWLAfEsKzHYlnbB
5Qg/Xsgnd/zBup0Ce3jlJzsVwX9Xo40jbUSnUwco2uZ00yKDAN9bOETc91zyMdIr
7wtxelUSdaTPTIlfQ86iL4R6y28XDgRMl/woRxnNHBz6nYqii6CJN3P8O/V5nNkW
n1ukdZFz6yds4UX3XT+mx2HvzTMTP21LTpgc++nnYFGQbo6jx77aDlH25aP2wFao
JPK6SoEBADh8F3iFsz9Oqhw5k1n1uVWgx2GVmIgFH6beEtAdaTuyHBPtwyIldJzy
IQGITWahPXPHo6xx+KgJVz9T+OESdufScw2twOaGYghFTBB15dGl/GrlglcMcJWt
T3Podm0bH45OMPyedEDz764BzehCWAqJeg7MMqxb7MeFcRHaCtRD3lSNqybBau73
4u4WfW58mQefHwsm6ngFS+qaQjiTISfOdvWElcl34Q5NWih7J7Xsyc7dAoW++KCy
Waj+Y4TsdgLfONsGO+qSf7A+Y1sABAfeQqA2gm8tZpl6uroInaB9pFQjE0JKwS1x
KSbr10TzgumOwJzMg8GCZwMCYi/gIeDnanEt7kXuzIkWIM3uUlwjil+/ODvFinPa
9OR7knkLRpnGaUdktPCGI25V0IIBx+Krze0Gth4ev7o2RDo9E3sV22O+7iDX8XW+
A/R7uYRZhdFxoNpygxhxGVdKkG5+N/BKQEhXLZjS77K7IoT7sIQE38BT9N5SvsJb
lN6Iu6obzu+AQW/Ha89sjFiGPhPKIwa3AjMyZz7qHzm+1lkx3daEYV+hpr1mzDd7
SLfyJF6yQQfVY4V8u7LKQGmpYu+fISx3g8aYSEi7n2AA+jwfJ+QRZal3ztlZ80nr
HsLblwgreKDcW5cKeWoPk0lXTAr0KXlzZqdKfLx89ncJWS0muz0ycpX+HPOBgMwh
YpGDh1RsqRpo6p/xSo1ql9gxKBg5owqVN3P+o6nteTdzGeHg0fu+Q6ADK33IXbec
OKLbCp1g74EOIVwr5+afXtnstpUDilN2m4NcremFqfGW+4QTgBS81bzgxdMxjiJX
ELnFKLn622/pNspRBa8SVJOBC5BXc+hhyPjKGLflOrD9KyD7REJWA5wW7/0sA/Yv
pJWYDm9yeE139sgZRRHRsUQACYe3iud4aSKio+Ll74q7E2YX51/FHOK3CDEkCGvj
10Zyg2bTKNOkcC/dzoB3wFXZq5Lp+I6742clzgrAT4ZjlQCDro8rLG0f4NKqa+MY
VC9Mf59KRQKUdBjTPDJRzf4stjc7t2SY+aD2u8zuEEnosjm5grj23jMmgSsvvYG6
WpyeHfyMwQRWzUArq/ZkxQamfZQDBbYBGqW8VYoJWxWu9yWw+5R6xAW4Fxt87ot1
uwQtHVJD4oFeTqlRVgJDJssy9p2T4ifqH2lLJYCvQ/jwdWR72A1248zXeKps1BcV
4y0udXx7Sr2e9txoeon++Pe2GySnLPt6IZGhB11V8BBA6Yc+XSltsdn+KwAyjViq
339r6g9v7/7AkqkpqUZ5WASTlkgNIz9QN5z8ch92nOq2ZKRJKZss96faJyF+aiHN
ZCV7FkwYqbhPR4kWy9BpxkumKqLkPYdC2ENWJ9r3SgP6Gi0Jg3FRsR+9lTKcdWws
IysBWLcbtjM2BfNU9oO/AxmzWcYeN0aQsfg2vPEVGOnSTWtdchq6isDzdwNK8Ynk
RGO97HLxfuu8zYedQQiEDrO50DoN+YfXirqFNch1VIhFvB23GnodCBurqsZlYh78
CIu+NKVpNLOKVW+P5Zfzw+D9ulrUuwtR5O5kCxdo/r30M3N1m4FlLqHoRc+CfjUk
a0I18JCp9vAM/Xp2PtUEOshDW1Wlgu0+mx01+Ya+LBRyMBDF4ez0TGcjNZ4h5vWy
JAgVtcPG6SDRwpY/GN4wTswEHJs97CFO2oWQ69GLKiPwkcgR0LBh7QhEGOW9e3uD
73OwX+oEM/wAcQKz/cHtlWjWLLwon7RDwn+S8Rps8YjP3TO81gN9eaeHMrHK3d2b
4wXYYRfw6Hird4RDbobp8I125YBH857y4pWtoIcmZhgmYmwFJCDYjVCUjAAkVMWz
Z+ued/LuM3YcZ8rmk8X5K1qZvRPwhYIWlYBHEsV8LUP6aKx1VbqhymnmyT2h2+QO
3GY0fPDW4KzEdzCGgbJpto4cBxn2Hyxg63V1ooA6b1yoqddF4mzOkUjpkwY52TUJ
oAQX1G7nhwPzZ1VAtX4+h5Nzicnqvs2bVxPPwPbipcgS4XBzRuJn3HqvgGO47jPc
/gYgka+ZpkkfUFfslm8ZZkeVdcxNUUvN6DZI9I5SHc/A281SKG1VtjzAhnJw2kyO
J/GA2vvuBcc/o8f57XfGmdOJf36/OdfxSjYs3BQ1/POqKMbyOylalrbOp4b+5N45
CrtPkhOYeCkqODMsiyZStknCMtOQR06nZz90WyuH8mccqsoERy3X8TcSstMjtGru
NEQD/kb16ZOMmCvUeddX0+Ieh93va4gNlBifB2urjQgGS5ijFSGw2itqAA55/ZWS
eBhalEYn5l3LbG+yNjnbv8mm/6ciQHRibSWfcfNt/040C0i1GT/aYHS5rhbyqpgY
9AJZe70/0y7Q7MkeJYs8mX8exLOoAm8ekT/8Qg1qMes+PAVN+ej84/9QW92qtoFY
AKTqip6zeQHwHar1buf47FqX1qOW4aKANpRL7RG4Ef0QbGKdHpl2WGafEFe3Pelb
4NvvCWiAG4S+mp4iNGjn8F/D43Fk8s8HP3B0rZIxin4SHK6jIhBKKi6zxDYox/OP
CcTgdqBO0VDX48aeaVs7JmTphQEpVeOr7e4kAm2n81o5ni3WVKjwAMRNw1h0IJw5
oGkDlWUq4gN+MgiSWtQ3YaaQ1duQBC9kdHpCrZR6XpneU8LynMA6Y3s/obO2TF48
Awm9UdOkw93I/93vf5Cz9z2ytYLTEnsy4Ez1D5UqT+v9CbiIOVAiDBsJtm08AIuQ
L0TSypLtG4Hp/HK4PpzOiVzhM+OgfwWe28OjCb0ldRMcjdyvszCegt6AarLK7kWK
Bmr2NekM0VT5Wem06hZg7e/uGhb0COCJondtRoehQd9zoikuuOh2zIhL7MHqi03k
thm6aRl4UeIt2FgToeGmO7qsOn0+34fT2iJCqbWmwSg47UQtlAnzIT6hFRoUrIXg
+JpPb1/HFedwnPSIx7NXji9HwygOzPBdX0Sd0SnTmykG46WZHHIIdwUuf/NsmFAk
jJa6iNRo5T8P+D1H+VRIi8GTJSRidVPf44jBR14uBRj9rbHk5d73DzOAeyXWHQxf
WtChkOjoZeXEfEo5w6kTx+kj1dGa1mOLNUy4GtdzxYvF4N13hd92zskEDrp5LWZv
ax4PO5LSVDRUIR1Q9zkwmbOPXemGPc0Lt1O0//sHP97mjTgJAOUeJ+Lki0LNHptY
ys8d+7nm052PW20VHsrNAm7oCJWCZJQlbMkClVRp1+LaiKQjjfNE7TZUlxKloODE
Bkh35MImWiUSYUV2m08lA5NZYZ8E+v6TutyMlcQeAWBU2Vi36NNg+uLBpKUcMmqL
ZWhdprMZjWufC8BD1c+2cLBMEuDnR49sr41iXBfPMRpYXGK9MuFr4nzMY7asAjyH
7KVh2kNQnEBdcz1uOyg+Z+4EC8klr4MUDZbXf64oZJqa7s5n+46RqaQFYamsxj7R
DIjpnjQCPH27MkFcPURB1w8UB7f8cFcNC5uvaXLxNvnAy29/D0CXDKMt5obbILwO
33K8aJBtWwevQskx4L3mxRE+u/qgLfll9Kvo6jIxa/SVax5ofCTCrucSGc8on3qY
q61ZftD1+RITlwNX5jtizgTujnYHoxVi/Xaf0edZNXKlKarVk2RbJUzD3cJsB0Rd
KUeIqF15p4TiyJjHsvhzT1MKDsOBTxKYoI2f6g/CSMHlLARsYhAS6ekLE3d9KMp/
1hyI0+xqh/fU/PcQThgI55Xg1rF6zAuh42COGWf9VOPKsGVKSjUYVld+u2dKgcpp
5AfFek0faK4DLWwWxCwtzX/Uxwok3X6y7e158S3C4p0bNe4Gp6fEi3rBssy2cWtG
qV27wzoNln5U7SHfwGW/li7UbZ42kdWlvW6E5IGhX0F6H5G5AsLIhqpXs3qcwkpn
duDA87UrtYLIKhPMe2IGw4R0IjK0EXuaQlprOUS83gaVIXV4LhTCIs+OfcZnAN4r
NLZSz2w4c7kNg0XPH3FQnClA594vFvICJsyyiOHAHWO77uPA7/V0yQbmG2uvkYAO
bwTcoNarWDZpUWJSw43kWdC9bLk7q3nCCGJ6PQVa3WqDSJKzgsIObzCYbHw5Hk+G
WgFMoihX7IN079M9tdASAaBKcNt5DlLPaClHEodyMSBdmkdMKH8WQKW3WG7Dcfep
iWNqdP9HfAsD7PHVv/BMO8MLHxp4/unHsgy5UbFrca2yvad4l7ILgZ/tSaZlT2VT
VAY/HwdKdWFmGdGgv3tcxu0B40qmMI2vZ4z3bzFothwIQVaGud7V5rcmq+IdeMXd
x5gEHVuC+9JpBH2tdYdqTgpXNSKqcWOjeQwySf7Cq72xi9s9ABvCC/gpDHbXbUa4
89AEkMULSqLVC25mbanmm9byhT2+4YYluI3u3UQrhiR6o7wiqwLjbnoxol8a4jWU
4+sF7lyVCDhFKvoNKfx0hTVCgkWABy4wM/PorRAUCngQwTMI9VGkUx3Ld51MydG1
n1D4rxilju1UlJimhHQdNhiHMbn+FgYYKE/YaMs6Ir54dMivGlYH/nBa9uys2uBw
Iox+PWsad4uIjsxcJr0tJfoSKXAwHvyBFUvgDVeCfXvTDvdQYSyLjtfArWwRACJx
yUHpQwQX55BZbZT/ecDY5p0PTXHPPsC5Rz6sdVgeQVKmbT1mGsrfBD7d+VZilK08
uc7aoJKiZ7zColDqVje6xpmwbkoXUcx43mRJjnAcRbr2W1dYYNl6kTlpTeV/Peo4
RejTsApCSpYsd+x3pM3KZlriurzxX6P+Y7KULPexswKgyFqEvWSu2s+n2hwm0NXi
6kUGCj4ITtrLJ5VAskIfwE8brUiNLvlZnYR2bnpxIAInXoyGmD1oBLrycVmYCRj6
gYCtZmruT2fI/eDmUWmGoG6zrvpBgZ3U8O9a9oBB/Y3l/iY6WYq70O1QkAxvrW1H
eLFZlD3zDE4OcZHdiCFoGSDv9gSUCeAVmWdZcZmOqFFQ1KFUcCFRQ1ezgn3KqHm3
iKLI3gii2iLwZdVpdkiuFnGcCuWVnGQkv+DKnv4A+tSfDUFEjLxKtBFkwDFbjQsv
lQ99p0MmDXoIvyQ0LoLrsYy1E3ys9vViXJAnIgvvID82b44f1JFk+ceIlMCyhFRk
PCEaMsaEd6ghrXky4L7SIPfL/xmyb4qkT3Yo72lcwjA2epoOjIK79CzovDI58xlA
TtDn3OisSMgO7h20RSS77vA66ck1C+p9o7i9q9jt71emHX9Vga6GpRzgKSV3+pNR
igdJZ5daKphr9PYzJ0XCanhKK58d46h6+zYC6SeAejIVEPDg4uYI35vDoeWrObq6
1eTv/yM2lOLW8YJl06GwiP/0zELuSn5CYnOqTfSbTE8RJ7AILH7nD//psM9YU7To
LTjKItMxHmZeLF4MqcmsRReaGbCVzd4DUjvBCwqG5kn2AVe5NQTkDU4b8LBZjBAg
RQy0C80dIjKiS7c6DwOjVZ55Wu1Mw2HAKu7mhc7+wGZfmXgrRLjLtIzpOQvundbA
1bPtzpeMReRClOMIJCG8avcOxDMCMkQCvq58PdTC5Ny5bQB16ePTItcgrv/TdWQF
YERgrVyEW9LuSbxalI9bOwVEe4QmtqyjMQsZG+s67IixCccz0KrLaG+35Fo4gNh4
4AI2JCz8BY3Ysw7PIluLRWdvOTrEAAV05eZ8lTl42AoCamlj5GqMTxbbanoc9jFC
aYkoZTKolXRh9teRPNG+il9a45kxAgo1KfUqSXZc23OYRRdaMo2YJ1W6kzNJGWAX
pJyY8hysjiicY4VgC6YyzXXYczNh4kMcpRMj9eNz2hxcmmHnWhQqm3Q/eu0PUbF+
Qq7d/84e7NPtKPDBWb900jn2xLUOF/NoxI8ME8CmTRnK/L9SuCtjhlnm69m5ae1o
3l6E4cH+ZIC59Gw5rnD6oQClOpzfOQNO+VX9I/GWbSxMMJjGnvv4iGBDs0L1EFSE
JfM2PS7vOwpAnJ8Cah7m9yyHxvspj6auKBy3JU8du4PI5FnBeEar6HJbvZbImdLr
qlxQrHBk6ZdSoQoKGXpncz/59v2r4AMjCHBwi0SL2eW0H5XDow86w2EwdhrB3/02
ggVGi2KpSb4yM4ioglWxJQfG+mk7hJ630uWUCf5SQegS+ghqXhumxp4blQRdXtsY
Vxk5pQzcYV5y8UVYLc5a4/h4CSdbZiVQlXhM9R1708hBw1isqiibgZ976XhWPuMc
El6bP3c3wGlwH6w9vLHYUiUSM+GrNJEVtBj58hyuTSntRCmVvo8wpuHL4AISR2lX
jdEqqV8hQpb5BTl7NK9xKYVy5RVNalFnAZAANXygB7tYAabvAK0yc2OPUJZK7XZk
F5kB47P/0wkzHVRX6GhQGBFk5E32HEqjrpoy8vnWIrtpDUUaKZYpUOOqP+5UedUN
F5Kw5X2hIAFtKXJzrzUcUhzM4rRw74QOv9edjtiG9thvWMd/RzhMo72zja+tce+6
G8aktfyxuVz4wYJQbAX0Wv4fELPjYcdTfJu48kc3DsPDVXbOuGTrsrAMi1ixUaYc
h1+brAO844QAI5SEyGihMuzaGTSWpQAMBlTeUVUhFpn8U+3xgd/W2f5mqcBoZedy
AQu4yEcq0Y0CGpRMKwEptfCLmiBC6WGXZICOqk64uoO7rwEKySPhzCSTj1EKRK+D
+VFF3yBt88fDJlEWiu51SlAPl8HjyOEYXG+Mvm3xU41mOnMCY8fND5ZzcegaiLTp
swVLFxuelqLwSYP1586Njs4FkLT6wpuNloODC8VWIdIAwiwy6I0kYKsqKaSqXwQY
bH+Cn3Phg8SWuApx0cMv5TJ8rcf8iftYWtPYQqN4uhjrAC7aW5yR55LW7pWtCmex
k++VGOao2uXqaXAemqBoP7n4ltge16ioQi67G0Lk+mpLAzrU10I7yx/sVmYBmRL8
nucebrC+2spvSdkZndhJ37xkXoKUgawxNtUrVxBogx8BNQTXmI7RG+VRBVi/XOJM
AzsRjc2c4aTLBQBEwofIVDa6B42ZElTam7eRCbAgMhfgSSZ6VHfRVLa1r7y3GZ/S
YQ46oXvX5qlOx8MDieNnXV19isOvcEUBlY3HlV+VtWsKUc9kqzL/HBpkVBqBqdWW
wXimEzWql/ppiazd47Ge1IOeIWKW2VebXVEQOUaTZxC/QMRcEUHH5deJrv1N5+Yz
LRT7+gRuTP0iRqQcnqOq1GsO8sq/ux7xeOJH1z+xtiGiji6z0YvOh6HRwbeYFwZS
jyS5HjCl65zMufq4ZGpS/qPFGw+hzEP0QwYwzhfwAt5tcpjJSuPwLdcC5pfCECWc
rDV48KzjRW/xqfFdwK1JdS/QUaAr37QEGpqIQ9etF5cB5LpQbb//v/KO5MMpXvuO
/9JyHKchE8MVWhechbldBnW2SLKu3wCQ7Kv6q/Ngixa3c+GM8yLuS6OxVhAxe+BX
a8VICVlhIgoNeKEJCnwPYGhCDi1IA51+LgvIP1c0goMpKZ4sPdO+2RUR8o32ng+2
oL/08Me22Pev3K65sawTRC20+uNlTX4wnU3K+a7ookw1/tJTMrvNTpt0nEGDj1zm
joPG2ezHeEJQGX/vshlkznO9LDaYf6mQA4u8sIPu6xEAY10Nd33VQUKwTmLxBhQ5
0T7+YHKs9YgNpCKd0iTaleCvSAsNYO02l9p0sVeDJ/1vrYOPEFoCoteI17v3CUNY
JZb8ITBW1C++xlgPODiD3x8NXA5aNlKqZKPBdn2HvLQcADupHwL5z2XunJ6AzPQC
dVsmBDzPYY0v1uyzdg+UC7vBayI19cEiEwc990WGyYUyJyuCIeeZJzbPKobDJ9H5
W7Pp2VgVWNtXN3cAV4BNtUK/B64ha64SsegEBVyW8+9+xpf6grrJwwiVlNm8/EZd
zngsA6zgwR/JETe2XJqNekuOmLFxwuKMO6sEqRu/Kiazfe1eCe1Ycp6iO+REtEQ5
x+tOqSX77ZRuV2gQiM+XEJ+ASNJViu9UWa9bZWIrozPIBK+J0EgvnY03IlQImq/5
OOcGhbkFG6Khksl80vbyeGIAZe08Hlcq7w8XRbZ+RJVdPa0mLn4CS3lo6en1d0vE
3LWGeTEklz9ozW5+xa2Neeky90LCCDrx8GFnfc2zRPk1jND8vhfTejnen7qc+3cj
SGFRXz7eHn2sWf4zaYYJbLxvMOc/Ig0kIcJvUVmS0NFfVYv+DKsw1g8cdOcMNxka
QKy7RCSqyJhkTZItfCVm8gVqjtrBUB4OjnguAa9KRbj5AGL1V39T659J0NIayBoI
ldkIz1EMsVNDvHH3dH/ivvEpnx534dStxfMbh+VzkkNkCf5mT2gYwsSPACKWVeBq
CvzGlgqwXo7U9nW/qTl+Lh6ZnmAp5Eg/0F8kjhCZhMdZAvh/0BHMJHvDjNVEzZ4m
qew5HSl4sQvSUGi+JFu4EsX6fXAwxs+SL4WSBQwa5ouN0UtOTOc/8aWjBcBpQlh8
d1pZ2l7QPOdSknNMJW8fbNrqF0Ip0xIPLhB0V3iA3QH09vpmedE0P/NazS9VXu7O
SwTR7JK5Udf3yEGv4UWtttv4ub91R+EZSKrpLqC0Ijlp1RoVIkG4C8dFpnl7lQ1l
bZg1dsW564lTwRk1u7FafUE9+d5S9WWnQ/5HTuwdbq5Yp//v+fClPbmH1Rf+zQW8
zs9iky2JPpAuHnCYq9Nxkfvm096hbKLWMNfiN6wF5XlguFivgFW62v5jd8uliXZS
sYE6X41/f8Mr/jogMip3PMf8GGE/kkj9DsaNajFyIs5WcJN0ARr/vsKsdepjzZt/
G9+v/iK7yJwsh4NKNxpoNbMXxVNmULqSwvR3ZGqzUiL1nLXcoSZkEMasvo1/mqmE
Wnqh+FY8LfrrZcs8wIG+nrtbWzemppDJf4FzZVBgLP2nEW/fNrdbydE65P3KZ4J8
UnjsyzfFGS4XcCJDjdVZn45aiV+wsb16rFXIA0xWRz1vo7DX1fQKSLXAooKLK72o
4Nk4bcCTws7OGLcYm+JFb04KnLuWJ+2vkTvaHIb9fA2aTatqN6AmoM1n4rTxJkAU
NvNWAzqAW/gaYih0CgC0pG39Nh2fm7sdFZFgcm7rbPQMoqw4Jw+HVmjSVh/UmMi4
f7Jm3tIZRVo7CCwibK/Fee/b9hb5rTIgeyEPKBw4TbNHH3hWL1vfSOHVe/54OZe3
wm0aVrg7eMuRDqLMQU+p6fNAvG1PZUKZbcbWxb3QHgYCUTaOrwBNTtLWmCWMTaWZ
jcGf0I6/rAz5jF6Zd9AlKMUaDh6+3h3SftJw2eDenr+pqRAKSNgi9hoxN9qqk1cd
NyA7OrhgO5UTon5NfOBeWzl9h7OS0dR8m+EP654XRyCUr0W7Q9XXeZ569pnjaKrN
Uc25479aSoHKHsD9b2FFenVjlzlwx/6EkQGZYumkVPXejbwEyYNu9+Zg9necgF++
ry48TK/o5nXvwc1J2O1r91ZwU3E383Cr5iB/3/9YjhrN2mLqUOR3zuhwwUYr+Bis
YwtjNVne83a3m1fhOljDPZ8eX156EiL1+kZJUSRJp0vMlxlDR9Z83dXGHTs2rX2K
lBhs8I6vATkjCpxjcZpf4mwZs7a3kmSXNcr2kraYu/LJMQECRbjoZyTz0GbyACit
SnPzsCjODFPHjbqJ/sD0wVttKlgmAg3yORBGQxZPTf+O7rCupG1FLl0MJ8LH4jbb
BzhHblKjssKk47NMnTQRZQ4bymymvl5eg7n7wRO8KiabMy7HvWgTx6zU2iFGy9vW
aQzi6zxzVuD3Lh1gOvhgeZ45qsqFH++kTquSyPnGCPp9O1fJigaYvX7CY/bK81Yi
8z367xVvSOa3cV28ymkpKudlwuHfjbQpL983fVsaIW657OG7Y+JIz58LBlQCBDfP
gbIlN8tmQSHa0hfL79UEPFUoR18cYuamfMbSL6MbS8oCALaB5LCRCiHyx81P6F8W
4IOys4pRzRkafKn8PB/Xi8oLHw0vVvdhVtbvGvHZ5w2mII6WrGHYvAAoL9JhVIfP
REZGSsC9hr7qYzdbB44NZBTzVCNLnD0d0iojOGEQPWTJBF88ncva6tq7rayvSh0P
9WUcYswR/PeGQnRJyaalYXt6A2fYgfGSHBXx+UWqph9ppV9UI/r74l8Z5cs4Jjm9
5KevfKnK93k2r5foRjmCepyZx/Bqy63MerAqyoNeN59YjFRlwHAL/v+ngamhYmtz
Xh2OAtY49ob0YyWw6wz+IVEdA21k5U0ehcquqCfFimZ9At9+En9NUixfXSychIEf
NPUXKXC6WORhnSMRuKW6MxVVC75VV/IUHEB8bPLc5E4rU0FF0LFnrlQmfAz7XnN8
ejauisNnuj6yHWLsnLloC9GwMUAbnSm4dqypAi9vjeSG+CDZByIyEqB5l3qnpzhx
i8uT/NUB22BvKTGC8ycZ5Y3yDs4nv27zfM0q1Ina9JBJbT7imgjtXqNx3+qR1xF5
b6RiEXDRFDI3L1N6xIq+xH0d/UzXWpNmOEDR0B6OJDnr9p00DvLtNi5kQDljjMiv
tLiIT3u4N2hCHMCNpA9vHub/hiFuB8caLbeOXiGg6LwAjS26DzmBwhrvuMQuQfB6
VkRtVVkn6K7aHoTSdh0MOHdt7g/A/n/lJEPfMYAwPuf0Hg2DDOILu3zFsvPVpkAi
PIqAV5i/NqcPLDgEAOVpGAZ1WQpZAeWvzgzw59wCOR6dSNmjE0l9Gzv4tOpdj88z
aGBXHs3R8zMZz0Bzwsli4Fqh0zAXsQMh0AaWrif86vMp0/wVCBZ0ZPGPqA07cMlS
Fl1fzJl9E214kj5fZgPgDYfol9yDgvT5cGpSaZcmZBowurzeZEJDS6ltvm4+mWPN
vowUQ7SjVwplZNFWS2HRg23AcTqgZq07I3e/gzTUzFErNaO1zJ2C8PjFLCEz9cMW
kjotRpUCU54MB3cl1XzqyEb5kwKojiQasQXhOdRIV0Pb7ePaOTzjx/Xdc/6ANTWw
9zTNRi+EPWaG5e02l1/frS4DMBYWt+X3QUN4DOe545HMi7aTkJ3ly9P1uIA1hJM2
an8OtTtQdJiaaOD/16SMgdt9FhXy3rQ4/bRV3bcLYp9zl7xL/rx1VRjySQBMOaZ4
pvssaamRaHIvRj2wi4PUiDynQJX5iemBB5H9CULmKUNuaQs6G833U23nsQovJ1Yz
B9OeIVXQ8u9+dqSxLt+0QaSaOjLNGhU49ItoF3aCLJKP7xWNrk1//q4cvH73mjxG
hI3OkXAsVFDJLNavDEl6CPZW/Jpvjekz7pVJrWJDT/tUuobdh7mUsNUDUbbQ5Upt
wDA+HiG81JNwxFpgIzR5BzDpsyRact6G3hcCepUngvhyRW91bckbq225vai3Xa44
siZhZ8P7Gv2XHh79eA8k6/lbZ8j4WtDJ5xJW/PL0qYpB5KGoCvt5cBC9sgWklb7l
F74okp0b1pF1dURsGXQZHZpc/NVhZI6LJxFY2jMwqYE0+Fkk9jhYA0Rq6dsD0cML
LceFBODHi4qkC2aVGNERBlwVY9BfmjrbQoyTd/exriXqY/ZNGpHr8rQOmLwgO4IY
Huu6FmMvatK4suh4TF9AA2WOUWJGFMIEWAFnS42paSjAGMp3aER33Z1LpR5UM3gj
M9exZY5arABXFy/+VljIyvgbGOBZ6ifn0cEpqfdgO3b/ef+UGOleq0a1RBeYWuyb
Xr0s4zJ2rvAyz1hHLYlO7S927tXJHa8UVx/zaPJCH7nQ+nLgprShVy1lLGyXCA+p
BhAUyG9FIK5PmWIDuD5jLvnG6Mmj00L3wRM1Jz52Gv2RXYm8Dw2YxmcsNL/nLaJt
BUHfJiHzD83X4Yurg8xDeKTv9GQLcxgKYwkzT/kmdVSnwNcnCz4gp3noeN9ZjgO3
QXpKRKk/mV3Qp7Lz5FyhCVrDCyiRdXHrjUspZ022ffvwN9LxzD9hMSNNUNuO/tY0
HeWNkSNS8sDfWCKXK1rpwVcyNOK0GdLUX2BeD9th8GbqyrDG4FB9XRYXpq5E3EJK
yJxbqab+4X+gIwdM4alSR+2k+4MGqO7DgKrS/Ty5TQ5ZluGVUdaq3de7UvqE8o4W
41Yv0fuxd9RfBpGiYeHOUSVExTkxa26l+TBLq0qSLNJKJUc6Ep4U6HGagyolSObS
/GYmv704TZ4IEU0yq16VC92B+GtMwSEWBsGOE7zchd43A5o+x97WNGbQdr0VSos1
7q8hnijGdmmpdFAlQDxr0Wqd3/Zk6/BP0iORfBpt+pA2+QErAXFyahUWTIxIwVLv
3rj794AWMzJXhe8Mf3aJ3M97Zab8w8sJCthIZKj/QdXf5+w739lTbEmFoOZVX/dT
Qh9WchV1/DlzDXCU+AoYW3o/MX3j2mwvktPclA+/7Ak30xxNWIZtqDWQrZJL5GLR
Qm0dFBTNWRmhMS2QBJ+3S5xiL85mgfYXhyEO86RT9xgupRFHCdzJ7LyDH7FydqY4
1i6aAorHQ7ojfY48EXCosYwi43mVnzNU5JqD5Zq4oboW66SCznxRN5I9blX6BP7d
jDqm69Yu+STfi41Zo+qRmltdtaaiIhLbFJpqEMOvNxMi0FQ9BZMUF/YtjzrsnLKl
O+7YU+Vf1KxNOlrung6Zo0kOiIZF8J1G9+Dqe3LnRe94KejnlFWS3MCOFOkAmwD7
az3J4DinxECyHpwofAC7qAjHMmwOv7KDc1NTWl7YlaFLirlG5o2+6Y3INmHluaY2
kpT/qyYmpe/ztwNqbjvDN7nbp664tQIOZYYr30lZ3pBzufg74vUvGYcsHTAUwDKI
jZq5btZxod5cHZyWp4g4A/dji56Sa+C3p2hLoppHEwmlXbZ6GGZXurD2KwF+OPqC
UGW79Np3gRVbTylBxx5nSdNSdCNKqOdr0WV4c4vojAAq2J3D9zPpCSVKaWRepQfe
6qLLxjCL8sdMvgK041q+JNsMIdEBVJ6+XLFNi1NlgI4jd/l77Halpdc5ON2oblvM
AwBi2WCvjYoBV1RigaVID6+BgL7Ue5+cpU7t/+JzeFbHPymLKdoKLR34+xzqxoTP
8gFqah+26PCvw/Kg7IKrBiJ6m/fG5etKn/NyPOZdHtyvm2MRHkWcIwtOVhvuMvZG
miRvNnOhxGkMeyTiBtD2XDsf02XVtgA/ZiV+5XPRUsP7zYYT6/4U5TMiInfbEZk6
l0YAGFqRGmVeCoNh9yvnvDJk4TRxQryWStPP6F3WmVvcHgX808Zu9AdUBXwfAlAI
atZjY0LmbdPmN8E7xqH7NRY4SEwgv7xAzFQrxwggM84fpzqg0xthTK4oQfLnBv3D
m0Smy2/NzeHFesmfz6CMYDjy3kH9k5wwnR3ZBm/1XPPf45DigYFcinN1c+uni9nW
9ue06AOJMwfuGXdTr74f5Z0r1mzdGx1U82WkOvQfxGDVQ6nxzLfYTyFIgm6t0w9E
3xbIx2JWUo2+1qJuA826jZmge6cUCHMq8appfNo1jBpXkwt6s1CKlbT2nWdvSz3n
jS4eq6/B+WH73u/KShcz0ayzA2YDpQyZ4oMcgGjrWxHDY+Su27FRIVm3Xie+lP4x
4/HpjXdusYjvlXHsEcFoPoNKsXk5ccazHs+lrbzGjGPBHG0k0gI6DuKbLHoajVez
sOVJFYqSpQnUgycFY7XbAKd6G4F+cPhnl1SV1BGtK8Bnc0Ii14lnH7dFLIASEnL7
L8EVd3p9kwdvVY+ZZvZj1mabCnwXThD5s/pgzQw/WgOEi61ajXijGma/JU0WXqZk
C4hhg0Arms7OWdkv8KMjak8PxJvjhjr+xyIu10LZyh05XpyVsHut7/QeMs6iEr6g
gebbIs9ztz21CThGkxgvyYuXASurfUxU9OEjAh8RYTDa/AB4rW8v21oONwV0NwkT
c7qWf7mmjAtBVe/nTf2YrqN2NGarX5QwYyPMa83Z1ff61FKpccW/JinK3ojt4hBR
tF6Bn/1GNvgyXsxq5t9z3qeQUNcIXSCL7hiNDu3imO89EY4QkDwBIXXXp9TftgFp
JYomD3IoLK8axkqpnZsItho37+lwlJrqMK/l7QDNyn4YUjZ/u8REbymPJZjbir08
tEO/Ehdjzs//8tvLJc8dj+C5cCkJOhq4VbTS00KuBztmbEPlm/PjEedOEe0ofugj
EomAhZETGnmpB8tPJFpb9Rzz56FmE6pw9oVMQ3fRoPeaYMj+gGbLDzJUxGRdJ6c4
YsifdjGPPYNQAKmTpkqMABZNGH2RMNLYxvG4KTBesbXqIvTJijbG9BkWKQOZBz6I
SPatoi0FjFYgiETTIT4QO4rVjAcTWbsdGhb8/QF7w1manL+AJ/6X0yJADj7f8Zmi
xtmBf1c//CXWo/20+J30TcybBe65HUDzpDYwPSez9lTbvdCMH+a6TlpUZWZk5T6c
vn/5eIB80riT9qDr6OVBJzXs45xa5oAnra8qFTv/45m7uhLPNyhQnDxx3KrQ0lIr
yp1Zj+k8zXZbFqLR9u2P1O0RicO6u+wAoG1/8dHAov1IrIsbGaiHQiYTliCm96BJ
VVFEoQXihC56N+Yzsz6o16gQmNRSgXS7dhvpbalegAe+K3FPnRbwkdXA7As/vPRR
QKsyN4TkCwFuZp8OeaLtvWR38frKI//DPj9yiDBwvXsXdzK4TjEyuVaNN0eJGay/
g68g5QUVZjADJKaCUDN2ubutVnrJ7FCB9UNdpc4vbgxddIZIDiFBDa8bxIkvWdMe
5uyYvqn0lHSRYql3h8wAGwhjDh+L25a9/dz/WNknOVifMyC0D3hEUpKz4QGRNHAB
wHqO/U8uoCEKThmzyLFXLyMWYBFgJOzHTz7I3gJ16SpE0gluJHbQmUy4kHYdm7Y+
UluxsZVmCJJrUoivFYc/+0hAUVDinjxpqw52OCXlWy6Bh8w7j2T+o5SkmHC7+/MD
ph57azitp83LTIN38G2RHfCpysW0VwaNoOSti9RDB4ma4Pu2jdC/ZE4yEktf+iva
xzJGl/buBSZWrBxHbh2z6+GW0bh5PS6sSGtqr2Ju7qzoAs1hGEyZJGPCKruSyLrZ
TOoV/hCY7/k0YF4Hq8xzSWru1EwPNXwrQk08TkOkxngvZYnjV5BS2u0bu/Jcbfdv
D5DufGqvTRWmX2iHnjkPhXwqzbTwWgfMd3rbQxWfMp7cD+KmcBT14zi6TlT0fsJ9
YfbMX82MfapbMAnTCRZjOKAAYx+Q0oHrmlPplBOdUkhhHECUG73oUoPcZIW0jj3h
0Vq5rqiQVm892xkH7R59v03fqQ5vQ56zfUUCr5n87y8XlMHauieKdIcJ72Hw8dUZ
75VmFXgu28grloHMqfLtpSP07rjpV3q9vDsJ34+cWhzAVXCPMvHaqbScyxxX7tZA
ieS8NUh+4QDKYQGwhrXlgfwj61FNqBZBFWQ1FW80ZDuQN2Ig6H25jzOIf0lfmz0M
thkK0TzmdGK/4+je8hP0CoCTPFWX+DwhBygzb4vz4ovBgdeZvzy6CG1EtuZgivx3
QPcRvorkQ9XL96m1qjncEv0N1ro8LOLWqj8rG3I3AHUbpKNtMZOJMhLL9sn3onbY
ekc+OUUhZ8JCsvxge44fv1sFZjnzz6JMooP6Lph25WN22kBL8mKTnMAu8leTZTD6
9F4MPgXs6OEWroyq9jMtFoF5JJvRhqhbekHMrGugQJYAHm6x/IEn/EjKoa8o47lA
4O1Eg8omalfhQwqusiNE6Tkf+xNKem4bAyfPdw6EmTLG1s0pXGxez0jZi6mBRLA7
Plx2L6v4EZN2w9yJ61E+IgcXdHwP7VqHFRYONqqujIM92NPot0/JBmhYAcnRNd5m
zcCHX8EhuGz2dhfSJgZKXynwFyYyPM0q5K3EMHRmRPP4jZXT0AQ1djteOW0nvh8Z
MYU0AswjI++4KeMpFaE+ulQ2QH5cUEHo+wKVu9qYzheQ4KvdN4eYKUufat7y2VLb
Nw7Pkif/ixfoat5pqA06JXw4PrKxDrEAyl3Vu/ncQGhXCW+C0s6D/mVI7/zcu4/t
gaL+C2MRCUBYZi44g4+OCcasDV4qBKZSyDh4znm9caYZjp1OKV0k8+54grgoSQcf
ojAi6H0RsilUO96IFzPN7uLVIHmyl8bWLolNnHhogOIsuhZI3ynPp8bAG6dlqoDE
euxtvUw+lyEXY/wvJCY3Wiwr12Pvzpy1ybclWd72ti8vvKAyshPX+PfAy9SnQh9e
zFszR3kjNDIciD1yQy0kD9qVF4KRZFqK+xESiFt5YkpXZkwDeiDYWVfL7XrQG8FE
lDUs7IxHJ/Ss56rQIxg7gIE9w67AKXaIUj7HVBwpL+ZEmsFCmQenkmIX2RFrd/Fh
4xzbLsEQEQr6zfa8G2aqRj05T9B8Z5wG8BisdI1y0qoPplp2QfOJHpUsNfuUJhNv
WWHUHTFrZgnZmvIerznFDleCiRprHSGL74ne6kGRsLE647JacB7XNqW3yQTlp8ZB
/lAq0bYYcArI+foSK141G5u57MSzL+CoOKQSzrQXDVgQusnhp4sF4H6Y/sdboaOR
W39V9Ggw0xfNnJAESNCREK/5wPm3msqcS8MpHZfK9fokEnIRhIiNymv54ExgGSa3
xO9NZpDjzw5FkuHT3XJLznvjbRrgJT79qAIdo3UtqwRXSiUechx0S07M/lf/kjE7
mzftM+1ccdqOEM4uChSfYg3RGrx4NlLyF7vm+EcOAhIRpwg9czmVaFsFwi05Hi+E
YTmDLmDVGRoNMzBpOdSo3ldrgOvL51pvJfsb4L14Um/wm8TPjKz6MoC/6syjR485
jV4iRleFgxpAuVz3BF1M2Cy7BOTI2A+UdH6CotEGF0I9GmVvDzMfYl3K8XomTOBX
R002MsS6rQjuFyOjIznX9qX+i6ipDXqNgdxMYRDUlO3duFcUrjbiJNjCOnun8Kr0
WoieDIxNi+jJjGo8MOS0PJONDNhCw2fUbAPTzIiFaAg4zugeTmhf/tPWO7dCUA3Y
OwHA18JzLqm7SMwACR/pyTSl0mB1OTW02rJq4nHB5u48wGQHDDaS+XO6op0MySmb
sjrYE2qY32MsYhQba7x1XW2IhIZZe4z9FCNHyBz8lS4lkg7pkAYuheQHfs8wCXEy
jdWDW40HXQEinTxVNgRDvZxowjNm7ZmF0FPAoqIIomUtCzmyU+wtWb2cCCrdNYtW
04/uQF//a9lomzSFR1gN+YhQ/YW1VpX7WkYxKq7OlVP8BxhQTL5CtSvAjbYMLZrh
rys1y1GQiRsmRDOYTysA3kpNhaZcKZq8FLZO5o1nEpzqOd0sBsEJSuLSx+nC2SVH
HqkkXnfRrCsoYxy8b7sNK+Y5I0aeBTnJ7znDdnUm5qsVa+ONAm1U/q59l3he1EaV
j8CY92rH/XzRhoyvj7rfzTZU/zBI2mGMG5gwDnwuDGLhHqHHMz0Urvv/DWNjaAIw
e0JVpeIZybpWRdUABPAism99QjyN+sw/jytbvjrBXDOul7JGd1aCnBCz8tb1uHQl
GejVIA/Cn0vtm6UKqPnycFrdq9jcgbA0u60laXKbDc8oV82hLQwmX3I+7N83zhRA
SwIjgPaQmfzyAEFZxjYVRrJhVb0zs3uCBhwabFZp21tho0RoQN4UbnDbfEI3tonI
SPmRU3hBvq983yQbIBCwvyPBSrfM911Jig5eBMTKVgDWw7HeGndayrRfALbdfhhj
AqaKZE+IU9mk7ZlL3R0Xtgiwb/EGRKKw3hBWbLs0UlBZStJEvN+iGzeQWkIy8muY
mSI24IXZZaR2XPT5LwcOxxsj2GDVFFGYQvTa6bTIeRr+zo4r29rZZvLmePwHVXKi
eR7lFCUKegJb0v6nSDnpUtPTuqZFcuG6Hb1FkJUhGe7Ya6PwnOnQO9Iuv8Y6RerQ
8XT9RCGWARgMDjLlKJaOYC0VgGlxGWV0pPQOE1qZmWh4D/0nUzYwMqSA+9NKKR4l
LhB6wqqOk3ULvs394rnkwIXX9vpfrRn37JfOFqb9TG5y7iRIqxamv+Vs84jrornp
ZfwG6B4mqTFMJGmDG9tX7wVU1nTYXvslp4ZSbC4d5QEBwhBekJiJYFE5fQgkshGX
T+J0ZwBinhyJm0YTBOQ30Yt9VOvCcNEdxTkxjBX0E4Fr/ggFlv52uO/oImXdRtU5
c0zwJD84kfF8l8LwhLWBD+l1UXiSt7x8QPnmcMKIG3RheatpAv2OMhf1XIpKzg0N
uvkd9KYqBE4ru4Ay6Yg58Aj8VNRB/3lmn2e0LA5BZC215ZGNrzzIrg66VCtImSpk
m833jTVKfS9U6L9y8gw4hphfjeULJYNUSqw49oZNXr0kC/vU2Wl/MwoHZ1/UQJRm
yQQiRqggWNR0EC29C75Wunp93XSFp7D1PG9ON3Ax76rPRyCit6GOsv8wcdY8e/OT
b2w4VFjZfNtwcQsfZcLvfiTAwq4cNxzmvAfrnSYSKIDYbjoh2t1uoPHgZV/3reqC
R0NO4WjET0pFnuhpRT23SeIQNx0NtzF6DgPOoVOCnktyjCzfM3dbzv+hlv+vBLIS
+F4594XDE8jD3C0I1PwpsQKPNutV59DNPnPqg9qy8Vq/Ee4OYbpAcqMJItLEm3ip
w1tAxgLf65DTY7TvQyGFN3h3Fu+QvrVHXa8r2wkZi/ymFF58TcrphJRQ3kSENpnJ
rlLGLj4Z1ywFiJT1mHTeSEQQdeguD5YT6WH3Qc9sMjlpAobjABhxNm7bHvRwjIQA
ikoE3drkEpDFguvKC9XyhK2yvexxQf9Wyk1DX2uTM376eiGjGaCj1iVkScYvlEqS
RnShVOwzAX8u9nRQKP9DziKElE5KUMHdiBTsRnynBYuyWlMk6gnRkcn7Kyzl2mFv
pq5UXifE+T90b7Xpu1zPDk7l0mYfBkf9wfgKdxQjiPL42co9WjYnl9KKT/QUMP0w
1+z2NCW1MDHcL8Yf8kW1iyW/wi/Lyw0JUw8e8Wfi/GGyR0qUfFZ6sYGDxGrjSXP3
MWMsYWofhGDHv1Rjfqn2ziezVaT6AA9Xe56ZcZm8j70qMGyOlGQVsvkXWNHQngrE
YZLGbWWdXNlhz4DedaPxo54RlJ+glARp+bLtKHLaFThUs7aff8PviM7S4oew88c7
HZzzmatbvhDOLQskBBMmvIz3mz35xxzEx/rUo9Hq0fW5dCo0zSI9RZCFm8SjcR5T
cRU+iQyhEwDn9Sjz4KcOz5duqsTSDDfVPCszIP26I4sDtzRPUQeV6eF5skrlfE/1
lGE18nJfFo9dtP1GFwIQxMhsOZPudPrkqwW79nn5X8cRt+gCmQicuKuxfJH6BT3t
PCYf12FGIgLKMXKdzdN1dYuLBd6EXAj/L7jlZOjW+SIclOQQAaVtns9qXYw9X/Vl
/oGxkV9nJnf5nuwzSXiauuIH/zpbEZDRsGnopx//49uonNrY7AmYRF2fzYc0Zn8g
nF4wPIrvudNa3Hp/LhJq1EJ4p2luUpkJWZilhXC/NL6N9nIE9/OKTcqtAVa+nf5I
LbIvXoTUkvikXV8gnP103yZ6obAl1ix6vMv1bnvzHzU1QQfCwygdFpk4voNtFV/2
9B2hiA8498kzIyuIkXx8Y2+I4PDMOTJG00mMYKyyuRzHnAp2FLJKdIiSyNXvIRYF
AMYHOc5uJbO+xvbZFU1VwLklHM2AmJ0UCLJhQzZHOjvSNfhl8nUlFcJMwZVdB46P
uCnh598EMQ26OhjYmXTizu2WC51WCCxemS2octbOZkDG+nlbZ1Ud6Zx7qbQEeoLD
amkcmK8AeZHsiXsJI615sjZBvxfg8dG0JySj7ig3WG+gHSEbYJDZtJmo2qmq5oXS
WkUH5m9Bf6H0UxM14f5JHGUSxXgClyelMYYqd/hK+WD+sPE8VdGp4dPbfm0zZAjx
t/ys3VDGIxDHkIH4fDRCqcPTtCdJBNGIz+z1CD6UirmQkv/ZrB2vgJbmanyeviIa
BhBQped9MCDMvC6QOhPoZ/MbdpryI0vjkveoiNtsF5HZXTSHwRlq+KCIFNwCXJl0
8iJkNlDD85xZPVeTXghRPiFXMVS0LKSdyU3RPDMJdI+pKfxlv3bDV2p3fXpvgXh0
rLxd0ReLMib2ZhZhiM1d98J/AfD/zn7q2CjBzEm8hBT4f2Z8cNU+kZyWDcW/WWpk
jwOA2/VF+dY2jTx6MYU90ug+HywBUPzqyxJONCByZxKBxOv9bsuCx33xqUexeZrE
hJLQ887kOJfh/3x4+7L44nJBgI93o37nXRet0g2nmDQCn3NP5IyQZj9iG/sWGa/o
d4AzHtYFT1lu5j8KYt6MiVqq9PTbcHUAgIYAethjbF3lIlSaHDNachmc+Aum6Wtf
gUoA44XlEa7NldgdzbODqg8u8Nzu+MCJ3+k/nQfAbCurnqNd7WeQ+z9hzb95Hr9f
Q/OzK9rA6/bWdCL5Qrvda0+FT+DhoiQfi7i6g396nw6JarVz4f6F0gGCGBifFhSl
sU6DmcMNlnIiKwSj8QnD8Dpb7jUkY9G0YvQM5QDeSaAfEC71GaVhc423C+lBNLGK
nG6V0pHyLr7lRpHZC5K1sH80OB3SLi0SOybbP3FtjstrEuFjW6fMVUa1AhvmbKDw
RMJeyNuQ9jxcao78nOAIFJPW3YRi7Gp6CbcQOSAquFZkxL+HMliO7/xLBnNyFigh
ttfp0LRtBVwzkErLsujRuSIKlNRvvDhOxdKk6UN70MPK7HoTq2fGuibaWnnJO66m
fkJuRUJ6LDfSunG1G/aFACmk3gd2ZjZtSlWE0/a+DOV1wNjcYagRg8SVDi0OdTDS
1ymINsXXJsSm5L2vbB7VYbXEsYtKVloMOXG/chKP3jLhVp8o3yCt0GkSTe8yQy+9
mFXdMIMSpedvM9AwtGjtgUMudXkVTAaNq8DFf7VubE5DC06TYCs0nwgj5CPqx3jB
vg0hh4cXz8zrsZ0EpurSw0vyoys3JfrWTwiF3Av6MqubvFy5fW/LoYU9WXIbdPTA
DDs8IXV/hq+b/wyaRsZEgGQhFGGzRzVFXcDwmZXaUoBFMCWQpkgG2HylRO3rHKTL
yVI+pk1gLWBNHRn4OUmYatvwUzg8rxqC2hYc88ffqJi1dI+cAjelyM7GZFCtJVSd
jaGkkNVNU66oMcHbM8w7HxvwB70Hpf85vek2D+poBnXqp7is+4loVPaqQyGfMpvU
UFjhxuXwsQxa9YZM1cXCnyVznJ2DwoGpNDY20FwJLpOCtxb1sQBeuhQ6CrXzqC+m
l7mBzCYEkh9ytscS8BhABjuvh43MZbw+zpJ2Ajn3/lYFzaS7bsfMmd8xMP4WtJUJ
/JOkwkDjK5mOyAVht+CPHCVPqB3dcpSMuMmylagIs2QHkUZFzq8yHHk03VXBcgIR
aCFp8Gmb0By3by48qb+5poyh+5k82dv3DWWcQZWqVH3aJC0JsOG0JdSHv1pS9v5y
Z8g4I19jZ7+3Yj3iMVtwGxmBE9JkABNpstYwNmcDtRVVTli1qt1k7DaXO1H/Brvs
eRNVO2txTokdasldty5WGguqYUQmcs33laBF9oINroHo4o4oiQo30Ra5DJSzeKKI
AIe+O2djoeiqHffhsL7RNPQpHvwbeLXhoAsBNpUM8PrPxhHw0aqYmXm0Hpd3WRq6
gOyOgjSlrpnX9fazLMmU63f2rJ5uiRCRq8jn17BcNKib+4u3dAkm1H81Hw7kwebZ
nLz2J7MkcXX3Y4jwDXvK9Wku14pDnIl8hoBlwn8EEjkppDMGZPqyCkdxTHwp2vj5
oh3c/gor9rycHabZV6t9Y55b0lwIGFc3Ut1FfMnSUd/xlq17Vap7n+wdw7h9SPms
6SUItZ2TXErDVvdMrLI5J1uUOubilNeB89aVKSakWsWXUDO1/r3fiZ/J4Uux0K9x
j51G7GTwrq094cBhCgs6J52bkNGjhTfKnFJqUaIbz8AzKtU4zfFY7yWBQZjcwRP3
20P4jcDTJcgRRQ1ITI9lIoWMD6oxMhHGg4Ep1UMKi/wt+hg2B/tPkcpJhzG+zJax
vjstLLdyCOgZGGBjatFIRggHrd1X+dC3DH1gNV0TIvSr9QAnoMIYZvZIpKuSv5xJ
rqO1mKQrW6Vndtn+p9c+PWjSCuPGR3Bnpzdloy3FnpPMq9o29CF8xnWn/gG02Fhl
aMb7oSkeMKukyMQo6Oe99el1/72GK5Mrw1c0ES50K+HWmm3T78EIAGYUGL82pDrT
HTtJuZ2MlHyusZjz9y2aODUShI2O67rdKIyWkWDNaTmZE9ntZnp0IUzH/LDLKBse
nqvPnF54l2mEjvQchQNx2Ptac10Iv/84ag18XNbab4ntTDAehqEvVhC2q78Uw6tj
G0BF23p9cWRKQO/GKfPuUhT2beYI/57T8geNLaJJarQxVRYOKQ5ryr7iyCAHL8XC
Q/axm9uNlXV2UIlzZCluEyiWEHrdwlx5qF2O0zelVjP8HxqXU7avkP/up3JRmdPK
xPUBaCsbBg+EVrEseFOpeJTxp8WBbdU4L3TYx1nX/xBkJ/4ZOyYS1sA2+7pYad5F
Hs6HRO9gSjj1LF+iEwOzbXR2B2/5sxePZHDIumv2WuTtYTZ95AL+DR+7kMefZWhm
tbfSq7iIGv/eykPTjSyfXl/TFwVLbnFM7/ZO4FTBq6rN58YqaDW9xULnH23m4GlO
5W8ZAX4qbsX+n/hZdGOqIJjYS2jgvhMwnxho2R35PxWimZhzJT+Abxt4yTwjxYtl
mWU0rFkJHpI16c57bXiEtlUjKtBwNiGS8vC8TlN5ZIXAArvwN9ET2z/ntNDRHkpC
VJHfldoAdsZIXn7t4nUhMCOTHTsbtydPfdFnAKWyIWIfGwf2DSItVeCu2tfB1wuV
PwlIq57WlyIR4tIuxrTKKq6R/6k7EoQIhp49cqF+O/MMtvWbZ+CJH2Bhh2RCgyxR
d/UMjBp+NDf1xjZfLMCRZKQ/bM1S5IWfbeCG4igZlwO07fJizZKHUtWYP2+G7Vlz
ZgkNZWEb5kNNKf/gR2ZWzoodsuzroqlOuyxG5EMLDE5T3FpeKuofGHlm7qwD1dKr
ShUK+loo+tf7eqLEJaBD0kjXmByEhFYrSv2Avj2CkA9Lh+l9iPOz6hPbt1+TI7y0
YxWIInE9/6Ckjrofr30tkaHVQZLrE/Q9OROuue3KccZ3Vz7xlmi4VmDX2spktmmZ
hGljNv3OBm6RAyEAeypm5JXCvODdLBpfVQBqDSQKqz/HeteGI5V9haU2QuSzEUvw
61BgJ0EbPWFZIMtzhIxpemwYEmlvt6S4V0qUFoLHhbWHblqNro0uQtBB1KDrNrz5
ZKhSoESHkdpHdMjnTyb9Ix1rj3wiOrrFvWIyfhjdLLacBCt8nCYUV+Dn7HtXbvQ2
nu0hETNajLLFhjdL6Y2LWwuEjbF9bZc+RsP0eoE3fck5klD1XgoT8SxK5dCE3m2E
9nRzBNxEZu2z6vN8T5ONv2EPraD1Wuljf7kqcZI28VTdJ4BQgliOKOYyaU6gpixM
HIVFbzUXkTgNFV/E1JCTOFIa3mWZz2NE2e79/7xfu88Rjs1NfktoeDHH+ayDn+uf
dsz1mVbKhPOakztDp14jpzw7vHqEiRVG1WY+eBPIVzeMkAIFD64g49aL+ZJCKpWc
ufSi3Lnnh0ES8EoUK33pUR2gJQKeMeBbyATi93pLflky5bKUpd0jJEOocq/4S47y
4vR+A0dmAYaseGa9uC+SrA6R6t6S8S7+GvAwKJUAQotVw9zeUCHtIgFAhn4izZ5N
QVCuZWPu0P4Of081hmcu6VlYrnzycI1iTe2QqXmCLrkcvZ6TwcLA9dcFWtquEh2x
c+oYoWzQXutC12AF7AH3rR4/BcICCWXNu4Yw8f7MQXcKbMEU/9uoeMnteP3x2Szy
CLAGpV9QhgLqlEn+2K8SSrPGdSyIc0tQfMeP9EoRgsUh3Ma2MmGntoCzHJ2DCsym
rQLW/yF47xA0kn/xV/GR2myNybDmSj8KhLPriBsQOy8acsR33iOUU0Jad6rxZ01I
f46BVaQoq+Sifo/2sBsiYDzN4YD37zZdy47ozlzVDoSSFedG1iH5jvXMbxoQxbPx
WW2uO3UaNS9rPQa8XGjQWKKWhzL6D4ulxVGD27PhUXzQ1qow9D5ycyjwM8xYVUOb
mCboJqNMJuIR/X2V18a/TVbHHKNj56AiPy9ijkqCkjD4ZvMdHcipfIIVxOczAoLn
FlgkKdravz1DCsaROttqHrfJL/MajE407Otz+s77KM4RzwFVz1JtfN7sF05J0mAb
wY9aHh+f/nUwsBT1QhHMeKabN2sojhOdVhQc2bEOtOxUVC/iXeU8ED1Axt5riAlT
rNd3o6sMpGUL+kwX2spVAZ3VVCxOd4xDOJ4r7bWRsUKip5JWgzZgWQKlRGN8H4pi
xwvCeHzeOxrgwBW94tvt0v0fxpbC3rerX0RrF6w9gIp9a4cp/ylrJ71GbhYBSOlU
K4YkHDGfahndBAKLyygq3EvRwqPDXICIGoiVFym5VI8aXmsqd6QrSl6QeMttTdxg
JCpALDKeqFjcklAIMiyKOhJweUDIPcQIEzv2aKvHz5DTwUoeVprS7Lm1+hZF5+6E
gSxXfpE1g9nkubbJnER7SNcGFb7xPAjflgroWNR9csnsUJh0Avb30BCpqvV09p7a
XXR+2QbCPX9AP4q659xCxfJt1SPjMLHpL3BKl2rldN6W4N5JRD/90rMM8/Nya7X7
NVfQxxYtJNlQmE14e1JxlbkvcjI7Ojj0YQBqm9Y90+XTzf7h1mky1ew5zdUPRnxM
stJvU0R3WNYDqPtD5QZhcZ72sluI6s51n2q5nSLCpaT/sSqeRC+YsprUk1zE+Tu3
xzhqQU2hd3MOkoWBeGGkUzcd2QEfILbebgGcdbO4t91Uj7X4MSRHs9opCsDFLaKQ
wwq6Lg6b1PTCLfGaOnSVGjjKO75d9navZF3Emghk2c79uZOL7hZOrAL9r+l8tLSi
52yhDU6b/K4Al6mrygk+tLPnWYrHli6gDXBHQlO854yRrqeNQZBVKVVYPcxOnsRx
Vhc6KMxBji3O8+dF4Y8whx7Qzt04MuaVDd3BnBZMOl2tES6qXIRWfuPoz8v6Ur2U
m6LaP8Y2lhoQxDU3/qHnG+UWoe/qTaocpWDxSzS/we1hLQGgVcU2lbpGrOZl2+YM
DvROCZglc4RAgqzZIDcpNC+ol1gpIBjx5+/JWmmm1Gjs+ouglqUEo9Je6CBWu3OY
vKOCt8qX9gTnlWFe1omTrsRPeet7MZN18FfKoCTCnY9Fku8yuomhtdWdpo/GyprF
tcO6dcpxFYs3MhTrg3FcKq1N3Sj4iSKgHYqHxVCHCEnY1LlOnfmWdtTRqxEp2HRS
jNrshyfG0BMwuEQ9YMDTzjWhbTkdVpQFHtD+p7H9JQFraU1vw+aYPGBEpPlMINp0
vPHCgPbC30okCFloJ7KfN6IjyGjCyB7542K27nzeY0EIkb/zh5cnevsfHYzOSzJm
bVj9rGvBSrYIrP6MaKQrxJmItUwcXYNgVhXpBiN2B28Jt2jpVr0DZ5/x0FmCXyM7
b8fDaXgcpq2T6TLzFQu1fuuY+8aQqWKNZVdHczn3VuDfTZ2gnKiAPCYpe80Gu6pP
XBxY14fFSyX7IYwBvpSt3iJySG3Up9G4JWuSrme6imB6YjzbqJUSWmZ7nlChXS9o
8tacqm/cYIlZOJL2OitzfWjZc0/vX/movflElROiboDufGLOm8PMZnr7d66sLzga
PVH96nK/TcbSz6dcWEw1B17/zWJRPWDmgthQBU47ZE/jCO2NF62w/UOcpjCNRr71
LJkTSet8dgbUKEJ7CpRvgYwXNTdwyjopXqvr+huepUzVX+J84zwZnMBTgdl0Xwid
Tg2vXquF6m5DcYom/J5D/RGtusun6jG8AxmI6GrIO+n6A+yssXoog5G7AiRVKYz4
ebVKB9iepobV+N8TS3oj2OICf7ppd+1YaA0ijr9mHLzUxTbIbVXJi0vXio458Ast
znSPKd7w0WaAaNvGuE1d8qnYcSf5eOoEe+luCyXdbigXc1pqc9P0PJzTvKv4dPY+
7DoCUVzxEUnlhy9JBGgB681TTOCSFKsMzY3zRI47aMIvXACcJR78NFKSETTsHsfO
V76bsJAlTK0adgU5ZXQq3FuVjf14WOYMC6XfG5awvAdREPLelPWWz/N4ezObzIqN
mwVGzL/5qOpNvIVo3saIFB+BcphmMcTsUGAL5qix+2GUizqHe2ytdEDO2eTSJCnN
wgFb5Pg29MUsjW0NZshkEY+yxwDbeJhm0+aqaP7/T7HQ20uka3X06GRagUAlZzr8
8Vw382jljgYuha+QqZGEQdHBFMTm0Mm79MrLNOm4WIIj3eWnfAKzpfAAeHmNAytN
3rzuL1Szm8qyPXC4FUOBez7H+h1qBtx1ymbpxIcZUh20Jbnt9TkJbkI3E+DWm4rY
XwFKP4ySXmZJS3ngJuhym3la0cki7gsmpbFmsuC/cEnWN8Eu+Cg93zj0+AQrX4i/
YPxoF52c/IhvA9gPE54kgFQWLngABOfdfyZCmQAAwhTkPGV7CG+EIu4fRk7hoCCV
pIdiVJBS8VXQPouVN1XqJpIPxiwg5Tl8b3Eh9GCBF4jSO1K3BPPLCYZlXeh8a+iS
ChfMBUGVnhkMe6dAlNkYnzseF6IHWp8UhJHHg1DCJVCkRD+kS0eCZpaZRKxTdDUR
5uzVHSxT1h3knXUsRnf709ZHIaat6j5ooSCYPtBFAzqL3Ci11icFx0BKdZxP2KY6
LlJ9lrYpyKU68vUBdmGr3thi5JtkBkQ7UDf2mBF1UkLdlUEoy0Yr1JPha9YCKlOC
nhLA8xrnv4ZF+jmcCBWI03ildG8Jh16AcF5aXTfKg6bJmR1z1lRfbMm7E0NPDwdX
aAYGamOpYd4Dk+3404ZzQOromkFfsuLPz9L5Ic50AsUDwCrWwLfgXkq8REt5jLlH
vtYlYe+M4D5tkrwxftw8kSGoXhXxe1g8O+eG6OXxNw1KaMItz32L5FrMTS1ZMvhk
E6P32TPIZKgNHAsHtssXz3Br/705cNjiddo3vYDb73YD26aRKAXsiSLDB7nnRETt
XFhcZSFJH24IyxCwwjnRXXdDaMeA810yzlYbi5bT+NVLuztO3KhJ1AVAZ6B9Jslf
Vqc79Nnk5ZK6/zgydLIwYLO4dRiVV11+zCKzmBTyBBmmBudZJTs5Fme4R+qYQuGG
MWDU0TlnlN9wsQ3AmDmWqOk9i4RED8MqjQQeL+X2EogHWuvya0P9OYnDyQUZy0Wb
BXmr6+XST64H06AMetpKaPyfkeT0YWZ7QrM/ckH7gSz9bMqLmekYkDO/Bj8EGPkm
djOMzLba4Q3kUEDCdkbjWJELI80wMjC+/DSWxVKXkHzWMii24vUc5I9qmm3/+IVi
7cd5I8PAHun7XhEGNDCq73mwDu6qYzAL/mngGFjnvAf39wTy4S+XzQXmaK4R3cgo
qLfHEo9PI+Ojf17Ki7oY4Qj4FvcAUdTXONFnXM5ZWrAuwnxOc1uIQW7BBJZdbZBR
9+FhUDsGE6hWIeK1UWBm3z2sColgKwI4e1MKTIkzmnzTehb6qaq66GsYB96RbU6G
aA5P/eKUJXP/ThfnEv0kOOdLrey4lB2pakOrtmkdjfJvfFj343ssTL9WKhlocqek
5xTX7+bqsUokD5+zMpxRfSSWUlmx1/XDSdlLWeToS6RSfvy5ozSKQILxcqS879Kp
fQwuLMDL8P2EVM2koPyo44QHhXIiHHs5du3AdgDcTDQ/RTc1NH8cnig39pJjBEOd
mfPG/5as61fLhpkhWVUYdOiarmEFqNK28XFtGb8vbFqioNC5kYYYX156JXaHUtg3
y1jaOFl+ycYTpKocU71Yj7ni9OMUttFHhqjCgazL415ovo/nYar6fZtv454TwrfV
yOeDaHIkjdVCB/aEgdfhFI6bAj0L0WzpnsAkbvIk7q1tOvYA/bT0AR8+nyrQBiny
dhprohQldX1kH99YODxqhdyoN/ZcVs63+wSSsqW+i3rRLEMY5QfM1KH8/zYSTt4f
WrsZDNgBfRPbLv0RA69w0fRUWpRoOTOoxFkSvENClxCr5GBMbTI1XW9xFwRy1lxq
DykwefQQnxq5ec+86KoEx/7AYlYIhjFJVWcD6GnBbIz3oNXdWqxV/P5MdwjhYHvs
idQb9tp2kbtzMID+iVgVIi9c76jjUUhRhlhH6UHc3Eywr/JHZxdkJchbIbtRH3yH
d5WPSxFiOGXmlbastrEhDNwHdDLFkskHxPoT3BmIHLBF7c15Q8kiX+6QeK246Fdv
TXkBndxCY/04h92BnH62fi12qUREJDxggEFWWB9czGlEBAGNNSejHbny/SpTaZ71
aMbkJUNs41oF6soB69i2eNjNbpLpIaGmNaOLXOroODMpyQc2sthghbnOEUqEdJ58
/bfVb36prKXmTB0UoY8/WI1PP/0aCyVYYlkFa3Q2c/SMmKBIG4VdtxgkzKyHiTCb
vkd4IduUoXFBURiqiaAtYzOKzigt7Y9ArhdG4EzWeSLN6HLSGyko2Dvyp/TlgGTu
V5xlFmTse5CTUKiEldubBGqIdcQOLRGggiMr7K6xhlniyjPsiBzbshmIRvOlfM4M
5w6ER7z5Ox/PzHFqjgy2wwGAdqQzcOeqcBtvOE/FQAS9pJNozLbGPU3bBJb741/1
NkddOtKTq0rKCWSaPQG3fILQHW19YLcjKjmWuWd2FC2mmK42+J7l81dUhiABe1hH
TkqtBX/jrVAIrbjE5FyY9op3SSZmmNJbWvqnmPIaEEAMbbJOWNDP7GsRFSjsqGnb
MUdb/w6GpSBeseYgeLflqIuVIJtc8dW/yaY0fkJR2k7oVIKR6a5jwZ2KuU3pFuFf
Hj6OAWJFqWZl5RbDCbNIMukapmJjvdmOiCcTWDigtmmrP6wz9J0kf6Lt2sRLYVks
Vb5kpj+tSRWeQhwG0HtO3YcvvR2wvVliXrwkbJjAjUyN8bEfX1lkZtWHYuVgYo7s
UxwDJU9v3YH6AI3jbhqYWJyoq4EtbYOdRv1KnWbXR1FtcLQ+mqmZDA6q7b8eVpq5
gTuCp/XlebSx08P+npWT4JNPaO/mRszoOoHag4lA/P+lr87iR+Vl1Huc3p0vexat
B1PxWue0WbpF8cUzegDgQj+a9F2AVKqmDWjor+Asj/km+Gxmyn8RjdA34OoeA6Aq
Bi4E6LdrTOc6Pa1Lv3mvOGGp4+eWm7zqml6SCmRhsq1mFnb2IHVyQ9t5zzWYLDKh
VLfnzUcwb9O1iGrOCwELGeEQVcTyhxkhUHeiYGA5+GZeA5UdbdFwHc6xwPt8HM0u
QABWfbjlVMC72Fhchx0ULVrYQhfxokIauXldKrzazFkhqPbx2f9lc1oq2yPS5+a/
CSCgJFH+jDBQsvmHvaiViFUWNWMTSnABRBTb4gqPP4eEMFjM3X2ujmAsx+dhSIFn
t3I05E86kcFInH5gxcXhUygEn0+hhhQzluw+nCY7QCxp19H9QIoHjGCAbfRcYlYt
s+UFRD4slWbPf7LCrm11rIQUOP48ZGYcqyrlNJE/h9RAMzsISx29WRjyFjCFrXvf
wskv58G7KIfXtG+46WJqxPGsNMrTkZLhOK+idxd9LX1R1DoYkzBWL2R29obD7COp
AzdBIpjQkpwMu/luQec2qsPMiGM3+0QbPJSSioGUiUUqz0xrJFIBKaLkGlrpamp+
d/n73ucsjr9qr7cZkMBLjh78mNM2jGRKz57etFNnUd6UHQdax0kHwSmyowbKw6ti
Uf8GRjAd/quC8szcpZ9l/ewaLm1PQLQoBfBadWb/QaADaaQkqxfH4zawf2aheZSB
CrGt5lbdVGrNXScA+AghQDLrc8X2e5g0gWEPrUfLG3ejsoixkmJlqM0NljT4ScqR
brg1e5WNnWmwJf0SWgq6u6uEKd4N9QNUBDoBJP4+0BMN2r36bu1r4DXUzu58jYZI
JHT4HTCq+NGCtTqdh2QQ/9trE6g8/JG2d0iRIEfAIvWl+q0B2J5kOjsJLe1GVa0D
MavtSWmwhf+mY3SxMbClbjrDJHUZzYBT2CjdBmXLm5Jlo81s0lFrIehkmTHryotB
LvNqNHMWFnMu6yPJGjxLx5wcoa2PLpt+boL+661r1tlRTCATj1sA+9Jn4kkVDdL2
dCB+Mq+Slw5ffprjfR2BhlijfBEMMEdKHxozmNavyrtnVOtDplBo1D2MAwvwGnwW
AhtNfS1Jh1t6MWROvd+VH3KaCIi+4dgNs/p0+8+uKxC4nIpWY5nbd1BBrrT25NU+
0Y0XXWizSUrb/MPLl9LLvi3tt7owwVOh/ZU8NW4AO2Gow4lGRzqO8QIeipIm3COK
UysmBSLlb5HRDxeVnShXMhF8D20Srblln6WSwTWW7yBLNrc+JWX7mhInfcN0EII/
gYhzLmw75RJQL4SlmqZ/LhA0+h08TNl+oLLT6bZvPAPzxDYno4mJ7SzNowKqC9+d
qtpD4hJvPv8oT3SvLrDXPT9SsMOrvidOqs5P5YVmWJ4voKxZkgCT2mlj2yFoFu55
FZjsH8nlTMg6mGkD2frKrLXjvSmi6QBQpVBxf+ev2b/XuAbugzcx8MlT7+CpxPvb
ll8VyswGC3aIzdkxKjoeYnTEPVTyrPRCnN+41CgyIlOEJF3vTzOIxTmQsGa7geI6
XUOdqDr68F6ChfjM0Z+nd7vUFQMKiAd+Z3geHpqldj4cnaPwtZVxTFO9peOY5JGO
NZWV7z+uvuBQGfKNvTdC+DkN5Pwu52XxlQQ7LxtDJKGJ3hBSG3IExHNrHGxSRj7B
nJT6qRFpsiwtQw1fgHiLl1I9UvYjaTNZ9OLIMzrAPDRQ+hcEoKEtEHXnVpqslvUt
WX+lO6AWnVkPcoqmYVWqPtzK9DasrFmp/n+WzDhF9zvekbmmFwQPv6v6lh5EO0fO
lyPcarTfA8THn82qjl6wF9ysfC288Tp8N3WFdjQJsCHFWZNA/gf234SVebjrDdjD
b30ryyYddVhS6wQJHb2PQA+p1S3ut5XU39jkcex7utz+s6DoiNsika7ASaMDTQ0M
LaGElPV9OwG0BKctSzSZak+c+508vqshDPWQ8aShE5XxrPk9rGDGjRWgJN06i1cE
7sPZIPXRfEjgvpwBNFXR4H7tuDywlliHiePsVGfMzC4cDvUwBMn3McHWTGh1i6x5
+Dk2uq3Yvn4971zS/gl7NaDMRp96bS/De4LhYiVK1hLYjxFo2EstihoCcXHP/0cQ
9/xLMIWQXUFPYo0dxrTlM0mfYv13ofLasIzlBJ/9UkwO/BGKRnIeOMQl8dmSwwDi
UgCXyiRDDLuVO2NPyrwARyAZLUmjffrjTL9oya6HRr/a2gK7UPHjKeJ0uEXdlf+m
ciRoDUAH/ScgemtZP9mjVlgeEq/GEE5Uaam8+pC+VQ4AyrvajO7+0EXML91pB7Jz
NqMJZnbbrGXKNmLNdn88RMLCcraF8FdjgBRKKRUHS9ZzIOfQO0DuTWvGEQk3eF2M
3R9YjRXs5zG3g+Uc+SubZjJAYznPdVGLDJ/w8eiaLJzV+lo5QJsB1B9ShGy1lruS
qFCsDUQm1nnyCUecQcZF0uEWNn7ffpGZOE5gaPmFcsRMX1Xofr7DaoCWvJsWJTKv
VFUhXPVECme0frWISPnWS+SW7lZT4xt8JtpyHn+tohC0zRu8UHTJn5RSjG/h+zg5
eYfpEerYOMuMbF570m4F6bA5z3PkPTfRpmKatsI6SYXTmWzD6m8rlDTcb/K9Ce02
tDLRAbK0fC3/ETXf7rpr94mNgIzbgIP4Goc79yiwLktH/h/6f8QoAYd1HV47IG6a
rm5c/ZAatNw61LHkrHg8ez+hRPbLwiH0evlWp5ZUaOnZTHkDALbQ4YossDJVQo1j
0SWm0rS45IYp44rTTrJzqSzicMRt+Ur4AYBBfAOzx3eoFf8f8G4DfyBRG1e1cInj
HNF+RnX2RmOUJn7EyjzdryzO6E+zoN0wrhqStLQtNJOEXZWm9ZLkQk3n625PHdwL
fkTG7OYDj8z8O5KlQgKVwJdppZPr9dxuTDiByftkEmmqrcl4ceGq27JuSsaY4iQY
tMH7K06dseRL8xAk6v3VupepUl2akkqVgy5BOFZ7OZqDpubgvlrZ8CMhWlZY6E/0
widgg1gtHO4wAbbOlU2Kx1kw+230YZT3o4JUQH0L0xlSD+JXF/YUVbW/FA7wPm+z
uAgOhQi3ONxnKZFlKw2LVQSYv4q5Mo5FZVfDitdOIQuYI++kjEHRASe0nAXGOXt2
QUU2/m6Y/t7is0orJdlRiI2A9anh940/MLU009PRtyZwsYDxIMhjm2aEY34Z2omR
vaUCp9kZWepopHThL4KKAuaeqJOBPc2MjL6AeE8tAnBGO1csnPnOPqzLWY9ZMzpv
5WlbmQ+SaUSBi9+1LX6N57RWRWvf3FjBtqpAF4zUsG3wF4lCIPWMSKjAFpNzi1Qe
rZQUznbyT3ThGpRNmQ+H/agsvNFPOTR93uz5X1qP/HcwuzgA+Fl5yF1PdxVk+TNf
JlPKPvtWpnck4Ugtn4Z2UiVEM2pRzBX9GAOtkB5k3kG7+WFLwHb2B4hhBjD0Ugox
kavwyp72wVK9UE7idpKXiC3Qz4cLW+GcT9D+gIO15+pAO486dgijB/4OElGy5u8V
EUM/u+FGCX5ztcl70qkIvfD21LFgTbqq/VM7ZeeWY/NYi9faQzdPQVG+DS+cFV6p
NEkbwKDjBQSBXFIjlEC5sL07fzGAFFdLAkYA3voLRWtEKcRPt+0Qm8AbO9OHR8ov
S0EgY++2Igsx6M6UvgWtWJkkBebtgOkzc93b0inDaClxQ7yUrDrzs/0YLsn6z6vB
4tduMTxFuyLYeLjF40cRA/mLk7XRnZ1gakyM11hddwXDPPOPg+hsdrvTWwKJmEBS
0lG6cxde4FlMxTPjlu3Vo/WVkJda9y4iaMJ1lZiIwD78y06vZTkfz7HxWroIPE3S
p7n+wH5O8S8l9goqw8V6x8XBx/Atdw/ENmtKklw0NB/tcg+W/6maFOuvlW9GZo/D
byc1FgUcotayIvCO5y6IHWQqKugbZ44803O2+580Q+619prItrUQW7mnh0VQrO/b
bFS4nftQJQt/zKBRFZdc3qReo4WJ10vM8MQYk0NKQPwtXqR8sfQsmPnOr55qCTt7
Rv4e7+yP/1maWDERgEnvDBKEl02CJdiOVkDjjQXCOHDsiMgISLka8hTFFOQN4vs2
4/Jsc4hfK1ElieLHZ0JmNg1x3kmD0laCFWNDnHV5bVSu3zN418H8JI6fdzJwQzGv
+XOthghuBNERpb7INesvqEuAPvIAPh4DYJtk1MneCU+1w9KWMnOu9YX8dLqARNY6
zXpuEtty3enD620rlE0e24WI3D6UNd+reiqi7hROPF/WBK/muuysEHg6whw58mzN
GJSaFFgrTTsC/9HjSTuWE1NnYo4AJ+pd0jaulVptewSsS00GlVrP8En6LvdrQsxB
2NuRIW+JIJZ7H7/if5xOSCIJbtjRUm6GSrbPrmF26r91vu566u/diX9ofdfnwnBe
y30v5rR8Vc40p81K0eDJUmtpWggm3TZ66GCLEhvoEBczgLTaUc5Wnl8dvK/FYxmw
gREvl72e5hx1e9sckr0RbY03jWrewSuIgYw7fTm1OjMGmnjJ9M3stfio84LIadUs
oAMcFuGLalQ0bzSvKfg2dLMM/WSmFh6Vqxaai4sV777dD9g27KJwNw3S3nORo5Zt
BttxyZDDYujA1+6DlIhP6DpE0mKiGdJJ6r/mbog8XXPhmFjz2bOWnn3X49MpqR3B
U4jc0WoSW0NXZi6fDW0uKho5Z2JYNlQvl7IVupLgjzqWBnO/EVsuY8GSX3J0cU0v
shsL92jTjy8OF+4XDpMU+DWqJeyHDYf4d8dLjgm/5OGeuBuHjc822PiR+sTqwt6q
6H9TSJyY+b4Bx3PyQNc5RdD+chyTemNyrvqZxbnNvZx8NJhCIQ7ixPkC0EzlqYFI
XtbJsndBTqSytOR16xcCI8kGNaUILtrBqAocDEUZvrqezlG4fy/jOGxw31PgblI2
+iNN2modSPaoET03wqx7TfXiPI+46bpyM5dTnMco8PzZfen9YJ96NMTudlrDGnEz
X/Q00Ph+dL7gjnWyv5Ku+ORsIvXnJc/50dm0f2JwJgmrwhHkcGycCSZx1HSA9dod
UjDMTwrtUfqa8a/wn4h1ECNH54mwLqOw2oB/za5v9onnAeV9zAFiW4gXt1pLEMjI
hKMz2oBG8Af5nduwzg9oPuX4CE3w7bwbHKJg387Er3dx+JdNLY2rDDCjHrjJJZYu
IUDiRZFAzY6tgMJQJ9vWQ8qpmWkEIWJn/iOd8UafKteAi8748eqE47uGM7xrtVOz
+N+Oh6rM5eBlK8Pla1TVd+Jd5xZ9aL05O49Xgs5PVaM0Y8bopGG6Hp8BtsWID/Xh
gpMGoF6+vMXhqUfGkYgWj7GtDh84x/I73pEuTvVE1MVRPRkjzMiiDXizcfa1Ll83
8YRRCL5SIFMjw1LpSOreET0vCqGfEL0cV4PuOKwmIDA6H7cKKzkKLd5XP3eYa/hd
SZ2Idt5YT/5RmYurMWUgyqYyDadJdpx1i6enuf0vTATF1B11njZprWUMajIw2nKa
C8uoY/OTX3WVUGwoUiKNk2jlMkcLqmNa/EnRzHtda2b/ogLH0Mp/NxnL0TZukw0C
1vsyuFcKMcZEx1QqfgAVSKIZZkct7836cduIirOvF1Nm0UUG1Y7fqgTvbYgxYDjv
lcbptcHpP9qWGGqQMdc/ncgriaadysAdQ7Nys4RvpmmJOpdjMmSPdA1i0wX4DYzz
WDmusQ3xZ6WsAINa52jvMB4dlU8ch6e3cI7iLb1dq4SOg/LZVBo6wHaoeshEacsP
aCJtt+eZu2imCP8xdolBSQd+tEqwOw0hBuSt/A37DSkk3ivUcZK7kSwe0O+r/L8x
zojbcan7dWYioSjdYVGGiMKs0P37WB1HPEeukRZXmdfGm9GGHx1MxmkiS6hpOuLM
Cr1wJAhm+F4pANzucILY3v2alRTzqHMOXR+nW0nNivGBVlyrR/VkB60aFvf3t0fW
a+jFWJvrWuTqR2eUzJZC9PYLuPDB5UWzpWQtPjdmFO7+e0ZB3MSYg+ProM32izYP
Qr5U7jWRqc5pjpwZR89fs+/jdRGd3BVuRw+4phTZkJjnmaNYFAHpgYXqE+lBrmsS
7lJ7wGpzrVhKoPGCduHfq5FkgfEVi9qJVTPc8+BJI7gOM8fol+lTkqj8xDL7XYKt
RqhQvyhivpeqE0bx2osVKQrrSqtkpcGjIb96ib4WKbEKvYr2lLJy/C2Jlx04ArpF
mi0s743nr8Lt19XK4JF3DWZT8BFinCmBA+5+x0i7/QKv/6LhX/2IYl+45/dhJkcK
qySpUWFUHHP39MUM1++fNPGG4sGH4IXj5eol5lQLrOIc9mAiSu9/9GC7D9hQePSP
Kdq3c5bB+kSFMcq0tyzW20rVP1qP1sqvL36xeOS5RkuN9vg4uc83g8z27l05lyND
5lzXkYLQYTIMUmGvZ2YxwajLULmmiTWz6m3UPYS5E8be0oTe/aOR4FBjUPG94Dvm
JpjquvWjbf4odpZghLVzHCEXWj8bszVTiRJ/Z+cdzESWzMDTgevx88WV2/vMsHoj
5bIKp0PfPo8wMF/3bcOCNtRJ3KJY/K2rBnb7s4u+nXtRrdsCYUq2o7vh4y2jSXbt
TrkR32uZw+22dkAKTiZueFePfLrni9t7V+RKolybbSvnhl/lhFO3zZ5m0joZpm4x
OBwYqwnPBD833DC7QqrCMp5FwTgr4XCS0bZlR63jH/uldyW9lWnh/yN0ft59ejLs
PHckRl25UG4yqd/r/wMbou1kH/tuPvkJgRZuLqg0tPbuUZMqJZo8UwJvbwjt1U5F
cvBpSVJkXDOsiTU7/wWAYd70v5NoCfotrUDwu4HZ/q0CkcTrinvwSTDkBNclsWuV
p2ieDxhXOykBfISfaF/hmK4NQCkFTW/DhORs0srXb4j4DIdNyZEijebOd1PykOCN
orl8Y0S15Ix6KzUw/kz1cfME9IWg7M1DgsHaoGOm449MpCMr/Vn/3YbgO9GmnTF8
O2Yvffag5pqc8nePU6GZVb8IUQSmCjXG7vmiyloVlMKROdKzTdWeYgrMH8ioBWBr
0yL+j+IR8Gz/ByCs+FSdP2BOb1hvmABg5QAlXXlmKieCfR6otV15WAjWxgxkHjn+
bMiXPFE7yo34fSMjBwBGUTs6ejyTBbDTjg9WMXB5HXzj1jWTi3gpJ5mkuePUcRcJ
zlzcFDJsscBwb7udZM9vt02MNA9UC+wbsAHek6Fb1q7vL+tf06Ka8ktOZQjHuqnZ
1J/Q8K7slyh+CF0EG/PuckN8bPYnKV2z5JK5DUVgWrYYEES6yjbya0kcnY4sKVlq
9xwu4RzWdyStlzDIX1tt4QU4CCyEORLtnWd/6IG9eEQ+LuBnnuLxjlnyUM7P/08O
OR7avd8FjDsjpQwn4FYCGG0W6kFDj5LzLlhkQZ8HuESnPsiwMlKndv50zUbcJtNl
5RnDG9KmtZndplVNlKjVlrG5BOBmokoKqBP459qhBH/o7CrfsvxcemucpwCvrc7h
EixJYjZegbfhuR49yD++Kp2mclRChHQjRLr9QKkDK6y1zzVePlbsQTQsMDweL+H1
x5zI9cXDByqubIG9/6gMdZyPqvLVamY7s5ZM1T2X9EvhjzDLx/0iJev8koRwgLTn
OPBP5d95KW8aIqxduOgPgtURqOet9dkr8LDIRmIAsUHeqStUErLSPW87krfjj+mY
IxwW6SjjqEy2LApJS5Na7tkPDT0xl+fdjMU6BEt3ixFQ7BKWQrBiyL45w09Ap/tV
dQeDblEPlrO/IfAuNRuChHDKn2yvexLNFtOIHlgz/RFB5yZPVH5m2jtKjbRKKa9L
lRrTHIFbGwowMIOFa9hDmEiaMTsgMee+sHZ7t/O5Xy4Wclqj7ogVRIx5fECQE57c
VjG1U33fkfRZiNEfGpUqOh+u+W4fFi9hoJ84lftZwBUrYG4tIeb5htSwYR2YFCRP
0Brd/+IOJ5udtks9z0ZIaa2/txVtxBLGYKpX9cj+oOE6IGQHcj+2duxxp8V7GmRh
DoLFf+6KPBISvogJ6OHfF8FHhla68i87nYOL19uCAHhRbDkhB8rdOWvG6aDDazRT
9QLskZULH9A0fyFYfp0TYRG0aeb56K+PInS0rV452ZZLzjmBqaIsFbNUl/3XF2DQ
NaON1hVxDTG/7+0P5ZRNMgMePQqasrKWbm6LabmMjLL2B06D5kBrrayJEVUjNzcd
FLqSd1dN8I9iDEaZMV9XkCyiUsdeQR3uckuyALs0KNQq1vaMUVmBso0J8IR7MKug
xQX+b1S74zYKprUQpxvA4WF47+En5/sopdUzHO0H4LhJ7AyywyTH5tPagjm83hVD
uh6VxX1EycB6zHnVpQAKIxVmsPSyTOjvR1KOZIXOvmt0ewOLE703F3iQKUXDLyv8
7Qk8o5EHeUBaRobPivBRzpmY3MiqrF+m57/dFmkbwiLI6F/LYAN6Hq9xSZ456x53
BQ8XGB/35kTBPQFabKqNi96sG6Hv6+7Mz4nhGEbEeKSRsxydiDpZDr3HnEJgFNyo
ZdiMe/9T5mTn9IHA6x9c9g18YbsT/hBEGMOOcEFPlqneS85xIBHW7KZ6r36VrNad
GCfgpXL+tc+nKk2dZdxISIWbHwQ4zrv+rmop7biEVCOaiVHTCwJenE1j+ugYxr9M
pqFhYlIbvbl7QEHJ0Pz0sZVlK57iLnvSEkZTwOolkLykv5UOJgjmX5lPTw8vXwqJ
710l74vsLBf8YQKLjLbPiHqk/5eAGjs919sMVtMJfT8eNZgTqrKs3V6clSIOv8P1
/8apVNFkCXJyrk5JPcklJ90K2LzKbtE3EGEt3HjPp8AMYThYvRtIqrOgIzZxjlrp
MW8IuFfGmUWeu4KKnjBfV2X4r7YMZcSP5Y6bdkUORge+r+jw4w6Lj0XRVPHC4tin
55jrcEypSD7ku6GVRm5HzWrT7iaarCLLUk5KIa1SItnP0yMLuKE9wyN0oRVHSL30
pczb+Audc5bgTxRh9a89vix9CIfDlC9WBTGSxxq+WW4TGi6fPtPyRyC+0uIdM7bv
nB+P5+zrk0GdzgjeloKHQSUsr25GWBKUHYw2eq5q3L2faotqEU89JAjrsLKEDj3W
2nlRUi1vxKNB0aoiiJnArEkGoMd2y0iMRR5ObwKGiCMQMLiCG65Tv71zwE0/0jPH
a1FexIT4VFP9zudTuWoazbnbyrKfeE/9f63/0eYECbCGAeHqV+SG4Hv62CvnARZW
XD0elaLutdhHiUPPlwmms+eBsEXDco6pvO1rNamlaJUWcHUvE5M7tkJNUZvqMn6F
YGat5yzBBSMtZ7bITvenUdgWLCTLMbCL/ldt1J9c0IZB63p8ltQnp6vwZ6LwnR0z
yCE8AdQ6q/P5+9iJLfcw4T5s8UisTPirDwHakgjD2p3Yzq93IXpySUFsnmH23byx
YFwb/QFX4s9NLCZubt/ytSWoBbu05VtQMSSP1stLaGg9ZhCgz2/fnf7MCwCLJI8O
KK5zx3JZd0KMvsSdRsqp/mJpvPXiJhfzRDgmesxS5UAAcQ3X1S2gQNlTc8nnLP90
AdT1P56T1bG4cWhHX5ZsfKzEx9Xzxarm95GAYGThHXL6pvIxBwC49CueVgO8koNG
M3kWaFC0+8D1TzIJrn7N1C6cqTDNYiL4Q3KCflhT6ES8qCmrhplQ46RElkX7BjOp
OJw5tlcNfbc2a9R2o5syJaS066U+ZPE3diqf++3s7v8TMtx+foZrMbwA0nKCZiXt
RBkP+u5flWPDJa6t7gBE6ooFnWx0ebN/F1gTtCxujZmRb5rZ4Qbtn36zSzXdHuMe
8fInSuuMJWWG8M85TXWgHtU1cigTbmPCR7AFbAOrBQjppr3fBbXnbJ2hFX9Bi8YH
u2qn7h+sB+/zC28A7VfNTnuIUUMASMUcMxcNQSke206xRslWavPECfpNUgXWqj3W
xfbIcBdX50tqpHb0fLPWdlezruQs1JM40I8p3aHd/gFRgtcfm7/KLie27qcCS0Q/
p/hoQNX3QLRP97/cRHKaMWxobaEuTXYpIltFhhdEhtYNntjW3eiROG10GqTsqQTm
VOtwDSoeiMR/NyOMh19sp/rUaA2hBUAWNLq4R0LQVHcSsdr8broMfxyDYPLZ9I07
R9rE66wlrLCwT4/Nkmo4E/Cgp6afQyi40co0E08C0o3uzQWs7cMF86MlZzQDkd1n
agI1b70JwfG1Q8j3X98nDR0fB37q1DHxQsGEs8PhZ6JNaS77z6YvrbzImruqIVl5
vDw9B/pNy+x+926qXFvW4ZyNKkqOJaT3iDLfSCtJmJYuVL0ezobMXepUjIlGK9ie
rS7PBhohb8a3r25TL4VWtZeBzSU55SZToyUtFuu7L4oDlvdtiH2tRtGsGNfgYJ2t
nnb0NOaOitGV1TQxFjceV4aw8eaXOq16PNmHZMrzMcjPH6Ob1o8ekDgfFzLcDuMI
W7VWEoVOeiKfouqXB4PEhiNvaTbtiMtpdFl7QFLsXarAdax2fA10/VYf+dhoyDdj
lXW+QM9oc9Z8ZoyhKkDJyrlu5mtQEXb6R1K8S7MAn4LRKBizt5m02MlJon8DpR+w
MR1YJ+caNQDrFgdTY5mbKgXv6aj9rZilhXkSasNIQq7cjq4cJ1g24O3VBBgphvbM
YBJbkYydzF4VWhfxc19qE+MFmrIcjsAp9caG9a8qsn5qFhIjJQBuNoxaZQbsZXB5
V2HCbhvsB/AO85PhmDXBBRUU/8bbsA6xvNX4b8acyW14juqq9c1fmGjVefQx/hLE
P66tV+sUZNfMoZo0keXF6VaUwS1A/pKWCHlymRbT8nb3XafM+LTxZ8nMcqYYOUe9
VhQsUTsNCaAq5p9YEci57QC/A+ls79s0JAv7Jje+MojF5uKfDrUTtdVtgV67XNfy
tOj9P9eTDThCrDJ2fJvRpoDi9HnrztMsWB1LnuYm/WnKx6W+eNV7L4Gi8f1moIRB
bZfe1Ery7lYXk8uTEo7q2sP/X4BSmojJpglceEM/UlSrV1+aHO8hCSjss+GvABGM
/hJ8Ti0qDdOH/F4dgKG+D5yrT6MU/5e89+v1lYGh9RzOoiDCsQpN0I9rFlXlZNJ1
hlyYMilkV4oyT9d6pYcnei8JQ6ive5vuHFlX8WAdzUYMzUD+QfEODBK50c8SQHr4
r965wt4xGvBeapYkR6bKmKoMdtcadHYCQrkpbs4kcNCVQYWYXXU50bF5LZIxzgmz
iuRI5IQlssze0Pe92HHfaRJxSy/HhrD0/82sl1xUF/Xa72CNqKa81WjUiIKMpNgU
1hsUcPQyC0lwJNke+dmAQ/t3a6mWZxuS1IkvujxQAOvcFkk33zIjM53Kr6YDomwy
emO+d0HaqsYN++EPDeGo6Y2QmuUBddLjQN6Sacn6ar7Sy9Z9POTairdgpECJNTVI
glWpKalTMOFgU5yqQj4u8wwsiwNimP2UjsdJ7kbRhsiLJZQsGvw0YiaR6mKKHmuQ
jiYstFW2y+ytg0IM7t6S2VSUtx73ayT1lOfDcn5mNljPnl1JL6XQLs1UisynBRRK
aTQq1288dFUwwn1mZCmZ5ySK2u1zgrcI8PvqONmWQRXjB1nFBpOkSdMf0QaRzBBl
qhDV4jXOAg++SDFDFUfEGVGjvgw5K0QBIB3hqaBVVAt18riJlc7/PnVX0MDMinp2
+aN04y1djypYy3kunI5koar/3T6fLA7cVJokVeyo/DbZXWCMTOeFrMP71UJbcApV
lzHvPnthmhZteIAE8ohS5aVU6/SQX3POm1Yaenp+QCv3WH9uRvrlgSd7lI6ElMpw
pLsVAfK92f0GwFjEbwFAThhUoJoJmlL3AImjpbCI+QZ3o7wxko7ClidI2v1gEuLz
v+XDwIc4eFq5GcRNF0qgqW7XzYA9EghvmqqLkvJ5+08AhPV599N/5k/oBeymi9ii
hftJFNrKuixr4roR8PhFk1FCGMrgOmYOA53x3hfw9MCt72ERZgFzU0APXtYhlcNr
6hbajF/DXFu4ePzlF+cHsPrjErBjzykxbS9VHtVX9Q5ijR+Gpk9unmriddlvXzoT
Q/84fAlaFSrt9RbSQ8dzIDULDF/79qf47seE+5s7AwxYajPn13k/rvVSEo7YnrWQ
riFawZ6SlVEAB+8zDx14XsoIznQ5E2s8YrGdL1PzliLXygWXD9Cq1oiLH8pR/BWE
mebtjbi3gOC5ZVeBzkpKoZ7FCMum95hr3CweHF1Ln4nRz90t958knQNeJ+PK6s8x
wZM4igRLxbaEq6ctDqhTouJp33vZ5PYVvT4/Ai6bBYLdNCzXUwDcTWqO/rD4g6nO
vwPwk0jx90F05og5NflXGq6AgBdyw1Rbuh2iRZKMAc9spCLL/kOfkferLBlS7ytp
M/WQ7679yq5OKR5zZmeY86oa468l7a6ASZOowprTRcrtTykHAYjBcdKW+WrjslV/
8RG9wDsputqI13NSpGzUZ3kQPAg5J2dHAsFI1amYbKfKZX0VdoZSZ73i/qA/sb2R
dOEh8pijBbPKd85MIYstSM1f3MvsiEXoSgJyiKEQf4UWroZ6vuBM3cPJ1X8eEP4D
7GJVM906CUyqLD6kUSAcsmkU8IMuPAmSWhg6bIydG+m+lQZeRBpedl6vFExwnPcR
lGVGZQyezTihmmP1g3OCy/5SkbEMEb94LB5H9JfydCSDkVPstUwpqIlJiO+Bewnd
oxspol6eiL8CfSG9iIoQaIcYZfKxyM8Cf8KHszdOgRTGErjgAFYIfigf9vc5fE0g
YgxSPP6sU/HqZmfLiUQ4gU4SeZweC2HAQJdgW4o4CDmN7FGjVpL/3xTw0Gv8Ie50
YckvRnK3Dszwa764BdQ3bQduxSdbU7zFj8wXp/aDqMa6zo3MauzcWCEVXAYBKqMm
W1/RRVr4Pp24+3vy8Vio8h3Xq7V7QLR0o9mhwd1Ze1Zfkmx71c8/0yMdRZ57VDN/
+GvrNEho0CvjJXG5uZLTPAZjo94jq/tWil/BQ/VNOTG4ZcO17kPpx97j4mKb8Pn2
5M4RL1mTBcI9TrxVD/QwmbBZUGASFLaHmlO+pmjQUde+Y+s4QuTVX8/Q1FOwkEU6
giZGZj5MRNnGzQud2e5Pw8ECEjkyI68tX2VKlB+gEqUf8+biMA5KC1iLvG1quS4j
TDPSn9u/nzYT8F3HP65ULBfsZTDCT5mjzay64M8pBzU5tA4UTRihsxZxzcHnsrFb
B4aG+KU6J/jH2sQNs86j0TVUnLkD1QQhBJnThWI8S5llPGtra7a/S26Xu1s+P/t5
ObCsEWAoNYRZiSbYti9Zi9308mmN25ozBb7g+PAn5zZ+aiXX/QtWcAvnTWMtzYNH
W6VtpY4uFwIzgvlQrIlsTRlqZ/jvX6W2Xz2vF39zV3jPya9nJSe/3UvMX8GvF1Wg
hZgUUMtvZSLygacmiybxNmR889SnTh2QQiSuCcgObyzQBovaHEH4+/YcdzZBDJCd
7IDbvSR8LOWrSp6e8U9JttwdRZyz4W5MB7ab1QAtCUM4ebsG+UtdZa5TaNvAubfF
o7fn180gT9/jqrRuZ63lpHJ3ibtqYCQYK/cN3SishsrECSPV89BkIo34DRtMbTze
oJdNpR9JDNBbnSrnmru2xcwHizqLcW8zXEem/KCw2EgQj27cqXMpjiKctbaAv/WB
86uxdL1+zutC85uWa0DQxhaxny6UDzQOZxDzmNeN6sOmQEoPzzd2C1huLTRSU5CM
jz2QAbH+XIprMph3wztYERYTqJ/yUE5z/3WbCx+10h6XR6hSmtxhFVvQza+0QuaV
GLIJrzsNHb01LsO8efh/eq/oYjxJac2i8Np4P6k/AbJ9zQ9NhvkpcZhA9xT/+oK1
mLbOFlHw/5Iv9TyZ6w5HANrGS5reSMbyS/0MBwbDp1uvkL9buDXqFnkNT4p6HqyL
Si9fNvdyozvlk/h1KxEQBWw17tmhKCOZsXquNXifMWIa7E5yIblWxdSWXVjuAFPx
jyG+bb0Ug+UN7kTX1MCHMBMeBfIRddpFoQv0G+VntS+7AnGQftfAe0rsa1MfPmMj
0vQARB1UeWnu2k60FY5tH+tLGe+SA3ZOHpyOuLEuiC2URKUVgqQGlICdOvruK1u3
hM7UT4P6yfPh5ODUq6uKP+s5G1JwLcEch+I+Viw2AjmBtkI742nLb5bcwLHAwum4
1VcWrI5AiktZEk6xVAsfaku77qRerCVSZSmJMFryMvpdHOBy+gQZSzfZoMAu6E5h
QIgbapxq4HfFjgnDO8s6yhH01ZV5Eka/HgE6EOSEdee2JP6uwePelqOznBZjCoLR
JN73AmwZ9AEw9LK/Xr+gVQ+mDgKHMQl8UoZuvRFKIgfemvPdSsAsB9cXyeLqPACU
Dbfkyysk/tLz+bBrHk+rB+/TdKAVeySIQBx99J97eu/Zw5xV6Y3IvsfrLdDBhqFq
mZJc/EwMDUryuZb2jDnTBGcUhHpgg+JJia2QqITUKeDq2J5Lit2Uq2+ux0+UjUUJ
I4Q0JMKkY88OIzFxYjvj1WkBqqoco35fpBZ0Cc9zPSV0eDHkKLH+/iKZSa5GCQhT
VsGEAdr8fw+dYY9qI/9yN5OqB8BaWN1kN/kpTBgi0/dlLDrsez2gOHwcJackJ4RR
/FMwwrz0abtgtWXhtvUjUWdkwMHwZcWq3CzFprR/KjP98Zl8kAgo7hx7swJ0c9Vv
FIN1OAhl2Cc4XFZe3zjpfpR9uw/gCBBWZmSFudbsEFFbl9aSWLfjq571WWZvTZR9
qoLwlNdhMgDdqUfC0rWzef9dEv8DaPMeE9PDil5mmv2NX1YzV7wfkIiUAXu9PKkH
FDVb6rCuQH/O20Og2VGFa4RPl9tHg3B9L1XWnLFWP52pSwiOpC0/b8R7OVcOdBp2
wyXk8BtcAWNvyZ+wKRAk7VHEAaQtQu2mOyuJJEyv+qQ2Tnk/CVOdhbFDQc8njZ3Z
pqQmGw31zLzki9NC2J+ramSXplBTLJBU8cGaEfMcjIxepH2NiJNZfQsBBXSSBgTi
u24+NSpAfXXUSNsupb+uVICM15ibZg67iGzIAILu/lGSuiorQMHkEkjifpArSS+w
vjjIjkWQT3AUNrRBcFF8SOfEQhbhHRQEtfIx8NsZP2TnsIIXCYiDG+vx6Ag+YA0V
0BHZ3TQXSNj4tYpRJ40kvGHPLBhDM6z+U5KtmOBWlRAHpR9+f1lx3qQHaEUp07r4
5c9q9PeyV1vrkRNIT98Hpe6RDjmEOQCOZy395qpfhnvuOJUuqXwkHS1mLJOYbgVW
9+caI0ngG7Z8skFP9EQL5GAfXV4gdbXFD+WsNjANb6FQjxwetvEwgGjyYinGfzAi
58o7MwNzJb9gBJlFszJfWstO1srnKJbe2E/URWi0qf2l1ORe/kJ94nab0pIKJgpa
d43hlIyZanP5jwS28bZsHQk41JWFepbFNn6EnGTAsys4QHeRMuPSMswzS4RZT2Jb
LwtyPpcW4Mm3Vn1stPIxMSJwwkrCET6wKaS5NMGLETdGb1lAS3ig3eR9rFpk18Ik
Q5IfLzyCHU3GtU4/VPwNdmqTDj4AOwpq65lMCReS4VsNClruA8sj+IxyTrMxecwf
zgROVenuEWE6tl59wH+V1wx/usl5v+Q0383ZVctO6c/HgjU3okeaou15BFXY9gak
xzGdScFX8vqx1WxUu40NUwo6qSczjUrjCMacQMsLYWTIELS3DTsFw+A5yg2SAdlj
WNGzoqjuzgq9EDBOacZturgbCP/9WRlO6fyGnLJiV0HMQfxfhZOjc9gwW6Tjj8yV
v4byyxDqOacTAHGhLYdsKIPOsytR97uXaRKGEmFjXqXBXhb/1E0I04dBDeVIvSFn
s+SBs7uVbtqJ8HiBO0yIha+iHV/y1d+EWQMFginWUquaCdxWHnqJwnYBtBbxCZdz
DB6/fQGr/PS+XNsIkyYGQ1ZmXk/Vmh8IP6T5eKdiToaS81cn5zaVEM1+b3k2o5qw
zbbuvMiCvAM/gg6NbLXXKFmutU2o6se9lVchlIvMWu0rq20hgix5iXnHRw59R7k9
dr8Nxq/jFgpfg4mLIwmVhbDPelrh2V+p255Y5hUWTpyvkpzm4REQoWZaxWiL86xF
fx2pwEn1W5qB5OPXBNCveKPWZlzQm155slChbiD8mSQJK7pA0My7i6dGgn4rFCZf
BBXcWZMyW//do2ACOJlQP/PN31M+pfZuDjF8DOYP2Iqho2YQfuNFapxBia+r0aX6
+LMyyUy89cYoVg54CScUkx+JA9+ocEcJuTue4nsh+hyW31c2NAqRlJe5FGjwB1Bo
hUSRCqZ3HMzMcUEPwt7vva7HQf4o7pr9M+tn3cXlCZEfXvIN8SGHW/+R5VwF+fP9
u5THdafygR7R9CBTGRhwZreR4EL50HF4iLxCLrHdnk+rLfBiy3RExv1O63AU+tWG
JA0MlHLL+xPPEMTnouTOx+21Xb3bl/uvBGataY4ZPnKoExGgjl8W4NRs+Rzq2T53
BGu6PLj7RR2iyr+5lm3qy0CjCZY1/kjoKftr1z4YbqM+kP96cPkzRzWmP1MbPkdU
SQdn5O7q5ibGU3HhHqrygbijvPxDdA85T8cjqo9PEtjh4SJJr3HB6Vsx3Eld/qYp
B0aGfKwoT5v/5UzYBFSvgYBgMgkcKuAQZwZv+/7Q8I/UQZbrmx6WFKt4oyBuHw9Y
n1D3aOjd6WoWwjEvhn6PZq7sn6M/MRo/lQfj5HHtnLkLrtxl9L2IDhSApwTZCMXf
jrzp1VI+giRyExfSvgPa+Y5hB+BKCZlTbvP0ZlBDIulENun8IxVv9VIvOQNlnNUb
sQNKtikmeYTeuz/sKxR4oLF9r+gKc6n5AKhuwlC0vbOdGwxbBmylhmhHxTfZU/Fn
XWPnkbBf9ZldW3Zx5jPvUA2UKc+UBa1nP6LwkTAp6Gmq7Wa3dv5N01krNH6sfnpE
57BNGS/gnb/Dway7PGRWeHsTLFWIFaG1dCDgFsLkQWv1s7WDvC3Kiu5vdK7A2ERt
+iG8SciQjW3YZvL+7AubOf2bu2nGDZ2+xupx0VkuGwafvYXmt7fo3eWrCuIAdryy
qMWS8nOEmtUPJmIg48gADCHxq14uCpv6VmF9Jh+zcGzP2Qd8Bse8JXNCNLSoxwJT
vsQG5uEJ190L6dD+8wBCNgCl6oFisXpf0Jx8OiDNBVimQzGOVNO0T9lFNj31WuMq
qfMMK/Mp8rTn2q31ipP/7Hk1l9tMThqjgizuSvgkMTYwki/XEoTj2VT0NvAN1bQh
v8PafQIcwKf+u2SJ4cO8Ktr1n+JMfK+MBRm2XVsbWGwwbvRALQrmR9v0wUvcpfHo
n7MDNQ7/Z9uLkttlvuR+kHgz+S6SBCGrfGyTVJ1ygm8KSnullXgpUwYeLaphiR/G
mP1YkS4HxMeYxWL4aBz2WhJMmwcTpmCaq1Rz6ha8Hrv5ng963qiNzQJsFeAZTK/y
Egc23E3eb0azbt2ONv9ngqcQeV63L+8+4N+evEqZ/UlsvP1H1/yaz/WZHUfqml6C
UL4IScXwDXBn+EOtAROovXTtm0HuGlOS1aVEXtIHgqZ/7///WqYjSL2gP8Y4s1UK
8N4J6Mc0rIMUNsqQo2AriMBfBTFiD01yfgjkmVygomgvUTwmkIDA4Sro7RGUYG0t
NfyIQcHWtta/nM7ObLVXjAXTLkMB2A8r8bRB6VvTNETkqy01yjvs3gtIVgxeAFxt
ugzWwEC+gMfJpoWcJxWpxgSkK7wloNcQstRBpWjdZn6pwNphpx+T++xxzQMARbBI
+jZQ7qYF2YvuGvH/R+QYC741aY+HCaH5IcbXzk7NL9PV4zZrc20+ZFqAkZdJypHd
PuX+HgvQBJ1anxvmArxMKwZQ1624pUSzvEthpn7ZKBksmn4PTyJFgYvCfRLz+yzZ
cY5UnjDjLL02rrmQ3jswi+2Lno6MIDbIwLKyWoUpsmcryiOv+y8eWEQoJEo49RrY
2cQoHcZ80CxK9uwHKVvvz+ggQjjY0TcTw+c7il/Ty2UxA2Z/AyX2muryEcz+e3yv
Oi+iRusxP8E2oYzWIKf4qBDsKl82lTJ3/r2Ddi4n37dUAFE12K3R/GcnQ3NlpoUd
2CdsGRqmGzq2BCud9RiLFBZ4Frum7GObB7NOqR25RA5CVo5Ym7vIpNVbM4ahT42S
hkRRg3j1PpU0mz5wg/KTWg/u0PxvCWseyYKt3gIjtloUjR3i76kHOTUmdW4zNUjo
AsqTEWY5ItlaZ/Mo4FIneOwI37LyXXgXEC94ch1iT/3JIQQwZzDXeJ+jokwjYHNC
LAywWjUkVxoXg2N8PPQA5wgmLY5g0ZqWElKgOFBzc2kBkFq6828/KH9hm3HnhqSa
M2czFYG9uZPOlSazgEIrf6o08oe2+dX3sPcKlQUO8gj+OAji7aCvl9xZa9bTQz3s
t8Vogy/bZvcI1tP6MAcWfA1qx6v2A0nSF7XMlIhq84qRTpVw7N8yHH7+v4q0hQxv
e6dtQyWEDRt7k2j+vhKqS7jTcaT8X8Ny1ueTzzELv5fZ5h4GxccAnbF81+T9c7Tx
H8gWs0cXzgedZkK4hoKDUW4g+QxgYg6fbOnq8e+eh5euUEKYd32/0Qtg30khIvv3
xWlj0da2avLH7TAyCi3A0aGgKYLdMbdWHtFx9rUzl4J+85GDD75oUZFrrkka7OCE
sffjgw1nJZVpBOqljOVwsT6F1QUrUlvzPrl+JR8Gzi1pvj+W9VEdKCSZ0Xadd4ZI
QhdQdzJDwJjnWOmP28LVPp1HwqRQCDcP9+WvAOhsJtT0k7uL4XFM9sn7LDY60hrM
OYEcf16HyNFJcnh4JEdgDvzG66ztGQAnfocfDyEpHMb6jxBxM+jaIu/tzlJV4Dcv
RAqERFj3QSGYkYj2aGcbLFWCStkUDe3eR3w2vL6taOtyJWHGZ5MdMxzpjVwGgnYZ
3otv4lC6WmF36uNWmswJZ9mLi7u/nJRrz7hBn/FbS9TRwAaqu4eFsu8CHUWgpoKa
+yvoOFKIWhjF+DXVTt+mf78HoQ0HFyeR7z9QasuEGtJ3N/KtsDRxa8RhqygxvVoH
BvqqBYEP63Oyl8KTMZ4FFlwqgeZ2h2hAj3K4nunqE5tqGpBaAdVYDoweC1eBzTzV
lDdpGT97vnf+cFgVRSigrIiwN6Vs0FUa0UQTlbY3GsExpTf50/z9ChhRsGiG6Lgm
DRCHBuVGzKVtsssIaBDGVMOmy1qz8puEdZOuzlWeDajnpdT/p1uN8q0tTA3nSaAt
dmY3MX+C9nzMtPZEl7o9pJyzp+HTFmsslMoxszPpn8F6jKejNP1lMRDSjkA1x2vE
BZZmRBVkxVUgJAYFfqf27cxy3JukcExIMGNv4ODTcYAGjyncdqgFykVSTz58Zg5S
UdjS4oqlanG1VumFbjmfCIj0BxIfZcJuEkBKaFmGMWue/viwt+0QNCVS/SBfevKK
4sFzr5x2QkF0ufovqpdfh7tSEr5764sV8EPNSytDWvXIA6qYfkTATFgFgnbDrrDC
Kms/4FAN2dtpOo89xw1xz06z4CchcmTM2V6oZGeDC+6v/RitQd8TUSa1L3g0/kpP
SIybJnOZEfBLRDICUI1FFA77jOj7sl2cR0M0ss7F0C0gyQapmi8a/ob8s2yk/el8
OsTEAIEufkRTjRhD6dpJp2W9T/TYBs3qCEbZVh6ZTzEEBlj4Rt3NHNk4RvjL/nZ9
XP/zEGBlKeSS+79diXZ1jL27GjPT60wX5g5WQzywpaSd0UadwJjfnDYADIMDCppG
rDV3gol2aYh4OCtW/fV9SLg48ISUxY/ZsJPwnXcs9pXgDW1sme2NDWetcS0QlLsT
cFxbNhuY/Ojy07gPLJ4evty6ehMhTxWZ2/uXqBWNFja1LIKbdSCWIdhHOmgNj2yf
KBA2yfHjXgs6k2LGIOxY9lxL8Jn6RzEQUEZXm6DLkE4W0dKFX3tzfk7ed/ffVWoL
3ua0Bq7PDDbcv68OIOVIMEYjcgFGfDpGWWEsgE08IsDiA2qMSwMabKQxb1RSlamW
iZNNdHtoK2HHTRwOrvz0Y2IHv2oqPyqGoNj6VExOLO8+8SRbSHqzrZJK40kDKLvI
6RnhtaavajI3nk3UJPpkjhMMg3TedJzoCSR6lVDZfH+JkvnLiQ9lVsPQCkhVzOdt
StKtrEf5Q+vKXOTgKDVntZhMpeK5v+RJVaNFbVTr6HpZ1ivsp54vZclaZXwkaq1g
xofjRgiZyvrAmY0RkO3xivxvr5sR9QC7XIaJD3RbwZLBwzPXrGyh1zfGUiyfGHmT
I7k57LKEImu1I3uUKUQDXRyWQdE4y+Ay95VsSVWZ8N35n2LOx1c7e7gBvR/oTFOv
QHbCmJIwUYXOIx+OixdOxyO4X+5b7GLUGdBkqYhP78bCEln+G+cZrbbvjcG56K57
rV/odkdvwjERyi+DKdzB624JJubOHoN3whvMNQ5ZqybWt+ZAbeVfzJe8W8tQDU0G
7guV5rfrHWc7lBzwFmf0eqyrNU0NAlfLnFLHjV0/MgGrVg5KZ+ZOfqR05GMXA6cB
al7avSobyGTEFRjYJjz6tqG0FD0/srG96lCJr2kfTyXFtc8sxK2dk9v+NEY/4aJr
81C1QAzt9aEtUF3UFQ04u4ufg4gQxyhuCvw1rsq9FUlaJRztjMLKfzhFM1l0UHnc
Xy4qJtCF2rPkpQTyEfh0j3Rw7oq+m/kY/25tXVVeI4uCETqVdMId2ltu0UdfS3BB
dLHe7A3S3o4Sif/LQylbEPTs38Nndfg+zvJPSJNxPvFYNXoqSdFt/3JQjn+eM9Id
ey4JvA4WAWBZ9GSVeZmUMvMDhlmqRKuNRg1rLGBFx2HmY36CxjGizB+lNrEtqbVs
FTFqELZm5P+Gn2JP0tJRXoIdvdRiGrU4NLpl7aDeB6vVWKjiePELqGSBLOWDjDjl
BmlQnJpoPOrVlvdb95/2OguY+sK6bcZzN7i90oRpjeB9FlTNkxoSfvdY6rtFXA3g
8l5Qkw9BT5eKCHfAWZTJMxC4o+4Cf6i2bfUZrqusEjQZDwVPNcDQQL3JEsa3CY4g
B6x9fLmvJtFSUMe+a8BBWdpkz+77SQ3zSvSQmnoh8qZhwoIAGNCs/RIuU0K3th1u
aFivrInxIx7WxbuJQPfZ9pCbm9uGXoRrojQdqJfWOulJS0+VFlyfF2Zs1k/Hmpgo
ezoJhCqRWNetR467Sy/V/c8b8RcZHw+uJ7yD/AssXKJLjc8sQCT/jSI5CL2lJNL8
X1uKeSDnB/Bjs/ZVfdNhny9RDhbuYlqblQhNImA2lU5A2E8/nGhNkJTuwKDzxq8x
h85+HkqD15avNUodI9q/vrszlFJktFhwtjLeE57noA7Wck+K5GM/aQZDDj84067o
y0NrkjGIKzZLuxFLwbfPCO9fNXNj4WNijHoYiIsubRjqggpzEm6B7+aCnefhWFhR
BTPjlXlc3TyE4PSXUBQkWwas3RbQvWNlYBiY+yqlafkiAoca6IZGZDq9ajWKr0aj
NgLYq92pWFlUJRNrIjGQaeqocgUwVexT9ThcGWUe2FBOEsGc0ImXLm5cYPJJqJSN
7TfQp7+hz3lO9lh/mqlBnU1taDbU2w9fxt82A+eDYAIAD62N0+oAuFWOUvBAcTW3
e+QgXEdzpCx1sNOtP8OscRIz/WIt6XPpWp5km4XVMZsy6xyNXxd51W6bgttglUN2
KClFcsRc///X+5k+rWIb6XTqmYPR1axGxcZ/0t5tWkh+F2x0ODmnqBPWkO4JGLcn
dT0lyTTa7B2+mi2a0QnfhfaactcER4c8tW4Cj5IJ6hZjXMWa881jZBH69yRYL9am
BqnPMb0E5W9bkzqNJuu+7A2QcQD9Fcx9339vyqJMl5KHK6GxyNSFNQDV33KENgQZ
B4XglPRzuJUuJsrym/fUwOGdxUtgtBF04mWHWhTwRYxxRFL0teLwZ8/jq50kDEGQ
NlY+Nn1S5fawNtZin0ngHNDYBbQOX3o7K7Oi9ND4P2hZRLvYtcVVMhItYhFs42hT
3rvR72gJEPr0sfgWXB4uFQk2sD+wYI+TN3JO6kdCw4bfaJ7c3cJWfC1eXv0eT8Nj
FFKNtL3rch2+3w9Z8earAeVFTZvrInxnQBciDFbnyk21xx6aUbabTE9eoGEO/OuS
ImcYDxqWP4LcnTHf23K5KsdV3+8BUAKBk1FDEae0JAIOjwJU4N/FeEIuBx351/kw
lzK6lmDRlY8pPVwVsrgs006vktDaX3X+jPDeUrqPPtR8x0Mr1rWVtw9x2jLArS9h
P9Jp9crDj9FvdxMiaCl2Gv1iJ1uXwnGYVvnb2r4DLosYdFpgqwVvnTA+c+sCiVI8
fP7AZtZFwr+PZCPvKaP8W9TonTjTwoLdAEdT6pFc1FXV32VByzUwQ+uyN/2q0SYS
Vp82hQUMIGzOjwvcNvartTIIwydckCMaDx1aWcVSO2ZLSKDvJ61V8qNPPN62BhF0
M1eGExAPn5Qpi/qXMy4xVCA7BISB4Aexuk6RpbrfSZppy4elDAVWzAilpfctWoIp
DvPXPWfSAmLtsAoZ1gpVhKEJE8C3MihIyTnoyLHWVLGVeyvs106Jk0QITC5Y0CfN
29PB787DLXxiuPK9bOBrKD94FjAetXQ3Eh4GX8YAFDsZYe8sG1oFC3KT6jm2HtSU
mtbugjC5D2B4VL8nNHXyspEbLsL/C2jx04zrNsC2z0yW6OPSRlUQN20Bh0h6M5WF
xri5NcuY6vkrpEmSomW7UKKGn97zAMoVh89Egf3IZh78U08xW+An6tfjjTK7De9T
r6OItEmv4GftH+5g7St4xsI36TAzlEs0e2Hjlao+qFmxNw8orJgRhfSCO9m+SPDg
O/F5oq/3vrMbqmohqVeCwZtPGMWZ2dUoB9StWUPxyIT8JOi+GJluzGk0dlO/tsOB
FGr3AkSpMRyKjqlvF51SOrU8gYW9tgwpjom9gufKHA7/gPHrsCMW7DI2juLLZb32
yNfYgyXyArW+6D+78Mwdei1yI6YcQZg19q+dVcPup4M1jpYMV4xJeREjP2mg/vna
MoVyWpi/wNOHlkb892aA1AgSQbI3XNG+vd4nkPum6v0ANLv2BlelvivVgBmvqg5F
ZLBrixClCoxqurqNT2Ibx3gA+gY762b0R5PgGlS5MrgG1F34+TPY4SMsgvYUCXg+
xU6BvOONQ7xLylkJ5/t789jviASWLcOJCtvYe3e2uMTQTGTHxqoay/Pvlcc5LQ9Z
o2cANi/jhlMzOR8orXEPxjXswthZXXCtZtC7wM4bQS5WP/VWZtZS+YxygdpeckCz
YHXSXuXcjlgkQVmJ8taNHd/Nd2BF+ogNVBuqT/6SAiYEyTlAt+ItJyFv6AX6H8oY
vScXqUYtpyL1qcXO6VHy1yzukSdhThCXke1xs092gTyXOxJ6M5XjFD+j73e9s54H
0MTbfR/LtJ/xO9D6EHoUSTSn0ENcrTFh4jlAElm+MmyqnvNaLj6Jk0h/9CaaVvDv
ayW4z8RHPdNTWDNo/1/uMlBMbJ+yXSU+ynKqSfTiaeyOyl6AUCAYOtrEGZL/lOAz
X6GIbYbSKg8cwYUwQ3T7J9PS4A6UihfKDDhOTZ244vSARRkA7FYXpKdUbLUQTMdN
0+JppSrzsyUDQFUK7IUwqSXJNEXC1IvqGAjizbzdd92tct9cdQWvnf4ukueJR3Bk
MYTuMK7MBnf6MJrLF1fu6gce+6t7fixnkL8qFdFG7ScNLL0yPdjiPz5UQYXQUpaK
bMuBpLMMeUpXLVCbDGJp7/APzOvoiMR5y/p1NjrOoCkQ2TksdYh/7z/kIg24H7D2
gla5EwrGiuK6E8httiKbjgP37ofVSKvDlUWepWMvyyVUtUf70iphfpGP3Fz1EjMj
Z4gUU2C124LFcK1uACeoevwiBrmjO5ZwjkEoKsL9MZMO4UiHnEowWJ7UTbX6Ikir
ikWe5RhXM1jrHQshZe1ITx+eZLB/8NJFkayZBLll9J5P1Rl3jXm30M8/s1gRtqO8
71wsk29uY7KKXg9YsuzfvBLKSbtwOCg2jdh6fsztvGriWwRyNaSemkZtCl0ywVDx
noUlB+j19n0CiVfl+myFbyqDobMoKbEs4n369NJc3dOSVgndehSe2bbmwU4r+8hQ
llYraHNRzCxl7o/qZLZ+fdAf63TPJ0a+9j2m4WaphYv2uSyoI+rI9c4EcKHsFkdd
OeQa660G4ViBJlwgu1JlmqYA55hwkZEU5WdexqBJtVKTzDkjr+EUF4cGAOqn5k/k
7u80WFKqpXWY673hJm6PKnQgn/5BQV9S9JcBJpxDpv1kjShvJw1Y/WURLnuXywh3
6rE7Vtv2bEvasgMPNsV6h7X7aiPcDpcQA90tiq/hR3qvCT6HZa6v713I9PVGDY56
BnU11l1SHLFhMlI9hgb3qMR9qjLyQgiZOkEOoA3q0VNzypI0sZO6Lr6K9o0Zj3yJ
3yWn8NXOxIgQWQcqs7XYJ3J7H72m192KWcjATmifSDugTqLjT8sLNkimFofSYBGW
ELgUEzN+K43CfHs/Ie9kNaxl3KyI69N4pwt8ZzwYwv1aui/ZKerqX+vOCrMdzgsX
+2RvkISwdpsZ0ZFL8QOdDHYgxPno1t/KxQr3r6dF9dBMYnUeDJuluLgA66zqjLzl
Bnny95w91zaWfrhbi57qVypLgXwjBvnJLPFSym7w2gqHBZnFZiq42T+X/rscxtZP
Sq3jr8adBsGQ9xiboWt/HgWEr9b2f6AHMLFVPxkfKHKAdmVIbx0bwj7b7L0VrEwk
IUpjPugVYwjCHjQ5s76tz69C0OppFXIpXZAHEPq4Ta8/gf9d1tO2IVursIq7eFxG
YYdcm9jaf3jw5F6SkH+kQtRRTDewLNRWphIO0pdFQ/SqJev+Ga/gGqhPgKyY5L9S
ABrPl8hdp71hxyCBliEVF0k8V8JDI0lJojr+ZUoVtAyJv14xevIeeWaVN5R5Vip0
p8Vl8Tqau2cfl6z48NutoIaI9atGGWqCELAddnRZ/f74wXYncnCwla1i6PcrjZ1c
hvkrwyP1SwGQZA4ahuKJfTGqCwVeve/g4VJrF5onotMlIu2nvawDYxJ9l0tTmdN2
hkhJL7knJV5p+99SuejaUucSG6yYKoVT9ASXpCtylSCrbhHa59VTxMxAXMAbeUAI
c+4ArG7iu0QrsqXt7QT0JrQZ5rlR5zflSOWlEVXggbzZm73cAPLivqI+1XjD6T5n
jYWgRT2w3YzNS9VCkTMnPbKupbJM00hHK2oSPe1s0EcY4bJcwS7O+VLlDZvtEZXt
PKQGrFlp/hpPsq9jf9XLj0XTBneAG7yECn63bwz2iuJPFHoS0jBc8Udpp5s3iMF/
8nGeHrYYs9AF4GiQHU/LcAXkKkJZwyeUBnMCJM/ML2Eju3AMqXfd7ixVNXLzfifF
X1v7ffvIHBbaG0s9cMec++HqegA4v6+ymHf+QxNEu2Ms7T6qP9kd0uoncoV8XfBo
ZfK3v0a8HPCkoOj8OOpIzITYTg4OWWzF8uJzJweCuEEa3aPTwU2U1Com40Ir0gyo
djS2Pzq/NnfntdU7y0eo8D6TOVRVDnyMIRQD3AvTIPgRrbuBGKCtyA2ewn3Hu8GJ
ZZiJAkxaCX1HA2HAGv6RoYhWjxSFI9kBbLLIrGPVJev5I2WBnMBwFz0inb/v88iH
dbVlRz2IGDvy1UFF3Oipyh1PgO3PrufJannZoa+eeIcrAfcdwWIaVpa4swSNbZc3
Pv/jsEgi9x7J+fogaGU46i23q26uDsqToP0vkUFBAU4ehJH2uLbpQ5vYc+GJeg7Z
bpEqTbWJrL2lTMipg6QvZ3VEvYC/pf4AP3X330/eso+RKgPEUE1CcZEErk5MOMte
Z/niN8IWD+2HX/jYZnQgJMCr9ZHXbVU9lp4b9thnI84XYOuiol6/YNQxf63g6aZr
4RNeAZPKrYTHoGfg45C3BIgiPyQFpfI/usAZdIBMeHy0O0ytKik0IZVNVrw7Ym27
NYMG8X8jnicaJ1405GHz24EHuFhTF0tVfe+hKT4+sr4UPcqKjUufGpH7uw6oOEa8
7hlWpMa4H8pNZMR23ADCko7YdEhCvnmlxNvZurWoM1jKQCKkNNgQULGbrHzkKP99
Bl+QSgqbOO2gds0qdB0m0cLNHAUp2SAi20NmWnupCoCLYnKtgNsZANnGvh95RDk1
YGz4IGZfMXH5tGt32mDKEEK5m6jtPrh8yojHB8+Vxsqfs5hUxXoCN8feqYvOmPsO
C4vLRCTNaiZ+8n2e3QJ37cUzNk97g47rMCysP2MGGlqMfNn+EfW6B8FT5FG9MyeP
oPWLRu1zB8RFSBMGAAVWD+UjnwLBj8Ytskhc6jHZ45uahq+WLa8HD3hLp2hdCB4r
ud4H+uhejkKFHGX5ripZ3eT7CUf55ToBZqGJkHLy40cSRA04GT2nDKlBjwgrXxXC
Ab5wuNd2rcHB66LySmKO3NRokTgr3vE+LJgj1On1xv57ADHyeiXPGut3/m6cMV90
Zdajb5hdWQOvrqpPym7G+iiBNUZuROneUq5gd//KJoJ6SAX/V9WOqkYKsZm7V1mc
G3ElHSaAjOEYUw2aBb7w0A7XdkETFFOOC+oLV6IaGLga9SW7JsWWtdwvP6Url4Jl
Xm5PwR8m38AoG6CSzUsk8rSTMuDQAsQBuZ8lgqn/29ekVWKvy7Ydm/DqOHHGd1wh
Rfx3S4P7i6kwsi32y7dXvgBLNuffbPulDzKIfTHWrlpTRO0p9WRMX1lNXST95d3n
iWfbsQuHEfcMMT46t6SYw0OQO33fOlgu0C85ZLNHAbNqoIDGcu5r8Dm7/4WUiQJ4
7ThMh8aUMydDzcvaPH7phUTBuKgbTZr+OVfOsdebu0fI2suhI4EwaiYRtrrJkpjO
rXRbYJMFLH8VhqIwnok3ogMn3boaPtFU4iZfzGfed+KevoEbKAomqpdbuvA2OASg
uWAOV7cJOgUlaHr6meu4PzFTC2l71zM9BvLPfFxI7eOaUOwaCMhCq/6KQATEOlt+
W0s2uJD6CSs2enGW0FsXZafqKVD1sjuCHPLsQqnzwJbv5uLorvoUGo+72CuDeySF
G9SOcFw0TcMsbQDaqDfBAD5tr/rvp3qEwXtbaE9cvALrNBg3+guYFw8h3SQwM2f9
jFL9PHxzD9HGMJGwIrzsu0ruDxYFyQrf4CJIbfApsEQyMCmr7EDFIrBgSN4SAkHQ
rIW8Aawo3xgIJcfArExJtsL28RGdYnIGpCayO0Z+EyRVxNpdAoKa2d0FodF+FPq7
h+4qTF5laSp+vDRA9JP/XKreM/liaJVEBxF9/jLMUTvaPgjtSeRPVPJhNOOdhGEu
SAXe+UlfmTB4aAXOWhf/serQO4I+v/l7dMHysH9fCSyco7Y/50oTOJzDag/mXepR
OLeeK+MyKHUBfghfcmwVwsuGNLkl2GSW2ZLL7xoMlgBSGCoqUiG/JKVtHhyQWLI9
SzqP1NUavkZau+2j0RGeAhizjdyq/pv9He7geNn2pU6dJ4pKNWcGL7ZPLKjNTInV
qpsPrLh/aSFmUowM4ejT9Mmt6Q6CoBwO84rNR62+SGvOtMnBN8I2KUZvR9bLlFKU
C22o0Tx1q3yOXp6iHrwUTI1RhxfsZRe/+nqhh+VI8oYCkAo6nj+l9KFipG4jaG36
aln4iGNboRD6VAnh0LrRN61ZRlB6ThzpxRjR9a4gTFM+6VqugvyaV19a00wUNv1L
mlyWkh8JOhuBvkll+lsqrV5jvTEOroSCscz3nrzsBS796jYAkmDqFgSqJU6MhbHK
b4fWHpI/9S/t+3vFMUd++kNUtU4YQqKDI9IW8NqfazZbEgdyO+4VeDPWRi3Yt+zR
aNhOEEPi9UTRD/50osVdzGGJm5lvQ86oDfdV2sSdxQRjqbc9Oh6SOkS6Qw3hbzOz
mr8XtbVKtuI0NFHkU7Y/rDOqgDhHOQ/L1RCcogiu9PG8NPi0cO8a/KMcWAgH2p+T
ZKykVBeiyLeb+JjPVWMmWMtV6SJG695MK0sOl/aN8Rb4LTVE4tHgLjMVqQYvuy3N
IjeLr8zpRT4/YLLAJhCUAbTRLadEKr5qgghNy2Ubx9zewu8YX526J6pnvgAdg93Z
aLvQdR65HovACyHXRYYz4u1rTWOWhL3TGT24HgxvoNizEuN17IB+u1JxfJFEBq7m
l5JmoXzCv5UtRhS8unaQk+0jVUhg335yos4txe93GfuaALxl/8DEOgfzodj6th/5
J+19a9yXwZ1OJXrdMkuynRHehCl3xZtnlZmgcmcSwG4czDfrQ05sTX0Q+4IHDiIz
6c6fAZYoUxja3/lwqOu38FaBv/fWCVqC1WRBX61seBcxcXWldIwUyg3K2MkdEvs2
6uKPu917uuo5X/tIZpLRtYu9ysmElMGIRl/OZxGHULovxaREyjeKb95jdXy8cL7u
q8oMGwQtYu8hnuaI8YTFaW0eRT5Z121Yd8GeioSqeKxYr4gU5y6tKJe1DNK/Uhii
7VFJYw/P1IR+vNtDSuYv9wZUr0AIg8XO7CHyaRBB3Na1zF5L1XOg13Y7gj0H+SgK
qQQZkRhx6LBiXiMfFjg4gr3uDbGUEAMWIvlY9zET4IjVFwO+q0z+0db4UgugjJWN
FrkwJgCq8qkmWf/whqqg8w8a9j6bQSxwBe6YcV51bwEUl9Cix6+isw+cm90YZIZi
o5pjkzdneQ3r/EWLPe4F8vJzIBLuKVrO4x6mhlf/XIbUWvynqBuf+MY9yvS1MZQo
7G1J8kQ8VtNqp3YRvjLkrsNhOmIa3mf+Ki9VEVFy0uppg1+8UqpZi30T39Arjg0/
vgVOaXetgHq+BWeBjUEQf5G+A9XG58DzbFDmT9UtzKqBhahkoIPDRuKoXxpzbeEV
A/D2yII1GRUU3IgxxQTzw0uzM03PpZP00vsjGrNciiHL/5qUx0XoeNhiAjP75pmH
K4W8b6Sa/Cs+jF15B8q/WbBbZMzYNdGAZB3aPVBgtQaoo/0fJKPArZCFsU2MVHZf
/oUqVc2JbuEUbs/igiOAMuHEJQvOnVIb8HfD9eyJRqiv6qSaVkYKJoLrZstDTFJw
7gx853XQxm31GWGX7RerrutdHnN2w5+zTfDo+r0LEVuHTkSQ7ZvccmHC1jt8Gpj8
TplVKFD4aeW1TJNQSZEZJM5HrgQmwbGgKFtkQLxuE4YsecUlW3GbHHYNo8SSNaSF
2kUSXWGyqlhdQWlDw7bOsWFKASWCUFyItmNbhcKSI3f+uQqFBc7cENttXd+fSWk1
3Uzj1dohbm3im/+vCBVBb9H2miVqXXip9fXuQ1mgoZh4LP2VciSnlsf2yiZnyz98
zpqhiGm3h10cmQrkj8CrBYZbs7Po2gx89NYkrrkRHyrHwqNDa6KF2hKKHOxwAINR
hS6A9vbV8reBqv8+mBSzJ37/gkpcd1Nrmw0tMabJVIrJYwAwK96AX3DP5wr1J4Z0
25Hs9WCaGfh5ivjBhkxY/o4JlgbqL7bCjVnwWzOzdra816zsCzcbNC8Us0MJnSFh
r+KZObt4Xje4Sv2Mw6+MrIUVRt0EAhCBXC4djxn/FxY03UIJ/XTGJAXAatI1OqY3
a7w204nvSu87VO8YeMY2uC92Ywf8eTDT+rTzUWEv/JIJo8uEwkiaz/lMH2X7bGAR
tis98GG3LZUxPbWK/1sBtUcN7kU5lHPKWLw3fBxz5wwbYQdC34yq0Agqzo3lccEl
ogHlqQd0UkG8mCLq3o+jBjgN97Hjo6A8NZeVuLodPriqF6NnDVO61ujy7tETzxxQ
pXyK1Yr9iBwmofuFm8zDbn18hTV3iPd8pWyN+u+qcirNKpSTgMV/lg7szcDaxEhb
WVf0K0XtNRwN61PM4SxUOhK95gqvJCT9TPQR34VI4SQr+uBu6AMQDsNpbzM20cuX
JpwTlJTOAUVj+hlE9ILGDZdN/Z00ZyN+IuZGCESj8xxUftF+osOOlz4KxhG6YYgX
rA6tbvE4wThW4gBxd4B5YSH9MRTBxSz1ud429rQr4t3X6kyRgGIRz/nJ7/ftvdNn
rVYF1uDZTVIdGhvWbkSXNgs50nJt9K8fm2Mzf3pgx4NtHqhPgkAFiaUjFbPgGfPl
21+R9spRAq4/UckPLNtN6p9owL4mcwB1/tWijG0bgd/l9v6HxLyE1yOw3kRrVIQP
a2GuoT0E9yfFoxPjO3HVe8t3eGuaI0w469n8aqnv2gVvrU5cGssgpU8WkHxQvVB2
/8FVCELYgFT43LI81ZNAHQAkMR/uW7V4B+RTvwIDsaVvhAuKQjiVc505DsUgUfVP
/boyw0hu88o+wWmJfkJynjGXK5kmHQotp8t5zDx5jAmTlJ3uF5cAsa7PNejyfrMJ
N+OUSQanWCekRN9So3emRpGIO+XZRWRk8PZKphchUrc/ZQytshOACsHPIY0fmrHb
BpK/+7oo9b3fZ94HNcIfOXYKs9Y/W6V98kUiJLp/nSXdGS8cYthgrMdG7IB20IB7
7LEMlxfK1AY4ftq2E4t9GEMs3y6F1Bo5Kt0YrNwCihHx43OQ/9iDRWlIn1ke2Nzu
iWTrudHvfcXFpvfp934XxeM+gF47Q1SAwBWec1otouGdORPf3prA8d6s1sqEND8r
BS0YF4ChPxDqs4Us7stDy6cpgc/0EokTcs8gwD3TdZizHwGfcVDXqUsDA7H8sEoE
azxwm/jYEODfo5aiMP6dyk4FvZmfbV2LG58MhYUfh/XcsDwggVzkmFjEoKnWIyhR
icNLY51jXBECZB9xB6h21WubdhOPNcNCAlNzBpDQBGbMzPlXqdj24OVaSapDYrH0
lt4H7/BTEjcuGb0xwtEiJ5R0XMaGBfA/vM1CfEaRYK58s79q0kgriEQv1quq0u9m
y8KqGft3W5i0AqaZUclZk+tPHuOVpXBTTl87OsLvHTBGn2tA8PRnu5dpT8ac7T1c
JZnSzpX8BpL3x7jlaG5FY8N+iDbjPQ1NoA+oYyIYrWmFp9lLMOOyKclx7ubNbXGG
W5SDmzpXH3H9a7/m9BLBFEaO6tp42dzKAJR6Nug6B4aka2cRiHUuZrVN01cDjFGM
Z9lNb6pIO9VKCnXNLr3qOiYaKBwuF8chAnsrtCcESzY0v/f7wLPPKtEM3/1faeye
Sa58EYiKdw3JBMa3MhF1BKbjzCuj1/b+zotxBzW6fF+DuqwekrKBi4YNMzotwef8
FFWrqwS1sPyQrzCRQ9vPqris6Doc/WoMLZzkC730pGsU+tWqWvOnXOYeUu2/8tsx
O3aMnbcVbymDpODzdmyZIDDMY6q0+3q99XOkny02TyDyNJMYIH/ITIR3PqrU7T6d
mfj7x4dMhjfdeq2/Ac8u4Bzwl4si3tGMNpGL+rSWF2Dim+pc4XyZRBgt6DoE99Oy
orP6RFKKCpWM++3ukXUNgt45X0haoaDlItF1VHZFE/XSVlg97ln6SPIoPybXuzIg
W27oIpuAFVI72C/7FRnbwBG98YQT4827Le5t6ZM7JqzmrgOpr4X23zwL20dvJ3Na
hepneAJDZ15ScQRXDE7YWA0qx/mDA4v2Az2pL+6IwNkprQSccmc9NTddULNZeKLE
KAf8GL732ubNgpe6LkW89oeNKlddV5P8zkIVPDLk10JODvRVNfAJax1ChbG9hQGV
v2Z5YDWa8QbtudaxnX6241Beo+/LsoyDudyzocmCNH2sBKM3QNByxz+pRVNRNP4U
57foptYk8jkclvGJSgUIvrD8cPw29iRKsAKBRS3yHYVzQdxPuiPochQ7XoLPK69a
GUvvcobONMUQCJGFCl2bW6sXMv5UvIol6an2xcvD9Jk/s4tMYMOrU+lmU//99SP7
czJgrtNYAcG8oKDsNcamdg+cmLAY66gty2C/4Mb5WbmSsQUYJ5yTSSCTxBydCIge
OSeMsZl9vjXnWep502HW1wb6x1XvG2Rc25Ec7c+PTVsWIBIsgtKNJPPbF+UcS6XT
2CEgzL3kSM+PGm5KLiUqRE8VjIqEBKgQNZv8MxSK0k8ISdD3N5FxOtUCEqoO6Q0s
y3MSYp8oDdn1LyziCccqOBct9TgS7WrIzoXsFB4NVHnj9dFlwYlHubO7pzu1JHnX
VLluKSHdxqc1Yi/jz2A9OiFJNyOBbs5rwKbFiAA+nHahuzVt3kiZ0D8Ow/3Mgt/5
vg+TXOhMG5x6CMrDucwpoowpCWnw7iVwTBChffdLSolLfoaehxFJtI91Nme8rxFW
b4z+zIHQVnb4Hvs6t5n1NMuBbKpqUudv0G9d+TemlCW0uz5UAX5/WifO5FAZ4ldT
kBgjSboXOixlex3+Xpf8QFNuqounFExPpBPzboq3bCf68RYK927vL15xexXrcQDW
jdR9AxubD4pAuesCmpiF3iI6qD/48osbvs68xtbY1Ge8g+h31v875+6OV4ug+Y7I
+AgF0/ZDc/hn22ygiuBBqCaDmcFz3D5fbixA5JBxv1iwC8kmN1aZGXeoqVesTgQP
0S5YZZNTP7BxPq/aRkWUOoaWFGSeKQEhu7GpMFltCLJXYFpko7OASgzLduF9xxa0
2qm6KPV0P9PPYGtNOg4/AuMZMJhXASD/vsKPshlq1Sf+veY0cqWAbiPhYfuZairV
ckzpfixsiXwOd3oJ4rE+fWLAKaFLsiZFWv3KK96MtKSGIZMk56+7qiPCQC1YQeot
udGp2eOVNkvKSSnP/Ap2d5WzZDIXoffBGNRAXbVqM0b4IVTlIuIk1n1GuqttBmAM
R63rFhj6LcWZK5egaz5JBGISjmuKDBT92oJ7mrMofy+BJYOUABKtZknPvzHm2WAl
71N75EaCp8RilaTS94ThTKNIDGz3nwJdAQUyBLFCo+a4s7bCniTWAq6hehZX+Pca
8/fA58dpxcu60itYQgbEInOlMvM6Y8wektzLgkNLG7JwpQBb+CZBJUEcOl1fytYB
pinKPzuuwEZACfx+nOoEP9VmEnvW/jxZ13X+MFSclegsNL8law2sIUV9Vw/qXKbD
DmGai6P0ulQBhK9mxuwX7QTD9lJP02qnK4wiLC1c924tOrr81akLi6L3diZQfeIK
Rx4S5SUe+WRlZzMzhmIwe3RP4xTxay8ngDhEbh5CU0wrAUJVE/mpVpmK8fAxlIDY
GJYhSjU6H0+PsO/258lpdv2MVxFwnnsfvaiTqe9g7j4P7pOqJNR8s+UHudMhxfm/
+OaiU7ueySSk694InnHv/Ca1awZYXq8Y5bMuI/MG659JfzRuEDVOQ998CYdHuC7U
UwtllCPOr4FPj+EwZ0ULaIrlZBdS1kTn6qCkHmWlg4JFvMIC6uhljFM/wBtcwpln
6Ak4zmuv2VcpujdsJSa5/W2PxFsXHcExw63CGfdgPul6ys6+Oer0nsVf7eI95h2f
iQMtsvmX8QueGd5VTfwTqGoOWOrugfz06dei+ytztzP3tluOGQldy2p4gN/um+KD
dc0AvZT0xfXDXPubq3TTimw+c3C1EwJs7nb7nYTbI1ENPgN49flNWNopU4mA2tWH
CEtGAgZg0im7RrMIcQTKKunKOjVkGRbjZUwDvsfIAV4ri2/leSpHq5stl0OWVE7p
3IiwHDKwU0WStOrQt0dbdf7ejj8nc7QzL7Efl7EjNjzqwBu+rZ/b/BXvyjpiXQbo
ComnQaCTJu8CcvgbwtlMCcDguwZc6LB+4byBaz5Av56rr/HdCXOgwFiLnEJ6LvNO
PB/U5B5QNJYKHW1mUobj27sqS3VTwNHNLnpU3sLr9vtOOgeD4EnX3AmX9SaZoX3W
7awPSZs51OkP044cMRDru1vyIGzQd0RS24KWShYS+wkA3mVxvec1NsmldVIWGSsY
Kylaz5Andyo7Bn4U/xIFgZpJwDeFOrimAjTbjuTkfV0aMoCpOZXl3BScY2zFJxkb
9P3tH2GFjXoUalD+EqPzMTUZr/fYMxAslHILLowuM2UYcHf7rT9A8Rjow/+mqE/2
LhvsbIa2AinL+dn4Qf25lOAPSMmNOJkl3dh0PnhUC6ZoLNHofYhjB2Siz3YY7+I+
mIMyIfFEy6fLO2N6mzIKRP6u3rd25/PzJPWxmFp2yf/j0jU54dbTV8yr0RabanZq
Wnt41Tc5wXFyybHdE9ugjcxl5o1F1yzjCzbAdaGnjxsJukkzOO4aNRsZD0K2+ZdR
i0xrjdqtjdObgoJRNm9KWHYDn0FRps/7vRk2Jkbt+BE19cg6+tgucii3ka7kcuNV
5E+s0AP9/RoMVTwitHwNx5jNwfIM6I2jXuF/4kXUMtRStz11gHrq/KlXwFkp4haG
N3TsGphHYlWIz5VEZ0dz9ggrujFwlO9IHpAOuglGku5xrIvVcOzgTppNhmnTwRV9
in1yTdpbcIDeqIOHqKXE3RjzLYIMsKi7PXK0hf7EH1Um3tsBPMtiU7ms25rrNq9C
ucvWYjWDa6+zbEY9kwglMm9YTm0nJoKwng1zw6eR6f1c7p0iPoVlGxfc+NWAiHgA
X7dhmIOl9K1tmse+t3WZGdOh2uPHCnRAmsMSfZ2AGVaynMOy1nBmPiCFG3W6xrYE
DSi887eZZ7j7dOCJvGVdFj+47MWHtDyWxrcwXSehONOkj4haMjOTJ+bEK7MOE7Ge
1RpmuMAPjq1l/5VK10rtEbKEBdN06CCCOg16rk8yY5Db+G0reo3zyt7y86FqXwPD
TAq36Sd5iK7MLLdK/bA3hQAxaeCddn7VwZfAQV5/pigx+IhP83zpZdtGCXTqSxWo
8RGR5WgjfDe69NaHJScD5CMASjFMSc9CxgDxz67pnbrpC6tyyenGnvclByMrxn2+
BWKJDAAcfQURJEREGhJqsSfhoEdxyppA08n5s2yxgnNslt6QzN/bWcZ5xNf2lCio
23ctyH2XfAbT3g4WilhL3rLTL1XM4w76PS7kntmNmfB29wRMeFCXjSrS+NK4Ux9/
dUbFKiJqKbMytSdrBx0hMgRRv8DTllEQ9pTHQ+gHsJJWWjSTPdpC1oTsJhgy4wHH
ayNxMv9EsO1Ohp45sJlL/k6agM33sVhENZu+LH/FflSpIcLMIay/JNivgqHRe3sz
FuNNUh1utRaI3/AO4Bgq/+1i06ZRVlmqx48hYCAA26SmfDqXavEgM6MloUXC7xNy
ThJOWy0H9hjyI8ToyuOkt56P1pQoyiVxdFWnXOJQoxQipTFNzYFmJchXYcFXLqBf
CWWJOMnpMYkjKEcAh4ak3jVXkyGvXebEvQWJqyTDiDB2djHXzxN2J9h+Dv4pZRcI
70mQ7TmwbhQF8Jifls0KM7rukMTOAxsl/2cs/EOSaW8rf4mz5oW7f5sRAOq9tKAQ
9w67YGCCpm9fAtaa50jnZSWXlT4NzCV1bfKuTKX8M4omUvoQop0uPGjRywEa60Uq
fQRKjZd5hgRA6dNPcD06W+l6fDcKEKnErAe9Qa15zxZ1BbzaARpjryeL4i38SKGj
tzaMbXM99zDFi4Ex4uAC09gfxnQvqSl3lntBL1vmfQHBNfUJSxdR+6zhonBBfV4J
tjf2gXUbefPF8xtQayUJOQOiE90VaWz5G8GPzLjJhCg1c6QWTamgQWz3wpOCUhis
oTqI+ra9SC8tqNv1aTIZaJaFMk8ab7n+/A+x+Js4D9bL+5/gmyq8dRkX4dPqxTl8
SqpSy8S/JW6BUhvVlU73S40OMvR09AYXRwQlhPcvMIU+C24YlpWtfpQDFChmp3zB
s4ZKmEv3/rtu9bvIrpOt6sMNaZTZm31FZqzOUEWH42AaK+4p38gncXUWwN0PuY90
KEB3EWGkdtX+dXndE9BKXq3ALNdlV6/2nBRg0ZFhpYnAKgUkkbOPaRg9TdzCMWEb
+U5UeEx98OTmzMahfio27RB4DMlleSCd4DSx6VPXV8ciXDhpmCxc5IOv/Ncw8wLm
oF/lCptROviXnHu7qHR/ZQsmf07NkKyDqYfO25K6go4GlXAVkaNE9o8GQ9EAchtY
8gm8F8gOzNCvSiK5pGhbP+m8HMr6sQBPwehTa0thB+Uhi3ubfoNuxfS+s7jzHu05
algfTsmWpOsw2niniw7877yo65dDxbOR4lBvx+p9fmiowy4ML6/Amzk8RmkiERPk
XS1lSsxsBFMM3FX/kePPaO0d/9nZ+3iVLRckRKoKSHybCi3EvWX0yTfzjVgmJyC7
jOkjIdFPfuzR7Im5XIjfJBDKL6aLtISLgQanYsoe4pKN51Kpb6Sj8uyTSimi+AGG
eyBqcAqevjdclqzZJBglKc/wE4P1DApP48Kn+xm5UftGTYRv98rabQzQI0dwkYWL
u6u8e2y+IKuD/EASBeaNS4/ZIYBSZOR4V6RR9R6syRbxngyZEFRmlLsKthXg0w36
8p5ynxYbV6TwiOQgBnx2fFo7dMmice8LEpMmQCWaMwt/PBYLPSLmfCdl9buo1Iwf
94QxfOPX+vd5nNA3ENBLv2LgOw3qR6TDD2vFB8+nj4YR3USmPjNo8hh5d8XUEpaB
8fZshJhquXy80sPAnsCj7wCOXZw5KSz2t7EhD43eHS3BxhBeyy/hdaiBVDLJExVQ
fiQlMLItjmQE81yVX69r7Ao8o3xqtthJL93Lb+M7DsVn9cF2Jh9PIFxFOkCEgAtZ
ELIngqXd5bhb8dG+OOMEUahssKj4YrhEAKIrsKXjNfMCc9mQLLEGs5tn+OgKrMpx
Q5b0zJX3Zli+lsfN29QgTX1ixmpi9oKcjcsWFyUOBnZ4lg+K/q15M2YIGLzxBv1U
4zkiTpMPwuzX6C/KgU2Bxa38ZYoUPoD427tkYQxq/g3d00nqgqjiPmsz+Mn97kZo
vUsF4b7ua4heQ0eMUIqAhwj/7Gx6xZazAe6LDRBUcUYjk+1Y1hFc00l4e6Z6XGkM
qLv3b77gCi5jftQnLBEydkzubd6kPRHDQ8M2+Y9eosRtbt1cXr8nIhugQZRuhxP8
JiuTi+nDfVDJwCajqL2wS8IVxxF4wF5Bv3zOR99yMljbSkZ1bm3mlzmE7fCMWF7J
eeaxH/A00/MJa+O8smfiNwyPNLpw93kh5ocv72lIOW6oWvx9htafiIX3P/4PQNXb
MvvzXnNbeKTpSB9MfhJ4D1dHS4aulGDqFMKZ0p5dzSeAv/AXzrIPvQoOjeotQY6i
tb0EqH1Wa6Fwb3hPNQx1BFt0ylBEBGnmJhZf87s90DbmRvcwVOpmgnY6+ul5eJPx
4C6iEAkGBLZ09jHBs6OToBIyALIJEP27ggIGstE6Jb9xcXLW7a7E6umwkFuXe/45
DDHkuDsZKfrZggqP4dEYUsNvhK0jsOxkiDMrmJf3q7MxIPmhz9Q/vz7KKD7497Vf
6bjHy6I0T4aekELxPmcO+8hG7cITEfqOkxcf/31sWuAJVLzr8GB4qY9GPpdMUoNZ
YiZyCc+3TuMCilIbYPaeuHHQK9bZYX0wfsgQn+v7nBiAIDzvA1mEBBO3+FR19aG2
msrUm1rvccdcIACF1z0LTHA22QkJ4DTJ9MQiGDfNNiTPugb51I0Uj0V/1s2Owb3P
77Hwtz5djAVhe3+9Mw4sCqxgSVqkEMRV/yDPLbZPf68gSdV6spCQiNYTdmMoObX3
wwT63i4xW+cLnM9v8cMsOaG49EkaR+FgNuWbAgq5XYca6QuJ38CqXr5yEiPlmIm3
HJ+dcFHvuZCrcaWVWMi+n9doiivPrEqmEHxlJyJNdj6iYPYIgKvaZxSDYjzxtev5
pSmYNMRsAaNM1lIXC7A+1JpIUghVQJozjBWUXqpVAKB89JYkQJyCR7BoyJE8k7Bn
rpeb1kMz3LlCgX7hfIxt0kdUJHXLMJfCUfvNmjFH0T9LdcRm4Bc6A+aJUp7+l2Bp
xzZ+LK+YJOgf/5SJGnQ76qHJ11nKR8nd/W+IpwNuEIHXE75k+AtiyLp3H6gbz2i0
kHALLDDSOxB6LigpcwRuYTuzd1cv2yzSdNx4DS3BuGYVBIeTbzOnAiE1mLZSqGAg
3CoAaSFgMPHKtuZ+ml/9U648NRZ7bfh6pltsnIsyURauFOiRXHNLFbxY2sD6K8FC
+S2R/ZRRjMN4Td7pV37w/RMe58tQ5hqpc6ykfg0dzgrT2QFoszwUqHZVIrn2gFy6
p5OpoR449s/EN1G5GqQFuzN6vmbvBZDoM4b1C/wfI1aa3qMF4CnHWSR/7jkrKwZ3
hPzIHF88shLW6wmWKPATnV05zDck2W0ahheKnsOTP5VVsGZIo6ITjiAkeQg0BK8F
Uym/462TQdnu5KyYDYyRzKOIUPa9VNWOw9ijtpTctZGnHqqd/ew/euemkeHmxU/x
q6Ywou9uIglj/SxlCOkmK5QGOCfa+FMJSS4vIJxlh/D9o+D3EP9ik/iSstbeQElw
rThA3041ghCE5SoFd/M73f9OtqKh4CAoO3HRaVlsvJv0nuHbFJxvZGj0FcgtPcg/
3QWsVQkzesa1F0eOsizXofXSnBc3J3/NDwU0vK4QW5JssedcPMt2QUC4FK0M96Ug
uapLgHtmUob0otr6A+7ojQkQOuu+Nye54iXcv6tnyonh4oG7oMkDwRWGsZmKfnmZ
dJRXL7vLYuT2K7zq3/pHRW7p7ObensONXM0z9LkGccceOGyWkGwK5/LU7lNq9Tgu
DayscdD7p4ShhAqj+02djCT+ckozd8lMAfvD2QzE0MmeKTERTGeD65SzV1pLf+bp
ge0jGxaeFFWAkzjI0QTd/WxafogM/dJUhuW6wPXSmiNImw6EnaEi+0JiVMkjgp9v
+saO2LFrO6Z3KMdayS4VSVZ+qjF/S7QORr+vWrydKChs+iN8dtKxwEaKqgNBQRuK
FctufqVlDsJrG7wY6G1idSvJqw+B7LR3MAx+p/YZENtpQDxDLPQJsNirEZdPQHh9
Gjzc71VUmhxLKYcIGdG1IjxCPgjbCWUYOe73AJX0PdOnkGqpvUGJlIjfzWeU3p1n
5eCgxlFZuY/3xts9tda9jDPLGh4G/O4ipYeaIIsmffZIJA0Eyz7JkmRIBTAQE6Xo
aRmFbchCnU98FlNmQp7hWPldhnL6PaKnrnFbk7qwMS4fsHC9lf272qZ/gkRAotFU
isNsK2DklMskWxG8rhsxDMsW6Tls00jGJGBIHaRKbeArhrq5yLUieqbb3gZlpb2Q
A/SGNlHCS49Mllium/PyP6/Jql5K7oo9dTLuvsapFv/IFgmj9HLE4rAp8SUoM6WC
FTOGRjpEyHSFaJDrjFYmGKbrH67oTTc2BqXfVkYmbcJjC8IXwOQ30spfo7Xmcr3D
YBb61rpJM/RG5DgymcEOpHxu50NKrhdrp6vhvRIsUbD0oTQxvvkrHPROcU82NRN3
4t428+DqA93PZ6RHWN+G4KM5O+ju823Ty1Esu4wyOn0EvrIV2D7sHu6bNC03j/ZO
BMucPPwhKgEfSkbuXdTQzTkinPZTzEWpQZpGcSUm0Nj9TicjNYviFB5e9hPHgVAO
uh/217neyk+LUam2m4XXhd/+3EEkffFl5a/cLyWVg0QVa3B9khrVIGAlYSTSfLgP
rVDoQkP9hj8R0O7KXx/AgBnILWHVR7jAzte/NRya4GWcC1XhaLDTOXQ+NuEsZJHZ
pBFrIcjdo5qUTUyuhlg0QLfMjtr2I7VjBdRRybP97K/3t4eJEOXZK12e+yS3Em/C
tVm55SzVuXQfCnTRQlJSlmA1EBliMGfGQJG527GsAves9lFL5qQnKwqIOtEFhxlA
/LsMHe4Vlc9xKKIMIRPP8tCiNEym+eiw/P5lW5Xs6yRr3I9JTC0fmXycYYgBexkX
paPRGqCKSaZm4fy27V//FeCmN9SVf+ECNagJhWIH3fbAozI4l48qp5/unPaXBc2A
6jkVRz58p68MRVsltAZTMKnR6MArJtL7mKhCi3GUFPayzJMXFphkAas5qAu8J01/
/NdacBN+zskpXM89gfwEZN+yEWOSAB5RRCjyoTdzMxgX8mSo0gTe83UZ/FIaekkm
vSO8sUp5pk/drfgHGoEloh7e6TOFX3x1SXBjdYmEoPNo2oqyPp4CFUEovSPEVLxh
MTihxB01yQ31sAUIfLpwsK6U0fWy4B0P+M/0wAyvP3Smyx5YjNGUSsboqgi0NZeo
OCihhPIasAkuDzvog7UatK7Z4qgjYEDyKdZ1OjuGHTpSjA9EqDrtiRBuDvBbQHF2
uzUwkoCq5URJ98ErVXE4gT/8ygNc7j0mtHjkfcHVceQx5LKDryKqo3td8BNDzYI8
/wQBK1kqKv4N5uBCC3QxSjddnpUYqwhtNWbVBx8kPmWVSorcr8tO6/77efqO2WP2
PfHg09PZQap1XTyV8eR3YnHX8UzffJLjGhkh4Lzxmhmo5De7CpD55nE0+myj2dw1
93wLbiHElqp04lspPsSKVCMVf6ajT3xrmsm6V7gWGLZXXL4IsaLdyx0Z6OqKB24V
BeU2f1Yuqo4L6+2A0AZO82glpnI5OaKMmqkJPVLwhlU2AZQ/A0YJtJIfqS9XUnwP
UzOX3aEeFpkIlyti6CjIGdHFr8XrXPw2nV+WpigqjbwYE0fwC9Te8vsO3GfKezSM
HRWmzPMt4ijArOTC1KJvY9mbrVn2PhV8c2JZd6BprVWMEZeIJ5I2PHApNGGWg/bD
H90s3tQvS9JIB1pfdhv9QuiQwPd8FJ7/AWlmPZ0MqDC2TpaDQlDdtwBdDB+rHEfq
Z/atpWWtV4weyy6rLRIv8QbKp5NmkgNk04x/zWGLnGtiyHn5L3gDMpBq9UyJl1GF
A+SDxovjOph71NaRZGTLKH0ozo/dTHnpFLHfigdQ+3wq8GEA9OcdFbxxkzHtSKBE
xXh9gHGSa91Efdlr0gDARq33ktXUsE+uAV5A3WoBxVUEtS0TXu4tt5jKToARTBdI
3IOklWtNFcf5fu49M0v4yv2WwMPbRttDfrruyScHDnM/UUfkXIUpthZ1HCYTlJRB
8qguu86PudywQwXccUvg2n6MmJcGrY1NJOWPQrDldskLjbSPrLplH+m1b5fukeif
1GpRLozBJdqawHhyVfIydCgzZaAuc/bsNRi3H0qKH9UMojYwl/nMjPLe5YkXAK/G
1SitwvtheJI9F+d0OzifLsrWRCER9XPdOrmZ3WiX99mu8DC6tbCg4UNNC1N3+QAt
J76oaU/WOIX/ZDlf8AioUgzsK3XjgLOXeOkJtv9V8UTap4lhiVCnTLlRCiKMyzZJ
Hxg/D4G66eZw0JGC0Joap09h71m2BlVm3P89WUuEQMZoW32fo8pym+9wQaqgp7yh
pwgmhzpY2fBw4k/faEDu3gxwrzUz2i9OvLtUL78IrUhSuEvC1OQa1CkZH8Xe5GlK
L1ebBZe78/BeA/jq7P8nVX+hO40EUcddonVu00BlSN11iW4zEW3D+qYqHQOUVmu8
WeVR/h3lsEtOC9WzyQe8WADSYqTVpyJYapsOEJmPBj7TO+bhX38tNwwi1Se7Ve7D
neAnBeDGblA2ksaSKUM7mJ23LCB8fJxS8WeieXXd5px7yp+prhdKw/UuOjQ8CdgK
OXUCKuaH2dbFG1xqkmfYMjOwzi9Oy0WZ7aovNNCDZxBmWopB7kSkkVBqIla2liO/
IN11sqMCqax9YLrCa0PJ85A61a7aLyeSvMwv0tqI3KjgQTaaBbdhaXAoBGAfTvsj
9rshDFgXPk+Nfve/PWd54wOqJq4+3CC5OomGCYjgD7jC61fTWQoeIrxUuA0yw75U
bW2r2smGXlVGDeR8RhTgaPIR3scWDYbE8XrMJoPyovFPbxdQvqf4aIHcIWSpQyP1
8XWI4tPZXMpv0YcDCWssmctUixw4/9D5irBk2yl9LZKc8iVdzZuxtpGagrzVKVq/
zQMZ6q8I70uV3kl9dAjB0nab1n4fDSCYwLYHJ7apmgF7SWvxZh90Uud2elwHld4F
VnMApEincNCvuuHLDYIMh9ELgb7P3Pvbbi2y+RRksH4e1/78MwSybdl3fTDVA6Ib
bfKI3/fIswGCi1sxJYeSCVwn/+cw7Ebde+tdTxZMdrX1+/rOPu4Du9MyVfqnDwBU
emtzRKpRly4I5+yy8kP3AJSwGOAvlx5uqSh6oOIqYze1Ln1Kpoun1lQPLEDqgabk
HwA8WLpv66gviB4v6SY1dajxnylBI9rIUZudKw03yIB87anMSmvybHfUZvyGRac0
h10mF+n3UJzcWbI4jiLHYmaRlBbk9vQldgnuvkGyV94/fjl11TlJMIHfSiGqkBnl
2p77G2QVt91roWzNjLzgqRdChhOdYsn2dhlLn4QwWwS1Nq1V68ByNDvHRQ7XTagh
6kmmMg5LKIiputGTPmJpIQgH0/BG7xgrMVUnN9buhqRbVYxnf5MKTOLz82rTDLt3
rdnUjNlHkEeY6LczMneYNRmEstBdSq8pcD8QVHmbDw+ehpatGdzDODd+WnH2uwVm
5sgrpOXtwneK3eB1XCulpSO7O9ygysV7OC0yAM/oiKkFcykn1j8K7qIv+Xwf/DOv
cl/usvL28D5VMswntIoAUIW5NHs65ZIASgIC0oN/EDHQX7PBoLKvhTbXgAGk2Wg/
pyW6L4VHq0MXSGDQborLbLdFpHUMcK/IaZlIwHU7kvaggHR+QJ7PWbEAqqTtbhPQ
8JkZ85+6T0oW1oDFCoRhO2hx8tfCJ7phLYJyWa3VXy4tN2COMiduF6mvq20Ocrf7
9u/8bYlbs2LkMul+jRXBXCuiGNITCB2qBjapib2ewJotXDWKbk2Gw8TnjyTwkLAq
bZDsoM8JQmMGRCmXsR8u0/hPoqMiPFNTYQhvKx8kRaelLwsW56ElbQQ+ZXi+2xqR
KnaA7yVIMc948OZeDWuJEYoaJzBx1jcrs8qYeyzaG1iuGhWgQdDGDpTrb6jGRVhv
+EaDJZBG/C+prDJt0lstS9t+8dzeCvAUqeTfn4aQEQdQOi8ObtKzp+dZrROQ0R5Q
9a3I0mgBmHUdHtPJ+QPFg4SN8jZlI+paJjDYHcrMgtLDPBIcUbQ7HzGI6up8ep8o
0j8L1dj8lGBO75pPl68NZ6o6InPBzgCsDeHSXuIUk9+I/vCXNVcMuAC2khPMbkRI
yJC6TFusDdDNmAbIMCML2Vv5YSLMutp5uvyQXHDNNUaMUgx9VjhDEmK+iTIqQ0un
OBwxcTvdzDfgRV9jLxdHBA5LdsXnKzYbhIzXcoi2D4eZPhyLA8pD/rgnJVcQ0oba
EMgKRTZqAYZbNVzOyZHRYIKgMmbWzQI2Y4AwfppZwsigdQFqC79EfQpwie8cpENg
6ijupnkaqBJiWZtky47W+nHou7GP7t7AOAF7HwV4hc3Nf5IrJpmlY0v2w2pffaLA
eUuN0FdS2Imy7dBLPevinnZvpJaDe4MrrnwjM8V8s4Dp8Zu2uzZ1s7CnVjFNXFsy
Bjg/JBZ+obUUICxxNxtCk4yIsYx81EbupHe4CWAPhm23X0Jp6P3eATAYgu/B8ZzG
zHhVsXY8VQ9tQSptVyr3PuamemXzB3vLkFQnto3L9oBWvzmfgkkeLykZPssU41N6
TGB9iCGjdU79SmxwSBrI97T7DrcEGp62Gbrvo2yv4SBcUoEIe8U7ga8pPjzGEtr1
t31f9D5dQaCIyojMSwZuQegmAADO7njfT8i5B5N+Bi7J/EsFbuSPim3vod70Xyvl
+gi+5DMA//K9D4EfzTJp0ZjeVnImNxYpFH6LJx5pAB+16LJM+T2Lpg6OD2aQRN1F
mN3cKV/80OULRs0G4vSsP2y0Cx/N2nkznDtEqUhxzRpglizD4AwsIaZsF4jgjIpb
sptkh6OXCaAWDWGZy1HI9cOoJ/b7iC8yLwuxsQYpE12QbrfJHvej9W6wiUmgCnGj
Q4kh34x1CjVfwyWTDPrzR8AmYh2WqPyRZfaRqUj5jdcIWJB8zKmyLFuigj0WEJpU
bqDK1OJPNC1+Q6UimvU2581f6WNhaKq9KocF24ZYCZiHIAmmA5kqB1bxZwu48uSt
VchLvmH8EV15isjbUQ8uVq1X3jmloe+Sjh1ybhMlo3h9qGoWDV+kFw516KeNsjh4
JMyOUyY9k2FwEbyfViiUq9Gwusf6IaU+tpJSn9xbPYJpdLAqvfcFCuKau3GNrPz0
/YhgIoehvjTTPddA2U8ThAV9ep4CYo3uOrS2NZTyWTg9Pvm13yrGDP9I4aN8h8Q5
3/9kobd6s3P3Q4cvsgE/+gHGPEPIeVKeFd58hWyQtra9NC8m3H0+bxnEjf3nv8tQ
gj6s1yPXW0V+lW3lB6qrkOr92jTtGZ68kl1+sUuYTa/76m9NxL1c3g73FXr7N4KK
ASiS+4qxXXzyjEEVUNhJcalp9vMQuNCqXtTrK9OxX+3RWL74UucXTwiAT0AaxjoT
BxPjrrSz/tiIc8uP5/BM0VAybpwzi8dDerfTfyAJelQmxiJQ9VUa3n09qxdjNNKT
fDmu+2Q4cp7uIVswAk20cPaYq6rHjuFMQu0V7HpUOOi/YChTWT2eg9fyFYeFFI9E
RoBpKNypAdr4X74mLu3mo4g4mD0DJRlsNxRr1LGleYXEwSJySIdCj15xEbGHPbQn
FzNrRSrlDJfCqLJmbXykzwRhIQHDVEThTcnidh7Yp+7qZtx4V6/XXDPR5bk75VAe
bOhZdGNAa8CTPtsKUfCAJrVGGjeImCe/v+4cgqp77cMldSMU1SczxeqgvPyyxvGs
hOqfHMSnns1eGt7rYfHWbp62W6GWYPIG0couLsRtf0W7gmSF3h4Nry628y/ZjRgL
I363ee+mMBScMVDp2opcBD5YQkfC9UwlppYl6mCtLPDN2Zk5q3zRRo8ixw5m9ld0
gAjOqiIQbT39ql8XKQndIyDJ0WxTfXTxagRsVcqR8sPkI1Q+8T7C/ievcG3kGcY9
CMHvqtkDMHa9fNZaSuFgYeX/HzwWQEwBl6NwweMH/zwJApXylZImi1QtvXRtnKDV
4+kba+zmgBELsjYREVwPSCiCyWKGy2d7dQW4u8asIFK3DbfDoYlqZIi02zPwVk25
og9oqdNukTeQzNC1jNxZoRcbR9xLA6+0K4s0IKBo6SNkJz3/AEcfUsXzS139AiP0
3XmPQyYtCvUeyDmXXtJW/zDCEnfVwdUUlZgDaw2A/0D5DHYzkQlcIE5qebTdvRUZ
VwyyfH9FyhKSVa/YjqMyvj5K5LIU2TzbJFAYGCBXyJovbnwiKlUsuXW4oA01qH7f
PL/GG0pCrTOAT6/F2sRV6LZmUtq1spGuvPo3svNy79C7dlK0uJ05e8sibxIjIB5B
ExIZl/wCB8CUl5+lx9MQLkl6M4kfbOuzjQcpJun8xBIacIjPU2kxSDfRGROwopq+
aGJUpkWh2W6jaDtLgwFO6a6Kzg3882ce9sOK2HwSPeSB6Fx8GXVb1We2Z9zKmday
JZy4slN4eOA1CvpKh3iR5b1Ezj74ca+F9k8aOjG7u3y6f83IAW6mzdNZuVYIxABe
yAkFHStHBWkMmssWGQct//Ys3dgVxus8+1oEnf0WHeFuFscxcwY94gWVOgjifqvZ
zQSEhEHvrZuuK7tpw+4cuhgcozVouEWw/1sfgFW0n4Wfq/47qZ3FFc54D1Y3R4sp
F12A+lZyvfkgo9rEMV6VQNZ4KRBMNg1XWWMDe0pOkicnr5lAz3w6fRUxqV96FU4k
SC6R6stbMMAu3BXCvRneGXUb7faYXUQMvbtf2VrMoOLm9fSDmx/Z2FGBW+wvM/zU
KKKkn+ioLSFc6+esBPbqsEuP8JhZKEEZxOye5f34asuXWAugrgC2bZI7Uq1H6tc6
a1ylQiO8JyWjKOnh8wMP7Rt04CaX88oKQDN9dSiVkPmVtYPDqHfIjFWLgn59e2m4
sbqav6mgEMoByp7aZeJAdPbfV7MgBgvuuyPzKqFOB5dbCKl3NEbT8Ats7yxTSX9e
DNah3lm731wykIJEyjCbG1USSN6pcEd2kb2pUDrBPODRDp4mS42SaTnE56HW6kZY
WTejfbYw432O7RjmPXKqVFuoGYZTGASF2EYXG7l5mKbLquzzvVCexppd2bOU5Jhv
VIKyQTn4N9voeLz8K26b5Pw3iWeQyOwx+iRyFGdpZqEiPxJpm/VJJk+tFIcxTXj9
remJ7nHZofnwf4qakLHs+d27IOnpYcblIww2Sq39Zys+fKNbLSNvCMFay2gJrh2h
lzNGwI7TvNqXLPZ9yz69JC+1HfNGmK2LoiJpOwcJwnHe1AJBpiDVKmDvdmQHVP6K
z1yMqy1d1b0fJD2ARwmQnSkbcOi3fwhDPhA/a5GFIm5B1BBa/1jn1QAtjQl1AJJH
+iy+B7njsTMQ/lA7mwnEWTdnZ4fX7R76WFhSoQLhWVVyg4+YXjdK5gZpBSWjlEvQ
ujIfrFVBBMR8cGHFHVZ2F2uNztw8TAB7+3KmL4NCdQV8qvCZ3Y/4Jdl3WB1PxkfF
lUrrT37YvZxBJ2CtVrmCxZ4702Bq3AY2/SQjX6QprlN+f2fppkaAttlzg7aEmRF/
5ivm9dnQ+A1vHMeOBOW0oxPGd/DDlGVXYC7qofQfQS9ENLP7rSNMg0RdbIJeSomx
50BVpDQk/uC98mNU5aHt/S/VOXLvOuTI3wO/C9W14eUkB+zwpSo04qTL+3XRlBMj
L5Jb+0s1xOi8V0WuR7hlMmhxoqhabVDR6RX2WH48kZI4urjcVVYZb+NT8aYLye7e
c6CdNtquigQnuoaFxFFql4i+Ha/3oh2fEpre4qXRcz5MmNrVyH+vy0Cx6xcpwz42
kjsLfWfp0IJ8qHp4U1ZdmVE9EeHwQRrrIAyf+kwdy8uPYPaMaVJWXM18TfX0sZgt
M06LZMXm1KsURRHYagMSiB/GKUSryRchfbCriLNh+OwWW+tNE6tP2LlA4niu+t2u
fEoCfuDdJKFl2bT0ryP3Wcdq+6fM5f7jYbgEKrdzvZfZYWxWzWaTuBg6B9bofXY3
Lv9uwK7aAarFeEwEI767WrWnUV3eiDdg2T61zwx1o70Iil9IHVo1/dS+qJIOoNWt
do1y2oZZKKGIbenzS8S14eM5otPK8u8heKiUr4Y0XzouozRn1aC/wktPeNY8ciWh
EwEhlQNeuSx6jEA9yas3yWVpr4MxJ9q/nyazyAiTSyn+6jc5VSiS6jglLVvmu1XF
dU4zDKKbQ5591AVkLlR0hpSIcGAGqulCP395CzPuzeGxPf3dCDxLZuxLcOl2cMBS
KbRVCyEgQl8RGGmQx5Ph7kYpno5kYUkPfwyfMjAuK9Y8W4pY31xrHyxXifqAG6nm
HPDKvVRTOvcwZKI4rmUw7PaJPxc2rATN9BKLODDBVuMMP662onrFqd2hWLy/5r2G
MnvN1h01yqtcXFZRTicaE+0eEwVTLd3/sGOft1gV5YQfWDQlavMLbK5g7yZwc1jc
RGvZvdTS8rwIVLXPvIU7267QZ/52M2Ent7mj6Cot9yN2RPyG0gqVuAJjrD+ZyN8d
a+PtnTdl2m/tJtwUlcL/kFtYOaeVvISnbEnmPWq/hb4v8GJyNwvZoE8Oilyan71p
bjXHNfiTPUcTDSjA1mUjaimj8G8+KcsrL6YoJke9OFe5Y/pkBJsTqdX4yIMRBmCa
2ekL6lvZWkutMiVOEQpHfk461UsaUCE4W4MWCGf1BvU14ugLCFb4Ei0WztUFkyuB
eSzE1lhd9QAY/PUV/tNAokmKIcijwA0RIvJ6Df+WlaWDq5Gy7XWdI0cgKYs0POPC
U1JHAt3IYFebYQi8TOkFnldtcLcwdyvXaUbPhoeUuhCC00V+HAAlaBRJ64qZerYw
5dqEcmLO/cvxdfhpClOVitF3QHcxyNGSpWJtn7NyispMDruou0wVj++w/LFYUwX9
fS+1ILWr9K+TKeQS2BA+hX/oGMsaF84NYfgdT/+lXl8T9Ime2r/6n9MywwALV+WZ
4xgniNzTfOMGWOLf2TTW4EWjmGsd7y8l82ShHvJ3Ur+9vmuDAgc1mk1JvBOodd0t
GTbHpO2aWhwex9Fl+h52CmYHyhWdJOybeVB3eBZ3zI0hIRxZdHJOxk5rD1e/PoMc
yh3gS3HPbj/tijOKonJLADaf2dxQwVUwaVj/nPT1m04egV8N3twtAvSduisaewCA
Mlgw+Fi6ty6CcbHSbmEOFCh1H5xR3yZHGlKG2ZeBvUenAOlSfObvSUjLXPsa01tJ
76fFJU8fhCduss7KYLh41wwUp2EvRyj5P0jdB0L8zEWQnmZmYiXf+NeNYujN/ORn
fP5GD95CNrPUPZd3gbPAvpa55bXhNy8YxjCFn8+b3f7DGkrpQc8kMMsMSftzKq+p
R24Bu6Pq+OFtDni5huw9Kei/cMeXP3M2DccJVISHchyAzj9WnvOCaYCZEqhh9rDA
khv/5fSMNIwMDMVJbo85lyZyrgtKym07FExS3wOuDIwVwU1Dmr90U0lmUHOI99Kk
TTad33NzLfodAcM3rIh0T2CDClp8llJUW8mPrVyudIdQhJfVR9+z+YozscB4Bebp
9M3jQGX6AY4GXb1HRwpLLZhQXlw3j1VRtw8WeGHrYMQT3krFbLIsdTlCeLJOWIMd
ha6FGx3Z3u7C6r1+r7UfjAIs5KkYk76W8/FQfQjrZ+4C1Pwbr7mA2ThOIaCzAHLr
omSl7vtHzCy9cL+i4fly4F870iZUfgkAfyhUe8YfDkAIqiF2HOKLRfDoAwo87H/N
cMBEVoj4k+8fVU8CFLBHU514FWXMicAIKHwDVUlFxG60iOMSDb/8qk//N+35AECf
NU2JsTfjIexi8mEG9smLfoVGp1V5sDnF9Zhb2M4j8pfx+/fbh9YMbdsmqpdkq+gT
GYU700XJ1CuJKtIuvq3Fwb3i9E8ZoBl+xD3tHSke3+v40BGOBEkZGy8zurvU6VLZ
mXyiLNJJsQxueVkYh+Cd/C9r7gl7zljWxNEpAciEHfzHKXzgIRaoHCJmOoFu4P2K
pbnAUHnD2Sixq6PlWYIREURanLj6vMND7P8tSLVc3Sr3cRgGG7u2DUbNJQSxcErM
BZGbjpi4e04zsiJq9zWfPi5fOGoVebM4rvQ7HoO+54eccbw4ov3J+WXFlhUg7lX0
yxnVW4U2mcv9uCOGFCeLl3nzHl+CsUYmXJqjCtIAc8rPczzEnPWWxxycGELQ0IAz
vEQ9O6FuHM6b44EBFQKANlZ87JrXHAEZ7zHpcD4mMjkR0nsYZKSUTQ373As/V5Kl
VFgE8gKE5OA9zMDNk746VOL6jWkDDzLDUP4LC27MtwuGQEqTgCuHwbIx27ybHQpf
F89R6uRV6+ICQmcMyWDkXaQRTn6xcUObF+z66az24ZU/h0bvgA/i+1Mb0LK/nsrt
XLDmwTyORoD0gF9EfdgDi5TOpjtBYQP/szB2j9yguyTHXXhL/omL1tQjqPfh4avA
SSTTo2zt7OJDBFpX3EUbpEtLYBlUmnF/vu7BeLYpCRi4py5FYHZR3wmHe+Bfaflv
++fRMLNYyUUJwZejNKyPwVvOVzKFDihSAUs/6s5jBIPkQ4Jgqh9fx2vTMP4z+5CC
k7FKT4l/H5ZK0bbAeEJsZ7TlH1tsGQkTTfsotF3lXMWp0CSoazm8a+PieBN+k+zQ
buKNRPzRUbNPJqtYaOERgYxah3frLD//AzDAKSQREcTqf97zL0NO70CYHoKJiZU2
BIW2+0ReLyhxw0EUDSWzy/eNK8t/QeWqN5CQ9kn1C1IlMrehW6JzlYwAWHVY008a
SiJtxB2MIhZHPfhJUuKUUizrwleYQbGG0r5oNekdyA7X/YWgTSvdE7wdxC7T2fVK
WX0AMBAsDGt8jbE+tqwrCyW1Cz2EQs3otZcxgxcaG7vRIj7M0lpaN3o5dprFvWFV
qTq0vGK+jlOj01V5tEfIfSO80BPEtnX0ZL9p5RvRAvBIFLN/wqz60oGYLbaUbvw7
KGw4ZrOYmsojVSI2hESyBOMTj0ImPpyPbwECLsC3WocGDeus65rYLvj1A2SojMWC
/q3jKPp4k/fXdl0ft7JMth9GBUOAxwoGUfNQ03UkYQf3OpxIYF+3RR0TlAJOdG1o
vhPBrFKaAUbLMfi3mB1FbmPZXypp7ecp2kIIhNU6F0qg8+4LJ/FxQevaUo18+78D
yuB/EwuSy2XIzujKmCEjZtzkqwIfusyHEUqrbUiYfdLPS4dK/6Rmpa3QvqdZZdGI
TUBInocfH/d35xz6v0QButqLSaD9MuiBWA+CcRxTH+R/fpDJhnLhkpbpY11QBhVs
7iog74IfeojSD4if2dRqycRWNd86NIIRb6XS7PIXi4wd/jRPdDFvJpoCQKWNkmLJ
7MOZDGUItJ5KncJMExaldSyzSeqpx/jBz3sGMUjLN46f+Z3wdo0p8fZ2svNiogJF
rWF1vQSeEoUNE2llYM1y1Lkw8n9pMRTSlLhOrWVLOauypeUPkeINhR7XQ0l7X3FZ
2HPBgq2RHWMpVdvv62kYCBae2CEnnLhlNNzuNIs7NrfLT3PX65EObXdH+76f8kr1
D9TeiIvsKKufpaq8sW0Q+R5hDI30DL+LPiUagfBChevXUncI/F7TCK+KysdctxEt
ofTN08cC/sMm/OoqeBAYMuCZMUhB4YRyKbGZB9xGQJlmCFIE+20X1qf2hIWJgIdV
rLWA9hAK7Yys4PMZ3OiSqJeUlzcqLUdfBCufkgYH5XnQobaU6qBNZ4GLDcHVGRAr
sbfVHBYK1mZGUMkbenHa3tDwgSlp56iCVeQ1Syf2xg+HHL9C9m252JA05x2WouuY
QsyFOarwNJ84jnH8DRwP9/sH1UUxiRQceoBjoLOvU8vs4EhvMJsX9f9oszQGbg1q
KB3aKfpemzY8ppHBkKlo1y4eqs7wvKacZ6yrz59wg/atKyO0Q5S7OoQI8QB8kfkH
0wlXegakX7gG8SzLkMUt/Z53l+WqUcyAfqX7Kauvc1JW1wYOcYQ77+KWFYtJHKmO
mQ0WezNzpgIujfHoM2Y0jI6n6zsh89CcmL8fXEdm6aXGZRVinaQySt7Mm235Hp/E
7g0g1rH87M+tM1mjMBc23GfUhBOVWhS7soOrqYdxs61NH3LDN91MUgscbH46rc/B
7FkqNHziuz8VAgThSyrQHXkPSWjxHnVrp6M3OOKeuDyjnduunVy1bUUFlmt94frI
hqCXw4ARIRKrKEkoAO1lGsPM91vzyyvDnPZNzpwCAGXzN4CgPTEFv18QXehTJram
Ejyv3OCylJg+ufRA7Bp5VRmaWC76riVaGtdc/MglDbS9TqCT7iDtAyaFpmvg2wC9
rMkxSEPJUJgAyohYQtnt3KzlIdWE4qllgKEvx5uHinsFoNFuFXR5RK8CBipDys8V
hodrRU8zdm7TD59Z5AdE0DIL7nC7josHYF3ZIhFDsr2CbZy/tiV1qMcvcQHd+3ML
hWSUxBEInit722iljRqPYKTOSwaX8/6LQ7Fq0X/T8XP2ep09Ke7Ue7bVSojNL0CN
g/l58PqD4IXiKghpvDJoeN+5D+Cb/U21JwjypalJjcPi8kpMUIDru/H3xMn6O4g4
CTPAHsN8dO+1UpzUcbGPUUIksN+GLRLlq0aCCnoJNbF0IGYmmBGUIVRD9sQzp98z
mFfdtZ9xdQFB92EMsm302xpe3ifcmOydQ4wQwS04GC7oHNLvVJw7pzRQIqznBvGt
a+RsiM5Tx5+X85mqH9kqMiLWwN38QZhxKn74Y/3gVZa22xLWdGvY3kUAyn+ARlwh
T+msdl3DJfaXP2uvHIp97gXnIk1shOJB8kSdtCkFM3dSc0p598mltGRid1Zbh76x
U4pxhCd57UozzWQO49v0xJD2bXSfv8PsPJ/L/eEaqt/bEQyda/59bK5K0JaPV7dp
rgEtJ2/qZ568nwMqwJgOQc+2aU33MaVSsWmMDHUkkv/eXcQqEmg/8aJJOp6AHixL
CbsUZL5w/i1HTQd0YSfmx2MRyvwJRegZfL0mZ9IXvww6ov9rpR+0phP2wCSCSvrq
v2HgGK5jKDBXzPVUtTqQx3muz30/NybINY6qzWdo/7sAWBmOCuJwI81/JFTaVkyS
mkZ5pHM1s4Foo+tfyFki4h1jBgOKadD8CX115fKCAZIIy/0IO8Y9nxbwqj0mH3ze
PjNdifInsX9RN01KpZoDUny2DCXfq57tl+HiTT3hrsuk+KJr7G0M5fpmukIgvdwp
ANr9wX8QOou5/nG6PDEK0w2WSaJDLJGzjADm1sWGUJeMXKV7xomfK8c5Z8yz+K4o
t5/x7I9FHOtAGCGHDDw7mpu3W5iqQLc8M7bzRKu3Y1cxlNeLjm47DJrZWmXEAkQy
xleTPUD9jCnq6YyI6VgO9tEm9M7UpKa1hlqu7GUmUOB+/8POxJqChAoEF5yDhiZ8
Va0RIuWOipYuKtAD2eJ2wIwxr4XG4ob3UWIycwXcjr3nK9QCd/ru2N43hbTPztB4
aULjbHB6/ku3dgmd1WO4c3urFYhiOEZ3Yqsx00rUDEd8eMmVeyI6WqiJJvo1rSnr
pylHTGtoqJZoFVkBOOgnFtGVAN6UBhyLCrw27hTpg2ZQ5+VKWBorfmbWn2nsCykx
78F6WDKgreuDLfcGnU+vsHBZf+asF84jOoKLu/x/B0vvwaewbSegtjI2f/KOosER
D5TX4fp9LuepGWveqK4gdU6IxfJ0ttx2s/FEBaf4rOiw/pd9isb1nEa0Rv9BKZUA
4PBZYvwt+FMwTmkZKs45AbTSw/VY4togqdlxYg1pDU+3702dpir3qzcQ5DedttAU
iPO+0Smb0coNz8YZVmKhKQLHxLGvPBRtNlByrQy8LVzTIk4pFS9EDVyjp64527U/
e2cDXikacGQURnRu7tjOC1MMh34p0nEWWpSF2rmPTKWnepi4gFc+Pp6Zb8T4qBqZ
5L9qXL/l6YpJdFeqrHZ1yTEKqd3RC8Ro/c81D2DASAGwNCM+eAzfNjnH8C6qcyXy
PqPsGZYf4DTgD2aJFf+/6fwNhoXAHhuVAVLDEsa5jNOfDShBMfl+M22kEOIVyl1i
SytQ68zs1IFgtveoYuKdCvqysYF0DFwAYwdl9jEPuOMaHZHUirJSX+z/pj7UOnFL
z/Pl3o5DpaFcuwTIl58XHA4RSoRozfFe1R4UiJqAKUYgaWaPUrEOLI8pbxB4OpxG
bi5IC0qA5GwVj7UgzOP2M1OaiwfVx37cGnh8NwPr+9xGvG9h7fAWOv1hffX3V/lK
z0mmUOYhJicmPcoY1gepFnO249rst65rqIKIE2+LJvYXz5NNzh2p/Sm3i06h+Pn1
1TtWEZdH8+SgkoN44sWwfi4na0KZhRbwNquoMXKXc3oWPw/RIjf8NLW+3k6MkDx0
EqulCrH+T2d5pnfi91O6D2dNbReDOt56HIVu5GyfFHQt9gyIOkeeIK/n3OaiBZaa
EtXc0nl8oBJ5EEI7r8qyXaovUcvasmbCfpbYnFY/3O7F9DzFvK3MLtoVnn2oPdbb
Wk7cvVDZw04BiDYf6dcrawkRGoBQSSQCxJKC5lA0V45b1RpjDisQ9jeqhOUWMLEy
bHiMVdK9fghDIi502GmQ0puQBxF8QPmfRcpSoAPJMst45fYdWaRAOciNhcd5wCWj
fQAnSYnDAVyqrztQeic8Dp0IPp0lw2nbFqeXIuGoNv/vtgY64qY1flnCM6kpO9dJ
nLBKMcENJpQL6TlaRNCLfJbQgqQW8o5Ze6FXHMg3lNtg/6xWV/XRqnS5XVMrsLQm
O0SzWT8FlviHzx5nuo+3RM9gFBKIUI4DUUWJHV1ksf2NDOhaijwEXCXzN6CRCsIo
ERdg8CQwM1ZUJos7u30F9I65sk77OAKm2/ft+cc83AyM+Uu0xWmV4nA+goq4SNrx
ZhQZCWKGLa2IC98TsioDOIYVfZMMdQH+fiTu2vnAuetkhTgtOFDHb0oG6d4t6z7i
5weW66J5h3NM/wqN4Uq2fPoEDvgdfUkHWib3DZbJwTS0M35M/aaP2otSXxsvSlzk
QP5batnGAn2xWe2fc6c1lRIoZCvZhwJxB7MpEaGMUVC6vJVf3n611mGpxjxM6wWV
LoibP7grnyocvQ4eGrOZMSprffG013Iyu160/UNTkcqN4PBb+NFwTS00Txp8cJ3O
yd6oc0WxB8BACDGT7TXweV0sMxlq5Jq5V6NL5BCafsQ5/LJpnv12FsInfaHabdWg
RqXt2B3CfBwxfMQKqo3PdAqfGb23IQdyvgSWpP6KWHhPziqv0+Yx7LjqTtdCxRK5
OUsZVEfGHqS58Rf6DStnKXGMxPP14haVTCuYqng32BaJ7FegSoxtujmjpXq1Ea/G
Erj5ucs54/H0C/HSjimRRm3cnkqz4cdV4l57bqQ2w1yWQZIL63FJmG/wuVzzJ7+R
Tf9JpWkkSABvW4Fta1J5KbqIz+4OGmzpX3lKGsSNJP25jEWdWZ1NlCkzimm4sY7+
GVFvps9hx8yBRP5CdTJ2u8KELPc44kHZNjgSmECWjPXfmNXtWcIpBjgqV4XI5dVH
Srvvf8UNb7iWwKLIdU7xaTcYWVM210fovPYgi3O0mmgq50ih5Bl7n+zQre5Zpnu8
rnMS7skcVblTmuZhMLkb5yJ7pdnQte57vEMwF2/ktc4IzH6xrLg39zfzPinmggWZ
tYfyKbDntOEsKCBtCwj49KrM0WZtD0hz6yR5kcFsSn9W93R6DwtHUwqwJA7ibVwj
Pos8CR2nq6xTxvaXDAB66TkiOjNr2rc0rZqQjpfnuHDNBrjJBO+PrC602iNWv+S2
ksORgTYImxu7RJko/C7FBrYQSKLcsLHqYaIzj+X2Hwifq18DrhGxHovt1RhMLk+T
IieCfU2iDZqhZRF2WeNCxpjnCKrbXgt9WlQPfsA61onyiMmEoIq2PgsBsJWSv1cM
j66m9xXXuNu+YDQrGpFnT7ag/gYbDLq70xLYZm0pzr4o3wFz/GF0Gv1Mv/Ss207m
0lB14QwxnrcFOA1WiOszmXpfiyuzUeTChTrz9CxHBQKCChqLgFkQm/qk/p8Ywu1S
DmqhJxKuKNxR7T7rBShFkQE+5IJGzuI5faxshMfytBx0awwLEwP0E9eMeO2tIfvL
VQcQNQA6Lof87hl0m0ugVLuJnD0fEMZ1PA5JyWR4UIpkQ5XYS12V3Mh7e9jFgXt0
FfuufA2Kg3dK34JXQdeOva+3iBRMoNWxPsgt7ekY0LOkYHQeu+Pupu/Qqtm5Qk77
FirTtl9KUAK3sikF0reEX36y33xGxBBK5wGQTNKCqR9YiPYpd5XkN1jQTE+kTrVg
1QlHmVAZhwTAEAqk/B3RecC6FhUWJKtCXzOvdbqniY/xzN8uY+RnwKdGbRbV9rgT
YaBt4+l7ThK7DlDXgokBTNXgG4uh6DnsjZYx1mDMlK9lCFi2ZIwH2DvuR2GvGIFP
9elEGt/CycKl2WRfRmHjiiCPCAUJcio/2OkSvETHFKQCbvIRaU20DZW4jDW6vmVG
1OO912kuYYr/3Dhb838LLvmp+MXfYUJ2+tdAYqNVUHLPEyJA8zIDvBtUHwgxPZzY
3YJ4P11j56s7I7YBLl+yqqPnOzZVXYTAOc8LdU52LHEtue0NIMieJUFRbiLd4iZL
BkFT7DK31vrKvrebeF6WU/tw55A2kEhR94uBTo5gsG0/D3GK2wf0ufrzwrPBRNMP
bUO64Q3/oBdU8ra6tFzidgJK/TddeIMNfIPN8NbfAlkhkobpcaAIjdbx1phQCrrC
ts1v72vzMv+hU/Lt7k453SqB9rmJPjIUOS4yPnJYa6JTx0kvhteqBD/WdgEptV5I
SbHIAI/Xw1xCpV9inf/hxm+VEXwGTPBpcc9o9eRCEQYxhfRQt24/ZBReUtxpL8mv
HJzKE4nK++vUckIFZtEVoCGmp43MKaO4bG1tfLIHXCG9t0Hr5lSLKUz/J5BjL/4Z
0lM6VPrOWF3P1Ktq6gPDH0COFWb2W4m0JIl/tBFPyhNTeGh0ayjoizf6qBPpKMPk
fpJxAyEYVPAtMMBmPJr8xwJxNbHal/rC3peGaNIpNADytn5PzV9f1Umu3xpHR5e2
DGq15xjR8xjUWQKaX5AjgMWtvPq4vYE9W+En0Xv5v+IBrot8mP9azQXlbB2Ce/iE
XwyA54FhwaK1xQXrMM5iA6pXM99QkXmmvIu3+KOJ0Dgn62koMdWY8MR1SJLa2lAZ
ZjI3BQhlUDuaM5U2lJ4ftlC+l/vHGW81Nfsc6vGi3/oPoSNIo9wVlClpFmuEXUtP
SEYoYRMrYDgWA1cMAVfidMlqawZbJMGPsFq6/xSzN1QC4twwqRfpILKLs06GsFid
qaIuGKoKIVKfJiEBaFxzdDPGVdplJ3cMNBC2iXG1NC2STTxwH7oKr++a72Z9HWfK
j1trrplsAF2riEAoXsdqdsgzWntFyudBTkqnJ/R5+gOHCKk5Y7v25e+NDMqeBSZo
LJ31879laWwjNdcwMM0c8jLDi4fLb42X2VEC/HEM+1JaImDDzu5Zv+WZY6xrd17P
0TAhNN2Cg5WeKH3ccZstJvqj3rJe6UiO9Rw937EEvQTWx5JlFtAHB2tvfzoXpYfx
4KlQlUfedCnJXU82y2DbM10hV5+AFXmL66Ns5pPaSTcOrrTyUVmSEW9FlJVDh/Kz
8+KtlaOhy0+iZzSfSQbsTzBhKuK2VdrAxojC3U3Ww0JDdvFPE8fjiv6jImfifEog
ECVBcFn8JTdhO1cSMbYbxsUL9zvjfOnniTPkiMCIU8mC+69R1qRLJEyLVZvvEaaj
Sb1OmtgR6SG2O3feyj+ecbyHlfuYrVcZoADpUOt2vjW6u3TxD2TQ5PJjf4mjRzqW
bjFesyytRjHpnaQQlsEePOGA9LuOsxTizY1YB65PL4PC1wIZv6WG6gN9iOEjdXoV
zDrkpG6tt01snTTWeBVz1+/ly+TUSWx62vUBuwGo1FyrafXuSF5yJDPNwZ9hYQa1
ZvIJsk0brdSk8xv3zmxGyjsHGlV4VpHFBATVswJZwginoPUVLl/kIwK5AR8gbejk
05tQGKENATgWeJguMsr1rJrpPulpTutH6NebKcXrC6yD/cGgM2zEmZomfWbdXMyi
cUMsPl/jQaa4Wm3XtBc7GRrraUO24t8vFfdASPGVRUJfra9zdpcWDwW6VQV/KrOv
rNccBdwHozlPPMADA5/1sksUGAH0elf7jLmK4L+wcsbT/qvG+6NkZQdKtcvvCQNC
djaFbOaTRGkPHjfXdGT6EZEBUk1w+n/QlX8ynwTwmQlbim8kg9XYQHcsLahWYaMg
8fxg4u3gMoS30Wd+4KcPclmChpzi9SUWe4OZeUYiNhmOFr/LeWo8Pz92Smk4Yy7q
0G668NePMHVzVhx0v1JqDzV1UIfGVSJzMvTupbmME05LwO3xNAZhON8rmcMLRBD7
GIZBQo7qk3vaUqa2SqW5JwyNbjzyRA7K4X+I6M5ZdwaOVBiANidQZMiatTLaDFo7
O+mCk/LwXkhYqvw4kKxK+KIR0yTHlp+WhvhA9x43MuQkG93u7oNJsIHBSsdT1he4
TtDnn+EnGv4CzNzabDhtu+kAtb352BrJ+VerGSnbuxIYJcOZ4kSkILM7LUMaLTH6
olYXm88wQ8Xi3oQtCb5MYdxU76pvGmLKwJ0CepvNinfLlkEr+8KbNoXF9TZcOnKb
lvr5MjliYOwb+GnT6N7zm1uiVvMFrhC5bepJ1SzlViWxEL9pXEuVoAYMCdR5PUuC
xP6ChuKJ/Zifm9uEsF28V6ivvByN8BnlUv3/kbTYctUXtHV106C3LXRNabFkFvfv
v6bjzCCvIwKB89XpYTYQ8nVrbtP00543fNzrG/hkUUKVFc0Hrdy8hwE3TSG+5WBL
axVwYlxv+k1AArwoptE0FBK60ZfHENjYV8y4/vMEbAdEtkVadGMJYx/lj0F0XhD9
anscJqSqk/06Cw+eA42R46SnUArtX6xL7avnR+EGJPvN6UnRGEGJJ+kwZX/8/ttF
OsAyLFypVx+WnO/ITuDajU11RKnJKtfkRVftjuBny0KdT0vC26aNQemzhCZa/yvS
FZkWaEA9tb19wvoSm/gfY1Z72gR9OXzX5xL1i563rk62ys/WEI4Cp0ljSCsFuuqw
7Byz2MV0YZWGbuJshjlXM1YFsrzBN18uSKfWw/LZ22w6lQkcWpLKRGBli/cgPAqO
g+ChyEqG8ZHPr4oaguga1xwgEvhG3Ybpk4+dLVcuHSYB8/yEwgwrZLJhppe+g3yO
5JKY8bfefNLLkSU+dwM4mOxTbYsBrfgd8Bm2E8rQG2r3vxXHTJe95AFQD20Vzogv
77A/a+hg5FTiZTaOM8kEIRU+2QUGfZxQV3cRAdtvYV1Tb4FrUEuuaJxLnq+/b1j5
/4GY1/wN0o3HEWEBMy/s18q6Ca7GflkzHFewQqO8aYeFx8vjafVQ0deldYhTMkSQ
wvBxVGBCtz+EWAeCgl7hSUeWwaWuIR2VLZKZ+q3gAu+UktZIBanCHLW/dNTU6KXr
c+fhwxasIzLNshN4dm37zWlhhePjlH/JN6Yr8Mt4PocCLOfjFIqY8XtkgnbQ7T8y
a0mJyOyzgf/3GZFJRSWFyveZoAopA5Ki2N0W+HyTuhgWiFbP4jirZTSDyjx0ZyUu
Vl3tzvzanWJGfB1pXXXu98Lc/BzdVwGIpPy5A/T4ztCop9aZadbNecZIG5xf65iD
l0ayt3I6I4i4Z8FHnyM33W9gW4+cnja9Z71fHZUTX1axoVoBRG/x6IEuGBpe8QYF
0ZgWPc+6gcqrlUNp3tnStEZ1l9BroHKVgMAjrnkzc+hX/sY007XXddI8QNPvvKZC
hbaQ0TcLBCecTAeP8SUPuq2grWSn761vbGy9ram00Km9/hfNCd7yTjXwW4PpN1+b
xq0jNYsS67x48c6xesR/iF11VKRXWByxtC+C1u+vDqoGix2O6mKMfEmqUHQOanNk
nFiUIrknwj4rvlWH6Q+rjj/HErEwkB94uu2R701bANVhzWPTnKoSsLk8fP5wBSZ4
+xtHkmQj3YwC+ttKmVG9aDTnRhVlCNWJEGt3P/aPqgCqy+kB+zsqMYs5nNhO37f0
Os2RB8l4ATM3lo5AWecVKpX5n1mmhK5x/ov5U3KSqg8Zojj93PfHBUBBwF6lxbPB
BwdztGVH3OeEsf5IRZFdBCcBV5QTs0r9fYIdl1TXHTgXf8uEs13+6BXAu8gfK876
bEhfBjaE5OiYvPEvg2Z+EAayULFMOIm8QY98VcCh024g6xpAb5Wrcbm3gG3KCATV
AKqlEV5aBJfSppIJTI7B7zKEZNW9qk9eSKVleO54RjEop//iq6FDV1vCAX7K8Z3X
4d+5/t3NFwL6n9sgsRIOWEXkcoFWUxJvCbLMnWWOs+TDbl5qVgy01E8MfLsOcn3X
gSL+rgBpiJB3fXgGeaX2yXc0ktVictJ1kuqkOH2IzNUgSTE88j0f8sspqwjhOeWJ
RLqzdnoQQpDXtiPMJ9yzwxDF8PZuoXqCmIDnaj9EAhpaC1lKjI12C7QMTRoEUS56
S3Si5AcQz0JA4l0y2ZpaQN/phQamt58RtXCegkrSl8NQwMmYu/yjqlSqH5cS9KBg
QhHs3FU5ex19TRMoNM1bswn+dwNjjTStN8a/WrHee7dn4BrID8mO9WKkv8RsgPhP
uaRBFCHCH1S+GmwtM0rcirGgNuF5AKF/nUkHDhHm8xiELupjf7ffaAhsYwVUhW+d
HKjIK8MEX59FhCr2mxqh6w0O4UJA3RtbRWbEzEP0dh+XWDjkATjHQApnerTXnZRv
rn+oZPrsT9zXDVPNTUAViX7mN5fno3SP3+HPZ4ubXyoIGatCCG3AFrTwuw8kto0k
LbBSX6ZLo4f6BJ4n57UZ1257IiA7ryu7tM23eL/aUeIVJ6vrRzmVDMC+H3y8bH49
15vfYqojhB3uiPAM30XVl/tYostTieta1Bldu32NBQpM6GaC/mzYJiEI6x8/0SEH
OVrwuQVs1z+LM9cigaRlrcHDU/tvrla4q6ud1qYrJi7EzQHHXhs8b1L8iKVqt4lR
saJR0sUpVmSTJrXf1P6KGR/41Vpp+/86tW7y+T2zNt2aYvUbxmm0V4W3mfn6yXFO
7/1Z1jW8anvGX/2mrMtIW9OgpdQCBDSrU9NaoUlxzTYv1d1VXjFql9+XL3/TDfAy
0i9urRyA/yaK5lseMrjA3XWWAcbU0d4dBe6irHKdqWv3XmT2nooQGjMSApSyN1d9
BGhfkc4ViT1S36mxPM6kkkfxGfe/exV8XETTTPtc0EacZGFCJ72glp9Lugqjmu4+
2lkccOibAIpp8zopZdRVfZLyoSeYl4WIyaTynrPufuwbXv7Bj4eY3nN8sBpVBTyY
0ZdDCoa1iKDvET8DHXHBrvuNbzDTf6apv7I6BZzeZS7pUN/JrM565pPYZ6h8znIl
iOFVkAhupTlzrkeJ63t0k3Lh8XFAPvmjP+MaCQhhwXqJ78BXIlzgx6n4KjiBubX7
c0Ug8TGcOh+cFtDN2wTwcwGm0+F5Cn/TVVS/vvTeXiGZkqOhPm9niR/Wct7uYZ55
jX+7ymOSTABE/nnRyFlvCOpC4dr8gXvuLmASg648ygnchgKDbClzUh4YAz9N9Ety
zmEDM9Rjc3/BF7n2D0wWDyr2dO4FjrC/tfxF+jn0naTrsFnKi3gWGPiNgTWAjwBm
Tyf5w6Y5Txk0cvpazZpl01tqT3csF9mjqvF1PExse2OOD+bxooJ6Q4OTLKIzxvbr
weF/fnO6+nWWIM8VjXl0tW0bOsakVKOLWmpntlS6z5U1cIgKP06gZ1KFIFGluQSd
leq+dXFqbxJ4vkj60Ovp3r8fdTfUPTgTT+IAg6elhtU4vyq/PttoEZwGRxdjLfmA
SuohbdEy8BZqpr5FIAChYuq4dR/h8udjQUFWuWvrxCdrxASzOPGzvIx5rgJaho+V
4LdTWBCGIAPiYtqToGFtzzirf7UY3dQAvg02BF+22raSxH+7gVOf6kNpXNzljZBV
wlbp8wTmGKRdceqLcO01CkMxmTF9aXoYeencWOYTEUWUK6I1bJJJ5bkc++/4fone
XoQijoe8J5kQ0m3y/Q6JAECOCZKgKFZx8K+P/jaApz7Li82fto+2Ks0CxU2nNTns
z41SH1d1DtVul3Z+yhc/za9oYgY9bxSYMectYY85250tWLY0eK6gPXFq3kOOKdVV
p/gYY0mLkMuFog7CMeRpM3fIv5jOGV90o+BZ2b86fy+4bSwdXGNrzkgqlzV5fnCH
iJEkek6L9/C0kDty8cG+qC1uSLSPxG/k7bKBrQPAyv8JEF3QPR29xq0UiqgUY2D4
UhBAzoSfFuv0H1OYfom7doo8C4eYuFfFpDGvHFZD4rkqUMD06ABfspfAceYRrZUD
lOl+Sx7r4LtFnEgVY5DhkrV2GriBMEyE32GHqxkp/5QM1Fw/QBqIychNfyyDpo2N
9z7PPAc40NXqNbMwTxyrDGCSN2b7+8Vg+E+YgiDL1yOQxDhZ4InNb5PQzVmN6nF7
Bu9/Uu4drEL5Eb6RYTtZylq7x92bO2xwf+MxbiP7cT3coBgQ1AArsjice/MwZIpG
ofEnVWrAT4eYZcmE93jY7ZXKo6WKG4+B/NzaEEkNk7vcLkk8r4cskpKFDmGBeBiS
ZEWQrG0MuwfuY7H3zbH5YNxs5a0jhESurKNURdh85qDG7mJU8NNv29rYymDFSlOR
xnAjbWGmgBwbpxlyKsjPOb5bHoR6Jws0qxx7wK35SNk7fRCgR2GUz3PK0vLeo4xy
pmTFpwbLAF9NnqTkTnvXo1hewFKoB5cQg/McSVUOs9LNyPhwpa58QME3AxV+DeS1
K5ttCu9CFjZz6D4bQDmGUAHJoj3TLo29PckapbQ3pldapTW9fzPZjkpZ2ev8qwIE
ceclno48BbsxnYX0u8y9wn3KaOfyYjK3Wz7gUtENPTClVg43Z7nviwWoglTRoREe
vMJXUyUXrnD4WxTmZn7HgF5fIJPDwPjroBgENlkpPK7/64YuWLzabPZRazKioMlq
sfkHXICjq4obgbesCAK1axqWRvp7aa7iHQy1OxP0YRL/oGVKnsE64VNPWC9tQvCm
pzrXAyM9CrlfI9Twvs5y7SAInjuhVX8zf96uYfrzhqxOSJSlPgQeDjou1y8ofOuB
O0QyI8qFYp8qIdG/ffzBcRox0TF6ePrtmAkd8YQdgDN52tZUVQxk9sSOtj0N9AIn
ZytxUyMMpSDLw9eeq3GejtL39/2FUFtbnMhxIbvGNBk4xLh39LiWeYheszl3r4KB
hA1ExaLXjd/q/+voS+hJJUCfNm/RQ03ebVPTaY4dEn9On99SY+JDu/nInx1NrxtA
7jzkEExktFBa+aGntjMfpXbc0rd/gHj7UvzrT4xEm8aBbxhX00YYg8juezEU+kTz
rf5Lhm2nrjDYXtiVTBfUZj4rY0Wq8i3ctQNRx7hWmBHevKxjGGsCvuTbZrRIVuiH
pAXIs+XiwZJ2/UNNUOlGwLlnEFR712MCZMoZpAV9pDiNvj0Db/3CXOibFCQLK+xg
F+xp43zLweRNc/9AX/D+dUOelM0A1ftMQ5qw9lmofemJIvRBY91AXnLyBPD/iFnq
LbpESeUJSvsiDEhrXjbIV9wmBYdn0L69M3CmLbKZ+DFRtlkMNZCysRWOaB3zhTae
37O4ivFKYFwyXvqZeFXRsl5GM+sNZQTF5YAVQ4l7ROQGAlhhQpI0XtNYHXAosrR8
CuEtkIF+QJSpz2th8lEmdIkP1A2y4CjrEy64EiIGusYtdsyA5OGxqmXUdCGuy0oD
OI1VeQ0fZaFIw/sg/+GiensxMPmJw0PFnHxNsfbuyzKLlgt3dJa3Zk8PpdFFXSoe
ZNbHpByznoFzLo/HTKOpdj3hp2znFjQFn47xnYmWOrlJkY5rX2oKewlAgd8i14RA
LszOoM84s5vLDZ/aJEnWeiL0FZfBlytHIOC7mBw6pi5RpmvRplQg4Gw9A5/FROnR
+VJtklGMoyidDCv6lZQN5de3GvNFZpDBI3qcU2cUfq9ER3K5o6aYQwKT1aTkfA64
LXYgOh2YQEBcSDwSSiiFfVb6atU96iq3P1HXGyLD8aD6zlgaZaFRDigjfxMc1A7w
Z14vhB7fOGldJeXSssWOmSiJPmeyBfxa3rMQ1TCtgj4Ikcil5YERyoFBnTzkigjN
WvkjSO9zxh9Qchc7TMf1coVzZs53bdzfhr2fMzcnIEvag6E6da7LniU+9toAmOI6
1GDgp/ZY5oQQ7X287XSfZRWd5w8JyU7PIkpx7OeOY22jksAzHK/xBpQRSpIn6JGv
w+gJ4Z3O6ksN9rIRYmAmAFtCQJAq1lBrjZAHYiX10XWUkyudcupJEkazaTxVosEH
HOxxQ3RncKf1hWtCUcLfIZB7VhYWHX7dljI2bh8DGVetzt1ZBbSt3hQZZ0ktdxw3
NMEKO7VARZlRd6Fy+rrDGUwBejKnu5ANV2pN5+XSnplypb78HtMkwqCbVVPg2BEA
KG1KIrrDCLAWZGXYUro73biX9aPeC3DpfWIU8BV7r9KaBIjNuF3zFLdAVOzZj+9K
waoMN67xNn0XK9/9ZVyJON376diXGB5eTtaAqEXzeJBikX7Ewl8+Cy9clYs7CLOl
EA5UcF7rEMaee7lgBmMwJM3T/Exl7OO6pDjukb1nJOp2Z+wDm9YRONDacNEZS+OJ
sPpp+19Rp2HrwbeohCc+sF0gAkhiEhl85v7nKs/2kWnl5UtPh55FE1iRcWZ3dXQp
Y3aiQktIAEhEgByn2b1KkkJjVc46qPcLrUQHrUqOkWy+Zzlmr2gDfRxcD9Mr5Ppp
0zu7G0Xa0qkbRMDl3VM+dZ8WuMKH3jtRx03OOyovqfPnPUljsd4Rp4e8t1DWAPFq
t4ZH29MFv1H3y8/8RqoRvlJWbwe/2lB+4EPUT19KhH6DV+J6CdSv5/Zc/KqOfUPE
hdVHnNuf9JqjO7f0Hw5PAGxQsVMtXH1Wwd17Axixn2CwWlmEVvpq1cgVloyJOlAj
FGpSpZyoChqpajA0NhjjkSTbjXsFqa5tMQpMiXpFRRQ8J1EvMs/fk7c8NH9vQ0FK
aRKZ892yLGEvCZscRsYVR88gFkX3lYKDB0Z3nYjpgIV+lWoS3+IOT9smLeGbLTjO
iT9MkO6JrrNgwI+0R3Yh0lF3LX2NquyDIpEurR7QHanGdj+ENtEz3280TIF0twEb
lpNbCrUIt1xHE2Ne/vaCwwul/nLf3Swyxhg0YZFuObb2sk1ke9kwMsHc7sj6duC3
n+hG3avBnXnMjTGUYZGoXZcZJa6u+rhBzvJyjxx8BNNhaoeazWoUhO+ct2T1KM/U
PY1FXIcx2QldW+gZNOknAs0Ifus2QitjQBJAqksxq3Ufq21IVEfuJgTz8Y+cZQsl
n+dHpoX3ef4Wwi2TkdHHek6PdYm3Qau15Ra/uR6oflPSXM3tm+lFd/L59xQHTN0d
bJJHYIUbgtFc/F+bKkdkyPbzZPzL5Vb4CL48cuVx4v63wiZbhBm5U4uTph0OSwMq
EZA2lYd2DGMSRaHPkNCh66dth0Fy1BwiO6LfyZUJHZaPjMljxd0scq0TlIOdQb1N
JU9AckZleTnwNhEb6gUNX3IquJCYEutIcCRPIJQTdKbxjEa3IdpKnxSyr/hsi81T
DAwAUn3eaxZMGew/e0JxQLc6W4TymPDmY9fwaRekWidWDkL4b/Iczrio2wHYHs84
GOZghn6zxRqLaxp8iLT/jXnBSBeyUhRMMTyQmD41OzuM97EV15L5OMP9Qli6u/Uc
12oUHrJcaxXAytJp7VwOS+3yDyTKHRrkPU75GRR+L1An4og9jhhhQeYh5LI+B6Xh
TDe57iQxkPLnEC8WrxecvAQx2e2/gjYMBeIDwzXRORqQPiMwChF9juYmEr6/ZC57
J4+Hq/iN4s+ysIgXozhgsTx8kuNWWhEZvbvDoJPoVUuYqCg3keXwR7l+DPFYyw6T
tC9MQBzXGIz3rRk3yKbRobC87tyyH55mACL3xxYpW85YeaxaC1CIoqVF5piLmvIY
godkQE2XJ3ny8HcP72/UHfBu4KUa+N9pU+0h+zYxMc5Xs5K1cOWLmHt/eb3lkXra
6K6U/CZOjp6283OdObLfYYJ7AuaVYxd2JlNkOszc/4LPFqPAuMxDgFz7hLcVgvHY
2eiEGnLWxR87ax+RBenJkxmIkZBwLkTaSc8bH79GiAyjovh/iw463q972NQ6UCiB
K0soE3v5cc3AilDuKX7fs8Duk59M9Vb+pvEhYtL02FVNZGcI3bV3l4TnXvMNbKrd
TUzys/zlt1tJIO4cABToOil7KS1T8wbHKJb6pQ5UX1DO0n2ZpY/U1jwfPBZ9L9cv
57kToFyT7XPliTeHfl7dAKoJoSP3VxJq/E3gjSOxs4lOLq4iLfuHiSA/HSCiEkfy
byjvE20cby08z5UL/uv6N+HTCn8uU9FjvtZJ1L0YEWNPHQxewpKz2TYURcRZnkmU
8+lW8YDg/SnQvPhyzxmegEGFJkOuScb4h04oTXYTyCOPtlCF71i3HWlrALOKsEKZ
20vRJqE5rNmEXgvrKuyZVpNxmA0eqxxMPOEbz19cnIQzcNGq8JK7Mg3mDAnIc4uP
+7tPGK8XrW7PjNt4zu//S0xn0rWxIQR7AONJE8BAab6Y3fqCaWNKyHLrEqJ24htL
IT+s7uzZQYLSl8AW27qtjJWTI5RvKzr5vH2tLRAv2mQ0YOUou0Z2xWntp8n+pTNt
7pyoZhRRFCQkTuphP3fu6jmMW4+W3SXQbTs1S4sbfIkndL41e0o5qEsxUs7i8G8c
NWe72DLUvBHLQk9rfHxrJg8DGyMKcxMusbrKTbR1D6Q0uK7ldRIpuKu/wO53nSYZ
sPJTDIOM1s9r8evtU74LHoVUmyTKGApQbR0vD8xCzQ7T6BGcL4HiyIS8429ApTn/
u94j+gH5/jTXau3PG/qNOIQFplFQINZg8LIhmmToWVRXBy3/xfyznXliJ6w1gHxs
XMiwuF8cIh0jS1jDnpgHLsSiHzl2BFUgLWvAhpxi+sWsj4BvNnPFhhgF9zZoInNy
bIPIFzWEXlUj7mcFZ8/0yFFhialtej9nbb4ijlxN57pmOduev+zQ8kQAjcip9GS5
+gNNk3lRT6hFyN/w9YVwRr2vxEMmuaq2Ds6EOujHRSGA+h0IBKFrScYT7fizniC/
zUQdAP28Hi5EPhQnNuTFpHbc2DStdRRSgxhZ1fKnzMMMD32U0O9zpFDtPIrp1U5u
t35ueRNolkV55zaWuwp+ksZz2kR+ge8AG/XVt4qZEZFwZfIDoQNpMB1gMBm4cEzv
nppk/N+3ou0NHWoP4G6kCBX2EZcuSaTLInNLW+q61GIDbalSO2qVWuzv1aLUqEYf
lWNYzMtUzpky82s5Pt9Pk+og4FHKVcdgpjJ2woRZ2VbkfH9OWzyg+Qqmy5AXpD5k
v8FZWo0iwjmjmLSAryhBwPtIzPzbutvuW0qdCY0Md29+rWLNQnz/2GMcz7nWt4NW
iToNkPGAdOEcvRkieVY2LKEWLued6DZMobWIu+Ug7mrTJvWT5fJJoNyAoxaoHEWW
PKfs9WljCBd8nOhKYnAXRUCOte1fi0Q3PsiUloQxSBe1FTwAZo+kMvS1REsEmWv3
qNOuwNsP5WZpfRqD/f74sYEwCArui46KJezznZGjS4py1Rczf3urgsLW1Nc9dBKG
m+jdQnGUoll1WhApZy2TXcxv7M3JGgnlaXUU7mjm/8Uywyq4j+RBefUrddlByNVU
rxttPUysX/HF/247tklSNIzaPgQzXxj5v6ACQgsTQY6HLM4mtg9Xzwt8tZZxm1Of
qO+DL8b+Eyy0S2HQFQVjJBch59z/wqVxNtxAUcGbBC+bKl/rUz+hw4h7kdhBIJDU
5TUK4cec2jJl0Fl+MJa5vVpqLNiQPlN4hSLLpgqMvFqiH5VLVu5YgRuRk98tFB1b
gY9X28NHXCNQ77xwNLAN77sLEhIMINA8tTd4EMssZtK+KPuLGKrcURZ8NCgtDc+X
gaAOXzkxf9CCPht4OGP+YLtfHnt/HGbsw7h9DzxOh7DzLGH9bhiMgAZSk4WgDN5a
Z/5xgMHjj6hDh2N1+gHOa2lj1qZ/Co9c9n0m9tmoBk0dgORafy1jg6pAgwGGLpbd
NNC60okv+IxC3iTfTToPZSBzp2gy5PoAf75pbqNdSs1uAT1svnqPdGJY1KGbfrNV
5WnShKwzyEBEvB+J7NBQiCib0g06qmke5Gg8/laABIEcIrrgIrCMsUDG/NyRTRJk
+l4ZUmBudiiKmYb+X2GUtxoQV7cUwPiIkVLhj+9LpHtRSibzLquhj2fdncn2VW9w
9NtnWPRHjUif1miEMF7r0RQPrOBuD39l3uIDn1Vwfb7eL0tCpWOd9Ykffa8iaCGH
8lNf3QjwtH0xqSgYgjHSLACGGoFx/UC5qwcL1wX4Cqy+eRFLS9sIEu5wZnKcKDrK
mrLg0RhEU/KZIfV+eyreuIvjmief+qjTHg3PnXy3ZWeKRGLSYQNzHr+jIXP2gnGE
e13GSEoEen2KS+nj9p0wXpdRONYU9ghWe1/nRiPF2Mdv6llDS5+mod9iX+5yDwOh
W1EERsiEZvshZHskVdxAJ6gXteBG9rUwHZ1lqYlO7jLIRVbgq1/na0Kx76SfXQDr
ALM72Em0QVNsYi+QQaOeI3yVseoP9E5z2WM2OfosWRkmIVA+wSDgCFDNc9/A8h3w
kwWebGkP7KSpvhksmRVdqI55YPL5LVsA6rbGPaF1U4Vj9Db+jTqZwH0txBzP70Bk
o07gwJ0g+hDdKKprA1SAgcUwAbNjsuBxUBQbEOEbypTNixhQ/fKASqyIcm7TaAOu
yqn6t3qqP/aafivEMiWsI8P0RdjixLz1cCxH6F5HZv/L3TpW0exOd9SG9nfLdvv+
XfShHhO52jnvUra59kHf6Xf+HLn/CtcQADe7LHqjInC5DdgxasY9LFHktWhw7E0z
ynYDMEnLazvVESUGrYVlm8dpmmIH6MiM3O/SnHdJzNBWqX5N/YOu6gya3usQ89dk
AOKhvDQAyTQq/5ePGVJR4gOzBY7EEjGSX0TUFXbRMy/TeoVT9OdRnnLaFF3J7QzV
qtb3yw35NWdc8agbimlhC59AhQ1lxq58VnGUmX9Gdf3L9ncSlwRZBWHbWVkYUWQZ
hFfzPoK8vEGitfIB6+kOgRs1Xv6Uugve0WdoHgNZpk+XiUAEQnEFXSaiMlVZinsS
1L4O/XtyfwfXu/ZSn75xfFhKHkEuXvuGkM1Bf7XAZ7AaWGhoSxraL/G1OprEh/sR
TWz3t5Voih3+Svfs1OjBF5mj80uwImLKJmJQEEoiYfCMzhb4xlzQm6Zw9yArFOD5
C6tC6Z/eHxLkp3OPruRfF8ifpuwcB9xrcm7PJlLRwKm2ToG4mvMZAtIku59lJ1yG
AVZ4hmT5PvsYcQO79qpwsx7b0HHWoeldgQTNBq+QvoJ99xixHCZJDBWRf3yK+zLS
iDJZ4jGBVofR4S2jvRcFY7uMvtJWK9FJ+LoykBSlsDDz4mi0MfnoQfoFZ++reEIn
qTu3vfrZU5gbLQNMHwoQc58/8s4GIW+yGYr/Ht+0BLt+ZQ3m95Mk7fEyZWBcla5G
kKCjRTVqyNENFvDsQmYicfUOOzDWh1iG7hzgxcLLSmzv9zjhGo2ljTCEEU1RGXr/
Q/GNPgU3JIanHEIDjJM3IkOpLEkSixSkMeWmW8/t6Z6+EnU0nVduGTgx3F/0Evg1
lvO3jiOnYen8x6JzifmyqxXCxAlLjYcwdyoH9zZ9/S1YXpNjVbfuJro/omNwTul2
dq4zZoI6rLBG9U9GcaTpfmrEWHbGNk+3XdzS2TD7gqfzkQ7gix1jTI+A4vWsAOXc
E710cr6oxN3XADqABdxVhzvStCnEISjTssra2F2remvDsyGfBQiprS6++I8nlurw
RX69gn2Ij3VOGncwpPNbBjauvlp2aOZxig8882rouc7oALiZ5uLQhzKOZa5kytoJ
ug9QY0urGXilrAuYRdpiuDBjonD25jy+q3+L1bdNYU3gZM0PgLsLOOAFxYpBX0RX
5sro0c7CH/jh/5xLlmsSpw24eOqp3/OJY98FUjEXCauVfXYAzaBD8vUvrx+yHf4x
nyGjxu7QdYDdrggXv2wtgixri315BFanwWNijp0hDOZML0Zw74aP8IpC/tNV6QEF
nLJxWRUiAHQ9C0Hzo67nT7Vs3a5wS8AJkJ9p6P1RQmeNPhDfihMOEI2YnGH4LWYI
fB/bK++ZBqQgLwjbPkTdf2o9mPbT6Rmb6v2SaRNgX0EiUVB1fClkIF8+9DGD7qYe
xdGyC3qROEtK7n/Lv7S3lLaqBXJkHQRLKSZDMNlP4cIHK7w9+i548Org+Sdy1Jh2
clXy4hhgSfP7j0ZVJ3aK7ASlq7cmJkZuJ2khX9NTkxyM/OsWeDn716cVT8m4AycP
sIYnHsCeOxoOm616ssf9sF+C14Ymd+vcx9BTHsKpV8ULXm5iMuCbKPACv4D5kHlY
/6ijsOVWknHbj+uJAF1ehA894Iyrz8HpY0WCYLO3ub1X4lwJMceNKGw5VOeDRomN
bzAoHpMkWWCv/dwUpXdBvMONX3ZzHGu45EMaYQiZK5FCXZKlPU7R1OXQlGBZjDxc
e6urjWqfubKJ5UThO8BTBPQez62agRLzA6MkHdrfTNrWrMn58C6N+5Mqgc3D5w/x
54Lpur0tTZqUewc/GZc/PtHT5wydOsgxAjQ0DEoBpAJ+DOX4p4iOz9cr4xuC6YJl
1Rvo+Lo9okMADvt+SdHeqAXn7GdTh5vmD79b3kkwFt4wZrwe+kXBsik3VAOlIwTS
JRhVo8RW3G/r3cQhemg6xWLwc+Da7ZK2r1xY6kfnB2xMxVMZl1+oWJvHLKyhhu1V
LpMPjk0Q0yhWI6eVOC413etl47l0kTGPlfTsRl5A0ZfgtwO4bbNXVZUM8SZ6EHSR
D6vhGWe+hLNOjS5UL1ZJQCIfzaqLstfDak9uJFWbd9NoF4erboOxnsKXcccpATeB
6eUOZx3sm8cjV8b6m2nM6imDhwnDwbaYFFd6hvRGmKEihW63EiPvpJFGP8QWTQ8t
ztN+OzxB4Cr/VKj1q9dcnkUZ0G45VCsRggaU6imVq48JFUhH6uCjnepkYxvJAfdy
sWo5OlkCQ1CBt3O1RMelnHNAlmb+mXz4CGWpsLhXY80Q07otT20sZyafmi8E2fOj
/YbQK+BgNtDIKcCHAuQ1ZcqTN6QttUduJvDD2SiAVH9v1mnQRqrRuqrHnjmRvyYc
F6LUgR4LJfQc8cu8ZxIs9OeM0Cb+O8/VphX+bVIkWQhcUaqlRFvPZSPbc8VL4d5i
O6kM+XJrTjTqTvn7vVsIdvfFj8rgwxAcV1i8p83O/bVUG6IG8nEHQvBHquYv79oc
YBLPYPr1nrc6c6k/vA9Z/u9NJEZzHdi2oDMugcgsy1W+N3LBS0cJRJr/R8CcrT+p
e+QsFtYoqMW7G2X89o3YDLKxSsSFv7Lr3AbHXtV1uvhk+f3KGxaeShy/0C/EpCmE
dpmM+q9DYV3CgQqzNWdOch6DUnra85Oq2APHyuz5gK8bFFZau3PbpRhdqScgvq8A
xRNzyzmSjpPmd+0l+aWJI4VGyETKot3JR00x3fjXu6xXruYreWUkBLjgfIgizp8B
ZVhu8ngMVDsxX1O75aJNVzn9b65gPDBxPeQF6LvivIFNpqj1tj4ELyYgzDSayDTP
ubFyolnDW91E3+U/sGLocc/Qhsf+1LExa9xO0PSFp/HP6stMF/3EuprpCA4GxVAU
FVnAhqEl226cJuAH6N5sqUNyh74lJySsYVZv/mI0ryXvVyDM6uIf5bcKhvsjUyIG
otQUbqqTTOcp42rvCnctI4Ucy98kjk2hsG0g9K/ApmPjS3lYntVsqRLfNjh4Oa2h
HCZe3p7tJx8CAbXK0LQgScrIzKz8hxmeyhClrCi6OmLbPVVhjggFCytqpmf2xG7k
F56sw8WaY0jvIfsD5GJb5zR+r3UIcFbTymK9HyKeMX/VxO+tuW9vljJSTfUFidce
U1+PTwxkhmhVMZ4b4uw9LMik/D9XDerrNlQGJVYKupXAB4m5sifURXtiI2gcJLIG
pwOnHQjOgye2sUEn0UlTHGk0Q4GOAd5INFEzgJ8O6u3KA0SBuANPEWwT+vDMOX/Y
4dVH/2PIApy/5+QJULDPRFl3QeD2JNnvdSoDjl0ZYvGtZGYEePghNn3UwZXojJk9
7iTpqWxxvX/o0z9exRBF+GK/JYNBp7zG6cylGPqUMeGQkIca7dyXEBly+MDEZGWE
Ti8O4ETtapvmlYn3FkdFf4j6a/R2abcqiACFsC1vXPiLtOWvG2IwqGka1VdyUV8L
3fHWAYI5xzWN++ppf9XTcnslYyG89oOo1CFzzKKL4oFFwoy59u16lnkV0Zeqor6r
jVkDsYRdx+JL3nWa4gqErNxyjmR3ik07AbsAkBXVSb1qRzDr9iGhg1JxsjjW2XRM
WBR6q+ENbg3/N3nSTr96Nj3/sgr+ZI/BkVmP6NvSDongGRDxKA/MWy0ohlld5Ale
XizwzRQfyKev2WuUyvlsAqMAkv/IWznNpjq0FZHyJSvXBIix6GAB37Eq3ry6Z/ty
aUr6eNayPfBGDJ/Xb9J4sUVYgWZaJQ9qrH7bYAzUaOeHUigAOnl6ijLcVMfS4ZLf
XbqJTLY75KtN8YEtcOCmZrMbLUX+lYQB+/nIUqPq29nlr5bBdgg9JJHqDL5FoJpV
2PNNyGozs0mMZhWVmMGX1nbc4TEr+DbRS1L3gbj6BGa5WlvBSIhPQeCf89aL0V0V
Bu/BGku1N3uhYcWvO0pEwmuxt/zGq6s3TkACEual/J6EHEdsLNs+1opVEL6sMWug
kdomZwSvpm85nt2EHk/5z0QWcDOJyTk+UwdOjjafkK2D4MGYAvIuHo1P4W1NBSRV
j5QR3q40K6rjypCOELbDqgUBTEJmavZ9fR2H0/EznnNUzaoKIbGk4fW235dNsbUi
HocPr7OdKfcTuec3Ub1qXANbAGT/S4pjcbYizDtJV7+LfQHAxQl5teWBnD+Mpyk9
wMEKiS190i5j+a77It6c2Tmx7ymZuzkI/02WBVfHeJ/aQvlKasrLZHKSVJaqIn1o
E8lB/e7fvM1YckEeCA7TelvTvl/w9+MT0/CtSSodFIwV3Ho3GzNt2g3RlsN6FsZd
mIzJjG45UAe8LqH2IJgjtn1vy723N1SZGwUx/TKH08RHvFkvRIx9C+P7IFeVGlD9
VxpopsQe0MeniHRRoghWpXKepLVHDD/p6GDD/NRMTh8he7n4utSOI0rjwFD3XqQ6
MIYCt64C9nDv+IGe4j34joynBLocdtXt04EV9BPG9WrXAzHogKeYh7vXp3B1sNz1
4RUF0yiN4BbQJoaRdm4MD8ZhbyygWjoPs8P5kqeH/e/GoQuqJ3+kZuLUa//YdSIE
3ANYuRnjg26U8JegIBd0OZLTkNWoVEoqx6i3GkISzTqiozgXCbnTDwFx44yPf1Px
G3dheRI+uexJScsiDBBvW+MP6T9D2Xo+3A3pu0Cs/3UEyMaG+YTMmDrrWygOMZH9
j9DYmoHgPBeMBSmKnKl6o/0BqCJNjBtMLIigPmMtra2JkMtiFx8jv1CmqGgsf3vC
KUe7z9hwAXUCyuevogmLf3x/MoVwNaY/zeCI9Uu69zIf+cPM4IQxNdAnXdKVdXRr
zxxD4XEOlewiZphB2wcwoA+pAK/HNvO58CmQkn6VKypHlRfZsfVVNqzR4cbKhT+M
PNYR0i4iW2Ps9xAmk7yorxe7565kRL+skNG2UzfWUVb/OfkQenX9eYa8GerT7gf6
rFqE81iI9WkUwot9yUfgiN1hf5f87ZsGeGgLdjgVedHR6vVbNS1PB15It4ZwWTgr
0dOaJSNeBLgV7s3AgNE0k4WFzxtu6th3WkxxQ1+JxtBoWhSH80f8bI2HaVKr33ek
t2jNKj/69mjWm3a1AsC5FX099MwaMJsH+SQAkhrGrMD0B2qSNQ01s1tbCAkkE+8P
lO6S1kh7+s+sWBRsvPddrnPckFuRuLGqGreH3vqNd/eH8Zv1X2QUgxGtBpQLcjVc
W8iJM5tRnZgtTkjMCoYV0rszKHjv3Roa1p2l13tRyz43n+nzxTta3WHSa4eFQY6r
Zm4ahDmak7BfMWbUiYYBxvA9M4VUon5GXTparyVEhVFSamQthVESpqh8dTJV6Y2A
2JIVrrdaWw836exsLVUvNEEM3AsZyoESE4qXy7V5ydoT1YMOxoX6r6LX1rxvsLC+
NgBt8mFjgEjo+04Z6wXmwnuaP7nXlpQVb/darRALcZws5f+3zr5vCi3YW5JN1YHL
IjvdxllBe/RW/tGUsOXANUnsJtXYL57HMNYXgGbvF5PIyZp4sGgyaFQSzLOI+3gh
6D23OpF7+GOJFecOWsNB8Fl/bF3TVS0mMcQk7Ij8LKt8Lm9aSjnf1YjZiyHRV7kL
4Xe55Tm1qR1NZpnu2MXiGd5eMPFm/y2XBZ+5FJZw+Yses98A2wE45VPrf1WzXGcU
8jb0vzbWGOJFz5GhNd7+sdWdi8onOoxwf/fS1kt0eHtWBhSm5nbSn9bExmDrB5Zm
mPQMZPpgTBM1Vg71T8Bljt7agmYnO8SSGhJ9tsIYo27QyKYeSfdTgG1u/ELVLzkf
mGlsxnzPyNhAKRqWYlRwoXDgodC2gZ5IcBcTcjGq3aKCMLaYtQUJXF+g6fJjeaMp
UV1CPZTHE9Sx/4litL3ITGYxXXe02xHKJJKLK1svJSKOxpx2fv2S2bgjSSkRJBrN
7MqwmZ2eoTthungwR9Hu/z8XnHkqtGSzF6P7TMKRhWJciNuAOI6w1bTc4PiNHTeH
/pqFsI6RV6dzmRe1XWduju/r6pKvZPweGnn1yXHsKF6EWObxBFd6rbrJcQTlCqeI
chgoE0Dz83NsJ+K8M2I4p0LynjFei7QrW+dwhoyAG+S6xTRIrbxYR6bqYaoXXx/a
yngzpG9fyRYxclGa2ysGJhAzwdhBGopHR4l0By+lkHiKcNyhcBjHbzlgUpO0+aIG
TeNJvY07c/WcdwhAI+abIPfPQHtLB7URoAkkEMQdF7Zhj0HuybrwlF5SXHmz9gVy
cVgJAD1wKq95S3zIFfExxCqpuWMLLqMnMnJ7NtKLw0Ltt73ZN6qiuOOyoGD8IqgL
cW8gY27lDZ60a8jB0CY4wYZgChHC0yVxzC/AUomoEISI9BaOBgaG0RrCnU39HgkK
hdSAHLpse0ILfIyx5xEK7nINrRZrxSz2P/aLi0NWs18CehPT3XEdcWF6eAHEDIxV
ayeq6E29szZNC312CjV9W/aCVC4LPgHbQTbAQpvUoPxpYRwGK2FvNLeH5dyhvxqI
JRhGJ02JZmahp8AdoNxTmNZuTUQ8mGRplIxrmN/psJS9LD7lu6IxWnXgdYclY/pm
BC8UJSuykJnCvRmGT40x5O/vegwf20oi3grrKFPxeZPjEjFt7QEL5mYe5w55rwcw
VYxg3gHU2BNLXF6fnSEU/h20AxPYOFgoKLtzkQqmjGy2UiGkKFYsD5oTlSa1QfW9
O49rmEYg5N5DtRL3K/4HzhekAz0e1xkHCCc+2mE36W68YBV72/xvM6ebseBAkZ31
SDhPuW9LaS55sSX2J7hSmmP5HaY8mvkbY2nmo77H0ugBXgi2N68iUloCMnBWeB0F
bCx+Yf6yGhphHu2a45sBiL+kbI0g5gw2IAPjrh5vSmz/Q1NFBDBAH2VYHtqVfa6P
D8ExTnpz6erKsAmA8wWrfSYkVnfMkRRmB7zKCsvgQZGnvZOazBX2zYTsS3Yo5AA0
5SyOdT2GaNUePSNqdZk9mxtiVmjrzzITWWDrcuih8WI/qeqRTwtMs3qOkFqlSI2B
eMpYTVpqnMR21TAyk4Y3LnVyz3130lc80KPZs/dLihEOIs8yvQO5gcmEVAZa6Okf
snZ9fcQ9BaQvLSRIKEIxs1241k9HFn9voPsBYLXvOduU+5F1TbkMIJld+je0jeIp
9p9kjG/lhdwn2viJlAK42lM7778+wKO6yGdUaHpXKFQqr1WJNdiOpeDiL6P4E2Vf
cdSBGIY2PkvCeNelmwsYmbxqUiPQQ+e+K0A2NyXNMf5GZUH9R744Oi/noUqlcZYo
B2448KN8pjTR27Vs5ze7jQoxyj6ekeLEhEqSkT1wngbVJIWyXwz06hybVbp7/DwB
frOic12uVutlt1FWuRxVJmTj8ZW+AC7sIJvKY0tz9JBTF+mUvbRBTTwLyX+PmzcJ
f3kJMYbqU4ypkx78ImoZEY4xe/S3M595oSsQFujrxvSrnxJIa8D+n1bdpOpGh1r1
X6SiWb4INyuhby174s0+y16Lo3hFnOWta2iJL6BxVjZSSAhW8Mv1ywXiQjnkwuWz
chPWbVCMutf5Q+isQNlRg9n9dQm/aBTwjW2Yn/83PCkUISLIevlFaMu//er9xkas
ykFEjxzXgP6J5KSV1mbl27Rvmol+bMkYxZDvEI22tHFAubN7lx0080WnpTfDBnFE
ijQo0Ptpr4CC6ZyHdGOecDgvs/Y/nlVwC9QmmRbtlRrdmGKv3RpfIz7pTOypaXpm
7sDs4hZFD47f7gLgUSGDQfMXyhp/nZhVhY58JlYZO10rO4yXflaqT44HRvYcp081
wJkfApDNYzE60geoCuENMqxD52Jx3Z5BWiRAL4ZmkvQiLXzFQN2Zug4zRMTjeyDr
tibK8Rl+X7l6mZifUbYnOIwtpyAytSTOMnqhU7llW8hMo5i6NkEsMT8TF1d3zxoF
2gxXNTZuOmJZeBSFAqMsnTl6h1o8M/xPqIQBRPvX3p3WlW3CutKoyMUXsV8GM2La
eDmwp6Hss3KkG/bhZi/Yd0JePZo1ATKudA4PYGGuI4cvy73JfTvNyWum//EsSD5D
nmc928CRhZRAttjneW9c+wManPd3JcCRCcWJwDv+2TkeOdfZ0A2Y3sUMvlAmA1pi
2Ym2CC05BJns7E2qqcj1Vl0z1xAcNdMTSao5RYS0+1z2g7Y4iigvy/T9+C7tfpyF
URa69Pm4IvJs5WJkc/oG/LpxuSAEqamDIJlqF9VpAZWmu6dDhYJrt3iA3KVQKvCT
T2vQ9pyj3bxdwZLzzITmW3pZCB+MthpetdiQvphkCnP92czqnfrgq4X+OWEUEpiq
5N6QOz5BLe8AxiSyduBi+v8Y3BEA7c8+wKJAH9I6vtC+TNKsU8L41gusQ/Ys7knJ
HLLwe4ZsZAhh6eUikgfwWL2pFCLWKgP0CqAF9DaobM9A5WzaotvjznwVX6JH5ILr
KsoIq/vc6CjBovYoEK9qNWiiydHMCqzWw+APVmOp7eA1FILX/Ngf+fthd2uGZuIc
KGW6sWxKOEOfP/+XNN3DvtmHb1X23cWNX2kxJw3BMiicsP887I0UQ7PyWPrj/Sdj
fK93kz/duYMCm0lZ6v4F5gK/vj7PV+k60BZdgHa9Sjm1PLqZtPkc70f/pZEsBwsf
J7aRm6fCPBI0N3WXgc8tMawtL8V0IG6utT5dgRasSYVDgh8cDd9xbBTqVq9Mx/MW
i1y/do1zYpG6X3ouNw6JmTCZHGQMUkUymBAP9TzwlbPRYJXcMyUgXA7ydUkxwPMT
/LSCLuATs2dLB+Jard9CDNfP+mS/waklgxHzX/Yzrlpy3W95fbD0StkXoZx9aKjd
eJQo1YaqvRbwEYEWQjjDHMSVammHWn606J4vF6TQiElWPPjZn2IpwuV+8Tl/iDzH
yaX1QP2I+mT7IcwNO6gPh0Zt+OxlBV9yZBzV8Qt+1lRO1CuFY1epe3WFtllo+ArL
RzrhKs2ImMFbIFea1vqMXPvmLZ+MND/lD/vwqVqJSxZQ+htHfkbp/2IRrItivPUw
Lp0XSIwgUwQgODSVZvXtSGasfKEgiOOkIfdCovvOoOdnarIb5TbtAHU2+73HHM3A
/ytnsbAykbWAcpOKwsB7PWPVXxdk0OrdEjfhCfr7wU7xgPJOURkGY1hghXAFCSlJ
VEm2IcK06K6NwDgI0yOtrEAzn++/6Tk08er1CbxmxUrkoofmgZTF+xAeUMeOIjoz
ijRt6L+bjCupmJ1BBH9ZJmr2t/RUOFs9y04yUWH810bcQeJwuoSubarX1AZKA9Xp
/fBBS/EWgU8KN7rAF97ItbwU896BoB+WTDlTzLtgF6By8sHKBtCLlv7CzF0TfVit
YC03TTTGjfBYGCGYBotxxPgZXbkKdwamM+kt5cI6FqCUWVk0wBmLjPBf8W9osOyl
CZBfVCV9Op6BS87LKWYWDtbT81L5QXBcWQuGOqz2xauMlU2CaJDllviG2sO0yk0W
Dkz9yexK/lJbIoXyZEyIdnfqWSbFSt/XcNZyDMCeum0qrjfdCzZsjX3KlI+LI+U3
+TJbTHj7WDbd79G1o8t9Rw9d9PDPtj1KSRZc3RQd3qj2djJ8ICkS/tI39zbcEUgl
pt8BRkIP7N2UKde5mBEHYk6HlEkz3l/EAk3G/Phyh7bsdiRdHpeSCXQuSFq2iTA9
V/op2akmWHRRMSaDN2goGLnNb0etAOIAeS0GtEgLIRAkw+Py3s7YBOPB9rbCjEBz
xoUIZ4EZyq466E3IwVMwNh2gDEZOGwRa3TEahtdEjaHFedTqx1Jm5BHGtASvStTW
5iB8LPLyZ+TgClgPSMCKjbUo+364RJlcXYUEoBnqGFe4YNYXO/WnkkwoRX1Q+lOr
yNvRbb9rpEl7jzpa9XwowsnEsRYzugdQVD0p+Cz4XDOYq7scwkvse20VNsJciDkW
SuzVsnCLfXVb7d5hqZkJ7bNqbzUwc+wRniNGX+kmGEMsCw/V9Tz3JYA+lHDy0VAv
jXGDO3ptY7bLhvBIUsZ/d+T59Jt5h923Xw1zAN6Y7qN/zKZkIdq3IGtmWjP+CS0R
eL1Y/bi5MdQIbl2Az1wu1jEzXMqPGfF3eh2gWutNNBl9mLvIMoJFHMD69vOf63v3
wJnQZniOxzLZ/RVI0H4pAEsZilMAQxv9DggLVYkP/6gGeSuJ1iijjfb93K/ALR6I
ni7FfcWg6KSpcdAkhYKANuHo9Cs3jXTJu3Uhk3l4KpZRfdxuQOR0rvaDfyZE6wyx
60jFRyenZ4DqJoAZ3zhemNsZsFy+D3yt2ZO3jvty0/NJ/sNLViypiLCSyzaPQR91
admG2n/MjYKeiV4wpxprUyw1BqkS14+5hm4Ue0pMoQytXGkC0y06ieZ/h6rjpDxo
gr5QnBobsTnyPnfMdE/PtlBxUmfQp7qxyUbfmTyY6dlQSvHI3j7hs/uWue9IFpcA
oAmwOQIoKtmiUrBy4UQRJ3649WeMbxqDlEivu6ZHLsEeVxK9/3vbuXaqgfe2OKUw
nqrPxV/IE4NeiA6rd5wwP7oms/PZzsqv8wjHUhVuB04AeWZSvXOkyIjmch7Zo/t9
r9/Gf/27trJ177o2wvYcYz1Sv7kYvFVBi8V6sygHBoFiRFfSpB8Lf43sO6r1Tr3U
/AHp8CDnkld8dVS7ZwqZPmO1Z7TSrfc7dfRiBEvgeFfGrSoxXNpBGX8IBLsfQTT7
ltCnXXPIPY259pwijDGzgDmhXk72Ouf/7MdxTZF0hOBkcjC/0NGRxB/Q6B/V9M8O
R3zVYqDVlfQ5d3qKgDCVED2TvG231j3WLnKR7ajGJuwN8URw3pfmeRzbas+CJpaD
QLgSC8fcMjd0C/CQfD0HTBjxGpVMQIJhHLyZkYy9ICtgKPe77R5HZqInR/FUnOAF
x5YMDQTvdOxPbd83gxu+tdbAOhITSA5YwcE4PUsE2HG/Lp6zi3/bkaKziJrZcFBy
MOADbJtGXwj0swZ1q1foHYU0VEkVGMhCfLjeh/1CVaQGYhtfioQx0pjqJ/i8LPAb
i6gHPmx4HSRGTx8osMJYkpUzk0HFvWBaKDeVg2TX75Pdb39T4GiVriW53JAxWOwM
i87pDpDA+ncri/pFwPcZ5lQGJvQInJiWsbp2KDjko4Y10EMRamLs1zOIjjW+uJJy
v0xcyE28SHzvsg4KCPxkUiH3DdHHPHvMGMfUtVtELbKAdv0ufBp/rLtr4gL2luCM
/VOKcWpMS+6ERp3ZsacYW09u9ZGEuGqxPmHcIOZbml1rSWUg1njw4Php8SD9xxjV
nBrudPC8Fn3+89aZ9lxLA1rmMIyE5YsDt+NIG7r4MJUyKT05tzdPsRmtxsrrVsHl
qld/lOMwK4XFczb5BCOE6loKCoTen4xRghZmFH3b/jPa2tfCWY3Pv0SkzkBV+WDE
pFloxX87w1es4KT5rDR0pK5qGmNmJ3fzdtb+8K6piJJ3NDOitB1LOsr5B6L5Ruwg
S4f403zTJ7F4SeDVM6KSM2CnexJbfeqQdtJsPcmmIf4V9xHgMtYyPQ9C68wHX5GY
h+HAt+GQZaGUKi3W3HP+qtU18q3GB4BVA8ZrrKRUj4PmV1Xnga2TMkKMYI+fmx+z
AgCkAOgh2d+UmrwrEh5InABziS8gt0Cxs1SkDPl03GxQmwT7onWO3dsME9uk5xQ7
tHllP2MHp5bIuFsurcNgcSvK1r104EmHSYwhhnzVrEQJoKFm9yDlX50vSQZ+wTXs
LQ5zdKZJz+CLeHOgIqppI/UenZRQca2nlXrvUUtOz5HsEY+5edz/YD6WHpbocvpM
78seSmTIWHzwwlrrRaEvCegWYuvJvKNkG2iP1FaeWxr87rFZ+f268jHEt4fZayYQ
PKBIhGxNU9MnXlMpbMkxPzCKiaGltX2ch93IiLhgC52RXZEiQIuTLYH/+FliEd/j
2+uQBQhdHy80QT8nxgbv6JhllyI6uldzPiVbHxV+qUJmSIfAf1UE4haSpJrl+W2K
IaDUkqAkJ9scXlMHcztLvw5bxFvvZWolNdv+sVO93ifAfdqYFVyF2W+3h5Z/M1CV
zUZDE2DOkjQoQ3iN5fSJrUPs/SCdGOjTooG0/sWvPxAXCtTC6IE+IrcMd8asSG90
mv0wMvh0f+zcyIC2pkSLvwxQE5YTBTtxStD97NGDe6dKa5dBGKPXWyJiT6Eg/CJV
+6GDSH9djy1C09hyXifFRTXo7X71S/khGCa1jYN9AiWdAx894wOln+k6k87ZIgRF
MJQpsI3Iriij9ICHBqeqazk7q/xuVH17qNTVg2KhW6Ia7tXrMTb2kATOwZxiTEd8
VK6vUWTqwaKG1SFkoxuj7HAp5DLZsoG8jyuHszmK9TT5UpZJ6F0c2wARUYbk7rGJ
5C4P9U7R+YWBfzd3g1ScqR9vj/yvd4P/aaOUX8BUnkcQdsg0WfdlNDeFK3E42FEu
etS78oe/Uf5eFnO07b5RMHkqQFlJTgurKH8EXX5n8VmNUxVcOwbgQPMNe0KtahI6
xJAmlg7Xo44tnl5/9AiMbt76Iz4i0ttDHwvQdWArepXmpRN3prNhVbYroZMV+XcD
4Lv2TmFEDtRL+p3LzIGB2/J8noDbo2oYC3nYe6DLFOlMlCcemJWWiQbAS8e96pgf
kUdqveBg8uXm3K1oOSHBVzY1TL7xaizmy/UQdJsfBKydkM6vOuzATserXvFOKfAN
FtlCOlq7P5bZv21ZjW8X32qdCXp27bQWJl12c/tKL0ZY8ghMWtnYcmcWcZSnNd3t
CEjr+qUfw377wq1ebgUMx9q0NYHcLkyFXtrWrU+edSLhCNnKIsXXyBF5u7xP6fNj
oLD/OpBa26N2ko4oB6XIxD75vXCtFcxWNg/6Ja5wdhYd53hYsfBLczvGrYnaRWP4
93nkvQGg35uQ1FEChH0hs6gtkrwJ1VP0UGByi/lD39npGXrm92SgNNLL+we7LmHj
5ktj6+OAaGJb3DawcTvlhZKd8VU1WqfXlNhorv+1NkRU46Opb6czRbdnSq5krSGy
/L4Qnlq5+0lU6PtUPZHu2hODvGxuqw/kMkhBej5DlLbS26vSdvwXG9eM/JG/itRp
paUiRECje2q/Lu5cFS3Z544TxfniGmSDOU2td3BlR4N+/dcJ9d6Tu1KPXuOZINlH
vpRr+tFEGC0fVdn28EIyjsKDS5hs7fHLs1iYblE6hpMyvPbFbcvdQRI1FnvJkGc6
OfWujZgjWhoNO6mP+ZPavZQw+pI+In3Fe8ZuapHkxuZ9cSMcrVZdOJMeN3fyPqgm
J7YjfdodfQsSvlU+xdZx8fi5/0u4uVRPmc3K5P+jaQTA67RnZMo7Lbqj4+rAydvS
KmwdmKT3NEire+f/GBFiY+GC1L7UAGy2vfhE3gM3CF0MFM9JePFi6CdWgNAHdUhj
ItG6kooTH3040INuSmJn6hmX5IN6fIRu8qspmM0ffdLHf1CSgHA7uDpFRq3iu6hm
N41P6pujAUai2gzZa3y82zXudFy0jyjjnBR5gdlVJINARqOQmc/t1Kx/NzyNd41J
NuCITewUXGCc3J41+M6CwelEB3AZodLH/orgIDVjINXbTUUvJkIIh4UapgzgT/O/
o2GmMdq8UJjimdqDAQJUm9YyAT8BkrFNfDUN05E7B0P8/4OmNeM7vd0o8BBGp+2x
conu6Fi2ZV4oxXLirREV2Qu/7+rlXBFm6cXyiNPTEfx1NJ6gOvUwetPmCgMmfHQA
rIbquHn6St1kpPO927m05RT58+5sWbuuUfjw+ETomsGjOTk3FaUI8sEZNaubxMs3
Upa5Ih3RQgktefbbNytM7O+AXf8idyVjrEFOEA2H2MWhfT0SnBMLgTRRqcEi1TsO
qiWMu53NaXvqGpfAy/h11xd9R8gKvDZVG2AZtJfGOOR2SjMkjMfwx2npMTiOmQ/A
29w20orYTyeSysB8uKwXbyhqTwYL58W86+wvjd5Tp62wtgiUNtUGuH/YbzuyuzaY
ADtbBjxrlmLaMPA4x1SZcM9IBqdbSunP2nrejBndS2ETxSmLRw2jQP2ISKQqrhhJ
ilfnOZR6uRKvow+7Elph3JvigkKpLE/CK6gMd+mHhUMGSvzmoxJ+0xCzgnqPFsg2
rVHKCirlJEbPuBqpnMlXwgM9jjyai/FeQBKftVzWMMUOUtSmCCKmhzrn+4lYyt0v
axvJs1i4BZhBZDoebFNWfp+dXW9xPMpZphMrtT4Y863W/oostZb30Cu22IYL+Mxt
Zd905tXetSMeu5izqTXmRjAU7TEODvql0SN126NmpmA0uPErreUNtE4E1g3SXyE1
QHYv36lYsYg53zR2FHftalZUcZ6ln147qv4JzbD6at+cubwyS3kUEJFXx/0O1G11
l+4jCXMPCkh51WRuPWnVO0vJuIv13z1U9bR9uRI1yVAXifSMebceTQ0xESfYXf/X
j5UEzoS6ooVfW8HklRUTxMN0ZhEq3nO/mJMmEi8ZEkhODj6GjtwLsR4bED/BzWqe
pn5xQ5Uz7hSXGWCRqxZc9VkAfcBc4Jlr1ff+awozGdKdSVrzxeVd1e/q8WOXdqYC
dHy/7DDvdN7NorV8eI8GrvmmCysYJzuCjLB4s7LAg5M3P3W06DOzybWYPSff1Jd6
0hzrRZJ+JsTPvXBKK1yao9tHM3JheRRU5RzUEffKvB1LI409iWVOQNfW31RdZL4+
fKHU7K9UAmzL4XqQeRYONOujT2t+Vf4FRrHsloVb/hCo3v+64Sr4FTfKeNKHewpJ
ANiBob0VNwn5Ho8e7ueE/j5zICcqN/sCMGyrIAsQbtKTbGVd93qbNayyJkG9mNAz
rGn836ScPEi37vcTkAJRpbV9Xmo1wcffpSYaAb0XvRg+9Eel92Xi1xHSrjLLmhAV
5xTx4sPc040gjvIuaPrPzRX7ORoWgVW935cflHXohnPbc5YUDYWwOVsqjabfE940
jlVgtoHjShbniBRY0h+l/qtIDKiqKSCC+DKxPPGOxa8UfJQJREIhGkwd8LWAmVAe
7md891wGehcUx795Pqe/BK5Aq3Ne2E4HRVdDMhTJKFNio4oqqpcgek8Xl1WLRFtM
l2fg62gl+MC6tygIu7T+mfroQurIYo+lj89jedsa5hITG9fjWcca95cNbpDJHTeB
4pXtO+FiK/Z1dwa69tMdIGCwMNZfuUG3IFeAjknYyZMOCw4TFDUyG+Rzdhrard9x
bjs+Ob1aFndfFO642TOjd4lxWLJCDpM4W3uFs3jmo+OOiqF01KAoeM1lqRIlVmn4
UKCrirIiQ5Sdovhpalj4V0cKUumLiwVgY05Oilz0GztISywE7nnlb/TRdnyatAt0
8ivt24HP76DU8b6iNB4xW8CH7kGWQ5Z1Cd/wVew4yTsLuZbpA5nc6Y2m8/Forn6a
+eYEdi5MHetRupRaBHbhAu/ohBUbFhGgBrYf0N3yTFMdpKBlb+JY3D7rbmKt+Pg3
MPPqIN2lZKsabVkWg8b2uo4VMw5fSvE8gYnmSSPFZL9w7zKQmmY5R8zgmKnmhfm3
F8x2BsHyc7RQYIADX2s4qNmKFj1pv8XUwVbrkgKq9mjbDn/KMwISvM8YnqfLSIvt
vYXLkkMDYz+qE+e34IRWWhrFwh8ZIxpdcST4r5SKdug9vmxzZSt7FK7Z9TbsnKPl
WFywyeMmbu1wCyfNt8ZI4uf5GVxu+VpTSR3EN/UY7/4+2zMp+YuJT7Awpw/DHmxP
qE1Wa77xkX+uhBGkZTuPU7oMbpedC0afxAS3iOj6L7AOLwR7uBX5usJ2b9nSp+bP
d/bW5gAzuX74+TPGzd47+Xho2QG8Pr+zgJjc9HBGY+FK9ige8Noc4Vlymv0EPym8
hx+8f7Ho2awtMgHhKLWu/Y5x7z3hCeYGx+WXplD9GgUcutNzqz7NhgHrheaYjolJ
uvQ8tLmVmPX3UIeo02WiQOQ3gVuxa+BXv4tUo23JPi9G5syhpDeJ1tw8GT7Uwv6e
Qir9uSnbt0rhA4Vfn93TDAPYITe8zUqyoFS28Ly6K6I7Ql2Uq/5DW2vTh2jXWnQ8
2x39MWG+cQBFA6Ku1wHj2S0C7ZyS3deI/xGP9OG9Al4neJ9twE7vE5ZHFnXPpYrp
R/mQ2pfXf0SSVBw0eqNDMiMIADCvAtK6x1x3icPSCYDwsr/hRghBwp481yBl9aRN
6SCgqfm5e2sfwjnarUNLtohysUX7kVwyPTEa6Bnb9wk/e9d3F+MeM5N7nxsha3qW
jDG3tKlVcXhtRr1jXkKUAxhTNfrX8g2Zn4rnmD6FBwBZng1Fn8/yOUarPeVEK1v1
DVX7ykdtGAE3LmTPRJmO2yBVcDS7/J3I3hUhFARlG/WR5h+mnEcDBzJzxeg468nE
Yl1Rjlu49VaDyEi/hqyHrXxxPaa4tS6bPUhtc7uX0pfONa0xLXCiGh//QmpDOJaw
HX9ksRtFufHbgalMjX6/5nLlBy/Bcm1Uitg63RFtEdn6vJ5DfXEn94YGtkjR9ImB
LeuXIjfm76lgVU0cYHnQuOAGsFkzj/OVWWsnnW8S4nLc1KA+DxYLxmhygoJ46lh9
4qUCnng7Wavde8qGO8sLVfqBtOl1aaqeaNpGyPGN7Ucw0XFGfEGmM6FSeZrvJFE8
W8harCRCOC3S+NbaDAyf32fnrE016lGim9cutOmBAh+OpZuqZqQRZAT3/CmVnhvT
SZT6Y6ErA3KT2frJvhajnDXKthoiXc6PyhcABP9SxVD9YosWnj0+UU4qRm77r6og
osiP558gREW2pXHeeZPwwBdQG3jw6tkBOZQrTvkQFk7X+ZEJ3dEFJqEeRiHs+PyM
aY2oG4/NelKbPUJ4sBqbk9eH3ParaFecSdF1GCBYHVVIHFjDZI8oSh4PBDb5q+Qe
mJoOpjdxIW22R4yb+iJorXxO1NGnRgt82C0aNFS+2nUt6uzek6cY67N4I0SJnz/J
2mFTbvdTH8BD+TywBdYZXtr2xrRVzMc4VRF1Lj8HlRp528g3aD7057HqfDSCc/lf
S/J0but9yqe3RAQ4siXnX0sddPwuPGyVZa3hMeUApISru0poyiM9sUzthq/oBNQA
7xzbJWZwLlb9/M8VIRNg5WVhTCZlbfOB62uASSZ0L1S+WOgv7jvUu24+P9LzBHOg
ZBofw09pFXQLdNMPTsyXdkBd+waavQsTgkMjkPOA2mqq/PJvBfBNND/icy+rdh41
2gJh2fl1erRyA8LbWKr1n/zf9+Emncm0lZWIIVYHozpRJyPexQRwn4S27QN6zurG
yD5fgyJDb10zGyTaYasseThWFceoUQudNt7FPaQAhRBDAxaWnPPP7fH3CNUcEvC+
+Re/ydKEDZKU7OW6/892buAlghFKROWMgrHEwV34XceI2Wn8t/cwdbz8/qzLenPH
edWdV2hupvmhzm/WsvFTdXuOwsj30JtQf+u5kZ49NuqVFiRPo+jrShsvpl8gUWJL
S7LCEpTO6t2Mjw8l0h3b8xPxyse7A6Lk6WB3q0Ao/tG1N7YuJ1LVeqmHN4mkswmx
HnBlXKLTWSZmDOlarT0aWFnLnzDr/2NG2YZeKtZ4X2F2dIzthwO3FMaJSZQ0f3zw
SkAwBqG9Y2Zoya37sYKs7+dIZK530zeZ25U9bN9dnmX78Tw2De0OJUjQU5Lbqcvs
oEC3MWUqftbA1RnZYem7AdZlZhVV+LCfwjzfMWVYfj5rH7EhD6psjFF7aiJWaftk
jCRHaDFR6P8CTC/lqXQ2k6/g2/muDZsSJw0uBqNMJ087StrnlDvOUIO/uikKrclR
ENRvyJdM8XNsUn/4+NLXkzbj7EL7DiaI1smxijhkZu4gakwLQ1fpaV8/kGyMc+Ol
icyNB73JB1rE1jB9aY1pdYKcF3qVSMuxVawJtECqIL64TSI/QQl4SUEuNoLxn2op
A6clX4LROvqdL5jdTW231kc2yerqUKoWjQ1cBvask1Y5ccPTAX3/lOZjNEeVoslW
hLfqdnIbjBg+VUWAVvHBQx50X7GAcjEsvX8hBDwLYSewbriXN/298kMVjuAmg5tk
4h2bxsPa+owBq6nlEuE0e6G5JaZTwPTSYUEzOKjgaCEIQRPRqpxabRhWuTTpvGUS
NIk+ZcX9MDUUSP8ar8hpKz3E1EmIWYHdFIYgHB2nYCJjxHvEtoWSf/p5Fu/vqCAW
N1qEX0q7vBcrEGIhL5V+FKGIcFIESglOw7ZB3ZTKKJ1CcypLtqZv0H9J7bz7fjqw
duaMmG1vx3E55Ze8xBZ4gwCq9m2Nwjp+Idsp5jxpU+MW/fLuZjxiPaDhhXUPyQ6w
y6Pm/e0K84R7w9tEycl+zo87kiSiCinCEbCENPb13lhcWgSbfs9CeAtGLGvTkVeR
3/YXADjZei1rt+rxcspXthtgkuL1XJ9MFLROWqg7TeyQYCXNLnTDNZ5vQzBxCheu
DvOPFbtv/kRAQn4IJLuzIvU4optSsOtfJdnUHDf+aDOd/m4YvAL2XKPx+3+YQrbL
+xY8+t+6nDHY2yfp+QnCi4aI69JQSs9nBsqqvu4EtSb0EfE2Xb27LjP26RTTsa4T
kTGGkFl31F1oxcANwE/MXd5Li9MFhB8pT/Grc/Fhn8lyMcn++bmWDzpVtbL1YqiU
ompRzq4PgUXMX2NMUdGj1yDciGh1aAaK36SlmgCFIO2HC4aGUy897j9JvVC6JAXL
bwkgdj81YbJnhu7xKM/L0qBMUWAYjtUB4n/vkw1EdErI8ZvRp8x5yKZPANonBkOK
iei4726Q0L1/BcF0XVdWpufJ06DY/CsaqE/2ge03oJWXDe+R1onsaIk2unnsHF2C
TX1KiDPydRLvZqhsZBQRwvu3dMe2uw0OtagyUTPua/egEYJ2T6vwE9g6DDIfr2lo
k5sOv5Kk3TKF1k2MbHUXg+9bvmasxz0xAPyQh2YZIxDLyQC6EeCPMdNeoNPL2EF1
Z7OFez9fR4MHTK7ojhtyCLKSVdbJpInCzMfn/N9XxWQ2mF+PjhNdxLvhN+7iBZSf
tFDrISPzqeF98m6e4U6J9qp5I6vcQK1RspBoELSKA6zTEN93ef0sGfuRJZDMKxgp
ITzkhrHS3BLRzSVHdeVrn4lOv4XFcrYaBRh1oLNR4mcDaNwmVjWoqwOcUkDNE3NT
Q8S5zyrfWWZvyMCeT9BQVNR6h06Zk1lRU5aY7oBbMpPeUwpHP+klG6VeTiZEpva/
bzlYUQ4UK3mjIGDJLmmbNhAVS0aeOMHOHcntctgHYfN4+4CJTOLGhwhlrtcZq19a
SnPvV8fULk7shLLb7SDasCsLFpUD8A3vjDVQq9L4Yj5NTSfD1A8NRihgqoEKAjAJ
X/h0yyGHApLOfRR4JaWZDMu/mp34mx3oL1QCQDVcekHQFWD1Nv8I9HcvpzTxEFmo
LnxWHlGn6VWAUfPDP3KfToJ5PWfog/pT53dtbHQ53H3u5nxM2VH47ziXeVuWQ/aF
pGwxQP1rzscu074J+4dO56QSzEuuny8dpgXGTdOn7Xd1JbRsmmQK/6MwVl2wOODh
1Uy8L7gsLou6riy/5zBX/c2k5f7en3aWpRW7aMxBXy9WGifSm7j4Zq2ZUb2dG2EN
mBGxuXgKAnoj+WINRzQanWtdguWtLt3an63sptNFAfv7tWVGZl1SInBYWXVElSDA
bnwFG/atnRx1s8PJiqLvG7vtRYIImKFV4BBOURu07xxiDPF53swfAJeffQz5puBJ
rw8alGkFhln8E3WkKrv2RuMSwjm8vKFCjD24dDfFWWZYkawK/9U0mGsfNQ4EFm1c
txQkn1gQH6wNZcGCBq6h8iOS6tMqRzY5KO3mJnWoxnZmw0FlcpPdq6BCiMHu/VK6
I6jF2f7p21M1RMPdvzv0JmrjWFZtb14hnl+5fPpZUk4yzYAwBMwcrGgdL8SDiiHy
5vZZl68V6SwSyaKSwdYcmVhlKEHPIhJWLH2Lev/foBpcM7YJRssEDJddOIvjtvBe
6rKHVRyDmkdhm22KtqN7JwdTEbsDrw3TNvppDFSRMknNjPgrhma9KrdUChCPntZO
2yTIxoHEhL3OIoGFV5vstqivDyGnEjqckyw/qAnRE4+JD3725jLf5jXzZwJ8TB3R
iLdz2t/T5R9AM2IQjQVk7VvhNEhDOtxCxmZRUvK2uIG1quBnm3JZ/7bVNZPgQtxk
L7Od+4kwQbG+AJn3y8CD03XgQ8KYdUS6cXmx52YHJ8GkG85FlxpQc0ddZ/2ZYM7V
nnBoVk1te+Hzf9Rpyg/uoM6uzPdBfwgR4uuXOLD7vTjb6xO8JpWDBVMaIqdr65Ey
qBeSJz/Dq43KEGnJhzCgJ4Uw8vix8PpFAoP/X9iU59T5J75CNHH9aVmCtP8+6wdd
9ut2isjncjjqhEf7PO7uIVDhde5Q319WEMYkR/sv3SDng9lSsDiPlXjpAfkMz+M4
366+KR7hweK6n0RQk6R1l7iOPccZdODA9gJfDryyCZx1Jvl+GfNatdXelz8O402w
1F9UXLrzGlisJYrKXGHXhGYKKlU01aAJRDyMFJTTUyqA/Ws5ZIuyNRB1gaiw2stI
6lM5GwYMrX70VmFJ72jPmlQVs/ZssGKELUtEemfxjk+DNAcm4Cxi0dcjD/aTFUfk
z9zcoo2REHrhyKOolv6dkLCq0fmYV+4uBEdPHeqbhIK1JtTucvMpVk4qfNkuF38E
CIiW9Tl/YGtCjA9unu2XR6+DxRtm44xyLGzausavNZ8JOnCKBr7v0CaiR/2sQ5nx
o7yMwi4VIADwpE19ZSKp1eGSSl7wPmwuRduC9jUHz0cyiyuXqVpoNvcGpMvnjNM7
EaJx0k9m/ycIawyOsSaeAqeD7jEU0iddCUTCsBXGIyxNfye5sW8FzdI4eCV57Wt0
amZrWPOGOsb8S6XtM+P8cefFirONbHiHX9afKs7xaxRXqOwb3XypvQ/vXySpYb/b
9Z0EvW72VWYAfjDHnTGhz426pfz/oX5Mwpwfnk59AIiDcrmFxXvCFAsb2MN1jTkK
U+6MfCxXKOE1JMlXfmZzNM5gtLCvTfCU3LiFCweq3nO/iA2jU92ZHcL+y6kkqj/f
Y0MNCVhUqWm+9ANB4A4No/WnVhwMQG56PqMEsXMfZR0LiuuUaiM5Esb9cQR4uwUb
857p0jZNYE6RlNqzut3lTYURRDH+8dbDS0azvf4lMbHzCh6rd6d1J26TkHS01F09
Gw8CMs316Dv14Hx/WM7yBl+sT3JLX8hBaIlAPcodCoRTNf+COCgeifkVY3Er8Fhk
mAEE1xeYf7v0qqq4P4F7syfJ2ZYEC/vsLR8WxWna6swtSk6KMi0ill30dYzhfbIz
AD8EdktleEZto+KS8v/F5lyqtmlAeDDAv6QQzR+/FlEqBjYWj7w3CTO0vmhJRLbE
zY6D5KcExEGfPfUdTdott78Vjad1ottrD/pLmX+QzYBXH+7ZDXHQmYFEDnujAEqC
ikTXkGhJ+dYYtev8Eb96S6Pu+gfpWNmmtXkBEd0RuMciumhQPEROKZc98G7GDWdN
z01+vR6DBmGVBXF1iZGmlJdOCGJFKpa7IVkiqVoEgN55RqeAfbly00aM2BT/bOFG
ZMnFqpwoNHrtoHBI6d+xjmms37SQjikBeHxAJq3Wc3BViPSEg0ums+o0eykWH3x1
Qbv9LLKZDbCc/R9Bh9x57AmP2w6d7S5mzMpAXk/wSaLciXFGbywvp8Y3EdnJYbvi
QDsQxlbLtOMkxEiH7Yv+tC7+A2g7K0kxaB+i8xgSRNrkioeKgODmZgIEvpJjBggV
3Mz2d3cr4BIEncSQ8ZXHIJ0iVLDzMpGAYgufna0KSDH/E5zkA3IqitaDTjcnLyJT
g5BBHdX+qNYQKtwKl9d2jZtc7lKLH82TMpY/++6ebmQeKo1rCrLxqaBg2tOsvBnw
nqXNRf7R1gDmpg4yCAH/RepTBTrlO64ibuH3GfDz/OZzPyqw0k6zkiziCiveqo+8
XDVOAm76wrCpaBNjuOYbKUR0bcoyStpFalHysNAkrn9bVtMIiOJMeMuwObMo2mx1
218cjme6+SaBA//wHYKe8vXsAbKxvmYuSGIny6LkPGzOVIBIk6Ri3IKj/GcLjmgh
AjlBNZVcMP0Pn2M0jz6EO7t9OXt065t9Gy3TR778lcJjmYhTF+YkK28KY8ATrO6v
LaBlPsppHpfCPHvKqc88lgqmg0Q2gtLOwYmMV7vbSEj3L7aWFY6NWrciDdIHBGu3
oUM2TdB9CDn29ZKJzmmviRqFMe7QgVoCKenrKkdRi0py9WS5NZ0AfK1XigHZ9sO6
NTqYu6oqFFBDIK/eTUOoiaqZZYDIZ5dapx2Xp53MV1pfhcsPiCKMSquYeIeGkjVm
hxJ5iHe7aQUxYPmoabR8MQWWyTMx7BsBuxQ8rcoxa9n3IjzTrr9fWR+N6d3WCNnO
ci9TDn1IRrgc9EowKu2OkaJPojJFia5dYwF9MjGt73HjIGmX+70m5o/KXkIJY7Hg
oPMbBK8XbMWqK1bRMl9ej62ghd3V9C+fQDzOPSsgIdbENy+5iBSKVTJLlWLvguOh
hpP13+ca6XAf1wJvgOvYJHCgnZbdX4I1uXOxEHXlMBOLHwc6etQIuEVY9l4sypyX
SebtsssoAf+dR1qep4wY9Pqul9fRH8SAHOELVjdxfmFtSVPwr/83VDX7pjkPCA/9
w+IjCcHDSaOkT3hd8Dbyd3e3et83Eo/Pkjtspacr+I/zMzPTespe0EQvIxA9HRSw
LVz1FzAMv7zUdcGX2g34FJBq6qyCziMCJusLAdqPvy8C2Bv3p/CaXRhVUSe6UvDJ
U7QxBplq/NByacFcP6e4WSusNwgv32Odu0W/R1i1LpfRZ33rtw+iKy9wcbaJ3b/a
0xyIpEp12e0KmMAxXjZat4GVij0Ttk7Eigm/z6lggprfZCq0LOD1b9cplnCbbvW7
p7Ryodcv7z7oWlLRzTokiMrmNKDYvsNNuBK1e3fFl2rVrkMne/IeKDore+M+r7h6
ickXPHXr2ZMlmibwU1G8nSVGq0r6kLutXXs1QEs1gk1qxF31falZ6ffDSh8sqbvi
0XjQzTaET36sok7e5KsDKqeIbMJ/r1spZzdSXIeim4OJ5hnHS+GGh0J+r1M6sfIw
Y1dpuePTd4INwcgLOpQS71V5hBZorCLmbQpIi7fh/FV+8nLFid0JELb2NpAYh+57
W+z2hBwjcE+g1aBGxD8gg2ugnspBuvDkjDcib5HclwiMcV6bUhWNyTRpXRwhccCM
02rRrzY80URfD1fju9Sp6V+6ZCX1OXrEB7ukI5xmqRiufrFUiy3PUH+T9NocbdLK
2ZfhD9E/hdSbbbqrLTGL6aUajei+z+rhqMkaWRh5cA2FlU6LkR0eD/kA4bZ89f32
E9AEZtTILsfZPSYJUzDqrD2ri0nhdcZI1sn0dKBjPpPZmRtLHrS19wMMHnHWVF3k
k2ILjIQu8nEloh+4nfnLqco5mY9I3l/sDNIT+iyL5/ivwodY/EbvUks1FnGm3Uum
0lCYMPlUVG29TTtUc+uzNdpncDucwZtJAaVO84+Jvfdw7JLNDHrNoLDVpBiQarfT
Jb3euF3lNowF4hOIcDg/Gow5KaBNF3/bq2q3U0aRMd4u94WlpmYY/4TuswXnfVgp
S2OE5l9BlKmNkAApfT1giVo3lHCtBTzdLbbNhM6YOwQ6rCVc5O98gzJ4ITVAI8XM
0Be+3Jlm93TndzXZQ4YDeI2coKLX8thWnpEq79kCoBzu4cp0HyZULWI2DKz/H8Nc
PvK3SUu2buFSVsiqm/apKRTpImQ2qs6dl0QkE+ES1jKUgjV6bVtFviV2ncOeLuQ0
HBHO+iZYGTreAHTEp7tMHz/zcoSideJPcIO5Lfhiz1FV2A9gAhdH4QK//3ixnW8g
IQlKyzAc5EfV6OLQ3dH7IfdqGIV4JZgkbTUbHgCSDZRBmufapp+kBCDvHPtLUkxB
SFrNoluuEzPlVgTWkD0iE0MDTFqwTyAjQ22CBmBMuEFK1APQ0K3aaRO4eKz6JZ1v
e/14AcVmLZIFmNbXcbKkZxhPgfMjOOSt4ntvJMJ3Ok6nyZ1up8YAlgul0AANJpEm
FHYQBS1IS7snP9Tfjjox4X+WzKzUH0Zwf2FHdtKkMT8ZmxpKp/TLOzAs4C3zKfyq
wlzgps9PPFzGVWcBmPkLZnPC+rB+EK86kM3HF41ppbcdwCF3BOtsXFvsw6bjujHV
w7A1fzWKuMBWPEmoUNLjmbMblf6rl5nsJwzE9DetaHy+4k56BmGrMzkywRGqnbFE
1knOglEuwDEMbmm2uBhjv2651BfblR8JYLjWowsLBo1I0ttOAVUoMkUSvhdhzl8T
/+CLeo1gFR7cYkO8cCTLF1lgJpnZlR3Jy4XLG6/KL8KgGgL+dMmNJKVZ5p0EOrrU
Kjh/U4ekBS3ofiK+WHP4Kc0Xw1FW4Z87Tw2G6MLDdKDuc1W3tmY7lTKbiDhwrz4j
npx2sQt75ueTiX5469HLgL1EaqmgqFkp8cxZ0anxSEYqOrQqSHHwvyLEclpawg96
dyH3xoua7kehZBOIjo1DsBbVxmfuenpLYyEX3oUQjV2pFGLSq4NyW/vmFl8v+0sf
ntGARfeKWbekxWrmbu8q6t/1I3YL7dEsxk+DMkym0QuTusISVpaI61xS03dKA6Qq
L+BgBQ1SD3NgmnGaGkTfm3G6MSu4Uv5evbkI1sTug6MWuE9s56tVYL/yxaZJwifU
5QuZbgYFsZNMu/6wweF8YFRlvEjxhk8BqBiBGOLlKpG0Hs02k1AhUALfXmSPgcFN
02sMA2h8g88+qLjUiMGFv+PiHwsqmiqsRBY6eIMj9t8bztbyKTILOIk/ZQxpIK5W
ldTXQie4wWDTq/Rlak3e698U8XKHdSptqEQL3ERVlerjOXkT0aOCJHG2SGMjpbnF
/idFJfr+Vd4ad1MitAbOGXJ6mbodjpD4aqC/HwqXSipk1leddzS6M1Ldl56Kj7Mx
RSTgp6unDO8f0SKCCwIm0/sjLiG1a3ntYe200SjoclzcEJ/DHWsl3hhVSY8FS9+u
iY9Z5EusuuthhMvfbo4Q//pXntbaWTf6xC2905rKEcSDDS58LeomD1cTom6vGFSh
kB+jcCP2vw78POC/ZPAiTLRXqWF1Audph+NPdydOtRM8L4rAMlDdcAC7NXMI2AyE
wM7XDrWXbdupSofUQeLGZik/h/MdPRsqDAyMhaxzn0Sd5NPrYFWiwOJHrm5GAUOr
dc16beK69jFzh88lu6UneWV89+glXRbbOjojDps3nAhWzFBTuKLU0LxcOU/Q532Z
9jwhI7u5C99uE+tSWRnLPurZZtPD0QDwL5NCyzAxLUyVFcni1+iBQ42pD9CZVe/x
ALM6umlAYf5im+Jtx4F4sZh+6wxBfXNmS8i218d48FAJouiZ5duiQL1eDG34g3fQ
fm53gOzwIH3lW4P1A82OLp79ETC/meLJs3oKO6JLwKLWA3VRTqSGWtCoB1qNq30j
zuC859QptzrMAmIZYkE8V9u0wH/pxoYSwcdIN299FcW37wveAtMy4LVa++2jCIuA
PBujczsQ1G9ZtigqILOsKNT18Ez41R4BXDSYDgRMi9sU2sLGYhJvoFz/sDNtfhil
AAQC15AjVq1nqzmEbbgYing5CFq2kG0T+8pTwndk9cLZIpFtuT5mJiRc+bPxbRR5
HuQQhk3C6k7HWf+5CkV0hoBZ8Lr3BB5GHG78sbD+4rOSOWAhHZwnYPXMpW5LTdBM
aW+yc1MqSyWLSUQBWP0uW2pQ9uY78LX9mjW8IDygRHBYTLQS7Y6Usioqv5zjSs+P
GEQ/PCk6Vde426LSpOayDFrAmQuGLVvBNFJSdQT1B9qbMMit2Y7LTpU+pbg/7JmM
7bCS8ZBuwqYmU7QoOmKbsrpAzDbrisjfk52IkpskcaLvc1sU7Pc0FUGlpU1mhm25
gTdGC5ItKKz1vuPCAvpZBPKdvvt1vTxewqiuDcAK0S57z3XjUKXQnL1heqlAstO9
TO1lPYoPuVM4GYsIS5h7cG/2W0tCOHK1EdcJhKNYjIAKTl2TGj7c8/jmaVIL76vA
aL4VZzlx5UKaRtqVmLOMuTVEm9D/nKFbkXBL8VT4Qd9Th5O2T944R1mptee9YlU4
BUh5V7m8bEHTgS8sdq56ByxRrRDOtVQkwk8qtNnKraRE4dkv9QqbuWxeQbDennnI
dsrdpArbk4D122pl78m8DbT+CKsfq4pmGFPKKYZxqMnNMzN5bvnuNyeYj8jvY/wm
h+WVhwzOZaf+yPDe3ZpuPcoOZuJtJzn/Yj90dHV4FTJ2KFSIVzIavBhbP2NbDaMp
vfDGdyebCxjA6sVuHVaTVQHA2OS05bPyDoejdDJt6CwcUPhBiZWM1XV0H2gTMApN
4Mzgg/R4pulMkBeJLuaAJP/2Hu/FqblPH51kBfIUJE97iwwdYcExmFYuNy7fYG9x
MClAdzDtKdF8b82AFqv1MdT4l+OJo3At1xPvGJLntOYdvXLy0k6EIwoPXEuYPXyc
kCcBEoYaI2T0gHJjy6hPSvClHRyq6ck0tCkhFqAXsRM7kLe8SFScNklunFjG+/0z
GRMw5K7ZMrhfxNcsYJXX/8UY9cMtmf9rmBN5r51kB8JlREnTAcNuxcGHiU06Z8tn
RYAOKIWNcd8to1UW0rET6/aAIstirYBtupbYSZef79rgC2AYixmSdgoxjOIBbV0s
F8Kn4jkOCRieeeYpT5wF6wwXU6yTFUPwumliQhWnIkRSvD11gRgasj2equ7m1f6l
ZDllE3zOxulXprS+fJxoSDof14GoR/iizlMWM7xHuF5ZIX3XVSUCHK612N6PNQOS
StfYIgh4guXKlL5BicJzywaYP0a+0IEptnoEvho9QteImZDNoFrsDDp1PwWuk0Yz
e+6HnNVfo6IuZrED3DacgEhpX1NyyAVef7y7bM9CZIF5jqhbuW1GREYoK8OrclOC
tMG9p+sFDD5ydIqF1G28M85A2I2hzOar3uhM92cW0yemXa0th2UUxhr82ewiEYTY
mhT2uodNMJbvnKAMriPnAXwMD+huvHZtEFamHnF97Afyumj5fMw80jRb1KAV/JPn
7JLJP8vYWDijIwgCeWXUmA4rjHbqhGd8wr4NRPHVEKJnCKHOQIsHl86YDksBKTH+
I8B4DDLiZ0THPVxCbULpidV/za9LY3iN6iKOdekc0c7G2f2fLrHchaAuddzriypL
SJ1ON4RiGT8sIsjzHNoErpZfseqWks7snORJx+kGCbZYrBhESMAWyZ2caofTTKYL
1QJa68TmkJYgXutja2OD0L3aeIEg05dL1q0KkdjS0FXTgwwi3FUn3/LaSX7/t6Ki
jxNL373svAQdSJvG+HUgg2PP27zwtsVovriSl5S9aeSN/hCjP5kc3netIxbVI5xs
s3UxYafBbTBwtt/DvMH14RC3nTtmcROBVMt7klVWL8ayiotI8Y/WudIwmsvedsz0
PQtB+qwhNALR6PRY63cKbadJRMhOfHOzL0up9jJaMdENiuzm9Gc/Cx9n1L5U149d
jcCX4tOWSBfc8xeGGnlbd8bgswkYBGSEACRzvtfp4ReS7N2Mo7hBAFeeLC083kgI
akkIv7xnL56kKGa6D0zlFBzW9PrTXOvEEozYqPSHRF/0IZ2LcegNgfAnkvfyQNpo
sY9yaastGV43MXAaB1hmArsAhudSSAVA79gatlrNJVsmdW8he+AgAFB7JYylcnwu
OZ3+z/GM9AFjzuV88QLDxhTs0izxuJz42wY1jJExEu/uAdmtJt0eah+AaMzkXLAZ
ySN7zk9QUuAeL91ZNOX/3hwiY8n6V3SpoSfFMMQey7eFrV75ikVwuRWFiDSTZCXA
qTTo6TBA1YhXBQqJm+mBCL/VyfpRAfKtM/gZSuU6n1RYAmSG1ZRzdAp3vFE3BVTZ
Idiq67zho9Nv+EDdbnf4TvwGm6AAaIrLNgWxVaj/hzgxXDfHwhDKdbRxg6wJuM3D
u76zVE854ivu5u2h6Cvu1yvpADMsaU8l35XMotHAz6VNG+bxya59lU75VcG+ETC1
onzjF0OdtjwH4KgwQQLMzYZzqqkEg6ZqrPxzlwO1vrUM1aDT1n8iu56RV1W5Bff2
F4/GnjEfMpDHdBPoDb69CNSkELp9IyMLSahzXR+y7syTZwJ7hnmMPA9qQXIEkauY
fcRpJKUbN9RrBB6DqtolZprffwV+n9AIul3u6A4J4XAuW8Pekqwhqv8B1Cl9AazV
7oO1PxUX0qhIIOKBZty7pTP1Nlh8hPCd+G4sdB8GkvdC3uLygYHSya6km6EG8P4j
LBjIZsxn/pw4YC9T228d8mdQc3vvPVrDwGzqahxa/HYNwr/P2QtoEe7issYCWpgu
GRccIJ5QqglXvzNcArQwoGeEuKAL+k0kDtr9+HkmuMW2T+zREfAw5o5u2e9T0f3o
3sFY99a45qBSw2XOlI+ed9D2Pwc9lzwvvDMXxwrHffR6Isnq0rJMBbaNb7dJU1Kh
dfDGv7EvS/qRpk4Jgsk5PHJ2bBG0X8klB6DkgieMPbVHk+XX2jf7RpRyxQCPymJl
zZ6dAdup+dQfXnw5sVbPKKwVNJLFDmxg53LtqABj5SW5ITOn1qba8/yqG5xwy25G
3kjY2QKG5VSykmz7hhzOYenBq3+T5TV8haPiZtyrG52i/U2SE6Wom0hyi80/jzT7
OFUUdHRhTgMmtcntBVDnN2r0npZr96c7t67KfZr75mNQ7DxURGGzFZze14aqZjs6
5fw5ea95l4trQsUvx8ll/eMIUJoUKfh8BD+QZ8+wXZH9Blct4CIwJL9nKlezzTa3
BPBL+7bD6Ch1UoCjLnuZmnNdtKweirXlsMPxyOSZbJ6aLKvfubmPPktNfwP6tvv8
Du/U2TsCRSU0WhY/qi+BNc+iKKOaAMefQZvIqXy7TbP4yqmwTSZL2metnhI282h8
25dnCvUzHn9YFE005rgjZEu/WSho0vFkKhDZLxyC5PDwtJ3+Lauyt1dbKS1I/V4d
ETdPcFs/lN7MQCdVbTASU4HKEKau0weo12PBSe3Do20pulKHfdgbn1ntiLMzjc+Q
ql1LNCm1pGGOcF3espmLYmd6rZC7ZAzV5+UFOATRgLPgdv8vpq3wfMkqO4fvLDRs
4o9rWsg+wRLJWFMNoqhyFob0tORvUDKHVx6U42xvPleFIAV75CrkZ7nDke0HchqV
90f5wGNQqAvdl+9QXFCarL2wtqpL+JyVkfuaVNwGY2b/GV72iw6zTY88p4fBDCTK
YujB3zYKGtreZuAvtmANPe65eZ+lBVdrHHOCC7nRPlxVIMSRSBppL6qBqIb4lHEt
06hyGjB0eVd3u8voj2F5xHCQ/9PEs6okpYjOpJJA0T2YZQl0LTl+4QKVBskuh5xU
H3c6c/Y2QG4NYBUqTvZu5IQVKMnBvduwHTaIJnabAA1P86664qbhLEwqeHUVxecO
s3RPz7PQqdkMU7c8F2OCI3Ace3H3oi2FgFIvJ7EsQTZYjHUHOKtt4vCvLWwqLyef
IcatyzEUxEaFXnbNDlEtkv+HLBLPxqEsZg0aUcF9kGULINSHSpDblf5dEIrYx2oz
3xhMa8KcIbf76UMwwoUlrtiNb54pPdUp21iVSpW1Cg+utCkC5nMPxmu3CNFr6Ve+
IclgYWE59JDVi70teZ16HZE2ycH3lSP3b4AdTpHeGOBbLKxW8tHuToqrdja81Im+
Yx8Bs7HJjt+rEcVtq96PaUdtbsmEBI9/uRj9VMDDA0/3tpp7OwTnZfL7RFmD6EPy
yGj6uZmdmAq0farBjN1ztvJyPdsL99RT9akewuvt95/JWQulBkUrg/G9D9A85Gp1
9qcrESpVWHGenwiw9wnc/LdImgLR+Wo4l1RvVJXEISpRHBweSy/er81/jOmUg49c
0Qx+z/kSfOKwWkO9E2Hn20IH2Ed8kdbtiXRKJEXkDgmYc1ebYxrvQQYjFPKR84Yr
eUtYyNNT++CURk6RqNyXdYz+vMfFTTmD6yAdJxpnWAy1nXSZHz2Obawc8Un/sLSu
vNTpX7PjhapwObtWv7W9CwDFOIsRFjdtYooS8BdqKaWm4tA0AnHNPqxmI7ZkFjLN
X1EwxhT2yFWgNpj/EbyMGd6z5JtgCxNCcTh5q+FYDOeBPx+A79pz58bpl7a3UPjz
eNgrOdP4llHE2C1dTX0XuYK9+QNC41dW1Zt/64BncqjK1ujecWIDsyJeNIpA4W60
8Fdkg8UC9ntb6hyug+gXSEKNEA57+xxM4Kc3PYaS6VkhhcMIOoAAKDX1MH+ks8OQ
PZCP9WkoMe1vHiPlrvC1vNTPbj6kSgAj49jV6u1rQdG98yqfaxRIA/lk7OcSxclG
+52zD0OJXeedsTgxbpazcMJAz4nuz8T42L43IIXID1PzWjP/5i8ga+A3Q7mlUIAx
dC+2nU0/Z5EG+Q5SiJ5IX5koXtP0mLtgBXCzSV2RFmaSwErtKZMXRRc6EIqxulVR
qMP+DSyhBLwV1MDojYtap/tgLJkKxiqG0OWlY8X7xaSNQeCtoIWZFRRsrk6Sh8dq
7WTZDgIbpIQer0cXzf6nRKNoW5hRZI8rKMEVSBfLtg0sDYSkp6BVmXhBAAlVBY0/
zH0Vf2EeDWxX0M2Z2fu42AAVZfS5RfVn6EYGEwgldVCJQxyUqSPM5sfnSSCqzC6/
13oHXt1ag7vQhiAUnyBryEkFK5i70MWguDqUz3YXFzEAc81Tq3pnMLxXbDjkZZQh
R+lYjRA8ee6BEBIhxeSr/cZICOZbPJeL7kc6ghNIUwfT/wZ3uu7lA1T2F+1bi8Jh
cD/W8FhslNcjey/nPRrsUCPCAMGu7YUw4ae5d66pvwlwgzrAG5MJCUIGOE/JYUOW
qYogfaLEJg8/nC1xZ/cXXo6d3XvSr2ACZcMDRPhvM6XGo9CeBbCAgqulCUDB+3n/
/aakWA8jbELTK4KXp0Qhqp4AsjEA9UMF5wPMYVf14FqwO2/WRXtRfX24bkgBnxuy
AVLpx3hHthiT7HTrGh00E6asNHINaPtHNhApEOYTxMbU/K4LzkzXo3dYZuvqKyMa
n6lG+NhLV+F4pMeTKN7+dB+0cvCQm7oZtuJBD0stHVYYkXtHtkaaMkfzGtPT1OhD
u4ML4TuJ23VuKxbXWosQ6PdPThqnmSpV412unbc4kRc6pWXMtvz7EVMzQ3jglv7+
SP5BC7Oya+JIlReEv6po9gPuqZY/ojkNnsS0ll5gy9amInVJreB6uzmxhmkODqz1
/Fcp0n1sITD+VU651xeNnkmeiDjmcgHMAFzXsCIXC/vS25YosUCBJtwegjX/uSvG
go/mhBtAeoQYvnxUfLaoKLXGoWyYuvH4Md3LSPIbWCg9wf12LqnmLX1R0lwIcTuK
C8bw5487eeJCAiBMuI4/gGQAcNM4fuQJ5A5PR/ouhpyGcpUaxKAATUtFO/ic8y/k
ZObkeJEQqf0MJ38hi2jWKQHlEZtntUJyVhNuCakcx4NaWvce92JVxEE2Qtu7Z57t
0XXCgHrWs7gzEyNAaApzVH6bKu/Zs2ixX4ozOCxHIR//mxV19+qQYIYsX1o28vUF
LvZYOzCTDESyytGeY/UtarxZB7/e5A3ISkhAVlTnWixKQggrtJiz5JQXoF7a4ueO
gG9N1XRoPWh0OVdQNhxcTzPaqJFyiUeFa/yQxVS7cD+SN31uxtzFAS0yLf4YsCpf
Yo6lWWsnz7OkiW6HeFQsSOPGpVTDLv9doOYcdlEoze283gNzexCv54RXpFuXnK3z
PyeBUG/wjr77IMlzBpqJvV2lYLA2hWyWJo4GFCsJGxLLC6TTG6qOssjgd/y8J8tL
fJDWW6D8YBpDpalAH7T56mJDjGGtgG8BZfUuRQpbjnf7Ih/6I3Wy/cLf5vIJD+dy
xyhe/u/lVvIWdnlOtATpc3tx6wSLM719Ymm29xd4gECC0BOn+hN9keQcrp5LVNp5
r1MBY44jKmLszSxwXVUE6ekpfbaPgHfRkSLMPeLhoswVfHkRViBn+23sWcv6w2Fj
nZgOrjK7QDANATQDddhnu322nCt7ONNNdKARsfnRMd1Bwzwr3BiFZ2XTUnrXLvqS
3U28zmYWFVTEsMk9NCvksGPopk7bvgbZvrTjRuZSXve4hx5BI8vT1qZWeSPG3QQL
fg+Ue7q8c6rD28YoMSFG/6ICdhBvAvMEKrVqQq++FmoeLCQlXw79N+PGgZidNjtf
Kab6TaFZ6+q0NDPuhBq0jQp+AS+X6f+tSH3M/A7kf85nBo+6nhwO4sPbuscr9DjK
R3pJM7f/yy0MZDKK1N/zCFbWMCx3S2IkPPh+4CUmX7wggvo/atcanhjLLQe98JkW
8I9PwbbP81T7RmKq0uAsX2aCmggPIz3tfrNVTVe4hEBQjRA8ujDpb/VGptNNlc84
lywVqYC8DYAHX3HmG8McCpx04yJQJ6ZaKT0SiqMrZANFyck61mjk9Mj+3hRQFNSQ
yY3c+jdCD/Ov3PlfCWmU+P0+4EqiQNQeMTU/DXlRSu6y/vSc45RK6C747/G7qK9h
7SuQ5fMdLdDfRMuGajzPe9q8/2dLEOrT46jkt60F3Oij/CF7sXQolu48IwUBDUEA
1FvAlPWnCfn8fTkdQnocRjE+CdzX1P4EgQQcQ3Dxd8QumcGt3eg3cFHABHOqdzxb
mE0dzOK6fVgxaPbZEXn97odZyVW5Od8JEDSpMAy+MjqIco0ag/UdlhiwiZONpvbP
wI/k+Hc8wHpkKO9/IgBmmNuiABEuaDxN3PfMrutM/wbz8ISuCXQK7uYhi2KV/CkB
rYTa1kSB7WnTfMCRj+tJ/msPsJVPH6wxJdtpPzQLO9Ma54vK0NjW87TBKnw3/dAk
BepZ02HU9gBDPP3QByaQRyMYwGe6+NlLt/zZjFHxZVdm2aW2Fl2nzgh7p7FtqXBk
F5zHezqiqTuXruc48Lnfrw5m0pZDGvvxj2Y67Qbt9xDSNb0+Oy+xAFsBgZzbM8Z6
nY81H0L3FizOHDx19Y2RyxpcJNngrc37dvUjKIHqe8epatNhIN2WPVJitflHAzC/
Ij22oeAWu5J0pkt11+ip+cWe4WPFDMtMAjIwZwtHhTUCcNiLs9OPoC38Vxrf35A9
fpnd2gCznQ5Si4cjl85cjgLAzSRp3LNt+b7/eKHD3MdWIID27w3u/tb2gHdBNYyq
yYVxkQQCr9FtOxnQYQjgKgW5vpTe+QlMe8e+AGt7KCHsV7rf1Kqm7uPeTty5fGKx
3PGvRhEhaTLQIJ2whKd5aJ9375DgZUXfVuzmR/Ltz2+p2MX2rG4KZm9VXRauitZm
r43HEnE/lGs03GPJOw7cLaJgAczj/G5inI2txtCQejg25/C43lCJh4MNq5ZWdwgH
f9tW+4tdyJpH1cQRw8UkXvZDLpf3zBI8ZWw8J3nGU/anWi+u5s5o6u4hLYbLSkVD
cYxrx3YEetxt4GkNrKNZ2HUl5VUivopf/ARQ16n7C9uS1ve0V/Xo1ew5iz/p/PJu
lGVK2ehVOChGZdr1tRofDyCQXKCkeKOUZM9sh/uuIaAB+8ikbtQDL4EwPk7jCg9y
G+7R0eTdx59RMcUOwCOuDZv/Eiat+C6BYbsCRAgtBoY3GQaWWSz9KSKSaQlGm5Pq
h+NyYydRM3dMJ1KR2p8wk/OqgjvmwaumCP/vd/SKmvTj/ZHQESX6a3pvlZujAT82
o3HqJOBTrH80v25BL4dox3yQ4gok6VSgKigfXoDhQ4wQcG57EV9BpsWaO1OHENlY
edyUnGLs1whvmP+6IUpZRW2chrjSj5g+6ELnsl3tLCvLLxtyXRQjD1c8X9IgxqHK
P7/u4KzGZ5NZNL4GDWd3LkBqvlRmZlkQGAXjQ+x7KKW8RV2UKkTgjd+eY9a+Cfep
TCmMRbvsN3STqWbreXOIcaGx1xwo8y++0VysjuRwoKTwBIb+6AanTcF4DdKG6dO2
SlCRByBL6h99eY79Zysh1ZJ7yX0pzci8g8+KrkOCsrs9lnB9fav1zM6BAMXLBPfL
0X/BLWFxmCrasN8/boSbjs6xNgDQCrglINkgtb1LP6rBYmbhQ9iIUwBvWYHVsF4E
VA/PovZral00e65mjC+rjvUqquPjIvdFEoxW954rjWQFKSdXo+xB6Pvx7Ve4Cxlx
GOdcBk6p3HTXrJUfHPwIV/ZufAg51Gu83uudLJyO9p/qvEXEnNmE5OCrjMw1j4bd
IWhHG7A0j/0CdhFz1aMgXjB+s2khvVKLDwBNka7I0Fu1IREisBhsLeEYtaNbJ0Pm
nbqe6Q84243ncBWqLTNx+jWtCyeoD956AtAV5G3k4PGdlV0mlCTb/dBAr6yaoyRn
4Yzh/04qt/sdOpvGsCFWm5a5O1Vf4GufgAYMqA+D+9UhrhzH1F8+5P/cFJAHV0Ov
RGbmtTIKkYeD/1ZoM5Pczk++8Gzr8M4g+h4F5xBPjiuJlfIhRXeS1F2nRiFFsPHL
zc0fzRRlKg6gNzgf25oNIIxhZimXz3BGRzvC6/YAhSFxxpHLbrsfe8EEirMCoEZx
k3JBPPwt8rJZDBkJ45EzZA8uscAtot9zkGilYfjgi4y+aCydV2DVGI0L7s1hWawn
BnOYkvlGcaUPEPd9Wtu1MbYQditOZOaABVuNPK2EEZgJmkoNsJqAqys9grsBFn7I
uVaR0XdYCW6LTSY7XS4z6/l9rAcsn+y2XPwnyZoQ00GTTSDim/bpvg5EGfvqRtIH
jusAkK3++HzauoMXiu4dZHl6hoKJH2JmzcPc1essVkZQlihlA3/Mqx+D7qFSN1cU
yhcz+IEXAGj0pmRTNs8BRenazUO4BxulmzCSQJpHXeJS8WHTG2Xw8FV27ZWAh6U+
gdXjEeiE5Bi3YgMAt9ljX/gK8p5D62JBvZwib9BoXbQUlz0TV1x5muPliVEgYE26
tnXced4QWwZIBb4r+lssIQXZiKcO/HWQagy2ObHZs5uMxqpYB5jYYmS+kEVyTYEM
5hllwtLP9dkuxS6GQ0LGXyH+T/fvoaEnDJmk3dOEy3fmJWrTt5FCVj0wgqxQywDk
P4OYLO8jg3QVOFJkR7nUmo/JKs4dmNnCGV7tjHYbvHIv8u4eKax0SyaQ59faFHJu
NlEDDeceDBn9sy2lK6hjDEOkECzoX13p0MFyBf1aBbDX/fik2CkpT+NK8PgQCJqc
aDxw3wNITJOkx+oLobJ/9COFwZPuz3tkDJUKRpasKBoXrA/69U5ytNg7ViVHvKqu
wpdd87eR8HjXCntwnp4mdLYuFUyYonMqpllHQuEaAqbPRGaAYx+el0/fUlCLn83k
VvL6Ymbogq+3udFkKpBBNLiCGs2qw9+PUSifmUwPuinlKPKfzTmKddlUYXEVEMcV
ckY/NHBsCRXPFIo9wimw/IHzY/9ifobIm/1ZkHVV+pyvimQc95s8cYxBaRwNKXiY
ymjyaG6rAfyCWhPbdgnquk49fNGfQwUqgxxD+nLyKY124NgvN7RyO5AUXW8WK03k
Un9xX78sDmUcOFDdhyVzg9RLU3Wz9sQowOrUvDC6ViGlGu7VXt8nzpMq3KoaPzfT
vCkag0OVCDGcgu0v6NV5p6Glcy5tuW/TVORsk1YP1hH/tHfqM6FJsWl5BKMhPGo5
h+P6BMX6VJc1DlfwzaGxg0sN2dOrMdYKeP95JEfhIaCSzV9Gsn/mS2hyAvKjN14T
UJIiIFs+tFUM4ejJRNo1vHMNEdrLBAXwZvIbtpJS/HHRhvwiVi8Wj4BIlxSpKMeP
Av0yRk/zpLxTfawE45pjtMb/ELgWvzLhaDMciM8lT1C2iDJ8ichu9DkYtrMUhWtr
JN+OaLRw9Q6yYvDvlrygYqyj220IcIBj/Qg627mD1ihmwEve2y8gOxSnXfmwpBs8
VVqZovxAWwOMDDycyUVBwLxSPoMIkiUMRIMkV5O6BIX15z3Wlmqts6oTzvKAF7ZL
cJxDdlwvWQOl4Dpoyc1tLWPuAl4iV1vq7Y8SCZA709WiKRF/WGk4of9uDsFsjdqB
15C0FPzetbxE7KNAHo7qVl9oJuP7AkcV4KAuNWKO7EU38bZHmaelnKqzEQCOWKvG
1A/A4FvS/c8eXozH0C2E8/ONUz6WtsHVAggBUXahtY+Hl3vVifaXN2x2heeSmr1V
a0h64wn1leiZB4RNGZvC9Ho7rk+qaVC0UsFIXWf6YBBsBV7SSkxge3sKufKVbuEQ
vdI50rB7LLeXwpCXS2uGQGOIQ5enTV8pH2MmDoeuE6T3aNb3+sVK+iUwr0aLyGMX
vPN1WvgowbfDka4xC9Ps6UF/l5d25FxdJm7xIito32ChRSBxaXqUTkIKWXkRdEx4
FcniNfI7hmwTS3dMaa3IDS5JzejIbaLE/5VhcNoip0ZZy06SrHtR/dMY7pHrUg9F
8GrpImFrkfOjbuBgWWRsnuNB1R+zmZaKYMcBjfOL2nWyPkya/uP1dhAIOyDMnkbA
vt3yk1Rbb/B+WdUSwwL1z1jbu8OLW/px6M1OTO8lKX3GjhWgXffVo9wORxaEROUm
CZNAHSAKgT8394UHCHcdoUwjpz3m9jC8UtTHqZ6sKP7JVjiN7olpAJcvv5GbNcUG
kENg/dPHxWVurTQYIv0ye0Yy3QBp5fHCJqBkCsPthmh6eabnQc8jMXZI4arFAzqM
jRXCXd8cvuf5ps94uDSSVMpAhoC6nuUmJsMWnKtiLI87IdEOMQvisGrmp/VVHXg/
LZaJGaCMDJ6ZTKSB3G9vyeuo2PESsUUbkP8kKjWbBI9d8w4L4k9LaP0DpgXl4QFQ
1rMZoXqpsAyzZrjBSQ2f1PWDNwRZ4J/I0/0pUq/OJrSGJK6Yjul6I0bT12Mj3H1L
qIZL+z/hKNB2ET9hpoByCva6UMUUjjruJ+sq7NZ7+Q7FmeneB1WHl9Qds3Zmizx/
i1kA6UDqCnFn5VuGTylkJb3WvmXdfxQC7Wljv4Xb+9kjrx9nWT4lF9PYyA30gMJ5
dqFl+hFwog9h8tRjiD1jtFmt9f3dM83atVLNegEAbprZspRgs7g/Ww75dcjE/gWS
NORg8ne+WHVo2nZXdd1FTeXDEQPUImXGY8aOboX98WwZGS+MSarY90mWwxH5iV44
jcdmJULwWQ24ws5NKuX4T65QV8GmY/tCyafKBZyY1l8sp6RZrwa/lrunPghmta0I
Jhs6mp2tDu6ases6Y0aHhlPx2bzGJzvQjcb8RGOEW3aymtBahTSzyfsmiWbq2Deg
rsjafHXUUGhhDB8uUhIi/7tkp1C1iV8HWA/0W2q7m86RFWR+Ww4Y8x2XMZf6gZGZ
mFtLjQ882E6itO0rIOXgqigQOOaGzPC3Tx4ZW3ARWaSUodXVzzDCZYo+TBMDEMGf
Nvgrzx0zBUIWZDoOeOJyX/TOJH3yU9e+qFL2D79JP8sCjs+4W/bcXPCpYKEHZqhO
jAZKcZnjgnqRGuTJ3K4oLTvWOdxF8MjFvOgYsdBi3YFtEKfJynUBw8smUbaxhugD
0qflymQWP0eA9vvHx+VSDb4h/u/pAfERvVBq/JaMhq7O5jKCf5826f92JQUN2Vu2
Wjod2EYuJrjdjq8YoKb7VH/IXxOTU4cMrp8QLlwLR/UmcqpYixXZSX1JkunJYME9
PKtfv1AflqL09KHmgWEYgms3ZX69mmqaXOJsVJGAWoJB/us4iZEpbF2NxppaqEC4
MrASxv7adEtkPS5oH3vAVx6xTlc1evodVBZhOSxOL+oxngFgVV+fM1MhZbMzgDL3
alYZjQIdIMK4cRQph2rw53jV5TGa+qyfH9JhhXFJGsrdidH8+qIMZx4f4HT3Awst
CIgQKQX2ulxorRaau8lrTvLalM9T1Di7OVK2cIo6X/HNgwFRCegl/J7t1STb4ywS
QqMM96esYkl85qEZH2609ybYdzC9o5H6VhTQBfdxyCyd2FrZkaT1T+edLx5TSGwk
cY1k0eHYOFob80S0Vhks8/KmHPjWIZz5wKYmuTQpjKAk1szTClcr1cAEE3eHL5Lv
NxmQcx81cYEM40gJj8nGJj/RKHGoBuyQTZdX3K0Pr+chTyLUvlag/hG9cUbnOa+5
jUmcN2ZWr3Qk5ERd+UiYNpwi5kJsuNNjMzG6dM0PF9s+qyugSbBJ64msXmmlkTeb
oz8M1Cay2R0VuV3RoE9ovD+qWcrx/zjF7VF08+uGZv5EqmVAM2nmMY1OCyYPnpqk
LmWEEI1r43JzHyMNgLs9d9ux+o63Wu4ixTsxwDYE5bB2i5lS9AYOJAKhgfNPNft3
ZwQcVa/giy7Z/kfsWJ/qBBdeKlIfYIV0+WsCzNj86o82ofRlhAwFB4igBgXkr9gQ
6KKDb6yhXAFMdFO5es2nWa3ZwTtmqYwwBW5rPBkOfVxd+2l8ad1sCDyUJ7T18GWT
gqxRKvW7vXZrnp0gZ1FRICgAA/pLJzJG1jWJKZhfrsA5ZgMldgAJqkoJLu+WgRmH
NQDYhtzLcwhsWqbt0zPO180nHAgv1F9NTyXa7risgbc4dVFjtg1oDYtL+qIElg53
VTjIzSh5SDbiuWBbzlnGkmyrV3RhrFOTRpi6WbNyFF5E+HKjCY0j1m+LjkST7AFb
NytOMD0LGuzQY5YL8pjP4mG0bFkq8nk4XrMZqAJez+k+nShDRZz6hlWdnjBgQ+mQ
Hh8khxxMvCLRth4Uib4GtIzmSoDTmMQqJ3/U4Ayu4KYU+CiqLvQmPNn+vONVGdGI
wD707Rx16XKPmZtRYneRzc7m1QL7H9Q3nOCSg+ehcizo/DpBzd4iO7nMBqWaJO3c
icVNTprWLzCGs0MQ8MY5yVu10bAf0U5dB0lDdhK7H6nRuTco+hxABnqr/ssazTfy
qZ+hSjQYeGQ7EU7lHfkY069tc+h7jOYUlWHa7Pqjbsns7P32qMwWYNsg4F42Y82O
Cl2sXpHGUbuNRGAj7gSpVI2CUcmR0IL6yRpmo+TY0MrD4S7VY4UMmDG7qg4PyHUQ
TOvi4Ob1deLQa+inYadyX1GLsFIRJL2o7hhtlhdtzTXhrmr6o8HcfrzfriWofmv3
4fOggld73guk8lfavPgjLpH1tbBsUNY3D2SoLigBghuZncu18eUslve4iK9KP5Sr
NfaaQgdlhVWcs60hrA4TsYJDv+G1MqmqHyGAY2NkJ+G900uytE1ziaZj37g2897b
Tuk4gP3fHAE3vV7cnZxcKMZLAZxrm/7q56TmZDxbIBqogUzx4iQEDcX/YWD22QVl
a1dzLTOU6IV9crfhFtUikvduGc2Y48BviyLOIG0GBTGv31XeGQSJtLO6Dla4sgnO
ZfGfLd3enia4BUcM2E8arBqDgZPh+K+Wu7bADtjdyC2uypOv0/m08xshfMLJKQFc
s6CWWrJ0orXu/JgYAEsch5sx0vK++R944wNbiXt4UD67VnysgemM8oA7z+MAPeey
aJTO3MitbrNaM0RKUE661fV03J6FZsh++AfsNis3CTleVViCxXI/wD+liRwDBJeg
vGJcfP0Vcvl9JvuwwP9+PL27/SImvPEPuMsmdke/DLotBatGxhC2sw6BxZSEmjRD
j19fWWvDgEHYx/nh+7tqEtBOxvNVMYY/hIKPK7Q+AqXei6dN/2m2A+yG6Pp9q01V
05XekF3UZmgl71M9gbDsLYiypPlGi84LNqbrqVlrJJjAsUcVfE5mJhrBhjGntFrz
knTzho1zT126rV8TSCerMHAgHkmwbgbx+WEoRsMLcWBI9ufetLXjVZcWSUhsWW7h
O4xi1YU4uyuRkSS70DoYpu8Ck05H4HxByAL6fAO4cNLyiQ+BbxL5JeyCjdZMZj8F
/M3ucBR/kn0SWni8qQ4u+i9GC5Hqtf39YISMw6F1E+G1jz5vkWRoa0Etm9Vh30kl
tAxWKHoPVeZjb9d+VQa9uYYUKAvDqzmsgxWzG30HJyMei+DQaZY+4PhACne6k4es
H0lPzieUMR2I/tmolpXScOEzEmJOk12ayGOAt83iFCv5C3WR3X4cCIpkwhrrwJBl
7DRjC3QsddyKJZ/K2vcdZ0rKmrgILlo6Ju9SojFJXvYwmyPm3KOUJhFbobEiXXAS
cAbTt3Ei9iMUm4jKYtsV+iO4W5PWkjbCwQm8sa5kND1qU+X1uDjVv8vu3QqAfRda
ibidu71pFWxEY7kzMDsMn7ifVg9ls6mEWzjymMyjhVKCLbvRC3rrARgpqH4l+MSP
swST49etWm/Ik8IKT7nuLX2RYigHqedQJdVu+geiizJYIPD1+1cuRgEHijGBNSDY
nD7DVL33T76kVvCtrm1+/8dRgmqx+XLxlPrTTSPxM/v0n69eC6NG9gh5Bz9D3UU4
kkiMUr0xERhsloOB/OKsIjWsVHTf7xem11ji+HydA3drP6KiB3xfrZsithj1ZuKI
Y58QIWJo/2uZjQG8cv7FqTrhq6WYUxsyhxQbpr8a/fHAV2CN1jpDVLBL8dWPCt9u
MRUJk0IGYUifviSBynASwWTerkAcKwCbHGzTpma1uFp4/dXha6sLC9YYAHOOkhly
l6lk/ec6yLOCzLQib93yro9BVxo1aHdhFz7CIPT6LBTHTz/G1S8mdB+VBH/e0dYr
8MDYGgExW6a32q8P2bBCyUzmUryGoQbiGyXOkgIAQkuorTrUi+JFR+TOtdMwA2yN
XFPJFzbqwpYf/FuNIkGP9RDANYWrP5hE+fl8h30CD6Jes90tYaJ6JnBsLFHr+9hs
CpWBLER6S40W9j4OwGdr0qJ2ffDj8mM8L3dvJrjpbiaquo/PRHLonYP85e+AJvg0
NyT7JMzom7f31u9MItDP5+t2+h70agc1Z8ggvIm8tjg4+MGFYvZz3RxNWZYUux9P
p+499qtcnVlYX51xUIVDo9OiEBNIsXgm1V5+zfEU/YLUdBAIL3gB04Xi5oTUYvNY
DZHF8QfTLjBfyIrkLikNV3H7byXdaG8UUauyWS9354dPw/rUi/DZoMmtllAsf4li
pnIpJi/zx+UiNdKejVo4Vu9u1rHY2i3gL/UzCZxy15+aUcMrQgI126eyhNU39GiZ
J1wBUgDnC6Mi+X0pnp4jNaW1ZcIGzKz3h3dcq9EY5EvldtJzznNakheSWzg/BMQ8
TO4HI5WrpOdwSt0aDnon7KvYsiHRa8P0ID3cNdoOWUL76OCS1qhqGiXdpIik4AKs
QCbgN78IZ9ChRlzpat/FNcPgWE6o39bWkbPd3+hsFyuddXdmcYAEl6y8peE0c5qO
N63v2AA/CATipquIBXdlaoVN72eK+iV6B+Bg1pF5HO9Q4rss8KJyM+EtNNmfX1W/
OLNoHp7gctfgPOF1zfTw2OA1HnnvUIqvP1Mwh7GIleeYxhQEOU2flW5J9wmVLcnI
ZxsYYuwubiqW2QGrkLRCZS3Bd38ejxIjdnKZRVeVhd4W8Ko3NlNWuHS8aixt4rWA
8QF0Vp5xqLDlfvQ3rQ+e5vZjm7zC0tHVSdDWkN9wXlBto0aFB2dLhufv3U0DslIu
KQz29LAzH7pMpsjOlZQe6jv5ucTeQ++NORHEZh6TN2i7K1Q40LXA15QhRgw28hfa
a1HRMUh3nYKyKILRwLJ9IeFfdCLJYp9Y3CX5UAvVUWmD+ARCAHlWBNuGewN4tpG0
MEA1MV1Kf3kCQG+ySwqcWvWL5vSzw5RqcJ+eP4IMSmwzgG4vimIiELa/Yyluvrju
OCedC86Et8Kvc6zTOYITnvfzNAvmh4z5Y8F6p2hTUKBdQo80WCiHvRKe8EvfbRta
LG2yiBiHi3OqQY8i7OScLd1aOOfW6iFQ6JyQ4gmYSE1esWIycrDgVtvtjZLMGb8Y
1Yvn/rYGnucsspGBWmvXOjPh7jbIalj58FlRoQh8aSpw92OGzuUn0Ky0JHIs/a80
xsR7rt+VuIxxrrU1p9jFqbT+/Dtki7krqfjDDM4Xnz+PoZsDSGVpv3F8q5ZsapAb
utAEZDi8EjAj891bfbCS1nYUqCRypwkjSoKk1UDprWpfcpJpn4Lj8BBnMJznPa1u
IWjUVjhugDAkojYTITPewuh0AV1K4MLSsDHElQlI9wqKo5KouhRyhH6DtFgfwcTy
992xbsYWSbFcuCReTQzysU9JDsjLvbHlhTiDWTSxl8Y67gzmkhb2b8vTo+Z+9ghG
mrv6ME3Y0evj3FUy47tcev+xGjOvadM5Q5/t1H6oqW3amGhcp76NnjFy0qiffiyf
o/QrjWAg6QOXHg1aT/LdyvfLn1qA/Xak9FbpFfgcZx9yVlWowAOIhjUcazvw8xLN
w1pKVLRxsXhYY8MfFNhjFqi7ip+GrBOvLHnscF4KYAuFUg0RUu8SJb7zlUw3Wvhp
K+SiFXyahQ4Alvjc6zeKbhPuFId3CfGwiohMm6mzWdiNdHBaikLX8Lh6w43ERuf5
bG9UlTZk4c9mObpf1r0PkzirJdgrS4rNO6U6ns0ju83PFrZQTP5uHJdvpK4Ae5IX
ItYzu2BmnRvJk4Qu04dFPu34B1fH2byLzK0Hof7w5gbi+mmIXba4Sl4n5UdQZXWm
qAySceVdiRqOzUtlk6Uss+EJ3IBp7/9DDQ8zd0Vwnc9PUl9xGr38OuGyfgfg+TUV
J3JreWKvxnXrD15AjgIx5GhA3ktxeG8mPN4MIKSMDX8YdKoaQu0Y+6vP0JJPpCwL
1iCjAUx27Xn0xDW8bu7ZrN8Dw3JOilgS7LthlSZIrPZ7s1WkI+dGprqZcXHsadHU
1LpnTc1ybTtD59pjhtuW29e4HA5BV2jniwKdHP2lEsg6nlAclrotH/FrOqGGxW1z
0ElhkiyojY38MVdW9XFC1jD5QAzbpEH1EEWFKjkPX2ejkHd162Hw1yAOFDC3PzFB
DzfIbzK9/VRAMKjCkGy5pX1AxnDo89rwdazXwDJ5uvi+vf+BXKfEP0dGqRerJsvN
tNQo1Hwge4//L/i3I/c7Imdw1IjBRiqvoUnBY4ds4OjuS4iq03NfEpF0dcrD9pUW
WSK9kKbe6pN69dicQC+ABEnum9xr7AWbsROSxcq/JqBYVr1+EJZgiPFZMkbPNdoG
KKVMXFym1r4UIaq22RmpRj+OZ0o5Lde0Z1dTbiPESdT5y8MjvJ0zWQ0QerqnB9Fo
WUsE5T12TQV3PztnOmS5Zt19x9VuSGwLpB/NanbWoPXuH0BNsVX40k85arYLPAPv
JFc156iUaOkSLqMEjRnwvT/aL3HyIy8usj93hW34uep+HmyFSQWuqIBUy7MZXxZR
tunEmj1u9KdXDYjPvNdFfRs8GfQGsEmXFkeMscFEg8cFM8o1jooV0G6LnAj/0Y5N
oEkUwU9DgGbLnUiPHNRdP1mbIb3Gy64LTwtADulZBz919EpQIn/lPbfm9IhnBgN6
tJO5bauwRoVJvrAdl7RVo4NFbXDxk1X3x3aKdlUWnQPLOEDpbW4ARlNVI1M78oM6
2PxWOTV5l5wa8Z2Vv8dP0IOaUcwTvvBXxh3VB5iBh34xFRLzhJINGr3LO0OpiUri
a6fhYnsKg8lNH+A66h6+kH7CGSZf/rTx0Pf4AgsM0mkgwLeuaWSmiF26OIfmSp23
4OSiNRw2S+iMpemUe8K1ZysKGqRa7YDi2tUQE70Sb++QwHrjB4EpBrd0wnpevOr5
ODWWbVo1vVghVC8RduaBTGhTETwoZcpS0c/65Ymx69g06xbfAx7oR2XbX2gmTbqn
8iB8tpfLbbLX1tLziRSc9NAoYa6FqDONZhSbEUur74h1DdUj1CQe+rHWIFo6uYDS
UTYVRZ2wbDn4Bqop9N5CGJN+rE1l3A+yZrdOdRxhQJKriqMTBgWffRgUiLRAPx+6
8a+ajXR9lI1GCqoQB+Wh/zS/ORZ5W9cjuZuIaOo6wQsQMBDNiDY9pMHmvARMezJr
LW6rzBRx5jil9H3xW36DUY/luGqEmz8HEL5ubmjNS8aLzullCjOW/Br4zz8W27zb
kwN7f8LceDr7jTTf4PrIGO3pEWGsdCFg4V5U/ITxs0Un7QShaUSa2ICMDljH0ARa
xYW6ejGRiC0OIkH1ObR86b5Y0/qxELFQl8aeRaTFE0fUuIxFLyWklXDSmhAvAi4+
8O1sKYAfVn/JCRBtJbTX0D47pVGpmH3jY7iujv6LZSwO84FmffKtwbaqgDRUnSWT
4jZYqefKZxrmk1xWIjHKkbuYZtrmrG+v36+z6fi/BH5B3tJqXuocSN3tiCm5tAVC
xRp6mwsAlSCHaxB3tFL64Iy9mqaFIPlt2/Uxk1e+umO6xeJ3uD6PsYtYsVtXwe6+
6XwX6f9qk4wFg1nq2G/Qcg51yb5kKtOwnRY5zgAj1mLKhVksO56/iXlfXWJVB9ls
QSsDWCFUsPx4cPqKB8AVCO0m6VtLoRMuHOiDUoRLcJYOaTwx1Y2o/c4juKpH7Q8G
ytSBvVJPgC6F/F74pGZa+r/N2Hh//q9/PGqOtKpkJzPAK/Mbqa/qMSjXkV+DuFcZ
Gc/jczmPg+PFStmHTrvxrRGa+p7rCFXwl0caRVs6Ywx8koEhdTfKbxNc28++RsSg
AGzdI/+NyTz3SEr8PdxcCJWewoCDdmmnyqQCAk2geoa0d430YzuYw0rIMTS+I37g
IQBYQ2+ZZFzDMQIuForakyS29VQXzIVxhv9KE/1ee02r1cn9u3hhjgJdZxVmFQH4
uX4t5Bz+z0QDLJhBuiqo2JUK/wOtpTfa9HE+9tpvji6Jy8FkLoMhWsl85KOXdF4C
TLuLgDsg546nGtNtGFxhBJ5nsnUkJX2O8DRQOZWz8uMpCWu2ahZcnuvhyCQjHB+z
ozt/gtKHDVlMgeWSto9JUoMrwd1PzQkf6hhCYC2+N7mTP+EFbwkFQRuWCmwWHsKI
CdwJBz6lK18p4FqI2h3byhxf0aum9iOGkMcvURZBofX7+DlypztdRsjg58YXWHjB
iwdmYq/oUyiuDmsIeRf9kT6jVrrKPBvzXgSa1iQiHUFqZwJdfXA6rzBHKt2769uC
jB8GiJcES9p4FUZAvzMcDxu/unkdd8vh333CaF4gkHEnSIq4D4XUiLSS4HOSdov6
bWR0anS04R7hRMgfHBHiBM/i0ZEoo2E+7cv1aMY52ztHnqdq8Ub7Aid2AGNgolG3
hzMYFt7uOCGvszV3sa84WNfSw/LYla+2sxNDGbAU7yUK6D3VqZWlekTjxEyOQbng
4M3iAiACroWXZm0+LV1HQRI23gVNmJ4xsebri1cBR94E1cF9vmReuCmA88hnPV/E
c3IjMjM86nr7aObUwZsFDNMYtirKeOgcqL2/jDOWHo2h53Yqt+zbBupVrkNUVSTI
WM5MaXktr7SuRFj15WQtmpdaNb8PecsE8sRMkdIBihO1ENwiWf90LWQ2h2Czai4T
Q4KTD0eWIv57zsm87qNzeLe1GVCQP9YSroNHb474XTNR7SSSNv3hD/IjQ9mhKWuK
DJBYLveDhuHhyB/TCq1Vnew3UltxtVa6U9HhTtVNiu2pngEzIWfm5PXG0ep0BHle
V3pFU+kC55LzaHJlWMePVmNwBE7NUj1sTylIooC64BKI7yruUhBLrssk9wLHfY/1
OCBsOfksJYkA7JfoxkgloY/2t8v4G7p/9MQNjyoPzJQm/5+sOZ3OpV6Nvi07om1Y
rCLDySt1gW90JYUtgrh2YAiSTBtfibn2YnJ5yB6TPHdUIZ7aHQ5a7od9GLIhx7QP
WFKTGYjOJCYGY7SqLnvCyg4CgitK4lHEijd0Tttu9DumO71sOl9g9w8RZoT+JsLc
/T+H2K7W0tcQ19z2TbY00QrR+ZU31WkT/ylIeX8ukZm45N1nqWTGZXF/8Xqzgaow
i1Ng6ItwB02fKx5PcC+z7lSeagvGOJu0sIEW/Xjk4xI7D+3sxkT2kznMOvR6Tb/Z
M9tzNk29O5eTrdBjK2cko3hP79bZO0MqURPxuZRgriUq0NUCuuPsSkG83R1A7ZMc
uKgIRqYiARa1Gy/GLH29EZzYQdqjCTyNFxSAIAcYG73NFmX40tJb9AxsZwTABtAh
8auEGs/19ahtXLcSF9TIGQRhT7kwqEjGgH3N8UJgIjbXPrZme9501Fxl6nQ2SDkw
AeGMUk6JndfFaz7ILKeYYtTRUt7e1qhpZlIw3GbvJ02800WVeMuZ9qyEUf10z4gA
QD1tHIA1ErygH9q59ll63YlSRtw9j7ngtFEhwCGeaxEgg8k3UFR4ycgaqlgb1P45
pwKis2UoPow2tLEfuU9Te2bIE+QBzgzC7U3s/yHaIIE3JaeGiBe7LznklocxOyBS
exmdtlDbda27IeP/QZ+PtkoVLlVbeX99Uctg7dfCO026rZaCV/851jPwvJCUtNdI
f80Sjr5QWcJRFpxql+Mr1LlLqdqolserS1Jq2nnaztKFsoWGCwuXxjmJ7PAxI44y
a0IAKVGg5+lHejt9SFZUyKr+4tZY52tbgF39I8kTHBmgbSyVVdQXjYx8EcenOhkl
9JtE+dPMtyMArAGryfEuV8g/WCB6Xvq8CqPTa4cFAVEfB+2Nl8h59Ob/RIUc05D3
8GJ2RFr4DygWpUpzUeOutwvaQMN5kdDP7rZrTbFZXaL0wr4m2ZTBTgJO27IYrAm6
sUhPaGCIB7m1/dKlUXeCr7xpUxfojMmezWcgh8ysQvbJCR+pYOigFq+taPDguXGK
OhXMu7y3t98dyUITKfuNJ0n8PTX9bcvi1b0gvISoj/nL0gW1GwmgJlbinhaFc8iR
cIu1FBmfw7z1Gxa+pTy3UJduRMUHGO70DQQ/X4thLiHMb4HBb5105ZsYJx/HUSM+
902LgPVtVzsewFP0e24UKHISX/n2Xx0bmq/iNgg5XhCgTm1S+OSt0StiJPzWfIka
lDt0FvsqkT+JDrr3eTP+vO6f9XrhCJnZVWEd2DWnV+5yHdv+ByfE+Q6npt1fGf/U
bpdSDLKZYMKrqGW94KPuqef7BqHe5CxtCuOD8ha6JM2CHzKdt0htKlLCb+aZ7x9g
mf/zwID+ombI4bZVqzTMiHPjqOfuM+uIJFPBmzq5i6YC4Cs6zYIWctkjKC4ms5VG
4q+/LtagsCe/hDKywAvQ832fAI+/Y0u6joptWoYdRfd17xSOcIlSzsQTsQJvLyQ7
q2k20b9JybyksR64M8qjE7YeiEJhq0bZiwckHh+3HWTPCjH/gC4Iey3IbVH0g5ut
EhdYWq1Z0+0MwPow3nnQUBJ6uZLJJHeAoEXKUOK3f/hmkqpplaUrM9r9fQGtgqft
lGna/NecD7JK7381Sn6VAm8qFc/rFeV/RyctcpXTXao/4yEZKAnl6ew318Z3E2iW
t9ltqixLcXHcdZJH3lZeuNx4lK8NPwOHGa9yAcvIJpv2b6ofvC7PeHPGFnpSdjD5
R+pDsPshxQjPL4vut2JfV+yrLBGN5j7y/HZUdXJEwzdKy0lnFzKZwNJpExbJ0Ibl
rCc4abipjgKESjPgTxl6EWEv54Yx38Z7uku20D8IZ8XK1g0PvVwl5Nn97wvR1D/n
27HJpmILCjSHl+3grAS3OHIm989Fjmd79FG1jEZM74IUxooLiCz9wLJCEhD4hpg9
sp4NZgO5uTehIJE74463uyswDNyFPpxYpAufb1qHiPVpf3I4Dl75gHz2E45M5K4n
n2UlqxPHAuJDp3F3mm/Nr/IfipaCJq4eNv4FD+3jnr2ViZ3wuFnjHBIF+fYgtxaK
Vm2PQM6c8HZS2+0Cm0SFPmGaL8DhutBYdiaSfRWLBjoA6hUUhcGzVklF96pLLsbT
ka9OO2Jd23+s5zHM+OnUilymaz6x+sFPSMA8xOjxclvE0DP/ZX+BUO7HiYmKbLoj
DhJ/xtbmmP8MCXWutyBdXDJEw+odArM1hyVCr0LScxh90cbhyO+yho1+UcOwuGFv
8X70U/T0mI1L7vSeMa9unErvbfk+XU/JlVhSAHssALB3CneB5HddQTSlHjPKJFdd
FvVJnAWuXbAABn7Oy8xBx3dXEmWGCGeSSIcKkKIlfT7ewXt2AuPrO1+lyTyzfvXB
57VIwUgd4AwHmrvV/8LueJ9e2yCGak15vOH2buC+DRE/HPvUCbau3Bj76A7Inf7u
0RCsrhboH7itjcGfRAmO1VvuD9bTBwb1BHMBCBZ7BBgEQxcJsTs6DGZeNMsO31UN
93QP400VHfffVWsgvrIWpJMbkiJcg80rs2HjA6edfepXd2/7LW/YS1JotOB3UD11
Ce29KSaFAhzL5AOVHfPapAmRFtPOR0fwswIjtRx7tbz03tzrOO1ze8W1mfvoXb6l
RCZLCGeciqMxEnrWdsXaknmbp82+mAdQ18DuwbvdG5EP4RVz5YvrK0VLf1o7FGa5
YwOTDjs40z6TGq4wfbHM9ttK3loVGvLOC/Zutxq1BaUdjVup9MtnGvZUztqPh1zr
Eh8DKOibN0xDKOma5A5zliQlK5z58h0dfyeYltQJCq1Zwd3AfVIA8/mq7cGE7ZrX
jKKnBjxmJd0ksqZIUWBeqlhux1umFEIopVVVuSSP8B7DCvK+eHwMNEO+bwIkfJzu
6yTG9bU2ec5acHqWCF8WcvdflWMa4WQc/TRjUZMu9pYQ3vTk6YItBNhbxMqlEJuz
q/3bFVJW68uzy2jtuimyX8SYVmyZDEpnYGmZ1cn8kErjRtPhWHX37TCoToGCwlMx
IFI6eRWS3G8yXzQYdnpxTAxDPM4Qz7hDNZbJf82wrqMLfg7j+8UiqZLc89FwVus2
SLyjuaRZXL8V9bsWezk6SRwx9lCwPgvyy+KHUc9+FND8TPk8mKoO58efnpHCjsQE
XmeICxxsyNFnZsnb/hgI5+lbyb2syg84g/VnKfIzj/hGpljoLj7sHVy5zNAgzZ+N
JyNBAixKnL5Cn7UDlZn6Ge6sCUPr01rJp5M8yVlpaXOcXu1yeWGxLGBeki2tIaqX
akdMKdpyaE3F5grG8htot96KUbD3BEuBuzsh3zYfTTGc7r+nD5IuaddOLTAzG7mI
qX47vrXHdFN08TKox5MLRumLJhCGvsVagI2sO2Xh6S4jTyWKNncqDzPU/jUdSj3z
7P7NA5UIEsntZAc8Uc7s4Jmpj+6DknnZyC9BNZ141nNnuWDi/GfuRTqso900NIwU
54B3GPPukIcPLHBSUsUU8AEkDVDF39U6wLj1R7RABoD5QKFMfEcWcdrtNAam44SQ
Y59TL1Z0Z9qKShTiG9hsvZzxRGd4se7A/jvwldnUVh1gO0QD/y01b/4P4YDD9KQc
8WY2+vwwvoykQw8puTW2GtsD/j1qkivlK1klUXPysBtE3PpoisjbTuRswgBI7g+O
wf+11RL1vBnRJS7nX+/BPwLC3LpQPrL4RcukeFZRu/S208GPpAqBQGle5J8l3sgl
gO6amtc1VbCbPhZ9rQIOcu+4BIrb8WiJMQe8C6+64k47YGryX3+Z1XDQ86gAr4W5
zkjd5AZPiCv4IrsVsbJ1PcCVbEdRp4109hdfoTnBvjSW9eeHNic71iJUGR0DHhJL
hUpiQ4n8R0LpjFqTrqJPqb1FZd7gpt+YJ5VoWQaOdra8fJ1FdC0EC5S1qozGCkCO
oNAuIoncXYBkr2zeSoEqKFUi9gR1KqSB/wkX2GBTD9SMOhLpEIVOVg2s7Tocw86f
sRtgCa9+Y/GyaoGGxyJO8FfaOAEWcbixu7sR0egBMdV2dAvtbtI4JT92fkqccU0F
O3ngwrKclydCmjk/wGIlpS1tSh9ymChPkOfh9FRYThDbkHY+2T38MTeTPOTHbMBA
9NNjWvj1e79/PrFsKBUXmqIPb9HC2jBDwlRXw369z4ADsEUK7U2hqbekZAclVsX3
eoko/hH8vjqTUeuwZkU9eBsE3nrYPfQjA/WqqWSHsb6BRPoAk2+DxVY8F/6Qznnf
cx5yHTC2ieYrXn9gmLAouYLzcpF2dnMplqLZYx1lNSIXsaMCVm84TcPbkATG3lSw
+t0+CweMRsVrEiugDxgZgWxzX3h0ZjMYkM2bvpEtn0aYQnV4970nP7QxCHINiqqn
+BcgL2NQkJSf+oaOwk2UnpXsPVfQyv8BVTBUhbSledJXQz+8In2ayKrk2WKJjxJ9
AmwUsSUiDSVlAtlZ8AAcbrt+4xPmAT40BEj1hQhZklzy1ro9WWm3EooX7HjiiuXL
nJhRxvxUbfznllrMLPXq7mLAsJlwhxf9IKqfLZgVFEH5gD16g2ly427ek2P0gOaw
KUKzOdYB3zz1b2GuDEXghPocPKSRgxAiYAKSiIJ7XTjLReRbh1hSPkfaDiwROgDi
n/kG8puZBEekuFHaZrUfm/md8i71Dv5OopbePCtv/cjF8e7yVgI1ZG7akgf0+T5U
IU+V+aS3OOXskHGVcH+6E3WexzvMCE5bR+4QbVclwky/BdlFB+W9P3TNXZ/Ds4wg
tPnjRYuW1aycBZSGYg9t4T96iql487H3io4kDdNPYf7QtaXsU1B17MjbYctGpCF1
Wuv9SrBWenM1BIhLZ8OUJ1iAwYPXeo7nJW1/JhLL/4FsJ2gb/JykltPtLGfDjUxr
MBrpSkNazzkzJSPKRKPd/baPRA+sOXhvA644dUifr96osdmTYeUPIgiE6YjaORiO
2UugQtppVoPxUW18h2x1E031ESVn8tYlTbjSWF3Za8NnOq2rPXgD7ku/3qRdNq66
KfTwIcvz7Bg5yu2TdG7JZS+YRnWRdy9rKChCJI6IOb7Oz6YLww8XdsWrTbe0yNQx
2YAMegSIaBi6I7kKjyzgi4iumLJrlUym52nUnQq/iUveX57tuOIATjTFVm/YkL2a
O5Wmon8mIlxw++Cabndg5F/D7srrO9af6H9LYlmDHDqIQWW53nyhnx36235JMF7X
iRG+oytUyLJuM+9UBnwYiywM3V1gdX+OtBhYuFOu7oKw/4YfezzZAmFLq3pf7/JH
iDW6Ds4GSYb62i6U67MXOwBSBCywjqGgpYtWs+06nej/3/gfIQLebQRPzj2acxPr
IbXxXDCQHnuQmwvgkbxb4qLfKqT+zMSMD9B+kT+FD989/9ae5co0D52rVsw2x8fT
sBWP1vfB8Mhi6VAR9UCUVmMLGHOCRoXGqYqbCwUkITVRilIhiZZ1jfj5sQbOUhCP
xKAESr2Rv/MaAwehBpktM0ybherkftf4R7l0jSkxwUJe5Req6tlkSi2ZkPa19Nsm
dhHk/Vy+ouSAsC6KfSxyMWUn80Qy8hk/hCiZA5OJKNkpjXaHxF0h24f1RkpEijF9
XVkvkAdfmyK5KRkcDuAG8qTucajjpmbwfNaqFcPq2+SoaZOo/aapZOU3qVLZREtK
77bYxKkdCy/b/+2FW6hcz77eg7L/GdiaI1bDh1YZsYI3RdsFKwVd6cMo6GMwydKM
14DpuRs5qBl5ZN6UYB0vlFVF5VBudoyeUc+Umgx1VBgGulGJqLB9mkotHLEWILPm
sWStN3DI1hWOHByj2sycn96bMmVkrPq9rREoUzbnxCDlNLZvnhkBS97AUx6ZqiEl
OXPb48FWxUpxUXOTGEh1tFmZeGHu200fLybdYR62CDwhWtU0E9A3PUJqKKXKdD9J
EwUCa58NM85bh1pNZ3EkhhoPeKScnKh/XTYs3/DUz2Fot92dbVyKiz6uJc2oKnMi
XhpwzYN6e1w8B57R+KZKoLvYUxVr2QuDOc/wkMR8c5TM8DKmmG8V9aSuOJdZeLXy
HRyE/2wpniTbZ531JioMh5aGzgObnXIBdg/jk/K3Yi7QBXx5pJAXwgE7mLfiBcfk
A4hU5+dGduqBzEzAU9voPe/mVi+tK64S2XYgdSWN4i055UKecIRA+tDDEtkMFbwe
Oo0iz98Bd+X0+vY/wo5kcVImsdfiifH1g1nxp6ycz20xJsouXOfzYrgykb/4/u1E
6clqBUrY6+1k/n+Kv3b70zV3EwnZNn+EbrVQ90t8cQyRCXcsRjJBz/MydLEgb16M
dqxR+j0aUvgaptYMoT1+reLGNNK0wWNM+5jPIJ12XrHBAVHnFUwH/KXGJ7RnwMD5
RlhsI8EHkRw+huXq/26A5qVCyVqZz3FiOhLOCuGZKBAi87U5T6B868wnct5BP7ib
O7oN/yaBbAFfW4fL+W/ivRC/6ZKtkSFvZjJhWIeAB8d8vwfOT7Jhn2dUqA+7h9Kz
WBkYf7N6duq11dpdsqLe8E03GI8FLrnrdznpnNkdwCWjXAqc+SMCWO6rfCx/fgTt
Tsmfdnt+oOj3ckaT9nsO/ZnZf68NuBhXBIIY73UjZv9uZfbqRdQy34BlSahDx8ZH
73JekL/nPV65KWceJBKg0Q21ZBYa26fiWYmbjK2hiBYp9fdoG39kRtqYnXbHo1s0
ZpCGhfpOvN3cXaSrjR8VWNgoxbBKWKOKwTv/eQO66CNYYRcnyzl0xDwh/MQZasaQ
1fvdzS0tSNU/Ycix4JCLTtKaWWJ+ZTOazPA0TwkevH3fgibwVO76ScmznUdphLmm
+BG5QQ7KsUhJAEyFgwVlnewt5AGZH+CknxUrZ1LMfYqBJ5n7k0bAWqz3l7oaENJX
SZuFNOtKttB+51P4dJIwi0QlLARlfRAwCCaaBZQnaBKlP6+tjGtA3q+1xxPNQmNZ
rir3erPams5sX/SEp+wFUPGf+ekOKUAwM1vL9nmz92I8Zk2pMkWp15VuyRvXlcox
Yo1qioiEP5zPGH/X2+1c9aixkQG+ACloWnjY3dCMNPpYTKrwXoLYrPeZ1MalS5jW
p8bzYskAmyCaZYkp54Fv8fYZZEoT6xEmqM9y9GmuGbwsV+GXio4j+zuYe/ia4TdJ
QPDXXrq2Fm0nCoTwmJy0mm5PK9ROwTeVyRNEe0r6kMmxtzmtmIwIxiueyNLHryYG
zy9GzcbWb/C+dElae2XamKFDavvsPlwaY4ViFv/Ah3vLYWy9E47aV8dqc9SpwVE/
RRp1c4cB42HzloJYBu2gRGu8jUD9Dg6eFmPxTKdHFWQkznukY33YXW5ibPvtDLke
7qYliQJlfSD2n/LQZ2+Fx/fy1sq9RD/UcEZgBT1XFKnDs8McNFDhww2LwAdnODQ5
W69RyLWAJ524bCTwbdxpSZ0Gy7QPvD+vKlorrUI7MevNcXph9Tt3d80gGqjcfcoP
IzmCFZf9rvVlj8Ehh6wFwP05qMm9mGv8i15nZs15sjhyZFTafwnvQqiQaFYehIsJ
qN0UxD0NrIfig7FX3mMpBiP7vmjJ1w7GbwYWn6cmr7n3A2cGeJLjFsW+ve6KT1A4
Eisypqq6SLSaLPgXj3REej3v7ybyn/MJ5No2eEzVIMJ+/SntOY61VwQvdc/USU2z
sWzLSMe1f6W2goEF1/0S3TYeoaVwTQl1PKwaO5VITR11z/cmJBnU9nU4h55K+CM/
hRv1vuph4L6nXDbvRLmQpOgORGfVZnSe8lY0N7PCkefMKi3WvWUV1OoEz4FvjBBj
Ka8dY+FO84/qhbzgOWWQqBL00G0Ir4+9oV6EyMx8tTmNBfcY/iR37m9MVE5pG23l
BjuJiliqcqUszbjFpanZlpzFMirORnXRgs6Kh9X8kQJBZvdMSzzzw/F0NG/MjAxS
1QiSuYU/yg+hw1NKlp8dGrTWc65cD+qlg99NmHJpKB/hd4QQYbnhVfG6cKNNGaj8
R2JD0dF3YyYgw2oKfeFlgvNEdrqcv5G/HUzRYeiMs7YMtogCPKyq/GkxrmEz4+7+
5ct2z1WrYLwiT05ho/MmxH/QNHTVbPjS7da1E+mXARM4Wchi99+61wiBI/orU9gf
E7PcTpoUexr7Zp5HTOOI3CwPhSpdhP4V/H6fwmbOi95VaOd/aJi+Y+lDm1C0ZMA6
1MdmY994QmPYVQF+HfG++OdA0dNjNVnxv8jKAo1P0TU4dO3HPX93tUwtk6t29ELl
NiAaY5tIn+fHpqOo/ShWILNNk8dKkK18RR3EPNvZxt2cD6lDC8QPwt9QFvU/3ehg
nJTIw0lcdmgwWOezAMRCUV5sEhQFnOXFPY+sa+corvK2VOwJIdFI9zjtzARaHLLR
wJvGahY9/7V5/qofU5Jt3VzDgE8K1xVy2Mly+GBlxPMMHsi2rzSA3Ipa5In6neLd
oj5AZRuI4NQD9iBR0p7Y6RcgHGn96SWxQsYBAYcnV8kV+SMUIEviYiFc2VA9/ShK
xZglNMeq3P+awHDpy8KjH8tqlMu7yDI6IQNGRWwN1L8iA+BiGgHa/w8AQBSKKiqF
bGU2h15aRIvDjtK8DzyHwqROaKNyBmgty5AqUhjWEiYlI5mMuBJezTWXeg4zzb5+
43WUnf+kLF98YavM+1B/enH9+aczt+5PyFntlXOtnzFOF55ahsA/hH0dLWZp3iaV
ZSpJOIx6O3ws6HZlNfouzxHPQ1X6JwBu1Aq+5FckPSSJkB3Fzf5vspRZAD7xCsEW
TQhiFjg2yS3ffgpLLX+cBMttSA4vD4JJ0Ddw4w4tgy/6Y8o2aQgFABXug74sV+DG
vsANHfdaSfs6CSYHDnuBzlYLDoTodHzsZ+TuIqxcGcvwQncNhDWSYxICjTR+dv3Z
oo/TvpNuYnsfUPiirGSb6yDaD4ehV17jJYI89VXg4sTntqHliTajlOlnoMgGlIQ+
75Kair2eTapl3eFJe0Y5Q/N5k0ArGgAcYO6ky45QbuTQPO7EZcUbAOjfMIxerKET
mFLVPmwoCbhj7uTObSp/vd6HZE9qQbRcyA+PLhr4b/GJ8SfV+8d7ioFZ7RG1okl3
ga3zUlIIsfvP4vS4/Uzfrtfvc/FamaWjvoW4E7wZ8c73R5qkYd6XM4/EemLvJsfC
qxdTZysTE8xKJvGAL70AfviJAcNzoK7IZ7AOjcw7H4Pn2zyTByPgMXtkhUiUCyBV
dryClLJGfO95UGIda4RBXt4cFT1JYTCNuQ0i6synI9YCKcJ64M3L5jGnpcjA2B19
+XZtryuwNK6GJUoW/Dr/dgxevqSTNYSTZX0HTgrl1xSqRa+BTX6FeajLO6e8BRvJ
WKqse5g1EQFB/4yKUQpVHrz2yRuefgLTNV7wAH/LF9lA/3cIo42vMTR5V/53RTfx
GAdpv80veNBPaskdhtp7Sg2n7cknCsUlCU95i8OnOq7EbonQBDtnXdIG9lJTJS4B
tMI714zb7KDKhbN2ieuCDS/Le8ffujWixF0DejnKMu3TCQa6LcgfLrSGqg3Ra2wz
h9rhTztg+YpusIaGKTHXSdUa3fYLkPGP9IpQJBsAbvaUR56vjzTTGorXBdEzyIsw
EYWc39Puwk80/OiCJ/IKlZ0gwjw/MC1HJiH15Y9OttABro1C9CqRQqEI9OgSpXdr
O8ZqYJppgvvyK2GODw3MvwytFJkYVeql5SPJLBvCfK9LV1jjlLI+gFP8wTIsjXTx
7p+G9h1uR6IiiAOUqgZZgqjYcw06+GjF49OlT3AZCsvFLDffzhWT/ooR8LxfDZYm
TFJ9cP/gpe0FgsVWByTzyrqg9vlQRjiXrq4UceK3DHuu0tcizZnX2oWNVRTKhTeM
W8+mXQdF4bMjpm9jPIQTlHimvcpziOoKwBPRt0NroOTrJgkmnDYMSxTmM5vR+0sH
+gRXOpymcskF5/w5qs8PqkCIuVO/Ckw+JwpLRiDUwygmGusNRo2H1PmxhJ9vDbm/
jffYE7ZHD7mB905WqRhXb1e5kC7C+1ZpGTdCVSKx0NhWdlsXlRGxCReo9jg4rJgM
XYhOPj/sjxnhBLHXAeKoMTNGaqrPS3kncdS2GqGTUdYcklzv35VV85XH19tDc/3v
1XorDDDeDwaeMyBY2MJck9AewZCWjZDfHfV6ojGXqvBGQbw7P8hH4DtmjsN4GfDq
aIvTXD8Fi0qewo+frPPRMnBiYcb3w3D8fCHPRn5auqI4SU2khdFEPdouVLmSsvFk
SwZW+eEZCG7YrVY826/ljO0o8sboKPhlI1M8s9ypzcNfJQp8otNVVTgHPkUG4vrR
HAdHhPUI3SkDeOH58+Y20x8CqInEAz+4Jtl8vQko6EL/tductHQ1l3VwaUMIEqXc
p0ZhbS0h+Pgi6M4d5dRSlaQ376uglCQ9LbVacL8b5zc+s+Y34Lrco4a9VrbktmUG
ROPgN9oj4ArV5kQzo8pSUFMgAAbyvj4EHJwKsoY9+olCMQYjfeFHgKxfPeB/xl7W
gnq2S8mS9YhwWpeBs8A26bWfAX+lOl7C6kdRfU2xVH8uVT38cy0KOV1ejXHjlhQD
q9IzGPrdlAKDYRrTjISiqM1lly/JpTwR6dgw7qxtJGiIg1ZfAeFJ9q6q/zLbZ1ia
hdWegzaEiiNLccta4TDZnJ7Ep6yFCOLFhRgHEEzBNW3ICM317ev9Qj7qZKXWdZLg
P7VsMBmPatATlwtfrke0NuTSAMDwbyKL6QSyOMfcLsv+yBcPjF2JUrmRDg1IK9U9
h+g+nkZeV3gk196f1wIuDFJDwui/D6CXptI8TSn7+4zIEU5DKe0tezsKwNIUy1uz
1Z122Bw5LcxGU3OaiMN9ptyJc0zv55DxcwvE8ugAG6jF3TXXU9kTmD+3iKUp972F
uSxkHvMENdn+56ykjLdZsQPeJYAfw0V8k0T9Azeva4b6N1F/o/lxz7Urm865X7tf
8O8DM+znfCA6ffb5qW+A2Ga32QUW+bOsbwU/4RXuHCzOxnZdV/+zz9uCKZmPYEuC
m11C7wEWrEgHLluU+kBts37IslrXrizP2eeolUENawSuCkTSgVUEtVB+27q4APAb
W6q0kGgPmZyS/1RH5y2Ea2KEbDRNzkipelEIw1Xy9MZG1PF0+oS7jCLFLiGwOI9B
06NXeog3uDeEVGHOzT31EPrcgKFok2VM1ABKTKk/BFt+0ROREQK3jPKZa0ggTce8
S7N8K9ljqTQI18inSSU1+xJNZ9Idy7JVr0QPDlaQoL+7wXvalQUnrD6pMUEu07zQ
uydi8LU2hghzEvVm7hBu7Uf9+1OIyZ5GVVB45ItlqdgLQzgnQkxJsVKtBNdtglLM
eBzZMYjVAK7PV8ot43mEF0iH6occJLPAiZyVETXUm7/z1YVU2kA1yB0bWjredtD1
1zWflRm+rdeRs7H+s9pjP59oppwmGzW5XXaw4iIn1nL44F7JN1i2G15QWz+Dy0Ke
SRWlByxvO7Wa35W+GJqBTFSmkr69K3jdH+sMCd6HE1KIJmU0rLZSdDTdHJbntYHh
m035aUC5VOo0/ueeZfrFOlcnMth0pwcC3cGZNcrQpYTNk1b1d0pw20pp6lYFgsEv
yolpgfEQFLc9OnyFQAmv90mfvwEBPA60GF5HdfMZ5yTY6D/nxJGfbQZM1OfcwOSK
3azPjc/gf8FpVIjzO4qhyxvXwWBUejJ/Nul2v5U3XEq3jALQzV0PhmqoCc7n1y8f
rrFW6F5s+nDp9LSh+1UGl3plKBPQA8l4DYjyDvxTsqX2NMQ3GJ8XDEFJnTJkV/AF
fDyH9lCg6kSLzrMNq45cI8pjBv3GOz30xcfMiJKQrH/xLKvn2Sat39oTJ85u3G6l
ND5rutjPHwr6SbVzF0gSac6GQkCxefsYzIgzlQhLzanFU+q0ac/NY74NZ1SCIxK/
GPVKPZWtPI6uQr+Y94l/V0qayWp4wlWdBXCmfEnzY5KgipxfFLU8zQjg9W7Eiuxd
LQvpuOStPRbw6flgyXdRVWr4rxOmel6OCpOO2jWDHRregjobHcRTygmZqELVJy22
/3ujHyK7kszSTlG6d+vIn69UcsdnPSzbopSES1kyLlPhzdwMvzGZFLMtX46LMT+U
Vo4eXJbz20KULFRYZ6vJMLt860H2zpaUhZ3DKVT+hdag27R3uQ+CBVTBsRICpVz8
EIC+5k7aSqP7jYDG3/fLjcq2OGqXM9ZFN/nuKiudq7wSXWyLNkB+VuR0WkdiV/5D
G7ayxalKrqwUm7L/OIV14k0gxVWmx6X/B4KkVqgkEaZavLkEx9XjtkrCzqVZ6Zag
+63R5v/fmIAg6p1UnZY30gLR7xFwr6so/lsG/chPKqbVBDIhb18Pyt1QJ3CJwvgS
BHzbjbwFsa+H5FdmFZ0mhmYriyniakdBaCuK0K6pz+M0txMKdpZWfiSpAFYbikz1
Ouo5dW7j1rsrhET7m8kzWTN8zUTfqGb9WMufPpvCMNpcIpZa3PVWgZAn1vyWqHB2
oHz+ZYUGDjWaCMvAeuEyVnys4bfasQ1yvrNE7k79uI+qqvpopVzxfX861mbMN6Nr
wvGzfs3CWnhJSDUZz0DUsv63YXnXIXyQpSt+CvKV4v0DqYTB+YO9efYAb7kAT2xL
A2aWhySKDhuzrWAbKY/PXltSfQizbir9fYmww2EcsogIYcpOBFPUOlBmwBm3lAAB
p+y6HaBE610nzWtaGvE0DfAF0D5j4ctXOmtzSlgNpu6F3anSRQYHGZnuLYWinhes
6j832YrHkC4zRJBr5w9vjY2+eR2TLiIsOUaVek0UDMxZmOhncHH+bVdu/bQvhgVG
+LYpqKwZYCTrg7/0Q8HmnHHPA8XQ5wjN/EcDVN/N7h76ee5HiiSff70zQFdjzwO2
jjAcp+Fp+H4o9c49+4a4YBlDZiNTAqY+JtJguV6MP/A6Nmj0OmESl6jer1kOfqPM
UFvcm+ZfX4gmuJ6yF1J8RdvHEPdC9QoMpWL31NoNgXTc+vSuDjgvmemmHwY/hEQ2
a1orz1EznCtjr+N4kmEXq+Zk/U4Lggi+HZiGkq2zHkWbtCJB/XXEG18o/cy/z+kW
DawDXn6V/b/9kHD3pLSfieQBGJkoUc50XgvOJlVqKsyQka1hUC7jqNP/yWIf39my
EgCu78JqiXEin0DKWRYnTR6abW8XV3tGMdB9RuvUcf+Tl4q41d6zNY83tegGeyj2
mZbtEYQqU3x2UVOdZ8Lklum1YNoCjhji6XEd9T+9N167I7xKWDmxcqjr1YXX6MU5
evgYU5xP7pCPkFYKeu6azfyH6THvnbu9QjlKhA12DQgIJ86Ur20HuGKM4M3C/lyZ
2QRYh1E5cif5bTumV2nXUY7yB5EpFsFlEE6eajEbN0DDqSml0bTnZ+Q9ls0MiI1t
jGDW4WtDb4EJxM3jm6/ebGdmahQ11VScrKDrwkL3aIIU/Cn8FxXWVHX9c+gk0Vdg
suADm6i26AYn+B764zoCj2H+NkTu0c5/VH8TuoxYaNvL1OQNJ4s3OqTaWNhhyB4V
ezoCQvfIyHSpQr9+CPV3egGKnhYLq/ZSE+KMw+ooWnyEL8AR5Hna459o73wJo+Nd
RNzn2eNSmf1OlAtW2kZ8S3PevrJfoBK+5zgrfevPN3qM/HelVmjrst6EncWmXacE
AKyHYJiWeDTqG0zB0EtAoUtMkGcDgyWbHDtNo+yHZvAEWxhq0BE83M+7nzc1iVGT
9VC14oX0YE7kcNqo2uwLHkhK1LbIxNf2BfBUEjEQd67aareZbWAGzQPzZb/Vu5Vc
7M17U956BgyPQtfV6TIL8Yt9KRY07ncFznJ+hqZ2ugCuJ5vnUH28/JpMMB+YsHNq
osMES7GuqDQMls0P0r3/xWu5TIPTxnbXjGvylrMtavzZQE/pyYyXmW3hH3QB5vqm
Zrqn3PehdLTv0UXx4Ysg2gI9xWgd5bDNnkXdwEr5Ekkb9cclcPFqLQ8h6XpaMm14
enGk3/dvmL2OcUchaI58ihxS6sX1/6l44n4tILlevOvuU4QadsQ5RkE+AlmuWyDs
QEfDLEj/TJCPG57l+eOyKZSMq1EO5l0XtGY5Dp7hF0nfol4xA3aCaEEVXIMHvSfE
xA+mC6wsyKBoGzCAnqg0Vb8PStb7b9R6S0mmxS/dHfgvfGOfnOXyj/0RB9IlDBzt
6NF2tCH4AlD1Eh0EHYqarO8d1ZIVebuYkaSX47ueiDHorVoPSwMpOvE2Tg91ZrhN
/YF2YaYJKy+0nnJWGripWxRLRhnboBjpI1SPQon/qpD3ug47Tz953iKj4IiocGyG
gaIAWkpJr5ALUswobZNiC9lxgnjAVqo595bDPk+gUpeODvgl5v7D0R3Rj/Nbh8G9
jHOIK+4QMxhmr/BS2cV0dZTv+G/FaLG/V1pCCL43yDGdxopfrFZdlHbEYn3ueoX5
uOKOiRhyJARzyuBDAnm+Kp657Pn2q4JnAAQmNMd1LA5hNsiKgoeX8EVSovoOHla4
Yda8MTYiC4n6pnV2BlNYly+F1IhDMxMbNcsDM7NmCjx2oBGj+DvnDXLB0iKB5HVG
9UQRaSv/hMunXPcjj+ZaGw9yAm+XWy9/MVe8GbYbOp+8bgW2zBKuyyViiPtyhkVf
usoG7S6OO7TotcI0/BD3zSNFP5aL6X/LCEiKDipr/Q/bcXf9xrXcblwQtVgRvGmj
KNOxBt//Gs15uS24AS7vkVBlTv00fuQBmHXXHSFFOR6Uo+a3QRkBlmWHTYu2RkRr
m2JniCjqWXQz0b9NUsvjlYfGaWaouhXSGVy7bD5M5IvBzTM30XOZo5TEQMIUzDfL
jwntMKZMUSyXUjbfGiCsMrdT/RqzSoJvB0d7uP8L45KAQsE4ZP7fNUcg/7SijUyx
+H7/WNZokUhHEu/XxkNvKIAco9L6MnwJ2ZS8qEZHFZxRqLa4t64ntz6XNfYG2LrH
9hdY3Ai3BzQfxo15yhtscz/X0kGtrot8BD9nfh69Yb2mCf0SVs4w74bo+ovQ77d/
eE5QwdCcitQEpG9B9t3ygjESJmdP308cgHCRrha6gsEBFmbUNglCiKSJ2SKZmOur
o4YjqE9TZCYDdwnrhAX6UStLPLMG2dTwkzJaoObIMJmCRVDFAnBaTSB+KiJk+WdN
p4Mtnf0DkCpNbUeJz82m7OQEZXzAY1Rr5vaSdzYolrgz5A/g5g5VlzwGiLaK+eet
H5xmL2nnCYhDIAYch85OPdxhIJ23MQo1iLqNCHanpNdE24iJ6Uc4kEoJORL2vcM1
nvRh5kPl3yzjGF1yjEgrkLIu3f81JKZzDI4zVDlCbAbHUU6uQbWjhQRlkGoj+viv
HNc2kakDw/GVsxf9/a7CGM8T7ccSZ2d3/HFjiAEmZrpS3jV1+kXVEyoedn3t4HwN
JWzZZ1SPX1XUWIxABeXA+RH/iIFWk6gPCyvxVQaLNzb6EskBXLIOprqyWJ46iF5d
3VdFohDNcJn8a4SKeFrp3/Wr5Y4cg2LmOi8WT8S2mwPBSIuQDdWzgRwlbqgnyX/P
aqcqxvYS0VRsDWAAMtNLfTr07WvVt9S8ceoojziiWbXVEuIFVmM3+Ll6ModfLQYj
0itncAlPawE45T1mYsV3sSFeVz7abpVb8L4H0tUJYfF7xZqUkiKhoIhkJ6bCRLTb
RtC9ywFbVk0jeHMfsM4fZmqN9haNg0SUWDUDgGu7+wmkneEKRdiZVjxrBK5Mg30o
0H7ZcurX3rss/sc1sG2UqkWMhUJtcavqjDw8rgN57eXvLvwFt1sDj8fS45SNF63B
bYhBphV6CgCyzjHOdn1Fui5e0UXB0YVLh/gMXW4ekzoI7GzKI9o+000kBy4SU5W6
E6uX6PwT9QkSU5E+C4k+CwXH9js8EMMWvb+I25MKJp/pivDY+IJbN9Ln8Ma0SMsn
sFiKwsw32+/wkTqiMfYmEXoFbgejFNbq1R/tXM965pWLdF4ORSgYEAdFeZr/btlb
j2ObDP8lQQsfGdEAOwawC8zqo63Oic7vdc6ht/ABab/1sZ5BTEn+BMZuMG4/rF0N
THa2C6FXGPWeqpQpNfAe4Dn9oGoAdQyzVwDaXTun1nxlO3Lryt0JS4kPKJcYDk/X
mlr7FUbZ/9yx9RnxCluXS30wrgjTvdeCJX4P/HFBBaXQ5GvwL7sYdlcoW1vIwTGw
kG/N0SLihXcK8ot+WB//J1wUTez3OVklROuEAqBDRT9yO9b6/ma8KogBLVf3dSt5
tqswgIoeBdXUWRxZvfliCjZE1GRKcMiADMHhdS2fEdtDhPHGWs4xmbO5OC4QWOAK
/oH15t9ueS6g0LnmQ4dllB4cAHhi1kVIpX9WOGR+pXFSpzfLcrCFJT/EW4rGVSAC
hrNORutdsXB4+z9nnpvkkt8L9WIQVUwapiuE1CTojhnyJVxbSXCRbUp4/XRi4zFW
bK5gQHHtH53AfAzjncbObm0rdDJoQKLp+l2V7w1nMNhUqozhzhkTkWhdziyMbiPF
XJq4CgyxW1X01WuGeIzeQm82Wm+15KnW9xzKQbwgo2PGhxZYSWYBVlWur8qe7Gp7
2zTLUW15tLMZ4ncSnsQB8UkpqZncoRxbzImGdpMQihqR17dArc+Sq0+r7ugE6I6B
+ZhtEhpCJuikwaCZs9nyrp5nUDX/DgYn6crb4udQ0jyR3wSdkV2qJ7DJZuEee94B
TvCvf9/mACQ1ggqg15xqaqGp/SsJAnZhu4eNLVuB9jlcJQU9djp1SAWvV38b83DX
vonLgk7lTEfMTzFLHypUUt4WsR2uvNkaJBlAjgnFlQ1SegBsNmHdZH5L2x09y+Dd
ocBTBiAHB0u3z8TyfV05WdaG50gncmn+fABYLT8Vv9nbGcijQ+8/VG+R5bQOf1Rb
qPvv10x/x3Y0AR+NoGozvdzVHFOEbrYFrkO0Uja5tGnj+Sz5UhQLaLiVOAcROGJq
qH8f0Pkagual7pOc5UCstmQjb4DFmKbfpAaglZJO3dD7XFxcNMAriFGx2GawKKEt
zVYubCMOxiyy6OgY1hBvUpb9LvePiA92p7eQbMxvzuQvkvVzBoN88lw7hwhHqpQ8
S6mO2TYoKOdM5rOVsnupjhpfeJkqTSWw41SHNvHMLWXSl/Cdyy15Cbj1w6YXclBZ
Rv0ZOu7/0MsHMefussBEe+EpSyReL4gz1RYNCFNd+5vJHq+YjH66/V+nb8QCCNZO
qw1lCnkFBiGtHgT6B/7yGDFqXlPfWDFbFOqLN5pSHjHuQAjuWbcx+kksqF7dsP73
d/ct+vKcW3WKXkb/q1lEATKDk46Z4qEobTA5JfnZ5qp6rephiRfohzSn2ONVS0vW
U1HOzeM9/Sn9tUqrnyNhF8jVwJUA+/Ygz/ZnT7gg9xu0b8VJ0iLAURVTStbKsRLY
JxakzMztfncgwyD3ths/7ZedrmJ8yHkZQJcVBJSTX6N+8WaxwuchQMblykPIQdjy
3GPzqVVNK5jzkU+5LCCHeaAemXY05M/TC8xQnGaRy5d1SIfmlQP0rUkK4cjgd6k7
PejcidkY2Og7X+TxXu1Tjv998cAspY/qZH0NCyAENMndimeojzxYk13ZS2EFkvfB
nWQZQrVoZoc/GLnk2ov55ChxUeKD7/nIECEVSV8iDI5Mcee7QQ7rrkxY6emMNhsD
RQDslbTA6lvTL+Kx+wj8tpFbtQmvO9DrT81jTRHb/oZmuWVMRTwhCAcyDOHq/87z
7o+29H7CJQEgAN5bUYNkuczL0nrLQ43aQ7kBl89XobcnhEXBUvzx6GNiHDwTRb/j
H3++V4qHbpE9KOl/FR2wrkbvk3H0YmysBGyuXwHLUgg0rXdl3LbZPUR6y1hXNKT5
0lmV/7kFjpDic5DTGidrwQTQMhhqKaEBKoOXml0Up5v523myt/fBji4VwIzXM3MS
kAO58R8Hwy6g9qtottGD7Sg3ATte5bJ42bwKSCweowSWt+RnMEaikeeQ3pFu4lcT
hzQRxGkWsDOIjQP9xO3UxNxHvNjL0jyJhrgYovj1FLqQZHVA5Pfv4sqQO31yW3Ab
MtYppPJSdA53X1ziLuFPhJyzw9BShrAFQ5EGcfJCaSUZvrvTGdLamospqK7ODNjZ
auDCbfS55d4uVNjrNrcSgvEaAVb0R1wpUrfVxgGJ3JGC3TFNjXsR5yWz8kPmJZFJ
Lr0Ka/M3GcqoAY6OjtjMm5osZeEZulzFzy2DFkTEnwg28WJxERw6WiGL5R/KPk9U
QA6K2duJpufekLNS+2y5cvkcc/99R1PqCZnorrxK1RMv+l9W2U+zJEn/tIbAdEH0
7ystWMHUgFidvxYE3FnLAbtSCRXgGsi/sPsCT9BZf1OS+Z2qFCgMBmWGpzsCdBA+
AUqNFdKPi9ngWlBXfraZ0hVZwTUvQkdGIZnBHC/NmyKvULrXoKjR53JnD8IHudwU
huiDNzjml7o/uKm9AVJGCQsrLSbdPgVoS1oykwtmeRwi1Al5magaQZ9uW640ukSN
6Evcdr//tim9/iFtDw9eAkrOCFA1Pj/WyLFrmXJuxqVqz0f2DuPvOjHr7p75pQRI
DEDl4JgUOL9rKLMJvorUFqyj1WyU4d5KrAJyQnxxqMqWFb9adKEJlOLyzbHSvgCL
K41b0H1cjabxXLPxtzr3I7EDpw1iVgFu98Hqkh2t46bzTIRtCYIva7tCNrw2zPhE
8nuOmm9VgnlpoW3F0gKQAH6Po+vyOUvtZ0oxfrnkLHtmbx0N7C6Cl5UB+nefOIkg
bG/CdicjY3xEIrF9E1RIGsFaaeUE1kTqSOXKrXXqqA15cNB/s5L6V/diiF3yA99L
OBAtABaDlr6z2nm+yexnK0FUCoZbvx7p5IcY0hPj66l6PIIPnps8gl9SYMksGbp5
qTqpqvWsfZxP9bmAnt3Ze57BCKAYsSJIMuq9Ahejoy1NmtIn6hTfUnAnU69zSZy6
X0dE6REMr04Qs6BSYixHUcrbxS35w8MmFUY+bVM/1QL7IEjSug6F9tRigsp0d0ls
mIaIl4Q2Ef3QgihsPGy/dK6rCdKKpr4N7HUxPhNASxN6XlGq7yEQSRDqS/Oi1Oul
29CGkpD9LlAJwc85z7N+SiArjKW+spp9ZjH+2crIHnm5aN6zIgaxbRmSd9npmgz9
Nlmr4zS+GGXBw4U+Od6ig69Uz029KmwZMWIQVS5z5AhJ8hO5/oSXVaW4ZP/GM2S/
YRK6/s9+IO0RbOXwtO4WwdGeWpLOcqm34MEUx76TowKzoWHa/MdxamNB/6hQH/1+
oi1gAYs3MbN0tqk9kXgCycIIPAPYs7p67k3NLHJUX+23okVq912DEKHpAm1A9T7j
FU7GGw+bt8bVs07AEr0W3lIsPZBPcpTRUH5pFkIUKeqabViL2GBcgoiQlMqNI/9J
Ydj+G0vZX8T4TEy4sgxbbMuIFATaZxcgCxrac6diX844sSbPq0k5NnCeLxIklWtO
eTivnfyh3q+HmKSecWcPS5aVxClYbU17t8aMiRS2fwTM6b9CP8bqL+NGvnyFqFJg
za4NDyeoDPLvxvEUypo/4qJVxBaIhld1IO8uuBZyc2Jo/A+IsHA41cPJCjSWmWeu
exAJPLYZ/CgEWMMI54X/Y82mmmj1k5LdZh0HrTM9anjEkz5bUgi9WAkqeMcgYYAm
bSRfGivbt8ifartMU5zlwkr95OtuHRjpzRood8KW7IpZzyZaTu8dWC8FVF49LNIM
DwUxYNeW4q4FlY7rdr0kPwW7Kyp2XSZdi40D8gbGe8KJKHIEK5yN7ndP0o7JWCU3
4UcPg3sbrSa+h/bnw+eGV8sqeFbfQeodktRJja9AcuGirfR55tWicDOCXopfrnGi
ZibbB2ZFm44YSGs6c1QQl34UvYgk5EHYlUP16XEARoBAJ0tpWrRWuH0uNoUlM0JO
uMVefNCGbG2yGEu8RqsbZe5fMzYH232zewCUJBuRJ9eGZ1LmiIDhXRbvg1gLtOl8
2IMbhd0p4qde6myK8Y/D4smJ6Rb4qhGUxLnJcWiCsx/06RZbLlckVlbukb0DJdUx
1QNeYWyzqQQtwYfBfEzbOWSCLZ4rsBWMJ9wPD6i5kg3UzBGRtgz8e1x3a9b1x35O
nOFQlNB47OHDy5V2ZYaYj8pFhCdq2ZIMohdiGKvRfIXvFP5BfP6+LZwjLMzYrl2N
e+QkdOICU2OodGb+pFSww8tGZvCWMJ/+PBffZcXmnrOcIsvJUIIIgJ20eE4OaATo
BLfEUDClA4QEO3AtA3hJ89lu3s+iUwzg4RDbSbC8WVRc1L/lzfjy0W//wa5TfF4m
jFlrc7O2f7QP4l27oqZIfW9mYb37mrBs0PES/ZYON396s5E6jEPD/LtF94unwn2m
4wJ5r1RnuBDQUs1MWrE11W7fdE5STw69izjSV9mvJfdMDNOv3VaJjx8PFPpG5rY7
7tXvGWNAqpHXzbBLatmTCJDQWeGuVe+7p+KIvpoNj5TWwtTqSiHSRydP+9aq1IuC
cFXGA9lkkYUaEcGAg+lpgyrAmrQ+EYwOVKie83VJHzPPhtFwFhSyX7iCoEl7FIXW
Auwgo9ogRleSdxUhtpRzrTYfNpP3yXn0oFAmWNUAFJSusIr+gxRx0L+964Hme6/b
/ceXJ4Mddo1obU1wM2S/Jld2v+/QNhT3YbO6SjmoXdnb88wrNDBQ4DRvCEsUabS1
8PpIyCyJ0xS8Otec3HaaTyFGosJxcid0uRK5qZnusnhmbIhRoGYuZSQ68OcbKiKK
oWT3PW92v1AVTVR5uuOFW2VKcNNsa8CcbExo5Qkz4785FIJcusvcjGXx/RzwOLVH
b131Kc/lm1GB3gEa43sTcXBSV8OlFzOJd5uNM3HlZ1M9oEfZzJItkpiEKaS7dRKV
U68j3kUnNx301jB5mte0DsLOsiArX6f1mvmJ8us2noHIugXJphory2rS7y2BJdN4
Tzgtr9ysQJEIPk3/YwZGAIq0YKW1Qfll4UxDNXMsT5b2w7ZzoBG/mvnKquTzW1A3
Q9v2I/iJu4IRBfaR4Hrufc8w8nxQEV1ItcVpM9IDWC7gQ2pt64TZ+7tbOBB6pKFl
VMQayEKzaqVRVtzVXyQCdhBPeKnBkHf+CKYeNA9QdYaWIAxoTs/Mk+0zHPUUNxgW
09JVXWqwdJ2HNBG6SFDdul+Y4+TKZv634yZ8jbjS1QBsnvpEqoPDBTs3pFChTo7d
EciBBMrf7fdkyoBnJ3OzJWbeTTYbkJg/Bow06kO1d2HIInePBLR64DONThoibEWn
FI8+byN16mcPEV4U5Y702GtPje4akzlHa8RfIS1bCruTzoIq3CYAOyQg4r33jUPq
FJYlOJUu01z7BUCBErVX3KFqL2qx8pVNHNXmwyspYc3RWUqGXZthucta8xvXQ5lA
aCsrgN+rLjyZV2dBx8sl2qIeYxkgUXGDm4OUl3MvRVqYGRp7YB2dk9WaJG2ox2FQ
rZwk+u57OX1U/UgrERbfOh1RNVTTx5T0m0wypkdzOUF8oqdkZjSe4Gc7v/Ync3/b
trXCcBMBCLcC76+FkM9BqZF7bdYJVgfos0LH0JAp0CRLapUl2P7QaeM1BNT6VDtn
2iw2/o7KnxF3aE84MUsXXP700yWIYw2Mb5s8kJythF2hBNsTnM1ePrVrHriomz3z
lqqTxzw7ccUwKEvPuE9FAY/YJDDmMk+s/KNctT5u/IRwOdPTIbITMeGpnYmUpnye
tUCgp7rZuf9n4iKTMaBmHXIPiRl1FLnw1/y2b1eApTk5L4YmYD11yFfnZw9w9t7V
WG4TyFDNOkxwD+k420PO+4HpHKVq6m9aKYqbS9riZpz3RZ+cB6OyUPmLpHDZXcY0
miDBuePaCziuXw0pVoc0GClOc6Ps87X03NnteEKCZo3ub3wnXSTUC3canReHnIAh
VjswXvz87euYX+2/fsjj0kdQ+lIDgBoifhf/T9fEmpMelHdT7uBBb8+nckCtiFgz
gLfNcPlfJE1Mk9lGfMwNk7xjEMHK0+mcWB+GShBqJSW6qqt4JISu9OBJKwDeYbJV
JVh9ozltz7DjdqSoxTzWCH0ArAJWZ+6FhEalgpGGkpHjpkJdZwGFTDmcBCK3G9N7
rJXrC1PZdBXJnFrn1tbHnKUiu1+jzb0dtXtICpbpFF0YxZnlniqWisbfKGsX5s4N
snUhZtd7Hfpc6KfJjimC0JQ1Uk/gAtSSnB5AmHxYk+1etRIaTdzgqPfvvG95/iSV
vjNjAX3QbL1C6pAHPr9H/VM5QKsm2lvnhogHk1N01IDqSkUVBOYUnLXVXHzhvq48
QY8LmUXDnxjN/8O56918S7tfC81uCU5ZRZJIDEL7Aacj4K6mz8qdhFdEbJCNAb1U
ax4cqs6mT17w8YNcGobbmPi6qfOAFTErdCcvtcFEZP2RA48tB1MEbtc51w48If8H
4p0wRhygwvCAlubzSsG2nUHy4mhY39RtZ4kf/vmUCbQQHU5q5nJxB8Dc5vxNyXgo
HddUvu0GD/HDvsd+UIVpI3dtq9puDPKIlfmPqiJ+MKIRolmkeVk4qlh2FPmSDK2W
HJO06UqYWolKjA/BagMD/00H0EYg+iYdvwykQLwv+D3D2/BYkXVQZ48kh1Djp9sC
1xoZGG5IYQuzt8XQtkb8TJ8uTEevuzSF+/nm4+hekP6kcVRWjSHKfRu12mhtr41R
dp1rIAdPuuyf/WXctFIXziBjVJ7VIqvetrtIUX/+B7ITg2a0LrmWNXMJBtzGSRe8
fKZxwUK890U2bUBma7fbvQFnG05rReCY9qTgc53nBxePEgGh9qnA9+1SblwCP6QT
rKEGJgrxn7tI2B0SIc+d41MGXCVZNyGYpMhTgxpvuEXsByikXr4I3AUD0qnlDLp+
muSS8V42oy2Y6dW1nySF2D3pZUx8ylB2UzPqErQwGXuTCpjPyEFCzauEOen1Qc1+
NDJ15ADm3duNU43zmY6im7XWI3P/RYXYjgZLbzy2Q2fjyomY4iyVOffe7J5s2X9G
RLS38Y1QznjncidPRFqfjqaKhTg1RXr3G4JD5sfImHnNE+Jx1LX2HYCnLJshswx8
98tDlT/LXwwLCsnO/sURZd1geJtc9W41biEQ0jYW/UN00xwU9t6HNLQN5wCE9D9d
NOBQEfB93R7lnQ1FVLaVctr65J13tY1I0xrNzYR7O2G+IhyKscOz36MmjvP/p/Rw
r5PvDfGmPKXVy3LaqNGMcRGmwQDxt1vFGYxEmlBXbHlj1Hvu1uLjrhssoQUIL+57
ggu730V6+Xk6rhdSjeDsi1jh7eXsggAbr06g/5AI99+gRsPkemCBQdIftMWV/Hu6
7Y6HPWNrOnEibBFjVbrI7C6ZQWT2K0LcVIUVT2SU4NGZ19QVljuS7XUB526zES+J
+Sr3QZ4yX8bYUuCvvZFZPSaWL/Pl6k/stayZ6r4Fw8290SWC/an9rf0dY7885rl0
OINabmUmlqLf/2iwQdko/IbmWOTDWmbiK6GEGjpolpC6Wakomg3DWY/VHi8tbUQz
clnp0U19QyUIPrBXl1KeYqzB4xAW+LuqUxqBTye4nFPHT0nkKuLf7wGorn/034Or
m5flwa+mzzbXZCe1EU2hsNk3hvKNkRxg6xEbSkzICOuDkOtGrwE5rHEqFNUzx9m+
Z/4XgiR0/feTMS+G63hZNY2F9SpAfIMaVG0Kp7r5Tdtt1kPCnOPAF89fDVvb6P0J
MK6mwX3E4U3K2/hlSn84a5YKKPK5p4up0F7NLtQxVPrHgZIoxFblVr0oxFQxik0Q
/OBEgUp2Ga/YML31duSzvoKKN3P0XDf65IuA2SdJoAoJoxTmONtbfOtCtA5aGQ5v
E0ZehTgVZKyEyC1IxCD0IwrA7IkWOWF2lBbqfg9vKDiPcWBHaLjBJYvaryFKyUbx
UGeLePFioh/uuBen0V6psxSj0KpXj+Dhi1ZKjiJXGvodgXUjFxoeuuXFGtWYvh34
YIvguQTUptLC9iH9MB2ASKvKNpddqq3Cue+gK+tkjS4Zb6Aoib49xJdRY+RlCrbX
diaOHQW0yewhI066M6lz0HnGN699aJsz2psLZIzQdfQSPZ4zrqraJpupDFmEA/38
ocMzg6NmEmZZ0ovlZoqjdtaePcObhXvZknpHcuq1DhtSpDe/O8xjGulQOS0v7q2L
yzygCyMLjH6U7ChAOmXsaUthm/h+XfHw04mIB+Oj+/rfDaix498BnDAJQYXXvaT5
ULzkDKeHtJANxU2++wx3S1lala+mCpC4XWTDa+tdYnLlfkh1gU43jD5lrRIAq6D0
92XeB8vCy/+ZiSYJe6n0zZkn9chBYL03UvPgqu2rVPCRcgt3Z4gxmWXEGXFXNbIs
ox30zdUh8cNvj02Ljch6K5I2vVEWZPW/34itqEfnHs3saT54d5TzaF3Xn1GiOOwU
objANM199tfiHCJmMF33w1YCyv/CKa2LngFrVcrahs1NkwcjeEVMqdmGVl3K9hZ1
tcqw2r5RKSnJNWNz7qfNZZa8tw3tXiKR8e9eJrzmmR80NZZZvJIlBpcBRSx11SMr
iqz3jYPSSN0r2TgETs7xB5cTp0HbC/p3iJBLl84DuXxdPqdIfN+sTRMc11yayPAh
uY+btzBnryKtW+F/MXPm0uLlvmM6W8yZqe9339u2VIfVF4RJr4MD0MD6FhDqFDks
r4JuGdYZEsAoZ+Gw39Uv1Z9L3cvtT16SwIboldD9hu41cTlMUJhp9Sb8pSBYopsS
AP16R8mw7wFnyugJcGRyjZF1OVpEMfPAXap72HXKGeLFWbz3yKybjusbrHnRhsgY
gJWY7NJ4BDy88SaOC4yMJVwGYOGgOsYZDOvRTu42Cb/WpTy7BD84iyYmNTgfcnD0
sExxw9YdQ33jl0XOOY8jGsMYB3//w1tBdoNvp6lVKXUTmkMNww32r3m0KdAxW0ei
7Gwu1f660z3aTqBbT8mYMG8VAYdlX9qAw3VBn/csmN9vwWnWl+OZcV0AV6G/w/YN
CRZjkQF70gJ7BDdkI4ebwpU0YBuc17aOEAFWG4Qs04B6dNcL3YblFIX9u/tsn/cX
LERe39vg4EHBS/zhn0stBWVihv6dK5fvLfZf7dAKOn9HAoCGYqxT95nREJvDn7Ge
wCPVMf5K1DOynSDlJGyyuirftDRu80r3JpYms0PLsKe/7ZcPgT2/9y+INtpEZphT
IVcU11PU2QGXx9FjOLrQ3CDJ/qIwm7wGbwVrdA7DzetE1pfNbfLSfGY2MIUYtttm
zSvaapm5ksAQuTj/TEy7KMHOQdt1NbC60iF55VRjCF5lu3O3/rA5ymsKJ5+b+ikA
r0WieJ+5it7jpgpFcHirl/ZaDBZPPazTaTWiZmXanCvOi29Gt/FtsPiVs2bkuKxR
agiyKKDQwGNBehfCSLDO6d2ywJhgaHzNIRsyZvGhEKXmoGKgSaX34Fz+3kLvSRDv
hGm8rIJYsHmwKknJEgCa2uwcSKXgQ+qZW4hJ0MdQOlOg5nJdIRreTWtlE51B6OZs
Sw61C9K99HVHEgXf+PFl37UdslRH+XuVx2pFFz80MIj2YtckscFuux4JBxN1xZjM
JCjB/2A2ysY11ci98miRrYG2sP9hE/rdg5CPO6U+w3FeOAq9wsINHmSLecqq9gc+
FsD/Adjp12ioAXfw2uRNzhybJtMsJY8wuWvVbxG7463x6zRHaWHNwWRF1Lr90uHu
PKrZDWDyJDTr2XEBTz7G+ZRIKSUcc6vLl08TX9JoccabHP3Yw0cpeX8dIJlKq/Ox
LanAnxQIhNE5OLtKIWsqFbwwj/CrMcn0IOeKGKTn7YyBPl/++ogQVKWhWI3qGf6k
655fLVUN0KYsEXAUIDtrb7u+sqK3JNM6PgJIPvfIQc87Zgkco9QbNqNe5fZLpnoQ
QJD+60kjAQpE+flg+tVgjkFVqYwW+HTUE9zqxNh+e66dfbdT/j23ohEqKyLVnNwH
aP/QQg/9rAgpzTLoYChslq9EPhzd3U4zF2iJ02AcxtF0GJYblwICggCKJ5v1NUJD
tkwn+Cb8x6aOANd7n3l0ab7oU4ZOamztkVV+XbVKEBXqfH2FFUMCw9yUqPNjEBI0
DPqeXT6M7U77F9rb8XmKNttMlyGpXZOoEG8QQxDazenG4bjBBzsih2n5LnVFCS00
5Fz8fa7xEDW8H2pBdNurryEJahwSUQaJwdiwXqFtug51FzHpQnwDUFehfcO6uARo
PbjA/Qo6cC7ndiCuLLiP3gmuOAtDdOK0uOSy8sQlIggurTydgjfbxcGp6/9nRLA4
R0/F7kF8CxSOh11gi0EXqzqWXROLd/oM5w0qfHUE6rTbuaYhlpNJftHgz7dzFyZ7
YjvaBXWVCbrcVb8QjzrI6/OAMPTJ1s7kQt3Zvynqq5gdY5a2rzH7N/T+gJ23SHmc
Qkn2CFVHC1RZKdryU8phyGUseyCE33xObqSVkf7UGRoMCiT//QrXvMAmQ+R1b6o8
RXtc3IPIkDfzQ5FykMWoqcByyijUG+v4YyMQ3YirZsmKom2447FQblxIpnzQc1C2
gdb2BW3A3kQ+DN8VjOo4TtV/RH7Snwzrbfe5Pht8qxJbL5FDSxbwynh4xbAiJwst
P8VBlFDx2PV2hrEnVVHcv10kXi81KdcJnlj0C04kBZndYoEQYT0iyCrVhoRFkS3M
1D4HEOfd9YtBh1WT3qjBrEMmxEiLt3fcNTRFchQ+qF22JBx1+Z39Y3tWfRVXWgph
OKsUub+nISepe1y81eh7OqWVplatPSW5beISshnllDwOaYE2C4VF4yNSvraGAGQd
7Zl/NRwKiScfAaeHu7zR8M2TFsm+n79CAiFl+iOrfkhWovuBtXvj9IzLxpnAQbiO
x9/eEGmQQtFZsYKczzRHlKyRaJmYQ0CauuLEYbmj6YjSkmbJYhFuVa8TAEle8zA9
pXokPGwb7fl7ipKLZ2qrGeGIJnMHQg9vPhI4OJN3GRSLDOidXULumHoQ5aLEbzoJ
9hKWa4S6TQKChW2VtKndZqZNFNvSgd1bws0XKzONE7DFuIDv9BtsIkTalmSZw0qv
WPwTKEu7lt9VWmuQ72SkebLKZRfJSGeAg5XadS9MGaOBePuldipVKwV7t2udOK9G
eN8bW31UcFMGx3jwQeAaUoUkwKIxxSIpiVua9Shn0IhCQsijPbLUmw1B9mpwHi+B
isoY2ch3o3UbXgFfMCRhze5RtrlB5lKQXJ+aNMiD0VSAyFj1LtNMV0j/psxVagrh
/9sqDWgw/njGk/t23axPEHKe8pl4pUKK1zqKk1B9zGqFmF5ToCcxDaVDv3kMrCEC
4bILt5+1FAVrDlJz9NwYehKqSgDXLXXQibZEbmpTfp4sJREuAgS9WOcH/y0BC81V
IdupRlx4ENXiFry82DaL3JmmVO4qTtDtfLlfCgaoCM4q1qcUNTgkdNy/g5FH5+ER
NBm31Ux/se1QTIMEvYPVQkq4Sv124dCEq/TPwaNeWGOBTYusTZX0uP74ikizrRQm
3pe7wRof1PArqY+QvVzArtwxQivEdYxq+55qV3zQtallyRKjWKQIv5InSaSjb0nA
BSZWrN4T52ioCOtnjp5wMBEguH09aQAHvJV3uEZfLd5E8geOV0lszIHaCP+VcD/m
ZYwk/LL/LxTB8AzSknPlr6/RZ/yBttgKDWlFjLIyh1+Wlj0aIJ+tBs8m7wDsGA7F
DO7tWeUrvDfruWROxyRj9qe3NsYYWpApkX3yFn7+TOodkRFOmxocGcrDNu4Tb6Xw
tpirIR6USC2URAbk70kiXxKp70D455emvVxoRZ6EiKCigC+HMiakhZjzE4Gg+fUM
ZHDyww8pDr1ydYglKmFQyOpXIobCNjYXA6bWFOhIcZ4paR3zRp2oYAqjm3Xg7GOk
IYGJZ1IDpEfg96hGe75QaQyQ4IGKF3F3v1PqiUgQsEPVWJszei/XC2x4EGM3I1Q6
IVwuV7WWD86fO48D0jd+CwKGOusNv9nbpZPn1PsnGewSp6azzp2PcdYcIBP1MX3+
rUFSDS9oTHmxfFtv0zN6DasE/FmIaeV7i2/Ld+o3DYZ0ljHUnEwVcG7C+HBRWjte
72ziHtO/XJxFhyKOpKrMoBm5RPtjZbW40TSrn9P7QkRYhtF96ulVk8bQc+zbPkX7
8e87ikIHv7fDaH18Ib6Y3ystIx9TVK0tAloDMLQzT8xw2hGz0zaX70Bwo0H2Lnrn
ff77abyZBrHm1eeZbcLnaYQuBq2XjHBKyoxKW4j0Ox/9XnpToVZMtrAP0eun5Yyx
W0t7v2hNMej+ueSYdI5MnKWAbf768t83F/UxiWkJwgH4SIHxJhMjpSdgbUCKox/1
K+I/+rGK168XxxUL+u+Vu21o0M5DX0YXy1AEBPA7zScHySsECAkCCZVQTpb4TIFz
Q8nsOe08EH8UFh2zhbLQhptUnJjRrpzH0m6ZxAM9SZFYs+wZVtNH8j+To79GYPIU
KYaUm3PVSzbRnAkgpnqq+O9iGnBR1LxGDIFqOViFQQRPb7sg8KwZ6sP+5126eACN
p1vkmorTMo6K7hVCQmenT6MOmZEhRdVX1YyITWxqDu8pQ/pdSqwp8oYzG1wz/kzq
w1rxdTyHEjwFTA9lrBDuk10mvbCpfa42p4BElYvL2PdubrSot9ziJ02zfih+rNH7
XhXdYtIweJQWa1ln7PyfIIuF4tbLgH6o1weHMZBlMRQCmKp+thLHCUh+x7xlkD/V
IcjJ+BQB2HQHjoImeodlca/4DdXzUyP8EZ9Lm2WDlXj1uPYyKvSMz3llv/DTQj2P
609DnqGVEYmEQ6HhdhsBiX/+fm2IPhv+qmfIFRR0uEYFZ2YJEBJ6Mz5OiPxQ6QbM
xZY4XjukKlanE45k0O6qYPnP+s/VF6kTRcMtJAhA7BJWgNXQgTz3GgOzfUXqexpf
qhD4NYEWtCXQ3nsRfnrZTyKnJyZk4BOgp5RJp8D+m1/McmqofEHa1ikDbkHDhh+A
eL7OdYS1X/kKbwhcCoqYSh24Mw9I04DhNP2sUt+nYZe3QbD2QucfwRCoLLWZ3zL0
Wv6D0MUd5GowjajtDkF8FS289mK2HNng8ajjr7rft7HuntgHergjh8NL6LxKyrzq
4saXJGHggFa4hby4tdKpKTgYy3JJhMcRMlBBdSO3JxCX0cprits8AJ/24Erk07ps
EXq67GDFQmqzCOrxi3t6PsO8Dc/flGDb/XglsiH17fwqpmR6gw+Sg+BcQUy/odht
Vkn5Bj6rnDU/nXA5bhhuBircsH9Dk6/RW0ENIMHUinB8hwO8lHy8itjYfn32HqIg
5ThmvKhb6jI3mNpa0aXpjnzllqmZ1pvfmk3BbJJYAvJF+nVWKf/lUo4W+plJGKbv
xyHTz2P5OoQBzqk58tTpiShhRJFvJGgSGdQHphoPQn3Y11TaUzAopfWCuoZ++n4n
pWcBxyO3Fe78FsYPidIpgPzCjnpR6rZUrUebn9QBU1NgkuFDnm6NyXzz9UUZd1wU
BsGzc0IJFPEgwmNelDAJJX4V/x+ofmaXt0bn5yvOOQHs0CQDRglu11HnY/Xs/iA7
WtHfl9TFL3rsnuO2I87WgO5vA3KlcApzThjvdMLf45EZO3f8/fnfxl3Ziuw3pJJp
fIHCeDHvzDa5UJDv3gCP4x2a33YDPjIU26rswz7EGhGEOP+TMkLXLIS4kB5nfpgQ
g7LULgUKIEfptqihoCT+dCzLbWyGS2exybKiAd9RcqM7t1fDOEdPXf8PD3/xSwEQ
jTmy1yJzqk2/ujS4Vbq0BDFWNyT3kj+SNREecluvSjzpmvDSru/mAPm3+FIuFdQA
oVx76AYr72VT1iRs185oTen7DWPfCTlQzK/ytAfVAv5DRi6phuz6FfCw53MpUypo
6O1bVO5BmGWpYuDhZa7O/TC2xpGSH1IUWe6gid4YUXjsb6weesiUhnCGY8w4AT0b
Qnf5M/VIexbUjnAOnbmm4UPh0YCnUAcbt7ab8X9Bv+x/My9qSqU3/SrcXqtiraaG
2KFEd1NK1+pQl5stoFOPUpWyrZD8kmf8obT+Si1CvpYmtHXdx9ANiXA0aS1rx4G8
+GtEh1y9Qf/V7ZAtqhSWlWiCBqCwE3NNN+LgA75lBzjZziZM1nIs9KfJYrhbcftL
AkY+GZSUDkurmoslQFvUAsamwLKKl6o6wn11+FBGuMgnLAOqi0RBHEhrZQZ3gRBn
ih2wMojtC1Lts3hScG/WOZwsohcE81E5a1eeO4Qdv0GwGN2Ed9ngEPm1BjYvMyu6
+WANBBSlsg9g6D02j3nZeRN5PGiu8Bu8fevZ0VU5hz+nfosGG8psHTYL3s9ZPCzo
6RGZrNDi/SxSN4PdM+MpoyppdVioJy6dDPIX1GiV5Xq8Vc+0MB/OePixhWxyqa46
t5uooDX8nLrqXB2GfDMqIkPRzdREhFQQZbD/UkWTMUF5OoqtCseWU3cnyxWa/+TY
RswubAtHsud/fdn88Df66g3zsW9R5LzbvWSLL2o/wZhvtEga3Do5BxgpgCeatELO
2wADN+FStL+zCuEeavr9sQ7momest4ElVVToU2Ux31hT4fnCWmdX1qmp4T8NrSXM
PU1RTZ+A4MWsbrtdgJF7kLK4/HUniiYLWJn02qrWL0HbqQTJu2pwegMbrDpy56+T
Ka0wbSPy8VPNHp6LwTxZPBqAvmvO9IsjZYEzDX8soZ64k6QMEeojdPd0hFSmutdO
19kcH3SGB1KVHV+u14YBnqWDUnXJTmXsmzKnbWRWLvooSLb2zX5JasEFFbEIN2tu
1Qu6I7gmlqaqyecBqDwqYZVFlfHB6dYx3YRDH9HUpMggCnriNu3jL+uizmsaMUjT
FvcOF/73lvEfAkZILXbSZNOF9MX3Fj+JFhrMtPQK0klJK9V10VeC2271R+8YrDiS
r1AacFPf7VCSzIhpHkVzKX2bl24R1toW6ywDTUEwSKQFYqFXhUVDFX5fP34P/YYR
RiWcJfBYLlzmLs5Se9mOz+l8ecwEfrqYK4PvyrTTqdQ4z7/0SthapHD3SK2dLck2
CJT9SyfbJWAAYdr0plWswm67rsEAJv9ubEEg7rNhAy8Ky/fv9Oh+sRrYn2nDRufL
7nV1B+J3fY8FaSVUQGfyOPelKJLSwag2vfMPhtxsqXKX6SsI8gfwYiN/rBKg42y1
3E1fdoHVe1++lnGjf8jddyyFYOb5HljGxFrEc99TPiOY0tZ0ZrrQQOv17ojv1ibS
7N8U/be3dFUEXx+cMjUh4EI5BbJpB6g9YXsSKhqYDn+Epx6BzEwTuhy8pigytsUQ
Hb694upYrdT4gvmJAcOB+MHIGaZoeVnjXtv3hilQ70aDczq4nzX+hqAIdAV3ig9E
tbdMUJzPfX/1kj9XY1QACQdMFsNABgu/ofwot5GwE3NbuW2Qm5hNAsPxuTmGkEB0
fdDuWL5u3+hO9yVALFSLmNt+MQ1sP7szgFYONnVPpaXb9b0KzNl1RU1XTJEPQW/x
995CcTHqIAprzsi/lCzRYxE1nliLLf0ninMv4dtnQZJIrulLE4Ori7i77gQlpMcT
54Dj29A5tkF6Db9IXCQ+rL0W+exNo2/4QBJ/SlBBvOGri7h+zBaXy8M8cHgDQ90i
wMKb4bJf2YPdb/+0cwhZQAmd5HMuNDGUZ3z+O1IWwP/m1UDhZjvXso/quIA9nXwf
PBpXKGr2oe6sNeKUCn+BxDmy4b8VuJQfahMlOdcg45BJUC2QoBbNMt/jk3qoy1sY
ElG2rXs9E7G85lFYisUyYZKI+ldEvfvyh7yPtoxrv4UwvaecZulmP4rTjPYcUInm
tAE1df9yQ/GZeCAsl2IMhBkTtSFFmob64Cf21BYOcichExsLk/O6enitoa7xcIXa
TWC2ZhIE7v9BPuzjRUBca39h7WkWtQungDjS126LxpnCBxKWBS/AhWWpXloJlDOp
OW6RNtS+8CeN+1vcXdywHpJMvj2o5EhiYqmSuJ6LG3ZGXrRN2QH7oLBr4bVCMMzb
TmldG8JSkLyhpkiYR2fpwpnuh6DNyUoXohq1/qhvDMizaJ+2pEhIkq+mwyQK4644
zq10Oq5o3G4f6n50OPA1ihSj3gNkogtnbhcUOp0u+upRpcRjmLvYatXjX0PmQubt
d5hmmsoWn6tX+80jVhGXSsqQpbEsEPgRm2nP96qQ8V8jkK+PxSg+KV8OiYkQEujS
Jq6OQxlwTMst1cpkxS2NATk7NopbkH1EbR1VfoiT6eIhkPTjpabPfgx5Y2BWsat2
YdqslOZXWjiBgz0Yvid8vWu2ADQOIHnpnRx1nOQ5if8YUAX2vaAX7MKAAwz+owjB
OpAPjiBveqNrV728sPzmVB3dLQ4TriGQIitjoEp83mLmlQy6VgY4XNNsd0KTrkIe
+u3AplN1CtJE0aNBEYRLlM5GdbpJBTgL6JL7/Li8sif80NA1bPb+RNqKsj2bq2k6
aPFEyHNLqY+suxEe7KjI/Hz/hOyfVRwa94F2XMP1K75MNNFpPi9I5KiLhNPmqce2
oaEd0Ciu+Zw7qzggS3HyDEdQVpmXUpEGeCdu7uJwYMxgYkX/RYa+G6GtkoAWvTO4
ZU45UNPC+8j+Oz/gyL3sjHc7BkJpJnolm47iMXdzIoQZRfS4n8RXOd88O9Anu9q0
ZckaMrtxxawRW6MTw59mxVXCeHX1jprCsCUQa52IUl0io4ZWV6pAvngQQfG6y2mh
SruXZQoOGo/lmTIrqiBS9xzYQnn7uVN1MslberUbHNAxLX3dgE0AD/8ENCmq4p4a
bO412hAscpxF50/FIIvB0hZg8WHsBw4OZjcgkr6Opsmglxeq9fiefSf7A0y/lJ8L
qJHLz5MfqoDQR8PSrkhjG425vl+1iawAZep3DPxAi4Nw7y3u8oHg1ve1dVqudPmk
XkvGPSaAQGSbIC8aracSxUCOEnp+rd0WUwyyf6dXuhimIKwwPSH7IZPqk+Rm5CEy
irQkj+Dn/Bjp4qpp5JRpsaFJv/QJphmn1auqnijPLqWYPp/J0krkJGTlElmkgT8W
EPBdBL0MdPlQrqsXz8ASfG+m3ICIRJa73Zz5DLL3KXFccJUChV5UYVuo6h+ofjuR
+pDANAqL8mCvhX/EQ4wpLPGXHp6zO41AIiVrGU/VFARyZvL74DbZnnY6ONqxmKjd
pmdMupEUQ/Q9DioQpbjp29MFfgdcVBaXB4C+pCPfBNuiboKwFh5zhEPUfqLcC5GK
bOct8o1de5WI+WxjwRFy3kCI845pW2HNgwS0LkFxoHrqATt51j7WCmafRKHVKEt0
wwGrVsLG7PD4bHPdl8eacpdB3hi5rnwu4EzXxPZRE/LJfYLG4dCUeFvQBxvLWxSF
JvFPr23treXmi+cGUsxNGnHTuXIslY5frmnzDfHbuqpy//ORyJKoU6cTcLAFxUHH
9XzxFGQe6n82Trd1IktcJC0wsZxbVv5/PaNedTUHQ2Z6cSoq58Laq5oOL8xX2obX
1M4LEZJzfpE7Htn9BANHvlNv5SV2Hb2VfuwV2lj8jqDIsr5AgLeYGgUC9RXymB57
SmZzfZgA+d2MdkE4CsQa15RhCkqc3jS4/b3lWKJ+Efc8i66U+tUvXi/lBGp+VorM
fIYg9sJiOJld0NUkznJKHHlSjgOUrUyHRUaPP2MifwMWbgCFjs017SZvU0Rkr91o
MB09ZXjPTYgWPTiHBkH1Y9VMjjMv+g/IyQDTU8h/V9yzzmhcVJXe/RHbc9+4HOg2
bNL3fgj74Ps6NbaApkgF8e72p5yaPA+KHuYZiu2mTFI305/WEanPLhcgir/eNUUD
u9X3ARK299KliKhBXwPnJ6wMeThfQbbwUXHQf+4+dHdzuNPiQcEs5PFatPlFLBMV
VMAwBiW7GlNZodjkK4iE8Oa06MaIMxe+FlzaETGNlQV8+6ykmxCocwCrlaGTDeVf
OL6Iy5RlULo2HS3rpdYizltfuOvDdmJ5CNxrI+yZ41fjAkXZZdUZBbiyRRjQEiZ3
vuXjmhozgNP93ROjSHLvHs3vr6dxJqd35rNtuSBgGVjvc2tW1ib3YhibHQTFphgz
Q/qv6qoTPdeH7OnICx0c55lTodYP6ubryuBy7o1yhV7HLxFJbRMJsiIvw00rW/AX
OkxqwGFzBjBkm+ONtYkPhEaLZqgSF4uDr0pRoOMtZP1qsfugrBSxwnggQC+hPwCL
uJHnyl1EXUQbDEg+oA/IiAo9nHRZ7GInm51CC5xsz+I0GKG78fPQK5dXQCU/BMD7
HOqwEmOJfYUWQyVrvx8mrkNrnEn16cxf+V2KGW0lQyQC3ncmmCkHIew3NPH1UVQ6
bX9hnOh3xk3uWoGQHDhLt+Lgk9Qb4OQMSiKZ2GH070owGXmrEWFbFafy+dVFf0K/
uLjDAcg2dlbYENex6GQKgfdEXF9PelJHOQfM81Y4KUp+uhrKT2FraaacC2Rf9g9B
ctHDbndqXDKZH+EYuMvu95jNH3nK27QM83TgRoH/PhXYaUl4ndT6dNGwdc649sXo
rz+FeHg7o4ZHZ+topVKiceyToy/XRNL88etzSFpwNYpw81pP4bBUrAVv9Mn4QrMt
qyvNjk7dCou+5ZHJ/Xc2Rhd9ivWzFhFOMitxgEHOjMkT9a5SqLx6BbectlKuQCn+
6ouorYkYvgQTMwlWXgMORpXaJDI7z6e0uq5zADTEa2xo6aHDK9oaNqRZ3mbaB4HP
u8VoEsaYLsO8SCrVoTevD0Ugikudpf0fLFR7QQcYp35z2gWs1lIQ7kYkWoTD8VKJ
cNJdGVxeEWMwMd8b2ki95/pshJLSb3Lr+X/NkqZ5u18kHJTPqqpUqNwShzRN6Svu
GP4T4BYfqn25XUhLoMgo5wBoEZpseK/ZXHkFaokzIfrQJ1QvAJbkOTVK76rVgxmI
/r0ORnaPLxELtIEZWTFx46/maZwEXYrVHEO8vodg6gfuBqATkB+uOXh5BVpfr63B
IVFLtHRwjwFUaCkFkl791ol6XQ8c+W4szygWq3qPH4i0V5c3gWQl36uHDgf6FLza
r8vEbaHp4hTTAF0dSa1wsrDICpntkXP2HWty0LKp+0QjKLJhbbOvbGUH/c+49ayx
WUP3U3AzptXvuZxIGcvPJ/RhF5zc5atlj9mSHsVBkAwEiv9AFYZ5bDJvnXXt6V9M
dR8RKBuctp4tkEqwThH5Hy3q9BRdnocNHlCIB6qTUg8X3LDBVPvsIM8KV8xuhiKg
2zatOrmG/pKWT8ZMZoZSOL1cGcPNJ1VU9SBQitc1ukBzhK7mikjRlplt3U2SLMMA
BPvIPwGrGhmw4wXDV6LM6gCFJ62zb7akjMhBgf+fgZKvzp2bDZ1PuBxJQngkG3/y
2XGEfN1eozKyqmb+26Ha7uGWXfh9eMgIMpGktZn3A2WN63VGR7DX0xJwfsbjqtLq
IH7Eo/p6VWllCloFhreXndJgDBciTQgve+6w2DpkbWiIG0BZnhWF36jM4c81DCrY
G93BS1nPhU+QHZqWLROGaVWif4wfGHfyt/AuHlYhonAfWNxuXAOK54k760nwF425
wxw7RmZ0KoiHlNEpRQ/0An44/JEeby37jJ216LmOvkgdx5OZUYE0K8dbShsdOc30
ZUcW+J2nz9ZGX5/ZpRahvzSf/EzF2Gp5W/UxbckEBUBCeseeG9AGEy0vsdrJweWd
wCnl39mKV9y40OfpU5ecoYV8vfnV1viF+TEeCws8xcNCIlMp+0SnhNNMw39LvrcJ
2X/tDI2zLLDW6QX5qFnKY3KD1LQHwnt5KKeW7Q0ANV/c/uUg0n1NRF2CdGZ6nzAp
itAPwML6wHP4EFb6bhONJNaTQSvU5TMsGG0g8MjoxC/Y+YvAuOsbOeLssaHzyBuS
I/1pVlp/glYut9zliwA/fde7OvV8GA4Em+M4pY0N36CWzXo9KTKwHIqXu6QDMtZc
wjjd12niKoXCFR0KnvHuuJfIHxES1s9600vVUjCmEXcmyB23zGXDGTGfj09k1iww
Elh/woREFVNdjHd4aBVpiqcw6Pt8+gJP4+wgDV8tXdEKPVyCIU6OaI/rpfOkEeE4
svNnDD52dRGWiTlzjepmbhSXr1VtR3Qk+27fpJUS90KdMdc3Dw7p60h/HUNZtNzy
vODHJBhGdo7K3Uiy8WSag+gdbDyrwuRwOkRwhAnUd4qAEro2BXVeBX7iNmoCEHC1
dP+FVJsHMSC8Qru9BtmFYJMVaJgFmmByIQXvTR7FFibrNcW+dHWSAfGppAwXQmcM
/aUPJi6WnCrlY6giaToO6R4LxzEHQ/LvQ5OrJDg/2c0+t6q+G0r6iB8ekMd+0GIH
eSNSFONDxY76+iCJi8pHTfT4ZlnAMjYnl+ZgZO3/8cFwqSB4Hnr/kI42/JLDFrD7
whk+xSy0bagaFEaItf0Qq+3K3c+Ed4YUHUJ5O4G/qQL1W1ano7MfbFt/89vNNurx
urxk+ko3eDiCsjXS6jI3LKG+DNt/52drNccyoyvZwk1caKRJq5E2xgiZZHqyBR1h
rhJAdFhiaGPrPAzCLMf9Qlog3MKNDMFduKrUD21TgO6vCBELNGd+7O/sfnu6nS0y
yxk+yZfNylA9vVvzIA57geL5O5lcCleE++LLVWt1KsZYP/lQnrWCTS4OuabuUqPw
sk0Wxsx76ZCuSSJCwv2nsXZXjVFTr1Kap12JPdkX2lpR7BNnArlCZJbl6qHKbqLH
KaNltn1nYSbKA3LQmu0I6dR12mswKGmOU9RXT49bHX5SpngfSWa1fa5MkWpWY/Nc
1Fqfx/tjX8CAU2d7R3KKHePW2YuYLrnG8KFqH4gg/vGdMuJAgq/KvBfqqieLarkt
yrHHHVqVjc0g7DxK8x5iNdPd+nafop2UODFFuzjRvW8DAubhfSSJqkUf5qN6Vgc8
hWxD/WlpM6jxJFOwEK0QK1wFe0Jk7NFUFHDDQmzHRzr3ls7VRQXCj1hIh77c1gW8
qJG94/WIiaBrVByzz78qOxaCr4UXD+OSxOjyo5OO9V6IhRRfo5niXc71jNTAAdPH
9JecPDy9ryOjIddrT1stiZLY0Ccq1UdaPkDQ1tOnf0PYfxXbE395gCteYqH4pyMm
4Gq5BNrloXMi75xnp7BpiHOSQ2HCFpvqaqcf0x3hiMSf+AgzECYurbYDcilUne8v
sdAMawrZuduHHQQJSKLMaIcxGV8dgcffPtGCSuKYTnhbiYd0QHo8qH6P0lpk+KVH
R8gdhv7uosS/VG6XZR7tVnzKY4vg5ucyx9zomiPhbkaLkV/fU6HhtZFQGYWQuw8w
7Ddw6KlcuRZJoWjLpJtFlkDxSwUEYLheJ6GiEEpYVlLkBRSWxJ5fd8oHtobu7WVG
ccxk0b/AvW3QxgUrkEVMA5TX3VJORLsWsSBQKIqHYTYdBf5Lv7W9SZyk9gTDH4/S
oey4pI2i2EYu5rzJAtbfVtn71/DOaV0w97Ox2rzgVGjUc3NY1Q6kFfjouHnnOGGX
aAeYi2pl6te86gRFTYhZk93rJK1Fa1lZK4MKNoLfb45F5Z2xwK+97Z7v3G/1WWMH
jg28cqWDumThH66BGyxx+M/EaHBIgfie2EAUp0E4GUTY7x+AJKqwjtCWHFMMR7P/
1jsG+CGNR9In9x1C9sw22v3C1Z7ebXksa1+iZH45tfz/7Qt0c5ozZ2Pd6ExCqqVY
AEmJwNW7liCI6ogKnGhQUy1h6cjf3eQRZED4kNaYN09QtAec1w07tt2HEPH1p7gY
HvbGf9z2TUoB+Nsf0A/zz3ADQaEhE7qWMcjiONAoC9HoaWGnmJohrc0cEYW2jdHr
Qf/lzJePabNm/fitieyYkHwnBfU0qi2GBI0eB4k/iPKctgrMGZ9NAMEELRjo0p5I
POIS01zpdcsns5L3HitTN+/dKh64EY4T9MsNLVCr6AwU7Kopl5Fo9vThMZ8zaucc
2nH2CKATWwYmD4QT0XWKgHMZJCgqsYRUrcgDWgNh9XZwdMXgter+d6cUWTWLGzXV
nm5N0O4ASkkIaKKAZZ0eV+bkPg2M165LJRtz03nywPe+08vvyg6b8z0qX9VHA5H2
2rinjufVFElnzbOf2Cg32J/PlPDufUBrweP4Pt+7+k5KoZfsasyB2oVTSMTm5/0v
e2juhVcLI3hyPswuojQNexcmVrV+C+PAAYTzNGdAUP/eJ1jVRoRrRuzkks1QD7uO
BNEvj4CGfYkyiVJEkfrPApw5WP9tITi1BW6VWtUqu9Hc2PcjuZ+HjLx34iS+9zLk
XhMsXBmRGOk06oBEINrl6SMcWmpCeYnijqGfJ7pOnWTM8kv0ge224xlAHVk6uY0f
9CKNYc9GVd5AxoGvxc5Ak3fRjBSnNVRFvTWnYz49/WqHpxByl7X75G1VoTTU8Aao
tvMawKpvsk4STHMiPTEQYZlcUhTOumGrfUEA4TchJriskD0vDt1rz8kqVoigMxK9
Dd8SL4QCnLAYqcVdCKqXJleHLuCdWpS8broQ9L/Uegl8b9ZOo54SnuT97ZhZnoqC
+4hPm1KcI0OOWKO4qfUkCLEVy9IJ4aMSGX0FNqCbcQh3XwVoibzDkKCvvlgynn/x
iyeu3Pj0O8R10U9lcViUy+z2rLkXaF00ITGQsYZBhfJq0Un4Dbc6peFbFiUowkdS
R9mCzT2SbLTNYjj9CzWqA59RtQVK90P5Z/2NbfvQEEFIyibVY1DTBPsRPtg/p0ke
LkY3zUCUhdZiExChMTR4oC2nXvqUd91NTfbfx5w8ST41k9UWKPyEHnN0t+BuiytK
sxkOTsFjXnRASBADUM7CwDnnesI1knSKjWiylQJSAx39MJZ7eNojr3b23oJPUCig
RNK0dpbQ3DhhyT1S1gUBCyIcbgshMrR/Vk0U9JDqYSHAHvwShxgdD3JfBe7KYsSD
UslzordGCJIMjnFMZ0O5HmTEEGgxJ9OwTR7Nkznf961S47fUNKt0OJheXDDdkS5o
8yI92ITdDZ0T+jLtD/VDC9ZdR4kjXJ/o5R+pv+JlEv5Wv0yuedJqPHv1XxeYDy5C
RsQ1KEvw3OuiqmFVcJDUA4Y+7rbPSVqCivi8Htes0MnUDZu7fGYvoJHw8ud2nUSA
y5y28XVxXhPfjduVtJd83pjkTCZQ7GbYUBwk744D41n1e0ihjwehEUUdAqfw9Vyv
R0HY8L8J9x/73vX8pFFmHxPtx3NIoX689uljOKpCKUQj9QsM2Dqdto2FzgN2qgX/
a4efasULQL5E4QJNuwd2OwT0f3GCQ8NCsQoJXtJrZwDXGu+DFQ4RsT3/i1oqpDjf
Cxre4qrPj3ssI97HVT/t4jpPBdDE47EpiCAX2vIkA8swWqA5YxsaDZeKsDeZ2W0o
oNfq6awuvh6fF/GqxNKZ4pFMtCJTT3DUvXDbZi3ic1U3+squXirlRPTRc2NmtjS1
97l+Q4ZVqmNE1gJl80v2t7e7Ym0j0Amfb0CchAYSJbJDHzoRm097nIhxc6+LvzUM
nMKctBHwZ7LmqsL0ooJCsRS9zUXE3ryjq97whAmQTRTHJlEFCE7bjKFNplJ8lAM2
Lk8EaYLWtRaRzu+jZft0TMP0aH9i9PuZvGn0vb1wj/E8OF9o0qI+4uzDPjj8afqC
pVQO6DkOOcc9lfv8DtXi0qV4tyiNv20srskuCBkNeaDZxZzYlBxk/NXvWWpj0YdZ
b2R+bUMZOzaMXh3BWAJWIK0BW15cAwhaOV9ScaRR8O4e2iw6agZMG58DliaU6Wsn
i0xvaRopTGAdM5JFF8dJcu6GLINBOnaA9gVt/ThPq4vGexXUm78ZQF8URvrmqtkN
r2kTZ1deMNZbnzf4YFjzJc3VEB5k3ptGf1/vXXsAKn9evA5Y+kWg/KkseRmOStNC
CY+t5n45CUQJm5Q4ggZ62s45blIIE+PyWujwZAwZ5eMIkTJ4n+SuZq1S7kzWjik5
BiPLThTcT9Po6vC/Ek+S8nu5j5h8JU4YVj5yhBVWxiq4XDLt2z5d5PKXVYzdq//U
lmKoVW48WI0mQyKhlxTWrc9dD0+YJiaj+Ys0r3r9r2pSMCa1JfptupHWI9rtvF9c
YWpZjrvAr9PbJubY81aw4jcCqARpNiqh46hYIH7WGcpptyVQleMiyL5b8dRuAYF1
c45+153jaN4tJkylyqVXw8K5UdxQCfoxdDR5IxW5LXoYBKHxxtAcJ3lN2YBLEcEa
LkX0+urF43Rx76XsGkG1Ddbupgwrd6n5+Cb8rJTPXRKR8juostIBvwsfEkV3jEKA
Yrc28QZkCGn/tCOuE3aayII7ecO64cAwnj64nmXaAA228M7SVUBh5cnRln9E5ONF
FGVM9YBrQNs/fM58c/EzSLqvvcT00JmNTEu55utZFTzkWkGI26rExkJrONll38+8
ForqZ0jQbTIavZDe2vJ9QPnKCqHvpwDOK5vqs1YbRCSSQm8FtZqY+Qjt7m4hHDE1
qdj6ynVun4Qcqk/GpAdM8UW+FHxE/L74l98fCoo7wZ/7JAfE7Nef9d7AxG0NaNbU
kwUwygcbwnJLsaCnarvp2atasqQsVz0JwUUvPqHWLB7b0r7giR19PwomShT6i1ky
izw6iNO58Rv4xbW7FZw+oMAtZL9UO9Bjkc5ycJwUK3eb7dqfxBQwIlas0IGJ1np6
erP7ROWwER6nyoY1lkzUoUWjLQZdK1NWUX9PdUqLrOkk61Cc4XwYHExZaYNER+Hp
doFuw1q8fWh3Sm9/LjdvoosTHkc6bmD8EKqXQgfa14w7gRpsZ41kji/InFWd2gj5
DA+S/WytHmpurD3BCft1vc/dQ0Xvkx8tG2tl8dwWSk9kSbS9qwmlVNNscvLVsNVP
1a06R9IsuobT/BKLDGpqTz91XFHXRsg3btIojadThj3qV5cKwolQNwlUVQMaqhXE
3mzT1yqE1HVUuFbuAmeMPCk/go+zryBV1B/+JKCkRq1nsGSNhSMNJAx+AxQC7EID
D6L8Gyubm82XLmN940vbiILgSlVwt59jFOtEqpbaWEgDL4Xl0OIH6qjTQMirsh24
jvoLXVSKSehuCB+6s11wPbYz0v7+Eu1+TcKFn8sj7bCZ/dM10tVHgz799ub8LvrQ
yAZfJzMMuTGAnEWKKpgHdTwizoj7IMbKuLQJuimKbLalvgp33j6LlRQf0xB3EEGz
0JWESFuME7v0kKcOPqDk6patLpCQKMJdXN2m0DbLrm5dkKbAwA18upNjE1bXyHTn
LQbn8zoqb0zArLsyAZiTs4jqdkE+BUwgyQ/d1YqpUgYm/gOrAbIJY4QFofNJCL0N
tfHSp33R2vaWdVUT1/BQvK7babyJPLyF3KZHpCMvmHogc6gEcq7+W9eARk/a4N0C
fS6ObOz0nSBSwAbpy2hmRvq9fRwRCpDcNSD9FK24UEldSz/9AlGJKvgGq1FXzXr4
OpwYUC7V7C9cq5Ie2eFqjmFu0QVWybAQMM0a/G8ClY/t+kHRewA8QIXvO5F6Af7+
QqCDzbhbHUnaGyUTTT+EHYuR6UvVZwigLs69NtlYAr0EUNYi0aFEWlctm21cDX98
zOSZyQ5tkiLmehSNxsNkZ63Slo2W0djr63kPPjhqNJ2aYJCznq0IBBoCTLg7RZdd
QFedWEa4ThJbDqbXgTKtI6EHsZ79If6IUahPfInSeRpdyw2q8SqdkHceoUmekKvN
f5nfmS1UwLGV66Im6RQmklZelc18zthAol2QI3SlSsK79D7TKwtrvLaHudO2ZpHe
SCHsQ1v+AANwvpXv32PBdyrOLfygyChX7cZs+kJMQF/rOaGDzj6K1znUpsFX0Hbc
Xl1gKg+y+v2z2/hh+2Nd81MNgcRe/uHzcE4l1i7Xc7cRLU3c1qKk//NjjEY0HPha
aZvcvKw53jZTLYWkMlDfz0lSfVOawVeMUQt5qxXvWHtxLBOAZDr7yB1ZcC1cOK7H
YOJA8U4vi+s/8Phh9LPj08fGl6ZWObGBhUbwls6d1ied9Nr2nORxQzWy3++XHt5B
MsLEeT6ulucB9bW3XZ+UuTmGaH4HXQEDFeu3PjM4advhF3tH48612glerTDnFdP8
G6rInaHMby+d2OnhxHvZuhVjvK4Ufd+3kJXt7fd6HwWujVVX8AOqaDvpRnBZLzx6
Y4zWV9O76xX1PC8f+VPfNYkzb3BXx9zpmQR99JlJb6zePdHtOvkSIZ4+jDkOXQ3N
eDoESBgy60g1Th4YFGmp6qZyV9sq6Wf2ZXD+jNH/tSUrOe2ElnLvXvZnyoxEbbf2
ampikHN8Fptofi5xZNtrcXrRCPCpUujCkRC1PySLKJMQfDssFc0N9jOnUgarlGun
ZhqA7o4pp9ljmkCBvTB9C/uitLfFKHT7H9q2RlAOw0vyA2ZzK32URsIrJrXso217
5DRpiv3knkj5YHzLjOSWxQaZDypHCcMveB0DLE13RDLKVpHWh1qTGsjXi9xTMBAr
/hCvAOXJ2OUM+ybPUbLLsd+UQLSe0tLnNHPDLr3L0LEjq/RVCRgYSclXw+kEDidu
6qbksF0zbrmz/4oIlWRd+OTYbdU/rxeti+7Lb3EIYAMw9YNKLm9frSYUuJhTVg22
JJbIQh1gdoFBYrX9LPsTtuJ5s3UgxsUbtuzMFmoD1/duwIGgb61WgTQC7nxBoH54
mKCTT+5c9NtdpHifHIJxavRyyid1j9ugAF51h18tEyDehVBFpdTztBMJznju+dgh
1fDuJy1apV3dM23S/z/yPN8jLn9HH+Syz62WC5POwEj8fKtJ97ksIftfzOJIm7xx
MOI40jZ1yq7BkCv7P+yZE1wUAk3W1hl580nDrU/q0bXNj29e5NTjGuawGSyqhcm/
BBoDAlKJ76GcZ5OfNbqox3As/XLnIPZTXy/QwW/xQJ79CjKoVuWdt+jl0UtmqYj5
q/fha/FlXGqSznrNF3lELysrsJFZybvRXn13bzfFuds3E/MtGJLtxpbjbNSm86Ac
SZPh0TkOCqdgScSE2AK3lHMAL+5LohHCiDdFHgJ8J5Z5/ra9MYA4ELRhLRZ3rWMB
+H4mB1T8pnBEo2CezY6KE5Vsky0AmQXZiFc1oE1BwvNCAN93vbApeC12UHMQaE7h
YaeHh55cPONFR6dj4RoM/BxBoehRkFXIH8Hko6Y87ZkYYUvtDTh5JflOgYVMtH+E
3/Oh2x5q2Zj+957U5s9IZxm/QIi2QV1I7lgpWWmdS/44SaFFG2JJXkn71KCU55Xz
QdAQpb/pUrycMULG89rBX0Iq6tYXu1CykffagbQC+wv9pH3u6TEuDrwdbsut+IBI
0YBRmlcAy5YlALU2tU2nYfBI9b6nzf79sZwfqaTJggaVf/qJBr2lIAHn+ed662XM
0I+6iC5TPudLXogYFeu1HjN24bP+zSSSSNxgH0ePtIScOc+Xo7OdYTsS/MyUvAWI
6Jzh+Udoh1upYUZPUzu+rGiRuhJ4sMSJs8itZVxvhhfxDoX7qP+6usc5ondmImsW
4B0wWJJYuHBmZWKXAbM4IIWjgRSoyVMj7EAttWGx35oZoGFUjhfIdSNZ2Bmh6dnN
Ut/S8BX/Gk/iT7/ivQ2qjjRJSPX1eItO7Rcq2UpmA6wG23Fw3ufaoec+rXlFqbtC
7oJxtcREunpLoFIpi9OQNgyOiFuQ8bvbBulhU6ZzU+plcZMx2NmEWsw4gRmSxJQh
RxrAJimRg/4v9KXdRE9re+jX32aJw4p1MoJp8uDGnfLdAPSp7/CeK3a90xb3fq0m
JstNaHxjkSMDaxin7R6tH2a/CCIAOL7bQSKXgtmPM+fj1A4Ectn6dr7s7b1KW1jW
Jj9vilA6TYn/TIvGCb1yxVD/QJH/Q8L5atPOcd2DPTg1XgEp7oH8VEhoqO5u34y6
z6U8bLhxe//Wa5wuyBIKYbOkIUOwY8V/oZJQ5ZuVxIHBPfbUnBcRerUOGOKi7zX7
luBf2OPR4QcFdPGiRdw6xdHM/QmsiP7io4OMPmYWKXCW4JUrCMcW2ArzIIC3dcYB
IsMd+5TuIBGEkq3AKy0kO8pATElOEDF0V3hI41orKoOB0NwEYXB/E+nkYFj7+tju
3Gryw45OE/j7dfbbeg25QInDeaw1WJl9Aijl/6vuSeJHsrLYQTQrQ4nAgaTv6BBb
YXJ93O4dQySbFCj1XehCdd64t8wZhrqM2b1CRy3d8RER0oRmh5Li9OJhN0/hLmgZ
7ti/caZZTtrI/G69K1d8d9tSp9Eh9MWc3Ppuz4Xzj248taM6yx9+fdT1HDHDGc0P
axINqDEbaAnjPrS6CvLXqrKq1vk/Zrgsbm5fDKNJoq98bFOtC0ifS7VGfRC1zOGI
ss3/WB+NN+wVPcHU96if1DM1f+5NMtm5sfg8zL1X2mnZCsckDa0sP3w10ZYyrj7D
el6zJjUwh6Ti0WuaXNB6c+Zlk+FoEAcoMNOzDLOMIay2A4Irkk+yyR4PjW+RQaft
J5C8vRCksnMF2r/WIcvdfkh15jtr5GQkYu8aFa4OuG1qVR5JfJTx2GGuosCTfj1u
NZKAs5dNm0/syP1fslUArBN4jGTekpgx2VyXpAYncAVI2SQoD+5OGAuz1W4tcgqi
8/7lljxizLSuq+jnG3SR7F+zf4VswUj17GpIFYMu3bEioCAJJ8AMwNDNQFJVGiKp
b5XOIdbHP/0nF4F+3sQMmdT0NE4xjsoctk4Ys6ay/IkLftnEZl8kgPfc8f1xWY3q
BvomZyFiJj4jjvhGhh54xDePAN4mj9QNWegr3SDHbD9i+4dJH6hxk7QKfn+Sycjg
XvRNoWMQFpLXIUHKnEsB7CLPtXy2xDR2qhg2fM0NTLEqsaOb5bI6lAeGo5228LtH
XdH17WAI72PGNXbWceVx0klp25/CzB75p5jjvV7Pxr6dIGlP5VxW6fF3ZkJFPKqG
onWE64ajnuiQNg9s9LK7fDdIcKX/Wa8iw5U2iUG+zxa4SbT0RMfMWglF4fzG8ch5
sMxyG/ifjeuFE+UP/n8dq/X7PZSCfNesFUBSwuu8h9sAtptwo9oC7EIcfuxxQ+0d
7MbBSpzASXKMy1TCDnhJGGruJO/QB6DvJstrkQ2JVFl+qMPvq1mN3U+FEZ9uQNR3
0grhPtQjF3wkT2TbqOw30ZF+nT807mpKxiDkucGvhV8R1FlDpfdaJoLHm6a8XH8G
kBKfLFvzx+BaBtd4bCfhyRUPqiCkMZNiLz26Se/0NQYEDDfuO3Ejrbs+nx/ERC2y
ZTQsDS3E0tlzSmAzUC9kZgNcXMxg1uIUmaOmkCdSXdY1e2m12hDvW2V1JkihC63j
HWyZGy2JbNxxR2JF91mpdWyIlX1Nup+8pD45Vy1UgMfRdJmE1MsgT1cKgVbUd0x2
nzDvEwHV3EboDbiH6UVu4GisqmbkOfQ3OqIilV5qMJGEIqSWM/xEkssLU+a6HQln
rjjK7wArjQHRJW3SBqgCRlsIjYH4XbPcBXA6+PZcPvMEaMp1mVWDifCZ96NW3QAg
IzP1l8wVA2EpRii6cttGl8Pf4X+DCKKAwlyiKJdO3k1BQSHB7cN6jrns3Km1tl5D
6E5puS6CPAmHnKua9L9QdPU5BXAyNzval7GaCJ/mD7Q22jlm5yZasceoH3HVhJp3
xMXmyvS1ox83XB3usczHykaX5gIBp0KvuouLN3ry7eaHjx3VZ7oN9EQSsjoYM7EZ
otF9Q0WG2KRqsoCqrrk7Uzuq2vkDxCzuzFDPoG4A1lmmnXGpi0yX780dck/tH7cz
9Iq3q0B9GtMR8oSO44ZiPvcA0HjzcCBfUjIwVilpZWnlgGH/8ETmH0yyI9ekNbjx
gOCpo0lPCivc51u7IHI3ZRUfePfqmUVu008+qsPB4uVh8TPMRntGbaI+hRDSWB6e
V5ERy99WFSfsPXSgEQX3A/2/KnH7I7mInuqEHS0vkJlAPwEEWWYjkkvKddvqAr/h
s7r0HwSH3kNbXGbMgapTO8IbU3lebobivCq24EfXVATdqGwZRq/JUmEE0w9ZX3N/
wP88YuYeheQFGb/QzS0Vlvjc1PSULZ7HKR3eIrSTAlHxOZR4cau4+8HjFJmXVkvc
vXjIohoDDG5yrM74kNiKLcFSDfCfgxNp48J8zqLJqiHr0f/+n6pUBlt5+LgG6zkN
VtzisN0Nsv0sR2ZiDaC8zNgmQfOji4ZyffX3ONvHkNmvsOYUCZ3re6w5b3+RH1Yu
3q5Q6cVwo3OQhOSm9OR6p5crz7Zydn2+N17ItID6Onol1Z4/xu0vypXIxn8cvP1W
x1kYdMJqJlvi8heIzex+E8cUT+UGy7iJ7MfBQfQNVzp9PrwVOVHEGOaM13bYkCuA
dkUtAZp8vfhZ8Z6sloQKjbbr2nHk7y9VAExfAZ/SAGrNCoTvGyw/jyYMQLqQRc/A
meVYeMgtKC1fA7S+GfIZUosNTGAMkGOnUVEe5UHlk8TZ+etSKTG2U4spwaL/ErFr
QGeWfZgvWHXYs9JZEQROFxITrEzV0pZ2I0KXVWMe3wdL1nKdK52KHXDSEwNgd1pG
nnwFIEoME/RDbIK+CC/1CpQ1wBiKKpOyoyeHUdTUh4rOg/8sV3kZ1Yg8ACNiXXVA
XHzKRHsJCE+p3dT8XHZjzNJ8Aco+P67Sc+jjb4WWMFdpI3nBAYO2XGQ2Er57p/Y5
wzz9hq0/VX84dr6PTqWQNnmcf0fkegV/n8fP5D51g+INvoD+42b6VLi/3is0bo7I
4T3VjWF1hsaQTzuobU6EPV4RxrOB0wKTsxDZEtKRfWRqjCeeagdez383UhpFuPm7
dsQxbWL05UfieEIgvwbe+9s0OpGHR2/Q9ADsUdVNKpg32fvygZJjEKAIe9RybvGF
U1EwKkPjpxl4PVGefVuvNnMdM0ruesCZuPRhWdY5ECpIufYI5Ye4Xp1lKad9tKiF
qj4hXPQ7uaaTUnyFjInXI08jRTS9FD9MStiR4fAm+y3pjxpjRA+Rm/JLSx1VE2tx
1TpkbPxb3+8CAaopqOotr+4l5zSvIS6MudYXsVWs6gr+M5DW7e2SWbNRTM0ADMwC
H7zC/EtZFryjt1ZBvRqMNhp5gJmyYmUlW8x+hDdtGcL7jTqQtxhSQ4O8EBkL6aX9
yQY6xQ7ONdLlYXXrYWE768i0PI5DCSHPR/G6bfeTo1CxlQqFa8bP76JE1JZJLueY
JToFkXscF4d1tvudlaPzvJKhWfoVWX8CQUU4OxnZGrORcgskYz+7Me/OQFWF7oNK
5YeNarjTrFlKSO0HfAcycLKv5oiRwgTVCnDYDYmBiQvONQGYJbHC8fXoZvXr5eX5
wVLxaowAdEEMfARYIApxtNdugCTLjlr5KPvl0SMODStsohM73N3fRexGtO813oDD
/XwTHNbJADqVSx7jJ4WKpPl9wGnJBnIeLGyYgQ3cTzSChqTHFRX1TfmgDDEig3z9
FLSblycMbccF8aELvZKAkLrywG/NIVsmivYMMSrUmzmba/iCKmGITjeYQhIY2XP6
sgXRjVR9ml1GRQb1vruJT7miMBRJkaZr43KT36Htp5M+QAsNSUKqZFZ4domgIkmn
jnzznz9ikGMWVboaaXGznHBQsu+mKmYJ4o23rgb8n7+vhz4QKK8WGlGeBb/96IiJ
eHdECnPqESKyK8Nd/8AY32+2+mW7mPiOoPVlGpN8+fvZ/PgfekrpW59AF6G3uqjT
kKOLBg9XfPV5MP7KunBIsoWTEYrksvjEQadHoa4Kqlp9j8o90q8/AdT+5HGcOGQU
Lj5//NEisdQjc2O5QJreXDHycxk7TIivHg+DBlnz+8gx7rJn3JrYNbc0yrSd40qe
Ski+2ZCiUKZN7eUu8OT+PTA4jzwoMZGxB+O8xuMeXHegjvvbGGVfgfqp+953kqys
DxbqzHkHvGL9mdFOaXDsX0B8DQ4a6iXj+qJPWIpmjKsgU+APmwCnrSHgtWMPIa0k
9aWFWa6oKv8lhduhcIXkjfkhRPvTeo0cLECuLPxXhBig1OHzWDj5q2UZjtcFszd2
9KUc7D9LQoCt2ZAVlbOMssqLVBQoXdZxsl0BoiYUL3tAhKn9zZErB+dC61W8B09k
YirXSRgoCbMt3fwb1E55qYlqv1Qm/R4XepDbis5wJZdvNJD0XoxjWJAHGMuuFmiI
drDLMLEs66+xwzA+O6La98dS4XMgTZgAYGMPe/Cq8smC8pH/3K9Bn6KZeF1I/cmF
odB9PLPMSOCxdL0fFjrJKzESrIF11j2UDV6Ls2i5nM2HITnH5TO6ZCG+NCiLIO8Y
+zIxX22Ao/iihOVBAicviG2gd6p9gBuh0d2NlJECUgv8Pi7OppYDoXj6TDIghNE/
eUDI1K4tsW0YxReSzzYRgGlv5XDC4quuapFRQVxLx79CMg+G2Ap7MxNRGhZQ454r
UEaBo8LTRBZ+0pwYz99ZR6zDS7RvkNybi1zEHRRiMIFi2jOZ4ea/TXam9dy9IhEX
9VhKqr1zY51LgFDeM1YXAGlLzx6ao7pux0T7QSzBjIYfSOwFVgxXF1Qq/VeN5n6X
dwOCjoxu7h9TtkDJ43nQXgPSXtXNCUnSNxo0o6uRn6g0YK/ovDpqM9RHJX7vWP7I
uV8LxgzL4O/cCaEKNxF2B2DIct0CSZaHrF3w9/16HgN73rQqvRzB/XzVHRmCgIIh
dsIGdKNBoupmFljo8BD742KWH0pCuz65KW6yOsfcGXAZsyfOSBxUdxA18jrz8/UN
b6W22EbHOwhZ5UYu75bGi3yM8mdXJuhAfnC3fBNZOAcM7UGjwEehtY+31G27bh2V
58PT81lWYZJI2SmYuDmvkx5hki9b/BtHq0FbfSilLC7vOKryQA3rzMYV9nynPNix
xEthFySxkxly9QA3eT/DZI62CWf5N4MnT4lmdgIyCJaQdzPDPkQNZZdQhwYYD6ZX
YzMTeQmZgqr+fTED93ZjNL1tKWEkTifOzOvLX2E19dn4qBW4QURLjE+kJP5oPKFQ
YCdGeSrueZ9F3/7DQfJlVMlvApumvaPACJnWc4s40mflbrR8GKbhx4LYcnX71pkr
GVgXuLugrqC8u7uM32GtGTR9lQbrwGN58NM0wQn7w6AwJwoF35be+ONufSFDTOMm
/WV8o5bt7D5QY1zUnPJY423kteTlY9hqKHb0WpNOLVqLbBwB62panG5tQAVDHuSt
vwN6kkWD+UGbt/ELt/Hli7QN20WFexaha7u+Nv313Daj5R+tNF0SHB2uv5nZhksW
E5QPr/7uE8TX4+nXBWS8QP7Hm/3K7cQ8U6xFADHOHMYv0lvdeE71PRy/fUKo+PCj
x6qPyZZ9icXy6QfBxyxO6jV6Ar+m9F+9z6s3ezA7MBjvYPItcxVsL3KEuhlGonoM
wTWalWvbiqCywTr2c9gn7rZFFn4jAlSd1VTKInqcA+Lup6Xs9IqU+BzzFIU1NAM4
llk0q5cZ3aABsznK2NyQpMhVZAZHqpcXBgc1AqmvTMmR/zee8f6URvneGZle89iW
24RWlaiM/NQaV7Qc4lplILRleHA22tFrE98iGfBUoumZf7AUMgbz540UKMlARTce
Z1sHIUSExfaBhjFNcNg4Mz6EJzbZvuCa+pi9911Bsud9JhTZO6/BtfCY0NNlCDPN
L5XWA24ODRWqgs3NyKJkEqWqSpZn8YJWFhv/CIdw/8qYYQ9XewNACicIWN2RJ5eD
FNl20Lz4IZX04WSGrSvb95QFytRszv5lyuiMlN4raiB5e4RmFRC/888nhfSp3TLV
mVR5K+HkgijihWQ/f346ubZVlofJy1/oRDBLGWCt/ZJEjEK4RxT2JL0GUig5UZgJ
EHhtN1KR0Pv1/NDmxa3EsM7DiVOC+AWxRbUeS9IJEwT9JsLlQP+hyw3EE/EQvkDL
ccWIedDyOao+WQlcONV8/Pu4KxH0XywtL1/XPwMd6m6IfKhAzb/8KaALna3OBJ3Z
UttHcwpaagLQ06f11puJInvd8NfqCELvUNnPZjEjyBMuzZW0njD9/qEqO0d8IDcm
zTMQ9oDs+edlburkQr2dOhL3zteEo+4qL7EZLmDcvoUfke6eYKsib9Zfu9AzVV2f
Ht0O7/D2x0qiDNLbJ21HHuEVnNG7FF/KCSVJ3EZN/NEiBAwhCL5oGblBkAJXqxiJ
fT551k1Z81a8Kllj4EFnCmPb5fs0nd6oS+UvFNOpML9onznAiD5Npsd6eXf7glyO
M60ra4jplHYrfMx68rIZB0BM55ULPQSBxmm8Yg3SCo3sVn8r71ZsZF9h8+NQFdva
u/7yLcDFYvauolhlEfOfgORcNUqt0zs4czbZYbHJdmqtUuG5JO38oOdK0NapbB6G
yMUB8RZ03ORHeK+llbyeVneXoEee6ENu+ImWF20M1w3g/Sjx2GmJw8GzbZGne21c
DFpKhvSIp1DQJllqSWMcx/l91DB3byHzb2unqLuMkFwpmpPuOz+xLC3/DQKqSWis
KeJ8bZHuf/LcPIMQA6jDUkU99rWmZTq3QW3kgfD5Ywb9SyuCRc59HLs+srSdowhN
7t3sFL799aLpu49/wauc6kVMNPS5gNjo42IrUGoFg0UFAjpY/MQpt2/SaB4Sk54f
3F+NfUYFq+QYAo2ODduzmU7T044AUKedJENac0ICOFkHmSxiUcW5Ch2dmrgDoE0f
R3pMh1gV1o9iv+FQzFlznsvMwxLOGUsoYOMAheMybycRt4m1g1wErljO6xMnDxNC
7FMz4EkiKCS2dPCCXZxUmnPldEweBSxkiZjSeKBAIv2dPm+QiPrhxPPy8m5wF/94
0EDNVNDqCcrKDN9GhfLEktQiPOKjn+F9XNF1/HJFSLunxa42aq+43+lp60HqFmsp
Awq5YcAdWl7tTRBEWZXzd+tHicL/kNvcaQ9b8MNB91HDZAEO8ehzHTqqtEOjCsld
osXr2klPo7U7FamXQhCBprbIUL/6elC82LISbtbMuxyRIw+q9/vFfmZYFLt8bNL2
kXzCLehmVWQt+XCJFMVAXe6Xr2PjwDrlkx9aP321yUE0REZjEd3v4PXBvfqPmhxG
P7loksBI2qN0p3q1ZR7lZw44c/JnPoIQPw6P3/YTan6TgF6uPRC/Jx1p7eMIB71G
WkMQ46B2zs/QP3jmTouYOOor57AcLmWHVlP+f5ZTxAfXvFkJ3pNhaSWZfd88Vopw
jl4Lvpr4hLbHf2UJmAdw/IvRlzVGVwssNJXDCGjYe+tfwubXuzyhbN10pglCPevu
IwI1ziITFjoL/yorlUH7E58s1EWfmTkg9oL1u8wxGOwv06frHwa9BheqzJwkOLtW
C4jgXC/oGYPNcxaA6sVJhCtFBO6DUxjB9XJSxJttvzyJElnWRhQpwhzFCqoUGAp7
TqB/X5KrgqhyrNsyut4g7jGyzJJAh8/1qLn311exA6VpEPfBNkSfjM7XL0SyViJX
Zm3dZVxuXXwlnm7CKc5XMiXD20qe+Hl1GCY6ZVRjTEeBG6AxGuFoZhych6jV3WXn
bFU/I90uEmnQlHIZqK3Y4geabYFoJoqjwEMR6esJzFt0bsQeJLLKqg5Zhl7LRApr
5CZ8Yl0l+cazD71stW0D5DinvCFKWixYn/NCu0otSW96t3UEJOaDD0Tb7O9M0PsO
uXhGK7Pf1F++rh++O4fYWlJ1SNYNl77giDuU+uyOcMGGiwd8D60taeE1yCcsp4/S
/BtNZNZgww/B1ugWtjM6KtrP4oJfr8+Vw3PPifnn3tI8cVbRu8wdXL8ELSgXMmHq
ZOWANq1skkP5ClMdXW74D/Xq11R0UoCjLHwSOZdkbZhqVZ8/MOLYzBSCOScAWcv1
Gxwv05yAeXIST5auhnWaki5BkW6rOtlla6JhhbGf81vW203+xnbiQ5BiZ85j812L
V4Qj6ZduStmDDDuDi9Sqvi/H+BvtTKn/pRXuZUZf0rJkHyZGztbD3Y95I0oGh25+
AvMZaRX5OOyDqq9f8Ps7CgrHnIYK9deqLvqTAeaSHMqUwbFT4I6Ot/BTn/CjSqAg
8dlrGe4/llzLUn1LPaNZ1fUWzmZMIK55UoPtYxOC4yL7Y9LIfUgjZtW9PWLIzrac
/EYmY0hM1rLIZqDHdnNUHQ75PPd6yFUBEJNjdlmoDf0is/sFSTBPM+FnkuWL90TK
hLZQnXap0Lv3wvi+LSoUv3zuHkQQIZvfA1aHjtSUn4/OcDWdND7Zz953ZcpVh2ZE
HO0K6/bnwNHGSbNK9U8bp6/YHx7h4cbPQp/5sK50JtE2pAUTNZtRw2Qvklr2CFt3
YP5aXVSDN1mS1nPcyh1KNpyvjNQhf/Dzl2gMZV7Fa6q8w8EzE8m70Tdqki4+6tyU
IzUG/XE4AV6T1M4Y+MMPAw5HPEbbY3yBxv4KWNDZgfOnV0AkSe6IP0FszU1ZicOZ
MsfZtfKLlGy01qXdzXVGeJ4AimlBexYuygsXuURyh7NnnFVEfdMOw3lFpJDRC2Id
k/xnls3/hB4Y98LIOGetAEx55XBi0di4PyOs0Z4W8IkQGVtVm3u3JgwnTqaSyzar
qGfJEc/Q16t0qUBxq+Bp1auGeFZzeAjBDVXXtu4dzG+CzhhrddLl+y4pDlZXV/k1
CraWi2z1Dw2AYK6ZcCn+ICqVo6X38Lhr6DKKp4qiTvccQTvmbaThRhi7r8c/SGI+
qc4nXN3kH6zcMrmji40nHxiys04oPqqaEVgO+zbP31NiB5BfMyEdZBKQ3JLr1/N4
Aw7p5aiHSFJve1eRlCtFJQiTIs9wO2ixx9UdpukSvkzkNDfUftnW5XrvpovUahFf
Y1Jtpu2vw9PfH+mopJJMBVFFhj+dKwcegKR+98KCs8oZ6yJPFhO6v86OnvFxxk2v
Ijnlwkwdcy5epeB6MBQY72cDXTYA+Mh8zLQFlXGcN3E/RKS4InnIKEYco7S0fJGb
RtrbvYD/CY4YgsNNKvQYOk84/biYizfa1jMMVt670PYRjeovJ6kpIwB5yfEZUxF1
LEdj1z9UVXB4Buk267N51GN9/4Vf66t/TCyYojKNb2CBcRUOFVSq5TtpKGTpkGea
qTIihBipq8OQ+5L4u9uzJFWoVagF7RjAuwQm9SSi7LSSsUlDe2TuoiYkyGYqQf4Z
/j0XirrUwVIQNlInUId8Dpi6iqFZTitBA0QN2nBs8gQKu1wPJ0tA9WlR4iSYQOzr
kbgtdKSR5mBRMQYagl70u3hGdl5ZdhxIq6IaNa2h5hPqZE5UtiONvi4/SKmCc9j0
lOJlHFYYeIHscQwDALjK38/8NC9SI9o73JM0TdYXCRUXMHHAFvPV4//9c/B1FfyW
20QC2ImFLEXLtwGLb8XCKlxq0pHatxXUmdX04ke1C8TucZdBv+5ZXCxlujwvXIll
wxXPNIZraHLFAakY/++Ga3KAoEvfM6Vt/wFtEEwfTRQduwP1uz+Fvo0/naZOD4IX
51b+L6C+wBDSuO1XeiFRghFH2AZhl5rbd/PdGm2s0zWLACuXzl4vdiBvYpw6bgoQ
Nnv6xHOz+s8/cTY94l4krrpLzxsRlONvEf4OEUR05TGemVxW6uMWlo063MZ8X7DD
AzD+KHqmLMXNMAZxyMMjiKT9S34AFA+PdStb7TbcQWlaLPqGknAK9YhXceL/iY68
CZjz2E9thHbTs3mkJZ4ZF3IKDumXcaDcw1OHtae19y4pwr4ioYUpbHeQ/LQTDWyt
G3ljS8fy5h0OlRpm3QRbl56H4UUpcNMItkkuzALhVyrM6YSnwhi/vWNuaFsKCHHi
9VjYIfY3p3gaS5MUPlhrOJLQx3BWDyQqmhH7CoPyE2l4G7zX6hudeEaTVBoCDHTG
sJ8j8mLsvhnY/kHu879G/Obo96FeY4Wg48gJMSNNDDQQ4bZ59wSBPgBnjoCdEstH
YisnGkRDuNgCmov/vvobn1iAnHM6RjSzeECGYeJGq/B4599Zw2TkiAGLC619Mo3Z
ITmI3mjjUFsKoPSC0y6I5AamLAXBVBgdTk7iBCByHE3KbhZJXaOFt7XHgvMBzrpr
bfpMKgfDCuTy9O7SFNXKda1f3olxijUof5gyvTs1hY20L/Eyg28KcMSjQjaCTpaN
etG1LU/uaJed2X8LZm6kzE8/b1m40UUnI8BwVgZOTuADdUmzTs11jxFYjd1pdmfS
BgTJCDBkhqtfvq1v3DWbSwtaakZQdNf3t8m7+Vhv+vw1D1j8Sfg23vawuuZE/nsd
DndlwMwcRaPLyp1Gqm4nN+13ltyALX3csPMiLbX4jq7g+tJ0a1qfySYJkhtkDXDJ
uu4qsTBTrQYxicYAWtsDVEqWcRZAmMMOoEQeZFx0cwjmiQE3uV/0uNHRw1/CzD2k
P2s2eD5IgaOdrOhYKmu3dbNX4eslwCpk2y5P3uu7C7C41MneiQFbFjtjZgl75yJV
hqNrlNR8lculx1u+fEcLkzaF23g51sGgYNGe2xuHvwIabss4oGophYMa+bRjejFy
PcR7lXJWn9WR2AylcOp5ZGua2oWC3vyPIEZ7G+hKZ0XsMZi6q0yABwrPOhjArq8i
2FEvLWAE9qxXoK+r2xgsEOphU2/vyGyNzyTQVehVGvZXJQSmsSJ9FspEA33YDNfa
yr8mQWieuykK0GUpB34YGIgKgwLdWnE7AYcGGBNLYpgCrPn9TTEr6XAtMzDEeEu4
DuMgYBsLrnVtNpo2p5QlfQoW6bPGTB9Czs12dxk9dCvlNpg8KeFeYUhl2/+Q68nM
xjXDD4h+tuYfbX5Qcw6RAe7OWHlFRu00TfiLJ3TQP5Cv4/nlerSMLZepNKYtBBo0
8uSlJYbEVUnHWsZ+Y9/UYWjJWQhuYj1kSm2EZ2yCSOaVcoChgVkGMAquj7BL6X6p
C+2c1s8uXXmxlAgl3IQUWj7UHnXmhmyt5pqXqYmCbHhMR/P4PQ08vFv4dYwR4Gah
SdApy4XJ/9vqU5aMm+ldcwEI6IyutKVEUI2v5IzmVWXNMaATiCxw4psPj08LTYPi
rxvpw+fyLbVC73inzwkOs4nBwO+RRL/ySKcbwn+uWHTRjbXM3jQFVxRt46EcVMI1
nVH89F244PFlWIFXDHj/s1WZ4v3MAvQPtiuPSPje7q3IKNxPYO4ek2wAEAbjgnQh
bHphxUBnfEsqlfiz4nxudDI7NimKb0DsVoHWRFJ2pbbKgDk18A36DYMNzMWzLTVc
Hkk8Yx+j2zkBCek1SqXSScrlNUeOEFL/qqWtm3OwQfQu0bdzfEdZDi17//MU2kgg
CBY+hDL5h0yYf2Hd5Pqdxg1Omzs05bO2P3zmdCiur9mJ5S1ZPipozTFa0lP9Pb//
ytY6IfGpl9FUVBHDWQDB8b4YbNXYq8m6rE66NzjlL9eq0vd4QmzwiVUdOL3hXYDv
6AM6QnPwlQQDg32oowY7NKg8GXyHXhcgkeZMLuwEbuvDKfhkqTx4TG37XMZEGDby
8jrPIHNbdDXZ2Wtwsbmd1p6J3Mo9c6raqXWEWjfC/EG+RKLMDzepPysRAdweBS/Y
aJFVGhwZqJs8COqjzYjr+yDHrMWXr14pFyVYMzbIAa9bDGEl3/VYd6mPTqDPGY7+
e5/vFk5oWb/Fgy6C91tnACcr/BnuXqzaIh3mY4LSsAStUvNNkPQIh281Z+Z0vvkB
VChDMA6z8aenWbGD91an85xPEIGj6IFzB/QuqgyL+uUb76uiMh3iXb92GN8Vion6
N02VsrPqedZxsQ3va/ZqHSCFv5Gd5jLNxnS3qvn7A8qo2JCoK8PxJMLjiLilSDSH
4XlON/nAfevVtDRDcMJxNWaEqVhcYRHVD0U/rJbob6uqmN9ElD/6hIwUAB7rs0SD
uH9aXAINcS/P9whOzfcllzyJxMZbP3m9J7P18msRjx1uKWaH4uEC2ShsPdkD9dkz
3jCDsITgLT0BrFqsDVqcyg2DsNSSSxCTUEBqyGvtenGf8SNkz6Qir8Sg/4ual7LM
wK/0HLwjyzo9LoIM5803jJZsyKvsElvNRsxjUAFKAYbHj6a/UAgQ57uPQS+q7z/r
ftHFCeK839+Rfrixf0oYFHY1lGMS52g1pzp5WrAmQiEsMQeoHiza/TWB1xfzOh0e
1rA/3LS0LE1zw8mjD8D4RSg1qv1ibNO5onNP4NDPfuhAV8Ytjih53lwbJE7vGM5V
B1W6ZbNPzWMRLLFoOvVpdpbWSsBMQ6waXt4KS+4we8Yzne//6Yy/kgUpmhqVnUM6
2marYJjffL1layFmdoKGwtyaaxOAXGq7oG5UbpQ2KAm4ktQyNB7jDXDZYivnuoMS
xq8bmeyyf3oRB4Ge6HYTe1CP2k+jyB9woTLSR8RBYjnfY1sanznSddOhav1Uy2f9
KaBKCFD50CqISsYgvw+MuPYfnuLAuqiAfQilY4kkb5m7Qz9/c/DHCsWW8KgkUSZT
7yGdfLH2qj4Bz4iKlC7wosNyohNzOa+e96ffSXGUHV1kLd4rB5//Bs9f5x7oy5l5
0x1+AhY1Ifms2qwQwvcCKdY7vHiEBVpRSD4Uqu9MBK2mi90QlLSNBYDM6ZXtMMz+
PLdLlUb+FZZ1sPq1xpCEOeqVtnSkAuXJVOMc2wduI0/9V1oulx3zTT6NgCdtMC3Q
WIHlKcyypMjIpl5UngRrdEjSdltBrFqD06eSXMDEfokA3LndfQ5w2QRIF4G5zQVk
5CbgPSgdm49tYeyWuS326R6nNKLYEgwIGckDRMJpH0eYwDWg1CcbR2WbEMp+9N3L
n9yec0F6MnQlFkpip5sIdFtrWwhgHOwqq5dv/Ri+7564Dz8VCh0IEofhe6rZjnuA
THjvREjE0TIACv4sNLp3A/VNmmTP9QllwUEca5AXWPJRS5rsZPhx3os4EW3XiMzp
co5XkSVy8Re0w2fviU7aTveNnvnr4P8z9Y6Y8RgaK52LZnbbR2hnYj29JzAuwiC0
ng62DeCCGBbAGbRfCDUmX4XRIIdWjvcKaWG0Kkf5umpQXZiyKTs3l2Ef6oYfsrLa
haUxxrsRoIltTbgxZHnia4bEX3A8AJmsPJGaXsbw8Zeehwv24vxEuratqocg+svC
AEfnbcZDDRkH6nUS5nSLcL7PmxqF1jWALDMppBzJAVGPhQOgG6Yo8/NzSHMyM9P6
tQ0CBVeI0+vhhWotxTMrQ/zBAml3BwPpKpAct2CAd3XHBKdYoy106CJ6pzGN18Lv
1zqorOszs1byX/r34uozR045a+xf51tr5FzLM6TbOJbOhvozcfiN4PRSS/RhL0Yp
PZRhnkAzOe77unfOXX7wDWWgZMeEzOMIqzAfieeo02pOmMWG2xiTGkdn3eoFImEs
xXEYfMDgblY3dSy01C+TMW9FSz1FX7TTTyIwwNvS5vVKwtZGaQtGdJ57NmwmfJio
j8PHaVP39bWNHKO6t9L646Srq/6fXPlISCPqBZwPPRVGSqIgCxilwLuuyZEVZ8ja
OH45WlfKevZpRhk3juaXm3Eg2cJ56cXq4ODxEB7WopxroR2rmWhiPDJE/UGx+/Bh
iod8AJRryU87eW0GNTFzmVFpl6DA7agXIkYQX7EQ6fqfaxjQLg2BSU3ukAX7HMKs
SXpZ12n/ATNoSkqAMFUs+LcWDwHiDS/q/oUrOCNOElRTq2DEeeJ5z/Eq4PxWIwkt
FDA0wqDUyjQ4cXUlzO0DPWb0+DU/TKchAKhB8GcvvaIcewN8vs9P/IOldSliCc1T
POOrz5afHss+B1NLlnxtuTQ69T2rmwsxS+zZLXriGuJgsfRR2vbTu6wL1/z3j0kw
70MVjwzeVHc5unqjZlNlwXCSfr7cvJ7EFh2EbLcmO60aEDFSnf0FtqQ8CBxkyaEf
wv1G0x9zsP6KCmyBYVq2fg9oRiQZcZq9DIYTuVwunDgvmm8cSzv2NeBAY14p2qnV
qEEuUESDUrVbHw3TegtG4wPIu0l9z2BVKziouAFp8XvjvQnzvTjI0UaKKWRb7oVM
SEl8J96M6UUSEWZwoJIaieTb0NnZsOUiY21EsP9vlrwKmPTkfnZGx32gVeoAE8u2
XocttKZ9Vfuu8jCSCaOhh8lA45CdMxymG05H+QAn3ka8r9bwGL1b3TiuiOjhe/qj
D0ChGLzRINFAkb856mTnBuns7JRHtliB71Yeq9Wjvf4g4OCs7a6g88yCKPist2nV
aMBLWeoJt7WvqfESkSwm7980iD3GXqxl/2dQor6cz7CTIax2FeXEhCl/CohhTJUw
Fo8z13vS1MTVlDWqmBEKTNui9K9YBGPMQCMBg4zdVeUD4LcVSuR0ki5+arzRygCJ
0GJ7vno2H8DOc0h5jfpP8QeAeMU4wKvyg4yMXFBBe3r/jWiOkCtmE39JNI2z+lTx
276pHg/VU+/SPzcrgwLfKTjSOLHUSi/IrjVanOM0F+Ic6k1y8f3goL48/Gt3qx2z
DGs5guomqDhAO5j7aMdVkrjgZQsYGiQzRlxmPAvbppNcMzdygPqcxA30tX2HO2tX
DxuJTjZaz+HK58twc+47nLUASziXNnAKoyEOEOYLPAp4KdgycT1c9qTe07m7zD6W
cOPssQp/XZlYtuwquYsreM5OHJaPx5FbdQLnC/D6XVy7iPzc1Y8cfkFm+/5gEbVt
GU+X3loH1D9p4jvXl9dZiGzi26NU6N9AWodwv16ZABAamiw8Y95F5P0yM7tsrFdo
ZkMrx/NR/rpbXY8UDUGPAldUI65XJNtqAqepYl4T7BWc97JeOKE+aKm5Gdcxt8rs
/UMjbs7H8+AiyTAV6kLFrGUqqtAeJApvoY8IWYKAX93+GC8ZMKs0HqXO8DuyoSjB
zdoqaXKcwQ+gLODHP1ipZcCCFvHl/952HvI5NWYob5TiYJiIeS7bi6wse7HoM1kv
tLShTiWItwdXc/gwWEkHava7HRTvDHGKNKq69sp2pLNA/ei9fs1ceVre+XRoMkMv
fath3usMqnuxqv7bUCQEbd3heNMsmROQv1HDCpnqCIROJCnpOq+85oA7OKq+nvZK
0+EtOKEwHoytUpuYkBLbiHHmKivpVqWmkyudC5++6hqeCco9dtpXliIiAPtnRb57
d0p3w3zQAtamt3+0RL/g2cdbMGGc16Fszm+t8eoARwwXGe5AIWKDwecuUUHnbLkC
SV6G5XXgLRtYN6TP9r8CgfuQt3ejIl66za+j5AB7l6pA64WbeqXF1fUtmEWfxu9g
eTUC16zokO8XcSbZomdU9iPFRN1sc8dQntNxvSdlvs8YdYlBOrqzBaR90rJ1x7zL
tveaC5PONYuV8pVTBzNhhBi1wjA7Hnv49hd1CZK1Y04CAXhb9Mxy+j6FUZu0KF/N
hMHB77NS9S1Z6qMIdDSZAaKJ7QrSe4FiNfSyKuZBbAnOgeBkpnXu9UAZmYumkCtZ
UCMj1okFMpg52ma46l4/9HI0rPzWAtuJ4nIut7zNPSrA7mVMXkRQtabXwILrwVWZ
ozjlUI0Mwej4s7oeMZsybO/haeYElB1MpTMiTQyN7bnEtZmgF7dcZ5Xp4927sIVP
8mEOmSrzkToiyBaAuKtjpibQMXXpWv/CTfUjexsDOnyAxKoHSxwcgrTle6VAqJjy
M8XZEYCLQ8IdZgzwpfncKsSObGz8Vyg/5+vXbwB9XA4sAp5j0ztwJL6ST950T4hm
yMtC4BTUUOldnLYJG6phtdZ3kOEdXcp3H3vSZFWwfxtC3PVtLX/fZVAX+1WlMoDC
IIAK90pVdBQ7c4I6q3o2x6giDy3xh9z4bTZT4Y1ryQSEfmfaPpEnixkXD9wNTpGr
uhJp9rr5IU6aobpLIn7bWAHB1qHmXcYSlbZwo0fRpOd4vr4eSCIVb+1R9Rrpts3y
SC+y1XuwQsmn+67FgA/8QCEfLffmqTJ98agBb5XvXj6+rN1XKuo/86I2ppwgLX5U
4fMUQvCJf5ZzzxTzXhVpVGQ3mnVrSGiEOm9TOatRb5D2rZHuSJcc0byXb01DsNs9
Hj01FrBOqazWdU4AP08YIYX1rvA+9XiIY571+6htAuTiFObcRH9ob5j479KDw+Du
EFuhOUKKgaWHsU5pE5gfjBCTI0Dgi4UBBkl+wxg1f1P2zrZY5e3H3VEMLVmEpLTh
vpt1laspwfISmCojDKVH0qXlOLVtG9tz9yOZyx5qFq/m7GpZc8EfvLqgUFHqLYDa
dRGntphl2yDvZQYO8FSV/wBQAZJ13CSSYGO2YlVz+Uh30UNd8AiU0oUtAtUjYCpn
ekTzFPx3irE1IafkAb7iMSov8JGToo/XbQ3DtBHf2Z+muwSrm/10JYu2orv8LC3f
EkAsICKk0mB2aLY8qGmLO3+F3b5W87ZbcBz2a1PxIFSxj2NrTPub9d8Hs7AztvOT
CoiPEH73x9UmI3lAW5cRGUPcFTQDp56Gr1k9oj9grbl6PMkVAUstmItB3aB0NJEd
i4Q4+H7i9UKQNuZvUiAmC0glUwfqRCdR+kakrKBtixIeuoGJTCcZa8WYarHNTq+5
ghnJD8XQkXRzKwpe499KAm8UE0ZhfBPiPrWnE8g8rl5+wjCFFJz0sKbLGh4pmyvC
6rdi1rRMViKxOloNk9q6s2eNiaQHvtRsR5X6DyhcCQ/oiqUEgIaPkn+3UjKaFpGA
Ubve43d7IJ4FXkqtJJ7V/OtbFvJWVuKV/5ONm4TTE4dw/utXrhdkUflsxd9ORZp/
+Bx1JfPwiO8Ffz9j2RKpOPaagKJry84jJY8pEu1fA7c3qGUviMU1xTnE+LYtf+4/
6xlPH193deD1NvU1uy4e6VJXkTbcknds2C65Y/m+B5jGq9f8HHN079UoND6r2biO
27StkEHQyuJfavW0WYMZQzBj61m7z2BfyGI5xfcQfSO4dE0rpNBR7de4EP90Fep1
AxwlBLMMZUkePBXCQghoqSaSl82bE/sw9ePmblOSmAkERvaHShcwr1wS6yH6qB0r
6cdr3SvNj6BbyIiY6a7jKv0/+cyuQIFgUX0heToE741cWLrLbWoEhwBL3dJ/l68+
bbOFoJb1CDSG3HD3/e6UUuzmOW03uTKT46GfmsVt/AFt5ox7GB3rGod9AtPaTm7Z
qfZ7sanh1oiilggKIFtmMjXlkNsHiMnXCnT5Y0jbqxywJS8lnksEgLlNWrEvl9mg
3LAW++L9vbNESARCOHesd1vqLUM6l/ERd8jIgxgHtCILc/eItaV/wm5HzG5o0wij
HQXH9Mu3otphbly/VJo2gXmllaNNf68StjrbnqF0Mh5/xRn2TgsBMAvq1iHSW4Gf
i8VF9nvWFt1VpzHYmr6ooTqCfgpZhob8gBBLUwGU4k0/BLWapESV4Wtl30SX+bFk
64fOgUVbOLqQmPOBbc+CfiSvQACd8qXs63ZmGmTSEPKMqolWw/zfmhLjYvvBKe6x
2rpYY6M4pPg/pbnKMyYGdnidfZuiseAGYjSR6eHb69AbVvvhhLcvW3K9bSxHaIYf
Uy8zRhrJ9OlZaLIUyegMzENGKm0o2Y+8aMt4JBEcrSo1BoizNI67ycebm16r/FKV
v0778l/kYbGLOlXacnIs0+vsAwJgZ6h+gHuWNzZJkzilvk1HRebT/uB5wgwnQzi8
lrzPLPRhadMIMWbTZ8W+bWXrkeDsIv38LHNvkONGIn4/cpASDQOivcSXuPcwcI8y
k6Stsnj8OB5HZcgDoCv5nLcwC6sHJ9RFe0GkX1WU6pduEaks2EF4Qq8MTh3UBQcS
aEa4akG6aexoTfXvn6yToCe1/0MpTd3sRactcbaLm0s1/mi1grO4iUz9P2cgKfcm
CP8NJsKO7IS9KDrx5St286o4bfVhYOTznqf5jCvvDodtv31Mve54lrSZbi192hVs
fdIiG101WpFXo0bZ9XZOxSAddGfFfFRxCuVSw3wqCXY151zGKMSkfI5vbxZWME+M
+aEMIHTNxa3VkhUZy7JN74Mu5AjV2wu1GhynTDAt2uz8a539zE5n1rpL1DMnVlxF
B+BTv09j1AYCJfZpnrLSON7JhNWRk8G7ws9+FBrnZ/LS6PbJQJ0jufg2qNwZdxQZ
yX02JfZaAY9FZW4LveoRyhp6sFlo6Ck2y76iJaK980063FJ8YhI780vW6ytMJkIA
boGAFARszBl2qd0vhZ5vCJ5reAka9EP1N9lyZBFhKI4SfYEyj98XQX2CWDoQnGyq
0aTlgjvXqYVgH2zHxBfL45r8jyH6nF5qYHWiywOPQYj6JumOn0NXkSoHPR5n++2L
AHdYqSDOO47zWU+cifSLohnqxrRapKFBtOysg/KMfm2fBswVUdiBq+izXiIvqdG5
uRVjaTYm3fx7mUYYODYl1ig1y2cJBtZE+0mondLMdmEJAP9a423zzaeOS1hh3tQf
WCH2/sWQjyHf9q0c+5Rm+tp5S9TvkbpoD50Xzpa6eb6ijm1KDzIL28G31965bOys
Xv4Qdv2lEzy6EwL+wp858YXANxlVAMII9FmkDnDmFudlTqul8TCAb8SrmL0FCthO
Paz3t8uWqHsX8HDD2r/gVHtvVul7Nnv2KZzwfE/jcOJxZYlG31NYm2MpNcjY7lFt
6nz57DQOMC+PlzLg/uVPtLSttEH2WyD4iXuWSnsMv1Ek+eEJ24Z5cXV/GVBp7WJQ
Nwqge98J4EBSycalBiFJwrhxeG3+AhAd7XD8zfbeVnLUiUFj34cwmn7W7Mh75P29
+FXeTq9IbxfAPW1jw4GvO3qbPw1aMNfiIHIk7J5P/JmRCNZKwFrQUTGp+9nz+0x8
/B9IJWEJI5JjEQ8ssMJ3zL7/RpUoTBEfB+fD52aoy/x0iTqsdYrmKa57Wu8eUP1O
T55B8IAP8FIzZb4aO6IfresLcIQKCQv/b6WYXaVFK8M8OirizxYClSYxYMdeaS/9
YzdGun1M3ewYpWu2NPPSlxplbFMakjM5QNLtn/iE3OxX9Pu2dpyrO/7lzJDnpeVT
xrZ7DxpRW99EevDOufKS+F1iFLOoFv5Uq+cS8zaTbwsECqF+EnMb7pbfaLyuBrw6
R57qDKLBoNIjVUM7G+MJ9PEPJMFluYe+P+pi5RFh+9OhXJr89sNrdwACsXA0/5dq
eGVpHgghA5DHxTh2NNtr6s5XH2kzmHAHUSxyv7+JEjfVLD3NJ3DYwiPqpwRJhxWo
Seloh9P+uN5uXIQV8+GQRbfsc/XGuI2mibFTQg8NutfHRUAutBVFPurnd7no3duT
9Z4y9UfnUyaGuUY2pHA95wjwNXYftjnQpkdeslphINmhTWxoF7/BLCGdE2exrOWJ
1DT9fDq1gKKOKFsabM02zhgzIINXhwd0PWLYKNMJlVdSRDMa0c2NdqOMyHF5ACxj
z/O4sHu/LQA0+4jVs541ndFxF+W6K6Cn1YxM00SXcEfxNam20qfyj3L04jp5T4W+
uQzdJHYoLDITdGaYum5yCXP+Q/I5f7II56L8Es6gJkbByRRalH1h7C9mycrvGGz3
ByZfH4FI/HQjchbmuDMK7IDAwfJGiiUqpouW/1cu6KYi3pFya8oZgiosHP4g9F2E
i9lMUBNiZPWngeptBdFtspU1UVcoErlDFIHB11v+4Ten8PaHw03MCxcLj2/z2PRh
yM5un9+EZiKBoAaHpVZvqWNZMed2qd8YT6aTLh1ddreOm80exayVfQI05IoqE4WT
OyT/BdHTEC545jWUZBT6fX4/ABSJ1zdYoOl6+GPXA7aFEs5zSyia8wVkYLO7vlHZ
nz6/TSvzeEAfeov65HBWnN8bNEEwLTvw4XxytzP3SBvDikwTwCWPQAJ+su3yKUzQ
Ms7LT9eew2N/7BmJfBMicbv/38gF9rTRBgZlVUgAThQr1VCMrRpZxnqQ9Ui52NBt
jIukI05ukLrWXANfxPw5/7ljC5d2shDKYm7daloc03FAHk4zVkfzVt01sDx1CARB
/Cl0GIFJlQvEvgPtV6whKjZFzmxXZn9hrNaLMxh9Y/MdjyHK21VqTHLa/KtrscJz
0eeUcWttlJXQd+jXsKDFqR/XLkFUbvuVq+NDlya/Dgw0VFOJkvQ/zLaQ/tXP+xge
CoJG8NqO5CP8OR8paSX+1BkyC0FJFRfbH8aaM4YTYeKQsOdMcVjIQPJNqhN3pT1l
mNFUYWkqJ1IUeyEWtcZDZSkgjkpeLUqibrJzlOA6MmEkpXdYGhFaDkK6M7OC0oyT
tAsadCf279uBgvXw4lFe5NEXHqc7ySoWpbCaJtxavYlzbVECGtrIdhyA+Ija/ssm
k7RHdu15D80wqipTums0knGlITyON/B5wrLAvTWD8s/g6LAAFbCoHstB9+bqt5e8
7QHA3xo1DVvkGUqJ7f5a8zBc3eWbqzZLSWyklxwwFfg6rfu3FPlivZNEbA3ElYmq
+4iAfuCgE5wdo4lkvm756Cc6npxpZptE5Nby4cWNxWrQObFG0eAUxEZzfN8h6hSz
3A5/k/NEe0Q5ChQNK+W7wu0Tusirn4Hmiqw1RYbcwEOumS50GYpjuvYsE+AsCGHl
DS3755BbybzCLUhPvp/cQ8ia6lHFfDF0HYv9IKV/Nhg4UXOQJcKhvDBYGlbLf2ot
Os+gGi49cGe4iaspXFGMUm22zzBUK+/84THFRqxONHJ7W/xKZmw03jIs9wQdY7KA
smFnK/TYQ2m7xLnDB2kaEL/GY7/wkgprf0/fPlvaL4uYD2K7C1TUm0637l2vAk0D
W8tob9Mu94+ujJfJAENjbWLZ32k80BJKow5FxNnEO+XxTI48gGLZ9B1LZsQCLl/9
Twot3app8ku1Sm2Ej5LesG9Csg5MIK/+f7U1DoJoXuj3qxifNRZ7aaG3Y5ROfbhp
CFtSmedzAOx+mk+Lfn8e0J7NqVa5MnWaNJrkoBuLKNz4MyJAgisIRgCYWWtrc/OS
Ra5bOZsEG0/d2FXGcLNqfQoIX+bmDJtx2Zs9gShpOraEBx4clZBpzmkJ2x60KVEE
+IzFsGeUpfuhYicD1lX69Dxh7aNiHrTXNXKr5hLMrxKzLY/Ec+v6xVilS0PtjyqC
YABAN8IDZrLCbp+9bk+Tr3MiVgmozXMzXa+RXg5DYYaiE6BG6GTQJuHnV2XrzCk0
6HT5pscjjFw/lBZ7jksej9bF1Fije/ScKyn3uqgHmo3RdSSlHEzCs81YmSmJTuxQ
cEXdPIPrNBSxqr9QmDirNDweoSx8/ahnxa4NOF0WvAcTxVu8aizzq+BCRo8Rxlx8
dMUHXMWjDWStC8okYmpoZpQTYYGRzSUQIXXDZKGo2gtbpeuwnDOnVpiZZaVZFhPs
eBb7MZwUQfTnXmrrDQSoxk0kn/ZQI/mOapVk+i2XH6X7AesOYHw+JJeIH0TrEgS3
AOcu1C9mfMtKPKMRWcfVelDFSJPd7KLltwM7xasmqU8qMAkCBsDBOTWvqQ7BEF2X
XWh6q7QNyG9HFKkgh3lITv/TwmLBgs9EIyFmN/5N1XMpp1ZgcSIpn1La3LW2Uz8t
RYlwXZ7QlIRX1NYeZdVLWqM2SxTkU5yL4JxggXh7aXJ4tzJL9NJFuXulC+RNPJgJ
PT6HrGGlXxy8n1k6joGoYduzshB9LRsUXYgVel+wum4bjHba7bUnDOrOL/lYN8fW
1GNnL9bhTVEQ3dIoveXvfroJYbSfD8E2fSYNrEmX87vfiTziKeYeyZt3NbduqevC
Am3Ijx69PoQf9oLgZqYHjJOipxTir2gk0MTc8fTAR/dFGt8ObVQlDZDJH1Uw2F23
svuRey6psxhZhk6mD5drq+YJPuU/sqgtthJN/1LeUYGDHuqe3ZOi2ueUo5JTv6iN
gc+O+jZ8/xNzWKNt/jAvS4Axm/vudy+SU0Wo3RiNuY9ZZc0OQYnazni3xSEjy8rS
NzYwat+V4KSEagzyh0oQV77yKWmDkBePQbfnghD3jKQl1Apl9aD7iBhPWq3Rvnu8
w1tchftCuiIrnga+cXlMrn8efyCmRZM1KV2zo7JpUhQAkzPb+PVqX63FIPkENSvR
mN8g8DxUy0SFk5Ygjo++SNos4NbqpPrkwre8JTAFTfKkZB7WJajrsZrI/0zbhWqG
90TgDz3iBEuijQQutoCifm+2hrkj3JLpw3bkmwKavM1RMaKIwV5ZRIdX0/CBiSMr
BeaPobDm+UawgXUdnMFmGBBI3n6PL3T2Nbs3UjmxBx13jvDjV0vCOAO2cv1oSJiv
9JM7lh044jW+tklOlNpujT4zgBQgm5SX+grk5oIDqZsD8wZ1JOCuod3D2OMCPMHs
vOLIAzb9oGQtV77DY9d8q0uazqY00YdSAGjn5NGStI+8q7Cq1nAe9Hw3+DVxjoWx
1/RE/F3zM40HTKuv4VpG+O16Gu/oT2tGjcaIh7t29AsGwiX8woQi72a7YVJB0CP9
K1ShUmy1MUiS0/GiypjLj/v9VFCmxqLYrhbkBzxLn8MF1ayipkkY4jeJ9W3OduPl
+G7istG+H2co5UlbnyDPkk8WvsvwvKGbHzZyi51fD+TdfHglHYmpseISGgn9/Owa
MThByECIbgmKaMOFQha+31hdW6FEDBzuWr0nwJW7De03uGHtqyfwJlOCZV3R1w13
6WCzUHjt469TJj8lA2+JavKhRUNdxfMhHUx5XRlgC2YjFJdOOgUvC+bDgsoCkPbM
n91iEaL3K/Lt/uC7Nb9l2tgx5PcXYJK89Xxw2p8LWvgFfPQskjGrQRdtR+YkxMhS
YWOfhe4fifAyjlki7HzPd2jzTxTnvAWgOsjovneYXUM0pjzFuzjcrWuEWE1T1DQk
z5z+jhMoFrChoBSGI3yq3G7D2TtgL5Fo5nbfOogjpAP3ZHpt8AKGfMCQ6AIK7Y0r
0mIb/Ih9VzCPR2PHmuAGgAc0vH7FmS9pHV8Dl+S0CcbDihaMEWQiTgBjDzEUHyXm
MjpuAjmf9cRjrlCf43/ofT2aZh6vUOVhyx81t85bxoGfvstdbgLonOstP0VPxi4M
1UZ/L99X8YSRdbMtwPBLEYSJg6LK4hAC/SqTFHXYr57XxDknaQBvIJbJmXloZGM2
hwCdZoDaJqLWQfC0uZWozCpI5f/EBxpgpacodNP3dXfqeTnL+tMYuhpvs4yjF1sB
iDGO4fIbC/pWTl5qfKC5JBvL3876KrbI4nLZhcIyjwLGjBO6Cbb8L42dkfW8MlPH
XLxhXx3pDQMfO1eFT3J6ndr0DHBCL7IOfiKhvYwNXqoxe3qJoN4JHZEVM2w5A0aF
Kja+hnxEiQqVEVgzEKibIABPmPA0POcR+q7TsGrAn/duxAJN3LIga8hkixINcTr9
pVi1HzK7xsoi52qgq/W38MG3uf8umErF/dv8PzA96/tucocao7C1/jnkoNekfArM
LkASQzu2ZKBx3VAnfQ6K49ATyWXHH2icCnlZsIFFNCikXKecjqs6P2UjHDJ77GUv
a2BSobybHWfH+P+uqnvhkuLnS5PKChdF33xgH5rBZ/m12aASCVplbJ6ulPqUE+VB
CalB2DtUs3AEJ1zCXutmab5teUEy3yInI2kiWkTmoFKKt/lyJZBw/+Lv3pvQ1JUd
br9vop6Iw419YG+q/MDwnanAaR47qAGrQFiQzeZJRJ9e4v09BTc7zy1K6uYB1IlX
PUSvqqeAspqWnF1vTFB5nkUBjsffgjKaFkDkVNWEGfglJuefjrb5y7BKxm2agsx0
yiDArAGNy8e9kPd4fV6/lfY6sdc2tVusryCSIHgA3vX0C1iKik6Zo72JUOt/bnFt
QibQFZYbs/G+HBnYNvcXwHINeK788kIp+ORuGXW7gY/4YoH8pGipV+PMhTa0l0rN
7StuMAWzn6nP/EEd1Q9+Jkbt1prsVHpD0WMyC8x8UG2dKVlsMC7Zy5gRp1MNC6xC
9kVQxAZNAudjUBPMKeVvx8AX0QY50ZEKuod7xThi8zssdhE0U2wYBHhTPrTNLeGR
GTDrAA97EiyRl+raw//evDMLpvH1WpJKiXkWnkCCUIwLMCyWY6FdbmJ/N9HVfrsA
KQLvuUssrkuzfHqE5qCib0EP3sOHJaDFCxUO+3O+7y4NmwEZz13ySGMuOSMeJoG8
5tSXH03SSG+yzTihoI41qJsZ5iphhBHYED1QzQ1FYtaE5hJgnW2PDpzCgG+5J8dl
6j2bMRmS6+c/aZsoOzQeoO0hALIoF6EBxuvQGCdJ2FNLZmL96TsYPDeK5Ogq8vY+
ELy+uniXxMDgdjD5O1HszKuXGexsyHJuzBSUbRseeZGiEcZBi75LA8DU8rhApu3V
M/s4G8YyGQFcFlWwMgpNAGz/kDOrcpiDdMtT/sFnTcqFe3HhihDTl5HKnHKNqvwa
d3uDzPATGb0xwkQPS1r4YGjQFX/55JX6oNgBPPW/ENbRRziMPcn6pfdg5zvY4oUq
zTHEGb/klB3UzPBmd+zcJexNCM2jYVf9V/CpLQL21yVQlLPw2VqyNngRW4SYzJTV
1ydWVUCL1Fp0bLdIc/Zjk8iMlH6ktSWK6oHgvwpNlnGZo8Ll+IXstlRSZWv/YwmL
12oGJoa++BXvI91FGf3yDY2bEVOnwP6sDyi9CtZtgA6EoULGoT+4v2mEucRwJiyb
1umeCpMIOxqzf20c7NlsIhIj/JBv2aCfo5lR9Cj19cuCy6hT6AmnUdHqzfQsWrL0
mqiP3LmnF54qu/iM9B99ru756MzVHMUngtasZtul5056iklSnD61jqtdrlUw2GZo
HarWjkEE49hzLNs34acawja21LJe1LrEcxPKRxAIQe7d4gf/Z4mHZOA9LGzCrXpu
CoyH36rruwgCLWYf+WoxzRGmB5odqpguFrFYZ07lpxJeS1QjDvH4GCtqH55PkrS7
4aPrQVdY3YNGjXK3a50xubILGdHpTggfhWON6cjc0ylDq7bnENkNNX4MOjNx3qew
YlL0ufXRvUAheOVyafm3MEq9inoGanY8ZMf9Ei7TumRpGwLUPPkfr1zDzcJIFpiY
E9BXqVX9j4STHqidpPxmLfylV5Bk5Ytx+pJjQSGlqsB2Ks+XgLS6eFPaDK+VCuFL
nTcwSgkkJKCyjRNDmxWAckO8eoaDClpkkSX47sjSoFrOwDuntoV+r7opR7RiTN++
IdHWpfxNEC1O60W/oVJ69/5ZcPxkes2IKhpqxUjJaEROryRXQwR70SSx5buEJOBj
VKUPRR3p4oUnTioauFJ/Kz1Ayo94VVsiUYWeqeFHKOMC3VGpkBBJhideWZecYyd7
4pCQZVgbl1lxe5pDgF8f5MGdEU50bitX7ySwEYxBEvIz5kYuTrFLtrcEvG2GMZxo
7tJz5MjiHZnzFkR8D/zJWcyjYtwE/kmlK1plxMik1qpa1NIeqCboevTJryZGZXqb
LZdBsoVadNePTLbfPZ9Hh2OB3MJKtcKcpcWoM6K1lWrQ/qduABb5yPaaBwX0OKnw
1t7m5TW9h2vq0/8CsIcy1ViwxJsPVdjEa+j2dNe4lyEJwHntkWHckLul754egaEw
7dpbG8x0rhObYXE+NdKuG4u47JD7o4tKDJL4xrcwWnuZkVlyEqNx1ZiQ+N7OkXKY
xY+rbRk82Q2PZSCFHXR/987iXD3abERBTdIz8WLyBkkB8NOkUW0Z6DydXf9PHmcf
ke0HR7m3MZ9/xDJULp8HWA1QryAomjRL5+7HKRyVx7fYgbx7pDpc7RGp7tNwK1Ss
pZSHq1ZQ05vqrFSsF/mOeOsZMoGCbO8YghlNiQ6abWMvNSgJ915Ay39jF3k4IgNZ
cT36dEcWlkZVA1loV/4QhCWQGUnAx2skBGzaqEaRim8O+d67P2ajSqzecG2xbKzK
nL5GB8G3aZ2TpFSz7d71H5/BVpyg8XLxaUqBqyqIo/wVVRf+sNSkDInUvb6ULyS8
y5DchYZyxlbKf2eHwPTmcIr5W37ohEfU7MR7Yy3kFeEQXUX+ih23IivImHwOx0ax
aDPWExWM63gS+ft+TpGp/nzXIrLHzXFhjvyerTwZE6zbWzJddBWPvlCs2sCKRRkp
XWFKcv0TT2JHfntoHXpTZNgd/PFvN2tZ5p6xg4eM2avLgwtffNWGdNoO6UNR7y+q
WVGmlbZVqSyyDHPMMBP4fl7Gl9yDqlw2aRPoUAAJnQP9mH5AfwqH/w9PbZMTeqqz
ED3MVgtKBxABcLESXxgjlf0GL5xYU+OEyVo6b187FdQEeTqHfnaYRgNMj+lPTeNm
BRkcHz2Lt92lEQsDBSzL/Qnh/HglXwfDVjh2xs2B1HCONqDIfr0+WgIPrkewwf3Q
K+UjoTWlKMjAZS3Py0GbH0q985oP/moA/U4GQTZka2wEAIsBP7t+a/vcbA0doARp
rC8l3QaXN7GoR5+3f0DxX8Ah525pNbJpicqkeNKMMuSThyYoydgzRooGUepbyw4x
v2ABEnf6eArbU195YldQdQ60nNdTFEENfUA3vUGg/P+kRot9Vyoh3Vam3O8h3ul+
o5r4q9vcrVZQUHxkt9jjnapueHCyDn7wSeGR9gLUzFgSW/3i9QAhSbVIxDiFoKMh
1KlHVJbVHLsS+5OU79zIP16rYJy4MtzXiM52qXd3RLMvpZib/2j8/hdOv/2Sqnh+
+2tRgIzjNNC2qbfNR+pvGYfoILECctKlxEMgH6eIqWwDZMTHahKqyEXXK0gx1Goy
q/i7tI0KWR+VzqFfXU4HPp4h6MGI77cLWGSOUycLsVUIiALjqaZ+hdr9m776dOZK
frN4OcAxISwAlkDVLVyEBtyp10xavw7RgAwhk88kguBcG1Xgn07yBTP0vqclV/TD
Pn/S65PuyAt8+LPZcdpQb9QV48TCj9y7GJYo5PL8spMIZJDAv+mFU/HKTC1tubxS
qxFDz4D0PRO6FekUhFgOIcXKq5zIQYjbPzKx1Mm9dKtMTHl2Fg66Lmx/zTU88G7l
R1Yve3yoh3NWVzCoJMjiCjqcWzuZsespk0/XzV5rJJMH8P7OO6n6dBBsRb4aKAKB
QQEwTx982M4KsOfIyMPdJLlBj0kmHM2l+jqthqnk1+XtCdMrwcBDngSTGGgUqlwk
lpv0gg0CO6Jt+6hz698DPyzENIwyqBpaJ7TYjlFl0jcrBINkXTk+t/ifxUrJWg4t
XwtoiyF7zNZqDGD4Cra7ku2QqJAo2h/GRCWdIxVFgBruLrWLGNcz5SjMOySyfNnf
fa7/IGNVlICnGxLBN6UAOoWcSsNTTWZCwTfL1IRQNVEof5fsJatFkYgRwXQ3SIHl
6fNL79MPCoWAuYZBlbJfs7L/Fs/F6F7n1wO8sGE5amCK1yOcmszM7XKf0iOJMCF4
quN6/se7YlkgroVfLMspzdb5MpuXD8YKLmwXaF+p4TF9V5Hvd8C95xfpGr/+e1hT
sGGM7eA0TM/isqgphiQyWoQcuAo9Dx+i9RLIsuch+XFMhhnU65Lgz7VD7zvfFZ4x
rDYiLDwL7FUqPtl5j4XTNhYer6GFljJBrv7R9Pk0AHcYhlsEeA9PedZkC/TH0RF4
wTQU3xIk4wqBdatisi55Tfk0mbGAUAB3v6lMb48fjvGhupgiiEePSgq9EwJQj7yA
lW0Io9jNe1FIN5f0heKpAo931OSCdkXIUPNLlysdjnQUrORFF8OM3LxdY74haoze
nmIguMNFKGIwhmkYnesC+8t4jIbL16cANzrAwsqX0N1paJZGPaYEGTOpjssAXp8F
OZhVIbR2zw1UCg+TbCvi8zisX/yep6Ht4Gk+FhXv1nPhUzKBE3sDrCNZMzg43XS8
TmeWqVf5aP8wcGTokoTa1ndys/pSCHgNoYgZPMgL2nXVyh2vqipHbeE4hYnknsWW
vOlkMPrR6eP16bkZiazRpCOC/+sNuiMCXwQe/68Yld5/mP60G9U2lyKXYO9aAjy5
aQeJR4N18A4lvOZJbkOxZzKA59roLxccLce7Z0ZZSKxGCDTt5EHLjwjqU+pu/Z2e
2/rwe47AKvDeqSm/sM8f1igkMI2h7Y/SqUzlPNIpoIah9HMmVzrShuyDJcAFva6x
Ompv30H6T0AMd3eCTw8apjCJXUXq1Xw8/r3GEAzwdH1YfFb66g8jwfP8LfAH6vxl
mrPeeDijOtuyPRTXLmSQG+QvUyZDxUGRNBw76n4pQ4C75KAc/4657riqrdaKdy72
0GNktvulX3BSovuk3IRYYkDwIUINewuBVinPQGxZCgOtEV4DbFheu25bQLhq33n9
s3pMFs+WQ2aqcbKYjHTXhuHarzuFtvKzk97sn1zXQDSJ4GJtzQfOFvCohsVCafkL
/h89zFa5jShnxP0YyVdgx5nGTzHLrJt4EY3o0/p1vb/yn2y9M2lbXDGy+lMZfjNh
vZRNMNpmDTfyVJBaDv549q+N6ZjMWgXQP7Gm8VyauLkjkFMJVbglSqSStF1SCRT4
H2Clgu6DyCymd046vJALs/sc+TG6DHD4vPRcybTmvJYiNAx/Yq4uBqwxo65dneAM
h7oZ46GVCS8oZ+Q6+TPF38Vr29jAJYGg2cNv63dPRqSm6tMigBvGj1BxMY7eMJJf
0p/WMoBVLkabq2uypgRAc32+KzhkTf7x0BFwr0s/XdikOiF52KOj6ClxLcian2B+
yvDo71x0F0HFzjjYTY7IfWxSxGQOJCw/YQ1H70Js0g3eQ0obZZC5fyWzWnCDmRC8
RNY4Cki64ZpwewbxCEjXTvI9vYo1DLS8VheODArOdAdcOGjekbAFIS6ZbcdHxGwr
qcILmUhr8jtpLi2BoRfFM6UBPXJodsJTq4cwu28N+S7rdDbfHA3/vnvwOoL6jObL
RaU8Y1Etilj233CquTjpTkUWv+slsz5jhTOX7QcoECJxh2aPIzJ+5v3q8L08GC26
OgT5JLRsRJF+J7/rl0eugXwvOOgF4toV7e2FK7xr0Tw9quKfXHFGci1k8xYNVpQe
81LhjRknS8MLJ9XPGznKl/Gua7rGHZUvFJysHbFX0Tom2Cb3JqkutcJdlcHbUVP9
raPYlYA9u/S/TNZe6leJRFVehrAss7nDJLbuzk3fSE9srilAoP/bZa1lkonxl5Bu
TFyPy+bCYyW14MDKy5KOp/Cv+T+aaT/iB5olAKsQ+qAyG4qk6eojqB2h7usCTiQ4
YZVJl7OTNIznzb7Pj1a0jSN14LWqOzjcP0TtnqCtkGk1gGuJZ+4/X625154F9XO1
A5iv2eaKRRkvgK9tv0Ug1Z51kcDytrCQZKTA68rFPPYPTHMMHJAJX9J0FFiMgrqm
H/P1rsWjJqhiO81rrZAm+KCPerFP5n5PxrWqhXwH905vtjxQlOwq25Flm30DhNMf
F8oJRmGTwNS8cT0u1EH7UcacFjD5y47KMu3/jzcSRFGeObwdvcbu+81IQDTph615
qck+FO1uRIR4iumVP4gUYDr4RtZ3Sk/Bh27rcd9mYyr/7tBo1UDMhT7HfzJ/QOBd
NwVAtUi3iS4pdLqE9smE8cAlesIXWIipwXk5Ao4DNS8TE26H/Tm1VXJNaFpo1oy3
mO6I/bccyObMbtowsWrcVkykJwrxPG+2mlvK4EoNsnqkTdAkLKclTAyZSlVRm7cT
cOd9bKXnRIYq6ewapFi9kyb+oMBm3466Q8V7ETMlYmX91HzmDmKS5XGKK0iP9kW7
m4TAKCGQ4VwaLjpG9tksLTxLSJzLG/sh33RGTG1X0axv5sdzmcivRdAX9//oZIRo
eSe6pNNPwTUzdJ4p2itgKWqq/PTTQ4LrKoIGAqLjRw4PGEgiJihjOGd4nMhMBFSP
pceEjmzPuExzRdHLZuMisb/m54fn6TcX/QPWJFmzakEneqhmRorb+MfxFBJmHJth
eeyHhpFvgtdLu78gjGyilw3de8moAYkWgpxbXySQYsR/FVpvuKMtwx+YNjLu1Xvr
0Y5X0r1IDvW8V1tE+4I0jJD9lJiIoJFKaXQ7clnLUJo4sXB6jcfzoOonD8aGRiu1
b/n6iWL2z1o6m6bV0v7IeyynPXl1/v/4qf+AcnjPwS3wtybrxm6cvk7sr1Z6IyBW
JvL96GvzM5+1kLUQfo2IMZ8txx0p8KLpF/6iuuMrEIn+u4CLhsBrIWTDmtZRSZFh
jYDbIzLVM808P8+na7mxqvJ8j5iJw/ee4/2EoiqZ99eeUpuHGB+rq8idAuOzPEbq
4yohOC20MaWBZr5YklxdwBKGw8YmqzuMeFJ5VyObFamYtdCtgcXqxGE7ARt7c68V
kb8+86dbicM3PngLt8NtiNkkOz5+ZBDpnxOrkJzL/KX+w/rnkeiLJkBVBH+rEaVr
7EtAF4eH5vP+JSByxq5uStgJFEnUsdD6aMv7+LLYPN9j0/XS/irlZLQmxYJ+TMCA
2mDyCUD7RE8Q3bnNoIzaxjnFuFdt6CBDQi62qD+8gKGAxOCzIy9j0IFkjIvSpZAt
IwW/DIjHw58Yx1101K0y57iHYEU3+cOenZYYUMLl71VgR1vKMxRspoCmtGDW7riK
t7pZHk0ugwpz8sY6yijpUKb6z/lkt1XOU69SooJyJ0yHE6Yxx/2R7DhhFWlS8Tyh
YRPEQaYZGuuIKz0NNOpnOXAvwQp9LHstmyPoP3+quZgLcO4gtqe/91wZXM8HELfQ
t8Lj33H66HczhUp2NTPpmZh+dcWYNjjjrnwomOLAvN9aJnF8M/MY1ydn3f/PnH8f
z5QIdTN+SIm+2dd7/YPe5ulE/gSVHKLQVrowRq4ENgCt5WsSJPCphf1FaoDG1Jx+
JQ3xT2CjZ3A/RX6JMFMP4QBrU/vBAUm0fBGDAJ+fRXBStfWra59kH5SBx1M9HOFe
Fyg7oG4TWFxfpMa2+wOdLRo60ThMZkklET9K//pw59M+Xi6dzr13R/3HLhi/sO0R
5/eRgnnxYL92OaFXG9KTCwy8SI9VeXKh3Kogbxtd5IfHz/Qi36mKz5y/X91KMQzS
4wUuXTqiQiOKJucYr/74glD5JCdtSFOto0m01McgSHejPAUIBzDe1bSyKoXkzZpf
fgAPQvEVCYBZl1e7xJoYE1aM/es2AiOA8yb9DxONOIEtx+P6/V845Tsgo08Zt8+o
QQuXfmIzqODX+AtugvrrBPXQHypIHPvxSAwC7IcL1kSkx2SWKTERZkiph7/mbup7
VvKVcConUs3vGIvfKORWL3i6GY2UDeX7r6CCw1czCv4Nl0/v1pZgpkQV9dvuo23G
87gkf0Mzaup2C7M7Pj8/3J2IYRlvPnS42iQ2VAMaYRL7s7qTMDg1vJWpvYs0VA/d
Ry7oWFDBq8kK/RJQNrg3Mf85+nl3i/MdhJCEXTo80xqY/B7ZUyIy5olsnQLEgAGH
sGQB9sRx+hN4auKc6pcNZ9AGPBp8CgtASZN7KUeIL7nZzHgB1x0nHkaIS3AU6pYF
7V15BmpGkVvZyO5C2ccTWXl0Qp45yignVtsu7w8MvqIyco3i7i0FlABuB6yL2leh
8RC22UTYTUcpawntKuFvaUaYV8cpDyv7IPTzFQ37eLM824128B5mE0XoYbzg3n3n
VlEMoL9yAHOEISAaXvAtkYZb8dQT30g5Sp9dxi5a8OqvhOns9AhZSIE9Go8zpI2Y
QorgDEcKUkvWy6CMGBCfSNFPnojeIh+aQCoMi66ekQH4PGDBcBEcy+bPqISFoD3m
Q87mr7+XWnqjRovwTMm8HU8HMac53u67mPsBwf+FozLyxtnDyy/9U9Fdz5xX20ZC
QI7FhNXRY6gqTM4ZhgtJ11Towy3+i/ouHTsro3BfFcnynMmrM5oPc0tSunybQS/0
91qgHCymbCYAsHPKf3VljgESO9oxRUcRFPzicm2DuIYEDwbE4Ry4Otvswy2jjhCF
IEHnIjN0++ufiB0weUsPx/ie+q3er9RxlU3fRXb6jCh0nAt/nziwn54oaH9eTsd3
8+8WJ4CykENRDXHY4Gp6moK1az5u6RdQfQ2Xflf47GVL3PqJPfmA+OiXga0Hk0eZ
gamq9gwigk1cII52830gOs/kU/kSmAGuLrRTSRGUCmGNKHQiszpzMelJ1fyotVDp
y0+vrtijfWjZjCk7DJ7dbwFbNKxvzSqtw6qY0k9APS0CuUvKjN24cSgziCiQNfB6
5e5SrCXK5GALu3z5BMXcqV1UU/miAlWhT9NjIEFJW+WSZeBdpvVoOcWQm0xpRZDe
FhFXO+kQEOqL4BB2Ei6TMfC9yraHQE6RdQyHA3ktS9MdoYtvswAzuyvJB1GLnixd
37cmXtyx+cyjrvHBce/WoApMhwQkCdgHPci44Ufv03W13TrWZdr+LuUEKeMCcYxr
vE78t3yYoxbF+35Z0T0/5+KLkXhbi8UENIyYe9ZnD0hy9bcwnQ0O5TuMMUXfyXxn
bFBrjNpu5cehXtOyxrf3sWFIhpeU/Fx+46JwZ7/ASE3tj5qCq+cg6+p2+AHP/r2e
3qlHInO2IP9mA4aVO15qfscggvaZAeBKyuxMD125u92ZDSMZo0EWHpJJ1LcOTm3z
HgNIw9mOJyXC3+7O567sAt0EtpX/fMSKFgoo1BMqtXlHF6a0iO7qC+W6zKJea0O2
tS3Ac+/r8czxl+KPffgnD4ksR83NfEoHDSqsFWk4apgpSTmD2mADhOgf9sjOcQp4
7R4uyBZnjjtOxEeb39OQWXknuA0hBWsDjSq9y0wlHOONlHv/yAiIj5srXi/qWdm8
A4HaytMvjOfhQT24nLA1ympduVRMjaOONtvdqRveDLB7B7ZjTRSmnrC5Q4VpNQgr
lm6vX6218SkbRFgzFQfFkRzJGCi2UI8zy504NnSsU6dUtu5Rj/l0TItg0RdB3+3z
UUoa77jegO7Mk4g1TelRZqaGxWtobGS8cnTrvhrKXFP6YBsA6BYZQFKXFsN/x+y1
tZDXKFOtr6AjcFqWxeZ/DljHR2PZVDFIfeOI+rqtAEaekO72u+39RcGukkE1exRF
pNXbcAxwkZVd1HYu2823p3ArcRHjyolVdRF4OsHZpXp7VNEHEFyb7GEe5O+D6nQ4
lVFafVG8HlZ2sf69iNKnRf3E9fp+APdfKbxtrvzJAWR6pryk/iDc3q1yzjdmRdgr
Mw9HbwXyPiJovYnq6XJjPOWH1YZtMg+x2YpFCgqvVxhp2YIKTnZdHhRFBKyPitPT
kH0UM5VpnByEASP9l9et9qsRRzJtLO/Cy2sdWJqxmI+JK8jO712/ygYTzP7zWg9T
ytfApVBRTEEeY8o5/mAWEc35i0I7uRB4zIGnYwNmiqruXu3vMqPgpatkkX7tETLL
1wibTYqFCveT5HtyBxIAGynNFG/ddzs+FjWxxSdTi8pT2mb6oJUUwOIKlvHivKPN
C30yNRwxB/7Tc8HVLFh+rsmSL9v/gyl3BZwnzPA765Fv5910+NIiCwVwaFtQqYZH
a+LXQdRRYHdGkM3KttrwI/1CnLG5ucWZkNGtbKQYABwvdRPhwKJWqp8ScInjwJP4
Sqw7rvwVry7kwrvqUS5c3vqRkSy3+rYEEses3Wan6vVyJod73wD5iyJ3d3CifxXy
DTZpVHXaC1qtbIw3epgp2Lp4pcfCUAqo+Ea4h5r4dBytGxTFDwrYA5wmc0oGyfms
RX5vtv1TCycf7pLKbmQiqZs+TF2Revdxgkn1kxjU1fGxXG7kGJrqhj6IbSyMN8dU
rBgMTlhWfKDi4mEci9AS/LagSwTAp3c+L9oV31brjZU7Pds/GSdgI1YDAWNrxN9J
R79BzVfQQlrqJUG1rP4jbJbAwKyCmFjePNi+gz9g3knExPozm1i89NFz1LgF4Jck
4lmTRF64u4EVounBsHR16gny2i0vGKQg2sTWngbipoVbI1ElxS7o9x/JxDHr1gfL
AZ3oh4QZAe6HPOqqyRQLXAOTjHJo1hX7PbSEn/PEqf/J2Uv1WIFAyKew5uwvSoJm
LBNr7pnCglDGA4Qu0iu//s5iY5afJiyEXj3fDVUmzyu4WxwJFa3qudSeG/IN524c
VNW9FYAjKjgnn86WOyFhux/MQL8qJ+REn2nac7tRZzS0xangYWHmMFx9mf+xffm+
x/iz2XyPZYeKOxK0udLOssZ5BhflouF7WPi8bApKq6d6xxPTexQw3bbw28DMdpzY
PhjqpRmDIABqQ3OIjBrlZEzI/Xiq/B33rkk9tw03fXaYtTOaTOSESNZsm0uOW6QP
tf/JQKwbBXJpqB1LoYH+Ll6bDTDj62WIKPG0cOg2O/NcSWqUme+xdyXOVLhInyWB
FJhpCz9CheIN57igQLmCFlk0TprR1CiL1hDhA2Jk8UNntexc0OwjHoXf1ri9PgCi
vtqg/MnBZeYbwtG2+jhPTrt3gDdoUtKkbYbABBymo8Grmi7Am69/Ces3pnqIwFIW
H+mSgATaf3iQnvgeqnE8sWfVx2WuON6jTY3JoqLQrUjV4H0du6R3YV64QsdM0jg5
fNJ0rAsk2hACXWRc49Vo+jto/6yjGdltU/SHWNwVjWo9PzGq1CbfrWs1GPTYYLwR
yB3SpTPjXScX6Me/obToeQtFWEai3WNS9oQ05nVbMTuSa3MSM2rN7Ni0DuyEPK5A
qHhbgHBM8tXAYZTSLyAYTjy8A0slGAU1Nv5gKZFkl974vG7XafsWH80e5nUGIkif
nOODr03MREBaeXPIr1utj51DWgCAWTXpJ2pvKr6EWjUp+UMCSeUzwrds1u2pGG9/
Z/DdFivkUoPXnt1sgYZk09sdyLXOOrJ2d1d285Mbqo6oy065fSFKhUEocXJP0uA7
hIt3fkchcyYqdq5mu4T+PDJdwz6zaIR522AUyiuAc/Hj0wIeSPEvY1g/nJldwQUw
AgmyLs/h5keBMr2ulrqFikwwBGd8UEDpbEuwz1tqxaqo3/yVvNURBATwL2nFzzVL
vdkrAfSlRd3yDMFsDafK7TuRf74LddRYrheiKihIwGn/4tKymDnrOBPwJxUslK6j
wm15AomtS/rZ1eb48ymT2tZ3fV0RqatZKTcNpCXBXFx7CKWH9mNvIbagmBwZZ3Qi
xtjTwxpkvehaFZF9eiQkZhV8Qq8TypxWlEwouMQen6I7T6HdBXwIckWcaM8OAsXZ
JSbAXTaYUFi0PV7b7PCLZoIFaupoi6IMLFvwelIZQgQcREjL1daMAKzMvLg1bhou
Q9W/ng21odHqHYgYhpW3FNK3DvzISLKmG4+BQikUGDvO64vqG/a9DGBh76ACciUd
/XTE47UAQzyqdi393hAQ6sXtSPx3WZGdhaSGB9JTIVT+F03MsqtkNA8brN94av6h
9twn1xav0sAnj55XqmKfVcOHaYvhKUXOfRZNj1SkPswBS1G8IPOdWHRK/4nBoTCP
LESRdYv5/nTFTdEAm/XkzPPm0U+hXmbfeCFhR7M8pwnhMdjO2ErRffSgeKbZEM0k
d3uT2y8tTi9JMy2qfVdZZBbJbJ7ftZXyvHOjF57Hzk742lqOezCFKZTE+XUOWO2/
r+zPGiXHCShZbMnYmbtkKY1HWSwnBocHDbfnbO9IKScRMHQB5/eYu3jvP+otl6b2
92SfRvRuDUlCl7CHp4D71THKYZENQLHTlKZdQa/PhTQBN3qx1Mh5NUEr10/XRUJk
1THLTif6iziX7KucYplbP8l/F3UTIQ3JmfJw2rz+b1mcb573HCV+eab1yljlLHok
rLqXDoLv8Qdn1FgzfNB550zalz4ysh3BmOglaewe+J4UJOO6B74h29+/6JHkeB+G
2TgO4IyxA5oenXdZUNB8K4tcrJ9Bx1enkb3gb4jIKZ1ryHXpbVQC6ZONsFi0Q3HV
vynEApWLoDLLRIHnmN1Ot/mIlJ1AXH0ZIK+aV6e2l43im//vnV3rMVP/AioeNVaC
6Q1lXUANWySkfzTRiUxw7JxIOZKBL4zDWQMXGzpJTgFFEwHW4jmFJvdp3vIUAQd+
4wILm6JXX4ePozlIotYZa9HG+P6DXVtMfKcFfZa02T+7xPRjs6tCK4vaB5T1gX9b
x0uwC2qF3HJNFeGMt9JhPlKfkzdx02fSp6LdQvn2g0tZVwdUNIsbP7R9LwoDXQaG
UeoKK6Szc6lABSWSTF9XGTxcpGGV3tsnHLel0lFPdXLOBQvCvroPNaZ49LM6ZmY+
bVTqlowpKp0K1e0QX12nj5HSuZKca+wpipf8GhxneO9grPDZou789zW01DNDyaRQ
HNqB26RigJmmYwheenuSgUS6t3Gnu7+K6186MTVpM5CaqFpct7bbytvkL8if+N35
Zi79HHMFBuSaYjglQ+CQQJtqP9pMnUeHvlTMNEorPuK8WIKUTNroCUiqvdXvQQV0
4Z+j/36W++c/uJyL9fTxIUHYmK5TCg8wg2GDD5mTBo5rn7tFcunEK+OfiudW0haJ
8smf+gmvbTYjKSWWKt+I84KB3VdkkV1ULH24Z0HCFrA9ntL0IBQzRmjb8b/4HBbQ
FnMxb8l3+c9j3Ce8uX0G9u9NacordtoprOLINTdsAIaJ94qeRtr1bMvV+LeeraHD
hvG0grLt61KvneKd3eL2EJKZ836NFaPFMg9blCVdOeH2z3jqlyD5o73igtkTAA3v
5zDCsyQIqXUIdTkMLL26alSCTr3a1/mbQ4kMqsfF2DFMQnSXDV4TU0m+dhSi3mX0
fqpB0oR41HkeO77xCwiz8yJ6EYlv3c0t5RjgGsGrMcXuTvZzRb4BaSX63tzGBXk2
lB1O+RmwJIgzgvdBKNJWJeV6NJ8cBs6/pmr9W+JO9p0dlBwC0ELIXmcJqj0eoXhy
xwQpPacTeHuJH1stG8fGz4u/o70j6hGr9x72r3IH0YQXZM9mY479ZlDrpHQ0+IUj
SxNEdXnLRP40F6dfg4qIC5jOJNyLGPRE/33N0IYzQ0shyxj44cTHSTZ9qufwl7hu
QH9MjILJHXXtlbn+Pu+DIUPm2jXPdZJRhNuH2vWBFi4/fQWx4AbvVMLYDg3Bz6L6
87dkwz2CHBlmftBlL/+DRoZjlG3YN37thK6RlAkjKYbKbzARKaU0xRFXX37g92qm
7pKiOfqo7tfThyWtMwoFfaNhyAB4agq6Z0In2pzFUtyZDn2SozyXAekZD9/S9xno
da4tlkDutWwB5F3XEBMyNpraGArKZWNJ6IQIypDjxYYWj5qJ9xcwgwDZzECZeT2i
4hrLRFatDZqAzPQNdJzplD/WFw2U2KhnBoYfszal7e0tzUJOmSzrqOuLTdrLI+2p
mMrVxQn1iXz2aT7hYeH7JtbxBAfBfWniY9SGCMtX4V5t3D1s0jfbUhohfohnjLBw
1pni1Fl4IJDj11gVI+UaRMW6ae1pQ909jPLCmjj/XZN0M+E1ajUsTNXUircbSHjw
O+dXBsGp0Z6iH0veV4FbnajoW3Q1lBHJVyE+oBzODj1hO3WSZG6nWGsho3NDJUaX
cK7xFAPKN2+Om9wwp6zrQg9HEL/pyJtCXgOHgbjWARlil+1IsPzZJd61jerL74SI
UK9WfdElKd+C6jhaVwUnZFjEFR9veoDAq+ryFeHKeOuJt97E+VfxSd2fE06WMI1+
adKhTzd6Jsss/QftYnNXW2+tYaXeCJ0LwsJbg8VjeZnhaYTWvgfFeQcwyYykwi+J
sDJxju5DLXf9NpMdRVrt56zLvc2Bch7xXO/6JkXF5jD79shNQhJUQH04JuIvMXwj
701vLKyBzMNU/aUZxujS7demysikaJ/RshJd0l54+mTcfputGuNnAcPhHFhDNT4n
pV7qWbzydVVUo2/YW4ACnYfad/HCtReqZu+AmTAIYKeuY9dsAaVJ869R7ZQREAuk
7gTB10kqDcJORu8MK8vKfB9qP8YQtCrHQiHd26jTK24RS5mbe3ldGiLOkLEODoHv
v0C1X7g2LpGRSDbEC1yzGHJu515Cwc+GaICZlZ/stb4iqeWz1WdjL4pnAiOWGr+n
4cDWrqTID0EFeQ81BnVB1AQke+/PPrs3lOlW3+FBXUwGGOmd/PiG5haGdsKFDDa6
soEf8jTCr7vHM03Pom5RuJy+JL+v3+NiCMtkq29W2FtshfRDOZFqC8jlzOgPeuT6
wyiucO/G3FFqECMstBDaz0KdNRIkMg5LcqRg5UI2had/invM5Z8CKpaQw8DU9r6h
2fKTTXXqUUf09pKoextiGqFBG+c5g927uVUQvmPgLRuAPnibsmMMTKRsymCOuriF
b9C2j4cZU7lqVU/7sxRftaEevXuiRdNcDu5iwfFaoTbtyoOJXpkyUtdMsTp3rQWM
DDDQf2smXJz8BG+En9JEZU2pLkWAynFPrJu/qp2RkSqWgeBCt8o5Jhjz9RjJI6+k
5tpurL9w9c/Cgkwlu045ATYftBjrTY6q+kYMW7JlEkz7fs/38JkabmmABCLyPHoL
l7a1kNq/02YVVhD0XvvfHPlOYQoEt6Y5tIzHCumbcFGVWJDsfohHQcdbXTSEaDXJ
qcZku45Bocnrxt1y2Soy31VQe/DpdihSFYAkQ/4cByNYqj/OfnBGXakSH5NRNHWa
9PzOzJrNGSl0dsVy1iLDmjYaXIjrvm7drgdqpBrJC/s24UwVvKjH4+WlJAs4PilU
/V8hzi2k6eUrUK6eAd7kKzzYB9N4Lq5e8sQZcYHz4sB6vJdgvCiNb1qjO/Z3701M
uWq8+spzmF4OSG9nMebz/k6TaSub3YzV8ZDXoFmcx6jw2D0yskLec5dHjlmYi1fg
C3BnzQY/oH7DCJhuVZgaVI0NRtax1z0btWnT6hnKv817tIcmXgE2aZfz/A1cDVbY
P/IHisGlpnAsCmGOcRQ9EOOFbn2mgFsfp5WiJcsGUdaVZFulYcBKyuOVvnJOBK/I
bFjNweDeDCSVQZKQzpeNMU/+UpMVDrvETqpPsOd+3geQgxLKrRRpkCTmUJ+9wRl6
UYs3pE2LHKAQKiUgcmzw89V9Nee/YBNP5nYQxeL/0HFNpBfA81EC445oCQ7M8voy
a69zyLU9axflgeLoHFrtme34lHLsYSkvo7CzgOUA+q+P9CiMcBaIhyN6VlhDclIx
oXQPS8sHP74vJG/N7+x7EWhyxLH9buA6W7XtWdZTUJCzI8WTYy8sizChkOs3C/tT
a4qv9wnw3/UgS/rTGb8xGYz57P1pvCQSR9sETGJj4wJiJVm7Xucro7c4qV8Zyt0g
QtLDLsandQE1znHp0t9WDgtcSHE4zEhT7HQISp8dxY0M/CQcbEWEm+xzrFcA2Bdt
rhkikDzJGE1Pa1d/Y6oMGGjZzsL1H8YV/3+XoXxaTP3ft06WEgxRpu+kNmyBkzj4
fgSKw1DifBK7BnEpvgN5T31h3wmQJVBvaQcztc/K7gcBqpum2yOywITd/cmkjx6K
1d33ySe7ZQnaJVIYHtA27LC8XTBj/yRcZ2c48iCTyJnnuLKbIWANlNocc8/XAqXI
kl2dlHIWo59C8d24z8mKNTZ3PYLo6Yst/i4P/NQheJww8pR/tv6J+a7CooHZSNDF
C7L6CdQaTv4QTq8ih5LbRlwAZ5bzv9BH4Pq9zpcdf1ECLZtiRga3PA8urdzDW41q
xEEzr8hR80GfiBIIYisoEm3sFc6vdyszgfTqM1tTZhFMVsUcpZMDOGkfT6IDcuuf
chVB21j1t3XkGdEB2SqebLWVLaDXIW+wUCItCa7BRs3eFU4FmpBopSvC4ZCHSR/V
LtxF8LbhdXyOAmafKm8ZpQdVsw5OEROJwkyHxW8dAP5JFYQGEJ97Xw33kqUWK8LQ
HWkulhZZ1F3f+UZgTefWXJ+n6a/tVcogPMwG/ZayDdzXH5AUC9+U4VEKV5hP7dmb
7es9EaWTLadKyh9UdkKbNnDFZQr5H0C3oRNtGZaD+SuX4aPEcCiQvLw694TGkVKi
Re2kw7EXIOjym5TaFK2oUC9/LJddIyDFFV/Jts7sfGFGEzJWzo6vOfs3sz2KHydg
mF/r4cocQadidu8kxbBmDR6vtY71yt2hNbcaQs89F8Pjc9gHi6KaQJhn53zV9Qft
4Z6/+P13WDUofHuDdlfFyM0YqANuyXXNZhVG7C36BnM/S+DUQyh4LHJIZ3ZQtMjE
Vc7w8Dqo9FyhJqTPRGAG3iQjSixHQeTLzUHoicWh4PpRIwwe6n5y2LQ4D+jDqpM+
yauC4Lf20M9iSjCbWFpdc4KfPrb38IFURX8ky8VB8AksDC8c/qjgDF2qU70i4oJY
EUvUp8fXN5DNo4H9zgj5o0ZXWOZkkkkrOIbVYa3BpGpeW+Ea/FZskneM3PBca+CK
ZFVY5r3ewZ9Tt06GC41Ynfjh+qbRypJr2mwsFNlCRaOvdXAtUjBe1jI+DUxunNC/
wzFfoQjzs1o7h4LS3MRHFxib7kjYKO+q1z4QsYG+Qg2nT70WSgtUmVgFrNw3u/pk
gEZdaV/wupa0ZyB90OuF1GSHoUqITlv2qGQR/hx/A342K2hEg17IJ2Yiova8dRS7
RxLOfrQEw2CzOR5WUFiHBmNtFBFSdDGYnuRc6v5TYfZOpCvGsVl8xhH2BXFmPfcv
mtKS7vr6PxuRaZ34gg6rlv4vGOrukm021ED0V1JfPoabZs5wmCOFpyZnuDcJDqjz
zhAW/4GY5tUY3oECwuZS2WurLDCE7YHs/rHRRHOQhOCi16juppefnv8Hegah2eXk
VVCaBvjRc9pjhJfjZeiOhsf7jlkqfcU6LZCSqeA25B9+nwAhNdKxWrU+b8a4sw9f
uuM+Kqbp4oJQBw1CGQR/mkWeQVgVU1qXTCfVaxQZomuhUExWXcEXWu2FHzvxOVXe
sVJFxqN8o1cDsN0+9LgTc5YBWPH1xQekHipeln1pzIQl4l5J9/bBgoZGng/C+WHf
IgHGRsllHfFXu/78MJb2ou/JHcM4ZYZZ4Webp29KP4eGM83H/TthzABgJGcRfJMf
AyZPVsxs8wXM5qoGdpOeOkJhdL5ushX1UF9j3JQaM8Eghif16l/VAm8nfVfH9APp
XcwxxsULKhsuaYi5gSCh18wfTTHp8xRU6nC7PqXuWRiYoWUxVeOZpdvpfrt3/EVf
63PQjo5gJBkUvzqt0dyWrj1SpHe7sT3hycED2Y6tgA770qjsypufNGU3FS0+gWQn
0FvZw/QNVJRwWVyzVlBRe7xSFRF0v9t60RH6tG1CZgbecKY3P//9ccIMKhjbUgBi
WWTULCLnjikMpznu2Q+dWs403b9ae1jo2u5x8fuOQ5fdIIHfBobSaXS3OswZhBo9
vc/VgxrnuCC/xvV7+AnALUdunV9e5QqV/Wn37ElutdrOkuns94JrPSZ4kE+bmTsY
8PiUWegBg6mygzcIyT3CZsJmz+WPS68O6JXZBbxzgqcSg374rl9FRsVrL//8bGfO
GZ4Q0+RB7bsenx3mbyJza1M1HgaP5OxEnSWswdqQ+yRHJ0RLZF97GpwXIWyOXGCX
6lNK/ZL6dA4Hh+Ua8vaCjAiVpBk2dXMiT68HNhrc3GIq0x1camDw4qX44wW1FvGB
BNAvC7jSw5Du/wirATwNwVs0MaTWYE5Z9jtF1hDL61ofnKhJILa4FflOYztm+Qz+
eF/efjelZQi++cRoCPpyrJ8tRFHK7KUi2Jy+ykV4/t0dI67xjsQqHmJNWijeHshS
bDHfFrbNNr2lQzVC1i1h0NGE124mYDd5rrjXkLmPnIBjF/n/SEDBeN1Ggudjo8hK
Wyy/4/uyxFfXxoGXjEiiZMiRRulC+EsbxkS1Rc6E9sgF34cWvPmXk2ARltPGLrAr
wt0slVPQ68uaaX42tbvsMdTlkJIzq40d4lgAHIXBZDJmfYHPydHVjqXrgFTDmgQV
bkNgXnwDtYvTHIqACQMlJpZ2nRAK3sn1Bi/mlWlQBjz8MboLc3R3O12QeVWYeZCA
TCi3xfe3Ia6lOGfxCTdu3BncMme9eqiOiLPNa8OhCtJbA1R6vA6acQ9d4UMQZL6r
RdPO20l2RXBTcSXLl2mcCJnh989DtWlN9YDXtcTR+iAo0IwYeCHVY5ktxXVndbUB
wMoztFUcfnMXI6WoSzEo6ZVU+pD/up0pgeaRt3vteDE/GzHs0cg2wU9lFRJ3sE1r
aCqFAZzO2Srh3Y+CJVWaucFH0CiC81qyWmzLB+QplabTdnh+Jcduhk3gfICPH/uR
UtSjYX9xAjE9f82owWfxtv3YtpiUpypgsp7cj93GYYidz/KX+aOU1DEoP1mXbhTY
oD62jIc4Ml/TZVI9JIrWzRvgr3eW/FPn0T6yYxE492K3GnuGddaY4tBORc9nikb1
QrSn8tkPvQMbts5Y5bSm//rRNjbt39ThcGY3j1EpKQSi/Cf7fhgHgIeCfa9nM7Fp
gmukpFOdVdtybpO+fVgyidE0JuoUtf48P0WInf+Fdf0mMS2E5h+Nff6VJGPoK0Bn
c/wHCpnCTkxlrMm1J4b8JZhB+hwsJhLlMM95DIw/MBRTD6BtFInsol61fAzQcmzf
baOvoG6M3muKgcxJxWGJT6tNx3pSKyzWML0oPd16oO3FSC53tqyuRcXSxi8kq8iw
nZxbLeuuZvukdthZzAgyOU2xVeSrLHwAqIVY6RWJJ/xibr5dFur1psWy6+jmYZta
VxsndHe61NC5OPIjKq7tnpQbSHvjkXGxK6/2+nfvYiVcwOe0YMg5Gi/cci3tkGKn
79cTh/4bh7lHP4Vs3l1npWu4Jj6sDktZHRvBrD1rsV694EAXxAGTMOvz7XShm6OH
VsjwkBPaMR1iFh/x/vNdF9b93vNRCrAQ7AZyki6nakagrHFWo93WNyXYAz2AM6hs
jtJMz0K5S4ircrUOW6U60316lKSIcTyelURUqY76HEKsmh5K/Mj0Oa8/xrhlFZr8
CzaHUm5uKsjdj/BbNAaMR33GVA0nD/+YfVgN6A04D98JGAqgCugfsvw9KmKc1a4z
V+4HYmwv8/xjM5fGqHkqRDl88K0aPgBOVwLsjJ7Pb9ex8Qxkk8fpFbJCCvcVY2D1
2embNIUadinhndpv5SHei9G3Dlp5H3klkC/ZS4/N7W5oi3rcVPAVuWBvGoOCjZwm
s1ikxS8BhtQfnujcLKuK6NxPnh/PcNkOw7VxhAaob94ruHJkNIgfzouTiNvHci9/
5XTZaIgkNiqyQrIOlDXpURAoRnsODqcDVFgmZPNZZw6cw9DM/ehpRtGwUIPubKdZ
lpIl0OFbJmikQTxUbdX7SqQK+Y6NAUSU5n2f6uegNMST5X2HZM/Ep5ij3RzhHRuj
2jswdFI3X9G6153ws3n36CmnCXJlj0CWqJ1BgCpfbgZM4UI5vOf1Y4e5cy9iOnN3
3dauImgQ4qLNKkZ1Basy3CVLMSpa6sfFfb43xLdWvr5w+pFN9P3Jzwjy+IGtqoyn
kUW3G9INyfsMrZwX+FUh3D3l1QllbguNK8DJQnC0E18y+45W2z60WCmwz0xz026Q
+haIkR4s7zI82MamF8S022GViIem4uwsD5bVcHwrN++mPmsRd/zzL4elWxUI0qNL
/tgcWQz8GnjFhmNSdsixjUvRS84TQOJN6Dj5uqfIJfqjCMj5bETmNwqnpVaxBauN
Opt5kAyuCCnOJxp6dpLdebVweLmJ+KFVblaKj6x0zPAoMXaQt1gEOI5zUraBol26
Pc8e1oLbICssQj/DjRlTOkpXbzDOHGOFIdlw1qBdRw0nV6N2tk/Zg+SXB/W7lrMW
SkzkliqdCaxGK1DIbQnpLESeCa5m2So3QBQ2vAtMImFeUMkWLMQGACO1IT80eEK5
tFpxN3qLjQlfEWB7zbI3WOGh4KLmV9iTHs2jFIgapchsJk1to42EH1vFisf5Fnxt
WLKdqhNf06y1spTaQNnLZLamZ9L0iaxd1cYUjCBF6nb1jIhmiQkIAjRUMZsKC3Xk
IiyWlUEeBn8apClKhqy8NF6dMuxvAUiH50fKVDj/APcwNMD1l2p3detx+XFzkX4X
6qMmNcxkdlXuBEyWCIKmHfJBP0ouE4/yuUtHzwPyokexXK6xTSgyUPFVPYm/2+ll
uvtoz9tm8P2kYTa5B5kBvoVEJx0Gt7U+yT3rY+BrxE3Bs3L96QMOZI0N6t7HlZd+
a4VqpDvIA+8FB8SecCjAAwErH+ujnqxB23xGJmLT4pqTXVZ2p2JxlhyzHVvGmTrJ
icdyAbOu+UnNpzMl5yFIhIKyldWBPvftJMSAnHmmNVUdpEmwhI6fqa/ECiOM5eOS
fqMfE5cpUQxd7ZLKYMypINhM8w+lTb+hxOsmsIVOFvMZntRh9RDmc0v04pXF3gmf
GWMeOS8VZD91qMUyJEYDMJXJVvXEWFcI0tiuJRc4b4vQcIeAnamkqH2EYZoPpyeh
/JnM+0XhNZA4TnEXS5wWc2dPNwdvkEUxT2fKeBtovpuJBaXDwV56XolBL3lZlH92
71aju0eiCBfFY6sFFOeG9AZqWwSvNk70t5a3yOwoqW0F3ZYOOs0wmFm8W4TF9d6Y
FpHmGFhZCxY4hrqR8CC7naA/kcif7lFhPNnUUR9GPbLfjlqZfsrhXzdhJm/P4qGR
E/udjtRUyxiHoWcGwSmMdv5dpaUgCpkT/dBXWrsyoyi+Q8qErQfitZqPbJQx0WFx
nLypUC2ajECsvM9/JVpzLOAU3W53Nk0gHK+p4tfqUVC8Vvfky2mqpw55wVkstaic
GiI0UDgUtg+YRplIzZhOFJTc91MH2MTU+AT/eoh9tcboM2JgiCd/Qj4b6IUyUkB5
MMCWgn+Q0Sthp7DQCIcfc2tXOm4LM9AY4ossFga2QeRmTYgP7nE70jZrSRPPOmyf
xLhZPvzuUMsNIa8Ttv31o8dEFXDqDGDzC2BJPvfpD6BTmbk3BQOGT56d2gI/C2x+
fExa8yFPvA/fY4Lszz9GyuMmn7vRtt1PX5Kb4Aizq8/QsAUmqkd6H071MnMqe6uE
EIC4WpmTR9qSoxVt6wRWi9c2Mer8sq7bhVtmdsinIgXQDH2M6MVyQbB1U9Nsunbo
MiWOb6WxoXXP2TyKG/rhHgrPzcLFZJZ3iCeeXgknyNdQHr+mnLuqHx//vz0056Z9
X+okuslAKrfswbnjoa+51fB1XzY1BuOYzy5AyRWz5fXvDWUnlbVyFnVheTbDfFt9
MNcFJq2RtgjdJjeI6i7Rv/2E1ML2J9JUKS07Gv8xeT/35WWYuYsl1++fZ1/A0g0R
I+jImzvTrsj5qvF6s3vH/As4tjH8/yaMCT3BK5PsW/A+BMZ++XV5Cx/kJVsWrVIp
DPkzPp7DjDUBdUMIUtHtwil4WjXqfxFG0J7qw1TlFFAC4LnfRGRUqU6Vn+e4jFwg
Rfb9JQED/69rewVazoNl4QSzuw6yHAykap/HH9zi2Z3ddgPrjXHhu/aosXnnT0+E
2+Z4lsuAC3jcaPBArC/tsf5QxfqFtBsOljNUeIK+FHrO9h0d65Ah025s86y+FKNG
hYc883BBqomhdKLQGibG4bJf6OvvDY8TXtQyoL+8MGDeq5U1zUXBc4+jAqqedJnO
KYVqwCrSLBzZdTCihrJG3eojzm2zwmqvdb/8G5HsngZFcYQbh1E/Ard5sNbtxtfI
S4d2Is9oempeEd7/L4rikItPYEJ3CO56EScPHzEE52GXDGIsRUtAYKRmhxOmntyI
vZlWcD9LNgUkDoI8fuOwzRX49MGbrXByLmso/xn0MW22YwaJviyDbeKML1iRSsqw
Fo4aYyQnWaq4eHa7hCb1X8xrhmfoaXvpUUtT19Umv5mq9c/OG2gUSUhKZNdFmBGo
8qH5KueBTsifQEQFd90XPga4i9pOKLJFd1hCQj0n5JUgKP+QYUNIsyZ6Ip+qzFXw
E+HeFFs3+pPL/sGUMgfSEnW/SjFOovB6ic/VDl7NgctuQ5pmZNEMSZ8RflESZf+O
ULcbrJgTF5Yfldf90AB/XqIhYKQZzBKwcjt/Jd2TgfAQ5KowR8zveSXVjVoV1xhX
rDeHi1siBFK0QKvfg5aZoqFPsKyX6IcDMzPSWYdapaa4XXSz3PHdjA/LMI5G18ZR
1vuzemrjEYSbO6uq8PljhtI5JkDqt4P+NE0wYA7LMZwXbc3yF7WdwHdRTcIOI8Un
pG/ttIKvWRwn3qFHtPnDp83Yfp/PDdJ9ZfpEjfJd9HFzj+NqyHEPG0aKJpiDe3IC
gk5dTNqzyNQVLr2S4tyLe9UAVQKuX+Ra4WJDUonB7TqADLcPLzGsSV6p7nEGG5uH
UX5I57hrjXiy3rvF0ByOPlwMR5+Z6Zyfn4r4LmUX7vM8oN+Qj9BxfbqY2SjxhDGv
Lxx2nkTe1gevCMdPnJvl2LlAsoQtylu10RXqbL4pVra5ET9aSTRdx6HJeB2/6xj8
dFSlDSDCt7N9h0K+j2P5XVDCbHMN9n+JxlZ1l1wQqF4LDuTV6xql/7jjrJW8s7Jk
UFWP5/Qd7C8ToI9YSeLlZOathh3nAjlLZ0R8pZJbwmUAzHnDjUtb7A1UhM+ow30M
Y6WDs+pvmTWZ6XDcyv+H0oWWcYRHS7Kl5gRF2s73vlAOemwrQZ1vbWOimj9m/blP
slxT6InSiTQfS1Lwk2ApU5HV76REPlZYmSvRW2SGcB5hzHuk9n6DyfgcNFzal00f
3JaJcqNGggVzxOTVwrafQ3mF9LS1KesXWQ+SZnKsOAHzUYAJ3GNaAJvlQLVo0uVP
/zkDLePGpdcxqTUiFw8bGpCo1tGugxjOJSi/S7THQpBhUVeNh3fbzbM8DQTDCT64
dq525gPv51PE27Lm1KQ3XQLZ/sgfCTL9eFueLgLIY2PxBBL5NS74zVUC8zsOp7ei
jNi6+WHhS6m1Aa05ZkGW5VXMdveipyXqy6KkwBgNdHkzzmJZtp26I7dwFuDepSp6
md34OvtpJYQYe42DRnZW3GG3ZOjnEYV6GcOxJN3d7ywJZWCh+4uZzW7R41FGlM6b
qafMaZQTCMTkmLcMtczkabyw9hvR+1F1yEzvIGSTAz5b7vzCYxhtqmxGMLZA3PHy
X33fNcs4yb7mJE9LzDdJgO3zZadkkURE5bKgL2/9qFgO94M1iVYFjBsirmIoVZ+v
99a47SR9C37YDv4OUAcO4vjOhcpvBbiksr9QByFnz5jTKlzb56Mt1vrw2lrZTvo8
leblY0dT7jPGhjhAIBARyHgT9sklLIav0154XAtyDj7tpaBsEaVIVNnyix4qbJHN
zwzn/uuUQqWMPgBJwEuyPmbrILYtpQtLx73BW8U9GGmz7vGYLEPPwHQRri5biJEp
xkqCNkSfshVu7qzcZYCaMeVMwVAqsBG/DwxEbW4cYHO+ezUxAzkvMOoLrWuXjYcJ
wHdONf5FpW+nSJ/Cmv6HdLiwSxlY9+IqF9q23qluzHdseLZ5V3Zz7wTJRH9ZvvRC
5pXAo/ZlvBK7kyNFJ60gx8iQM7ptcazxmqgUmKALoH5F168EyAR920yPnMPufSjJ
qZtd8aOl78Aa+t2gXttilE0hRYKO3XfFCE8fb5rU5mfo96HzJ8ZFP2GfnkOCKseO
vMrrE6y5ilQVKlKlYg2PMdxAbkIReCWdlUz5E+P98QQHLaNoqPRafJqEpcqm9tDV
jjyHIX35LW2jwfLtfbt2FVeMgScl8+QxsgMy1k2YPck9AMH1Q5KEYsvFB0NgQ8JU
ROoIUzLRZHIMqkHC6aCFQXVy0dM/xQJxGjsAfhnMEKeBTQ8WQgdF3P4Zz8TEA0fL
HL88tKt680KWF86Ss2477DNbYGYQt1thJ7O0AN3t9sNdNHejDkrlTz716hFcWazB
+y25jqVxtwUToWegkb24Hu3fCI/njxsoykAgV3Xj2wSomGvFEvBE45BDOX3WJpGu
YiOJRX200X+3nYLMdLOpieflzSDkn0OPRqdVxYABQuzl9+aTEwCUA9MnGbGPDlz8
tZ5++prxgTnQuII8yi+ZCabs6ehzoDV0ZmMMmZzV4oVbQtI/7990pFdzCX/7j4p3
8RzKSvQQfarFn2Wv4Z1sOUXokHbk+C4wv65y35LBFkpiZP2A89QVFkypRsD5ptBH
x+kDPyhnyh1rIJ82eUnN7RxYRDNF5uagHrHoJ04vC2QdQHsawbtv7PQTARQZBDvL
Xub17pHmxf5zFM2ZC5hvLXL6tETS/XF4VpcrqcNzJaziPuIiG1emQIxo3UsUYxrr
FVgRCZhVXGSUP47MlQzhK4A6bxA3Ih98R47ad/M0xYZZt5Kg7oG1DZh0s1kqkrC+
U7ncciJnDj35xu009j4de2rDD8yqZBktIDYG2IYstHmfxlY1GsRf+UQmpudDOddC
1tm0wmXYQXqqMpq/4d35k57/QyF60XPdstCoh4zNXzfKHfUUiqnk+vZu+sSuHc6U
1PXAwPhBbZpXuuPNPe4gLKu80b8qtSjm5edJDBMFW4STKfNxeGoY2siPbtSlT0JX
4aX+NIag4P3WArVR070oNoGHc6msMIEJlD9AVYSCsvfLmGKPm1WkkP060pJzrVPl
d/MPGBaT0CYMWVIDEwfx7kRZwt5J0pLDXVuXHyK1pFyccYddutM0oQBI8R9P3uap
acHZyF+RUphejJspPsRuzUh81Ab9IxRco13JAFxH5T01OtlBF9xrdLPjygTeX/8Y
nHrdnlqQbVWpGRUOd6QgTF9WCFPmVtn0jSp8T/FDCzRyZD54cOOTj2aYcYeyQaH9
qQwOkTaQbAhjVwNLsrdrwJ8VU+UfJ5ftjpBkc4J4gFQAIWf4Gz/phcKayHzXdCdX
T6MK1/VCIXmHRByAVRPm0vc0n8EgP6a4Qf6QUN/n5DHUxNsgOrl2WxiTFNLhoOil
0wvTFCI2+9qpJd/LEm4CHg6gJwAG5PWGA8k0QIsEtjp4YPsGFnmZH1PU3AF3MH2n
wy97erXxbF5B4mq1mRQELPxw0zTXrdNJv2Nkt6eQbIpke4Kgo1xkZoWTooOkCNmo
o+CzX8lJTzC18BL2PVlK3xm7c+Glw4eJjqwc+T44Lbe6rzRMBwAgovKQ8XkfYbTo
E2ufLukTwmCEouR8FqFC42MD7knWinkVjZT1WF8qOIuWZolN7uI6tBT0/YE4WCwc
l50V+cjhPhQzmXjISL11UgJwssbfGMeU+uspiE3de6WJebs3Ll1ItWeI6JxL9doe
GpuDaMBqV85gCxLLRGcij8vlAI5DXHpmQnKOi1qZvQY8/YUGI7eXYRP2KKibIOST
ksZrprDHxiKvisPtcZQk/EZcJC7HmBfVGQZxld1huX6/tSVsguy1a3Kv6Q8rmlgP
IivuXErYejo5yndehId4FiZDjCplnka57oryYHKhqkocO4+ZIfgNb3R9TGW1nIjw
LdsKnEmfNifPjSohXlAhwO6mUAlJ9DN8GV2uvbMWUtPll2oK9nldWKvRJY+v3JMK
eHX8Wh4ielMIcrukUmosLP1DPO4Cq0eP+dOFfabu9LXrbqNdRT8nJcMvUw9duuda
eINPKbQFpoxJm7PcmZgNd9kfrjHDQHvyKLAa2Gf5VAsJlh3FDFHvHNromR3XE1N0
MIaConjfvLGK7558p4RnoibLgQe5+gkcmisdRGVWvASeBc73AE6BL2E8JS7dz57x
IoUVmHiHelogNfZNleSrYAePvWoMs5moxuWttULPEp/spatrqLl1Rr1ozDPAvuMH
HyrGDSXgHElAv1O1/PaXvHJ6kkABuNYPw2xARZ59GXZOiA1e+83Q4tMaPzOF+IEZ
oIkD3XhIKPmmLKQEH3ooGC3JPqPqTwaUUpKU5glWXeS+ALB4SWvPEhMdd5+7mwZT
sY3kE4y2LvrZCnkCf1Tg1Gq717aoF/B3Sxg9xWmdgZJKXElKuYcTvMVltTQ+WNSq
ddB9jSk3p7nXKK8Z4bqQ3ai3oeg+UMFv9zwATNPyqipv5F/A6N2heF1JZ9ut+68a
jntzo7FYIWuLLqCZIkcNJhBrtgF4dZvMC7H0wU8YAYb7WR1T27vGOvj2zfUKpio5
JV6K1bgDGwuk9uJsUbX6t+1VEJUmGH8cLFmg/u6nixKgPR+v6+lIUHN87s/FLU21
im74DvbU4QrvBVrLBGaakSp+88y1arcJV4fro3hh8x2AMHCnEETHZTW2Kb+rVvOq
fEKIOmwt2KLD+V4MfgF2yQA/cODOIbEztNh9483PwhH5sybyqej3ORdeL4XuF3Jm
3XGGZx79krGDxNcGpzmUQvFgFeSndZwsidJWUMrzAfAADu9Zpbh2LLxpELMOntjC
oDYWeV1d8j6V+8LVFmn1kMKrWjuWvquvWEsPgepTmU24/Dsy2vDqXqYhayscHRHq
6jXcOwOPQamIvlwU2puRXRTZLdW6g+yyOngvFUtdtKWc59cGe4kLRTg5uNMwejUD
lGxjK6R3O21u38Z6jsyAcMajBrO+VZjGVmxAUSRAw/ATrr3Byd6Wpou1KoYD/juX
whSkUAuea9w6BzIqb6U1VsJ4XO96rPNhJS/7jRhlPM4JpqFU3zKpw57mrejBVsU7
C6rLqXKbKlXQ0zN+SQ9T/hJJ5TnbG7P9qPHuSZcjL94Fcfnd7T3SlHnNcYkgPVTR
VZAZUz7zfceCJTyH+cJyqLiPI6UWUCMGhljAtNdRsCPb9bTGFfcJZH2OLkI9/T1O
qSu8APQvDouUIJlmoGZsxLj6DOrjZLlCwuYm8iVzhZ58QOrKudGDT9fPU/YN55Se
+SE29JA2iOvtK41dP0wpTcaH7Z8ZlfEmUjAoUNw7qsqy+FtWBKE9DzFkAXalAnYe
SM620WbxCZbhRLI9nzu4bd9qpN/Y0tPSbLZpWEKDBPfn8+NF94+ZRF6dHXjajmBI
3DLY1m1u9xfUHv3NWLZDCJkVkokrAnK5e0jwvmtDBDQkY3LrgrVA4wTqgpIWVuYS
iiVsg4zuuoE+PN9KmHD8m+6NanIxyy7MevdWLOuIqAZyHtQXQS6Fd6M0wmo/X/Qn
P0qquQcsWGfBpgEx0PhbEDF1nX+n2ow6+RabJBDPqtyZKrpL0mY61NbJY7Nwla++
PYVC+KYBUAtKAgYnX4A5AlTXzDtFmw64/Xce0GEXYL48GZ8G8AM/P6rkWcEVHbCR
/MuwIDPs/GiUVEz4rDEaYOGhWIY02/zgEaSLxOLY2jhqfUwW8ObEAdmmHo5qiKlT
1llMcvPZXU9l8CGKZbkmrU8CUWEXwpRIrVnUhcTdoa1C06jyJGI36WilcGeWKMz8
MPd2ZA9mDo6UbjzNPi6Ly0zyZ0FqVJiUPngWBIyB3RcNTjIBclvnpq7ovE5ydO8i
ciHwhLj2u+nvBrD7hLbSpGtW+CX/jYLJHR8Pr1KOk6En3R5D5VbRDbeFY44lMdiA
p+Q4ZwE7BiAJWlAoDcSpbr8KcTz1U2x/tE6sFYskN2piZEF1UsbuBnr89QqhUAbn
4hUIHbZUXvgzbZP0G9/DSX10uNKaRmz4HhaThMgA0ZJZgcVWt0tt4Pl5vVAr5qm6
YOxWOpxBwv6lC7cNOFlJjc8+r5rILgcm5K70Zb1cD5AVMQndKEqwVhC97Xfip+Qf
bd410vJ989XPPR8aU22lTvVsICy+cth+6e1+oYp0KgqUBPSzJA7WfYEgS5L8Pz40
S+dlVjm+haZ1L/LEqrWWLTGS9ugkEdD5L1YbmjT+AxGRAHkaZaGnkOd7vRrhp5tC
HRuUAFmBMYv5yXulMvFiRCGR3/qIhg31ZLhoFKLI+4UhDEKRBDS/ftGzkp5KS7Mk
3RTpmjkfzCq0v++2HKoqkPax3aw1WtDR+yu6ZPZMjMRAz0DBTZmTwxk077bTx+S7
JMnvOKdydu0Gz2GaI7Qynns0EAy6gR9VgfLDovLJ4FX+U9L4PjlRf10lZVGB3xBH
ZjjQu6KIngm7krhPx4+VBez4XPfP7iwVkiz4CK4tFCAhpIDsFNGo1d0TJLUJgFOd
96ukcIVA8/Lv1gz9lEF63LKhO2gwltb6DyPNCEy2TTPn1hK4pc4fynj+oz+ahE5P
6SQyqkV+r3KAl4/uanOq36Ra47uM6XJtkWv8nErFLMW8Oov1UbKwAC8ppZ/hJzCZ
/eufge8r27IRRkpCn3GCxIEUUkTCF9mir7UVtk385RHTqF1mc8btbasL8jffvkKH
axNHQQhoTiyXLy1ZdKV0pbnZADdXgxFOas4HNuPpE3NI4K9vpL62dI6lUu0LDp+S
HqdHRpQuzsqzwBn7l3GJD1DUaCESUhtgzHqrXFa9gKbNL8WMR5P2YVTHBpgt12Xg
OIo1QKmm+Eeqe5Cm+i/nVpT8RKScS/irp/tR7kpnjQ6N+oJ5Qqi7RAlBEfbZAErm
N1cldDs+uG5h2YoYIQleRdjCc5kPNEn7kppaTlT0QgiWtymVJS5tMs/3ZOk6Xzyr
C7guoaBDDvQX0XWNglG/Ccrv1xy5IonGzmFOdZTeysbjdySU0nAxUd9zOFKwnN+i
7ooBS0Rh/vg2ujyc2aNFVvG9WHjJR1Q5XL2iy2qbsoO+Ul35KgU4VsxqvfGTZBie
MM8v2YmTd2378ZuYjjHoWX4LF+aIuNhQ0cymMoyoqkf1MhMpJo2Ds6rrVZyYjpQm
ngB3wrdSTEXArtsO/llJtQNP1QEd6u2e5SWJHgIZ+aGfWSQKYKY46k4EWG6Cijia
2eDZd5qKczERwrse5smdWeAIGI+CuCw6L38w6h1/s8DoU8cXneIKrpyP5Os1tvwJ
ZJQoSH80tAjbX4Fn6YZi0fRGgH3GuUuC9zowyL3TbU31ooj6yYWCFWlgo0tON+WU
XIdeYFfZ3txkBRhitFJF5hHvfmSAtg5EPLD+6alfLOp7p6s6dRlX8ELfVLEyluhb
KEQjFCrg7GgAAj/AgfL1RW7n6ld5Kk7oviQ12gbNXZ/N+j5KaT4S1bXmLGtD8Y2H
KKhaJbcCwDzlLecHYBboN4swb2qmkiR4VyFQ4HiTQGVNBtpxi+Wc9ProAsEnHlhi
NudXC1fePB8T5UXXylMJYG0caVOrxthgj7EhlmuisCNfOvSmNYuU89wZrb/VWFa9
cyhzF3mKVlY1WyZnm2ESForOyGNcTCTY6A8ObefYRiLP5Rxdhu5s4WzysTKSbG6s
18Z/R3n5dgoLEOFO6CtKhRG1RMAhZ5S7RAQTnqMV+/xTOUtZKbvflECwhO/UGaMi
KyZOJm/HDtuPjyDFHMQm0s02rhitRQcingJoIUp0QmPrqjGiYpWIkV/T1QFfoOCS
yjrdY/vT86ENV6/0YiUXXWi9ZQBVsD1Z1LFOTplgTz0SsjSnQ9C8nOix/68Yd18R
Lx8cUEvh7ax/HzXFfIigWWYpwwquY3Pg3aaJap/ymQZyUHnro+bsQ1mqD8RTKi5J
82OK8HObOutd1qdGyEH+bv3CvVF2BHvMkctdFTxpwgcnszN6AKESqLB2Td6AZq35
vWlHQo8cGjHNSpis43TxHsFcFkQ60gHMwPOUcZYGvra2PCFXZykM5DJ9daL5f3IN
5vjJ8WP3l2app8Agk4Ys1OFZEtPjm82VFp8I1HdkIw8/QF41XGBfSzfoYZw7RYFx
KyOgXLlooIOU+5fKHzkIPAu2Qny30M1Pts2qSDJNNEYh3bDkPROpBpSXenOnKnAh
3PD3ncGhS2UwVSgoIDQ9zJA4MCgsO72hCJARKfrJJQvSn3xqHt8/f/BUjOfQe3EU
SgyHdr7WoAR8NW+GRLNIsdkqN5FeaK2JhKuHC0uzpyIEByP2jGrsB5WZOTpQF2Tq
LExiXJ82+/7lJIE3/v7rAV3h75K+5ln91XuJdzZUa9o19n/wZYPOSI+Q6f69O9RU
T+MuKt7HXqAKyypzI+Ic/suSBaVlSJ/mwIQL717lbSo2i663jss5fttGZtoKKzu3
G2htFTmHxQfjnP0geg7wuP/Hmh++q5yhsVIdiKRhBZQFIYK4fw3qhCuEnYa/Crjr
ZdgcahV/14Sfsbo09ewpz3fmiS+DlUiNA8UyaLU8tIMXqLAtOS90li8XQuu4/6Fe
BkTy/FmxVpyhoBOp9XFFCe01QBGzQHKAZ0BaTFKWLJL6eUAEMJD/Fkv3JaWpfd0X
Bu6rPh2kc2aD9VGqyVFgSSy04Vst6AH+I0Tgf/NU9vS1sJVmlRiiOkX8KkGVqX08
kRTk0+Aryzt1KKzv+ZO5bVtr2rsQSFBRi0NGOTHpit7A1yqxiPXJohFcKV2Pd7Za
94zGy9YGyA7pqQleP3xJLgE3x3BMfyCo3av5ilkS05lSqcosG09y08q5KZ75wDcg
4UGGqcqlpQ+ZA0WJi0yOR71r8EDiGlCZYEfx/U+AMNdXuSRQZZO5vBy0iPOkFKk6
ri/L7zphPrhkOQgzVsc5WzFO1jnn8PSRzZfIhlKw8OmfOsVdAJhNCvJD9I1EahKj
tGmxFUkEbRMjU+3L/8UD9VMKpVmEFYZ9Gb8Qu/rGJs3mLYTmqXhezay6JOoYGeBW
mZLBLZahf7/HpNpa3y3fSh95eflus5aHQemdEHPAEP1ncPVZVcgxpARsTYBfQIce
Iz0EusGl4fk0VUUeqmBhKzUWIDlU93CKjlln7y3wat8NHHZ/OLR+CWWNbDwKSIJX
0GOqlfpGkRUKbpYtrrtvBTexnUHdrbJwTJ+es8S4biJdK1oXU3Txdrk4TIZHcaCq
zpB1eK2dP+ke61l/j03krw9eZ1NJZ45lGXRmSSsAAF9grHc4PwL+FkmUyS9CuyHB
gij9Vhfx93gjxZjHGI5oWnaJv9BR/ttjg8lV50OgUN+jYcyryX3eo+hKmuWnkott
xMMyk2EKoeDuhLb5+2DE2k4jehPp64EqTnzwRI+h/naji7AeZmdGUvEVNBVCqwMT
1ByLy8emLsNKlEEoShP35FHTJsEbUmALvnaJeU/ixc1dfIvysoGmWtYUEGUKmGkZ
D0RuHGG1i06UhDzGddpIquIGKi9ccOJ+AJUkT5bpzn+uCBEvMS8oXBmXKiwT8tY3
e2PnWszXEc27h4DyjuOvUUeTNsh8qVCCAhhhB2YpNWWW7QnphJ6vU+TsXLw/dPFI
V9tjCPS5pX6jvWKGxntsu4slqPvBJXlYwZuCv087+BJZw0rlycHbrTBlM/Uns00g
ujNocFevFKPnrioJJTzX5JGIrAMNVgYWgTVyETDzEaZ7S9gzlGRkgXWzNdcw4mjU
7Pi0KmYritH1yJYRpNk9l8N0sOROVw0qfUwyFZMXOf2wBbQlAohBwcGFrKhpENxH
LsyFSXKcR/NwbhRCPW9XPD9kT2aSpE52SzBlBDARPSeeD1D86ywR+LeTvWgdbBOc
2ofwPFpmMgc1U95lhqmlXfK9P+Gn4DrR1oXDLbMr6uX0pnDyTD96Fb/K6DF9nDro
0mQ+cMWU32M7HjjbplCWQU9G+MsZ8h9NMLCfnGKcwPKw09BEPcFhPQRUAjmCZjzb
SFaAUc+DlcWVkKb4vVB8GinFQYGYGFzaY8L5oFQnzB+Qk6lqEHNWtNmQDR/vOkxo
L6h5bZnWxeFVL0+kmKJzIC1/KqnFHI+O5o46b/D1L3Jcy4r+0aeVZnTU4ci0uusG
x+XYW7GlxodRpW9HaHklNxpQe5NvgGIODU6VnXxwWV7BAdqBd2nemCetNVzXwT5o
El19vW6qso3UgLSfh4rMH+Dv8VQG1f2JRH4jpbkSEAyBfb0MoPjEql3dSFMMvQ2O
iKzcc4Y/VxNnKgTrKI/KAeB9l96rDeDjl8os3SDDvC5KVMhJwaHeFW6Jtk1E0U6E
ATGgfpZKUHLTib5oqPXkr/s73ve+L+zufPBH9eCaoQ/bPpKRewdUbjwBUqjxX+sx
MUz3kiB9TgNz5VGUrp1Dy/rZ1lpP9Svok33rRmfgwUVlgez4nlf3lw0qstPKoeHO
9aj1fFbP5CUFlX0IxmLfbRGci8mb3P9VJjZGNsJ2H/DRCMy7yQm/2FbQCCm6bmAB
aTgB1Z47gEkls/RhdHTwJoCUFD74FP1ySrKjwfl+7UAtyO3+/UeYkxqBF8Lj3Wje
H+05PrGrzTmk539s5ORJQjDnhVXzveuugvB9cy/bwM9qkjk8oZBRGpuHRE4QJ2K8
35Qts2YpUYJ3nFj/rSQDMTL1t/e+lNjW7vSqgKSopUDUzy5Kvr9401+ElFaTmxRj
U23LHZca4TlDVwBCyaLn0VhaApLi0hSd75y3cTEmoIZdEKbFX8JSdUGXVnPlPrJF
mxt8fMA74PKzX3UbbOE0U5JAG79neFsdeNZJLVUiqYIMOHWs3LLTJz2UEG5fvztz
BmC5nlNROWdP41Ta/ZOykWYksvZgnwG0FjziKfF+XlDBRlmvHKoNXV+ITwmLeOYi
XPjr0chfYPEZPi8thzNfeA7QwyoXV2FkOeov38KFy8wuRc1RZ3BsI/UjZQCcr+Fj
6aetiLQaQtkDPqm/mJ1223nZQpCMF599IJt5WWKtbeheE45Jyaj8f+eWc7S+T5XC
iTByRCxMczmhFQ9BKIPTDkvM8F3DeO2y9Q78TGFcZptGmNo3o5+DqODOgFuDc5Cv
3Cvt3FCu5KUuoBGDIYXtXeZqOGi67mYlNsVABeLxcP6SmYZxG+CYFoHaq+uBPZDJ
SvKj0iB+m/PE/ZENbpUYTuIt0loti5VEv3POrrMUPYNV+jAjQ6epfG5lbJkj8RZl
lG1dk2fzlBk0x2tO+P5JVwuxUDFZqnsXiXlP5XvWZxZWmhjWo7xz3DuTT0w9BMjL
SlPqCzsJRDjS+P2w2qzMH7cb42tjvbzXSfQ6nmvGBaP/tfZhHa6AUZpDHyFKz9bg
Btb4wZY9Mrt9jpCpRmNRrgJT0ION5hpBJ7Jo/KEi7do1PLt/+0ykdV9A9Ydb4rA3
lZpqh8HWpnIFEj/OoP70CsmVxZVM72jZQNXIjVv/iUjO5zLA4g8ItPiYMfx90Yys
9G4Na7eMGBlKsujJ3XbirCmW7JTTETk188zuDs+bhRfVJWxeEUxIhpMxMN/4I7A8
AnABTk0NBfcrrBpl3Fw6CFOmpOw0QZqE+BovvBT2xTeRR6iPPX+nSBtPtyq+gT0v
IwLF3D4ISwL5idHOF2M4l+MJ7fHkBCp6qRGrxBtOGIC7JirPXDIToJkvQmzKESyc
ulAcadcROBOJSZeXqYKj7wvi2tW6Sp3p3yY8DNl9pYdLX2Zg9tuMtctb6TZu6nmK
TUsb/PYvMKg9y5Tyyzf1gJfcFJFswrJU7Hz1WoQEeiscL6RPXoc/CB61lxBGbRRH
dSX3CQpiV3ZW0FpN8FLluYKTGuOIdTwWWuLJo4StpoHaJ7HXn+LS3+Z7qgT7e+b4
DS1mJqGrqIQBOW15DPXrqCAWhzdwFf77Hl51ob40bW28VYEGq4J0EIJSpV+cvoCx
FiuybVcn8/ZI/NzkVSObGjqpP1hoBDloa9hNVRJdVsWMW7epdHf0IqER3f8t8FOS
axX6YRv6MfaTTplDSF02VSkhKui2UDeu9dWEk4y3Hl2/+TyERGeWbJ5bgGZznek4
zYBO+8be3hyNBFs2bstDyWnteILtPtLV3ijjV8NE6R/4fpbDL5uj+fvS/HrlKMMN
NPrfugBbpzvWNJGyuq/s+sq4bUBXhc3BlyRm4iOZek4OJRbb13cdJxjvpXQqzc/i
1SWqmuZxv0Z5JzeTu0PZhzwxbYHRSjZcTevER1GcxBHvsYsMDtAGEkS9OG2HcI+H
GEkv2GXUAhtHRIASj8EzETp1iZkheNQjhI63wTUkDobB0q6bVaOBEedjMGraGqiw
ECntKcqyDXx1v1jDUmGh4Ej1C7/VxlVTAn3iFZfy6Dz/7tsX2QRGwgWsmvEZfBx1
yE/fCSrll6MLxytL90F/9MTAPC1Q1kNOCvEnB3YwFhbpID5hCNjrSfmTu166mmfv
QVlGGZWMnWT0a2cskwPM2dc4oTn7JXHSnZ67f+DlMD9OL8In+CcbnfPmu3wurQ+E
TH11MdR6dbN8qHTN8+N046pLJxm3GWc4OOKd+lnZf2uPnmf7fruo9IUKZ25tkMlJ
o2LLrDNtTXNsCDu57xLwDg+p4jMwts97ShnHcYBjWUi075QislUghvS0XLCAHpX0
z4rWV9mR75RE44cZeiWzX+s5mRSx8mftU0oZF6uzFd8xClfJivFeKyZsbKWgEDp8
bEOTwzvXVCuIv0ResPQS83ZTmFu0g9FcDONaKfCxJomGu7sGxfvSxsRQQZJou5Td
b20tijNAMsW2O4NEeFwAHRq0Y1NQuj1mejDV/5OYxwc4tqt+vPSsh3fy3qUz2Xv4
XIQ1+TxPgS3YUwfexh7f5mLEzFpQCzwHxpsVNQVk7moKwlhQmr6xFr12MOQ5F9wY
48MEtk3geE9MJcblBoWMHtTHXW621pqlCUt75I1drKQF+22o95FomC/5XqB5Pcmm
13CNXOjiO2pYxuGhZswKMxFqv/YFCC5aQ1T2vUNTXVtYUpDzp9uTZtj486PcMQSS
KJCiBmPE8t+4oyUFjMqUSu6Iv7PNeG1sP2GqDnOrBH0cSGDvb/bG6EoK1v549VGd
n4xItE7iZLHDnRufe+XxjrTdpt/nmNaVUz+MZpViPqFyxLQvJkG/OtG3IkSMY89z
yHxD7+0GG2ZGBN9N3JXbPC62Akd+rxVLP8o8qyaaGNv1uGMK9UjzPAGwlzcWUUB7
KhXg3ijPTvbMRiyrtm+jjxaB4dy8sRZzNQif2/VwpDnydsLAm2z2awCJI+PVxxVB
GaJXMgSpm3PSog50769LqvrapIkqotkjQGR7v8nfJayJ3J9a3eNAaYQYbInq7l9G
vu+Cpq7olv2xUAsB3nLKzaLOZJT69Zywf+mxDb+JSRzYUg+CZNiDQz+A2AvXk/Yw
cVxX/z2B5iODRBIWl2UfS0udAuXhfxR93QaDVylJA3v+3pCu4c9Ta89a3UF79xCY
ew0LU3CQrCey0usjYS5gkd2V4CSKXEcQ9E9gCl+gW/8R8HFsz9bg0y/Z2cn/7BfA
bXE953EikA4j8x0gPcEoq/GVBAf7P7ElRUQ5xCJ3Z8EBkTXN20X074/FQ+Fj7IVa
oE4DdHU6H5C5QRkbJQJLi98q4WlLNaFBdaKB24wUakUgTIud/xf8GEFvUGR/HQ9E
bjOU/hDTbNVyw30RNRbeJL+2/B3ipm1kei8DzEhdA9bpcWcOQHq5YD8BvcXgzjgK
mEyhioxvIJ7e2YjgnpcK1eKJCOcsYdq7Y71pH0IX+TDB2AKCi04m+Nr67WZgqdZ7
EvO7nCS/1bCnfLnLpFCxdm7l9N8CE7LYcimMA+A5FyD+aTEAnZmM6etnqx38uzED
ugRW0xPhwEHgdtTBNZV8P/gQOixiL/UYyPkQctFJIXovdbGfUxY/QEaP0eYWffQh
RaDXRITwxI8BbKKdvTPthtNcMQDD3NwQP7mf8RVcJ6+doUyrPUL0I//g4qBdx8LN
7QEVSWFh5Hf0W44Yrf6JAGqFOUA8lbbEeekqnciqiVACKevlqYly4nQFyxBBj8ga
DcoqH6V8WDOhMkfAxgJpmOa/CE5Okg8ZoYvlMI+2at9+sXlrW/6eJoUXHxlpKuGT
vLz5jOdv0XWk08nZ3vDEXZiQLt8RQLGOvMZcrDuW0QyFFVihB1nwzGtmdFBdEbq+
49fwzw1UBSYSFgFIFRAf8B5BazTKbVva/yAqXVQyf7RYrLGZfJTuQ6vPabpvRdA3
ZgzrCwDVuE6OalRVTaSheqawQ5p7itdCIxh1eC1Gsw3iO8N1hqjq6q+VSIrslK9P
tPEzqMUturlr+h0iwOymiGs0Oow412XqY9Q9fpcReumcYD6wSF1bbDkQCSkjS6YU
tDS6PDAGU6Xyekb1sDN/dr9UldZH/giX41Z14LfXLKnaYpLzrwnHYuMDsFlhjVXO
DyEXBsBOM6Ub9UOw7BcaPKOj/d/FVKQl/fGZ2Rfk052bgQjzZtYypaec7aStP5IA
YxmcrstfLrircM+NsZjqstA1B+Ae37OQjr+drXLhqdVQPaLYhHbizLL3X76nV+E4
ONrp1OQ32fQeN1DX44lYOl89Dm4tV912SN6t7BhwMJ1jDDEtp6Lc3tGBGDP2PPnh
8+b4L9KIL3mjADeJsp4y+igu5cXYZPSLio+8SiACFUwmiA13/enEEmo4hPBx9QxV
A809YdnjsVYpT8QtdeI28wYJNRWIXBS58JkOtoRn1Ibf4lpidR2hl9ckXOw8KBzz
EE/vbC0rHbnk/E23kukoGwR1kZ+0SskDRpLcCr/RT9CaxUVnIUaPcHRUqlCIuaHi
na8T2R+Dn75qKKcrchObImq80+hZsmLjNRBMMrV3jA5ZuwtBBKTNGRqOhRLsZjCt
HzzcQh9DYdzcEBaG0DGo1DmSYtBITK1SSlni/8J92uwQB/pYIWBLWKUtCy8OvXOo
kS+jus8gQLLMoP2oLCLz2P1oTi5AfRtxU6+601G1ocOaXk4PNofH/XRP+l9p3TOx
YSVKjV4NqqR6n73BFcXhMq1Qz3vjwROE/XsLjUJRMOwH/w5FBxZHy2nDg69a7dG6
UfSZeK+pTDchYRZme4pzXAvhcMlkP2og7bUbfbyHnZb6IVfzcLVcMLyD9RwqW5vl
wNonRDbN/pVDzUF/39hNTH0KtwDImYzDQtc4pyYyoFr7GvUFbptd57XVEESnREmJ
1oeMOGeeve+5yVkPL9fO6Ukp+qeR6bDe/c/VcBxzojf8swTKHMuiJpjg8pY8J8sb
0d2D2KSs5RbG6uWf7IHCIrM+rJkhwEoA70cRLXgfC/qrZapydScP4T9dhYiQHfi/
YmiwNw4HzW5BPir7Hz0Tn5pz+CHJPwKYqeJ79wSIhPmQaq9ysajDHeixo8KPWF4W
UImoO1PuUy05qktqE2RrQr5kjXWO+MrErKxSTNmT9pXanLaODCMjO57VROSgL5U1
Fe9v/0hokODCO8IbHyjFo7qYiPONhY3ZDhUszQdqCbuCKviWHUzoZ4FQXJyES2l9
xCW1qskV7TiQgmQaElR4jGcdXl8aoghKZKX0Cyk9LIVIJQeFuHv4PBYNxkiTT3V5
VGqRvYqL7aJkyT9QtSdY1lpldw+uN3wby11HhQCHUEZM+n34zxpjEn4Gz+bbUIoc
y1v7mc/YILH3MEyZ5rpMdEMS5KAslum+GfNk3a+mbQkRpn+uDFM9g00r7jJdawTR
ztBCUmKJUHeUQY5TtI+X6nCbMEGPyVcFRJFC+w/xfH1KtuVsszujb/JCCqsLlhHW
fScLjpXKQkujbOYjwQ+bsP1q41l96DNR3yreeqEqc5vm3D6H298kXUCwWHmNUqCS
7ml0JUjdC5Y0/BqciKEjfrILH8MA1rs/PoZzOw81SYrcCvwiJzentZUGpx47fqjv
kaIoaUoCGQZWvNOFYEqNNaNsLFu1dM4QQzlnT8UqqrIr9ArqyoqRyqMXhMncB/7O
jaZj+7TKkilW8gGdVA1SGTKNoNLPme6I/ySK5M8/EkMxnmriy4kaKZPf4bi/vZBQ
i3iotD6m9/IGmHFz1jc0iYLm26Yc2QKVol6gRomhzfsny7SMt6lt7n2c7TrLoC3d
bEU2LOAwtkbLpdh9YvcWDsCowWlAlMA4+FT/hDt0hvKWEqwvXCdooYhMQD161S/d
HmyGHCR+sSxS5vS6FKztYWi0dNA+6hB754zXfNYWfnw6fzCRRgG9oTX3QJE0WX3s
GhHeCBUVuEpsESIhvZeQBzY90dzE9jGbyApB47nzIW92KfaSaGZvtzxV4x0Ox8eb
q6BT16beAxy1XwMK5vCQM7RbBij1E+hjifk+jyTG9VEP5EMbClvgElonAd5IJKfu
NTJA/4GI50s5nGnSAjme803l1MIMokaQnqgWa/33NOJcFo/w9jagy4asd3mFBH5q
xmDCpqEapRUqNaqAmeE/yodFi1ATTaf1b1c21cyUme39X24XFhBVEA+5tRvqMFJK
Zff0WreIMCHeOqxbJbNvXnyf5Kml5N9C2kdewvFfV+k+GqTDEpiFFvols8o23Q43
KsDb+nJ56IokT0sm9Rih5Md3xLjWkcXSOqaJkAm6W2sZpdT+dSFqetfGKbF6ADqM
NJ1rilKi4VhVv0RZb7ssN7b2wzpJ+QQwb79xKSKq4Q6nYHxcNN6r3uGt5HsRaRWZ
PtoigjFCNaIlemJs7Yk4tYYs3BGG+9nePyyNiSeNaidzTEFBEO6j5MEKJIsXPZZu
HVO5/06e/ADGfxqcOuWzIyD4qhtOMMx70xpaqdEGwxIUKGp0xjOK64sjDeSnJSs0
Hj3hkYlHry1/VFJztncUOQtejGmHdqUbe53m4ROPTcogiqtNABzKgQzZDjDtHUeX
LVDiwJC3N9TnKTl76cLrP0VAVZhn3y44fUukmuco0TLw9kh0IAhLSZaqNnYZXFk1
zLEHDwjJUfdpKahaoxjwf05qrFRiZupVDXJQiskBkNnAz8bgfW5pABvs+Wvk0J8R
JgclV8QxE1oBXZ4BeFwtz3b4ypuPiMpyJznsHIQ3GX9grbdNqh/3QJ0HDwz30OQn
AYT7R+ioo/5qXT3GtoFg6jaTpGXeFwWU1vW22l7egDSC8P7stehG9va9GLRIniZ7
jJxg7npmplgBJJlRrUkz41ZhCAoOrXmgdmzGP052yvR0KP6Y8vLbs6pRXz8sfjre
KtA2HwEZEE7FbctTCg8kifzq5t8J+gnIqSfmSwLVWse8rxyX4oqZ4TpiG7MKla/w
+tHqEXUcdKrVznv74T90RdQ50SItuBcX387nau9FmGribdC2tJMVlWFYrFTe9WeB
3JwHdTcm6Y+4WYRP/8Y4toveGELVKL7LMrvb0+p+oqXoupVMcn/ClZ4kjd9ac4GZ
UxpYEuxapB8Ec2aCzMbyzgUqVWAZz0W7shAGPdxmNfa1UOroYUvnZ2oJ5968wf0N
jW1/6njvCP7YnyXnoMxhhIxWx7rVsZ816MqdJSCPUZXdm586X10fOj5fkfJm+QkJ
AmgWPyugjuMBWEiwi2w1tcSrtLccBfQT2dcS3o7kOverv//7hy/lHWgVxmUfW19b
Eq36saMS8Qca22ckxnYD71mZNMDijh3wbhBWO8ytwdYo14+aoUaIppsK+MNHBR6P
aZVBv34q79WSk2tuJMTwkFoXvUiGGhFBY1adLpuHhPr4PGevts62lD9kJUAT+yHU
FPiBGUreOQ6sYvdieQrHyOE0Ft4ovCnS7Zpaz12eKL8hEf+VtckeaWXWM4uASiiN
fHDAHumFhHX0v+1LNdKp0kX5HL/OajT61wlXDgw5BuvG+I/4ew6vGNo+dfUEMUJ+
f5WOznSIAYuvdT/k5SdMREBd8xCGNqgoKl66jNBO66Km3cmaTHOykUmjj/h7+rwe
vMRpsomThVY4IaKQUP4VzM40hUVv6mTqR7fI8hwOy0LbyzGiedaIcZT7HUMzZPbx
EyGXXOhrJVxJGmnOoyycTw4J5U1N5nHEorzzzyyU+mxaahLAspEBIKOyzIYDpPCj
KArJEQo6qY0U3MqKc0pA6RDNjn7NUy2LsU6mBilXERsK3YOqtZ1wqFu2Y6IsttQm
Jp6z75ocyBfMIXcopaiy4k8UzXlstkIFaAu+CCO+gFMuh7KrCNIa8TuBmq0C0Zl0
Q366Qnt5RGniQzMjkWDiuHwkDmuq715R85QW+xGRXFx62Jm2USnKm58RD9nNhYpH
sY0y/qxY//GDnvnN0sXcsHykXSMVtUK3ieK1nCW+i2vykUrta0kqQ7vHB7rh8e3D
rACVqsHp1whLIAoKAc9x6BYV/+MhpJ9qMJNwfRX+uiHfEmiwK/o7s50j6NqSJT8T
jWAsHJXidAqmlhV6Z8yZa5A4vTQtYv9Ea9DO0RhekCrKoglTxoIbLAD3xpi8VdsB
2asY2xYnvhaVKgLjj3vsv2UWRtWH5r23RPMRBtAwZ6JYTKqbvBoawlExcP9MBQjx
qMrULItT/vC3oMYTtiVGeVnLqaSDPcz/Zt5KHdbm6eUx/lDOwBqlTiZXu3FytSPx
G03Gyrzl557JUmxDb8ev8QVPX2UCmVOC0eDs6uDHzMfTN8v0X10cGgjlAIM55fb/
5W4+YddRfhoFhGpkOaosRIeJVsyU66uRc9TgwB77D+QzX78KXReiWmIDt57G1OyX
2YTWQrVi3iBCFkLSPON80ZGVIenwevmA6hj8m942L4TqGbngTZmD6AHGFYdwKd9J
y6v9Yf/KFxcjJ6dbjx/f/f4aeUAAgELic4TxhC1ARkihNIFAtVayie3cwL4DJwmo
/g0TwTR7IzTeq4lDLCYyheDatIB6tO4zwj2v1NrpF7Ew466+9nq8I+GSQ6BCXs9c
q+v3/FW/YdqxBCknVl8QSi+VTyjORGi1H8gRJqCCyj6PNuTgLbjpaiCvuhIGXJdq
FWviyy1hhbQp7fMzUu3YZxikuLwnnTwEt33kBsP0g0o+cPCJddHFzKHKlvlPp1ef
I9GewRptj0XzExExWl3/jAEvXIke+e+Zcz84BtrUYL3e9zY8i6YqTw4jNJM5Y070
G2OqiCq/Wk1qWQ4+QpLunORF8f+0Qhwk5azIWSPbZaZfOwNY4UozMz4wFZgMSLgR
A1wZuqVojDbIXc5P90g+0sCOI3ubLPU/7G1J4j4J/ilpzjfomG95hipkTfwifIQq
6/P2vpVlc+7uL9W01N8WeIx1zw3MgNb1eegAYIN75RA34DMcxe22UrFkKioLeeBJ
aIx7Ks516mTc8We8gpTkSvt0ftN2OUwOtlS+Yo8sRZnzBowO8eJQqNKi/sVPbvou
JsTC1MmwGXtO3EstFiz3e6aBqNV1cHdH9UlvJH3RM9t9azUO4q6VHgMXr3HkVgzb
Enewsva4QeYdGt7RgfPU/C/C1CW7rRVV0sZiRM1yJc5Mk4d2ndcn7doI5ZBHD/Ki
YqMPsnCf2W3X1k5EtyX5zvj1jztL5UXlDHQYWBioQD5Fn5B5dG9uVUOhhbVaZJLU
jfaaCRmhUyLadyb4vNloGm/WvsDKvQ3+Bz03j0VVfiw4z3UDVtZz6/O4w1sDe7x5
07OEADm0cPMTAeBhg/BPAHS1fNt1jOphs4hHLnRE43eUBthZeI+/R9gbrMWPPoMs
cFDcnaWl1rzcA1MIh0YBDoV/OiP91RKKQpVNqfML0btufLt1owpkqQWSXRJZ7C03
yVbMu77muTCDJIVJscEiONarMPbntrt19+YmL1p5aYMPB9Vf/C2Zwzd+X9JuHX2U
JYKm7VL7AtTlrpkzuDYzS19sCHvYAojupEdSn6dSq1fk/jwETbxZl622bP+zD0WA
zjcB0B7ovVkWddzQfu2l1XxW/TA85OCAOiCjqi6Kdj33HkWDBsfETJVEM+zoAG90
gShI8AIZ66/eLqUSTlApwjlVzFMWNs4oEEJfBbNSzQ+OXGuCC9snD3SGFVn0el8f
ceZ3wh6EglGfyCfw8wcjY1aO88JShEH8yGb6wNrubB+V5jEY/D61jqnRmGGiPw+8
2dpB0CkU/HNPB+qXPv3thsYkYOPa0T/heGYzu1C5rv3omr9GUvrdFj083e3V5uNV
6covlHf8rZZt1S2tr5GKhIpWZCC8ZvHVt7tmtHXfG1dLHGZEQA8kbmsU6vv9SZGT
8WbGv3hgiv59ujhIzNwJDMLvNWIWIHvVniADvWTZssZvDdUhmVXUjpqYSlpiP79p
tTuXCQxDCQdegkfvM2/Rok3L8x+gpwrnsQN6yG9LqJAMTQZndmHcnO8znClOTZFt
qoGuhpL88VOdGgTw0NxDNsbVgdpyLBX6bBkItko7KGk5OfSQ/0EnduAV3ybh7Cce
i0O0K/MCH7XohaZmA4cpKUXnsEp6xSoUFUrSSmfRJayyTGejh+FDFMNkJE7JKeBu
J0b1USiN4/NstgxKWv5ilQ7m4zV4R4GqC90BSqYGS1pe7MsCWyVJeiz9eDx9J/RE
3BWMCFNulswZCEeL62L9K0ko6B0XqzZrs6st1TTQ4a5q/I6vEaBMn+0wFmKkt9MK
eIQQ7HfTWKxJDgtyeDRotoKJWKU47dTT5bIE+aPZHNW/aGD90kT0By5bLHku/29o
csivLbasruk3MMnhAlkbgtldtPdFdTCoJBKAcBfy5bxS0g7eTFGg9lJy9PHIBdu9
2u8jvfC5LOIOIBGGgRUWg1zCXn7MD0vhmI6Z3uWXGl4jXOTsJB7qfcAKmHO02kWA
CiQLS39vElfbDKXD3pVa1vmUVg4UrSu5Jh76h+RA0J5QN+MyDQDxJUsFOZZiIxUA
KrvoCAt4gFG6DfKJsOadtgR5LN9YrGfdjNQ26TA8XWqE5qKOuFRKUVhbJmwm/IAw
BZ4tlqbwJyNsxLR40u8EGwZ80FWxZ/TvdNXJbJj43DLkp44UzkOXOINCLFqgo7IG
aJalFEDfnvzkj1Ah+SCsK4E5wuKZ6jEkBERFWObXn8TMpgt9nfpxYXPl0X+L3BgS
pVkIIDxKifzmEna8/JTTbmpqTjRwB8Y6TOBrv59tG9mYevEzBRvfmZ17fLGGmopw
TEi9k2GIulKY0x76r87UgIjXH3DWWUtbYQZaTiSRNXxb3Ys9CoIdbroLmi+DYgJy
TZfFXD+0neR+6VGHmlAJ6VYMcmOu2BQNjSknNuc5WsLJIg2ftx9luEGLN564VCVE
5ffeDT7hSaBg92xXtqv4lFAvM1xxIkpD1AjtPmNI96qYe3XvjSq1LscG5P+hqBn7
rntJ3Y1/RFcm1orbIOvluvoZAmXZUsOm56JGwLq+OWe9KtcktIcK7gIDBvXcnv+6
sZkBxjPzj5GvNPG0th81Xlja4ixX4ltuG+LcPYZtO6UmXsnmkrOdDKeMpROKwkhv
UKmWuHhjnsbjRfD3HuQIkIV1nZHyjQW5Nq2J/grhh6xZ4NHroqPSxBxdjQBRBaLp
NGpiXs+AasIh8mY0YaCsK8FjTN0Z9HIKjAfsRCrAahfqJUNgIWKwFI5c1/BCG757
79gMVa6gRqI60oVs+pJVqs82BVdxk/LTe+PWOcPmfaa5UU8uzgr296OE3JuNeHsF
KGRbJd9nqw1ObSZFoD4Et3/C7PYhQ1/8mf2sW/9s3XhuQ75B3CxtkO+oL3nWtL0P
3PlBQnwW3LOaHjUtntJcQq73m5W56/gb65fY77oHRmWXQGhdDv9EQIzk6U9478+/
Wv9IvJhbWAlkHne7aQnEreNZ9L39Sdivoej3KY0m+ylXcDU1lIWywz8NVUQ/OnE8
o+71na4MamCkyz1oBPF4QTMgGvbBmjuVz2xWcAN3lVXruxZm1QuqiidRJCuGtuE/
TOMacqrZlDp5FCf3gkY9IErdGhKn6/2sST/O/D7HLm0GUJDLSeLsbTRtaQmhr/KP
h/OK7V64/Cu8v0qvJChJbPrHJvIKuXl4dFyM8U+Dx2d3T/lNFX/TKZQhFiNIVTxx
fcBo1eDRGvV9bd/IB6dJFgl508fraBKZdVzSxrNuwPpvBMS18Dzl0/YDEdRCyLvQ
p2l0Llp+A0jRYlR8W2HPKgLDcVuEbF4tlPHkEPhBvRtPA3qpmo4rk4s40fom0UT6
TOhTc0NBO/nuHo33ChGr61BTgQf2kD4ZWadIVAA4Z/wli3JStKIYXJb8+WV6jnqy
8cW03U2UOmqF+oLu/Zy6uLtEQqLZa/tI85iklsNTTqrXfvzpOcO40UXK0rN4aon8
daopBp0YoYMkPKnUiHteLXJfmY2XDI2OSUKbnnlNOXo7KblYKfbAeAavv5LjlTVc
1pEgLwVbanmTcQVT8Q73kPPMG2kl34Ln1K5qeq4zKbWJqK1SitbfWdKMxRdFGUZu
B7943dN/2Rrdjj63IEFVgZboa4YZZLZy77QCOla/hmhR5L7wtsAD3Z6CRqa1SRNT
8HACVGJ7eu2voelE7ev9h0sAToDv7nxL37AU4g3xFajLBvoSkHLInsulVtek42B1
PlPotUAavfmB7wGweLXX0a6U5P5595gJa14E3sKk4Lhi/OYTaixSZDkNU/q7W7a8
qodLb82PFxLYQbMQMk36dtJsTRoW80vUeSktU8iJ0vCa5AqFMUUKSEALGVEetTYu
BK+e5tL7Ucj3YfyDcezTvWkmnhLxOlD5fslKqo7u2UfLKVaAtGRwTq7i1oQfGOfE
1Ppo8clSenEW3GJi4LhYkYfwHhOch+eu3Oh/LiMItIuH5Kf6Ai/iYZA6sTEhHOeT
f+F98zRBOaE9Z0JpOoL8fzneuE6jRYjPC5hgbBnFU9tFWjkIKeD7O4RkaSCm3nyR
TiFat9HECaZT5eNFK8fDN1gBrnUlmrac1MM7R2PY+T3ZDr710unKetcZTr2LJJXu
dYs5cbdESG/pqaFXbN4F+xbCRgQ3KIlKzdIHZtfepY5wK1jcwKS9c2E2ANFVZhbo
cdki6dtL9IOPmPsEMXK752Ne+CltjF0UIs8+umrdL/Go+9xzKCMBcpMIepW3+CuW
Q+lqe0xofRQQRs34kyN8ea9DWSijg2L4q0FDnBgReYzvZV/RfKfiG/eht7C2rLoi
sSn1N+9b3+eWf1NfeXijPAg/R9LTPIaYTgy81OTodsoDX14UXQRwo950oJ+ol03H
bnn+PYldL2NrLygzZ4L6zC1ZuPicfscPeygwR1E+ZJ7vqgFc8NFKEb2r9CXLIor2
CS+BVcSXa+dtKstKHXNV0vghj1ViQ7bMEunSM9QJg+cQ7plW0DYkynIN4AgX/PFN
yt2JEkbOoscjMcJA4b0Wz4FRM1+F+vd4qqqIOFK0CmxSgf5o2QsgE5N5kiU3FSVD
8TI+eTe5GzTokeJozjH84iAjOUXPhb4w3n73DKQemWksf6tlmrPxZIM1W6/O3786
kBr07avDSBAIumyT9t4baIslTPE0WvfISd1fXPrHIyhshUBX31kkxwKRqxhJRFH2
q+uImKLhTFXjRFCJOPG9fbZrunU9eQdNgp6jO1BWDUjlK7+sTHi5OwJ142xl+YGb
3Avd/yt0xXepcrLA+E7fFeydnP1pNSwma6BmuJBkAQBqw2sUzQDorNE/xcSEfdt/
r/gQM3pjg8/OYW4+aBCILS+yuoLJdJpqLxNUM3cI1iPRcM5nxM1qFpvRv9vdZJtP
7bzq+gFaBKt0Exf17FauKRifCDbUj2zUV5oumlX+xz4wzRgRxc4c6WimWHShsVa2
jCPuol5x0D78LhwFuwMMeHqLS4x3pYnEeHhFmgMPPAnSvmmhE9eTCTwIuduZh6Gl
752n/P6aoU7mdA+IAUcHs6iiEAE5DwEsB0f5kA+dDXKf6guW7mQg8/dCpHqAL8wl
3xfc8+932N8qQZvQLb1ksecIcNhxJj613cbTacqMwrOico4WhChY4HO4cH2TLsOW
dVIzb95EjCN80TQqL3RwwdBPTar30YBkII3OHf0l/pJYSicYbD+kELntvIUuf/nv
wQow7Z8W83KYimLUJ/7AWiIAh8ZGjjnpeEIMj7hzXfdfaRPm3SB0p4nPr/+ezpYG
syXa8UPgmgdWWPIQmD8VwHDnDTx3wy0/ZOZuiI2t2vuvGBaiWhY1heuwAHAeYcEB
qsVfTu5kWKHhZe3xBF7dN2NKb5RocbUzt/bo0RNhP1xK4r6wYrlgkV7WWTh42NJ7
iQ0yNkAKy6Rp+M4dWogrtD5pEM4nBTdpwTO8ahEUJvgjJpdigjXkQ19y9oU94v1s
tDgF/cIi2fbeYEX/2yGBwh/rmBao8CWG0UlLym6eXMvFFa1kcHx19o8q/uLcSlJq
YhqSASwtFsJ7KTUPRIOBEKU6XlYLXAT9PN+gvH0wvVAWEPu1TfPHwnBRCasp7Xpr
JvWMkYF9z1HX1wMAyul9CAKhrfwg9mNWaaAHF+ae3gVim30arsIfgU+jVWX9cl/a
8g8LfhbuLMCJuzrLdhPO4TPrI5pHh7Tm77dxKqcFgBHXl2Fuo9qWJjqKmlBNKMuV
BeC56AYQmY0jQE4jvftr3YYP4oQML/94iJazEMey7NiQCT85TFKluGh973DhFgSw
vmo7/FuNSJgxAWPHu1NO+kQ+sSuPqTWFqYxyP3y0Ps5GyCCkdqDYjkYCr0MWhJDe
54QRMHvH8W87xMnY5ThScwnbDI+R/l968mTr/2VV2OQ+aA6dafR3Ep0t+/u5HCKU
peP2Z8ogYVwkekDri9Mu8z0qED75wylYZDm6y+39sisQ1IPog5nksKQ627fwLMP3
OLDPF94BpXrgX2/Yhnh8xgKBqbkvJwKQNhrifHi1DbvwSRA6kccu+Nc1aTvuNXPI
S4GVd5IGBT5GF6PTj7OwxzDIiCNeKxweA/YXP2xy2JJNHN9u8PJMXEwtqKr1uvp9
5a+Mzcx2BAKwrysqmDy8ulO0qKEdREOyVY/LYKz5stlBPfITGE6Q5jkF1rOrzVKp
OZK5AVBswn8kvJQo2IFVOUTT0Wq+h3bEn78CIVKbFb4xAaR0LXb72ITVIWxFVWPq
+12z4toJW9Oc6pGNkCfyHWHaxVf+qoIXuBsQyCSw1HdgK5Ja0tIIoptub8I11HTI
h79B7aYlggIj7pq6UQO2VTPcOk6FeyDjy3gszqBYYT5Eii1KQ6NxGcyDbgYQnUfz
I9lw3OAYUs+fYe/j8LJjxt8HHOd0/uSmpNb9rMijcRrCU/SlE2LSt0u1rRkDNiyP
8HfuQt0PS5ryLgjKNQVSa1qDoh0kfPoLBqzzKye4veJk28JduwGCcpLOxq++uiXl
LWxAGgKjzhui4IVDBjIZu3C23oPOfe9WnZitR/d48zMJtPMdkKZGDlojryxXIQEI
4UwvVn2hF54k5guOeiyb48MEmkgzpjSbVuB30aOMpECYkcZyYqI7qxED2oXvYEVd
V3S9t9fC3UXEgQ+Eps6bieWd6bh4VZlrqHXD8+E10bP+zUdte0BhpqJUv7Lyqkx1
OgdO5wyg4RaA9HXYUlRP7ESgDFclKqt00NiKmW/UD3Tl3oxvQTmrVN9iR9taasOQ
wswIsEiFfJUnQene4Q2+knO3ISzQjw8jS6xTkJBiBWc6MaZZtvWRaprFvO2v7l6t
TWkVPSM8SnejPJep4RS/07OCP4f5YKhwL98B+zZCkV9Sofjo4VRVIxTyDd559h5c
G32gtqaNDPykSMFRBWfIV44r39Mh7jMRqNKhzuZpyUWCSP0x1sDgkobLzXc6Q68w
eCj00w6UxEhiMpAEzHN5/0UHzZjHVRhc5nScwYg29NW4+fcLBkPvkgmONbBU7fVx
8dIAzRwhRfOReQMD2zMZFrn4KRQRTHjmDhNwgVJ4xcpfApJ0K92O5Wjiv6f4C7Zn
vmpE5GgUy7Os6xrAayFko+HTmWmx3xkXnYqy+E9XowLy8yHpUZVLGAnluVxSFDBw
2+EWDiX5q2R4L2BENYbkuWIfVYD5U9XnJuyXnOn7fLi5S4exU4YYehBMBoE8hIec
Y3Bf5vECSLoK+xDMBYg2TxUzi5czuIZ3oE9I8Z0hemTlFBHMImxdQ4zNXvBq6i+6
yjbzVgqRq7wCJ/CEauijPlWjRz7yK0Yk+IwYGjs9i4+ZgLODlM+dtVrtTei7AK+4
GSjD+7wmQoSNP8lMCnz2NjpZsr6cEysaO/qaw+vA0YrsahXIJvDajngkOVMD8/lK
Kd7yI9BdDJ0P84jqZhMlec8pMZwN9Nuwo+B1C6Pav889vqqtR/3OhUGPWYP5xrlj
GcuRkDteWjgnFnUjTPPAVc+dPXmFJxvHw+7YXLlcMz61WEtu0Uy5YoLnctQhX1qG
VjX9ljsZ3cWmbO4jvRE3UmmcJ17YU97EZJ9lLdAahtOF9XHNSOU1iKdytLNaaoQN
rbLyUfOgQWQ/2Zgx9vUzWY+BPkUq1x/F4de10Mv9CANInXDG5M9BN0fS6FkBQG5K
ogGmMaIz8KMjUrjiTtZx+YPfEunmALyzt+vMvymm27UA+QgE2Hzd7G7cVnTf+Bkg
Unvm+f4OHjdQ35ZdkEGg56JByPy7GDBGJNQnVEbH8xy+lgvgpdtiIuyrkzxz01om
3Zv3dFBGt6CKCxLR5bez6Regj1n+TW0hnsQAl4ND/AITSleXktPp1uC4uj6PcN+/
kgqMXtSF8AxGThHkSqs88jjkL/NM1o4sDvgxcNLM4jf63L0joZyd4RkjyBXVsIcj
Dpa5uNEWYBczsIUStkyw318kqt/lO7qw2Rmuevtd0cQrRbUMOMuJv1i9P6YmvO9n
T3e1R1Kh8tURa07ZLebceY+3m5uDr+g1r1ZaA4D0LCNOSRYwVt/PsbDihe0vIqv8
+rsibk80nc6TCovKpsX5p/RoJBv+5zgKNarMa6EbVQJPSnnS4k1B9q1lFNCqdLR6
p/e0mSYyaaGi6vfhv8NrbYyF/RrnmWPSj9m5M32vBI7ZmhDAGvIIS2x5I54NcQCd
nn//LEmIi8oE5OmVJeyEELbNQP95ewwyIEqUPFUjiTPeWCOVC4kPUrbNfz2sbPyB
luqVsGN0iutz4As3Oi/jnfipxDQnJyFdLyeNnlSIDwcru1O+sluCXqUapsg7wKpM
0a1ewKoW+sDfebx+oD8O6j+GGz4RRRR0F3vzCSinG+mbE2Js6fLQN1F21bN3OmSH
gDlvPuLvvb8xztLmtzrlfKoqqi2hnyld8IBjRSdyVHWGyJ0FGaRzPg0FrLPSE6eI
7lhKEHdculJM6d8YGQt6cbGSARuo6+E0i461RgDWAA5OA9/sW+TVen231SKBc6Vf
yXN3DQSbx+LhPj4FXOv5QIJitB13GsSqy02/LuNUtKRl1zp+Txnor2abY1tyTi4I
XhNEscXM5eab+1ZJ/cr6YUqTmQC2HZUSOSNl1Yv4l+3s8DbpB/6RpTEoX77tUXF4
BgZfelyXocIqsp06RU/Rq+iSphd2F7EkM8l4xHVuFEE4ZnuwfOas16v5cWzWcI1+
wtHNovHua4tdY+MSar4krsfiZWy8+6Lu57MtVyUdMf6HRalQn3lSTjQJNiDQK+eK
pksq1e1TB3kAL4SfYrSZ79V2CO//AZOPAlu5mr01Xc1Gs2JIQKiQSoyItsFLQsZd
jQhb3Kf2DgiyhrgFLAHWOLJv/I3sZK3LudCpKKS9pC5mSUUW6GxasYSu8a5Csfgu
law8zb0qqd3OkyFxG+QO7x5ZAJw4jxwU345CHV4Dkbv9ifodRFL0i+A1kjv4BY6y
rt6JTnco5nR9g0hocWDtbsIkK3rIL7i/yVFCYCATNqr40KFLEfNaqLy2RLLG48AC
2InRMtKiD6nNnT7PzcEM49dyaqOToWOQtdVApKqtO9KdpcvUkgFgBolKVhKlwbIX
4vyrPy7dczY9+osFg9ucR8kuf8afWqkZ+79Dj6Hd8YsnlfM9RlQpqrL5mWo9S7pv
xenImmdLR0VlaGr7GmZQ6LpQtHZz+uL2NEK9nuE3e5IrorgWYK27Bn+1J52zCLPC
y9hKS7QFYIZJTt0in1IpAP+gdM6CUMCbGw9Wy2CLxEE3otom1i2Ri6Bzlio3+qaI
MJh6tnJSr6TlHmI/6+C9lwbjS05HLL/a8MepizHLi7x0itqfzyMIrFGOh8XCpbIm
Cw43TRQS6G1jJFKV4PhyjL7y3+Om9AuUGj0WTDvbtUG1s3ygl2dpthQZV9m2bifO
S2b0uCwN6n8WXlKL+mN7udT9/oiz0IoaZJgmYKH0gyhCVdWeIVoAOuqEXkiflaD9
cEEwygzF4OqnRecU696xIyVAkHwuOL1O2bi2tLRkVLtKExp8VS2f6YTLyZdotLOo
sst35dmltTvnUTbcQBfK69wQShVoxe/8eJB3S1hMSnW6CHRRNVuJho43akCKQNvS
bqUmbMou3aMd4LFk/gMSdosebwm8cCp2P3e8DxZO9LcM3EoA5N392J2mqZrS0Ll0
T97HWGoeN2tK8JA/joYqpfpiyIg7SHSh7O2OaJ0DcS93XMeX6gMI4bakj+BHg436
vR0wl0yOJ5YtXLV3To3xZJC66RPsrkZqFbeuD9r/zxmYzMsbR7kAJlrVg8Axhq3D
8QTTgk5iFrgS8pwbNfqurjJQ4/yjPfHd/OfEqnhC3VG9pgeg/PXAGMw2QOVq5sm7
HHZthhCLN4HkF39qjE7kKCvZRwTes+Pq5SSceWpHRBd1ILJvqx8iREHiTJ8np6JN
2A6zvLlH7/++XSAQx4pfDEvx0h+dtx8MSfPHGFEGnXCL2ktMGUPq7CARlxUkyaif
n03AnjRASuCAAPj/gK2qbP/XsT4yaPpGwE0t+7EUtAondepPUbFU8Ti0Mh7HqrKK
4JeY4ewq4xy+Br86pJHGk17sAPig8Ds8Q3TiNunPvg2l8IxJ3nKmc1PjLkYzU6e6
/K8/vADbm8OO3Hb3MWFK6Sv0bT99k1B9UmUWiWdrGVusr2d7HLBPXVHpGXLMqPgb
HR9BySl5MHrSfXrw/0GzqBCJa7G49tTWHWjbcCrBBiNCZLWprgftihO4eXggkP0E
ZYZv/CXk9gwZPxbkZZ2xQ3bg9lbirWB8vHgVpsgGCYnUr+4NV+HzJdbcFxTkGNFO
MdZURHoGcZGoVY9/eUeCcJUTtIdDh/1qz2+VF/EIX0DDJ7jFN9MNmnvGllF/UzT3
UcUQ1ToR4nbGOe0+FvyNsHZXp/SZBJihvxbGxzXcaIBHL3rRxtgXviEDsUin/c1x
hUM2LF9yqyk94Ri/cDJsu9brtnIQ3nr3114tHi/yURTjIVC5Ku0Tzxgb6l3tRT4R
Vpw98n0VWKWEjrIDzu9T3r3D/pa6yyOD9W/tAcHyY9lhVU13P3aRZKCrcoFhayna
5sKXbTLJ8/W73ez4XnabSSMN8hbsvQkX8l+5AGL2tRZey4W8fyQaLGf8ZIJH0uZe
mYfuGRmhrkB1ayxqCcX/+Pe+RmgXSI9nud46RnabBJsoeeMTesdpWeSf+7EUViNB
AGNJgOSnVqHkbJRPvduTch0R0w6OeeJElBb3VOyIrubyPz89j5EQn28vcxC4YYKJ
SKN6CTUqT/VjD6XPGeOgmLib62uImDm5hBjORBPtKpmcGyTJejLSAEANPW7An3MV
Nb5aJKv2Sb7vxigdCqH/mZsdZuxFU49c+Iehv6/y2TwEy0Rfjx/Vk+dEhNs3bq0I
9xtG3ZfF2BVipl0UsngVO095cCH8dJuKakwn3BOnkWjd0xLnyVRHac1HlQm0Dsou
Lh54ClxJPGkIuDeqRGEzk4bvnjDbyuMCphPmJh1iZlSSq20DhFnFfD+69S38ALPs
Jv3NWQga4/sv6Q8BKwRS2I1SNyEsMUuXFRse4RTVKp6F2uR3YZuzBXLj39mDjKa3
NXl/KNREjqAb1St5ZA1eP3GctMZ7nnUFRszjPB/Nt56aGFeoSzOZzl31/wZbv+Cn
n7bQvnsA6z9tFWlv9VDIO/trs3cUKia/LL7rloi2euGqukll4+/aS42BVDJ2z2+T
YaSdwEgDpKgH1i4QRkLSz3qxMmWJPbdq/f2lhhVic/ZE4kycBgkyMFcPm93Oj8Tp
rzCdWi+RyVVTJxOrzB5/5DQ60PBABe/55WJaD9HvaCybKPpbCLsqZTBiYT8GJeA0
wd1IoHro14Cslba5VcRhD/7yqjH1dqYUJRhwuRzYAlCcWnkRWyasDlfwpp54AzT4
oq44WFfq1DWI98R5J/c+kCWUBdsksxM7RRLvEETEKh7dnF9dLSHzVqcaREf8Qzz2
k+nuCz2wR5li5cfASm+3unJIh5qVoao8buAKoeWMGraEMEMBUdt4FAkK19FLq+pp
eulkZHP18xpHlk3VJyf491FaZeqO4cbcrCRMymZqtySvyAx6GDUdkYHbud4xYI3+
Ups9N1IZaV43CaLZFNEiKmLuzdPswfbJ+bAyqMVHKKRcjVLR26F8ZNO7rLKb70D2
yl12ajordONAdnxVNdOK4NzpmkFohTt6JOGeiS90sA8o7nlXb9rhZNGqW+oa6P9v
rD1S07aa9IHvG/kLPIfryYd8HOOf/KbethSI7ISmZtQ1FZv2YVA8ggjH/6GGTk8h
403wvdpM56Nc7EGjx2aR7SSdb08HtAhK+NOLRV7zorKqyjdK6FhuuLNverEdcuJO
WW6HdU0s2CPwzjfGo5j8CChxgmbQSO89hyGIPQpr67CGjUI6NHj//qFfQjRnekO1
lhT+8Nz+/vjggm9q6Rn8xzjHOgcCSpYfw0socqF7sRLXRbZ+HNy1plqfF5uVBotL
mCOtDvx2y8dRe12oARiOuxUMy1GiRqsfkpC/RDqVd+nxusKwF6pN7shqjqfUG4M0
fahnkscjcyXg0GAHv2Z2XGSo1veHje2+PFt5R87e+afaMl787C6klPXFXrVIXIW7
LVz3+lE+F00gj5y2TbfnLAyAYZK6LeiSyBy3vkVIuuks/XPJRTLzgW/TXpe0Gr2x
t7bU0hHPm9XdzCYKfENutdSBkk2ED18da9X1rcJvDt4i+OnsbfMuia3ujwZ6Vl1n
2ax7L9T3M7F4CPYsG68PZPSJ+1ivGkYSxVxDo++u1uokWBklz//EHrlidimf4Df8
9hhtatrkz33pmqlBPtaqHAKcmJ/BsDV0EMQx3aEcTKhYSZAudOXvhUMIgL7xYLzZ
KYkeyFuIrHnSmJ4w2nsDOhr0IW/Ua5JzAHzKGSRX7yMrP5BgBBQ4a8ym275Fd84k
++v+7tZvs3/8v0ivwbn/PgRI5euYoDMeDhmeH1gTMla0C50CAD6fK121NNUSoi8v
jU3m2Eh1DpyOrFxO2JVbmzRkxYDqURvhZHvuRhWnKdaRvXaOiUIaKLHN/hEDrFq8
MkTjHWxk0KDgW5iIWO5beD2rPsMCSTcpbs+GGJp7e+N5FJPIBy5cd3KV6BWkjlRq
We9LtYZp7OYqTi1oxfF8gIAYsM+hfudgxWukUGLjsH55bh231kBDAqMkzgiql9Yf
0rE58flG2AXjIpU1130a6A1qeBY94mYjT/aNqcR4UAwvOb3nM5k+i6IjOOwGGJje
g4h++PKqas3kZviVvVu6gAZpemsUQOc+ykckUYP9amc9OBzrmbuvHtnJKPcD2xU1
Z09yMlgf/uTFU+rzHK1kmFB+0geZ2RvbyOwd6owk5DuBRl7ISlKr+p4GdUH1B2Iq
Jvh3Lv4/teqhc/vJz3N7kqZG4DCz0ihfx8YTX0QPvdHJLhZ8LWqPZsZppPZTQPZA
AKjvTGvmSTQYU9/Hd1jlMD2+BvQmV7+Aa5jcLd6INHmW07GtEhPyX5UD+s5aoQTq
tJgqaJnscMT6SXQ4XrGA7HJX0RGdONjYNc+sQNOp4a1Qi5ix77jWVrnzf1fiPsZ4
4n5nyFt0pwB93lwPK3FJoRmNE4eL41kDYodzODkzdc0PfVX7zQw0nzid768EWeHN
g8unB3vs9gJJwwWdx8EG9rOgF728IVwOjZXelKK9tMDA469d9pgUXD1GdJi7PFmY
Wdw/bMPyJXGZZOdkxPym80Bipa3lOr60qU87DVuHKon9IYfzaSVCE0BD8vvImwbg
k045dMWy8GTwoqeFqa+8uVhMl1VZsVFKRYh+YArDotFrCMZhsYrAbcYzedITandv
0qUCd4SSdOm1rQc48G3sdh5Jzxj7HhT8EDULLHu+6EUa/NQ150yuBxMYruTyLY0U
kD6ccvcNkvWm3uMay+8xhqSi9gtEyebnJdcgfQr5Upw0MCP/BqS+7Tr9O/VEWGzq
qmkk7Bea/rfJyqgHPwzNTmMwqdWu+V8GoabMIt14qgbAqtLuMPon24Wh0vA6mGZd
f5sdIPjsus0ANvPpaT8aheSyea+IodBNap5UUXm5VGgEuzlCOZBQ6YkTTD6lma4i
OE3lCWfqpWXQndZr/KDkj1zkg4AFLURjzekKF9EJzkpc50BhYDhGAZy4hXhiyHBp
vYnywzfXpzzHalke5h4+CxLcW3RNFKdXhxcBGdLKds0dW04xqoShTNzx0RIvr92o
SBdRgZNgzhLxyDYPzzqKt902m4t6gLAkbRqdHT5CiyFG9FmcuTiAmhcVmj0bXDZr
zrfv1MxI7giQojNrnJCFqNSfJa6WXHjFNMzc0YvQyPAyO9Tx72n8Iq7h1oDoyvrO
KRTzWQyJZktkB4SAcVVBJjfaGvHXMOu5pHFvVQ8PXBJiRnvt6uUK64/d/HONPjmq
5CnLThheQ4aVvsWj7RC/F62o7IL2vUFpjGI4JYHM67LQc5L63hHmTKvDve0zkGCE
yJfII8PZWMtZnOnfV0Uxgg/wACQ7IFkFN1c4T9ma+mQgK5zb3QIsKoFNHZ7DJV7j
m8z6sP7TDUC6RBNkBrsHoQ22K/HqnkR7lQTMZKNH9//kxtG9Y/v9H+bshHm7zcQn
/T/FfAyueSYcB+bCxCskX0fohrawvC0gvuPAjrfyr+vh5lISi4+FrYXeV1FpqvSl
knlgD5/+zvvpDvWJ9HFax+q1B/LaD6Wb+tWnA61/BZ1BGv6a3cZ990SaeFs4qwZ2
5joAVykvJ2qMDdlhD5eKL5ebTwj9vow7eAZMYB+nzP1NkCMedoLMB/yEpdzrU/TK
oyttxoC86ywzN9xW8bZ3CmXZaWMVFRWTgjo1ykweV7kUe9ERcZdEamNa740Fxv4h
WAemrLlkKf9ANf2Tvb+cfo8L5CK0N95mrfcCCG64ACIJSg0+MbXWRI2gwFcdPZ+8
YGxnc/RUFilJv2r7M67C5ClWbtiYdz6XM2vOiNQxlyweP0EEfNXVZV4sYdSMm2E5
x9EhV4Kp8FpLXNIKxhd2BZRoxhn0FVlJkjXEQeZ22PfJmAUZtSdyd9adwzWFAzFw
G3LTA1VM/rBUWNHoSIAzj95PuFDUK90PqkvN9UkKeWoM3Eab4K1qPkaw5kTMZ+s9
ujRp2VA3uEzdNuiCPbh8XCUjdSNqOSVooT2iBu7LA2BX5fej5wkUK/VT+HF5hfNf
PLs+/whsd9QKrY+W1WtEsoUVixazC091WirW/ebGy6uyVUKWR3n7+VskMH+K7Nm0
ECtNhTcymcmRKXsMksZqzYDBGycBbgzFYmGdmjWDx/qHrWGlPHsEoZaCtvq282N3
3+h4rSetDnofGrorAiLmhONC2f3IuRJ+763zazoCeAwhWgReCryIT8KNbHvlFW7b
soF9ffUvkCaSsxkBABwjlBFBkX7Xe3qOWui5fYXQeMbjyzecc16ENjl9vO3ogGW/
cY2XCcDAiBrocnPDGPDat8Oa/OGWsZzz2PNCX8zrPhCYkr/9vwdyZGA4+Fxdbdlt
TvdIPzoyG7B9Fz80mq2JP22eXIhM5W7QaqRazyqi6Yz7Gaw4OtJy2y2cSrztlEQX
Wj7Yx4+1Wa3XiYULV8//q5lNnMhai3xl8xbt9Mxl4W8jTGcrYJzBgDbEh4ZaGN28
JBiL0f2OD8j/1HkERM3JF/89GVAiWCB0cSFIz2Q3JmN528I6SnY7r3tXuOAunpRX
IDvzAeEfYz+sjzda88o+YJha2S8nAYf8aBCWlbQmd1xHETtieCUOS8AujJXtXkwr
aeUFPCx2r4aCO64xPk2IoYVkKbIE9fD9vDQf4qnKAD42KmXcke5ySSfZfe9S3+Fp
4qF1K88JK88pQEszbi+F3vHJX4RwCtgUeMe9hRsnWDm8YwrQ9lqH4GUhhBRkQRpX
Bak5jwHb97fh4Nfy5zAS6QFJ4M4gZNKYO05l+KsRjyX1mIFKzG7t3PgaH4wDNyHD
yIK5K9QwaLHgaCF3dOCqo09UKgzw9tJQuVvAqJ7XyW19AOSjpItgyieNPEUGjChx
+u2aVc1PN2tI0AnS7vaAV5OWq18ZKhTexWoFPcpKHyduZ5wtlLL8D9b21CTJ/2/+
UbNqoC+xs8uvb2L2y1WzZIyUXhnKO5mjIxn6bILgEhvZHeYw4bPag4e+U0JTUiOH
J63YASdbi1ACxbwdRTkYePF6/Id86lvswueUIVHMu010tQ0O/+LyPZgxOtdgAxXs
yRJavTrKGoqVjOLMXWg0ygp0L9/r5nA4cH5N6Lq6RFsD93aMVTiKn/Ek1fb4mDXt
VPzb9znehmhFeWwFi88l5Lp1vBF2GY98cE6BUdF3rDyVnIzW4LliXlxXHX1FYc2L
JN/Y6bOzM02HJqLw+DI9PCoiCFLrh3ii7c17iUQfkZDDihw11y+QcBC6HuNe9MQ9
FVHEF1FS+RGfxw8ogB5oVfYWgCUwvUnn9pOcvfG+8nYzrV0Bn86wtS2v0WC0zPs/
fM0ESd+pZYwaD2w4i9t2hcklSDxj2hno6QBIbKowl4wdYQCL+RMasjBduvi4MTMX
tONvwyRTEoYRNa72O0445QAngh1eIC4klCXY1m3v4ikGH0F+FXBcTvXjRojMDEF4
nZIjPV+tGOUTYtr3siSMW0kxUDLB7NbDNfpmPXb3o+93NXlL4DPRVysDjmypdPOr
KI83z0zYeQ/m8w3S+wvuSsmLH8pR3TZ/UFraqm1mcYFh0/wHX1wEOMUC7L7jF5v6
/JfrptXYUturiWlPCGxw9Wl4na1+qK6ROFHTigBxyzb/5UGXw7yIa2g7oXa7Tw2o
U72U2vpp1Wf8GRdXxJWV9Ukhop/4VPdAGs8G47wMniXfJCcG98HvukErpkeb7HAP
ybvlCn5/0j4Lhn+3KHkjFH5/CY/lzT6w+druQktiKmlIxma8f71SnQZv/aVwCbKO
85jTPnM6w2FCucZKeiZQqDpPlJYc1oa8xWtvsqchOj0H2OqerDzmxzlMZ/Do2a1G
CwQ1reKAlpMKydsUlISnyOq/YddW6J2BPpiniFHDjdPcF3m/s3z0UTWEMbs9l+t1
ZWeB4NBI6rn5bCBOWoG/k/MzluDePaGgKBbaz6eElX3v5Ck45iFX/cNje9ui4EZE
b/b+rBVHAxLm7uqYSmK+/qrfxNmbWsADUrrrJFDUmhNffRaqeiOO+B6LtVJSHE1m
EY3oAoKgw7f1W41ZHoGsSpyw+RljKgmHdWfb6i2Jc66mjV3/on7eOi18rdGe1gYJ
OA4bpm+NT/mjYtMvNlSjsZieIa06lru/EeALVvKf39GJLxD8i9up661CsDCaNLmy
T6cZZ27RNj2rMl9n/mB2iSvawXMU12Hk956XNsjs1CJ3ywYccF5pAT2zugYO/6Bf
icSwCGo6IW3CzPq97lgtwuxNMQErA9d1BddqKkKgjZH6kpRnavSmC1/qWe7beg3G
gvzy++7E5HlEy8oNZzVBpzV1fsjb2GEdcutTSF2zG/lKoqAksH5SWxYb0R6pfyGK
qGi3/93LJqdopsMrnUdIyYHzJgqMtxoCxHD+vCrnSEmmzSBkGS7EPcJixXmYzmfy
CZhBAQGCkMT55R8dfT/LkQyAFDW3rd0ppk9rcI9FlD8EXNXM/n6AUg0U5qBb6Fv4
HP9I5oGKu2xyUu7Rn5z6SegooE1t6yqmmmVJo6FGh9Aw/nukBl5q271Nz4PRMk9T
rs7cxZ0JmCkts3v80E7vkHiVoaS6Z/kdFDY1wnVQJbEjtvaVD7p21/Vm61c8aUVt
cX84kj0YdMnLvktL04Q/grL0OaOag1MTdn4y9GV712aD6LaVgAaC0FMt91MLeGQ3
WVgGUegZAARsjtAubYygNh73wuEILfQZO6krv7iC/6ieU/VKST0g3gcpAfsD/JCA
GT+zzzEchpvIiZE6HpoO/Qj1vrUAzVA5CdxpUb21KUenFTzjMupvw/30XObtsstx
e+KGU85fFtAOK8oUu7r08OVWUlk1yuZErQQTgyK21V7Uh97oOWClEDFw3Pyj5JL6
7gVH3okR0qWY1W5bBmTbuqmrnKIbi3BkkC2ng0ZhXnbBqDDNow5Z9q4cHqkD89U6
hHIR7EsmWC0sx5VhQMITQ94IIp66dBuaTeCCWpTgBBfMbA8MuOVneDP65SXpJUpm
1LTQG25GAXG/g5FS1yGSK4VUgUY4txyQ/qgkWR0yMo/qhZ2sSZ4ZROO3eZD+EAWn
0osN02v/jgejVxII7w2hEUQ7W//Emt9NCJWkeo3beGVJec8h2OcA42T/i3lq51BD
djSdUslvLvSH6iphs92SlQBNeqsa+z3qNeqBOpDiF/xA+J59ihelFQ+JjptoSM7L
Dcu0p0c7HDF12NEq1I51/mTKSRBF+qXeRXmkr9cULNlxATmM3fS372a24+sqms/m
Y9Tq+MK+dmkhCPkKjtp/iJAEA5eJNzF4OGcUNhhBOfvlrIEArQ5cyJHhqbPJEmRQ
pslMCU9rzWosfNzdNsf0Ig4wMayi16vCYmcAyQwgMI4Jmbs4q6nIGvDxLIXNZP0+
fznfwOgPbsZX7hZBDjdxJH4vXumoVdktH9k2tMkk/CFOzrkY5YJ89+260vT+C3Z2
peAki6MB1zDclqnhJv2XqsFSlMX8no09R99l0VvCYQbgBnO0egKXyOtccEZKiwxw
gU5CvMm7RpIUemcxhNEvalqOZXE+FYaJ6AHHhcDh9AQ06/0/fZmgDaZVp8BdBxJg
cawJDKRbhweebBXfa+YK+h88LwhH4QCbh8jxnqxqwaaM+KVM5jmbMreyJuiXB0fQ
hs2o3FHpsb3oDIUTezY/oX0Ko2yuWXQsgPqpuf3n3uj+mfADda3p6YCyATKe2zP+
hceFLDBw3+uHE+gv7MOwIOVZ9aT7fW56dezCz0A+iRerWJNIN4RwtQwAUvZu1hqM
hDv33cln3tng0xjK2UZrTnG71MWwCi0KoxKr8AZMssqk3C5iarab6HH/hJR9R3N/
zXwg5aXn1P8bpsX4QtcKuLko9uWOKbM/5GX8/3v+PitlfIuxElATwahNMz/XDrHR
tnDcIRsliraPKwuJqiZe8NGXHaXwVy3qJo/Ai5h29UXc/8P+RRIz3vq5s/P3WLU/
d7BuC36pRF8u/mweGKbV6Gm+8ZbT8Ac3/xXhMt7ha7xZSRykmhKjIAfFGdJcAFsX
JDmyI5BqZzYghrJvU1JVJQXzN/nU21GDE6aMTwVruhRd/SDrXdOGJdLAxMM4yVUO
xjazkltTfeC70nl63MOJx1Ylv+5W0DFgSmipleC7gReVhfWiHGsZnh7FVgWnx818
EmA0OtjhVzFpplLMfL2TqGDiAUsA2ENd9FcHjVVTTxcik/7CrAhT76PQPvBa0SIH
78/cWlDG/hGdWHsThGP/0iB2nJwI1x2fztiIW6IoqpIkZKVsTPfLAiMsT14tuwQx
keCyKPc/m1zlzV0XgQm2wTmarQeySaDjnZfdNFUt8G//jJAs7Tsbiz88YuQSlPgs
U3FC0dW76feP1TSkpujVDQaUzPzEgpdr/v0KQ9Q4JVHlqvA/5K9HECbmiGh+aq9o
yknpa5+wgjUCSC6ogc8qdkXT00O0NgGZb6wUzRICRsN0FuqZQpG3dnnVh20tRi5O
lklTmIBa/+ON86OoQK6micH69J0glTHyj7vE+9/VRd5RSiw/iOm0CLppCyOCemHd
0JaSD3s0DcwLoV7eoiHjUYduo49cJVTQ+i3ZwgioQtAwhUdkzrEw5I8NQ0SD3hfR
rBtyYJj7i5uMCmPEpbUeumbdYwHSKJlkpe4CVf/hrKmEiFFINnbHWTzGZIm6H4Dp
mKUWWBm7VrK8+2VuoaYNrusDf/gNXlSq1zzGKtszB94jZX9j9tBb07FiD/AgQZIy
SpREHbTZrm+we8fwKPexzGleMi2lXWelc3kEDDbRzi7UEeE5GvEJVz1AdLzSjpnz
AeWpVWxH3lW3I1fOaqopURcloQjOkpY15nMAXYmAekdSjrBlmoBSHHqMpxzgTF3C
uGUL898pw0HVmZ65jOAhY7CKkZ8Yy47Veq3f39uyeH1dTMYViYOuE+6QIeAa6gjd
UUi17NAkGJSyU2AZj973cvYZu0z+mtGDSC5xKhfYxPHTTvGd/FExr9j0+JLMpNJJ
NP/XDnw0J58d+4kLctJgA8z+u0fZNkmg+1um6Xm3R4j0XvPjttc6FRweUit7fDOo
tqE9CO+VbMDrim9tehVTkjRntAn7YPQu9xSHvQtCuyDwzDJf73YrcfxdXL75K0tj
J+u1ZaIGsd7bbSsVrBakNQ+8SLIcXQ/9nhPzJYYv1QxHGKe17Z+S8IyVLynaGlkC
d2bN3uK6OxXULb/IYJt+iz6MHisITAd168gJwa41y8E8jIzEAiZcv/aWLMa6aeCW
VmOs4a5LFn8+nM8donjLXQrSNDem/nqM8o/r8jRa1Gq3RPonEIjLF05UebYq9dHH
7rSS8IHiDX6oLc5lNw53WRoqTC4frpPd9FKTaQPquBxYdm6yocO8eBKAi0SWccuF
ydm1f2UTceOhNaTQzxER2VvjQHA2jJDonvqMfSwnHacXtdGP3La2ZbQnswG4RpC8
5KCzaObpX4xnDZ1O7zcDbMVoDuy49R3GfFgbiiHFxRkFRl9BUowomF55BJTf5ZHM
ihHoeyvVnxuK+g/hGJbFsw6uHCdN0EBDv2JPe8Cek2m4fOfb5hhrxbKjFlwccqdS
kiLrJapcVJi/kXF+yGTU8JWwjtjnMIKXIObA0pCRmD/asbSH+tsazRZvtBBALbei
RvyANdgoq1m8XhU/Cduv+drW31L1mvvORXaNFxhYBasw+YEp6YijvuN3WKWELDRu
Y7q0dUXSrP5x7W2DsdXCdF2wPJgVRxbv7xR7QWhZ/wA37laQy/CTvvlgrr2t10oZ
lbmmbyVHVzfUt/5cpjEd3sGu6harauD3KkJOh14FRh60KrpKyLzqBf4nrfhsly3K
6hMxqT3jUEpNxZGdLv8SDUPzIdqgUI1gRQFFrOBMYMHITQbGUieWPWnGbCCtrhVv
UK473CEmGvxNxnGMwgg4AE3dseIUkM2t3DYxpmDaF1EhndFnhZTVeiWqwx3flzSL
2JdpfYdTcjkmLEvwC223drhkJk9MuJseBtVyAiXhkxzY76u8qnH+D0O7qsPwl7KS
5DxCJSKSGIgcIY2uoURewXr20YeatGfGCdayykvk3pN7RfyBrov7cRm9uv9THSIq
NSedygIu2kWgHzmR1XSUqdW7pb/jVb5MJ68A+rumDG5pG727/48aY2sv6AC92+VJ
NeqLuRvKgVcuH3m2JNn/BN0A9O2D53Yoa763Iay59gZycWmSxrGZDxeOM5rPwcoj
BYLW9VE7mRIG59lZ6vOAIhDNpjrqfniiR0z+YXG72qvNck3SVeck62qaBWXqK8xH
qptFVenrjA6jfdFjH5Y+sA+FilWuSihhWGR7k5ys9Z+l6N2HH1tiVKtc0gOC2Evn
njvuxmAUbPadShdyXpfK7tf6PF/55m1hu/GerMMy3UEgrlZmq/kU6K3UDGgsj2Hy
nAMQZ7187MVnuEyCMXfMY6N2S0ZePAjWCAeWexQTbgj3kRvhA81Z61bGDfBwiiFL
l6Jdbp5DHsB1m54rXbae3F73mvayzUfrrzaSVNncsvHOXMictK7gvgYKaiZx9bAI
QREQC9mpp8gXV6eK0k0ZvBoDHRE4L67no4TyrwITibBFxNOlDAupmcf7SRMdDKmR
OSlOJh4dfYsMge0+XBxY+tWlXrKAF8zHtg3FE86lBYpZDEM8tjW9tu7kbbPoFaRp
ad3OONv3K4+hjeWIKZ91n5AQXFhD9RLnHC8qggQUbrkUtKyYT5x7Df2ytnzcF4ND
fkdVwHJM9DVTMBcQC6lRHJruZNdPwlnDTc3BnkFEe/5Lh3fTQlGUmsn394QfnL2I
OiJ+qGhgY6J1p0Z4v/bh+6+TvGYKHG/uav6dlGgdXhwWE/PcTdmyRZyEUf/+PxD2
Kj/Oot8cIGkkscs046MN4HgJZMtfgDqszSPnYw4ozUxLG+spff163HF1kwUPpT+Y
9DaGxS+8kiLfh3xeMb4LDPZM7JiNN0D2NnLX9kFXtlaYwcAJ+OaSDWNBfbFYNdUM
2YB3IBYElX0m0kjIbZUmY3Ct0HJu8D8/Ut5HKD6YTEiqoJqkh+fI6zQVdJwbDXwf
tCz5WXfB8on29habz8e/nS3FerHHO2o73ssqcI4BezFb33iOhC+GeglmD2+zTyxN
9qP/lmdRbCRZCfYZsOYB6eENP9sZJYAs0yigLcAlor9WhB9/8+ertYXXbo9/KsEt
SNfu18VY28sxKe/Lv9CPxtmJjhmQQiMppSJ9NWG67tMOukNDVQr0RdfNWRlelfYR
AFr6ajo2HF1WAMg40D4wYx1Ga1AlJnb4mTezz9vpQuHuwdOMyixeGktmssxNfsD5
oDAkfEkZEGzEzTOWT4vP2VPDCUJf+h2DFpWDSYEkGtHwFakfKrUuDb9YJ1sIgE8N
OUU7/8UhdRFMvFLItJ07R88p14Mu4wXsIJZJ2tG0XW5T2JIH1HA5vffdYyAASHqO
rnwuhwXRH9RisAeEV2SWqXoIY9EVY+XYNZhj/Hu2ads2y/O4OgWxHMZcErnAhkn3
Cnboo0NLDShNfw9NqOsrDgnVMMLu2CnArf49HzqFymzDYe9B1o4PAOLVRohZF5KU
JMHvD8En56dxu/3S6Bl21b2tTOVkJAbNxfOsxuo13OfOr8meGtcTpO9f1lrSHQAX
Ng/qsI04kYLM08J32G2cBLU8GFPKo4c7YOX7xcC6yBD6vJvtSyH/LtLhHQ0EKc15
KJlPYlkq3PnG1SbOTPWzKFvdL5o/SPcFwFJqhQPMyxd5yzM0G7wXPsOIVtxklhkh
LstjeB3xsb0YeiMWelnRxZLqmcCuiKqUGDHXQD9qy21s8bZ38iYjgOePtzcW9d9l
EAyhDxYf2R74fnhVm1p/yrj7bHbuJ6+vIO8bdzghvjwSXUJxH6J6flniirPv5u6L
a0tYXeO0mHAKwCFeK0dJvE4JC9eLFNqPzyJa6U1NvdUJ8vChGIYxqFPmNxF9a5z9
xl401fL89EhS4YUPNEHGiFCPd960/YlJLBq8BgFhdJFag0ynyREcW1ZcBxb3+tXi
TuxQjvgvciPXC9kBDYQRleJUT3MaPEPFBvZ3IriyyB039KIxdgoyynYiw4LYBvlo
3HqMAS9hF+sP5F2BcToNh5TsPm8xlrLd9EUncl7NALH8YUp/EJda9Z7C1RQpywd8
jx/WkszRfTrfc6IHVTfb7AP6BVr6xf6zp3gtczOC7d61Ni8d2433S7udA5hDstSO
y3l2/QTdOu0GMyibmV1efiEuzims57/tDDpwFdpgjRE6zA/220YrPEB9R1LUnvgC
G3t0jJsefBS7oV544/4KBVlg3dhMT4069vPKtBq/LZulIKyNbhm2NhNMrWDCineO
6g5zkVOJwQbiOmxEaGAUGQA3HkE8rYpXZxM+VFvJyxezPz0mcTrQAqgN+sV3mMhp
aq/wjOeNHhn+TamvJT9BYDsYcbHbQvqjlykO89DKcSNOeJasu24XgZsqWw6jd+Zr
mmTUTOEVIkDxCzRJ4zR1NCy3mnhVwvPn5ogm4kwHBnk1paoiRcMOTkaX8uwb23bX
D7T+fhkrlLoy7KniDbIgPJVO3zHcLHTwS8hVdKAfBwEPm5HDaWEVw3LsInqstFDW
7Pfbzojuee1t8IZiDzOH9lG+2jp/URtpbECdVaGCrFJaHLLRxZSsOpiBl5IqNmu9
WoOZAEB/J2G5R/Vjohvgyh1w9k7tNY3b5MAZtTlgkRBcAGRJAg7qRAn1Du6TmE4R
Oxfq4eQJfNzBYmvmjBHTT2sfYq29+Xj4bQbrieLVGMonZsBJpA5hd0UaDnrz9rYq
urbwWvadSZ/Fyuem/ijLmKbZ5lMPuRBKZKh2du121brXKeF5Lik5LnqHtDc3mQwp
ctEwc6Ya5/FjwuXJTJZO9b3Cb9GflF2vzyIWZReE7h9SpMkUB2wYoRjbrDyT8f3j
heySX0k5phdSbUkM21QSsT6UDmUbeyNdHM0sPdOayJ7tjcCBu/MGrAMiImfb5rWe
tE5MPoU0ZrsJr/aYcliVJfA8uf2rcY0V/7Es2LwP+3LQgjmEQVufupqcs73HyTUj
ScF960uBiZ5/zUL5VLtmxp71WKpUjtI6GR/D9FDMIynVE3HwadRqcL8JK3vtlgoe
MzZFpfpZ07OpQl9eP7TB8wJ4DzpmgBicx8JnNYBjULF0od+u/snk5pHoCEyML8ax
0jAeqO4PVp4e2fp2SqGloSLf0pSaTuR7sHPNb6aIJR8ZkXof80Dt1G3NgfSz44k6
hmIy0AV7lHu2C2xUEGvCLLLGEdqPES7w0zeNEP8AfCWs2ZNnHzWsoZ1PRQYYLgSP
CvRT7F/I9dRwBq/OOgw0N1MlfecUi6tWQOLeSJrIOEhVmwwpWrzYUzCVRUiFxz9k
bnjr90d9+hla3LhGsDp6vnu+jOFTp6/bHfnzYw7vkUpNkTkes6KlRi8gl8kVa8wG
gRJ+UkWL8C9R/BZyEHiGsfvK+gukFnZLTExTizkVwV5DUkNHp5R+ZWcVvw/gwNkZ
YlZXEriKkVfm4u7bnVvQjBMWu/t3pLl09MCYvPwE1X3lTwCj18G92ZprJ1PK6aWo
kIUHHf871sJ78qI6qO5fTWmkcSN8Rx43sQoVXvDhFNEkiE3s1XkC3M/cAXJFGw2A
OKA2ntyXmO+JBac0SZm4m5pf/1EgyzV9dFpdT7rtn4JFLrHOBp1pbVNPnOmTw3ke
czq+Or/WglWcmPPMR7JEkq/kJzPjosKEoez7MIQ4er/W1P7rF4dWqBFN9OI7M9Gi
ybAFOvYKQqYzXoOxzGMOJUIaDPhF1JH3y31KJi4avzzkHh+pO8lRKNVQnkJvtFWz
F8ZuhinGYUM29P4FApgwt7QIras6e/eG0k/CR3az7xUqAOKE5slqLKfCiLdW5PMi
9r3NGerNBrA759IYUqD3NY8nzCjOFKTe3t6LInC4aMvo7J78TQx5xovQFa+v67N1
RMncTONYE3GTPf2+bfzpi4eCTHhqEcWpFlL+tCQJFgTtaPFHHi3TLAelZY9JaYXb
CDARTfzMWaMhwBzHjY5o3Wo/nQwDOgtVJLUc4TBQ+faHsG36Ova/IvO4x+iAEQPA
oA+ke0fZqRUwWQzv3IxXXahOMxgv+8YyfdXaDwwSrkh54U9wpePk348PBvk4dS5E
z0Q0zEYHyCA9lwSJH9S3/L8QJve1HEm7uvzsMsUgr9tlST9hn7bGfMiCNLinRt5C
/rXaGVajWoBRgIOTdB6Z5+Yspu/bYOUZ6ANuy7QUnUr0RmWFpqghuyAjYlvixdFo
BowGYN3C20EXUSOMxqwnOEBwabwreropTUAEOD+Nyh1wrJOr0VRKoqx75jDIWnhl
v6SBAnmctphv25U+h5GALqwJpGOAwVuI7PynC9UC2FmlVAGmSCYovevviUiA8brk
SvBjbInQfwYLTayIn2QGqUan0pH1i8c/tVIkq/y2zXYWHE4nT+zj1zhRT4kNU1rY
B4npOrmtsNjZxaZ2MjJewWSL+bevdcka7USEFMk57n4uc4Ku5eeiQo9qRRtUyBOj
yxeN1a3MxDJbupf58sQbwPMVNEPD/mv9heV2e6D43zwjA3v0A5WFtpVoTSgJRMaQ
ILXVPVT9qLqe2HNLyWCG+3cLsh0F4P23D6UB58Y5WMOsecyzTXSxcybDtR3pSDxV
rp31SzkH++JiE3/ngpcsA3Id1pGlnptI2enFtkmD5U33G/uo+03qpIRgwUx6u1QT
+NNxx7APuNjZxQ0ZiXWZA2+SCNatdYPtaMviqNYhZjr1iXV4E3fYmaJtSN4brv41
AEm04cJ8CFs1yWPJtes+2SodIRAwA8Xi0pyePqHL2f+3iO1ve+e3gEsZGljUieF3
JTSmUR0skTOSPauCLn0LTHsWuTa/BSw8UbwekDhpZMVbWdwtfV24nDjvS6EedtHk
Oi9apwlR+p39fdB73AwxGIT/KH6dd2d1/AJru8sUyOy5lT5U6KhviDn8yQnEZcPM
vdH8OlkoU/tZB17glw5OpHp8clxTnVA4WvY8SYe38LhRgSYHgHM4xK4uyTLlZm/A
ncm4fpxuGB2uWz6lEWY+OEvqqnNXQeeLE965KSauEbUKS2CjM6Whhl8due9x3dYO
6xX7w8qfVXuzedfZFsf3jdn9+/gZ1GN3eKnhzPpx4abgVLbcfD27sD2XkNeP8LH5
c5fgrwJQyD+19U0S/Z5yt47CKtSiw0zivfyIAS17egZ7iHuMboMgcKxWkzxxUtPm
MgWNmh503It/7RZjbP3RrJx2v7F7eRtFhNkZ0Gggp1trphYPUm5CpuUv5fJPE6F4
6LjwOgLrRRVCRYKQPChOwJhK5kLenLqk97HEANnAISp5j3aIxxdXFhXWPXBroyeK
AMP+lYzh6c/55TB+dR6J5Lw64iQ9nAdaIDE1XsSp6BReemw5tZM8zVN17XP6bOrL
fVfOjcIoHz3mRLN+2rofvkpMGbr/BOGuDIHYYerRl2eASI3EbDybCl8CL/r9ZOWo
xnsoSoQsGZl5e4uod/GhitxNA2q8EgCv6QIinVpX5xbnSmdvdhGMgeOp7nbP6uk3
qVFIFP8FDF3BPEoV2aofASoKnTdl2Y0gv0tWQMNsgKDhRfbHiI4T7H3DKdVMJdSQ
sZMZWDFG8KTYDMG2ca44iJgRA43VsWKC2xK1AmqOhJT76/v7HSZc9yqhC3a6102v
c+GklsORuofmaHlSq9niIC1XShHkcDlxAfgIeIpv3b6Xsjo8VT9MZHNeaXSRLTG5
L2x1gausa6VxElCesxaAPKOoZv8OCSakB4XfBppnQFU4by97tltL47+okDZLOaXH
NIoayhdy6dIqKDj929dkrB/QHSc8qHECuFzBI781c6ZapOERffJx3UgmchheJ5XX
ki+ZhA+0GnySWoiQR6X3BLIg0cQt3tE8ffz441HQDAZ0Su9sefSGEFOtTgNhwKT8
fIUCbwEscwe9q3at/PXw24CC5fVM3N9dtokePk0DP+FZkSVP9XMUy15V/ReosNuG
r9kSpqlPHNzCuEZH2haEeQO2VnW9LQQvBz6NgRh67HpszX81Of1m3qQ5y6m7Iplh
327LCD1SxEaX5peio3n7NasRRoRv4gEkH7CdvfAM3S89M8SEwjigfyNK0seIBO3w
OlsSX1lzC9QJdpCC3HGX4wz2XjyEGU3Htywce8pvshEii9lDmE3xO8xP0yMIxThn
Ae0jZ2bFHND8DS4XN/H4hNBzGNCK510L1DEdhPdAtlRSuFLpLjijuabpLtz8T6HU
5gXEq/D/v/u2E+XjZYrT2/kV8L1j6ZiIZ9ll9jJYrpdy73ejUKO3Gsw0WccdwD+M
pW+RrTyC7xmWdF9VrvAW5RFVWJUHZXw405KY+NZPOjVN1wYgYubkytzN/aYlbhbR
MoLeAQPT4uyVhOp00H7k2Zo51xpiuIkmksM9udYxpJHugOmIzjJXhb1/9jtLzW+a
QrKW5BHoa3l5FZrsqT1uZVYhITHAaRR7pw9IA0BDt/7yGzUo2t/RF+Oz0A9D761T
ygsf9CadiL678j+Jof5igJO+OUzkCHQXbsEnYj+RrDJHJPfohR1BxVcxYYZArw9k
ghcvkSB5O81eUiHcX46mNgbXnm2adt1EuP2izciMizp8ZZ5UAOr+wW06DIJzn37C
jmhewuOQiY9RU254PLi2g6AS9fqX982+IdvVpDW7X1ufaOTSNFqwVmuepjpFncWM
IJxRxhXYWxQRBcZeFxtUP+rySr46/e3UV+BaoXbpJztOgkYfZ6p4CopD82BeaRKP
fJC23jgoXsLC1qEkjpFXti8TgK6L1Ouyj/qivJbFQ3MgAScc4ugBwHm0G6qtrQSm
vIvYC7iHI79x24mChpq06J0pXOC+nY31qBqacwrpAqiYUy4mE8sQ8/66fWniHMit
xwyCzR/clgCf+Vd1r9HgFIeDQGYsjfkz+SgASsIAJ8H8CdN9hKMhBy3yWbvoakQ7
AUR4VGJmuMOZHrs9vSl40ZAZTlbotoHRMNGUiiCHU65YREFzwow0VG8EBpM7EHUD
R6QM1VAAnoUwgAcBF1yrW3t0ZK9zznVbNy6aFJuo5I2WXq6JOdHVgmCEYybU3wrk
g+GBOM0ymf/xgD57BBcnZyTYv2oBqZ8Lk5BNYNtgnWYc6VFLVlFASdLqtM1Gg5ax
TJc0Ac3W98/0pa4hnFA/YcWppcWzJIz3YU4gJ7g5yvBrkpbEJMffdhCnUrN+2GZx
VW/D+ucLkxf+/GHlw3UoyaLJTTHFFC8NEXlKTe4Ovjy4Xob7RIAyB+CxAePdfONp
w6q4ceqbyallAH2VhpxTtR8LV+kvNIjEaHyjXAWRFT8+CDGY4ag4DW8V1dJHIoDD
//IUPcsKQtSAXaH8mwZm0nyWk/aDupc6MwXqZDb0dSa14roKZA3e2pr2ov17DZTY
xnX6bFUOwq4lH/cVTzf6VDwUDd1VF1FMY2mphVYM9O9HKWzGTNTes9JjPVe+eacY
6tDR9GorqrD0fcpbV8/06tqtDT3KMySZ/koJLILxBV1EltHvto1GnomNPIt6m5/M
pTD/zRzNr79CNtOf0HO+WL+NhkQ9OVGPXCOaTZylIv+EBsGVcFTYglVJWykWI27l
Tmb6VxGzQPrApxTcib0lHgO50M+BrW6chASb5pXfoEQskea7TZuHbU7hwaSlyEUz
BnDulEaQowE9PFG2EjsTdaUisr2iHIrEH4EiQ7B0ToRlbB8l3F411GVQY4CKQ1mf
vTYfjcBax24PrT6Ob6Jd53Vlh0msuT5Qqiamxvw4jy0ivvVDn4HAj8T7tdDfjaDn
oRqUL+dvOg7HutOjdr1K7FaiXIgAFakpaG93P6a0eh5S1DQaK9CxSj/Mm6WkHIo5
sUVMQb1lA4eLcO1R6xrJP184akmTtJtEoTgPLH2gRvTK4F8MF5zgAm9W89irmOGG
hmYlDK/MNKh53UsvgpjR9KwFPfvV//vinGXUxtKVzvGnICd9r1sDGbX+49SgzJAQ
X6vLZEkc5pUv1X/ns24c1P3Vxxhw/2TcPVyCe3qbeOv7npD58mYvROa5oktM5DIC
Yn0iSg7dNCnmeYt6IDHG0df6yIhiWLiR46F+FZgIsvh8p6DLDSJU9fPSCpbU4nUQ
lgh0Sm03P/8N8wi+A0Bumw+lYZgeiWuvETpiHZT9NXqXfnHAABI0VVSkBZOQ3C4w
pRDIUx4yatjwwszjDiJHoMAHQszkPfEzUamaBY558aI4Hd9haDsvJnX30hA3rONB
8GvJo5EggS4yHgrbwbYO6gjd+HCzz4HHXyxjvmLbgeV7YUdDKXZ5+mjKoKDH4N7t
p2OWZ2SIDiOYhVH/opBgCw9YtheSoi0K/jcP19buWLcW7CAmssQgZile3FjfsIXf
wa06INaVPQQm0fCyiEHDXiAg3zJsa6piXYmFMDUx8WRf3SqwBFk0rgPQoAdIbh7d
RGFeoRI6KbD2+rLL1G1j3smLMSWvh9LbvRUWKan745E/FyM05p8O2klbX9aiY+Dx
uchSyhMmisaIOHm9gN/Mii/CTA1LdH37zM74It50DYPqEMEm2Ov66jm5+blbUkBC
bXfmw33MWW+MoBDaGoZeUH/608JaHTdkbnqKbmRa1FgBvGCceJwgrSFuZv0iNnjf
pwC4l1McS+jDnp3f8Dv5hq0BJ+yjHFwra0kkNeXX8ubqbJlVhdCA3zRwbMELEGnc
LhGgV5X2VoP1qepQzf24CSHSPMirqTRsaa6gmeHeKZmcFmgHbhUkoQsqBj2aIfRg
XuDsZ4Kw5Z67E4aGu1JvMy0DOT02yg/obuc7BbeZVJzOOejrq5DZDUV7hm/DIw6G
3h/6piFk9AeaYH4rBHKnrC8/C+pT9CNZkH5biyX7ElGvdXfrBkW7ISyze0qGmHXN
R6z1xh/5NUyXYk1Ae5SOEcjgxfNTN9x/L4p9m6hJFU+7W76s9TubSa1FWfVIgHE5
9Ik3b5juhMB4jfupjiQZdrZzO2pB8jSB1OmkEbMqOLY1I4nI0KtFEjoVhxlyB3uV
Os3zI1iMu5X8MKuxtN3LKATBsbW12LkM0dgua0l8AuL5zvh3bxtPTlxDbJVmir3g
whwdw1IAokntiNUZtY/gmctcdvAgF3gnrAsILyUGOKQrAdbO9yEMzd4jvF7n6wBq
Z0aNsBsydShYR7NZOWt/lUclKBmCPyk5/YhVOk21GGgj3NtEwOZ2hERt/w/xeXNn
WgOarSoygUW09pygYkwAEwdK2Zd/5UVMfGQOvn+fMrqS4IB29nfneQCvpZ8y8a1J
aXJhbY8xF8a5DsBEYbvrDh2pESUCCyS8TBAQoHrfUk/A3kmG/D6ldex8Q+CuiWnx
lb2s3qLuQD6Yyyai09mBE5cJy5KdLKEA+fu5a8XCd/FiOPUmgdjx0Dfyw+Q9E/Vy
KwKAV8zd1VLPUSafOsqKUTZkchLIOBXEolhIYboncThtugCkvvMsXjrtzwhqqzbb
z80NZD+TArv+jL5Cn62yX1Pn3c95xu4keV0qZOuKnyHdOFrPiRbNSiiqAMD9TmRu
UEdeWbxy6G5bNhN876WGZa64YRk2xsN37jyi8w36hF6VAHR2CemDAVoj5APn7SLb
/hZ0gT/xDpvRsMTjBZFYhlco/YZa9yGo/iBFml5DLm83uQrmn0hMB2XesjhAm8uh
XNL3cDRSrGDfw6XHTCwPEFVfAuQ2eys5STN6PZSjkg8T+Vx/qrf/bY3pi273UoMM
RVYrqQLEXa8TiOv8aVm9ARuSI6CBEfXEi3NLLB6pdrF80rqsNClEVfYXNaEx5RnF
NKO/vDJlXNntWDq0wLNnsIVQOutz41O8UIgamQvNtSxSu2DpdBGZiOr68g+/4/CX
gg0eNo5+DZiVwOplr89oAmuC4QSVO8m+UK5/v7fpcCZjthBN3h9Sf81jV1gLY9Ko
ZOR6Mnm4U4X0zkDKN0ixtqnnv/tt6LgUiPT/5fZo0Jg9eIU9JIACBOJfju7DY9K6
hLPnzh30N/PDCaBHbxw4JqwoUdPm8X4huicIgTiMJf3PIZNy0YT98xzVvW2MSrCe
xWoNXvqHR0bWBVxqgSrh2J1VV4yJXJoX1t1jzmcGC5OatiKk9k28ydFmaQWX5yEw
FvlsclkhHOErPpTtaQfWZOABFqvHruM/0VrqMxIJNvE1HPGMINjNNZq20bFdj1hM
75LeLhSMMGS0lMzfnS+T1OCJzHy3sonnLLn4BRAfU58BILgMQsSOZhS1/NcHGWmx
Vv/VshTS7mgndL3Jl90Sp3VtXToW9T6jsiKbKI40FTtOTZPJJExoVke6ZT1+tduZ
O3wo0KoJXfdQU5k+4rdG+cOafNDXIgKAF1t2foP2boJVFUBI5FKooWS28JJFqF6a
5dpfXEF8P8/279pWehPEdG8z2lDWYsnagWYVJBfF7oGl+G/NGOuHC8MWi+iD9m1+
bYSniJzgaKO0vBdjlon6JuA2myzbUPMhDyHWOWzyvJuJxVHCrp/PM4+uI64Spzou
v3OTNjBYm3jbHsTEm2tq1+nX8teS405c+LMAVYHMm6ZB0it+ChIBMW75ZhEVrsrg
QIRoaaX9GH5d5+ryyFweqg02M+4XxHxRXHPHf+M1jDF7oj06QON4teSeCGdWfCnb
fjfGG9y0JLQlMnxi1Pmx6oRZ7RRbP+Xnqj+xoCeo1fS9X+Q6OeS81HotNk5TzaXB
FWGPSxuBKLFdbVcoWaH8ZEIOy287LrUyyurGWHioxIzvQDeZmu7rqX+Qg0oKCfFL
m4SaXfSTIIsWkoGyeNYZW/nlGL1QcYFDvY9wNyBaA+kIydsue6sio1TAAEOZ3rA6
XiQANwhSeXZk+wDNRfGfNII7MYKg/q+Vd7M/ya5pBY2s3+3vKwhgONwjczN0FnUg
X33jiX5P+rhMPPl8Yecfz8/58TLNbjaqVn7pnvQpW/H1zpyZOzfKV6AfuBltnlgx
jn24hRyHrvnWu5jjsbOIHxN/wP0SH7VUNK8HZB+zeZA1dcPET42eda4lNvgHTiQh
HgIwoIs4RnS0JnfmW+DdLFzR6pu6Xz01RbQCuWG65m8m3FPFUbiiLAObBojAnFN2
muYQqpEA6wVlgOQzfK2BRpqHRioNRNPjpjrsHDOp50kzt0db2+9jtMUYaBDfSbAk
ScTUGEvU2G6StDgwHP/eocO4d+nJIXpHKEDFUelZ6CmFWN3uUTDp4eu8vTg62JKA
2QrSnr06x40ZoRo7XJMvRLDKEFHCMD1I14Mz3v+piiw/fHgn3Js2rmNhKULzO0tO
3wNppZZWyAJcxq2JQcWuVAobpmHwVqpRGtoGQ6+zQRQXLrE6l5oQwuPj1cfsfryQ
BJnf42xPUdmWZpMnXYKxyVmbb8pr5oSJ7FxWnROVtKVDOjkkgAs/ziRceFXfOp9c
olQAC7oXvP0bZJHti7EFsN/OBWpPqqCbG5Zt45dvWT/l1NvetzvnqlEW/ZEYRMwk
aOTGMNHpI5338784ZvvLi2WjESPPOaVMxVuQIa11xXI6yD0UW3TU4eO8phzepaMk
pTER08g/qydI1wfvGvZLb4E68y5KcGv8hJ/hYaPqOIjrMybFQYpViO3pNPsZtjJD
zH3NBkntUBfiTdUvq6d3QqLV0L6iSIItUu9d5blY+11CTkGmq7jkXOktol3UOEvU
mr0oVtI8pvWdK8SMPKZQbIItarB2SZt5CnZ84ssNq6DFZI1NzE1QyWyL4D6+Q95d
y+w2Q6gmi44Sk62S+yySZDq6pcXzdzP+wLwBTlNWhVvgEmHqt2FJ/mZfTzAu/U4L
8v4kxbkSQ+afA2Wj14EwbTrin2BacSQVYnaSVa/DSIqt3+CjYYUoQxxgtE0w2B1x
M1/+ABY/3l+VId4evw502Axg7XZv+jy0rA7G77GC45gNw5qMD+nsgRWac5Tcyu53
S6wyH9Q7HhR/a60h3Axf3HqtWbCDU26LWo+CQNqJuil9mrCqAxEUmOq/5YhvJA8f
/xQ5Jf08p1xzO6UrzIs0YLmytmO6zO7rUokX3r/a7O0/H9ocA1TCAI/UJtjA6G9j
SbRjBhWmd5cgJz95gCrpvlgiX5egLLW36vdZqLYA2feCA8TUcCjPp5Zo2ypuBSRL
OG6auFGXE+rt5Xv1fD74l4G3cLYftxIsyoyjfV1XzwbBCXyhSInx0HcHzPH/Gudg
NjLFt6VjV/V3r6eOhT9uFomFlRSUifSJxenuU7prAEshEzHA6DPqf+2BYCTlHvG7
vGitnBGl82PpqIVELlPq197ugvqW+5VP336+r29Tzy7CaZTAT46UhHDo6hU8l/OV
dOaRHN/rOfUE6vyIGEORFsrqAevefpLF245sqIcOJtE+IQGiPZU4PHwoPC98PTML
ejVbgoM4pCWLWCm/pzmWmwNo49Kfk3Yt31KZ7SMaOFJ06LTn4BXhWzdu+5ztRVjb
58/4hIZJrNz9IrlLlHeNMKt0x6shUovTcK5j9RzXIQCkvF5A25esNzqzPpyXVP8C
Z2xP9qSyp9YXbL/RXnqCrRh5kudZDr1NbrW7L41iJU/5LzuP5E/pz/Ul8Oyp2tSt
MlGlZWOz+31qhZp8tul7Ddod0LwkiQp3ZBZkJr1Tc4PMzDiviej4Bo8NiYGRDh8i
7YyL3vNw2xlt15IxWj4/Sb+W1BhtT+8ygp6QTQfJ+tqbOkjloPCKXAPlOzthRut+
ryRcKPo5ZL6XoBlv2D8uMWKruEjyIezWioM9AfoXaMEvPutLUVhCbgA5qeyn+pUn
FyT1ppVa+2844ZYAxxjZZsG4VWYDAI86otsYuhjzciKyYDcPxGNmTU+lXEZefTfX
SSIr/A1z2jwLTEQModf1rsNgtQq02E5AesdeJUkxgeb57JOS/h3zBzAChBRx5mw9
Myi0Wc2S96WcLgC7Hc3dOKpOosrLRuwZpLBtZGwKCWS7t9FVJ0kX6fa6v5oeobfR
M5CgCJ5AHX/MwTQZZ69xzmlVU7LZYgVn2ryKiHJnF1zyEMbkSQYj9PuqMNllUFS9
BzVX4wJ1524SleDCAIp05hEpxfLWtSLT/oJu/C0sP4Kb0EwTC0mz5Z/3k1mZNCBM
H8e6bL4v8AmCi2uD0SnCyl0WfGUr+vnDkNGN/PE4Pf23cja3ehufKzEM4ENyjvAz
oFCwj0q8qgpqsWObLx3rkGI+MKPNSBYR9YBktHQdfP7c4jdFZTTDquIEXMvTnCw4
z9exP/3/E0wjuvStnVvOnKuf4cARYlrOuTGQUwk+yWmK+u8G1VFSfTPsQckPhYF5
as2n9KU1sSzLrwJqxbrK2vP0UfNw/Ts1Yd4G2zPQnYBNOzwTfxJrkPUGBuu99/gW
EJkorvf1c3bHkTOowDcrMCJzKaSDBZorhIBx0gZB8opg0BoDuHa1Xa8oOf25GHj3
3kFrTDvDpttBfc1vdWK3QjX9mBIA415lfUL2tVNAjghZVwWT5CVxeykFgWoDREpl
+uhCEaz4DOSw3VGR67tGO25iHFE6VwPOV8RYng5OC2npSfzhkhgpApXMr47gyELZ
H8eOchKeClcUr2eZXSHRN2di+uB6SR0pHyRue9lJ8U5J04xmJ0iI9SFs4hwhk7au
rExpnyde1/TvFhawPsYi6B4OkztKZ7uJt6F2xwmw9ydE00nWD2NVZmhGJCJFwsLY
FYb8+Jymik+T8vWWzQhsysWheKX50yJcd1yCZdOJ3Kt7JetmAZG4xIwZw8lNGXcX
MVfwXdsYb/FtYwKT2VsFfpohO3we/x42Zp5HF/GqwdmAU8zQmRtHRhq+ADB35WZy
GrYZkz7ucwMKjro2MzQ2Y/lMrJ3yRvS7nprlYMTiGT7ZWz4nW0YW5XL+n0cZDkAW
WUzWs24Ket5Xo7NODMH2LD2uPghJcgHqK1/n0jsMrZXvcKuwOHYl5jzoNZbO6+sa
qbuvSc5TPI2Q5eSqDRlOH7cGZUCFpxisG3GgWIxZVUxKeNCR/k/1OW3Ybhz/NJAF
+a0jHtpDzm1fCdmWPPuzst0qHeBBu8gthd2CZA9ve7fghyripxlsQVULQL08WWrq
KWlHR1AmXiMVbop6auq4yhmZp80tG2C4/qkpdrfyOcG/T+bMQFPoOae5p0112ApS
TjI5PMMQXhD50Bwu5n2oyiNvFYGYgtqXz6hM/05SNXFaK0a9NraMb8qtKXn4yFzL
IugpHFapW5+HG+tjya1sxGJV+T1ulpTgSKoqoOFWALZIBOHrb+vKZnGEwXSoy5sY
VeqNGWMiKoQHk9byo/xaI/KOKQoBAlXy5BiXyr7xet6oyG192PYmBZ90dMChLFUh
2LId9txkE4jHCpCiz9mBX2evh2dQXJcfZntcRLoOjE/7+j8ZzQE8Jq4VnHpA0MYw
xFAApC4AmyML9y1WM/I3Y3FaqZErYhN8591VbiAGoCJShZyjoqnCC0hDkPF8LLLP
u9XHRs4C1darzyKePEGUnH2gW7Mf2+zlRF9HkydQtsdSdiS2vRlJnqctzFol3GYx
ZTzWCLkmZj5ovsG44clGM5fHuMnzy95qdcWQIZz/Sg2VcM05/gSpu3qA6d0GXcBG
C2dSQgXW75K+k7d69ylqbAV1W5v7kpvVPxPnjSp1wuSyCIC1qrsdLr0oCSSnm7Fo
/zySRlA3pb5RVAuk4zcMQ1SX+EexcmEAZvrbXjD1exmb0zq2zjWXxmbUcZxpNIHT
Puo4tRpuxKp0MtgcWpBuovuQ4ZcZ0BbGkPiI37gpg7d71jGeW2uXKZqh0pPA1Svr
qkUTB3SPSJOdA8jVZ+VeHxiYVAcT1lu+w0sdL8ZHfWDGq7+WkucNzo99tWK3ts1F
46129pLgZ3WtT2aeUpTIvFdJv2FLpPzXqVnRHc7CdGqGJdzWMHg5NcnE3di1pLfo
TtizoHm7fYsJdUcqVCkA3kZnnPgwjH9bZzs8aolqEVr8/nb2GiYdhQXuv0DmwKKx
U6Wlktb96w6lvCkPuvZ6EWHZQWiofNFVioH/t5MJEIorQ/iT7hazGlu88aeNws1N
2MvnganZDWkIJEpRxnXbMiDiaG5BGuNuclUHyyewNfBntciCLuMKMvZ9hAYY0w1K
Um8yiJ18Qbwc39pxeUEVgREgeBQs+taD9FurhMv8mv8mTZHY7AD9hcoR4iyXIv0F
A/RyedIUKa8Ep1TSyw9OGsX6XPVlskAb7S/afNiKJ3CSBlALBue51H+ffrar8eaU
M84JwjSG0VIXrg7zzCIDsQdmFndT5qSnqjkK6JMHr30a6K60l6hFGPmmvYkiGxMK
KFpKzYy16HNOjADXHEOhS3dX6A4TmK4nAjjpyvZKuAByBckLGQmNSg0LdpYfI2Va
bAGRE2RLLp4PA+Mx79iFBHNM05iQvVwtE5d53A81GvAPa0WX9+MTP4NkQJioGNKi
pZ7XqvUFjjYpRPEAseYMCt513cVKDuImqw+Pkz/p62JFv9PnODef9FW2CtDEfkzU
nnp+bNO9GNgZH9q7AeyzDdUe6Fse/oolfea6/K9zRiv4M4tntncFL5xqwzekU4dC
gQTa4wLR9PL4UXB/ip5IFB90ZI2OG/w5LQzAyGjH14RyL5V/QkHmIUwCj5U/qpUE
hL/o+rTpgNt8hpknlaTVccz1qr74krZIoMSvAn4puqQ3vxvQNDYqOX/PgXgjsQXr
wPtBKY9QrgBHpJlNcWDoN6Fa/Jw/qUiVbN8OwKQwfJNjXeOq8CYwBCJLJ2KrjnNq
dBKTrgGqoUyiX5kpxiE2mafoQ+GW4om+pZryio+dm5e9zJFo+QyFySF41i2SCov0
Oz1ybQSHDqF5kP4kCVY4iia7Q+ChhCGLIJHtGe3aZOZy4L8GZqcwnIkj/R9mkDLE
X3UGOBUNguwylj53bvnR1vr99p+QSFj7nUbvwUcNlfu0gqlb635GGYX1Z3XdejWt
ExCQaOApWerZbdk6jLH0cjiNAT/VOuJiH9AgVAR8Oy0jit1ANgAsca4F9C71VhKw
iqrc9V7i04fJdtgPtahNJsa/Dj6Jo96/4Yit5p+hAYuZuoBaeKlOSwM1C2Jw51nf
MBC5XLQ83fCumu5UI5M3I7NaGfOdZZJsfYwuxGN9yBkEmZdbgp99KrvOlWK+s905
PrkcDoEHO4SXUNWZHVwIFScborC0+vElOFQZ2OclzgtyEMZ9su8L+d1uzPyDFwVK
V2k/60V9V6cYqZiqxbAAviTPaMEiV5IgG8Zl28TxjbXSVxa1t53OtfYIYGd3jPQR
Zq/RzaJPQK1yj/GwbBFge8MBJlaWOwQ2d2l+wl2Z4m08dweSy7azCUl/xm5WRXcr
HmiPLprEEqFjKlV7lE3yaNqUw+QhgFXYl/sVLZ2WYgzccO0TjrxgUCb7AH6xhpCp
WPQIjc1XhBt019My8OVuSfMOOLJaZ2fTMRa2KvtEb12Eu0Ptem4jjjURo/y0YWqR
59n2tncaQx86SE7g+SiOPdvOOml8exW0x7YY1bUBUa1l4ZmX/TN8hYV/whSEU+Y2
arG+vuNXFFdB8p2C7nsS9QmASVhnQjAhJtr3YKb4DRWcwFlnfartKdBPiUF1dzms
DK6wIJOIg4ewNJmVKgCoEYw+YId2fJuRyL6CMJaa4IiijcUgOe7BITeLlWw3gAgW
GrRFBdJeP3kUzs8Cl6vaQNfffsQrxNeKkbmgNsqHBN9MQTHNrkzBhUzt4k7XcSMC
OjtUs5RyA0uLfYpYn9NdHNl79zWF+YXJzK9OGWCLiPyiSXRdEWoKauzkZX4ru5y+
hfu62Bp4TpMHTFSwrOVxLmg7Zl4L8p+Ebi0U45dF2gLoOqYIw8Rxf0tWeHLcnLSc
f5nFfmQIJbzB3iTzJdEwzOB4jkuqRXV0ppTTQNAKcmN8ne6EAmhjBGKHbNoylzpK
T9nwYVgH5jDP5/3k+z6urJr5zD+rGVkSzOsnkt9JsrAvvP988DJalLA+D1YG7t+T
0MV2W/gPldnf/KrrtrgFzii9sJ0Th302qgzTioEdtYcveK+7N9PH6dwf2en43c64
aywz7G2p+h7/rcbTmq9fjcC/Fr/sH2dey/1PUpS4zXrRxLzcOG3IXo7rQ6cGXfuf
uzs3I3wnlNpF7KEO8IXxSwJD406lR8CJojT4GTY5xK67UN0IJJnuucYkF6/EFBja
HCDlJYkFzs64AYkgMgddESsciOejVkizxBJ7khh5Jrq1MqVnO1vY/HDx+u0MGLl8
qDgVCVcbJbhrNzZsYQln17ECQTnkPmjh4UlbJANUypqrSgyfo+SQhcMK0sE2YEoa
GR3CYobDjTNM0eX0yktbqAC9wvb4tDk18TamJC60eFmhqghBY0E4bhrg8yqWpgr6
h3v90ghHxQRM0ZY2xIr2NaI/C8YtNNnTHU+cerFtjtAwZI1p0RL49mL5gBscb8SY
s7fETspcnWNcMm6hm+bxXR6dp5iCbLC/RyDa7LHtjhrIkP169+AU4nYPMlTVpoSk
taUdb8jUgaerVdhu8XeMHWfiHm5BPCctanjpeAVUmgdVXRWh4LLayuKAiMK9Uqiu
fwV9cGCwJG7y8d044+F+10imdYmPIc3JsAwvs3YalZrAzWs7DmObY3vm+2+yXyHf
D86ZivnAdTLflLqMU+0igsyNhVZFsHzMm9KOBc5FQmPm5wtJD0kBy5RAf2/IfXXI
wAZFuktHiWqfd2ySL89zovAlzizwDOkmRKoib92QNMeCuhUl4Aqu4DQ6A2asK6Ob
E4ypY40n1Y8VWcTaRpe+sj4HkIWw07BInqztAb/1KgviPGONouTmIMCgUOEjsrgg
CXqTY3ZsMeCqxO8MNzuzR5fDyb/0luAAgRFIFMTmCFw9uno41BeGEPF193iH4pVK
i4jFeS+OLY92c46ndlBOoTaCymsORkVtzuwWqqqbeGrYpH1/2tFTAvnZhvMYlk6Q
kuvQdySPkoXSaLenIvxbBvyNRsMGUrNnF8WCANkjLf72LviJUEw/LxNXf/mmx8on
pa7Pp5ooNflQ7MvdWQMan/+6KTeuTqZlCtsF7At4ByX7oVYBXWGYIzZETIsNFAnZ
Dan8PDEgAvAOXUxR7iVoQ7WrZATJD+huS66sDyk4bFXNbcsxa6sb/LBpzCovrYac
Ooz1wurgcYfU74YVWGVF20zn1HUaP6xVVIiPhenZ1iq1Uzc+ebqwk4zAPdH+3/hl
RDu/Cw+wxKSEoUimD3UDLI5SN4e2CZ7KAtGgFNX0OP30MobHgjO8njb1sZFcR33+
k+Bg43sAeYAdB4iMMzzCT9RUF2ubtfDvTs0rhwHIg/bur3kZQSOTKczuHA+6AwPI
CEJXGE5SFEoZMwamaRoWmkKQfz15v8L7sVKbyMrTZgboPzPeufgCDKlbcRv8hmUv
a6rw8/pybYAeKsm7njO8aEAPUsIF6kpeihlvE0dWPjRwaONhQ6iPgY9cBVajUBjO
8VQjbgQe7wR/8jj8ES32rG4y/vQr+x4EYalOWM2qqfE7UX8awEF6TiiHZBkyzcTx
Oexe6YwcSrmjrFSopATcM9MjWHdoj2OMXQtYEJx2Dy5AEg+q5Ms9b78OYurzTKOD
DotExV5khf4Dm83rrxUtmozNPdJlfLvorempl0dMkeKN12qkH8tfsLBrTzn3VnCV
7g9oOqed2GqLLtaIV1SwqdCdyf+c1uw0nm7p5520dvP0QZ10eADyYjmY4Set1NUT
YcF0Z5W1duXO5Ze5uNC5RjgUFm1mAM9Xu3nJbdfogPia4NDEpRlUxSZ9u89245EI
0M34JcL9gWturfotH0vC3sJIeB7kXBEjyjvs7BoeEIMCMv8Ts9wLmswajQ4rptCM
UhFx5+w8NO4TrHnzAq0NW+4qcK9FR3XR/8q8vfTjA4t3FfPLOElHrcM895Cd5ZiK
SzEyZPO0kvXXVPEcnZxt/9EYXksU97eRyJlI3KPmeQApn0DnOwZ5eVFjoDwvvu+w
D898Hr1IN66JhLxqJpp5H6S8LDvT2MyfXFSqVSsngvU5yuDKlrn0Ha9bibd1dXZa
6XQEl8LBmBoGVB9sKMirHMGlk15Tb5HcE9+8zTz7Ezie8lL9NoVEIgy5aiXpm497
xMN0DH0k8K0WbuSC9luZ9yydSrAXKTDZFh5BOtGEZuIJ4QSSPRMe75OpNwIJ7kI9
tmGHWIM2XzTco3hiZ+FF3QBvy8wI3HnTT5LU8EM85wMfP/LfPYvU5ZB/Mir0MHVa
9iUWGECDoS790iSn5EFy9cfXIu1XH9Scnj8/+zAqehCEk6TXp6adtIHlHhhzJMdp
tUz2h73jvxYrW/tOBiWfwmUYFwUbjUjBaiWr9/fiC4TS5+soaAiH/dIm9EFinht4
j9Lp1Yqp9nhOFU5fInKbd0xJpNuewwK37rzhDDgQRSDuCmECW1loWJ09McTtALP5
N9t0g3QkUi/IFWLCn1p4dyoQOkx5fVmJquEQoKbASmSiN5VwjCUB09zS45GaZ0/I
ISMirUmtRuedyh6HqU8uFSCQM6F27VM02sgoEZTh5ZJK6DikvUSlDQvz50Tfo/t2
f06gBi8I/qSGQNXQh/GRR9KtDSQ0T/uevHDL+5rg/3hHynJC1J6GnsH8gPY7bnEy
WomBq3wXWzX78sPqw6C56/kesjjh+MBJs9gqUo/b8P8o7nRxgfrx9XsgD7Zx+Jbp
RgejDGy3FEc6fIgSbHbVMdsiD1y6rN2RcJ4qWzA95qsM0hPpveCOirwfTJ8sYNY3
JRdTLcNQWWpNmk6TYeMj2agO/91svlGhql5Y7m/r4038e5zj2GPJkqa7g/HI6YJr
NxKljQtZxr2gmVyRNdnGYxI+Ql7kkCpZGYAOmNTSkzQdi3tE4Mas2uImmyLK/2+r
VHyd4R/sP8tKF3ayUT+/SJNXrAeu0FTtfNEPMQJICXYIODVv8lc+U4H5lBLZ7Sc6
a/JAtLcc3VkVB0bCF99x977Mi6qGPd2cMZIE/2/UT79QrBUl4MZmdSKnX9BpE6Kw
DukluxUVkoNDngPTYdFBtBby7g+L9Rh1aYW8jlqs2fYh0FUcXoc/bS/FgQv1UNYy
qCWpvILE/G+xciY9tsXGynpnktI18ddE+HMj11PZ526xH24IWqyai2ed0ioyI2Y9
V2qCHJZIMNQw6qZWJ/COHT86TkkyZ00d4Iz17qSr5txEs+3GA+sk2k+zTB3rbPIW
9Iw2qNbBYlS87bxDfZ+iS0pJtubNbA5r5JJXpHork8fwxpbdXTeqrrecs3Cz6s8N
9xl8Q2+JuaDwwmV7UnV0TAhvbUGjKwSd+u4XZdNIjhNW++f508Odp2Zd1zMbbXlN
UNJ/XE6PLk29b0Tm50VOGG46+z4zSlpRE+k/Wejouf1gIkmRGcRjMaSjUKcNZBuW
UCOgcojgoe9QcsK6NHobUUmN/G8uk3NbG3MCQOY7OOX078yqTMz9VaU2vsl6RMnb
xOlJaFJgO9yVPBieTiCEvQ61hOoeUbt5Ql5VzqUHeGCSOXqR6PAkAZXD2RvM3vSd
gEsYyj+f0MzEotzxxYp3CqOGFnBwwROWtWxayNT876SB6Lje1UDDIaRNqH6jegoZ
DfOSvStYJ1vziEenTFEG3+QjDR+/RYtcVitdRI4gnbX4zNPhHyoPOvHNBYWvWLGM
VZeLddRzm4UTVQo+rq/LD70borrQVL9myJJbSFXX1FgFCLH9oNA7zHd+oRhLjnlj
sdS8H+jw6n+gRjRja3k+YqZVR0MbvFzXcPcRx43vFIHOgiyMwlUCIXSRzBMqjyv1
UHc6f28CLnHqxHf1Zd6bSv6cZeRARMFNzTNoXXbd4d24zndb6Oabvk/Mc7pWaNtC
kxZi22/9xZtrR1o4MGtS+U3lWVd2Fup4sl2nCikWAwCLbICVrhRNBqRmme70DMaZ
Syjqkl92wXAezRh04F2sTyDA7zlIC2X16V8DSURdQBN5sH4e7QOhsJ33WTCERD4Y
gYNVL0/SAOysJVP8Jx15+657C2AtViYScDY8Zj7O7GpJagKWkNW5JsVcY+o878tI
s37sTA6Kmu/wLDDsQLEgkKsFn/jw7EiF+TFTmbj5uU/sxNVhPPsmiPNQ2nKTriyw
l+AVUZdj0/o2/TL4E7P2D8Tz1vg4T+r8XOMSgsO5CiN35V+WsNas1CegrGqzO0Iz
Y2P3XqGZVyOVg15knKhIFQPQqKWMkxquEst2uigu3OFvzXaZfnSzZ4Or+oc18SOw
lSl2xehGbuovv58Mi3Ka0BWNMTBPd/5WDvmv15SQV7ZQKGLNYXSa605bEv+xoH4v
EaovkUoQ3Dv/4gZc8KedaWbFY7NuXfQGl0XenxUQswIvGJy8UsNCC68rRNFmzfL9
wTWss9btNgq22orKWBFJbN579OiQfLZs0dkxcUlQ8lnuCWTSMFhBdyCzv6Z46h59
riSIhfcLPvEvji0qE1OyE6KFpQDJIAtZj8hl550Y2+z9vanegdNjSR/0MJ3aGAqu
pCp6txSSzAP6BWRUSc7Bu5Yw9nPIlPpcz4sv42OTz4ELbs0vqVdGTGlYCMe+E45k
aJjyTgwCAesI5VyKtfC6SvlVqHueQV7kfTbgz1xcfsRNFsHBLYMT9v58UIVoRRfM
8gvtaiRanwsF0voNZLA5SHI/mrHaFUM28MdmKETA718gFwuLG59Rhuqx2CFAHKZB
EbBV+E/hK0KIKxbHPoDG/mSz3LPfGz/plrIdhT3qGFU3l6DpkjjEG+/UJq3w1ePL
0tt0juDVA8qDZ5Se4dPNgpmABInDGEqlfr8plUJBYHWjm+mDxEM84WI+qldI7wjs
725PmMSKhdbg0r2A5IoTtnTRcsxr1m5/aM+4s4ASZxEILzzdNtSz58rtsJJgNlUi
6T/duoeSI7UoJyegcAYg08IXelY2kfTE4SechE668nQbaCd/HbD2h9egj1cVaWNs
26M+np7oGeHAqbT0n00CSDIht8RKa/yWD/VhUY5JrVAQ9/TzK+a1BS2HERtOXE92
uudnecAA9gikDz2PDpP7jekSI40GC6i79B1j7yrmG5t8FTs0o0r4wTzfXj897HlF
G+S+Qwv+Yz8st4NmZJqLlotDUBJ2xbxXEEbxCG3yrcA6Q5Yng2O3MJsLwQJ09AXz
ALwlMX/5KepK1gNql0norzNw9zPx9ffmpGrBxngMA8tv9izdXbhg7iUQJGCplPQo
BMqCoL/f1PWW76viVsaahkg37KxspkDcftpBuYtuCUrCDZuWnwuKkMLKtGkqme1I
1PCPU2JxFok4rOkC+K75ug6F5UUM3/CPNkcuRSa07MxMrxN83HbO6OTFRYPDa/ch
kfHNrjUqsnl5Vn59hx7oCi3Rx4gOJfLjHRD5ujZKQlvlfJy60TJLKjLj0NuJpCjw
p5QULbTboDrwcCMyiQw8Pr109r0RbvHZzKrrVpTKQaFtM2C3NqpmjDqwVqgE7Nsg
9md/W4QpYSNOvRdPFt/i2JUDA53mQsZhOkl1x0628Kkn/7Gh4aTrKGlvxRXdFvjt
po/KMmwg/A4r4+OKJUQlsZLJZVnuFkurGxPY9VtgwOHDEOMc1cdbfTBOCdwkONLT
aUFbQ70Z6zlAyWK5CJ0reMS9LSyS3BsY9Ib0iAEYNh5xJmqzo+J6z++5VD3JMYHF
xvZGHZ7BAHfUkjdawT8kWaDEB78PsieNIVR+SLcj3kGxymZdwfSz6ohrcqyOCe+N
m0X0diJVWJIKKr4aXqgJ5sd4s1ADtapoT8fXe77UYFJTGZOBc9D1VtZgK9RC4jGj
iaaNlTtqVYIIbUE/v7HBQNfue1ayCE+2X1OT0Q2C6Nj/Lg+sV7G099MNZYfhQaOC
LT3tqnfyIxZB2X7nxn1d0SVnnkaihGUq0seZYqoVoYINmRurkQ6hd6YhOnBVT7v2
O873eQ70fXhwskQFaHmXaS8YHIU2Ht8TAV+XoqqY4RlNaBQ1vjQMWeitxxG1Woq5
SS/cszLxbVI46vtoMIMvwU+sFf/7mCGQG45JFnPn1kpQiOyM0pyEn43h7nIL9nn6
dusElkFbQxflK1os2nLqEQ1peaInLkTjRf3bEz70Epas+YYdzW7YSeCz5HtNGAqv
ngf94X/dVb01fz/xc80BXMg1BppWsyKV2uBn+OsmWZNIei9Ee2ln3GKKXFIcEfKE
7GGgmlpqkFMjaErKBqh4qLDk3zP3jFz9dexnlMpRFBkgVlFS+FzgGxVjt1mjYsdg
00Pcrvy+R+LwntZE9c0+1nZCZXrvK30WN7uyVcSsG7eKWVgk7wSCtCfl+QIyQn8O
wYi31NLLscAoyVj8oy3MsJa8TY9hGbaXPktib5mVwduD56oPmDRafsAzwlgSnRys
sKXoAtxYVEGB6fqWgD/Zs60txgcaO7Mw8AnbwyKfKxJb1F7ofXSMp/TE7yNVbUr0
pXfRbRzzkqzFE7vB1mW6BoWthwey/z3BlxEJD++QKNIJMhUDpUsbUrq6MuLx/crR
0/jrimxK5pG6+6G2dW629fryF6s3K9YN00BXAsyHZT580FyzMePRrfGfks9tdYBl
BZmTLB1LNxprEA1DPV9e6YHhkeLzvKRPYIx696bMTkPxm99tEuUNNSm0KEMDd//K
sGmQJw2i2TBQvcpSCD8rcmnS0By/UyGV/EOBHnYbkZ5wQBq8OBQcE8dpe+Ml5Wz9
rJpkBYYxKNwIQiouP9DHOi6vInCv5jE6ZzAa/vd+bH5TFG+phGYfWKARauYiQx+1
OGY1or4ZnvXA7K2Wl2nWdG2ox23y/s8v/J46SQo1X1+yLlmJrvjyRHlXOiLxRnVU
ZUeWnFcZLI54wITnAGUWbpWHzY4xeiWPYE0zcul0w3QQmggRzamED1ZUrdFgNg0u
qtDl7LdqEI9WDA1eh4TsDCpROaOISFDT/K8msoSa41zUVH0YsrwmU4hcd9YLq6he
FVPzqYFqAI9RCavXNz3hzr5gvxL0reynl7cpFbJ8apL5fqF6prGiV+19pzNS1Bdh
NURiC9nndDHgg7ubJy6OlNJcTBl9jRsIKKfRsJSJEslk91Nmlc2XLRg0tedBWraR
ux59AtY14nF1xQHX5DSKnZEJd4Sxb1QGQyhWfdkBolVzi2erNaiNGXGPi96KWJvZ
OTMQ4nyr6AYl2OZ/LtG15KfRT1XV+C0raOg3NV4xBpA8kSNe9b8uRonb6LkOAWEr
dn6hG5MKX1MLg2JQlsLFdQhTy4ai42AnSmkRJkLPaakImDAC03LpSGvtqeHQ/W+2
DhD4D/IjDDeEzxnI/r6j0PeTkYw3IPDTcmeUWUnoqol12IxX4C2S68JxN6YbapWc
ejxH33fADh/SekVe3OdhTebc/kbfxAInVKTOvSxaRJARWbSiZhGFmlNi7b+KsCP6
4Xu9cZIvnDH7Nwo3hC2Ss04zEpm75IfBBnnW5Q5TcyfT464gf5RwknaDgwCPLVMX
LRaNzW0g6+gUzXTWwzELmmq0jvdfcrRndNzXIitSx//ATwyLKh2kmeCCJojnQB/a
HJvlRjLbASVdguMePacUelrBax7N35ESNiQ1eF4ooLmt98TulltsxSjRpPtHZSpj
LgD98QY5da/eTjfSB7aS7HfdC/yiYkRUYQ8H0MUyhwLXwSSOD0fAcakUMFCs5eTK
Qp+w+luWC/Uh2Jv/HqGKZLpnHnUVNx9wB92zW24bRUcKE66ZeO/M00YCltAA7vkB
1V7DX9ztmNIw2wLASpjVRS5G7OhRtySNP1QzQmLWa2y8ePdvjtNigJcY62DbmVNc
ek+ySc3Dhs++bv6W29GIe1ZKIGhiH6hQMDZni9L2Z21bvR7y8JUHWuP3i+3hVtIB
8E/nx65Zg9v/n4PSn0206nEqs8+7l3os3xph6CaZRBD4GupSs9q9tFFv1sz5FJgH
XRWOeS82Zxh5g6mpn2w86C4bUmOWerdtNWRwOjoigYxSlzBn92Khe9RoOp9nq+Ip
oeIRZC/CsAGtnCtRXkad//tqTI5n5DOP7jPhxwHFT/pSN6dDuU+HBzpAiWhndf6K
VSAsOrsWgoY/TbaEQWa0aZTJttzSs9kIq5XEUebYnjk7raM37wVkZee3roQdGtQ8
cJjXAcOcjGXIY4ljEVl/kWW5vnZO0CSVbOKoDl+2LRs+4Os2jTIRMf2J14D751RH
Q7q2BogHSMStj0eUI1xoBagevxw1r97/4/thw9zo084+FqiB0KAChy+xBKNThDuk
tPuq8kXT7OGHDVspVBShdZcZgPQs5Sl92MF11aNNO1Zm6yI3vrm5iNcurBTwy7RT
uYXiXp4t7ruVftKWurncgdzoHX+xUBKlH65OhZKz0G9iVZ+GgMuctN0Cvhje/1S0
uVavGHh0vRv4561oznovBAgkdowKGsVsk8D6ZGKcpJ3DKWZDqr4k+ptkzA4lFuzq
KwE0QznK3+nbtmqiTV+PYueMs+jr6s66WmbgtluYoyrM1G0ZGOz2WNlEwQurrstY
ind+mhfk3FeJSM4QiZGUqQXEEz3TP1F9KNEtGzEv8jYno6vdrBt/DjB9/BYU2i7s
YlIBCQMFDb6CMiLNW+MAJcNpyowNyn8nBYv/kmpN3mRii7exc7/759+84WEvPK+T
8Y1wxHFpdRNqCsF2hTxoxiJKrHDoTE1ED+Zrzio+egrZrn+7UUGy6F22ZQiriEVV
du4xxjvz3L+/nC0FvgO8p8D8BBOBlk3m5CzgSOaydA7++tbH5O4NnlWDF4YPTA5L
rFGrcQQyoU2dX9c8lGmSiPwJFtfavHmGV+QOZyoIQHFRUourcdBOdfgnUXPrKgDI
TAdfR8hrfHgZQq46PG3C8pmGoWakdXk4L9815+xv4Q/nTObLsm8cLyVfDttmh6+h
28HI928IOOFw2uvyzL7r+d8y3/j7CV+u8tdnUwy/WjeRxCl4gEGZJHSOIT3ShOeo
3zFwbG/ujsBbAZs3A1k0ZtkCU8yR3y5GpjVg4kEk0vj7M7niSku/1RB1mxHeB8FL
srmYgaaivZiB7y5Y+gTcVxgg7/F4YZBHcZliFXlHhC2NE38IG6E1q48wV8EIlStt
m3baeKR/RH8fOSE5mSpNrcxoRnYqnLqZ7swC2XBqK9mAXT6uR7a/TiyKrxbOXncN
ZX1jSLLj5xvUzEE0q2XDycpJWAXZJyQWC+t9KdvAKb9M6HbUKmkzS0kGQyK46lBs
WTsXPPyYJ9O6H9Qa9Y+PpcKuvpCuUzMN7qNvlAgzcprCoByzOdSlZRHrAhmhMQSO
JhcVMyAOLQsvnC9gMddT76DTp8X3H6g4yC8DxgxE7CDqxv0KqQ1mqfve2lnZm/6h
kCbIckXEIEP0a5rCXuOQzEBl9H17w+gxOuU31wNkrWebpTiQjJ63rDq/GU2hcTdd
z4scb0EYsBDE5JRkJV49/ubEO2w8j2mQDNFX/DNEzBe7jHLsGI2dsCHbAQ3W7m6e
136xAw9M69nnddsRQTlK6URlkGMVXGnmHyAvndJgFSz9+ggNgRS4/y6WfrV1oLa/
pQsVwLKwG+hFHaM8ES7AEoulVfQ+Ft2VUQksDy/XpcTLZ+itiPEBE3iGTkJBKLWK
ZTlz6QrOxTJt5406G5a16jw1JAXYCc/b9PUX/drmk/nCtjL2P1PexCtXOYgsts1M
+m4xwq3UgxOPoXOEHyStMASkkrh4U/Ugv1mvf6J1onHvH6IvbJarNLbVvyDV4YG7
tAlSpyPdesrlbmFQuegwJb7hqX+RsCNq48l9R5E1XVwNl2YuwLaKknVsw8v/ViAc
TwWXegvYDmBzl77X5jtlgTxeR2HyAKu3W5qqGKRYQErJTi9AnaVYgrD96gyBt4d0
g7zocjcDkjoQ6qSkm3rJfVwhzpzO0wbFtvF82jkBX9CUhLOLGz6cOKTn9EsjKk5n
xZKy7h8/PMaB0NR8YAIgOjJI0iolw+sRQXaKmXoIeUNyTq9askM4vtlD0z4JdP0z
WsgP6BtvCD6JPpltWVSPPXi2DnZwnfWX9yZhVktGWgLdTQn+FFaoSuEmIlU1fm0S
pSXwrP7ibrF/u73DBJ1r/2ShY0CRiUTVzIKlB9bPHJkR4xKmiYs+YMhImHG1e8bc
0AGwlCV9Hnjikj6doM6XZOlgoX19aVsRBX3pAcciCZbuQ0ayZ3mi5gz0/QS/6Jvc
pYv7j478rZbjsKkwhKo04sB9fJ9mo+YpOxjp/zFM1ENOdlqWdZDeGDq2ti1FIfAm
6u6WfynCXhlmSRtQaJ9AeoPBaIMnRxlFgtiyWZL3FguzE20WJpsU3HKVUZBYCEsx
ikB7pZf98AcepoOOcA8SwTh3dWvlc/L4I3vEZDmZ+zgTJOI8BUuOswGGZiv6JBFG
GAopNocdMfDCMdHexcfjgXqqOuHPTxqNmlcithwgwvSdR5myy1T6x4CK76zVy/37
f2PmLPtWpca1Z/qaP9mHkYCs/3BZcHHFAsp/zodk1ECMTRNT+cmj8BtbOOcx7JGz
4/Sku5AQfts71KzcRtO4cCDpIxM/0yzbpTKzk1Ywfxgna3nyQKI5uJ2mfBVK/jTF
qDB3i6PA/U0WLFtpLPlbrDBRnvPQr8gv6aRuKp7uDqCH44D778/ez3ISR+3GdmFn
nyvJg+tjMqU/U8XUUl/v0asXhNkuoqiM5Iy58H9POC6cbZ7ppi9v6jg/4+EjhQdu
jk6rH6fnut4S8t2zWKSEBsLLEYhywgUCNRUpNOI/sONzleOmdX+twBcnNme0tSyP
leIy0mcntJFrduA6ONfOzFgIi77+YfkMS3Xi7YQOuutAxXbuxeIGHAofNlMkaGyQ
Y09HwbepNDIfVGeTbHOx2cVJhIH0zbY3FWaUYP8AAARKVH074+OdDTWVdl9rYr4W
RH7u0T03f8/ERc+jdWuc7Upy5XPp9QOqsu3/BsgHretvXZ5ydTWx2ndnXFtjjymM
buavORIEwHlbY3N81/SOPwqnuEgToZYOhiw4mSr02bfRS2Yn8FA1oBU3qS1inSH9
SKAmoA+uI/rRzIjJceRi4Vgn6GpntBJXSxcJXY+bilY+hpJaVpZU2+Z1VX++3eNl
eJjglb1g5RfJAqEZaPhytFKrwOl5XfPfWqeLV53vq+PpcAwzUJd6PkGyEZyYPlZI
8crNSC3vkqWfUiOXUV7pZkDKh5WDjmFMGeGVN6w0gQRtNEj8CF48mvuKFPsFMxHx
A4gAmmT2Sncr3yD4HUiiiCla1QZ/aRh/d85HIZ4VmR07adL+Bo6cXjF1+E0ANOcA
V1wPj9+fRlEmxKv5Fz/gkhhIokqCByXgkW2KJn0wMdx4nQ9ANxq9TolHM0LIpxBf
gqSh7dRg5KRvzmJY/M6tnQExL0RMSxc//GYqxfBPNL2gzqVD81aiSr5bl9utl0P5
t51Cmwuk4cc1aqT/hHkKnD4/ONs45imdE3nrA9Z0j6rlCZ7IYt/jFyvXPW0rDjzY
483thX9Xu7YTP2sUyV48TUhgh5sPl+wEg9xNTAyXUrpqX26c2RT/lUgAGdYkxEHi
dfL73Zb0X71w7tJbnNg37t/Wp18yqJ1/27KeQCcUnrzK8iJU57UtfTx85ZPgZeNt
lDH87dS/Ox8gdGAFvIqLjwXQ+7pqDrecE5Y3QZNQJp0BcuRxX6ufcByrbga+aMvZ
wpK2cxEglqz0IwWBD3gZnNf4gdi2EkwxGE0Bw+A9N9KeYO2IUzWWQVhCpoqMy9kk
ozO3f4cTSjb+hGS9lOMx94k9CK7qwi4ISy/RUBqtzanSQi4Xsc8KpzP+rLFKx5g1
TgcEc1+0tM6yT9y6urNzBM8KXWCxrG8+ZJVCvtVXxKaRcP8S23lIj975GgKhTknw
wvUrYgnChhfYH8Ldkl5FLp4gBC73Wf8RdqsxVqxk/WVGyZPT7iX5cAbsAkCRGNjG
34gTyffGmUkL+uFdbPd+ufobc6kJocl30k6iaBQjy3nCXuTKPmwBnhtEDxXHeSDs
k5z0X3exvNCbKNgqWHCRKR/kGjbrUWMnCoomAwrofKdjlMUNIduGV5TXiBv9nz/x
NgGP4D4WQoN9NNbylHC/K9u1zvniQKXx12cYgGf4fSqcIO/0mWX3c9WApj0ruTp4
nyVrAcswxPirWAtQFdKgW1p1ldhHPKLl+QaD6EGrqZq/A3+8jcwQfiYknYovUfsm
1pqWiJvnzQsi8OfcVIWoYqW5ZBWrlJIAIieDcjw44LylhIDHbPw9DJQ0Q4XYoEaC
shG9wxiI3UGJa3DNFRSlJmmVfKvhHqZonVu2jw1DlksGBopoJNPrIg6NvRqgctUk
Xu2Xqrm8aq+mSvv7+/Bmwfh9SUjncL/HramZw+jUFl/mvA4wPBDWmRjAz4kpqWbo
GQIgeiRrARxofus5B/TAbKTW7YL3xBipIywB4BOUJ3CREi02MBPQs8S98R1iu2dB
psaemyK9ICwwsGdI7fNUEKvV3T+glqdn1w5JkCe9k1Vtpi37pwu//VZqQZmEe7RJ
rQjQ7Bsclyg2a2QRXjuCR66WymKtkRxfXplLZOV7LkT76SwxpvcIYwFEXeKJEdGn
O+p0UwtvdkcxRyvpwAKdUejB8EoAhE9bqQelEKyKNqqvysUiI3n0naebuHZBS4/e
Y62+DQ1gW+jMtKOT7+JLxDtdaz8FQz9nOV77au77B7cbp/HTSRDXykBLi3y/bQ4f
knZtZxVewdZufYVCBI1HWb+x3/WohUsFRSh742sr8nFos1szheg0TcwDiOX8HPC9
QUqimE1clOgEdCg5zxxbvn4jXSbr305VpMRCkGGhNLeHKUkNfQ8k9Bl7FSo/wviy
pm6/9GUKIFCnW0SeHVjBmXhppTUqpxH+wvslriv4aO4fKwjWO7poN+P5RYmuyx5C
8gETYG7P+2+qdE4HWbgasb8dTHJwMrx7JKePmdii43MzjnjNFbXLNVZwUQrYcM1k
XgyZAIALeIrjJv/elp62f+Ash+5M2mfHey+tpK8kgmxFjyvFep0kyRpnOXFsktmj
Tc6zyp/vorF3wYQDmLX8usSPYAddDTrrhVFidunaFISzwQqrSOdqRzVQVooFDOu2
8l2v2JAxONE8lLcNdk8uyCUxmdc1zFWarvTKiiG0UqBPKnNvyTnrhY3i/1MP+X+A
Lvf/3SUnw27HI0z2QAkIIIIAljmtAQYWVHFib/h0DlV/AvMJ1P6M7UULZSzaIdxk
ZmLGIxHHZMTQ9gxO52T6vR+9fgyqQ9FelFrOGrWHel9R6IsKL0fbT7BggdVUNKyO
dqZEqQ++Yxvwm7+sIw4RD6Ri8e1iWUX40vDF7wgTQaIJWTyQFAD+fMxMWLujl4Ca
83Qsq5gEtQeZ9t7hDGhfNLel3izSzr2ywEya+lPIMbQQYe36sjxK/bdswArSEKN2
JVUOGpxZYhB/thTynrCZfiuHLrzmrjDYACH3gCsRS//nu8ST79w9Hea7ISk8/iU6
Nbru3I/0mAVMcegsZhKk1gExyyjfhPLeTz0GgIph51sTDXPKVl6BK+ecncW+UuZS
/Gxa5XT1LFj35QqwafVXXSbcKStvwD/8wRpuuAoDYBuOEV1zADSD3NxK/7VD4q3a
JluAozjauuxkmW2fHj9V80jjWqszRHU1axH6tzBbmdMnOEy+jxERVAA7lpxdKVfT
zVlGNiNeZ4iVSo7CPfto1gjT840txQrd7fZqJ6NI2ev+rf2t7ac5FTOD9GRb/rGy
VXG34i+cLquZLFIZzdzIOnWYJTbuDUNh+Z7gvbzMsvvW8brWv25s+WbB6aLZ7inG
kKO/rEywXQ9zg1XCzLbfnUw+XATBlZASb7ZuO80YTob1jRQBpBnmA4cDNvM7YbVG
5XIzV8+gWz+ftJfKPo2VtZSEyW3tYXwSGp2DpmsHE095aKsMJIJvqZ1rLV3xbzXL
Z+Xyk32+Evjp0ip19rAlOppqikC6O7NysEQuAQ0rgfNZzCJrKkffngwPWLAmthS9
qFomTJ5Yzmx7YlVI+y0oxt4nCq1dD5s7NKjTlT+h7s2WiQTHTwaShfRg6Kk1S86K
jxSzZ4vzwswotWQzpw3IaEswQrkbQ0JRSZAFc0nu5AeooWmeA/GK4R50EeoXYGVs
5QA6plsIDdWKnAg0HWlhmMomdzDSqEucI17xtUo0aFY/6p9+rWXJgcqsgyIAUOFn
bb9oTkndXsBPpSLOftyIFsTaMnsEjZradzBhPAu6p8cS+p042EoR3PbDKFj+q62W
ZI38bo3fPTUdymOq7a+FZJE0zchKkAOsjg5GCwi0n+f1ySsi8ZP3X9Klh1T9b+xI
u4SsNwvocmet7Un2Yfr6G1j+9xwS4ZFd96EFOWPM4cBMKwfFkGVw+iyKoqizvWCf
Q5Zs2NJq01qxoAwHA9UVcD8JaiECUSzUtEfmmLruBZoembsTzgAoZ/1NxNN6NP2/
V54PXgIVQuAOH3HcVdT869FXv+3/tw8DoC4aKwoQPEaBFUaYvi7ZWSS/BtTC6zZH
uljXeed0hVBwSBQWD16u/U6rr8kS3ZODNh8DsOio8MsHPwgf3MdPsaiFavrDtkGd
i8EUm7nT1MThaqU0+VwDKH2badGSadl/Igi8niQFL2InGu+bg6TJU54GFUPCwDko
M4DVUdDqJroHkDK5UJzCjTr7dMuUopi6I/ju54jQs1amlU9YKqrn8tqMugJ2WL0U
ZXxMo3iWCDyPAP/32lp0N4kFOpOU4exYsUSm0tcW7OZBUxJKKpUrTNjVEQg/bNdN
BcBfN5A7cIE727xRo4o6SmrUtXxu/QFA8TDgUn8v4vdSZUHToOfanLhzznQ5AJYh
A6fMVh1g4xQ14mcQimzzur5uMnZWz8s8tPWZ1BV/DElTVkUHAorXQmXZx5F4Bu0H
jWhNmjwYCFcVgx7CaakmD7Qkkhe9xSXY74cP21y0yz1jU3FESb0BBINpn6DCYEWq
mzrDz4TyE+wAA8VdUFBIMEQ0dyEwlPBLVGcHpMP8Rsgzqdk/k6Oh6pPA5JBzCR02
yjadWa+i89HZQFvGTsMPq+LKno62ObajcJqIQIJvizFK1Nk/i5iXQELyWLD9Taxj
lHDfuCkwYG8pnzMgcEKI+nYX4ibV/sdaYQ2OOV1MJ+TpTMDY+wr3RONhP4AUbihw
z29T4VmkUuT/oZpQWZYrR6RWsHMBREqDioyFEcQRQbQEYXf9nChdpZGghwAgXBky
JR675QHpYPvPoaR0CTWaxjDnDVBEB0Pfdf1thUwt3bBn9jRw3sZAkwRc5/NgYao1
I4oqFlGWMB73cwGntzMyfHWthxVWeuHDjptdwkNAqWnpJScrHHJH8v1Sj/vuWTs3
Mbu8LecsCPZgQ2LNnYbl+ngc6WcaNGhOgI1KAY9/lPaYZXQJQ71LGBA8RPUZfk5V
pxSZ0w+ikmvzNEb+i6mjRwbBYiqQeFTmZMh8Mw+by34DlTHCn7088vSeUeklHC0Q
pZ+p5fkUYwri3QdGLeOOxTlk0iJ01Cj7QwMorCYQXSCWDhupamIf7Ai+ZLKtq9b/
natrNEG2r5nYujPSZQ4ec7zVM0qcVhiHcNulpHrJNNsxziWNFtPFJbKiX6NvxxjE
Feh9o9kX6pP3jZM4ByoIKc/dQcVosnd6Wm/t35LTJGz0AN3EG9qfQO45r/xsAx2G
BYUzHzKZm+YEvIPH3WQCl3Su4LRlV8/8SL5xEEK9h/EuJRvGKDEVer9e6ceL9E52
98FNQ1zl4DMMEG5lW6II4xF7g8kJYj4mHgAt+jOaqfIA96uGSKodu/bpulEyLvrW
gS2AznG3QVoAyiNYSYhqsUjCo2NW8SuLJeI7OGgJKdd7eZiLBv/x9v8t3GUJGSRX
lNubiyrzCwCJLS9ngVFJFfKAPmm0hQp5q4u3MBOV5Q1M+pVv69WkJaNl/Mtmk92F
RVkjPSfOw1jM0TCfIXfKLg0Xryxcwau3Kj9i6EfH49eE6n7kNI1+u+5SXHgxsgYd
9KOK65W/wNYNOA887SyOBvwduYOExkPDfTRLc7xjFXzYSQuJQByNGNdM5YEw8RnQ
Du8UkDSEHCF0lwDw40qRWXIg0KLxUVNO5Lw2hka8ZIexx9rWXcgyGeycuub6xN5a
T/+1f38GsM5A4fPRFPGIdGRBRkphKzINi5FUhRa9bN/7v3uvsx7PIrX7XNyHt6kn
qOus4RgFVSF0hXJ6UWqUkesRiYFzj8/0H5jD+xs7JfK1Xf8Q1Od7os0ReAYkQqAN
x5aHgbPXmR6GJ0Sl+BIspXGVjebFWVtE73T2z06B9mFS+8hwxrt/CL28diCqW9W7
BaIEAmY3IVrpxhp3/eGPgEh2HG4I54Y4QxOf6ahQNzNgMae+h7JbrfW4jaQjfgnO
6oz47T+0FqF52hU9STTd5mHtTnU9BhTb7nmbxAttQOc7klC3qGfwYU3xQgPMtN1k
QnkRk/eplWDzfhnDI6aPtweafh66cKeihKAN1xEJtJZIJfKoaZ3X6V2h3ryKUQeB
vktghwzs+nEngTYiqajH/bXfah1pH7RKMQKlkbxJWErrQaQIF1UfT8EXP6hXvrGb
ncQY5dBO50IuBBGOH5y47B4iFeih6Be2ZXYdIj1lEp1+N902Su48yEXahFZ6eGKx
/W81v/ye1YfA+vg0Xr9RZ25fVF2dRWthwVeLBqdwMj0gCUr5WnvwijZoyLKDB6u/
Vcbgl2TWBqRM1VFDOV/vm61h4x9DguNRrLR/BwG6W788fHNsE6fzZPUjzE+TYfHY
i6vOYuOr4pBoRPy07s8pX/KqjooVoeZEJMSC2iEqbxwAI1lgiWu0+GlyI98xGnDC
YJVYm9n6Ug+hZOagzeqQIKB45pTZ0mZi63yQZl7Kr2uRbyCGYo4g5I9hknJubHIR
BQa4UKXna7uzrkwzMs3IDsEmCKjdgBVGZQRwAZ/KZAc2upEXGkrNzJaJAF4w6p04
oBb6wY9KQn2laOeHWB4RC9ylgKXYl0mqOayY17shVD7FudWAS+aA2ihvRY2hqluv
bdA5miZYE6GnvPNZLgFdXrpdC/UhNiaC4ku23U3VhnJR6VLXb974M5k4ofmhtVQ1
PsHDJMkIwlVTd+mPslkO7PoP7wJGEzdZ2fFPnvxXYyCQzbfg13vycWz94GVyN1Qb
mrz0011JNTBv+6L3/V1EriwWsiIe+7lnTZQV6I/ApSeFdp3h6c1JyK20jWmiSmH1
jCWC5T48Cs9nOmag6nYH9bV8t9ZH42piiMYlp895RvPBUgsxX7POBiiR2BKxnB7Y
1hp1b1RWffaZ78Bad30XD+6Kj2IbysIPIFyX+zacBHn/ToGzOZurBMZ400JTg1+u
Wj6++nloAhpNsRvTu0XQRUQJaY2WczjwD9jT8awwojIGd5VICM+QofEiF7rSeF6e
425/RNDYeOiPK7c2Ff2Z1b33A0ZTG+vFMJGsdW0gC5ZLo2n+Ci89WE7zujjvLxKq
HNXXbY3o8Uk0AMgrootMEOvkiU7YqwG5vCwP9vqQF+QtCYU/tk8AI76dKPh+fNSZ
xfBXEo1nO/QRmlPYSz2U5fLTRUYihJFax0hlSu45C61xuHWMeSNrLPtcLxrbqd7i
HpVhkrmyIN5llARQHeUJquvB9E4PPKuSO918wMW4x0Oq3E8vUOaIMrKVTy7SYRKN
u5yuXObivz/WVQSjGkevqFYL6SIMY82uNeKX5Ne+EsJD1wSe69fOsa90h9yQQQIv
N8q8zp9W4ALZnpNODxIlwa5pazmF5HxzdPoxevyOTmam42iuAfyu4ZLIUw9NZmyC
tfHNIoIBaCTsohsUbstvj+T5kX5gwzfYqqnQx4Tof89v6m/+Px8vPcCb7n+R/VME
I43Ve7PwBtnolslmN7bOVhtjvql+6FcFKLpy3SSYtg9eaOxTGSVpuceg34hMZnmZ
aO9OsNAfj25ogQFMutp8xWmF8OvH4DCLBwOWscxe6cUcJliTlMPhAiHHCm4B/pjJ
tMJ+DO7D0YvyKC2ZFvJLUxbyy5J2LcI0oeJ+v1giZc+uQjtCDmqblQsTjZOKX62f
E6nGc0PKM/6Qoe5Ij1j3blz6bX7XFeLmY2SqPRhiQAsLexcKdZT5FVd0aJmQBfbH
yecluZg5gMz+NY2w8z/woWGV1w3syo0L47HLTTkyf7j9SXwUKQ3ezIXo1NSSL32x
AEBeNvl9eP2orbMuocdFncsc2s3lG0Y0sNb3Bz+AAl+WryWbT87uzgxMjGMNcC0z
ApiQUduzYdWwDBYMMEX1L/+g1QEFbmEsM6cOWNQlZ8C8kcLVl0Wts435fZIZK39V
+PWUonBZAbHcN9NzEROzGGvtMXNfYzX9vkGUgffIHxf9bCCpzxOeILvofNJzdPcc
Q+xMMX25aioC4DxJcIcdVLQyOeaLZqgqzV1X3R1wzJsYHFjjE2u6vkwTMXzeEh+Y
X41oK6AoNKrkPw8kEbDDKdYj/Lmvxxi5nXn7XLTWh/UfmdXaonDjRTtQVYFRRN96
Q3LB061VVFZnlHAtyHbWAfbFZ+2Y/pQmLEBHAK46TS7tpstO7YS/2egMa4Ps+YKC
6s/zTo3WyMuJCcfUeJOjq7cRTWIGx/qcNrqcVihK5YfGinXUK/4IfmJxLW5ZKhlz
6M5guK/DsgcMHm8YcTBRpweMYE1thvygi98rJ3inCU1FPlSaM9Gc0fAtjmaNzUru
FZ/pAMuHUUjpF+CRz3YGMtRTaqATMxAnplGpwdoxO7qIK3Kzh6byO2veybeX5icb
8t/m5m7zyKWXn6vCif48rl1+wPvaMZl2i+c3V7KWFYHl5UzcgCmhV48SPqGL4hko
Z8EeG4zoV6Je1HTeD5r4wo6xReSHt7pcVi9V5DE1KBsOILLs4oWvRJ+gelEmlD9q
o1ickGNzrQ0naNPVms1sA9fdgu8XSUz09UelNo19DkxLpmOvYV0Ad71vvLYWVx1F
k+fX/QjtbDPGBGw62EBSuKRT0JGgmP3EcPJYWqO6j7/EGG4bMY6e5MB+2qodulUw
28P8D44oJ9e7rdZuiAWWA+QWNdgQ0vlhkZwli6s+hynMGvbsbB/579t7Hzt2Exha
ZcWFdU0cHjkTXFrxWUjK3lLphMthbo2texr8lHEwZ+Za6/geFiKiiJPFiD6tyzep
Q5wUZ3HCreG7zkIa8058zImnhArfQRcadiyhA6QNbTwBjVi0UU5qYb7uW4RF8wdp
UyLQNS9IQiDW6VEUTr04Pj+zfFaqnjz2wAYA5FXuvWKir2lqLcRZYLC6Y4s4fmlh
20vBJnLpQR1xi87y+fSxW/AALkEsWkcvfKM3V+fzrzrMVFE3MQ6HjxJeEHWPZLyy
hQtbgiRAHMayvw+RnyWPGeFe2EajWfr6iQXrfZ9Y5SYdrOB3dkXTX9y8gJUFu7fX
+P5kIyUc1z7DszyOw0MRy56fd9GZgND8Np1OqtnPuFtd4TsQcwfS0MqabcKPdIsE
tAsIOlCayZDpPGUcfzJCbwqHPChsZrLAbC3lHPEhcU1XAVRjNLhcFN2AKA9WpFgy
xPyY5svXVI0j0minudZhy43k2p1iWLkzBnqOHD7UMURbThFgfXXeRgHpn45V1dyg
eYfpoaq90CsCcPV7X0/8awiX5NtfLjO58pijAsnsZEgzMWr12ZT4IaZzV+FMOj57
ISHd7CmzvPn1w6bcQOUfZNJGbUS9C+/RIjQtJLIdBHb1kwMY2gNFYgGIh1saCwed
n0gz0w2tZ1PuQydk8238e7FHkd7kdAyf+ojr0MPwnOhfpCRFp4xOZjNCE6DE6nTM
uDi7Yf919k7Kn3Ahuqk5RsdfrdJ26IhWdHQriR7gK+Npm5K3yH+qwWSrWiVCLVHt
sZ9vZIE7odkkUx/mwb9hwtQizoEKTJLU8y2g/p6lZx7U25Z/Dppmh2FdNXSfzzsS
CyX6iSViCn6GPcUDs1d4LRoKUvdyfm06z4sBQG/Bff4KFkSAmSmQ793QOSqAD16W
QTc7mKx7TGQT289zsweHvatkbhDQFR/9hIMGWHM/BhDOKHC0nm0OPZdPp2g7e9ab
dviD4OJx09g8pP+/ePWOyenKBqesUBynSvAJzaOXftKXUQokGb3K6AmiJK91OpFx
ts80G/Z2pbiw/o4m5XtCULrAnYyT4ovTZeU48IMKy/4mPKpIpIdS1/Fs5uhQtDCU
/rBCjI5d/7mstTzubGd6pZyh8k5V/38burphySr/GyFccGkMq2OFehYmVnfRl3bf
DsDxNqmzOn4GVRaNU1h+2JbhHFCN+kKrFupKWMwHgmBKJAalUf7/pT/rr7WU7ajd
XM9W0S0axnlqoPHo8ZoVJGP+AsA4dydUvbw73EYIxjVu7RAUTYWT2qKelSmm/mS0
8L8biaymWsHZzs96BHWZHlcWXlj2X+9GkIwNQmxLqYywJzhNt1b3z4YUQHDYE7Jm
HvbGpbmj/HsjjiccZvpeBTW9e4ALHiGDM3OfOkthMgEkeFv6M1oZY7tf8/2+f04Y
QZdVrhXLPrQ+Lny8bakkIMy64iOr2qCQiN8cRWji9f36rCN0duh31qXmGrOROpwK
vjciUYfUuYboQioMrM6s2r+g2K7rXJPvrpslMX8WLfm2hL3bE5w6lSUYEtS66fw5
ztVpV4GrtqjY8T+Ioa1mwrytToVUovYQMOVqNodmv+pm4a3gsjLlI/Gpu/dpv+G9
6QPMmWuKmR4myriPzo+8h32nrnJEQ3QVL/35kgjHvhOmkwO0bCHJ9Fa2xuA/Tmda
ikKH3AqIb/cYsiRajsFXre9ouL2Sk5/GsMLK0vMceBHEAFFNBNIpJK0D9uZ4vKFH
5WgPE4o7vt9ujjLoOfbbMQoTDGzx15gz/cGr188Sv1U8Nn8CnR43bKI8j6KkxP7g
dJhqXPbYMUfjV/JMUpiHAqVRBwf4qRsnQWXD7R/kTB/6ngUljTu9ey8VU8tCq8Ok
15Vjsr7RNRoXcCEAA4M8UdNLAwEbG0nS269KcfnUWVAKCTa0fwRNIKhARHzetGDT
SFY2/v+xsEuAE7uulpmqjMfdhd+FYRNgxhn93EDjEzGQrXw9l3BzAJ5DZRjiGkN7
CCczF6Z7bSHEQHQpD3xdZXfyMkeD+RrtU2TLeuA4d2usRwZlQz7jDyn+6jV5DA1j
o3McGecVnyYX9aL9AMM75bILEy+jYaT171i+rWj/TqWDIWm8FEesYLIysLEEupKJ
Gl5fnd61eWhqZ2smSBTYgCDzqAkxS2VAKZCCF3B23EiMfGVjE7/2DdjTWrVS3ch0
b2FMms0D3RUt6UoBxEvRRfL42DEpL77v0S32E9UkmvVktJOsv8NbvTnlqBV0xs21
XdwlCdqIMvBH1+Gus1v38T2CjCx3Z2qe2hifUensJRmO2RVb7Q5WuHTGbXhYwb7r
V4eJpPY+Y9Z0neUe0Bk4HkHO5S2lFLF7SKtObs9yVPWxoZHS1eE+qvaW9gryM9EL
hySSknUfpugYrQ6r5cc7yoVgDj5xig8eJL20WvH+ollCkU9bwTPjhThY5VPGmicK
6buzSjyVxBEE0pY11nB7C9kXRnF0XQnOkmlrsw9yIEPh3sp909kSEGAr6PWaqSBf
XWnnREDZdCbouWvFwSfxTOGaxrNFJJuXSNgWRNvxYEDG+JQYvrgJnFJARdjJnarc
xX3LIkgK/s/0ju1ZKxrYXnH6uts29vdM2WsYEMTrwZc9T3JIRRJn5tKfyHTzm8PO
Y5zMMm/V1pGHUtjl4zVqeHM9AWULl/Volf5sBb8yc1z8kPDW5j6fE71lj1TkSLLr
wQ8qJqOV8JQafijGkxu5q6pe3FatdJdlR3ymHPqcmVRwORRpEcveVendhMVPVPBI
XH+f2/3+9YBIedXluKrwUDk+Cn3+HqeLrIROWBdfK0GnnApfngyCCNDKCIARmaFn
/gG4mJgov98UpXsXkfxGuG6Xwviy1ylX+WgMfS/NJMJIFNAPzi4DvHTomJ8Zi8lY
L4+k5R8XcRxisN8a7KoJYfjtkBLogsVVUuEVXq6LOaVD7zggReladnaewaQM2END
ooJ73WgOD7OFbMJIBpKDbtJSqkIf1rGXfm1X7WyZn+8cSwZUUGhIkHsKQJsC5gH4
5TzisqQJb+0BpRSgd7pwJt6FCvhY+7moJ/Hw7ehAMLG4rkG29WydoSpCpyJ/ptu1
gkBTWJ7XENpqECvA5A4RFjmZipaPl/MkeGLMvzlV/vDRD84XUSCqNCzGSFtBr1ph
M3HeMgvCUrEytT6mxV6QHuDZGgER3Qg5QYPJ97CJWPnCMV/yRAIEEmDhLssDE988
IiZHVwP2AYyBpnHM+TnA0QPJ4P7rPkY3nXwl8YnV3nwNZ+fT2f5lknU1zXxGaJkP
H1IkI0kI27n1q0Oa73tOPkWyAeBSxIuzfUno0bl/T6cAoBSKdPogSZbd5Hqpoqxe
N9YyG0GjTUcD4oLbeY9DlbuP60xErp9g2UExrpISNc2f8nPWF7Kb70Nk4nWXmrpq
GLf5gAGaeu1FvFNi95PVROD8TNBvEu1VP3IhBMeT2U27oN+Hxj5h3J5IWy0Q2/7u
DKqjg4HH5MP/NSQg7qtnFmCykjoIqRJw7GMm8WhYYHZzDnsm0++NLz6WTeVnUxBI
9lR3VaVFVzLNSgJFeLuhfcaGrxT11T9u85qZXNoNsW8UQ8hL2pIpxE8KtvGLj7q9
U8T98tWFgOdR/rn5MZOSlJmDIQCxKoLiJJ5SC1P9m9F5Fq/8mhmlnBGmELBupcr9
Go7vO+m9FrDwirNeEnHuRwuatDf+g3/e1Ku3ts5iD/EWrZ2LY3ecaUIpeMXHHXhS
ZIvVg+1ui02CZEzpRVN8g0V+grCVFKB1IKXzrNfBRqv4PtJTGUZ9bqzTspD25/qq
6UFd+Utbsdfdjo5vCQbKessm5tnSOIitbCyzUjFNIA+Q2OgxHCqchF04EmPZH1Dj
s0ecjqU9GME8ZhA/AW/4xVkn2EsvpR1I+K1ElxRoFp+1vQlCx8XelIQV2uRXH183
s0ACS9vA2LvyYpXvA3dLvINsmzgtSSpc/N+VLcsWOHcZzh7RM0BNO3CQysHrKuIQ
OUXmlPpOL0skhn4RASMQhbfqq8GO4bRaYUEtlFNDgTyqS93U63Qm1YhxH+kKkHwI
N06JKLTNFlmWBPLx2sXIxX2EDwD5++DlUz2x610zjCC9OmpZr60Y+bJcSa1yiSkW
LXpi2V+JMuB0lTZeDHK6gxxqE8PujH/MlqRNTv7WhcZNBGi95uk2sBFXgvwhh4Fi
pGJVUr4PPRyD73qx8d4lkRwbheOaeNZAJjLsW/Fw5ISpcMvm3EkFqFJs6zi+YwXq
AhSvM1GPHlirDsx2BABh+XLp8DjTz9AcLAgqXtMvKiIvAyH5Agfe+5UDnq6XzdmO
Qt9noT47zCxMTMf4AUJfazDkHOamnHJRRh95p9O8E+rBo5yyQh/XGoBG1lXMCE42
E30bMjjqFx3mnhbB9wixMbJqAY1BYAwrWyCobeeSUk0zFI/9OwVGPgWsqmaI1H9Q
nh2DVmH55J5mtyfqNjlP2L2T61e5Hzoifhk0jkXefo2hZusA9pyr4N9ncal9Noxq
eXT6TzBeulMKFJURHfbzYoqzhqjBS19pB5a0a+euVLnyImZFTCvUzOtAxQLmFqws
t67KJSOsaW4hiaSPYe/vweBIZTXOE3e24n0w07KB3gaGb9Jlyv0zrMSmxcY44920
A95OmDohKCYqk/k1lm2ICAgcCjAZr3hXmUzf9ucf7xunxjny50m1ZOtyFahlP/CR
Eytkwc2jnMMtryRr18m38cs4Gyr3zdX7PfqiWIDZJ0al9xWinRuFePC/T7jBC88m
cYol8X4G8F4I36dA0YIAB6KrGSV+61UQlNevLiyaTOEkguGdjp5xHL5FBup5PYC0
8Aghq8a3dRlSHhlGWT+E4nO+SeJC7kgGP/T4ew+aeCZA6JzaQgRRRadZ1Qf/Q05E
b/o4pShi2acCRYPMv46qq67EBj2LDC6XywONZSdPyf+wEWEGmpL6+bzK3C308OjG
2EihN1PFDmNKLQGJyGkMZfIu7kh1a1vUjhiSFb+U41PvuaHXI+h2VFTuILECTpcK
OxN1xh6QTC+iVuqK/5kfekDFCDVkGzvNvyuy/QP1XANBCV6dZHE6f23I+6UazDW/
dTXzedFBC4pPJvT6qwI3s1hFkskN62fZcPVH9h4sCntFP8gJzxlViwRc9Tx3pX3E
wiNd9u1hiENNBcMfXVfawt1Xo0QplkYBtc87yzzem1aV9+yyMdtBckdbTEsrBQOQ
BCejuxxZiUwamtRhO0a2E+nbXsaBkwCZ96Vy4vahEJx8BzS4PTGO/RS4sjwWWW8f
vW4qxJjk1yJ+2sOwWUg4I4PX7WJU0ZlECfRw/Kwj/z3aIGKIVnoEvHnD9hufRy+9
Fqn2K/AB0gJUapF0TGaz5I7UGBXG+nBZZBnshXw0eLxhzFHDcYdYcEjd11Q65V/+
5jAq4kfJaf0sg61TuwIxkFcAY1LsGATiGNfZPAg/8gxBL9lXwA0zOdV+EAGKpbxG
GFSTvIdNWC0bCh85ykq847YL/KxI/NfR1d6S2rh2Fqt5BAAobIq/hvzNIDoJFYKp
KwNo64eD09zOT3a4nZaBBom68eb7gcrZxEpka7Y/yTgZSk77I2ip+8TX/lVipyPp
tYm9X7y7bHtpQRVfAy4z+1j0r6JItE6TA10v/4l1HIPQNhdBppu5x6JRzSiP7eb9
h/j2lDb6GzOVJ7hkHXwv0IhZwvup7nJX3jcFEcS7GecPQLIrOImuf0gbxOv2gMVa
3+X5Br3OZr6RR6UktEQWu3sut4zUfu35amtGBb3uvGJmAYmqzg01XVaBcVdLczE0
5NevIl02IVaJZZxX1ToC/y9hbkhW2wU+dpx2ISQBGuBolCGwfilYb6fiQ0pS4OdZ
wv1KI6XUvg+Wlpmp2gi4lRdflbaBQk5LVzt/uj1FBFaIFH5FDfctrm0+jpqEdXcm
0aZYKTOnZP+hBIu1S6fCqPdzZlWrx27d/xLrxNfyAzMnsIbz7Gn5vnvP5yjJS7YQ
wdDMYtG6rQKKXsidNYORNg1+JuIz30GQcHX83ZlYTxSDX0TenM05VKvf7wK0xfRh
0lFnm4HdRzjqR6CrMpTnuay6VS1scL8Q+G+F9/czhcUkNB4+mOLwyvHDR4UvM4WO
uxAaZdr+1O/zAcVYP893nS4kxzq+L7wAcXXqBHpOupTRMxPU2CZbLtzg2Hv1EtRk
knfZCdrif9JMEcQgcyUQQC17pxyPUcP2Yhr1NSAqYticnGwQsNBOSQjQdCUnQojI
IKBA4CfOxrUJ0y7TvShdbLnTm9AMGYk0FR4RgQPUsK1u15q9WyCdsPSo0QBvm7pu
9ExVD9TE233zxFJSAYH+MnhhZlWRkmKhEcGhBJRgwacReED0mBOjrHlxLuvStLuV
hHMIKEtfvbC9mDXMBOtpSSaOg5fP3KLTEI+nls97esPC+g9HaLB4jFNE/x0x28yA
jsvDqOB0gNnp5yUxYy903gyhHrFZiUyAjHiy8PZJ3DHvVq4wy8nfTLKhNzln/NN4
HWPfD714S4aBuZiCSwZMuuJqWhnkk7GWo62y8ADj1qlWkJEOTKzx6E6xyG7SKpvB
f4RQcrA9TlapDzrANhb2PxeV64kO35wMxAtA8Jy0kumf1hOICF7xLMbVHM4edKJ9
2rrIQIxtNmGFGMOZv66Pq37X/1T/kc534caIbLWPEarqk4SLtJnWfxtPFO6Mqbyc
LJHZB1jYZuXik+mMC4zwS4sOUVrQMyy43ZHARmabLIAwqSTOb4kFYTMB3hF5jAIb
ATq5Ljz8RHRhKQf3FxavkhkF7tobkC+p0QGNfPo5HvZsXIHZZwpYZ5MDf2R3M6p2
544D5MThcbd+XwSJCDHKiFSASUx9R17qQy/n+Ss22y/oe407rXipAcCl9/kSzZNw
T0v6jX/zD6eOVR1ScrGzxr6XQoDZmCarE40z/SLc7RthbhFrGZn8mrRw/5856guX
PYxefUw5YElzEEA+mcuDhl7fk9UbMTA3eCK1L4LvpI82JRSV9cwqV8rh9ux8Q7Ph
kphQOQ4St0qjeYZNd9aWHYF2k3v4lBa5R1qWZj5GT+PE2I58lb+8CY3fS6YllvZB
Wj1u44HnGViZsYzl1X1rLBDGY+KT8e09RXLbBXXe6H7PfNfuzU6pLETuuYcWeQiL
3uGEAD9kwAqU4vK3R1f24OBCm/2tcHE1KjscSp5FhjvMLzMWXrQ+U03PYEuvgwQT
Lr/mYcEurEqTsE7gvIsooTjbn79RFRngo8TJWVq4bE1zVj+sQf3nq9LbNUILfE4j
Kkxf0xCb3hN85iG9QriaKiqve4F8XRPjguEQ+Rsl+dZu4c4FUuqmJn6R38xQVkwh
RPNLvYGssodkPuJ89jEQr1pivVw0VZ1S0fwSMk74/ckcObqoqCkZAWAQq1ADAvIm
aEahWYb4E76jH+ghUNEBW0mPybHXrVs2VFnWqfxYUDkLHAcuIe9UMW47eGj1hACo
hE9kkx3MVzeSa1vcit0/C5JEm8VhSkUlowfzS/fUs2032W16WNE9K67UWQwf0Zbb
4UFMP+R0Rhd7Jziull6lx8QV8bDNlyM6+EQzG6Y9y+xEqOIiTD/hbT2KMcpuzsPM
/feOma4kJE88M8V/XPzJXBAVMaeA7lKsNt1wq14RKscVP+UUh/Cpd5x++dIvACtn
ZOvgkdpfKOLMaPALD4vNh10hiq9d1OuD5tSsSI+/c85PUN2PFTt6da5BeqBOqhmy
+dZi3iLcrsyyvkws1bKgQrNwdUu3+JGTGYL/NHnVQVy4klAzEijFWMA8p0kVCcV7
cCtGXsT9Z3awN0nWZ2jUsGqH3foljNxDNWzwJ2Cmep223Gm8CUKWXkPvR9rrP067
BnH3CaERgAhJrB1H8xOF70xlmi1io+IUgB4GKwXMcWrYe7LCKdUWRf5Z/uzY8lj4
su30mxmiK64OO51iUMftLyAYeazzXTP3YisNefeMmyESD/BTI7UdZjTADwf75zA5
13BapE4lRP5AYD1IT2B/jS6dk8hpGLCZh3iadxneKpWZ3vqWx8k1LsV9qRNdABiZ
Es3hQewCFevYoYbbBumPzNvBt6LjlhbvN9Vdnve5pd3xLkShAnD4s76qGALdJpvE
Pgyal93g5qm84DLeMeMYI7WPUfXgDnV5FsiBUjDrvmUrMl2J/ltNpW8xmTPkBur7
xCLCUndzOduqxAHj230vn6+EnskQWxYN2TbzVA+79pjJoSXKCtdKs6VprdYYstJW
EN4AZc48z2saYtJtrpbZYy9V+Omklsoson658BHWvy28UcrGQ4M4zuDTbKlLIcQ5
1q1bEKhfZNjYbpWwj/8NTSt6DW+ZwbSK/XZeHzbZ+jTjAFPz/gY2mjuc/KHHZQv1
v0WVSWjF6QeBeAWEY4I+h5fj3m+8XFvFnEc/EKQ9f2X8kwPESoy2FQXt0Vav9TEq
g/w8sCUadPM3223v163p6RmfxAqhvrZWRJWzlNq0twmDKrFdQsXXcL6hWio8PPq5
g63TxOzMYyveKIgtSD06Ho+pBx029bLjqM2Ow2mAqjnd+/NsTBFKNb/PXMGTbpB8
3bQiY2DOwsu2ARBS1v1IQSY37m65xSqdC6LpYI+05ecayYfhXXvTAIUeCPBKlAbi
4zVQIrlMZz1Eth6XdSdG6gNepLc3yzWZ/9TqRS7dLV/iCWEucSEqrAgGlja5ZZ6k
3Szfz2v/xVaeVJyoovybJgnnWL+OH6BL3T+HwKQmTCUyudKElYghzAsWtdmD05FH
0/6VgPQskoq6O/u5EnJrLym7NMe1a2OJb/AwoRp4KvlKy4Ki49wsk4rDSEFFZ957
uMUBTXF74wqru8vZBWFOppaSawmbDjCCCsgf/rEVCgedRwAgh0AHdhQIoQIspbjb
Nvmy4+hk5H83DAADAXD2fePrMiHH/uR5dqZ2HqANGabYjiofJjVGE8syDgyS/N3J
e1xtOwWaYvXvfntxCpnQqUuTahszeq4ep2wT2wf28g51Boc2b3vnHC+mT3ECivIk
shBCDZrov2o10yLi+At3b0ndHkFdELW2ZqyUgNIpJE84oqMHs2JEALM0q0EhY7nU
P7xke55b+L51KAxtAm1/WRb/lPLQsnq/rRip1fqBl4HTJvEeE9gQvnpkbncxufvr
c24XBfZtwiuehNWmWLLsDo3+RH5LLR3AxIwFU5KUXLU3AgbY4EP6OIvT1uiSghoq
6tWNCHSMXMhGDJugiODyfwMeC4OBzVJX5WGlS/9Qei+azAGDzYkHpofBYsLKXEj7
vWNbI55/zDYROdv+jKj2zOK2+UII8jBU+vjXDgJvc3GIcIn7EUPymkTOmrPYGX0R
5SP/HW3L5Ff2Ksd/OHADzW3QGFPZ/8XbLXLADHIkh6U3YWwTsL22LeK9ee2Iqqg2
QLL3ntKjzOrLuSO2pKBFK/UXjMxDC+aMXb9vx7Zv+FzsLbOzzNc+98vS5Gb4dReh
gvi5PAdodoyKNDro62bA0LUEKvTlAfyiRqVPSAbPmZ2GflHC/ioGKxs6lhXvjdW0
FfPCpfruo02cJwnlya+/wvqVkqpIZz8c4cUDEskjUzqxnhOg+Cje0T7FW1sJTa1P
w9Cd0EimUgmlF2kdErFGv7GTN8szEcf2mHBp+w5CP1z4aBmQU1ULnRdq50+v1e41
WHiZ1Dyni/elNo1iz56gV5SZ85kC/AsuiJ3Rqc/nE/7Dvv03sqFEPWICJQ6VMkqZ
TZrAfRjLP3KguhOmvyuuGkYujbjUMzRZSyM3h1PQlo6nS76exThbCEMzqYw309kR
1fnKvxvO4stywGjRWJyW5Ga5ZuL0XxJ34O2Cd6To+KXcZ2eu8ebeTwacLvu71x9/
Ff+GO4w8FNErI1QiPKHuxfz47wch7PZk/J25thqj0QXPG4pbcPbYVMSHRpf/bP/3
OnfLPuzYfuxesOVARurufIk/ITjVawMCbAIUbG7Bw93htuKQhoD/eI0GXuEgaGzg
XIBqmxzcpmZfAbed/25YOP0Nx4IDB/Vw+sfi/ujJZ7Q90t7WBr79q4AaiAGulSbp
HdKOMjc88TWo+ZqM5HqcoMIW7HKd8ZBgC/P78kHqczO/P41Enw4Le/BMjOEeSfCW
A8OPGK4sLfLNJ/4843mZaL1GJUHmvm610p8ahTX3p8kHnP4CCDGvPt1VckeTrNpI
aCtMQL6mDtSBJhL82ZxBM4o8MYZg07qoZPC3NnEB3NHcM8hjWMtt2i/ptBtRiPjx
W5THBC1V/JDYwA9oI1TqcQClwXbcWkQ/DmqGUSHfJR8dqCvDVYa6ZUv6RiCoDDn+
MKBTYAgr1RJzITBjXLEdmHREruJXjbpa4tG/DfhNjDOSPfwcFDOqmy1KCfOBYqMj
4XQpZ6GU7OywLtU5gUYAH+aC4MwqN7LUsvyCOFlVOd544W05++7IMejFSQinFrJv
8YOKnyWs6seae1IqlR6ovQ1FQJe8d0mYE1xx/bwJ6oZ60jhxRgYeUlns5JgB+xzj
Zt9uKHNGHMVlJqbpMBomGsB4lX6Y+rIgPv3qr71k2+SVUeEkVpfgrLN7rqWjHeOV
AxksUv36KGT8GMKKmBzDVBXkBiZh7ImOlpIWu4aZYYs45NpB0PN+vwrdyV7emqNC
Y0nBtWn6Ccx5WUcaqOLSS2ZZ4B+g9ErqKYdyjvGzUmXECPUQltflqDSUbsH0Jw9c
0xoyASq46erWNiMcnwHNnfjm52jBIbAovJoNIC+z0t9kAiCU8w4GOt/qnT0TWJJC
oc0eF0byjV2RtHuRETUACmR6Lsx1VmC5UaxYGwkwQVoOzGf884WOfp3qBiS8dTjk
UrbWRlQaymj1D0+oZo1h+ZmVwXI/KU93JP2nTMzRHT446bqPsYzyhS2Frh+SRu3X
4+U7k0i4uIvyhIP1WzPpaUpb3tIMPaRBHM3qLK6/NyqiS0+YTsfP0Xhw4mEwmM6U
clnqg0pscKlmP2ovF6K/RvY/9uAdZJTS2PqAvE6lmcm/Frcdv9XzZihn+hXacTzF
pcScIvmj6pebzLZBBuklSM3o8MOcXoodwtGtcj/vYmZeGPye5mCbtTofYAVsQLuI
GWOzzQscGPdZwB8NM9pSWk0Ykfb8hC6xMdZMwDs0jts1NepnAD+9deseMIwYVqta
YpV3jC31Az48hpwIA5fId33gleooFnBaBTJdIkX0UD5mZFDOg0eVgTu5MRz1Yuuz
iPWAPgHbr3WiOs1NWCcDoJzJXTEcPDDZaiLoFbFx6WKUsF6nfBCiWto3QzhJxxdm
nOSjE3X8PEU7oyP02fpJIUIek6edARYLQVDRiQqlmc+QCY/vs3uFfwdhqVxjWKkc
Q7BQSEvzZVQOM5A3AM+Bd7iy5Ci+Io1AJLHsxkpeUm/sTd3lQwlHV2/TOZGbNQ+0
nSLgPVLmvOMj3zQLqNCkuvhnKPGsqxvDEEIrxdTvDqVIc9NwCXuV4NNE3xz0uod6
gEBuqi2F+Co0G0rVnvfE0umgBFG/OcGS2N6cc1aW9V0/c+RRnZalQVUduu2fl4Bm
f4uKQ+a0ZZBQ9Zw1vcNFm6qdOqoBc6hRN03LSGeqZBJBatebP4cHnn7Nmi4urADB
IyKZIPyjIXzqma0ptuyHuoN8bb3JAoOvoHhGLw0Xe7BzR6dhuZ+XneRa7jZiOs/U
FRzRu5yap5NHVptDQcmghczyKPYx45+h/0foXgrHngNFQb3rMZj6Z7BM8r0YFl8j
nNCbOsyn2/tCHBApocNnVpwTCc2IJMnSUqiV/wDlbU8kOI+MpZdWnx30jvmB6vPq
rYL0wVE8FhwDYJ/TPsLsWEDmgzyplSKLOgIlc0jVq98mqDRZHJ5OTQp+Q71fulT7
zwAWyYveA0FptMuPNilXzKytgU3X02PeARb2+46YRik+wziaPkWifyjtiGiJSfn4
pYUWuGg9tsJVxP4XP2j1AM1mMmQ+BvSwQg0a18EjVwf4sAgJUI0+sicxE8Tql6P+
H5kUyk1n9Wct+1Pd+AJM3DwWWzKxAd2BAfBBl9QXwI2b/CJfjdRlDDQRD65buYg3
PGAphAq8lPPpEFkbI695lSQv3Ft2q2ahIbMCPlG3i8/8wnBJExlcnyqgZqhdGvWT
IStX1YpzhPwnispPpHh3p7XrThPziWwsGlRxf7U2G0TM1Z0X0z8RkgS7i9/yN8bo
hmzAvYyukfuwmASC9L3Tz45QUvTLH5BZcLDXP+g3igef14zNzURojARgBN/RmwcE
fYPNs8UPXREZVfmeRG8bfzTx9N0K+yWPWDrFkO9wP0dsqh5dblzhdeodSuaVtM1/
RQisp2QDfh73mXWuPwLiiy/Qx3XuIqPpWplKr1eXCVOnPHNIVFJ22KWh0gwh4ZEy
MDE4pqYzcB0a085Yxq5kB+ejfI0XM66MgJxzTzOBkzl06XKLWvNwHhSf7xlZnUJf
60hFcCAviq5NatN95jCghdQ/aQlYwYTDOW0Q9wzuekTRxnW6/523pKVlnNhlcKfm
Qey4EOLV5rMNwolpwNaT1C+ENrdJ1B5WEjzrKjcH3kboLVC2LDfNOXNcR5E678DE
XW6EMsifuuDZfQzTiBTDedV73bjsW7pmQ4iDiC19M0NIlenZ4kJ8tWHVcuFQNos6
Hp9BP5V0ijMUjA1ldwpLbhSrE0w+opSvEQpMsNVfj0SU644eTMVdXsmHPPw6y7NG
wLYxN6qgE7rnxrPjh33leQRWhNSHDc53IYN3nFEfQrzzXa+lYJ0eg35gd849WAmh
OKaMJQ+KLWL6tVQuPHfSPOVr1xx9cOBWFSANJZx5uL2NZqsk7NPNM2TGvDFflUWs
BX5bxHgd1pW34XwuI94+Vrk/Jxx02N8QFpEiqsKI3UTSvwLb402sN+epA76Yk2RJ
lauvp+5NojztnbgSJVkW8Q2WtZBXskFkoSfnTM/wOsUYx76/vXU/xlWAM3Vtnyo6
d6wdvorhqZvGG1SRN407eD3P10ugXbR6N9BV1p26Rab/vpHdBuypxyyP2CHOcriM
FwpttVuIIJ7hbhyGzld+sH0n9wq1u52GyW0hA08lKXh23raUIx2LYoQDnjTZwRDi
bT02+0PzT7Y/hT1ibf7lW0Usyn3iKIi1b7vz1WXXYi6S8IxNuoP+DUha8iPJob7N
ihUwXwzMoXuGUWHhFg9IVP7vh1vZzeNQaXEgh/IDvCH9e5wmPOHcaG6GQCZRwfiU
TlLTkyGgBWoo9rSzi+TctIuHqjAaTNZ5jAKnWcQbfWeGIBPCA6b88PCG5SlU7Jzz
rcHCV9188RubgCtvPd7hdGt+sMrzGw0NoM7oBK/K3flBreXpZqIttg8d/yFT6mbM
NIiuggPGeEaE1SYNKXgEfS3R5aBo/D7qzrtKIBmYHP0s8HdhnXvHhEaTjg4Fv69w
rLmeU6GFNRDEQ8UARzcaAQ3DIO8nKeTdntckWYFTKRHbT2envl8880lY6sAacXxL
EuirSfK7qlL0eJq0Xc4DbE9rx5QtsFu34Ggr61aFu5Ntx+8E2GBgVqDqyuPBBWIj
AJD9vD0x/qJIXPynjIgbp8+lPS9C9K61shTXK8WHYFlJOnOMR/aEQ8g+Iv3gzCTD
UJLe67721m4yuiU9hoNyqHaY91o9MQbp5R60uoUNKwx8YHM7PlV3b1zyheShM9/X
8jNOe9awzTFTAkxoJKS4/WkfsUqOJ+fo4op9N1UcroABLimWZZL83tf2y0Cshr3I
cFx3Fg4fsKOLzi0crPNoBQR71TyD6wSFD3lCDuJ6iQhYd5PuSOWJcMCzTIf6lGg7
CynTJ9z/W5DkLD7h3aqWgaaRjRQD4WyKiBX1yVM9VK/f28mYY73Y15mwxHTcRc4Y
uzPVOjhUvsvb3cPtet0Ux7DHSnBykNEZtAiCkPbatPbzq1rxhySUWKhbqD6CcaPu
fJvp3Fn3bRIyavIiuq6R7Z9IEDT3gRVOiFbpiLXJne245PMjnDW4DYg8UVY/N+NH
yWXor6tGN7Z1XKKBDaGgJzt5/ZJotMzkaNO7+OfOLK9m9MrolE6+3tfyQH9fZnoI
DCiPiU6jbPJzoGh6DV0egi866DUH7t8vYFCMX0UZ+Jt5qwgobqIWZGKL5benNOYh
vXn+wmbMmcOPQNOPA2xhe3z4XnzoI+dseW4Ny+wbhugbzYQH6N7gdzeESZ866w72
4PVP0ugMCKotqbnjyDEVoj3ts63W+Z1TCmwNHzsXPZ1z6DOmSlpbWRICVVJ6s021
aaD25cdgGOHZtI6X5NJCwjMeh2JymOenKYJ5p6HGQsNLJQBHrRV/ko+CG3+6NCHO
33Mn5Us9zwXtwqn7MtyLegILQphS9lcyXBf2Td7KopOgj1Ry4f+iinuOiYWCMTtQ
Pm2bmrVtwMyPxHhqN1SoUVh6pmBizcD1tW3JVW7RkU/Ims5zAm9rq25O/yln+mmf
Hu8Qwx345WwfJJjbieu7Ow9fcD+De1ZICdsU3zF0JvUyxQ+8OEcCJD4lLTFywmFW
HLD1ZPyCKAVtqb9gbIV1gKplkc5qRYF9d2GC4MI1uku2n6bjEupI/M9bXLgAseX4
5exCMBYJcwnFPrB9tAv2AbVaeVcTbz28GhlKQwLq1U3Hu0oCCZqvSA+GGjtzRrm7
H4vutAalvad0dfAiqZ1aEiovbIFBpe2GbCQKQifBPAm/BG5dEywDyVTlwUadoPeC
qCofoeQxFJSTr1APXZ8sDU59Y7aA08df8gvyFWEKI8hokWNkwh/HocoTPdFbi4t3
jfZ869OQJDhiBFL3k+9ZQtxWb2BhG8i3rmVXzUfNlvj9JafogvfGGuc08wnNvJPw
CeLgQhRI8kP+XICCWnTrIefsnj2QS02GYi7SXBybfJLYwlC4xTXwRM7WT8fCKBaa
eiczPCC0wWhitKBoMdYz16v9iSayo8X2wuv4vbcatelwZ9zVQONLrVKGb7qiKw2g
QMkWzSdbdIW1SiIqSNLO5EgK3xRe6v/yWy+jTKsb6TB1oYVpTxph4bMJpRLhzsD4
3hGnl95v84KMce5iqz+jyFFu/Yx1Z5KWTuCmcSPABvgyRRWAhCsJQYq9xcqsMoHI
zf2GjAMB2FFUMJFEySECIC2hs/hHdxKLMXfzMRBURdT2f1zjzfuwx3IRZz0kYhCr
tBqP0M9kl/cx9j28QgHwWgY0JdVZAeNmTCPMxtPXJukf6xA9WLYKEmetiIxAsNkR
DaRo+WQ+iRiMdSf4V2Aj4aPtdgEtJqvpChyX9Jqz5vcUvbZdtISrqy98O8QfQtIg
psfLa6IWcHHVx709Nn7mbSCRSNOtH994zB0ZsHyhz4II7KNIxK9FMcHAktadQjkV
iWMysERrGdRZ5OO3qpACNyXUKYG2WzScazX1tCbKIBAv9UUmiZP2fZ8VaZZX66l7
Kv4Ce/33ZeJ3xLeMZMblMfj/w1iBr1yfsZM9xOS9M0rcS7LKOGwwgq+GLrWVpnMo
hDfRpT+nOQvhMEoGK2/Nf6G2p+PSJ9jtN05zcUi0Rdv0FsuHlNUUI0Rlpld6MXuy
W1z4nPx4aOXZpTOnrfEARSCWSbBYZ9/XHnsrSCDjis94mj7QJ3hSy1dhObADFfZF
9iEuT8BRHxD1xMNKjGeHwPFItnI3D84vs++JD3neMJ/94/dyTgyTR63pa5Q4LY9J
2HIxNJCjpDzKs17651/WeW/DpMXZf43CZBiJEhRizKIcu65j9jNVaW4XWwIsuTsm
V8agET12qIhVX3QWrhqCffPMqEM1UjkmlMcmi3hgGoEqSXBn7xl0cqWpWg0iNxoW
WDkMpA3hdWcgiyo9K9+R7jZU3DoHUk15kAa0PZPRmEZcHtG8GXkY3FyGgTyXBnrI
hqb+GRcc8TElusE4ZF1O+vStdMsRUWTa6iSjYZBKnvmt27t9ypHgq/UjTGRNqaRM
uQEravpGXz1CtppFpD4sEKaOmpzwy4aPNibUXtAdYYMrDGGGOZAL5IlzkU684VB8
cD2RtuwymKCZPDW4kGTS60sMdqCzqX1dixHscvvlQv8HBcUsW8Zhmgr5oiEFQQoe
UCSrPu25vF4d300HphPLmpkARVopWCrbPdGohm+9WxrwfyjvxtKfMpwPv34QQQQA
09P5VxJSnTMcnUy8RO9v2B7SvtOl6SXDbLFc6cfXarlPPa4JwRuYlDb654XrNV1P
JuM+NfbTGz7bSrI2KwjNMRp634rD+vemmxhCvlVzyB5Tdsa000qLpv2UOBK5gAf0
NwWhg8hOKWMh0WDpAHFwb8xCs1302ogP0NzP/vtTenchyoFUqlvC+SiB89zB3lXU
rJ+Ru2kVSsYTiJr4tGJpYEX26Kwb6PSOJvLZcm1vb0HH+EylAs2wxSUI9f19+HlK
xUjFHVrIZqwkUQQKERhrfl9JQtKYlRQ406AoJlPyA2YHN/WBEBfoiJta4qiQXQmV
px4Pz5QnmXwW+2tEk6EuFL9GUaGuLTo/3zxc0VrW+iAkS2rFphPMYwOOb8ZkvtSI
1ikGWLt30t2NtM8bfBOhEEUfKiv2wNLxinhf0EZymT0CCVyX7/fetaBZ46g/VmJG
5S/6N8y2W+MjM+okXEOfndYIVsi9CXY40FktUBlh1xouPq9dbbZk2pVyc1CqUTg3
XDScd0EfSu3AOTm02vLNmroq0pYA7Af5cjmYhJM3JZxAWr/XgcD6QKXHdPRtDv8E
Dn1VVUoQzP6HPwot5Hn7AvcUAFwz2eudZYMmJ5zzM8Xe7RM1WuircgMzInVgsXOF
Ob08mfk++8sn0WRAFiZ4IYIckXyvoPxABgUISZE11EQb23zanr19Kv8di/Z7fA0z
o2M7m3DEEQE0/Jb4tnLboHN4YaBBWY7VSScagBqWHATGMvNl1x1K0a8gywUdhs4Z
hPJyNd5+aj3JnuJpOipRSo299WkQzuFj2YUPVojkWUyhd3CuCNDrMVNPa4S8Ldup
FtoPmf9vjlQpK2pC7Os3xeYdAezeUmjEcYxHMboEoJ10S2rW+eva0LMv+oJ46nuO
vquFjllNbbq9+PbPJmqN2NVZEeEKdyOXxGQNscX+vnx6phEBxxB3IWSERTRdmEji
2Uw6dUJ36epCIJ7BkPAyv03B4h6NoJxuS/JxqRE9JvIPQcK2J+dfw1FJ77xL73h0
f8gQv+OyM60NoQQD+PriRKrwCGXHDFpb+eyCF/S2T97AyGAyk1ds0g2rmDdbcsFd
ATTebxuSG8V0liN3Q76X8mXuahKec8Hl8o/hQnFXU3weX6WHLkpBEzh4zwk54CMX
0UzN2JLbLHqzWxgwDK1Uo7Bz9aWrXngFMKLc42WgMOvccAxlD8nhsKh6K95qhmNm
EiWpstAQHZPNKUZtuMsZlMMn4mDvXTTp4O5+/fpmUQ2sZ2+gUy3Vf/46EJ8oXeMm
RT1bTnQy5U9fW+AgfJBVsio7xlWcp97cxMK3IXt32ChFsMsmWDX4bn5OQgUUHIrV
IDTRY1riiQE3yzyKQecn6yrlzBF1pJ+fYiXm5mrfbsS+eTcGJC9eNGllG8aqyT+p
t+uMUalMGGT5gW4aqBYv0Khnqy6pEQCRF/dCzv9JsEDKc9hezBr415Efln7Gl5mM
l2WxhtTJr3JIw9ZOkIVPSYfQxXj/8BR6IDJDluGlJL8zNWHZAlzR9kI5nPiwU2y5
vI1tG0YiT5y2kX4YlI3SBmTp7GFY7lZXDNyG6poB9TYVONjULoLLzmMLcfXKNQym
yOc9jxcDg97hP8fsoddpfAUiyu3nSuFxjKOaFLMJRhfA0TV4t4aklAdhF3oJx9cu
dCeemeVWtCwU8lkt+Py4YNuWZr4DEuCbanXXO0RrIqiTEk7EyKgzMkptuy+hcvex
go9rpsC25urjAdHwJo1OQLCKKmhNDtT4dxoI6TwqfJIjiGl8MI4eqTqSHoxY2nMG
Rn7AgaTmPlPOGPTfnzMsw+Pv7SN/mkWqizuOdvuzMmr9kBU9yHQXefORfyLGMBNy
/wBtm5MUDmc6hQLlamyRuXgmIxcYhGmZ5mva4k9yIQBOavBVSXkbEUjgqbEhjY44
UMDNkd9KPfjcaX62tAyPIIQiG5eF/xhDztmZNUU3TSIX55ux9/DO2fQfAq+nOWEK
q+lF0bxIpv2G/u6IkwA7Kk7OWh0S/0p7zHlDrhB38CPELo/Xh+8SgB5lFo4kSWAr
q/Hd7oj29yK9IvTKyfPfq3yRIu07Cph+VzcK3fFJcyPR3AJJUaOujgVuecrytXwH
ekTmMXOjhTZaGrlGFhOz+I3Y54UXGjfGXfaftz8cfqR3HAcFnJ+CAwrTVL7yhhUr
5bIdAIIWlSRxTG3lhrCpuJmTAS664Ie8pOe+X2pRGAXwurlLu7HiiIhoR1s/H40J
8CwXjSpMz5Ab+Ud3kzng76q0nIurJ5CkPQFfgLMYdejV/jh7xa8qS+Er8sOudOMp
m4EdtNTVOoTxoX0pZQco5nHg4VIB2RCEwL6icsPuIfeFKA0gFyQfdW1YNy6pL+w+
nG4TDCiofEgby34KLrXx97N8D7YmZmoI38K0GZqslT16jEvTlzeBUpGSqpbYjF+C
80DFYW+rDRByIwqV6Z5eo1ZFeXpxs6U8BgUu2tBis3Gr50Vq7MyiekR2yh/EyftP
FVhYYxJY0foFt1QGfcMEZGjoHhwlhNsR/OEdppc/b+YhntWpLke+1btlZ3gA94oI
wADAtUMDvb8J4Iu+d0WSYkkWnpuxEj92r8cqd1fjq8evXuzYASOIRRL9E+KqODgL
gyigOe21KAY5jCgJCIZm6yIG+HtxtifOBj7MailXTDcTzvNoI7W5/SQ/mJxSg5dx
NVwCUQqulwYlVpMxhwiOqWTvaIN18xHHGqYx4hp4jW8e7IxyLirRdJqJ3doR+3hl
hsU5Xmr9sf6yZKFqWzzYaqeLGReEL8bCX7omDRVC5jNJZ7sXyS/VAo6tuW9WPyNg
2rWHLeaZ88TL8lu8E0HjuW/rBdI26p1Y8PgNzoVVvY3D8tO/X4AB7PY83JTXLCe0
JLCm/L+XKO/KZkkr/dfIJ4Mz4zmaWhddStPnGuINC1pO6c6z/i9h2j41s82dehQq
kBSB318aVFNWR5pgdsNHLVvyRa4ZCz9iXnh7UDW1OW8Lm0GGz6GJe0jM8wf7MtrB
JcBA/n0ZKwnzAWXJYFzWLS4bu3frOGZNN5INBI6psG+k2r3vaHgFt2dwFhpmFwfe
8SElEyM1AChjQ5rs7OEcCiZ+WUWNAynLBd+fbk1cN+W5Bbo0F1apQRDwgoKyBskp
w9f6rFWMNC3nRakke2QFKrZBGYUhvrW64idxW1MP6IVNh5Kvi3AYB/Q7eq2cpBhj
piKIwlzMRaY2mHm1molr9KGbQVk7x7MMK4zzdNIU5Os/40zCEUQYLfQZo9irxn75
95tZKm7Sm/mL+sqGLJ6UHwPl0AzIOSCxnAhmpGqHDmvTRBWVA0HOBSrBqSDsCEu2
GTnqIQXgv5FpWCRmVqAi++/8XoUa2CH5OZqrLMJ1vvbMV3ygDrYW1Ajo+BKqGunL
MhjjoCT2y68tXRtrcNP0z1/XctdLYlOcacUQMJiKbvKlQf86bEhPLnDzXoQlaTB1
8LsccsH0F7HBmii4Hc0hNdIFoFJO6GqnseGrgKSSCrjdpjK+HgHTUP+z/VJgTmdr
aZ+iRdVXyOGa3tFIkNZ5tIJVOAZziUOfG0gM7JtK4/hRbxKUXrA0QqBFTB5nS+a/
3t5Pmg87D5mzRnmOKCFMyuoh7dmelEQuzwYhKncrmV3BMkO6rjPJmaidOR2+Rg9T
L7OGGyR1v07sP3EPDqmYYdrxts1TNVg8PfhgzbrODC0fGwgD1k+5D2OEJ7eYllCb
WlAK4anvb+Tw3IY/MviA4RsRtjQ+Uu6MbhfIbPNl/DmZdSnkjeXZ7Cp8P/9jc7iP
0VHwcliV8uqtG7uw4RBoxXSUgNm7eq7wbWCINwTunnOH0XdybjXJQm+tP/sVwHdD
mXcQ/6P0yFccJqeFHG6pkYNgxvdFDtC+GRhZesVSwFX5AWuMitJ61rEx413RVdZr
1RwDFYRPYwrGItNlWSatZjXIW0rTxaL3uDiJB7eaY/lItBU8iT6uLiPW3FNw7rv5
1YeDXivM8QYRwZO7nmLx54wr9P0N0x5UPgzulWV49c8WEQIEJM+89CTMmrKjm6SN
NvVByJSoddqrjyLKz+d7KjDr+/H9w236wTzPG3KWNVUqBy4qI0nYlGFRZXUbEbFr
P3qPRUG+otT+sYWvHYLXkPU91yWDXmXXEaiPCQN0+JL3HQoa+zuWQD0Kv8p6XptG
fNGu53eKPAew1/QOuXxtIs0CU/Yg49Wt4kK4IKzM2Qi4SBfsPwETct7PDwqXtcZb
JDi11d3Gy6eE/0vKc/fXC2DV7Y113aoGSccaJ89xu0ZGKTTi0rcTIslH2xTtmKst
tQc3u7eqMf5SYeQO5ScdxdcswWhXNJFSPoki7wUIAqmEQVR3uFb4ozSJ5JiEgCcR
TuSMPmQzdELCJrqQNjGSrDcUJnPFVuXcosUJVub2RxnrB6h6B6PeHN5UksQDHJqP
s6B7ontkFzYVKVb7IUCmUksAOtt2bkqfnepWqOY/evMsLqWHEOp2qEwWBUE9RPuw
b9cchTYrYVOVPuAPopdSIxKluOhnohgvWYnPfff/ZjZDwg0KejGnUaqKWV4Zv4jp
WtV/AQwqMSc+ZgBoGJP7ONopVwYfoqEcG2gW9v+1j99BDoPIKTGM75BhgjOPRQFH
YTzwiOHxujoTVfYZaUZZBBSW2DlYDaskNdt2oFY62DojbuqGot8tutrKxHLe5Lib
CltZdbMpcQXHibNcHzlQEhu9c66HDC400sUwLQ/H8E9iuFGRuER/E0Mq+GUoBlXi
j27FEHORC09ZJPD9SUKVnrltlIEaXo/0biAiZ+TZkB5RSOa+QI01FamKxybs8gxg
v4rS0Sr5y1wNss6Mn3jxxaFZ2Wv3opU7OQgvQ1R9DHJsmzwSVvFIHcNRJR9adX5S
eqUhosAQz/GXIxMo6qs/BBXsOt43ccSvX55/To2aPm/yEgIiTlQMvEBNng0Vf1mZ
4sFfLNp901fVjDA7QqzTvhtNIOImxrpT2Axg6ls7Ngrgs/7AkixdnNz3D6RYlDLX
67/qb7gjsiOLfVIhoofCypgP+tmHdZndNUtxzYN4gW6213uePq+vA8Ds7tp77NtY
OiMMTHZfzVvCciwrvokUoqz5thco+JQjTIllG8P9G5vnP7xtT5LLLxE6P6BQxiA9
6Qbp4J9tnIYqOveP6izbIckn6VCeKwnwgbCsWAedTyZuaFXMCCZKcXcCRcr2rLnQ
Z0P8EfdVjml858L49GoT1BFizd/DG28MB8VE/L76y3gU6s40v0o0TOiXMXENDllp
gUOq48kF71zhC8S9W8+k34OjFyfeZiuOn40D6PrIdXXNoIH13VEDZfTE+mJif03o
+E0zmmOcD9MMDv0U35r4K1wKc/XH/fw8e8AR2RY0wr5Bvj9mND4K1bWJNxBQkOf2
feSmSp/N/TiGyPuUnKwr+s1qPAR1dBT+EU7Wet+SmIsdvcY7pjBhukSOqpmFBFiA
gdR0WDpdgrNJUDRfvoEVGU0Q/lU+Q6pl4GHjcItN9UVqWQRBmbs/L9d5Iv9wCoZ+
CLNwnDbRaEoSkZdTt4Q5ECwpKvZ9rnFi3CVACYU9ZuCq74QC6CtuPg2Pa+5Wqmi5
o2ajrnCTkSH2xpPP/3EQupoF3Wla6GN16QqF12gIv//V7Y2c7620LKjqmGSKBU+j
dWdcgL46hSC1JHgEJJh4JYKmUXDgXpTpiGUjOtIGOfQ/XUqPY8F979TVAmBzpUBn
6nrsRrLMYQn2jMvfMKblDILzePK19bpnRvWWNMbNaaEXY4Qd07ZVhxY5PjTmh+zB
lE2regRdmUjK45oRVdL4OVuXm4gsmCe3WO5+tJVnRi3MhIiL+Qem3VNcncU6ICFA
ftaN0B824tSZUi009byZo7no0pYnKKa9kvXZ1g/5UWbh4AJ8REhdG1RRaH/yBLbM
bBiu/3Qr4GGNirH33QYe5L+IbnZXZVXnFgodGbHotlFVCJKro0TlIW7/XB5PmOtA
UpMz3l9Ya3Wazllge3SxqBjbyPjo+OTEbSS8nruYMGKseKDT1M8g4ejUQEqQ7KB+
wS4CWdkBbtZENp98RXTSX0Cz0IMwbsBaBUBq+r8gCTN0O+z+fF9UGdfGZ/+rtK3f
XkUWMJHR5BNDdnagQRKVjemMqcUSctsv1WYK7cFVfm6ZzXxu8rFRYVHRtlw5MfqJ
/B8QQOnv5X/ja3dTTO2BLRkJJi9iC6limMhN5EKr2uHltVFpKXbMQhctrwW0fdOj
/iBq7/c8tnkJD70UuII47U+QfBLs5HEZru9nsv1yvKv3wtJxld6iwfcbKiMl+1fT
WWCC5zIXsqM8th+mQCfOJW+YCCf/C5UUIfaEwjoZVSsyq5dBV9lNqUCxRgTg1jwu
cdFPjsSSaYY9SmxeiCF1sGe+gNifSQA3fF9jZRYSNwu9g5EFtgxx/QTbaV/45AJ8
iOFSA13/ihUrl6KHxeSJ7OE0oWR4VTyVxAItkf2NvOxPR9DLFwEAq5Gw1rE3LUp/
COb8LlIPzp1T2IHT4dlqIzFtMV4bAEMbf1vsPWXS59tCCVK1Pas5gqXtvC5oYaNZ
VJF7z8nCS78MUJ3kFflJ38LdcGhEK6hgHXb04pTVRd6TcSZcavIJb3JZDbt1nhWs
YxO4gCDJnMyJ3qkVtMgvUR/ebq1n6BdS0Yt942N1syq2b49AdU9Vh74VjiyUZwVS
cksErau54BGarjhew0jD+qRNAcE7Arh3CKf0jcYcH5/+pp1j5YXLpxjEHCrLa1dr
oRxRvyDvmCXp9XPJEfwvp6eJIQzWTbGIn28skGfNUwhH56rKIYhV1Ob1m69MQ3Qz
7SdEXw2a73YCXzmM53ipDZkIMq/s5NdrO68Tu1JYQp2Khe/+7C8eKscbds8cPqdx
vee4CWwQTCPkE2ry42HFIPUn+n8m0XWZEk+2J9cyzkggRdhsAq4rpqIxBQRNwp8s
gLeAL0Nm3DSSQgef0xcTcHVZNONN30C3MnnGUUFV2bdeZ7xgtDUXeC5A1BLMCQmy
bkArf2ApaNle/4pOHHXFgNnoit3OIGVB4dhq87oPyfLcRgBDMWWX98ar3bQ8wEIp
yvVeUVqXZ8nROxvCoUn6wSvklhbu1p1EACwvq3N/rXiTeI3u8bgPMdMdbrN1unci
7MHLcTPD5P8LiPzmJWppTQctaUb8XbK/JgQWHQNPUgP2dmzDB6Td/R3KIsLkpVEm
zYUJDu51MiseCbjuf1EELprt8TojWE0WL0dZToLAQjid+wmGyIaC1a/0Qe9CDeiJ
cioLHBnbOwDQXr9AkHHU+hjOADM3aysZum/juGeLGR1p3rG8HifL3tWArL0VPG+x
nqeOKx9hwBqAQ0opFA0IhC0DrONMSVWiW/er7jyPJRo45sqApVlRdts6xSSZOHKQ
4l7AFjuC/F3ORmaHvQ7rF5CW4xNtCap0GqgYTxAY5830CRdY4NRKRyQ4sdhI3GPC
xxQFuxq7gZh1IsX7I6eoPQDPO8IWYnfTlHnfzFcR/NJX95C37SVE5BEgdhvMCRiQ
vBu/v7yGZp2kM8z3mna5mwQvJix0E8P2YTiSO1etg2Bt431hu45HiRaYE/4gyKw1
vEtDEHlpn2XVjajfVNgkTOL/JcRaig8bW5zNKDXAAI6UT/mpYtmb3Ld/q5b43cEW
83RFbdc2uK30p4F3NzdwzTXqJrgcq76CAAbd1Ns8Y7pNx8kjDVg9U2JDYc5Mvt+N
8hxoAXdnefXHOpKTVb5CyE41w9+Y1h09dvV7jz+cnH7auHO/JduAM00Vpu0hGGjr
xHxa8FkHdqgTPBPlDYO+yEs+tPOIds7Inq6DBaonFmMq88lh+bP/+3jeUYA8Fjc5
fPNQs57OjZaveJSTW2NsUM/d7hHITF422QlvyKJEVgQxXjqdzImbVHd/+fP6+z3V
xphxiGH7ayatf2QB02RnL4Tn/ol7dNcySj//GPHyh/yqQqdVObKKhzArN/bJZuqr
JO5ti5oY7f9ZRInQ9qMaPUs8/os0YU/M6TOVImFI0EAJLjCJ0yPuFUqgE56J71zw
qkLXvqjXv5nq0y8MeancC6UgaT8j/5MMBQSCSsFKQN/Fszl/Bq0Gj2nqt297oQum
Mv2J7o21OfVogu+gV33bASXvsKjLlp2+cOIqEk1W+l2RWULBD1kXnMrNDt3ZW08x
jzGCnftbr13RSgqXy+gJf7xqg1wOHKcWRRYCbw7QlwhyO63ZHdWPyaJ26AZ9vT6y
5cPzMzt4gg3MfT/WJfBtFqvSixK80DhNRwUU8TonG1dJiRQFz8L40CEUhwW8eQap
D1/GRO62VBcQmqemUheKW7XAAo6HtWJHx684TaX7C/UTha5WP5E974J0f/5cNM26
9h60eUoTRWizels78ymCpFGEA1MfS5W3kCSPLdxeLeRvKZ1oiQeREovwPmeJTNcD
r65iWSkIHqt6C4/xRxLwtb+JUl+BaYATiKtTdJ9CVBil+G7DfQZ5zGBW12/XLjZD
wjnLRamauTM3ntu5vn4SfSqm02+l1T5yxumg791svxGqa0XuWmG2F+4tr94ZoFGb
ShGV/o3sdabrs8816hBuDVWYUuNNUZ/AWzKQGmL9mCkyyxzlD6VaYMrU24cGcuqf
MqyYtrn/Zocpm4gMcYUuVqGDDXBU0jQyIo7cX9OXCw+ycFFwbob4FDym7xeV0uX8
QHOVYHuaRxT8DSw8fwtly7ZgPl8/iSV75DbZhAeuuZ+0373bw6x7dyYHb7Lf3nPv
FRouuH+UdPV1UI1MjRncgEg0VQf2a3TWx3+NH4tp6zvpfohCNpOSltjZFDlSDYjX
5pBBM3NX+8yYiLaI+9VWFdNjULaZlFxxCijn+Oy8FYO29DbIJVth5x+Hm9V2UAD/
enuoPoVyJ5kPnHOxI3Yk4CkM38JxXWpWAyDmVW14yfTPGK7cdEatbCycKLHq/4AG
kEmPcAGzOwapM3zTGaAVZybuMOD3JwebipRorsojrKcN61C6Giqq64DaXdc0bP0E
Wmh4MC54eiQ6bSk0Pe5VJYmqUJ4OgU2Ha8RtB/EZsax8vt4Wx6d0LWfYpEqWRYxx
LXmFmu1s8l4gAObsoolQTjer/qvix0R/9isZRewOgenus/hEb+nyiZE7HxNcLzjp
YWvR21KHbv76GDvOlzNj0ZruEaXFux43THKjByWHJqVbQBlr/eS69GyOg9WHTktx
Kn3XA9sYYcSXPtH0V+fJoPcO8mqWolkeeSfrTbXzyNoac64G0DwzvkVrlzpzWk/p
IEk7arG6I45iCWi5Dc9L249DZdvrBbdktg1snfiC9jFKuRLEjndJ35KzZglA8qv8
QK/zGZj5Y6VtScTIMiZXv5rYEvMONi79xv/51b4VC55TKwIgA9klm5UFTL1IV9te
RwL0tlI5kFulbKiclgSaVlW5hhwRRlWspyUuqtJWs9VhYM6FExMTaqRy1QVD32tc
V/8AVVXT3z4AfLXUK6hw4yoHG85lnPZOAD4FRwIkwK99P6H7KajUkl0YeV52MyYP
CzPQ7H+CJJL24WM2gHuz7bNv3anXSHSySDPxVmNiObZ2QxnYtHjMHqSgynzxEtCR
n/4Whc5oQxvldGEiy+ckoiuR6BjcbVlj8HzbN9AvnKHF3ITT36f3589xDWLKKxz7
WH7lXB460vnY56nwhmKc66R+l97Qj1jdvV89K2nPOjccLvnnu79uPfB7vV85npve
kO65t0NPLCuGHqx9XmiIDhjSkmye7S7QIwzcvhEtEpPVOBc/bBdEnaIQwxPgVFD6
t+lztUzuUAM5UHg7WWRdvTyv/OaelW/Un5nE6lo1s5bnb7IfuNhiIYbM3KQYENil
gIlbxjcMtm5rizj2uwjqk398gEitPXMQx2eTale3Xvqha5fE5NFT4o9/LsPunCqa
O6iFT/Po+JRHNv7o1h7TK+8VhjhaS3PqBRn1yiPZEitL7HD4iHG5XmDwChpCawGu
d9X1nrYg0sdLCkhbMOybTZOnZNFGE6hzRD908pZzvj4g61G8bDdb0m1OJ/elvyiB
CsC7AL9AKZ2GOVozeYQeOWnj8uigRSNP5lbLdy+fhKXBK8aRa4cosngoi5JoYV8T
HMuddIAP+pC+p76O3K9kPPLEHPWNOK/p1/p/XVowqb1X+7Nb8OlOH4ShKvWQAAdE
xMK5zokuKm6eaUQMEa4Yb8GsREbdQ23sl0tGZ9c8QUgh0PucabRJMumjeftLt3up
K0Udqohq2MnhhviwMdWy8vIVmaM+nKZENQzYNMdvYDl8j7xzrFfvGvINvrnv/PP5
QVeYsCTAw4/cKjKKEPs2p6GxfM+UAdQTU0zShTjgh6O6NCa6qjwhNStMu4dmxLAT
0Gm8jsrkwsNnuf46zQ/QuvkSXuqy0aTIuIeB0mo15RZITgHScs7vJEBcObXBNsK9
Mapg8F0P7oyJQixEpLE4m5VF5VAvDMn5EJK0yM1AXNmQoVopUUpIZlJLAzfhiJrk
emv3lr/PFh9+2QtOa7SwHN4O3Dyp9aAYkPR2Q1j9T/rBtZ5zpA90lXBAupJ4HA2i
25a8F/2Iqeg4gKeiaKwHoLs0RTy7Zlut83PWVxq5jj5Nx1ko8mts2ZTjDk0Nyi2C
YD+Gq+vusfxo3F4JuRfwVW/hyZZQFsUBfj8PJq3yi0lBkHaiC5UD38oXcgxr8f+y
QN8aqAXGeRJV1oaxhK4mf0Q/QWLxzi8gQ+6PNagDg/tiNdpMiUiBjPZraYLPEEKt
OgPHn9Y9fiDg+X8dkgU9oTAPa/vWYkpa2FngOOSKNTWuNS699VESiBfwgJfX5YSs
kBmNXDuRZ6HQslG3wV9o2o0j5kWg50exf97a1oD1kcWeGIdSJqJ8BUjH2ay2Qgrb
mfks2M4349ZRJqki8wEn7U8BOb57YTIeB3kxIKAWIKBkcSdfmnz419ao2AKbcAdA
abzVwvrajd0nwahSQCJu9OP3IzIOc3mhhZTgo4j4zmusw+abEf+jerda3paFf8nq
VFkpoNboQGRM2063hAo0FLj8m4yB2h1dk39UmakSBKB33srV/58hXwb+qC+Vjo9+
fhV+RQ/whOsYgRNOtgrOatiRHXAimRhOeWwUKhLyMymoXHFAe9fVBWFk3GJV4371
i3f1U0tXtz7vUUXf6wKpIZT6NV7Gc6+Jj1zRxY16BcsZy+oJv+PCcpwdsKOG+KKK
OmHXip5PAV+PpeAnNLIHZeQ2d0thYPij2VwgJrgIP9TS8u3utBI0/tA0ongYnpiU
JmBk9pzGZrlBgbJ3gcYXtMN9aTSqS2hzxBIrbzHGouJnEiCD2NljS+rZwNKzHeMb
6FxkZxxd3buUcKT10u+RDFw+ZSbRuhYf4ogqsZltQSOAhEIP89Srlv9MXuotGYQR
J3FdEfvYeNwjj9q177076aPendXPTBpZv0vqDibZFSNTON3RBOetXFfbSDfcb8AJ
1NNMYlF6QeedOlqqO/dvLAfcS716Gu06IfJZz4h2+J4bBwNGIY6na1YksjM/q5mV
ocOPrN1PpGeGwHVPtDmlU3jGj2J6exLktWQVwKnbW4nuvyqHzdqrsp/ZC/wdXkfn
HiZc3fDJm881q6bqYZUDD0qTLilnM48P9GC0Tqqrhr8ACFRHC/Uw7fYwl8iG2vJs
XGonAANWzDnVLtna6oHKa95qnMNorpaIPrOHH3ZYAnre55N4DgO14vhz2xrVqUmB
ezUySuDhOVRif75g/t2CxO1lJXnG1X9sggVADx5n8ZKJDNNqmqLwLnFTDa2ZpPeN
WW18y1VQeiTcPz8IudIZAxcvH/uD2tf+pzLyarcZhW8P2daQSAMXVP8yFbSHebqp
xzh6XJeFQnZAhwx4GNSxpjr8g6D8ly55IUed192NwtFphdfI5PapQJ1hIIxWvkMO
/3GHxE5fPVbhYVUM781Jk6uuThsXQA6Z0nR7tzpTaRznpIPX6UQ7wyaC2nWyfgoL
fTcvync+IPmVeBdvOXUNYnoA3trm9OFS/VKYEy3NXIOhhiq+IDuOc85NyMNHQiIg
J3nBKHAoiAhtR7yyt0fNJ4zsrEsZhFS7CiWsD4YxyHRK8l/ZrK7x5BwLzSkWj6Rx
ecUMohXH0SL3gNc67hQludNHOLxoyFL/6mDbIW9dmygKFAs4v6x7hDYpkHeBnO23
wv2+I5zVJRyOo+FqhPXtsvdcxrUkm0cPoRSouAz3cnEJGczqPdtmHgKe8mwV8Hrb
w9Bj1LbTZkHPsusifCR2kM/UxkyEHZl+3eWFWQut2sUSM1gxX4Gx9NmptsLRyQ/O
7u113qr6EASicwG7+8SYkTY2f9h/30nLXaKzjmo8gy1yBBN3+xzrE9Z+805Ffnox
2GYuYCMmdXG5iDoqI01b+UZM48QEDuKxxYDjZORNlvmEgIpoENEAcWtcscyEPQ2/
y/4CubxqugMajSRJjsR6PuX/PAIFHb1FGrW9hcLjyFB/EQp8XJ7wa0Tv+8ZXSrFA
wFmyEFvor1IB7IFWTEN+ahgMyhRQb+OoVaoKdviT87YwLWDSf4rYDUQZuSe+WHRu
kwWn5L2M++K4zZQ3CNlM3qE+ysa0JwLNoiGbZpP0NJohk9qUxmu5w7oQIo8oAiL4
+BgtycQ/SxrueP0nkWEqIlDOOQRk+v3T4OtLb8zY3/SvTysV6BuXIXNjUPoIRK93
g6mVFRJeMmi9gGXTkgEpyd6o3akkY7boPOU1DHiDTqGGe/YCLw8L9m4bo2foankJ
5f9SpczioX2yIDNxkeuhjYwmSaaU8vFCXV2ftWJgh02157Se5FvnO8NHppIl4PtJ
6wW3QiPhiU7SaVj0by/tzc8yXP3Ia9NhHlBKPDQmPGq1qnVZzhbE4Ny746/Hpg6q
wxie4wwuJ0S9qcvFKTOZ/lRqovrbAWxlE8ErBcT0Hkt6kS+j8//uuCKF8ujM4doI
tA6TAxVk4uzlWYR4fQLRmCPgAgoYy0HDSSxL7V4J8BTGVA0dQcF06vPwzjoupHOr
U7AJmIZmmdpH+CpgbOmddmT7U9yKLW2HF6MLT34v1ZEgXwm0/rke9bzz7rgTPHmS
dn+0tTXCOOXyJLxNkdfeEXEhrRPTpqmLzqLu6ylC8J9eSd+cQXPQEw7/eTtwhxeZ
zeRUv0EjryBM8Zvc2G4OaDWPlwNaSgh4YqrmA//W2i/0d5ibvEyahuUR3UGzkngW
qHVv4CuV2KUjKqOnl5LBzHMcvryn/jUGBHh048nWiPdZ6UUPRASa119/6xitU1kg
Zmafub1towypRHDX731Tzvyd4zYVnSHc4z74amiliNEkLjdpssM1F2tCafw+0lnI
cetVr04afCj/KVlatMYdCFGGdIxrKk+NxHGMcNQJcrle3aMmogjo2YtNBVR6knFg
FO+JfzB9rLpkPK9zcBgkJ4EQn1//walOiyzfLqJ2ucPVXsw4/Y6sGh9FRf8do2lY
MhRp+4rFAVy3pB4/Vr9TP30Rlwc4z+OfNcYPCV6IMOqxYNydW+9pbAqf8PiMfecJ
ARCe089T2wNYhCQwigovv7JRcNKjWxtF8ABBcTU0Yi2cJIpD/TDSD5pWxQo/X08i
RKFteImjoZi6pWRKwDelHFYKjavse6/S9uZ98HRXyxbbuqXvKEuGrUiI9y42pjZ5
3gMEjvFlwhNiO8lKfYBNJtykBTZQ2x9dU9RXBklBz1N0U6toBTm3Awhrtt5JtEQX
hMRJX7K6i0Ei7cb4FYvHxyDhasveKGFqYCE52ua9+l4OmykAqdATONh86/xoywaQ
rGaHgJstIU0CZhVck0wjEN67C86vHOxpjpv9Fn196kFxh/sm8qFq+d2QfC7WmG4s
DDhJyxRZd5qmuI2HWKELszGUm6fvzue/0Mxn3Qt7KiUffRkZjSEYcvOKtIwR5r+m
VCSfi/tu+4CWItB9A/3Kn/HqqH0ld5gSh9y5afEe1yP1kAf26CUJ7wnEoKPcF3H7
YXcou5E4MGUPzWRXubLpKQaugqeTLZmcPh5o9WbcOTV/Agz7W93xFtCG7x+KDzHS
xkHCatigkIU6Dx/1+hwmSwJwYUsA1mueOhWB3JwuQknnFxmT6gjaGN0AcCL7STfN
HfmBnYSu5YWD8fsjKFYVyqLDI3K2cl2BsSv00IhaZfZGmOQ70rtGHo8D5DoHXtXl
LT4CRItS4qL6F4/cZykmAK4c6SnSQ8Lotiuw1genx4nzeivwv1z0R4IyPjpiRO4M
spuA8KQVvNw7ae12w4JCgaUgPdeR3JWgU5INOOmqFwhDpTwVBPLwzSKhPKkRZhg3
TjS6TjeqMZWpyst57Qo5xSYLeN7lm1S8QUqIrsGMMC0Df0bHl75m8mUQYAKW/ikR
oYleX4+vyAMqareDG9wg0yZX29OpNQpWBL6Tgca1zl/wxa5xxEqzYWDf5dOPXVYh
CdISAhRXnuwCt67qZvLeQjjtujXfjz5lJg8aaF2QwNR4+qQpEnm41iHmPIHbpeOS
QPVaQ814urLL4bnnN1p8z4vz8RqYS2hypBfZH/lwWcacsaXeaoGEBOEUt1Z6EZyt
L9b2YmcV6L4HyGM2rCTzVgVSX40VMCwriWiGLWRdRelaSI89btKZuehEVdyqShvJ
YhnHDZJUAjwIB81cUII4RCQOo59m1gFb7Sh9NrWh7jyE0PiNgOiMhhq10KP/sXgW
h9RfHXzj6TE4ADkU3wYgSAUD254ycSls+A+v55Wa3u40LolhyDqkL7wfH6IfHNWf
wMpYaY73gFR5K+cAET5R1SYl3EBsY341QGh6cOui/iBaLNXTvelWsaIprL3nZbDZ
pbuTQGt0EhvF9kOtcW9REufw7cyaBJexpQkVtaXK74NqmjkAe4mWGeulM5iZHgxj
IJ5wlK1rpTnDoxpKw3X6eJi/s4VKeTurfgCpbVXFtX06M+ljqNZB90KP03W2GpP0
Wh8Zie9G/jHb+78zkCgqZEMBazx+QRMnNKJYdAOQQq0SKD/TQVqlaLvkmf/qibPZ
sY8GoYF+FqvKaFVYWIG0veqOjwWcNBzXIaYvK2AX3/JqUquoRnb93bka4moFpRgM
R0xDXhvUCNvLjwi7sbadL3SKWKR2d+arInf4M949aGCfvoIZ2W+YeG09gyPzJBpB
6E812Cq/Lqb7Hkh5J/5ajf2F/dgd4q3N/sBCoOD3X11C7ScfMB6J4q1T2yQ08F3T
k2dlfkEOVjePDVL2xcHDA4MF1OqR7ED/001zxoWFV1s+AauNLbOa8O8vXaeYHvWq
SPf0TDmbrGSJt3j+LIo/BEbftxB8XnHfwBig/Jxlpqm2zybpUmzStRuVu0BZw6xi
aTThAruBKmTGCGE5aR4yli6Ad3+ZphhfFrIiEHtL+Q5KzEFyDFhWFDp2RiMKEpm4
6sj5dqg3vf0O+oF6KZm4rxUKX+iiP0LIAS2Ornbm3IP9yTVOySOiGL1hN+grtEh9
WoZq4e/GUc7fHsXYZnI+1jlLOfz9P8S8qnNeu2BSRG6C4Xz1xbKu2DQLAMaVNmyQ
hWsinrDZwVcMEzBA6YkmQb8eh/PxOzu4M4TtZmO6n8cHJBG6Ie7gRj4QCeto0h76
ImJnxoSFpdWllKnSm96Uquct7/et/jDQerf8FmcASu1BOwglPBQ8P2K9kZSsy3FI
fnNf3welLhDliChaNdKBTBOAtT9hFsur+bSn9QmUv9Mu/cdiZKliIw40/5GMsQbH
Q3dVLtGA+7Ajso5uREyQzsMDgeCWeY6Yar3brxJSLbnFDCMxNWApEuqZMe3QNiD9
t3C1Xlj2CnbHrfqQzclIs/Q2NipNiY2AJayA12X4lX5VRmIXvOnDoH8d6o/m24X/
lBHDswfoQHuTHY2ECo6jLcTCj9u/xeptQkB3sA7eLnP7uHSGz/+W2+43AQgjFzwA
A1uuAi7V++Dt9f5636kcGC1TM4rvHPMH5bXPV0b7KSZ6OLSQIv//ZBrl3qdjpbD7
hjhF8Hsoz00UzcC17Y/59IkLuHvoKUcdRuNtHP4DVC3bUsHIUUizXbW8UIl0D5M6
4O3AVlfUCINzjRDYjidiou75CSaGN7t3VxvuM6r37s3Xj4agcRUbgH2RI0HlBSM+
wfCEspuGh8zwMwlfHAdNZbKCzX0ArtURRFLb+TVzlALVHIkunyWLoTuyfstVSfke
vWGUx1lSYwzUxdannbLsh8yoLC/+m2cirLFI8581KfUChjck5fQpYN6bM08q9DNT
5Jjm6+pZu+DxxVqDHWgi/25fp6Pckpkx9JiL7sxhZGaGrc6X7ZtS3s2x39EE5N8o
5qly0N2hbX9d6pwkdE7zkiR0acOdessulbIgnpj5UuD1ve01AOrFvfFZ/eKUsxLW
eRQ0agOg+j5Yck7yJaNIWgETND6cfFxs164rzeOaLOeguetybRVShB3/K4Xg9W9E
hHeIth+Km2FN4hLTpsa9rUOC0c9GA3FxZ0SbeJeBekD9zO7bkPXY9oJe+LdPkMGA
Q8PtGEwgRvLK570S5DifeVqrQdsps2ioW9fOB7g1GGpiyv+LDjCuniDEC7zPwq3f
gMb4K8U4TQm9YNZlVdyxwQZMsFnbvwDswu3zUqZTi4ebBr+rAnQBU1fnBOcGhnAN
JgYEP/kA6bBOba/OUeSFEOC0i5d9dxYx24t+doNkJ8V0djaZKQv95iYxJ0q7zIOE
P+r55cOVzRcCiqv8u/4XY19L6uDWUcy9RA+GZmFCRwwWXxmaEvJ2TVjzmIsfUP34
PN+tp1Tdss/OEa7QK8U0eLpFUKmok1Lug0j4rqI6or99M0F2yMHZzE7F863fSKcw
mZtrb36ztrky88Nz8BO+8atL/SskPCIRbBRmeAudndlNx+cyVIOX3A2R91F1pxrf
o9gyDGbZ9rQrfEmHw/93qR30B2tHJf3+LcZhQFs1Mz2Cu6uds9gQexCps5DkL3YU
Y+hro12qyI9zG5UQB04VDoXrkNBEEVdqHsccdeBBKsPPf8yVIf5xYDZtYRHJCFy0
tXS1qSNQliR/rRVKyfPpXleH8dxXisXSbqiwDQkpGy4WP40XFNKUmZbbc19AHqia
VLxNtRBsVw64Z8TcvxzBbQfBa7dz4+/T+xIuapg1acLiFmcp+ojS3+4wlEsNJ1UO
YUZgQFvCpYzRWaGx2HBEzsiluwFNM/5zfctblabxe5vKaNY9AvDRPvLBBlee7zsu
rhcfz+Mb7jdUm/xOHu7v7TK9UEwjO55cv9e6aB4KJApyvHLqh/Z/8GaLZt302MTe
mGIqWgM6gs96x4dNxyuzzRO1hkKSpSiuBFkihFcXe1dfNmCa5K5zeCekYIp+k1xG
ocBG1ggRMGSSgh9kJ9rXhLpdoDRamsDubiJoUT93Rw4yXnIQ4l6Gl13J8hdy16L9
sDUFXvTwjRuh9VLOQ5xn94vpT4JzSlCr+PuQg1Xg1ox9KUuzTuEifmM6KsMFuQxZ
ANFuu6DeEI+YoCG518Rk0kqjUILzncAsOV80eLf/FvBwnNIq+KEkCOrfPP7vgD3/
jdE5z2+ct+UtMwHrPFxWs9bvEkwL6LGnxjbIrVya4AVV0Zh/33QHZjEg2kr+fkDa
p54rEZJSv93ZHjMV4z7XhAxSX/R7Mb6Pa/R+PglcfnCrtcjy3EGV+LTczhY2YnRS
QMHhafc1ScJeLCuw0jkwT9487HEenAH7SDssmwSpJJaMFUIG0O5RAcPWvwO1TRy4
78A0oHLgxvcyzisZGTQtbCidYbDoqbP46kFJwhiOPg36u8B958mBFPqHBHHZT2m6
1FT5ZJnbOB6qPliR68tKwlFsmRmXHcxrlkgv6W9AzE1883zTWXsa9nei7gIbyy5U
KY8in8R+FdjKoi8n3xVgNM9LT65crwS4uqbR/7WYXmnnmzyv71q6edfuIC+fDFfc
ZR19vGLGt7uNFJfvWdVyBLXb5lKWdzrNWVvhH9rEO7Eb0NnGecn+hX11AEwk8p2O
jlVmoDsLwKHv7p0QGmyf6MPudDsMyGXroCRmJQlLp+Ci1GVK1/TrWJMPn95WtqS/
yeSMI8PwG9PRXNjfTr3ZbPse77Ga6qF3aSKEXJx6DndaCNrs5kv1fLFXfqq5xolX
8KViXf2syLQrcVU9pFwirAyYycvgM0NJzvKu5mp4cd6DOhkzkLteoKgFJGFpN2Oc
fiC55IfbDj8W7IlIWkXnoOUfCxtOJ/nQcp83Gf921W7v5onNhKsp1t4uxICAd6zB
71QvKK68jioRNXvf27k7rcIK71WbKBhZy6Pr648STY1/GOtWfUfrKk8r4KeipN75
UwGYuRxo8VPuoTum1cI8qkk4qoow4CcFMvl6LB60UV2BuSzPVAdOfP86CsW2owgc
5cCxiYS51DwQABl707fE/KwgShKFDh7JwDRupLxOIPbp65H28xbU2ucLTTnXdWGX
/JIgV7n9h4fA5Z/Ri5tiSh6Ck/aPmxlilVhO8p6HK9Ae3mywr1RDZqsvhvLaL1Ym
K9TVSmsGYYnLRs/0iMcznOV76JyuuPlWp74GxbxnuHS7H6qlhjv4JoMg9xGEMfeK
1mD1AiVPUrI5QwSIJsGTq0DsNGjWFkw9cC8XN8gey1tKV7PQg+X0n2X+1lLAR79S
LdRX+wldf9Qn1VdVjkbpDKnGB43F/z3SKsB80vGQmDKpV7ZtIy7wSYgXXTpak92e
CPhq8ukL0socZMIxIxVtoKpBlWxFiYdXQI7j8SKOQHOGTreyJTz3utNwaM6n2dE1
QpK73B9ShUqg73TcqXB7uIIZd1I9RsTC8G2AcdrILO4mUfrIUhXb3ViCKhBEb9O4
drIQrKWw9VCbmvKOyCcoFUZqBYWz6MJOFotm1mwfbDtrjKn/u4FhBByi3NUQ2lF+
zOnuhX5xHwBYurBy9M2UUFefZzp9hXplhefj4VxlVlu6xGyQxgcO+zLGGYoYNsqw
94BE3fAagcObmpPH7KwzZlIPBqCprGYy8a0vOOh7vThtg7hRfbmcZfc2hg5MR2ut
8VAYqOvufNON54G9XYarVPqu7/IVmvln5hC+hWQjsum9Z38dhSe45wbzmArCRET9
/yjPcghHz5pAo8jkE5j8htuW39Se0tOtnHmDApWdUy5M6pHexb2lAiFxbA75Bafp
/3ZkuwrAKC6umaNk0uduvxI6rPkjCX/dPXltbCFfkNPG9P5EJQ8X+8Q/RmEEWGzM
0qUZft/hht+IzzEvn21k1cB19DAjpWogig6QCHb/IZxeQbXQ2JbpfVt46qWImqnw
nzg9mC+9BQhuhkphYnh//Epr4otWAAbOliShEjB4HPZnwI1hWQavvxjoR6gd1BEz
AGtkNwU6h47Azmz+CLeCYNtuDnarnl5JsKDyTnWjw7TPLWMmk8gok6B2Acx8zNcI
hcq/nfBc8WnjuZo+2VcoR7kolBqnz9sxjirQWuZKBOCeeF+FGA0Bbja3MOH4TaPm
eFuhOC2CcDe42dL9G1sw2FeGe8yL6gTTYgdhl3aGd9Z9gKxE+ilA6YsF8N6idHnG
0e1PuwLpdz4/Cs3fsCI6Y4IUP2yu6mUoUtCrwf4txJRWM5xX9TiLaT29J7/uROLZ
SA1v9F1HQyISjtyDkJoSQqiweN9TM4VG4YSyplqFI0Vd7RYiojCKsXdNOcxk5Lw1
4hCxcd5oYvaAu/PMVCpLc1UjpnWZQQXrvrwuGUa9+PwYCBr+FnpwAcoLGqiAdXoQ
rTkVsOzrAgRVchhLlYb41nAv21dS+i5tyxK9O+khC8Onz/ofM1SsFLsGKHZKqTN2
K0uCdccb49kaZMDuYNNHda/S2TK4PZy5cvi5VHQwCMASJyFi+ZFDg1UA94T9wSkA
ksiF5EE+NCpSsOdHLrTDStmvt8VuzQRu7iFUphbRCCMO2z7d/jWr2OV+10kBVVEp
ms4p6PkuOx57iiAv7hmcWjuRYf7ycq1Zj66feVXSB90evnHwYXw2w55hpPo9SP8D
c/xUg/cX8+vz2Qc8qSIp+EsIBd+j14vyr4mD40SNbrPiBmPZlap7lAFPXCZnwpoq
ts24nl2hsDGqcqUfYF6Z5qT9qYsEzHilOcC7CxKSfUMBiFiiTlRCyJh/SuwQiAdg
Siaw/c0Uy1KDpVnKlezgljxV6vUXOn7C4p9OADO9PI3pOIXbFJ0fx12Bmnkv0zgC
jGrD57jrklBsNX9osphfE35+rN6NGgD2eKBsXa3vsYXgQDmAyzNwNIxKRrQykMwR
7V1X5ZJ5TRu04IS+odo2DAe8WNHUfgc6H6B8vJW1KvjnprQ4+KYpqwXe12hogy4l
LcexjiXrPnukKsTjmej3arjE5pbc86hCk7fFXdSy+OFrsv112xnFrqtbCqpbtVHg
9drY3UHn6cup0aGuDzixrDBmA23eZvw6yIo6Gxt+vGFk3r9wkp4wub65AjnKG8k1
iB6fStyk6fTiTce7o1vF45cqWr+hoo5PWC+2QKo7ZBZdkaFBKiqvxMQDYo/ha8jI
NPSQfSxTRqgX88PEDC93JRDMwQwAfXMR7OkEuysepxNsJjPb1rGPAYtNioJaVLYD
6Z0+BSV5FvJcT5mZrE922jKMcP4RxEX6CURBW9/lhKKPcFvxXPYsJQbBesd3I7VD
wsj8Q2OvZDMf9f6mt3OpcOZmEOD6149pywTDL3N2t/VHpVeeLJXhTyUHM2IWMqdR
Bc5RA1M4BSZpcZ2ECC+Ju25F+Ubwuj87mtKHP5fgMn04EynlbfKjZGiRs3QE3UuG
OMeCe37Av4BHbOVXKFYZjT1Pz41WV27X2TYUav65qMGkgXQlzsor8Vss9dh45eqP
6Yl0R1XEFOb/Jbdt4u62/pFN2XGfPnD4ve9lqU2O+ncc7fl+FFAAaypzMOzKeuy4
Ea06BYwm9sBg5Tup5+/AdpkrXyT5F56y0m/DmUfyHSFyvpXEIDyDXcfTv7dqdWb6
mMIiVjyC2yuXzUL4R1yXGQMfo+h+8J9vNkYI+XRjIrcc0zm/KvJ5I/2kuCw3wdG9
XtsrKu8VPMzwyFURRirs0FinGPcOYll02fOcMe2U7vNkUL3EDEKesXxvWu23rwf1
ql5CPzg4v6xYSI9sSAwGTsSZz2DBFiB6XRNOX4Kj/8QUJrkUmoLO2mzBJmjoCWBl
mTn92Tnrqc/Kp4PKtHUSSLuJzVGC5ccgLVMxfAUHKhJdTP/xWjXuS0PqX6sMjP2W
umdwERTUk9ViUIWIt5yZpaFwkTOb+LBKQ5/sI97CjPn80pJB+Fk8VR3gyhdWwqr/
HOZ5HhIEJ+o4cBrFFKbQbBjIahBJ8kXCOvSPrZC0ljukURC2XYHyvBiClUsoc4EA
4Ex0H+qSbG3Jt8sfHmBAlj5HSsCWhdsyH1hPDNUkHgbKEoXyXSpZXnX/jbnz2awu
VYcSFGOxQAjq5BexNzbalyZqZLFQ4QJ3az61B6lXDXsWKnvXDTg6BTgfTqtDRAfw
/k9sDhCsyFm8hKqod7is0/fCeby4lK2lArwBJ2+MOukCrk0jCHNt1aaUdQAFlxh9
kUkX4soVQjWDuvmMvoKP5+SSaE06YDuP0KVMwNV94CgfR6+DySglHH9AmDwXVMZD
mhONeiuB8CSOAVCvevyJ40oOU9qM7Jn9xHP1q1J7k3HdJcrbZSbQXS0+apmyrJ43
O0EJOp2P1BCYT9SQDdP39KQhvvNmTDalH+/9xBVV8UWgfZRnt9UXt/uLYWdzAHWq
UVAOJWPWQH23MLCyPEJMw31oG41tYE759cYEflTTmYiqX8sN7V/wux8kBpnJ0bcJ
XLvs+0HOjJV8vFLU4Y8kZEu4o5opnHu7cvieOxKrEf5/YdqOePamIKR1Qbr8vP5P
tbvWp7gMyg1EU+mW5dArl3Cs5JfB8jgCU59zjGPw8RX/7tesdOBQIuga+272ugfn
uwRq4YjVIh8RAcHZwSFLAYQtJZx3EBN1770hIG4ckRjlKoP7U5dVmLi0k7fv8erP
T6HRBReG+Al0vCFKYDtmVnlunTjkc7ijW1I8ErKmDIBSut/UQSKwHkZ3uHTZ5dOe
5z8cLy4a4OkOzSYVKMA6qRPGrLuc65uJTWu9pxxe+LmVVBwMBUDfKvEZyAVRE9jL
7BB/8eY0BrkGcVQJqIzJtbCeRfvQEEAl08Btc1bl1V+gVVXZp0ioMxeKYHBzg3kG
1Aa3pYxPiyoUieywRSztQSx6FJQxf0hKubBx4aQUIGvm75i3MOO2GRa8SgQNJQTw
f0O5jIxkTSxfHHlwvbL6wc2AigrKfGJ7wp6VOCyoTRJS/V8PM3GjtXcTX5BAGWOS
y/a2Jje6rSecCEQ38+qfGvi5gSPcHEocVd3Zk2v/1xRC5Ci8wTr03HG9B0yl3gOZ
XCrP9PnCt4Tm7UOL0/fHWz/ErF20TRfYUxJIELK8HdpkdysL2vaUzvmMRD7LaLF6
6y4iGALGlhs3s3FEyyUWMzogMP8GqVmRkuFknKSboFfc5O9v63E7yXpTw1nTAgB3
A2M2ur/jUz/FiotSv2XpU5bO99Ixj2RF+BwZPqibLte1sV5tv4RKrljh0pzuy9U9
FvbyVl79aATEfno8KTjaXtAQibgTKjCSouPVrW9PbL7VnRME7RaNME1MpQen9Mrk
uzxj5iT/9ElRh+R239x0jCWZTDRFL5XXwZv2G+XSqEeLXnYGs6V43/JxtvBo2/yJ
+G/DYSxiP0lHZRs30DtRo6EHwI3wkAxDJVoR3PFLHMTsz/1kFUvu3CvwlcVhRpPP
ijKManpA101uYtteXZp4aeeQLH4FfkBInGfpzDUIbAgcw1WlEZ9iWpW8wxyarFnC
cU1iFc0A503++2ez1uQy9mNKFQ8Ta/8A8OXkpVv0pTx/WfjPpEJ9AXfWy4U0KdzM
VAu7u3wwFKTj+eAYiffq54Zfl4aitIyHV6bwEQ2+I7bfyNHSw/2bCLvvA1fZCsxz
erCBZk0HPgmoXco3GeHf0GUjXo2oCOxCWBkqlhnc6mfRA/mcpl8n31tfiKg7/CRv
/bNEx+Bet/YcNhTyvDA2VIAP+POvnxG2aHsYx71uPQK5lO+vJmrpoqEjn/+pDv95
l5AFdSpYhBy9wU4Xqfd1THM9Z2rtBw/z9bZlrq3pKhXyuJCRhen4UUN2ewFebj9p
etZzqvD1sB/kcmhOYwgbeTKlcjrHnEwbRM7rupWfBvIH1GpmR9OiiB5gINIVrT+d
NnBbwVeXpEqJ7WY3/9CRtIpfhtNINaCTD3f2nISuZOcM7wMseu0u02NPtLh1/C3J
L6jrVcvTli71FDpcM+JI0t0j2H3sy11g4pxAva6wA/tmlsIgSGl+A7oZ23aAWrkc
B+3DzbqApvaiZ9mOkovMOUTMUwys8hQCHkzJaS74jeIT7+LXxd0qjdhFrdWAWJn4
XYfLhsbAYGYKVrg8Iy+REs+qpyDuifN3hHQ4oye30YPZcuVtJhRrscXlAOt6CJZ3
5kbEb2xF6KqVZ/a0mvSniN7Y2/WpxsVSX6k7LFPPOKbKveKzzItN6E9BB4tZzwYB
unk+hlCnI2uIDRpRBfvkU5OymuPr/0USHOZ6XhMJL0FlPyHdj/ULYKWdvHiUauu2
UvsUyUJQTzdnzRxVADE/IUSSlg2w0JEVBd0fHBjDG+BKKKJlrDHlxqp1KsIYBE79
cYXLpHqnl8LDt6irRmJFXwf5/i6ZFk27kzQNULCh4SE/FHVBa4ZGEPVQOqKNb9po
tcqkDUJO56H6MEVSO+Q3/NS9cp8cgxcZVLyf6Mi5ogHtfB4K7ITi4Ns2cEE6MOtq
YTOloOwKt6ffZ5UnQv5d745Hp5S1Ft82+GFAW0iMoNzkXXeQ0fL44iLIAC8JEYvf
inryx6/6qStcfxgClz2k2ORSfi+VejVFEAhV20/b3t10i4zayEEp+7gndWZQxWkO
8TRdoDE4m0uKlyv/pxep0M34c75yFlFn4ALttAcEL6X6VQHFRQjVJ9mtQcA9kHk8
bgDieDgUoyH0pK0P0h1LzzL84s5PjBMYg4wddVQ8ugxHCQMRwNBDhj34CKWLO/LY
bJVzRwoo9rST7BGv1z2UHh+AQI6WMY2+1S+A0DR82afWTRo1tCayhZAAwbToh+lr
QsdmBeVDyWzVcWYbVzB5Al/lSAnGZrjegTeqmWgy+LtzecF9e11n+xRLqTVuADeX
4BUm/1K/8ESm9YnW6zGaTFlRc/aeTso59V/hPGwn3DFgM5SVUN8Akn8gukBMHZLl
NoBgm3q0Fo0kbFwvoLCY8EtiETapgRMsCasob6d+qAOWMPfxY2r+6sfeewNwJqeT
EalgYfuxXT+7ysYsNQln+bCG7+pPQ2Mk/N3k+A2G/cDF8ciiahSjfGPKuVmcWKpw
8LtMZSNNY/SN6hkjQ6+xahMlfK7FZrgHdLceyUfg7XFqRY5k4ld/NlsQV3luCPhM
BiwMJaps1+QbaaLlqX0CRhqayLn5Dhg7bcq7JA/ERgONRgWVfhXEtM2/PhLncX6f
6r1ZIyUJzDm/aX6aJJSySi6zaB9uA8PvAVSmcSGrJwcb0CGLcJ9ecEVdaoevSUl5
0f4uU0RZhFgjzBPAlDniBGif7O4rGUkzqoOI/reFJfhsC3+aPr/Vla7WnaY1CE0U
tnydrrUPY0EQQonBtiR4kiHMoDDpkoxLvUjSuOrBnr3CygHgtuDf/T/hw6kxSxI9
iUm5jSjJvyZR+M7cSS9XnAc2ODzjirXVaPR4YNnC3eLFc4VOqj75aQSiUnignzsg
jaxDFf4vls7S+JvzHJQqccsS7faeHadu6LlQNG/Q/7yamHTYfnrkzngLMHGtgog7
hG5/NWDIzvuVlRkmtnmyQ6udqFdQu2vudkGmaP8hb+lDBLrAg5uX+nSARUdUhq3r
08N40az3SJ6FDyB4sqyL+pHsuwd5qDcJtBMjGNOSYWm/B7ocP54Ej5isIWPEP9Fx
f/bJeUWmGdP448Jca53zPHgO9wZBaYSkYelfXtUetp1bt9ZK5DzPcqJEe4moT6G4
MrYwvyTtAOMijc84vdhH57qs5YlWgOS8A88HDxjkSf0KjXbh0VHEnd5oe8+wPOC/
StU7451iK/T8PhI+MA5CngOSvyjfpZQ0MAYqEupYHPMxtZX4rKl640JtGE8muUKA
lcuu1uOh8LneVlTJJaIbfIFlrr1XUU/px543McznSh8PWI2GP4wvsLvalzgCfVVx
Si2IyD5PefygJ80jaYZj2Pa8t/kDfhKUohYyF1w+VcPoXvmLYg3EFkgPgsduPK8Y
gcqiSoOiDEmJ4LGzxPhIv+bxiBuuDZ8RWlfA34QswCgfCpzkKX1tqu6t7Wpl4uhJ
kNNGUpc9t5jZZpB+jxyHpBDHzuOsbK93N09w/is3PsVSZB1ULx3Rmk9nVXtSQXaf
ostn8FZ7f1M9inIBSpmMC26l5aW5mVhSH4/pVZRGvFa9UPI9V/m2Xmlid3Qvcmgh
ksP80bZqWZVpHB3tNdo+1riDXVJvId+j5is3HSjnEJhVStTRyT99r4Q9Yd4xSI9n
GkNh6NXN8eMiX7NB5P9i3acpeMzqwtvHG7NIAtO3Mf4Eol52sdQLW6YP7i/JNbmi
S3VNzou/IRMO03a4JSUsTmwB12b8Mh+ImU2EHCYTmgxkmTQnZ68YW6AiBqVfDpR9
Tv8AM2KnQ/dQM63l1w6XJ0NY4OdQfbcufmpiHeL589qwMnSQ9LX5z8BwS7cbhOgW
aB8U3IkNnp9+U0kuNi8NvRar6C+PUOwZonG0l2U/B/Mhujtc50kXxGyqaEer4MNT
7gPrafk4BSyUcEOWzljUpTxAe7ELk/anRuEflJ3RB5urD8fcdLcFLpYMiDtYtWxw
4j9ziunM38Qv0ypXFZoWedpm4kVpHhUa+OYqU+N2olSubqGE7T0Kb+zr/9XiZaSN
3X5RxL1YILiltzn8nm/LQxA+7FpiarU4HwHML/WokYBCuYgRBEd775xdoFZSqkF2
YVx8iVjJAuvr2LYQoKAe3pRroDZCfnAM/UVCTyBdY4uOJf3Whln4Kw44GTv0bpeg
atkx7YlSj/bJ0nTFBavL8zp28rFxpzYjJFxdB4bN+90TbOenLULNVtb3np+aiM1n
QEN+lLQpNsQSyLSAPWMFiYEY7OhF/jHSU5wARUBKsim3iNmejWOx6otlqmY2co/X
S7xJjLFidWr35W4MPqbLrXEif59ocbidZcrWJJ3tVSx5WOo2OpWtExllA8LSF4J5
6kfORnPjjLRLoY5EmxTivNVVV9+0HPeA9x1dr8fh9dxKsMSG9Q4uShBgse6CnqzU
Rk8og2qkehjRylWzOGhp5Ec1TOHlLaelbiZNYjkcXErE0Nc5LV596TLCdCL3dXSj
KmyZ9XW6doG1+/F4KU7X6KP5A34BLyYCwaehNsANVK8v1fekvrbaRkEwGr4uA/zY
/pj6plUTyNvGlluTiZK5RK1qoQEeYq0uSBbJ2YdgfZHJIAvx7fIpfQ0rHbCVFdZr
VBQmyV+nz/V/299iABz/w0XXB02dNFFAUgmIhrVj40yc/8AGoQcmqHXN5weJrcNL
7fLgZR369Sae70FiOsgXbQ/MJF1k9bm/3RWqSXd1MV+JAPyab7Fyzmb1ryehwiMX
aUp349zfRqylIJcDTfrdH0GTyOPysd8pK5O3e2M5RwOJBpR6GgXWOcMe+qUJCUex
OJHmuEsXIY/wjuB45nUNtCNC33xD9a4rQH25OChZJTOJs96ATTlqjVuglE/+En6w
g1WW/Lp80/5tMK6CKNGMlYPqOzZ1izq0M8XTZp6U7ostsrbxQPbypCS8nOxOd4sh
lUcrpFDOmW5emWzoVkaR5sPY33LnNxiihSpNR0EASAeWGqUSd3bptcorH3wgxPr3
VWqHkBcW29OaF7dvcrkMGl3qVYI+smhZOhIjMlO5IZRcTI6CeC76nlXsO/npOkc6
s/7YrATCKMGsLAVwsR9tNgRpFPTOgwuJgle7EczUa5qquuoJ6JFd92ghCXHYCEZM
+a6mPsRaDs4Br6kPcgUv26faxulp3V/gcGZ7NnPg6RunrosDgXraELFC+7cwbidZ
puBkMGOBbqNlycl30lh0gICoFYg45G6G5xjG0C4cNtg4HSfKPghVekgSOk/9S+H/
eeIDEq75wEytVgpbS493nQUiE9kCjuQwnU4wm4q8T1Jdcz1dn68XCQRK20TpDbxP
YKgC9jhd98AXBkJxL4oV103hVooBvKSxwr7iMYrbpWtuVUg5Y7G5EKJi80+yKgIc
c4jmeXkpV49Y7qAy3qfkIOAewje8tnYV68GM0/N7lsYYX9d7eJF1Nu/vXxHAm38e
hJJ5Zh04KrCpcs9H69arfNNjgxSGQxpnRyzaRBR1KBOMer5G4KVeZBQsGAL8lPib
kynXZypthFKdWLZfAI5D4PpeBGSAGLxh+lw6kM8vYPZSI1edtP+wdXCNs9EHnYhQ
acD9dOWLce7cZJoIwiyovDzfixDWSq2mXP7JTjwHTausri4LGDh0Rxx9CGDi4492
t9qF8n9gTMZDPuFGdMGX0V+tFhSMmfyLKsn6Xn22JDOytDb+GngeJ+EZN9OkoNyH
nBD1utcCcyRqwrFU80F7fvvTi2+MvjF+VE1vkw5XQTuo6eT6NOLNx4pwIRWfsQTJ
O4pnf0BRldYN1+R0AT26EBW42GB1lw7t0hhi88AErh7Du8RKGUxy3LHK859zZc5u
EKV43b0gZ7l74liA+k+ShpTQOu8DYOLIQWcHdD0GDNp7c2nTLoe80s/zbCIO8o7j
J4ogeikhWlGi9a0igwYGqzq+MVcPMth0itnbPo7ht6jvtkN+5LZxne9XYQKrOXzl
w7uCeTxpeFSJ6AabfWeVTrh2glkUUMMRVUrIoxEsvJMFnV5fiJ41NOxIRQQvPFch
7ISVbx99G4MAocTi4GUshUfwK02TFN/YN2+AutEdAZJ0hO5sN9L1S4liEwyFvIpK
RTyoYgAFnPGDU6sLT4MCjdwFzFSMArf04Mr8umMnBmXMc7txqONVRo3s75yyJhcx
88oWdfenFtM+TcXXJ236Gu57eFqwjO62/f1dvjW9EPiKJtXOXmLfMVvz5Nla76Lb
ZWkBC6bxmgUKCqBuPX7p/Phuptl+06odtzTsFM9goEkvEaLOm+M1s1XsKJK/Ao8H
1fdFshzh/AabQv9AawY0JTZQhP/uMblBVxgsh7gw5KpD3s9Xz7a8A6thxy+lN4aS
lGmbFkY7VF+/AeB0R4LXJBTaDVgdiax7gAaG4+k5tykiKb1QnVE5X6rw/0x5ZKL9
WutKrD58Uzx4BE8I9a45BjSsEgRhdKqKQoIafZSpnEGFjN7ws6RaGR8KrqKwZqqw
9m7B8RSZxbgbqDAcUT7FlrFUeo2Iv4dP9wHJx9Nj9nvNVF3uDan+8G1DpvKG7iay
xKB5aJKKGzFkuhd6UuJIXEi8+F29DGTW1b7cXYzVzKDz/GV283vKw4v4PejOdnbs
hGmYXRj4YaJ4e4MxWvQIbUd5e/iIDC0DWTCwtnSnfu9VeC78KDRzp5pLtlmu82OG
bm6xAuv4OyO0oDLGwLc8p1qUILs7z/aE/eru8/tj23JEkJNDnQlGUYjbQWLw6vME
2/jFz5Vr0Get1tZlVAtz8snIOlxwvUJes852xOr7xPJwB9mj2LSM+8qyhdJklMra
Yp5qdzfVkr0blTp4lV3nzNLEzPOopU5Ba+yUEyPGs2XlC/bbsfw7Tebdy7AFWRXX
jkQ0qRJrMyomZMXqPoAKqDkWKO1f41vG3+KSTa6ZfJwFi4gXfJxYMZea+TEX6RnW
d0ZUPki5nHZ9EiXuEAF7gIgtTpoea4oqpm0HolNgBFBQ7SEDk0zXLgEylPwi6JBX
PgUfB1mcDKLyDfhiWwxzyQFPs3XsOOzECDt9KbHDUaDorr2yr9CtnlzB5/J5rBPQ
/uKFiQGQ+CEmYOaxqpwt156K86WylajXO0YubE5MY+bADAC0D73cM/JkuBbGfPft
S4kSzWai9aMuuQPIXj/kbBnpHcivFrAbfU/8v0bQ93/1nPrAi6gMMlp4WLgyi1Qa
KHGAW1hGXui3um4rayRI6uocaZoDo0/PhmXPHnT3UJBPw5AKtEye0UgbWduxW9UR
pUtdxSNxBuCRmBHpSKTFvIbxWyfwzpxboqUDpTumLzahD2e1ytp6Btw0khxKCyWN
tRtG9yz++KeBKjkuEMc8xrDo5IPrXocHcTt/1dT/YJhgkZLf4wUXSwO02vfnO+gJ
UiQ7YYHvpRwhX903MmkU5JjT8mxEsVw04KbhfZA5NbmKlHn2grC6zRqe9Zr7+/t7
awBoJWQx9oSfwSGLU8js1KyDJ1H4Up9+HrwS5d+fic95xrBo+xpA3colOzJYULie
0ul+u/xQCtnW/wRlTWIMWVbjnTwBcCgyX7vYRli9bnsY2pEXsqkM2WIzRtapupb0
O1+1I5oRJXpm0YF/kru8PyL+KOeAjXLSInDadzvH1ny7wyMpnW1yl6GStgZ8Tk/1
6CxfR2dqMvX84hfbKRHJ1x4IWpWSRBMzoGXS7QG2xwke1SeL8Txu0JTZjgorgAsF
OwU+2d2Uw03BGB7wJjUF5LXRuQC23I4Kbce68OJob3NWBlr02yatDJqx3ZQQ4rwl
eOB5pQo+akZWIM2S2Hy5JnTDuVFyMd49oxJNDFn/JIiiSoRaphp33l6N+GEll9+u
FoIPGUthYuM2c+iq9pdk0DhlHrzyW1W6wFR2rDwO+G/iHavKRgYHEc2c7ngptMQE
nZa5SRRz/xMCrDw4ZzbGaT6K1EPG9BZbonZL/vrZmdaB82DKqvj31mc9Roy6gW3C
QdS7kaibSnG+eQknlHt3RUQvkqGpihHJ29Gez2ptDJAqU6oNrc2X0vVRWv1La6ZI
P7VUtmlnFHQj+dl+hubkXUl3niHKhrqyfrjxPwKRSZx3vWHtJuAaG/W5GsVPUApH
ITl4wZopYIaYK5x1SbzM5BjIuzX87fUYAgDnrcraGiN9dOjoFZtVJBFZrd0vG9qx
qq5Et9CoctTRsb2w1wTNl0s4PEISGIjpDEuuqlZ2pXSsiaZ5tBEl9P0eUEERkUQF
HSVRr1MMliLGnJyWCxz4S4WKgz9SmGsQQRPiJPaQjZan1gNAlEzvP7nHfzdvP+dg
pUicPPbLM54DDLkIm4hRL+kQ4ecrFsMiRCqaq972kD3ZGL3Pmw59/7TbOXZVRU3x
bmvJOojQLB1GzwmQzSA5FhCJiXEBfr3nJdY5DC7efF82dxXN2qkhiYXIgrvkQN7A
i4OM04l43xbatAzpFtMzgUHwvtpX5QoycCW0IhfREigXMhjiKLr+qusWbfaUO/0z
aWAcFyhhrJIbTO+UsA+Uf7nyqU/JNF+B4hkGQgwXcDDIeQ2YMZM7UxLs3Rh/7V4Y
TGHjHkCyrg6Ai0ZDnz9VhHwRm1LQBr71MUAmjPEUHI0itekAFCJBosvZ5ZnElLIH
RJe7QJINU8OtshTNPEeOEVWEXrELSjXU58br49MFtz4MrLYA+kQrfGQpJBew4JUz
9h+lrflw8R4Zh5jaTMy2gpNFXPsUQ8URuNS7EVaBcSv+RE2nHYjVn+z41Cfx1LTT
ne0CCMkR6JSvpKwpnC/DLd8ALkDj1Mkg9UbFcUCMALD6kim54jz/QMYrmXQ2Effl
lIc857MhON2PkZDTbBo638Ax41/1ab4rfsLIhqTMdh00XF4WK9vx4H/1hj2n3Fgl
Y2RlsMENkyRQtEuAW8MImZLyOINctFz3mUjxTDgx7jnYqmfW2FXsr5AhIc3Hv7yD
j7ivPy04xOwZZkcJUFSZ0yK0G/ZV/RJVQo+tbOhjz7PFhOKM+7oz8UE3Z+BxMXfj
pDorAezaS2u/CvmOXOsarqw31JYcN4BdKrLdio73MIP4AHZ1uGxpjHyFcI7aB0vV
9SwJad4Cvgd60HRLff+ZX6pN7UN6LyzQMUSDjQ2oTLtnn1xOizHoBe/YMo7lan1z
3Mcg0JbsI4I37F5CKJyJK8Hpnt3eoF2t0Zy0jSkghkv5A32spfJgwNRczt/VNzew
CQeng/cvelNl1utwCeYvcDNER6lgRF2v42xHafOuRiejiSvj36s9EVFZM7SWPry/
ziZvpjNIR6I8zvtQcnOAREvGz3VVbP5hD3AZ2ByQU500bDqEZWKEkD8R2dwQkbC/
iXULtPwNGBYSzFX5EkQIa8xFh7ypNvyijRC+PlTcJHaEM8kovS8E1DiQRGlPP6yu
KTYPILzZyuwmdB+CSKftaYBf6k8ucnWDL7gD62OnLIW1gegzFAxBjmM+ARy44bRP
kuNzGaJTdB1Qf+Q3LzxJusxCeFi0qZLrbmJCn92OX/LcwzIHiPiRaeHogIPDBnpG
MVtMNkVKW3uLq9EJ1FPMOUkrSQiiM4Y2yRqOlKpU4RqNYmXXR6/Xw6cCrUeEnwUE
DzermrTdaifHU+SA0kW8L2l52e7V8fXUGg0WBy+6XaGlfNV/yhItBbsS459+Yl7X
45n6sRR9RsB+y2FdZSmVlN8FVVs+HKa5nzLkaeH39gzCbRO1Hesv3qLoh8XbO0SG
J+3ZO5miznTtQ049kOHpylR73ydPX0aAcdA035SiMRbQSyJlpf3+jRHjwUdR+QfO
VBlpX8ENoEUBS9UiX3KQJo+BoFnY0oKliPxPlHUfov5jK6V5VkJj0zrouODfbzyl
ScnEHS8YEE861z8H0o8nRbCzkbB14Mfj8cAVPbxcTX96P906/kvC5HYJXDFW77fS
12u3gi3iOwuzuxXCAeAcmHjQVOpP5VzEedIE0ZI0BhX5D3BFHa1+t6HHkhRf7Xrh
uklKpmBK7wIf4vTsH7xbACwJIVbDMMdwGlcaLOTHXyFR02EC96kvqXEmdzn65+lR
A4Aq8c5ta19qQsSg/uk5SHyPTT5AO2FRyzCnRsWYhqs5COmiRAubLhWcDxB4on1g
/1q823ZibDzoEfSLUYnTRKeP95q12tYdDMffAs4T5ypzaY184lii+8AESc8pC+xU
3LBpMMpGi4F7LAGpdylDm837ru9Vy58OvL1XsJK0a64AD7Mkx6j5Tm3zGBvnbicz
i6EFwNK1j2GTNbYiVgJuHnThuXIVDg0hzRfB1ovuTkzXBmZNE5VFea9Llhm3FhJG
sHlZlxGbpJI3ii+gv5ij1cSY5mwFT1P+mqVjr66XneUEWJnrACcvlX/AlX+RPe+C
FBvEGBI5tCDeF6sYA0JNNSu0nJ2Cj5x0ZY6pTvVjP9W3YU7DMM7b4FpQ8MHYcas+
CdoLkNEbgc0qKDvzp8F2jar5KO31mCG3DPnxlNqwaJq7eDwnYydX9DURcpsZcDzm
+H/xXCJewWABka7HVf4tm2K7lp1EvqJExKzubCsP+sBXa1d+KKsGgDzw6mjWw8r6
GqZN0WnWpTCd2yQf9M/FBjHhVVxUcXZwY11YHbwaLCQtlUHNz5umQxWM/6LLpKNS
BzVdsNViItLTUCzicYrHFcpOiJ0C+2yTTMU50YOGDF0mxM5kEr2sbjD6yJ/dlUTm
T8FG8Ou0dd18BO9zlsLJHmcpOwVQGrob2JEbmVwK1dFK13MbbUMWP5XTrgef+bV9
gWTMsSKQZu1Wclgh3KQA2p9llaC8w5bS/j6uSSY+0ABbL4q9nogJOYGRIeYypi2b
I9i9BIh0YYJIr1UGP7N8VGqjtXxGVx4i4PLEGy0/46dfCm/r5w0EWbRRWgMUzjpI
2HHip6WgLxuADtX/3LFwW9zD5NtHgybzIDdKBuCh75fIultyb/EKU9WenKabPR92
KyyRvLIUqLgh5w395B0v0m9WmTUctEgJ+ApsvCmFbv6FPlwoezhRxEYvG0sR5qan
gdKsr8zwo3gcrCmF5ISENMB5+53V77fRHrG3SKRNCmDthcrDNJQB+2mCwGEUncDo
zW4YgDfIaus1Iy4DV976hsxnRtMbV/aY1tp9CAbU+lIj7am9iZszp/sR6d9YVSx6
q3sdpc8gEY/ohHSBsaenzHIz6eUX3uYUApGX0byQbKesc2f9HlX0oMpOl/36Zfct
JgFitEWZumgpsztOSsIJDdxkW0HZC0REiNWq3HjVG+ycopzZ4jpmFgYGpOHgXMty
D6ZuY/rz1FBw6CIhHnzgqOm2u3vw2QuwAv3hGI9QOgy8dBpDiTLXcu586VAQf9eZ
o3T1hymaYyb3llEIXhOPPmBEACgu+tc26v5yul+6FHmDVRKy7DVfWg+nlifx2FLq
EZtfjIQG2HHw++FwyIaqDlfwgfN/OFGBgZz06mRXHLc7mcHxcSyfNHHBIWAYPl/X
3DMHi8T5Y3tMgihf6/Tki5Smb1cvFBhfy+7duNAtFV4ANiAID9gXG5DFkWVYEn2k
lCtbv40sp/RCci+0sSoSYgGwF7ucMHaFyJIVF6nYNomgB8y2wtPePb72BRp+HM7S
p1AI8DWVksleHEHvH7D48s6wxemCqxN4WCPaIBVwqt95lLkgKj2cP41e0f5ern3j
zDycs1lSYsIq2+tGXLIKYbf0Bl4TKiBt/KVqZS2KqFOMoZKzL8+q4d1yAlblOuna
beAQeBqFFO9JKb9kSa/4wIsKBzjaSUbDe/sdKN8Eq/AnXfE4R1NWOTzB2tB8lGty
pJ02zHdwJzvyMhF+jWTOCVmLQ7msRuBcvrZ0JDm7kg6j/D5OSTca7uczuhKS1Tlm
vQoPNdQ1KA9ihYCVwgh/lMmA6qbSp6yYCe1W9w0xiqA4Qz/AQFjOZEK81aco8kMh
DSS80PCTcBWx070FdcbuncFkrmnvgUHMOptNtmoW0dADzITjvUkgN8bmnWvKvsrT
PUtvy1c1hKwF91wFDrlrhIrT8Uu2DZJ1owVYyf3ndy/LUxBimqwe7HIcYOB/BvJg
zY6BRwwwpu3naRW45O22IuVOREzAPWHgSuCpyfwsb8zqFINsGVC9YD1T4kzght36
72xXElqoyceqa7O6DrCEHVVy7bna+PRoUa9ShCkOQu8/4dgw97NUeZ1e/hoAns4z
enV9/Uy8Hb+rVVbvOEQy5nERxSxma2VAfpnQG7Zk8/pRoVWGuRZ6rimnHE32/7sN
FCY3+DU2ASyQt5qiTMPKxRaQtyMFWUadyZQgZbFqd+sI9DmV/rTqiLFQo4OwrvTW
WI7mUPIc+acKQOqCSExeHN+5d7DqvKCggtl1TRfliOCzI/91C7hTSn611qLydZoz
Xijmd1yKwjFSTwSr+cdodTFzIKNuAFtwfuRU57mAWTirtasgoqrUYbYcoxk8LuLa
/6Bo6NBGmAKwhKGKHL4L50JDD5u0Mz8CRwViOV6O3v0fYnF4xXkFs+Q1lljsCMoL
twhHCuBiKuBs9QpEZ391CXKTsLThrvHfw1XI6GeGZe461ilTdFNgB3wNFhU8qFkZ
A4TMmiukPI2jms2dja7eI2lv3l4tcroCeEKtSRKOGuA0jk3mc2xO8+TS+tA/qlzw
18a9vRjJyCWTLLPpylWx8W9q79FAxKu1XX/NsRCDPlWcJ0b7szc6Tpb+7MpoC6Am
skUbXndJ0eOgII3Bg+8UHFEf6CR6GzUoVFJfoL5YwUJ2Xq1o2ZKGm062bceCcwsG
Df4blHL7UOSf53mDbQb45uMnx9dRtSJG97V0qCMWel895/XdFAKPSp/pjfvOn4BJ
EGDw2BvrPnwr+otVg+zaQlIYYGpWzXImjImbYI8Sx1jmCFA4eOoU/RAerDqaAhfk
k5p7uBtmElZv0Fcu6WCCeMGICfuHN9w7eZe194cj6XNXo89ynByA8ASCSuY7gbis
3e6x0Za85puzK0NXrDDfSProCJkvRdLhg71vZoHe31iBiVj3jtTBNcG6T/ZXjzYT
gPxt6rvx/1Omg+oYvErlhvq4R8OCSo/ZYsrrEpVlwZO8Vm6fQ1eIMgBbVHiO59FW
uldGiqmFAr/nlh1VFDqHtahDf6gjQQ47rEGL1jarHs+K/BVl7oA0U0EG7/iZKA7U
LF7KUMIyWwH3WrBzSihbbGmNllCYUghTC41nbqEDWwhH+Og2Uu8WJA9GsozgVWmR
FApfGj3wnU7eY0cKtNn+Qoy/RIU9JTavzU0ECZTQ2rFm1rXOujoiDOyq+tb1zdlt
hSXrhLulcOTgJEs++eAVXSna46de5vtuGIJ9PIQsR1W+GqWQc+jJ/voEidwQ0Y60
4HflDxrdaqSCE40RcrT7S5jreixHLsgMTq+6Q2XmiTy2VQSDJ3i2EgM3klov3Wvw
DG2VTs7VhFSukQqwkYt7HY+uo5X+E8CVxi1mRIV4DHVprawsXBySNrneouKMiTzS
WfzSRhPToAsE/HoJF0exu80Ji5S4JQE30z7eUbNQxfhFeAPdpQ068T8XW3PuuI4J
8jwDqOzm5ycRtZoODTeCTbhLkOuVqMkQI3AiJbUMpNvfFmBptwtMrVjV9i7/OywZ
0kfH3v5fCkaqJO9ZTDTr9a4NlPDdcp9O/nh61xgDyAu7dAeU7O78TxdfZNkbrwkW
fgdU9j64r7BG68oDW+75YRo5K/BvvdA1ZEh2Sbco2lqlMXNKI2vxzX05du4fvCaB
y4tGosL55HOdXMCwLH0G85l9zmMTwihzlCj99Uol4QlLFiHGd3YoS/Kwweanz9P9
vYRp8TB4RkRt1gLeQE10n60UEKWRfyRTUcMmn97DCtS2+WIINC8fYXf9ikZ5474Q
juW6CNP8F3UA5nVojgmOhpfX82DLdQATf+X2JVOoAdklFT9eudK0ZxxnvUAGMkSB
4n74pw6YTlTRKwSzjzcx+WJKJeglmQdrukqQKap3dw2wIfkFeiIRF0JX2ktwsStx
ryvW6BdUdo7lTAiUjCkw28PvOcwZq3lEJ9fu82SKOkl9mKyhlyG3VfIieOX89op0
zEXOPyP4edWTBcMEEFvJtS1x7qS0lAVpOqoLlRy0UCKlL5f+Y94MWPRxGNNY2Orw
TBffGEWhRNZvjEN4MOLxL5W4h96nDF0Zl+VlDxb/GOA4asDb75UUKA3tLMNR/bUK
o6kNQM69nV3hbYD/1/xUz1JjWclOMVc3Xk+aIPZ5slyChfSLGXd+w7XyOxuirEoJ
5WJosycja1f+EMNKHIddxAE6I4vVtswwer4PDtaruUtlw+cPjSbWmdubKSf9P+kW
a24o1RF8f9ovDSLRvgzckR6JVfMoeJsWF4i112El3tb1KeyYQ1H6vP1+OZKx5dtQ
AnIesxlqZGWFN7aniZok4nziR6m2wmJhjjJATFA7RcO9iC6XIlNKhbA6ow5lC5FQ
giS1mVwCFI9E1Qj6yUDrE4J8JN6sfy54naQxzJEO6HBFr323z0aM2ab6yy1xCPkq
wO8DhvYySO2DUEnhZSvsG9itWY3lM+xUi3OAEQt1dPG8VUY//3g0lVjgBVe91DAF
Jbz7U9eGTRDoV36e3+QR2n2+xSICVBQU2pLYggHFJiIrF8LMmz2ZQrRxZ52SqoDM
ZWp2pS6rFqaehHib5lPjnQrm5xKfhchIozs7c/gBaatLNLN9jgSWgQ8ZkZ7+CrxW
D5+YwPKf2V4vfqn4+ZRdLauE76uF3hHv7PmRwwsB/b2OCf0MViiarwhFxo0h0gG9
oX1f2vk9vuMYEQAKxt7ctuemUgijE5bR95tvB3twniXGhcVoS4jYncAWGoUl/RlE
Iq776JE2ha53h7A+nv3ASWi4+DmNs7YZvFDx908fc2NAi7I1qAzMX7T9byUJLDth
CIuyDHupgPfAPBn4r9TcXcrnLBte8oS9b5Wv3bsNHpmkNZMR7D8/glkec1yZRgNr
HafiVsYaM6o3+EA2dOIyLaTLoqHeKNdgKHjmRIAX4lOY2bUSCyPs6JBllJZpkQqC
bPrOjcSnPyeNOYvIJHYqRNN9UQ3Mf065lTh2O8xtwQ6FooY4JpjK99SkUjcXzfqL
nqTsPD31xOrzdiVWyaTCCCjIyxUpDgL3FhN7Na6lfaMMoOlwyBhmk+2Ul/0GHByZ
oYRQb2UeWKPc9r94+0vN4TFCAO8gFf1xgLxmZ8oCRhMr5z1Jlty6oP1vuSXNHQvt
6faVlMMcCCHj1tIhaysMl1Ag/Qo3FtMsGfmeTXvboi2rhOrhy3at7yn3aN6GihHS
DqbS9F9EogwtIoi/66nCQHk2syLmLjxN+vVNBvyp3eypL2b7BR4uCupIt+6Poty0
Xd2FxJyC0CiZID/LDzXaA0Go10wunaIx5uonXyJ768sIDM7UBCLTc8yUTgl4ASpb
UgUkDK+qdl437RBUXXvsrK92R3/j2ErRXu966mqwqRmSwJmNobPU1ITce0LGPbiK
DMf2w5vdF/DsHdYCiT94IZO0IkNO/7jqqw8Saxv1N7V9nXAhZS81RqzuCars+t5Z
osuF6Qtrh4cl7fFQMsxIHSSeBeVQla8ALgRaXZ15HaemuCslVsgB1/fzLkbuOAqw
ggSOcFTtiYGsZUySjfyRSTDBE+ZEpC/p/yYgGIXVNes/nOlosO3TYUiXu/Gqy052
rFUTX9OVy8ofjPw8WhXvdFdhaiHORyd7HBAq189285lUNGId/SFTz9mQ29w1dFKP
WMrEWND0o4CMoKIS3kPcp5ZU/3KpRHjNL3vhkC3AlFk6JZXVNIyMv9XFe8xNTi8U
gClSgEMfXaiGWLhgGIvUKnkPez/qQJFDQHX/GJlDePpvtWss3WVpITKxu1swrANz
bnoWurXD7McllCyX4By9jfK9S1JZfehDIBnjsXyLf8HsYf8QXFYmGF37F0PpoA7V
NdmvcbXctD1ZiflpcjDIEg+XnwjUPBV98NM9kosy1F790errtZJdxjeqaNfI7jOp
WXZzppYUfVfK+uEzPbyVYZJwQeE5/hN09f0Cpvro2tkiMAFTLZqtUdUmyFyfJfdw
qSoThvmA3E5xd/nMYEiEcT5VA1xFxXEoHVRmdXTvcZ9H/dkd0w0QaAIT7Met+Fj+
bTiDRuv1BNp9nNuWqQDe2fESwYd8KUei/SNH9QMhV9nECH/+NeQiRZ3l6t38RcPV
Z+9HCJsYc2k074GFHS+AO025m0CbQgROIYfpwgv52AlLBbeczqLXyDCnJVofhLc8
RoeyBfxXg0Q5VfzjXkDalQvaASFMwLxnCp6x5zYTU7hPtu6s79yQy9iuYmM83k/k
hb6FiNomZvmELD+cu4i/sxrgCCTu3oSFY1n/DfOw36LTbPahq33J63o2BYhhxUBy
dSlblegC6Uvnjd/d3bC2xsf185ST8fkUZCNycgwwZvWQL2HORBVwUtxeGk38Hmlb
esaYRpFOIXqE+X9MNdX6g3onu/qiNMYamE+tE5BCVKddWi4WbxLQMV8oxUQT6zwy
VrAL/qwSmn1smo3qvM9IMotfTnWd28FMg4HSrFjPCswjWIUqSkZetIW1aDEdNWzq
v5c8X7Y0pKBca0iD1ob83nREihcfsu9H1Yv9qFczGVHH4HTVoNWgVXYDEClfLlyJ
hyrs5sB/kdPrynemqRORZfHXYED8WgBhBgWoQRRaHheZrdsTRJnJdB7WRyZ7QaoA
CY67yvwcPAuEFuBCex2bt1NpwSh4cvhDSRh3/jQUpfeNaYEymVDyQv21B6e8FMCM
/0JznXq3mUiKP/6WihD/kIFBLNhjJE50D2c2zF9g4XrKxKCUS6PIpgEPWR6gtzKJ
rHLjJlmlNgo32rpmLIXPi/165mM0cBo2hIh2WyJHq5QI4NBP2WF+jNVxmksk5z4q
n1Fu81IDEY9te7jWNzNdgg3bNtf1iFsunxow3B7IfHYkDlzXb11MEXhMXgemhGvw
rLzcVC9KyRUvi0bF9JVE1XbpSezPX0Y+NEdsNUfRACTS8lxVi7IakfO6bfxCOG8i
BClnEEIZnjRayPpUrMf1nC4LiTPTM725t0OwHc4kbh85W/yS54dhB7r6KnpJn1G0
CRfowcejOH1raXjDVBUf+85iVY0O0xKt6PU8KHGwXbN8hNUz01THoO/aUu4Ln3qx
zRh+0LlnUk9pEy162cGD+rPZWvlj8jrNBCkqug318GsFn565kOH04fMAkUyWJ1KM
piYICD26z3BtWnK1Zb2bSDjQCSzzyK+7v9diBBx5QCPbDuLIMQvr2YHEexhjn9UQ
1Rcs/tbXd/nhyv2873THqzf5gEMG7mLpsK7+Q2pdAJOJ/cqE+HshCIvqs2gpI/Qa
nxQQhJgvzfbQPHMYdVeFbO9JwplICQ7/dkQ9AbhfHb9HyTbK6/CjuxAB5ROT9BGH
zcAEyT5Ww3HJU5KNZ+F1dEOgPaIRL/qellvmOUZSgZy85j7gS1BGAiGTPAm4iE6F
oEHGMMMl7KTzrOUMryWi1wCSgalrd3UBWFm1XbMDDO1yfMFAoJ/3CMLP534y1Q+q
7OUtrfiNu6QO+SGySC3t4gVZbtGquIa4VhfZiHv+4CDj/rO7k7lblfTatMlXW8WB
wEnjWDlJzduHXfdkvkFxkoj6OJWa01q+02LM2j+bI1bATMRYhN0o9xrop9RAowOU
uJM3FYFZx9192jGFcazpKN+zlXGdGrUCpDpGUYFbtV60W0UdyaGMJFD5z3KWlBz1
vQ295XJXX7wTXyJfpRK3/wfiK86qcqkvatqB0KKuCAI9reOu2ab5vYYy1uHmHMyR
iIr1+rPkfSRYltEKSPwbY6Dh8YcPhMz19XNsCB+QVF+U8TmDuYnwS/8V2XSSgFnN
xWxRwzRTyiwZANnrnH9OMVWnGKanjNKmRHQdjoj/rbriHMDZx9K4Xn6tgUScg5eq
pNIxM0644vQHD89ljPCxwUh4KMthAz6ctgLrk5hdo+CNDq+O6FOZ1/Sbr2s1wMgx
V+Q7yLu/TqRII4HrahWjEoa41Lx1sBCiL2PEMYUji9te7g0/ZbBY6whBzPofp7P+
K7MiasZdkaGc1fKqkaZ0BLH88gsfWCBn2/u7XfSw5Eq3xlwXnjmslieA8qi1ZSpq
FWfk0D0BODVXAJjcFDpw4TS2XKPuDIS9qgBWk+/4fuCjFM6M4PjaLG+Fe+SRlx+3
Mgl5denD127m1xSSib5eU9TIrxpDyNgajPO7MnAz3HepydA9OcPHZjq43INlAmkW
UlUf/oe0PcSWprSXqhOGmlZs/Mwca/BhLhDmOwZMZS3s14r4YzaBZgZbJcOUJkzf
IqVvIxzh3bBxdMyXcoYQH3tQoJHFdyzM7AmTUPcvsTCpBrRKlKbVXGu9xghTXdDm
r/UtX/cxgsqWLhxpbcnHYNizLvziclZTODJPCroqORu8b/at8+sULKzIJycAp6w7
ZLMTGe/sgvgYUnw3VMoDiYULZWAAjlcFY02HJkVc5Ins2V0XrrYrRNwiJ/Knwgzr
Ss+itl0mBo+8gjkoZCdzs+OSN2+4HD+bKtrPvYRmbgLW8tobh0XPkT+3AdAE5UnC
5Dbw4751J67deUU22MO+1CZ88Pns2I693Cue0AJBvmzRwJxNYOoGWTyl0DAZ/wP/
42KRx5I9YZZLWKNzU9htf0/U2aeAt7jaVyQXtty0xjLNoHxTB6y10Nf1XXrl+Kbq
4FQ9PmtaUDr5PXPe3CR6m4b1l5KJURiEEFJSYxqmVEPKiN286rQJTp/Xv6W4EW1L
Jv3J+Cw1LP6EoN89deJOsNFrVaHTnUjEpz8BrPng4FUnYagrL7q1RVo2tOCT4R47
YbJItpOJaqz/B5BPvc1Bkv24bJvB0wg0gEsryO0nNX7rEO07iatiuY3I0JOgSXkl
OkdGRopOQ1wZFXu+vTy5bTE9gvtRpsGY2KXOtA2LU28i8sJPuNgR06HCd/ro2P6y
KxdHQ8Q8i2XJSjXHS57pepQJ+zKfcsYFlEYSHvjGr/+aICLvFnbu79NH9uoovjRJ
OO3JzloNQeJw3xq+NpNGOC7zekTUMQBg2x4xWphIHD6CflFFRO8w/uA9U5rcsS5Q
tFDvb/tuTjqXiZnDt9fpfx1ZyDY2LmuunGCa2lbhhCEeNRc+ASrmIVlas3LazHLU
9MvjIhWhmAykMeVoex3+CccQkdjT9yLTDs8Pf+eFNJ9PJetUw7aEWPSeTVVVOUIr
LNxZmkumnvagC0CWS4aHoupQ1pRZcwOqjgrATACmwg/Vn2mkyCDqmlLz2V6dmeMn
350Jd8lX/bymoq32mGIHGvEx1R7XNyiGbuJgg0nVgzqYy82CstV8QoxdUUHli4RB
5aexutKPcU8cps7OJnk0Z82FojkldSxzQnwdt+h8WJHRyEBk5TqwhR4We6hdGXPn
RgH+sLPrEgCMRfUz4o/4GQwWPSaWAQ5VxbFiMD2F3CpYZ2PeqbbAc7lOdThXoF78
uhsTLR+0R8D8sr8RA2RgL+bOXhw824+Xdjb70cYVK27m9IzOpJfj8G9OCiHMfnoJ
Q8SObBx3DcqvGzoh2yg4uKE7jDfgrU2jsyQIaUDlzGUPJNR+wIvK5SGpKoFySuTD
8i2CxItrSpXnB1qZKMni/JeOjfiRcrxcEV39ahGBfsJJIijXAF4rzzH0u6sEDOuh
GX5ViceAFEvcIE9gQtS7oes48K0uHJkUXM83vULdf+SFK9WcsDyCwjkrpV00POC8
C+XLp/BWsOsGSTs0RFAZm1hn/8ePvEdIelYupNvYLJ8AG/myVrmgeF4qdiE/ub3L
d1lr7vJEHZZzmYbtoGsoyEecIqc7vcNEjaZUKr3b8PlFZJLftlBlqr8ol7CqoHAB
rdDnLiMN1+DcjNhztTsdW5lDBs8rdQjmf+66Jbe/UwrPwwCcgt8U7ESxNVULYG6J
gSm27vj0tBnkLNJb4VubQOkf/i7VtzkU/8AfJPKbZ0P3GbEIZFV60P5ZzOZ1+G8C
czEkH5udzardxV4r9Kca1nYkChnMd2952vICfIdGghYX8mizZkU9K9AlvMClpHJ6
89F+5b8/jCK7evCgsAAE3DPfL5E/WTWFt41y8/Z0jOmOiS21s45XbLMl9cnipnWj
bekDg9LKXFUCaRl87LLzh0fyhBDopJvsMrfz4VP1MFOkTYvn4RkEyvB1gicC16RW
0po7RN8FGz7H21aS0HnZ87GLJInt1Iskv9ieKTjZC80ebDOeuLo1Ww0hfv8q5Zes
tibaBwuOAjaLsK03h9lyQR3mb0b1DsfER7wpIkcBkKmDbHvCtp44WtbBBGl/AkKJ
9x+t3+R1OMfAOoGCcDM63FsbO564rpAYTxURU7oaFLlTSsUZhJWLSNYL4kHb+IEv
BiIa0tHUf9zwpdfNCD/lgLKIk2PilWyQUPrt8d+NJJSznKWLUiSnKsnKUZADI5df
8kfbeHg1uJY9YDDjKeNQVdHIlxqTCe0BBj1O7ElbJmuImp/sc7SAMlAv/L9RLlXp
vR2yvvhDKDok7nkmGtVZl0l8oGUsvX7YT2y3jKgJR368EubNn8OTwqTfGedb+Lxo
tPdf7abN6T2opd7z7pfNOu+LMre2ASz9ln6NpG6Nd3W1j05MhXO+EuzcAKTybAg3
u/nPDAO747btpLCIWtKzTnkBKXlV18PQsTQI/ccOTidJjBbnUVboyj8AMwXf6XZ9
iGs4APWdJpsuFI2X/sC4+c8EhBkzim8u4UWfL7hq/rnLpBZxeWx4mqFi4Bv7t3Nw
+s+Y45NnvPaq7Sv/atw9pikQUhh+yciPrRj8Qqbmzlb5gOk4S6/EacdOwFJ5POxy
9YtWnQzyMzZ858q9+bsm2WG81Aqf8vqNvisoUm/f9fwfr+AFZW5E0EFoIoUcd/gg
Ebtgmtwmzk5y7Pqun849DqR1Q9TXvV8KCeEZcjsQDYfQTSWd/dgW13HBGWorkuov
V3HA+49dQuSciUbB0ZVZ7BjAIXI2cwImIWe378Qai+wdPbzP5BxB0KYjB8IxhWzj
iB1K6R7O+/dd0bKOTt3AmXzMqMmvx7r7+KkzygCzU9s5K05QCG0BdvGC66TZBAQ1
S5qLYcYVOqi2ndZ0nKexkqVMHrilbC1PKlIQG5wuDbJ+jvFO72ohf8hc0evva0Q3
HfVzMLofv9eppweJqHi4h6IJ5SMlSmPlDERW17oMIdcX48UFRJfQ9nkzvNkjIPjU
B5ILCZo/aRGDzPhniRemV5FYwHquhLcg6Ke+VkWjeDjfETzWKKB91MIu9CIHRbQT
P9u2cr+hzUFbHFeDvF5aosPUwOvDFQYBYjMP3ZgYrFP3ljpFN+awPasU19E54XLe
1v8r1rSDZpN7jCdsCeGEDp4iFBZWpw6fFYF5ZUoPN+9Vkv9LxLea+NOiJxjuUM13
TwymcsHLLZU9rbioyN8+6K8GwtArcqMM0pkh8RCe8yDggCw903KYA/heJHy7UUhl
sUjVp4bHMAywNLGnrApfYf0drg+TmHKFRSQVM2306W5V/qqLq4SA0KS6pvU9sa2e
+WkG6SLk0mQETLiusQyZzNvmgDKVz6mn8sRLFx8ieEoBt+JIBYhVC5ahfX+U60Fh
1sRDYJ/h5QPq7zqL6k4TWVbgmr7YyAVZHIbVv6QRbAw58vm1GAy1+0nCB2qkav7W
m6F7iGwUrCMMvvcxCgOQO5W+/nXjVOx8CbVq81ARWgeqZyoKT2BAllMB9lDaN4pv
1Zz2mUyrCa8vKwjiAVmNT74AUJKwdYN1Cpsm77LttceIH/SCMna5hyd+8ZHT/blm
tBuKefuHKaSDRSxGraaolgS9jkxOKDGa8KAVbEH4oxns6PgjTO/YJ1NSf5EJUcGd
NHRw8msRVh73UEnc36K4Xxer54F7PuiJBulth13sh8WO0/JHBCO6MdnblP52GnyV
Qn5RWbPKH6Qo6MTXLFd0FFqJ90XbkBA/zl5PAQM5qy582IQK4DybRJmvlbI5HIQj
x/289wZRZ9E0OQ2FjJF6C6vr12BpYxp9EhRFEtMSwP4ng6R1D+mHGsEcb6OFZQuh
3FHITOanNzyLC27UdiAH/EiDlCaQHY3itstQL6OxAcbNBNMQnVgcgd95KgKQhQ1d
vWEQm11bfeBnNS+LQqzOC3mY5bA2fnLUhgAkR8b99/lw42FtWPH+mLtHgvzILL1w
zHBulcjjXsC57iN+bwBxC3TrVSNH7TwX8IvBhXPx2vQYtYc//VwqqMDFzm41Ib4H
X/7fPyl3BO56xuVcLOE49IYGzfYxkdU0h7QQ3zpVs7fHFO4HkFFNtF0yUoP3TKaY
cFI6RzM0BCqX9gpajEutPK0+dKnDo8u4n0nrRlkEEdMXPseUsw6Rz+Vmo9nX/fYh
ueh9SLwHRpN9Wmw8k6AZk4uxYFbWZcL0pi5L0sPLsYnDWKulmfh1flteC3Wcu3X0
P9E4SoJC9LImhClfa1T+w4cIq9WqOvzD99bFwdOSdSbWXs5bebOkhG2aXFn0MXt/
tXRVmebUjKzPoyaN8gcpMfNKEeDM4Zhq45Yjt7nth3rVXs1XH6ANmcRRDWC9AMQF
DdQ7wS8ffAyr0nJVUbs0yfCSxfzrUq25q0zjYwPDUA2DSkW69Lhojz2WE9LQ1G98
hUsrZRgq1Wg/BiXTgqYE0NHrECdjWqeip4LBCnm37ABoSCq9wDyd1pARRqO/iT4N
0r/MJwt4rbO5A6qIwV8AvffvasyIWzY2hmKUUCqrHM7zankJgGadNKCkO9TKHba/
7FGnAJYrhTbCKdg7T8Peig5b4QVaa8FiejfnhgGosbTxJQx5ia2mOQQZj/Hd4wla
3ZaVAPCQBMgiDrWupIOc5DobDbue4LekE+IObhrNc8eSnm7PTrnVF2AXaRIwldhT
SF7F/JINfrPi5v+lAAD5Pn959nQ3wuzuWRMkP4TBczXa4ZLID+E4MAnlIiwBj7PJ
pvfncOCCEuqKqj5wlpQn1zjzdrgkjUeXRyX6SLMhuJI/InXsYyF0YBfo/kYxNyT6
TdSYlWiHM97cSmniN6BI1cV67lIbPSKWS1APbeGAYYjSx4G2uZ+6zUwqp7ge/cYv
zbRRze1quPQDOGbC9tDVf7Lb3d6gJ/l1V0ELZz3CQdCmh5HCsef4CtYrx4NN6cRJ
OXQt5nQEuXidz7qDzfjap1fS9QDn1p1O540drhi7h9uWP+LQlqnb52rtXdZUXyeA
FbVRc7s6JZW/RgG2+7MrEuUGF/DMvRf9wVIro1PbeUbu794IWxTTqqxbX6dwPvpX
gz2dYf6LK1nlbfI6K2qmA9TVdQjfCjsveq9GnKUX+5SsrzOwLlBksmuXGgurTnt4
5lZJ9hkaZKe9ahnwbKasBXxID/aGK6RCCoSDQsmT4uIH0g3o8oTtLTfxRBq4rYWU
CNcYUmW1sDhEDALQu+bTn8Ly4upVHi8ky9skAc1nlXfy06Gp+xGAFHTiHSkNG3+/
txSLxSYUjJt/Z2LXWLAhROLIy++uJXGstQxaRMYSLpgbXmtzO97AKJ2IsfAwuZH1
cwOjUhdz7iUXtgDFYK1OHK+yuztQfH7zTwT32U0WFgXYUL3KmAlTMlH0IcXT224t
qn3QReZ/0XWkZ69YO8eeY1FwEoRyK2xtym0idt/2w/4GadvQ9QVP+fZY3YusHFcA
mIofR9eMpmU/CHETCN29LrTEDnSp+udi2tITcUx7qeCXbvgpbTGt9q7kamtaJLrY
+ewbpyV//6jxq1jnZM0JLLiDMGgbhh7bmWeS99OO3SPXyOrfhSe+arbbpT5N872J
0B/ETwNYBeMMoPuH2bAyxPEuFLxnin+vQ6+W+uBIBDutp6UxsusKAeP1gB1nImim
MaPkcbz07XHSDf+MUZ6WlkBpZeyvw2NJVA1dcgYjGY9pLjubPcK+IcqiuVgMeIZg
Hqqh+r61BLlbWX1mabEkgA77KkjCT4wylCaAGCx1lse/BT6wstkzaZYl9VA1475j
ooIssEIKUx78P1I4XTT6DDnNCtCYVDSpsfwUpGoYun73OEy1XXKv+hLZ3OPhRoXJ
KSXmg3c5MLQOjYhRWlHS6IE2d3XIcaojYo4raWw0Zxmt2kh3iBVAiCNQfDQkwVzc
8WQsVx0Bntqq/tZ5b2Q+uT5KjfvU+6QRT8htONbxa7vzxjxUAXgQPCe+ocl6OXef
vSggIbCaOVLbICavx4DAp4QzzwXErAPQiEjB6f2iSPbqSjv0LwtToYNQ06c6tgCx
8tLfcUa7GpxOL990KRidRHoYaSFEsmKE7vsSTwSPiX+ixxdmy3siqE0ZWfcpJThy
6jqauQOeWlHfLjKLG6xdrTLsP+8R/T0zE3LVHCHhduyedKkc6Fm5iviRz41Ke9es
TrbkNvqKdqXCk6pu4F+6MtFbPvC4PEvsy5CYGSjjlBmCKVZc0TaxWmXKvfcjdQ6y
P8SsTGrPa7HW2+yXZT+QISdHuePlw3Nojn/zjAzZB/QTHysecTrM/CZ3AO+5JiRM
nbsn04y95ZujQnXaoLFJOfe/UdbNjj41t/4jnvNpkA3M8LsaA87LqNpCtJWAilxa
Vi6+Lg/QQi7GgFfS9ZczP3dtCIqQyhCD11lVRlXHm+6tYu0HWuNQ7BrTkJmPK9hq
7DC8huMKPcwDnE22Vm9FUUCIemYHHbDQqoRQf0IojW5JSuE9FDzY93jXDjV+RLba
5q0gUM8L4PeBNNXPOGjeb8ZKFfwzWDFXmKpl1+oFFxOEUw1RrTvQzSFuyJq7G5Lr
lkDWZHB/XRxzIypypPuzAg/bGxDG8+lvICKJkTPyeF1QgtCN7r/eUqefdQSkLuhf
RQy0Sn3OnR8nTLRUg0mphfkK9DJOcB87Qayx76K65ohbHv06B9rRsOv/ppzwaXF4
Aj2vFj2Lmom6XjWJ1EMfWPTPciRoa9iqZEnmknz4pMkviUmyYH5OWHfQSV4gnNgK
qqq8aIchtbUoXH9C87G7BxWS2FrIsIU8R7NgqzE132SRmEINTniEiA7zea+fmIIw
/J8jZQRNHYNqw3rFulilox9L8NEfZ6bQwJhOQ3upbfX1zQUsuQbbB0naIHIiC6Ee
qxqU7oCEbmeKKa4tMt4hTn+k1d4LTTk0BW8VP9h1bxQao71t/94Isuuo0WqfKmV3
1d+FM8GUMu6GFnJarqrDteFbyabRbmoNm0XGyoC0TLBRH7ELiLUszSVwTVatVF2g
L9q5e5+6mOMBihHBXhDjgTD8WA9c/OjZdQ3W0PSej/nRJEcqjZFQUYfhdQKT3mB7
l1dVevPl5eGeVyGFXHP1Vle+3xIHFuCW/MDT457TgF+ZcmcNYnBtXjbwwj5fJcQe
Tsnjrm4F8A+BrOMslqmWHOhUnW5w1e89rsEp14Quf8cd01Rw7bKcKZ9PTEFgiC9o
sG7gZKSHuFFN/IBBPe+uxEVszmoxqNCpVzRfXjhE6a737hz18YFhspfyKl+R+kAT
Xb8Vd5fsl5VavRejQjH2osDzbYeYb8+MZ6OqlXVjTboBKVrLceBH56/Ksm+zS/HT
obRvMGUTit1Dj7jKSJI1rKglvJaSID1wBPPg+WPH8LB1QQjyYoLjjbhDR34R+hrq
SHGnKkI0LHq4OQnJjFUOCRBilVT2+0EEsNd5zQy2suPwBDs8qKbzR+jExuFaHy2K
aduDK1GFcb059hh4lLL8/wqZuLlrTCVL7QVBrcVXiBm5/V+3GIIPUuY9iqZUAQI/
SAW42TlVEiH3LX+kqAO8b2AeHpGJow/Z12EV3W04g2Cfim2h7jZqwmotAHn9rz+F
IxiE1qjhPrKIaAifDwmbPgpNdaxy6jql17HCX9kwfnkjk1IHZT8/755B+SWHW+1k
bugw9Z2qdkw65SxN6duW+6THhvP0KS7gHkpO0P/NK/H6aFvDJqMFChextOnS8Wb1
+CHwh+Muuc4CaPixjewpbBW0id/+taoVWZr81qbEOyXu4aDDCrI5MtZKXUp7Lb9d
XrOTbHZzBcbjAnpGXlwOmHZ9UdD5uhgXkXxYWzRuXY+FVbe5e4geqQDNqjUzGZDY
04ljWn6LscXJ4BhbDJjY06OudUFNJoK+Tm10mf4yJGO0hQi9DfPMfKuPiM+ddDu5
4uI6/1+DWkduny/9i0G5kXmm8UAHvTO3vOyHnMEXrcVzU/za788V+hNCDeb7qxv3
agp9INiv/zDxHBYESSp4NX28AKE1dcpS7GDIy4dK4RpAC2DxhVycYRfxXCKRn7TX
deNel9j2+i7RkS0SthfiPR0PpFeaiDhR65I8fNpGXBeec86DxD+7kzmkdSBuNFRG
xl3SpnYubvb+/w4zbEa/lm9gwcfs1z+IxBd421IvFXhtK4HkrrnovsWOvDXZFymj
SuvK17Z5bBtSdwutLHn9VPm1+1qypn/jh2X8/VX60Wbu72S5zfnKDlsh+pcWBHVp
8rV/LFdc6Uyb9Xv+olnXNe9ae6kJoyossKfe6f+MyAzKXnVp2P1vCDF6RSfmVgi6
oQSLJKwlr/sCmkvCKCDGlFbg4/fNunsFbDPA9f2v6pr3R2nmtc3NU4i/O9SKD7Gp
euxDsz/EENajMKrh8T9Nsr+SmfeJ5y/+KfIYMAjyB9LN4UK20ixzGK+uhtEnWtVU
a2r+JwScMziKf2M0ru8jHoJSParDQKm+KK9SvaYc3wI3KLZzsPY9EF46DjIuTJHf
S2LY42/QNO3DYbSR3o6+ugH1QyrrZuKD9mkN1k3FF8qhr0Vh1Mzps6fLpZc8JHIM
vTO4Wu37ScgY335a5EpSVnWM1ULBL/0lTvt9WoeedhFq+d9OLdt9eK+32T9Q1sNf
VyviVu2Pcy7LPgarrPmdTz6ljvrowvSVl+kkefSCsFovhc7kVfHCDgq/sVhQ2UkC
tPbTxZAXDeHRBeDDBOlH4ZIbvdgKtWOhQupKSMnb25+2OU5V7T/gt8sj2tpVC/Wr
jwPytsZL8op7GUJ8CsCqNB1Uey4wgjn9srn7icr5EFJ8MOexZfffC3bLygVhIAUN
6V45oVSCTCkpzvv9XRGkPIPopmdDmcR1nv+xjanMQTEF9J523Wla/qGi6Gc/sI0g
8bA2BaittVHlpP+3QffgJe5Nj2UVU1H3H+GFZx7VdC1S/BQr+PKZx8rpO1GMRZVQ
2L6VKHLjedQstIgrj3zhw4RqWXKryQAw8k6fXONfMXw3qunlGUMIzarqrXOZp5ZV
gJj2gp7u8mILTII9e7pUysXtkvBCVX3dO0Koy2Kn7+UvVYG8KWY05YjwHFHtf2qV
prhX1mqze0hNNuG52XtI0q8IbQNvY8p78TBSYV0RLvy46YtjAM3lf487yDD94vo+
FSxoFl5NjOhm6fEkX0HriugY4o50rDfp6M5YxfOHT7rt19vgQXaj/lD5DYeWLr1W
PaljL28awPzBcGfvw/3eYZg0c4d3fwwPtlD+0SfIaGQ+QvmRGViN13sKEcHxKLdj
o138VnHq5nKLnwx83AF9Y01H5FNhtjZOCtdUFO3KX5+Rdr/u5hi/TpT/OyF5irHL
nlDc/Vgr7PGfHUPdopuOYesWr0V0gQ1NKHU/8bYeme5ihKLKSmolFlPHci7Eyklm
DPbvyXCv6hmyNOiplYoP9WeCfKyNVeyrlr616GSUx5FlKFouIe2CiLi91fbnS2rX
L3CLCNGp8hA1C0bw2aLnn1RTFHRFlryqh6tBzqbE5P9Cbd1/KxIdGhtzR6J8aHi7
YdmGLzoDfD7wJzeQO1U+6CInKV4IcsXCFidl/QsLjWoEr2oeMv6cMnvHjKT0DJjQ
lRAXbDz0+Y5Vd+Xn6xQjZPtvPGQyk/aybUk0s8o+iUsnJqBzS1xrzSp7hzCYkaV7
t1lnfojwvOIVG3yASKUtt0EVULcCu7cEK0LM100l9hDHgtcgGQKd6XH2MRyBHveQ
y/Fjdx5vw6O0VsSjqujJ/bhHvQe5V33eNM2fxGjCZ0rlmUNms6i/l9sjRA4eKLrB
eJ6fSDUIFJ3p5xlG62ltSuGdXT731REA2fk+aBiMkTTT80l3cP0o+al0/3SlEl+A
g5UhW24lLTw2TVZ0SrjJsTIBAkuZ3TPIPV08qW5kWEBIkOcOf4sbc1+4ZdvFFHBe
zHXCDcB3r2sRUmHyHUaqWtt8ZAYycGzTgxOpuU7LLQFnGGNSoJb6w2Vo9WHJSNZn
J4X09iwnrC0VO7nTvB5w8ISKzjjqDHIhsCF5z50/fpY3kZBA8jBG2Inij/TbBOgc
4DE9Jj8P5L+Grf3Wkce0JLR7yfq3BtjMN1LhEh2OFiIDl0SvtpaLuiuF8emfs4CD
O0HLu1atWFx2AcTN0BC96YfF8kTmle4RgWMQSnF6CxpNn8wVKIG52bAjbwIkJiBT
owmYQrcsZt3+x7YPUcTF17LSzTu3gEAbu1iB6qT9Chq8wQ80fXfwkNsJWeYCcGOL
u/LJ0rTBIXV89wXFeyShOPKiXj8L+/2Q70BUixQKsn6jydKxEDY/j3oevHFhJYVt
ew2mJ47tjG3TpfBgY6AV5gz3a+xcIWxiXKrea+fK1lQy0+WeTUn4/nLcu0OOykb8
xQ2udFNwigPX80SJZ1q2HP0xXgWnwZV7wkeXl0+2mxbvUuUYoD8pLN8Q9weAgHI3
KPkRBlHVo1fU12GUrBsGN7S7BZPaOqdG5VDClV9QrJWD+IZ/oFYTLH6+yJF+EBSG
eHLZ+lj/O3AVs792IzQhKKIEeMe8W7RjJI/hFAM6VEAthWtt4hyHctCLKlpzC+c9
BdnJII0tA3ejTY1X6fts9u4ulS+pIkVaYnW4CaYSpEwN2UzQlXvsMPd39qwkFLyP
QWYsEhxfQ3XnBNmzXfvVXXDVQZfbA2Z9hwH6Tku+VbNS4SjLcMzdgcuE8xS8+/K1
E9LPIEk2Casn5RbWRQKkshL2kHGqVTe384XZGlm4sOSUp6te6Tmgy3OtoQt0Tc6l
+LadsV4dgU/aeL3fnXUIFGg2xVk6ssAT5uKifu8trUGTsvI6qkjUiP/+4+YTkigD
YrxcLOd8nTDFjR4wPUkB0cUj3dqb4QldzApHNQHtdC03lLjCMFGgwDpMcKvE+nDs
VqKhC71MmAkdWyJok5Z1EmwpbKRl/a07fsqIDSVHh1zdJ0dUoLVRPakZ4HhnuSJS
eqZe3zNVIA7C1vXpxGgyRdDxp0g35UJrmaqB8cqcGhgG6lNwvk7hheCnK6ileQ50
aeCVmly1NekSMG5WkOW+Lp7CD8+tvIJl84nP7GNdhlRez4BFElVhiKDBwi4UGc9v
6RB7P1rHFRBR80me5DF93TcFv+O12HFxPy59uFwM/XxR4fVmwbghnACKKR/P+Uo9
dXzmBIK8HqyWCfbbldINHlY8mV3ldennY5HWa8BcJiMKts/sFUvRFECn7A6GTMiY
EY+inD6H+h1b67PdlFDb8H/+9Yv6OSGlb6T/Z7WU4dTR71f8autXJDaYhCuj9k3U
9avb0a+m7nzhdTNeE/n/4AvPCn6GpKUg6vcGKnlwLDzIE4nqPzjPt9jyEsVFXDOW
IyL6e/Z9rs6zZzorgTR/6SpdMM0XAF5bmY8xF6Mxf8BvTlCpdGEdqb81ao+bywr4
G3ue5TzjBt4cLpRhl4GizlY8SjZcOeUEyL5Zk4SRCwE/zzXP6gU+oE4nL0TLfoVk
KLMrifShUf+KiynIoBRwXCJvvlkgpDwXjpwwHq2NoMijIGk/soOscntL9VKA7M14
U97LuJI5FYY07IUl7/C8ndUDfWIQy8sP+VpoCafOxpbFZsZXKUwqvMKf4cEUTYqE
WLNsngez8FBNHndmre+LUj6+EqKAnOzsB6WLmWz9Y4bvVx8N+cz6PrtVFgEUFZ83
qboCM1O4zgC5G9BTBnPksC9kRIP5aRULPCxYcpDkIa4KxfJD6lNdZk5U2q+64rmM
alq2FbpoI1iqLl4ySJWYxFpIbwHu9T3W3dkQMJLJgMB3MYtGU8yw5//mgGees9KS
URNV0MIK3zJeMvktOSCqFuOa0LvNGs3zX6D3T+al+k21ZtVWaUowaPItSbosDvir
suyl8nrora4WYcXTdJCJJlrUbyZS5s4HES85LVtbQJSr1bAuIindqsKtePGbzGEG
UypYXbc2uJpnMLMCrpUiGSyZLyEiYDe5ziNGXVPtuAzp+gk0uWz+GdzQdQqnMcGR
LsgdPUZj3NbueKY/yInJiDbXIxWhzKz7zKFtCf+8VfIfZLZ+fCyPJSugKx6xqc9F
zdlY/P1xDhJz1R4SAFC1iPeocGdjwx6p9ykKf91bTF+FgVk19nE9hHM9vPXaakAG
HITMUGWY5CJycoBwV1AYIbN66rYnBJGSJchrvSkd9tFQYUI4b/pKpC+MTKJnIITW
PZoTA8uDlYIvr0C+iNM1JZBigPHalnnIKw6JaiJnmTzU8KDXcw22AqQldi21QTZr
O+X1Tqt4TOJdFAFPpJ6Z50/70EtrdX4g+/65gk0SEsTcGD/V1s0mo8fGseyoC7ph
qdQzX5U8NbX7vAfu4dKDq2Rv4nVN792uF3ONOFn9r8V0iTMBD3yPtBGrlUT1dBBm
gQf5y1ZP1fuV9EGJk0coC9J/MYsC6nsP6NsFazjmgSBVOE4ucJu7/wtc5LU8mZEr
pOBp0Se3kz6HFKQsxXpC7MmoHP0hxWH5x/G2NopnIyb3x7Segz2R1AModGfUwYpm
PsdnjV2obgvtpwF0YN0Fza7UVk+fqpF7BMM6qEPbkC55wA9A+SBWzOhzaCckRjBX
bFTQsh/p1FwQ+g8eUMVTT7zndlAcwNMXEm4QQCc1t6KeeCL/7oOMNTcww4fYOIG0
18AoQdg1W3p/rUmc+Qb8SzU2ok70KqHYbpY6W4hP5BYCHu7JWIMQ4dhpYjAfmRCH
Hp69gAdHQ+PGEwxRFFE+9k4GQBFcsfcMwQDRjYMzdfF/ZHw1WE+2WH/rXgb7IcYQ
ZmO8yOlJfN2jaWkZXRlg+ZDHlz7ZC1PxqLni9AiUbnjTRMWfGy+zNpMJbrcMBmoW
Ak8KucBEzKpjWtjTbEH57159UlAf70JboV8tz8bvNFcNv0amzVeXltG7cpdHpdy/
BtEbLEOsn03DCNtH2F9Tri+uPuiQc9nfP4207I4CbNbA8EO43o7F21Mi1bvHJ4k2
1hTYEblPi8gRQguw2ZV7bFQK7AqHRvkUWJgulM+hHHArShQwVf2/LKjJL1/CQfZe
Xwdb05ruGsO+IEJqkrN/Cw9LWzDUFVMPQN7q6MHp1yqD9vZxkEp0cHnwJDJTW+sD
Ubrh/LOTWidaRjh5TkDeFRJFB9Odnrs7/WN6HlVU0XAfky0fIQalZWj9x1gIvjHc
Btvq0pKsyo32ajUXJe9bfGmvozeG78KIMvCpvWdN1nX5WBgxjOBMiPiN8m8LKCoq
7T75mScZTxBSe34fCKYLoAqUnPhZhK0ltWuxmtmtnyZfHYxda3wryMkYhoSY5Phg
x3WzoD//sPM7VwHlNYTZ7XDgn/gEQr5IHMD2JTWdA8XJ6oZ143H7UYjBbkRlG0yp
qSnuPz3Uf41/CtNrD+hVXykDxpTaHUw5NPxQnGesrFDpTb1qAlNIvFoZkNfY/n9+
1fEKYNtRdkANIFSR8fP9rprq7LFY8u9C6WDwHsYsWG5QEUejbmW65nPcFQ4F3Bgr
1scIvpcu/hZetjqCRwIpT3/cNfLo744j1SttBP+PV6VJrEqDEW6UQb6gsZt3w6c+
HrFb1oNCbWC5Y1+kfw1TAA2DFgQj0GN0ohYWke6ZdTnHtg5G/Mh2yuf2tR1xiU9V
bAOCyqm7clpqmchZJidNi+vOAgF525ans5dAK3Vmkp0N6Gsk89Fgn8B/trTDMGRv
EkVSDCN2abZ6skQ91V6AVGUYJpSNqmpv2H8J011F88xZHU/4iQz5RZdT3xBpf4+N
y00rYwgFYPz5GWCWbF1r/L8dOrjWP/HndJAl4IPdSy6Olj9CfrOm5Zj0A8WmDybn
w2HH+gWpfkU6Yb73Xzo5lj8SHZjQurWaCmYGB1vAOh5FYf5XxtliaveFAVQzbpHn
VbsskmFfopMWSXWm0aIkV832cQ6fU3XxVHVHhugFSGsrzEcV4rZzLLT8dLNVHmfO
dPMU3VTP9x2rHZ6EiSLY6giMQAXYFp2SFud756V9sYzM6/9BQM/hANDsoFFaLQgJ
6gqJH5ja+bE4/r6d5gDgowm+kjQHWoOidmukVwLy5IBztxodV82kHsTyLRrmJ/kO
R1tEYXnwccaqav2mj1ulsQJ8eDWQDeodNsBTFwC+/8bPzFgo2OAnQ3lY6/7ULX8m
M+X5IcN+QGNyoQviVpx42Z0+yH9ZIpUPJI1eRK+uCZoMfAUtNeG+ya3+l9c5sMwU
qiYi+zUCuv8GMstb7yAID4JYy2/kJRZgGZrr6TwhmZFbhn8iAXBm06p10jQKP5IG
EwRwt2rHCRBbFdm0NHgTaMfhEePoQbLT0HCBAQP6IjqJh37wScXo6LRRC1YjBCtA
iEcOW7RNOtgf2qkYnGfuJ1ajS4YSwWkF+a149miKEse26vGmmLpbmYuomnxE6HL5
l5Z+tt6N5Ibbgcg+Mhj3zR0oYEH2gA/efMehF7mVEbmceSoZQmOXaadL94kwGsxI
fb48GbQek14TEWwhHP8McRdoXfs/FavxaiTryF+JPkdUh8bxfulrBBEMO3Ze6fRD
juj/s0aQ7ljEHZvX0VPi38e6f6xr30dJ0QLnoYhL0aYS6PJzbPjgb8yc897Q3PQq
PKgcz/FTwHAphkjqIXjDZwotqs1nIpKnKwlo7voEnP4gqZSk7b0Q9Vy+rgmIlBML
B38gJFdYTruDxvmSfqhWmYCOr7B3boW/R/ruN2/IMliQHJM950TaOMcAtUt16OTD
gg+CY6QkKx9dzhdJ6aBV1X1XpTxb2sBhgjEmd3s+GSnm+CLEQHSCZ/cL5huN6JVm
NeA/OQdgzMVoaRg6b5pY18g1QFGt9cWkQcsmairfMQAi1+jXfmIPpWGjNDVfAn4t
CpiNV8Gj5HUERjj2Q3Hd1L2hY5WtTCcwXBSKFUD0s2MfNKrP1xxe1Pki4I9emVro
hbr0rxmzJDYOAezbntIH6BICrYFXmm+1l12suSoRMa5ok1nQQ98fUP8dgKrhyN6P
UAuHAZCVW5Bo2w0A63h/dFBXkfnqrNZfS8DAF4HUXzt4u+D8sCsBIyCFPOg7RTOH
kNtb/EglvE+joihuMfYbevH92FJkEy0bWIgUhOnxmPpv4vqdMzMk5Dhx4utsZ+Bw
T6ZzzSqWfGfk9EfSJVrb5nLgkyBzM9idPe+VbNqot8RDF+ANu2CljZejnMRbCWOg
BzIL+fh4tLU30yAKCfx1AtXW7HsUi+UHHyHx43hvEtvp7ciCVzm66jeDnoKPjPGd
J7p7gnEYRyjw3ZcYp8/sCrRPtcSnMY531fQLryQty/AglEwTDd9i+z4AVUuJFJr2
pCioTCejBPYvVAzYcZPHtRwsxICTTR52TQm++Fxzj/z67Af4nYu+uxjm+seOLZs2
LQCAOGOR1+ZEE6CvyFcCRD3xsBT9xg0pN4cUock9hc1pR/576dFSLzs2QNtRFPb/
p/s4du2ZleAz/9rQeSvsgUg0TU9AaGuROVgx0/b2hQnZ3pawr1dGg3wCgWUeY+P2
W1g5RSAie01IMOWKXCWCyQcsB8dGgzocEiRhhNTSvxWWP+G64DqnD2194Q2pgxTi
ju2vxZdyzW7vcm3u/dqFwFJViIa/b9AshaHSdj1CrvLc/s+EwCYDpDCxTUjD7+U7
KNri9WA0hDruqKjC0kGJkt7LePGgp9eq5lbvi42XDxXpDzdxuaJbO5x0041HkK89
qPTPsvD0/a5Sce+bVBcbSVMDFUy/6ykPlWQljrs+iehoft9JkeBmPCwr+AbO3Rvs
1gWGQVMRxIFnwVJJxf1cJxuLmKXie374jGduisstBBX78xQoEnqxQx+VsYEoCDAl
o7EsQKJT9hW88wh6G8IAc3gZMgV+jOn+sglJHQqk3fAjFHjeXuRp0seGVSFFZBA7
0pRloCMrzBKRxBg7uoOrjzFs0YC8ZpSvZ0GTYPRCr87qCx3PrPOGRib2AMsOHIOP
KpV7jmjaMSIix5yqOcmma+L84Ar7qV+3j6bjAMDX4GTOBv9kcAUhR74gICN0Gest
Ww4sZAegmrJnbLle4x84lVzGmCk+uYJ0Yjw4FsS5iGUeMNA4KQ+DeSnYHoPpHWD6
L6Z5kfNHsJ2Gfbl5AAn3z6ksRGi5mbYX36izD8IDA+dJggeCIf+hwkzTm3xPS6kP
vwK/9PltQYxzENsqLlNPP9z+Vh1oBjL+tIb9iKsJkm31BEGHCoGxb1FN6cIGxtH2
l72IcwZRg6NdNrTgRXnHOaU4xYufZnOdzqXtlX5EIymFkNEMDc0IVqtAfGlgJLX7
xe8N5G5LAgICzWxM0dcldJMhrufFfT/8YqqLZyYf3JOmlltYnf3DTv0sylMtzNTV
BC6kuO36g5uDN8SMDmNp6Kp1EYuVN92MRdTbXHCWJOsU+1o2RFzu40l7/t+PUg52
n56ZGqNBkkrHWnISGwwL+hvjBFWsFYWUISgarDR6t3XJ62Ef/j28PUqJKtXX7RPO
09ay5LIaoncJIuzwqdZQ6xHCy98OAPIFMk0IVsVvIr1K1ho4FNiXzsjDkavZtU8g
ojIq3yqnjFhv6FgniLrUHkrArGyGaIzj6+92kx/87HP4O9elv5H/em6plq+N6ov1
NdfK7JHmZft2W7ghODxwAyelLI8FGvLnme8QgkAtD1Jv0hGEWBUJWRTy+x9qKZgL
0CujWkSG8N31b1yZoE823WWiTOvsRzHaQTTZTuKp3lZ+KCGOj6vDezMU5YCe8EB7
ZMAbhVSbZ3rCTCe7MQgl96ETHE17QNeh/SqLIG5C6SvPvqp65msoMxNp2AVuf/F9
da01m+SWb8Hqde8ohBiUiKSEbUO0Y6Sfo4G53M/sGPE3pgmC6kL/yIcugnBsWVa1
vU5NqXRe8tqgttbNrHcTn9rFCrUqhSyCey7fV50loekt5Ya+xFqkacjQKbXWqTj/
eSDaz9+c7gPFVPndF2qWhIsSfX89j84d/ZG5MOZTGVUXNaF21W+nfY9BI4cGsvfg
ibV6R8faez40vIp8U0MR/CbXevawkX0i/XeLx0KvqN6/kcdla6fIuua6SsoXV5e+
AkzjEDtwEgNuMxla4DpKp+WgWTOQZouOi0V2TBnSNBrw8NcwgvWx2axtoJi1PvZJ
op+v+YVnEzk0ajZxhUxOnjeJy6B6ci1bnLEtSC5Qz9SaChqnMmFqhW1fWVpOkwRL
XqSVY7AqGrUX3qZKbA4dZAoJEEBWi3ELu9wqgQ/kJTPfXGoe/9Lre2F481RBZHTH
W+ZFsWWRRznbyVmpNsDroA2kY8rsdk6c/8qFOK4nvRCfuXGR+DU+ehe0e6ET0ZHA
BQmbazRPvCnJk2x1v+v94ISmBJSzlccMkPE4C7OKB6q95PTmPepmMNz4XoQnyv0X
8/vC8oxOUWTD6Sacj7HSfVbsNQfnSCu/+NSYP1I+qZaEkqJpL7TGiSYCPdvJN2om
qI5BSopZQPAUnHvsyISwB7qEjAkNJvD2n/7Swjj30Fnq/X2Xn/gLSpKaLi7g3Y12
xKtjFQ/Ylfd6BJ1DHe7+F9bGjxym5nZ4k1L/gSmohyqj6afKnDwL5O+35qF+dFXN
Ra+yY/99SGlTou4Bvyo8D6XNDsUnrgGvyvzzGJk4RUh9YhszceQ+cwsRfIOdSjSL
7t4FKVOaUZ2tDQlhaCVtSKm1sKc1xAuXKS3Zo3Io2ySoQsuGOW9WYWAAyXp7rQ8l
Dk6PzDg/Yb8xl4GBuwy3A9XLskBda4lGblQ/p0DxCy2UgleFPiibPlmitNkAD9bp
RUBBt++/YHp/CkrUfeBeCZiSJ8fp4XhDxFPqHMTu19xkw7ZCp3ElvGzXfLKwsg7W
aMK7BGwtpEJ+sRnAmjPtxSMfJ16g1E9p9hK3OqL8tMOpTP6jbbCh+f1ZyvqI0Hr7
bjDSNayg4abzHeubiptdYW/ou9PBpwSTSXLtqzpTgYn0s5KuICu8viZLP3Ky1c/k
PqvzWM9ptWaetP5lXTu73Nlf9ULpy8nhBCH1CGO8KopIZb7oa3XMSVJwvgFbVJz6
4rETXvv3UZiUMO3EKFtQQLupAav08D6J3ipQOWAfOP99XAMYEB5lCCtqsTb0RhwX
Tgi6891sxADlWhSosfOqPXAv1MF2MDrgHmld7L3EsyyVAbbs0md26QjCANaYqEZh
YZuOP1gzTkU0VUhyYUfbxm3LxvKqZh9fmaLNgL7TqHBQHM0Ft9pojBH7sEVZ2CzG
MYJHINlNeIET3Pw0+44aixZn4wB0MacdAjY4XikAE9gvDvrVptNJy8khk1/aEhe5
E1Y4zbeUO+640nY3hea34+TG0dWL50zmoh1+661gz3hi9NSnPIL7cJgJKEcZpwX0
IlIZuklSNVByJSa6NNHTfFQqUOYHcPIhvoojxGeTy9AK68m/ELfiGkuZZIYAeTcG
VVNd79skswUyT6OqCtFqgwm1cAVgG8xJAEhZ0eBr/iUWzYZcTznUtfnJYtzovkzn
hKlTMgr8NKra+LSK+MmCBPW7AGahJuXi9TED8JTTIRarrCUcvOvgSH0biNFL41iW
l3+Oh38yT1AuK9smFsO50V04LY7LHrVM45JOEAVryaZXfaxMxg4u5U+cZ8QjQ/MF
ZB4Fm61jVJzUWu+A1LdTVJDNfMWttn8+LC9R5Uqyj2R4tOOA5xtpbkSi9Fmr6NzK
X/NXvw4P78cB7lLY+LMGasXYnZ5I1jqM/9I4M0WTmWVQoAnVXhiMU4es9lKxk7ch
n+JQXpOM7i5+skVSAqLELM4a/cl652aW5Qh8kbY+ednpMxKj8gmtGNuddzH3IdWX
UlnYUmXG4DukzsPM3KQjS+9mAyNYh/8fhmSUUJ8YrJUAHivwbALEbglg/PaOg7VA
TYfwRdf72TtjFq459FAhVoLbhsi+tjzIXK7gxWBfqegZJDIW3pXakjoAGH49Bfv8
C81L26T1xt02/SF6QL6+Pb+wE1UpbI/JqIDi9xIKx9X2dQgADhNhxdz8nKxPUiBy
RzNBYixpBV1nbdKCvNIrqUs8JESlvyQon94uvYWNb/BSBVQApcIWrOkL5XZ99E+n
tDP7j+r5pr6ECiRl24wEAZdCqrxNz2EeiCR2XeEDeRi1BnqOYHLeVJICxTMuRhSt
tLe87egwivNFXbvxPvoUu8+gTeXS976kJ8eYSDqyUrshGu7okSwiFVVj7g5U24Fe
f9+UloZSzC0hEfZYS0ZthrqGQ7Eifl6fN03aLANly6nOxpZgMPKYYUr9APUmTcgh
/isM/YUQOOgHnxorrII//QKo6mjPO7DjgoS0agVdvzSZC17zTht2tt5KvGG3cK4C
9Zpkoxe5i0v8z2zBjRGst2vyKbvUXrc1ft04VYYj360enmGtjnyv+Tc33KYsTUmZ
9g91KfD1IIHMtEXU7XkO4SvVKoUuRtumg2z1EiWAtt2+92ZG2SQIU2xIQP4GYhug
2HvHUtux63ODEo3k2QrCgpG3ZFQh74SVGcTRbQNne5zi6v+Gpqg49aSOHYbeoaTJ
rvevJ7qIWC4LwxVg6f7Y86D2Z6komtcxGqkefBE9cpCArKam+czv1K9kMKA7dNNg
04nzRrE1FMtyNGf/T36f3g47KP4447PDXac2USsQ/Fo++4jc6qelLpPA0VZpUn0m
jWI373BeyG/oJRFbXZhK5r+3WgwqIH6Cpc1Bj5/NyMR2xHhEIcriBMNXMcT7Mc+J
yj0FJ+2kxtdHTjUbAggSln8A7x7UuUc5AzHDeD8909Njri8pw477xLD0bvcpVU4N
QfRbO0pwnikNTa9LEkwYLSkcZ1Dc4EjvZ+ND9yKHc8gNlDV2bHX+ccHVjdMSsIBu
qkomHudZrtGRQfeMPhxR36bZHks3ujX+c9h8KWcKVca1rL6rUhi7brJ8R/HbqQqS
6T8TYGZuTH8+0lCD+pakShetgh6n39qtq8J41fATV0lyF8bMJH/N6fgH+D9daX+n
+Dpndkwj6C1HWDdglSD1LMUp6xEJXmIajbQD7nXE/gFanf1eNUM826e4pm0PMMtq
zj28vG8yXTUXm2XTHrgPRlU5v3Hn7Q7BwkDHDSwxeeMYQFGnC3vQloeE3C7cyIbx
EYieZk2/is0RGLH522Qw53wjpnpHqlK5WvMtpPMy5OQPTdbFsSLRZB2bSX4oQ/td
8oYGG940OTB1QDCc0IszU60/Wr0fwTauRRNQK3lI8K79SifweVtZC/iZpoYaVrQ+
1CTRMCEUZ8Lv6BY5Ry3pjvfH/cew4FqtOwTaFKp2TUxMmAZiZVTKqBcWQQRi/ubT
i6LuanEuUbMwT8j2zAiNoKQIAaU4FBsI1eiaR+x3a4n9r5/HVBbLeDfCiqzV+o6p
tUrl95s8fE7SD9exSjNzi2LJAD4YMA22tp7B7gc+dgu+4bP+DF1w6z3ADAkK+xO9
j8AawRL/keTxcavwuE4eFFRj00uECke7QLMPhi66N+C8TMCaZyAQjtwLwHLio9iw
FjA0CTYWwBUhX8Upf8OHI5XO93E5VuXElty7Ci4SZcKDsrwjkdVqLYDo7sFkkz56
O3mP1badf4CHmidoU9wBi7Z1fuSisCvi/wuR0Q++lcHu2L6S4BXTr3EoY1QtifSO
TPG1FmaK5mrhV73nMQqpXE7MzqdYOR8N+VuBAf/OY6Hko6qHIM4SwbrxdBAnW9Wo
wr67ivGvC5B5NBNHCSSaAnb5KH2wzGgFWM89JyulApZUQNEgupgyQEEuv3Uo2bwf
CnEano0BX/8tPbbK+XLEsCuf9kPY54mvZoIjPICBmxaHA9Ns9naNDPBaFDy/5CA5
+RJTbb0TYdvXcJ7xCmKdHO22R5EAiK7ckAimWvt1anNe9LMQCMpymscJLrf6o0f9
Ot4nnXl6MHdki/3visaWdJjlwyZKwHQt5MSQM1+TOsfYhO1NUw3zMth7wBmyf6tb
Sb/js49AyYZgCLahKPvhE3Nktv52xYjGHJqbYba3xHjVy1ePGRKM3aYyktFeuwIl
xIdlt6RB9sbuJknp4i890vq0QRqBenINxz3AxiGu4an50Mra8zhcbrzPklkub+3v
SDeXDqIv4RukOjBbhwESmad60hQ2qASSmvLB64CcuCdo7JnZ5kONTN7akPNvRG4G
bdPB1Ky2Xwmn3Xa2Kbs2/E103sNosoib5IHDRrPX3bdATO0B+OzAMUjUAmLowNUu
6UkeEh6RuwMwG5ZO/DQBa6juNnoWynDw6uHa/w/UaV/jbwjO/1XuWjrH/0OVFqSp
S03jycW1FnFs8MrKDgc8ZW+Qeh3SBXBjz0sPrp6dEX2foGIyPYQ2ONCvwTXBx03d
U9+E6tbY2mCklhrq79zT1l0dAkb4hixAW392qSeYOLIAJb/Sgt38uMW6H/31w8/A
fb7go/uqsvyaFDIf8TUFFSWlSjyVMIxgFPTDor/Pe1i25DSQHyuhck8hIVM+qiY2
nwlzJA0eF+FFS/rfHuVpMJSrMzBiGHxxsBspphH0h4nyjJ0s5s7I4w5P3NCASVDt
qWBC+Ky0KUF5In7iM1Ahk6McjGY031MCKiB5gVTRr60b8iTKEfCoy+uflGWcfpaO
Cywa6ISEA8dPAhnr/oGCvYHn8ZBG0ty4l4yQUrIHiZt/AWb4t2sQWHs/w8nCeZoA
mkKrqJkRdOBG4baTACunguf4mY3n3X9i04ATExMOwTGOielozxsP2kZvOyb+C91Y
VB85NU8JIV+4zGi1KEOytvx+a3VDRn6KKBtUhSCTTTlv4eYYQcXFsUJeuwat0vGV
135DE13rj6ruvZ4ohJTmQfJGhTUORk/EUGlvkt7tA7U0YDEnFbio0nOaefC3hudz
AZ8ZwJqtGLriY8xmnlCfAhIxBT+a/WeSLGumUm3KHSkxdl0DKor5DJranzfVN7kr
HNgb/0Vah3xAVxKDfeok2661X/GcgEi+VC59UHfgl0ktZc/ce88pJy1YjCFTtqCz
UGDDDYrhIu+6RvpfQunbdW4ng90alWJfAVvDBz3ehYI4XKbnwvtvU+FBS1TXPDyZ
rWw/sXd5qSRTbIwL0SHvqWJKgnhiEnhb0HVUCxYa9IJKVhcYey8YYPR9DKGOCPmW
PF7YNbcBi/hCGIg6DQWSasE66/onjbkoRO4LGwc1s4I9EqBXUAzS4rjngMWup77d
3LIOtNP/aeDFaG9Z2UpFvDBnAmsX5aNcAWGvC8miqs2zmp4t6jH15VRzhQ2cKUa6
RZ1GTol83EUtU/Ee/x0hZNwmg12Gt3w/hCuKVCyhotrouAi3RbrAAXV5sW0/KUPr
B6gUmREQh+e2zg2T3Rhqoq7+MEufqmndbU2mYxsuzOWkQIncc9MxBNnAIx9yIRIR
lzccuj68dxBKXpUHCndDuHk3ab13PkConYNrWBZ5rgPqtkyj7YHFWjd+1w9N1bI4
7tXtgOXnuVDngradan/XnpgRKMK4G+rw1EEk3TcZeK+hrcHcfeA/OxXbUa5I7mwT
B6HFSDMEcsUQFXScHX+YFnMR081VIV/T22Y9N24WAhZ9P760lhjdEj6Sb4bktJJB
DrYASun2BKGElBzNAyiViT/1WnwqTNOuTJlTet5YB8JJGNWRJMUI7KVpyDUrvf2L
PWzF0d+P416Ve9fQksIQMN4/YfOxhIqMuJZ/eZNk+bHKlqMx8GaFH5/iwtQG1Hbg
H8hFBdhfgHtvmWVUosqo6qVAVJ743DEllGdH6Dk4dNAm2Ry+W/2eGIB2hNncEGUC
D5cNJcD/tjijtl0oIaqpbz3RG4XL1jblRfhA9HgBBoX5jYUKlArOxjrM374UVrtZ
bKgGx7GGpxpZYTYcvORIlXR2kR9Sk9BYw4eV5jzhRHvAYwCBM3IG4R4HBOejozHi
NLL1dWpJzthBTiw3rjgl16C3a4/+C2IKzqVXuxMAewQAObX2KhJFEO82+jaW5ppM
gBYto8xOtH2xHCXCAUp/5BY872pgqMwsUkSlUW4GdkmgMS5f7tRE8vdpqjnsM/O1
cUZOPwY+spjS6NgV3aZNMjNSO5V3JNTSMeVFj9d3Pndri/+Yy1FAId9WWRD14HDA
bDPMkFrRXyb3TWrLxqLyVmVL2wXTScwZPjBw56642Yonr2uDQ2kv2lQ2/qTlrbEQ
14+0skIrY6elHq1vGEQXAj3VcZ6Jx8+mdyBthwPNfyFeh4TZC32uxfq5sriaQOa6
hLCycDhtU+ZoCRJz8bZEpOpI6JvYmbqYQt+pHyA6tg6bjUbFhux8ZvA+vH7ACL+R
ukyxKk21j5J58mtceRb1lEDJOUdLTzKuAE5IkeYmH+Wh82ZGiFfQaQhF+5kUc3Dm
cbvVhgCUhd+c34V/tOGwLLoWKKhk4Ls2RG0A4fte0a7rdS8MGAsmiZPhmGOP99Oc
FutyXn8nDjCo1qeIgZAFfqXcDEPWLisscCEyyElKUy3H0SMU3yNk8y3u3ZCEzjTA
XFZgapRLNWBYc1FsAxG980WiK4IZnvi1Xcd6evGbzoKxKrns8ohXHnYcGJ0E/qsk
Kuq+6LJA2tXGED76wCz14n2P9KJGqPkCDXmvV8yOqNY2uZCQMhuFcPu/gqeJPpyg
GS98aYIIwKmlEXnpQ5eNag3J3rcO7zEPETi2yRn2Pc6QXNKmvVnGVGEHCu86eqAr
6XOR0Y4IDonZX5kiw37AHva26XS2DaFF1jBBak842ECCgCISuN/FOHOqrNUj4D1F
e3eSlr5ir9pvYjZo5FshtnlS4GV2GF30HxE5xnkEJHvzKcwQ7kT34lwmU2onN5Ea
WN/AVcxsYnKRUDrlBMdE2FanHjMRNCdKJs9GtGiBYYTT+acaLIfn6bRwyqDSjCBm
hDY3XS5RdWnz163VR3KHLfYX25p7RXLIhGNiWl8tE9ALynYN1y7kuNgihHO7sHQW
nyG4WNhLkfVWHWjX6kLXsT32imdU5r07g74WjYlQ7SmBhOc80ttmq/TDqUaHUShd
C2mLFAyn1nzaWNgoz6Xrk3T1NYci383LFB6Hlb5zHASbHDLQWOUO7fNPy1sAMu1j
bYqOOc1wJGqpfVkd2gKZr4Yvnu2JOCAODkUgnStaJ7PlrmBO8genIj2eXshJC5zP
7zvfP/GMGF/iI3nmg7nrbwvYldMMMZgkQ//y2dWjVjH39vVD+Ia30YRk2EFsNC+L
R1i1A+MbhB21hVHicaFM969mscE1SCIGxgvtsKzFnxWMgLVVQ30ky5JoQ3wnoBwW
y3wwpWmsZl64aiZPoo+pPcIID+RiN+fg4WGUbshxWS2pSs1nRZgUuDZg2w9sVPTY
r51YlBWIZztwgzkvUFgwlRDuZihiWbZV/rtrKweZWdWWC5KsQ8hqj4JxEp9fav97
/9psUop1moU9UqkHeWuw9VnUSiKHmRNenLqZbT/8js+Mkgq6FzuEQAs8du5UyCi9
7ONnyOlk+KLmsVR4SiK1zGkCvL1nvXAj//FW8HYlSyYyov3fy2qodYJn5yKQFeyR
RmamhL1ty0H8/92p0BnfFum1e9TNeSC5xYIEj2bfz5HQXFmbKaeHugajonT5bzWF
3TCYFxG+J+fvLwU+HLTpe9yeMHaGnHG1h3IQSD6e0pRACYopHB59zMpAtE2/Aqck
0+qfdQpjPnb1PSFG9lCfo4LQ7Cwl1KkWoxTpdMFVEhiCZRHqUyEtjbSXYqXfgFAL
3Td66USQehnW5+QbwVnBm9ikbBaP3WGOihKipl0HudWwpGmVYkrF15yVOjE8qokQ
UPH+fgNEJ9rSaKSwjuoxeTRzualasvDVtyuwr4AlAj9Of9GNLE04IVrV5C4txvPz
8MDOyZXIgT8cKmVRKopa4627BdAaH9Ngix65I6q33zLkZDDgJ5i/EAnITTqxFMLU
sOCgFvR77z2O3fuYcZRFBmHj0AiNlKGB2n4jPWgo9nxdlb2g/yagfh3EGPZUdg00
vk55Bexc+Uj+mXnEtAQgxp4To3cIQ+PrJIqhZbq1DTgMY0jzQeY50f/LfELOxT65
h0+3K3f1xmqC5R32ruTUfXY2DC5E5XRFpdaxaVB+QPidOj79dj27wf7cjbK6n74m
5k8rm2vJ8zSsB3S8ftmzXHDW8jNziNpbVPlAsGTFH02/N9KH3bOogdY+Os4Q3EH8
ePkHNMWCORj0Kn5a0RTh56uDZSe2MzQb2d9/iSuL4hY8smhlQb6covkBStuvSu9U
zDju7mj5859/CRf2lo+lXOrVV8R15E6HsKqDE8bQfuW5+xKNj0tV+rsdy/7GFIsw
Yz6h3NeAH8LOHvJGvJ3nov1q5AoKJIXjXX5jDeMMZnxxoSgG8ftWBlOfXFMfLF+x
tPyY9e8e54dTSgHfx7BxPjqDGyrKC5F5moghcMAh1NAGr50T6plGogXwxMiA9Ff4
BUVdSj40l+4H+3NsOGa1OLDL9kgvFWvvUYOUs/RjBqv60XPBFOx02konRiWZTRtk
NPawkwKR1QkRpJ6rpaD56kwAt9+pfXXu55t8lT7fpuds4yPXNfdzvpwVqddVKidx
4GNyZ9qbPH8h2/DWdfjVLCTRYmHaCvoeBq2GuD3aMQFG02/3XCBDATyMdwAoVdl/
sDyf2NmxFOS9RNtEbSpeWEaT/XeUgt4EohHMrbpyxCfCbWu60bsu2DXwje0MpxYE
6m55a8Gv1//qSeytyCV0YFpsN+PH6k0PIiBoRvV4gxmvh+nW0aIU7120hdWUu2v9
lt3tas7GzR357WSMp09aQqmnSN+2WVSl/rozmHQ1+l0HtxTwwzWYL4tKSvFkgAhm
7Ofq4XukWAI4ClOIjKOVMtMdqfWQj1WFUYMPNSQgVbKN+s51R6kGMSVE6drcyTeJ
yNlaYlGXPDzwRw1m+yLNgT9sksqzIBuDWKL1d0FB/gVUlJAOviig8eAEZTjawTst
ZPKmS67GnTtOkk6hkxGQcvQx19koyrRyoBqphetk4Oz0wtQAogcwjJbWXEDaunCS
QnOcTe1aMIJgyglv4Xarzul0hL5XnReV6M6FdoB5CZOKzHv9T+T6NiM4rznJkCFM
iVyhjXwvrccEaT26+5vh09pX4mcnFZ2IUFz1xcsyq+zxPKDjHDTfvorLLI7F56k6
p6G4eXzS1PZEHWFjYrg6eliME1TnNpCmpP4waEUyCHexP4BJdVV+864KCC/19AR6
WKSRLwkgKJEQf/cTJPj7W4L1C9fksQyRHw2uDgISPHh2jeVBCCMPkogioX20Ut2+
yHOSVazSLGgplgZzDYIerwbgchHyvusl6DPpT5czcGOMBMeg2uirauj0IOEnCY3Q
rxrMReyNJOr0in6qF123j+AjgQOk8/GvitQGLIxSAkhxJ+baaH45Bdpx1nZ6X+E1
f2wD4+U4HT9QdrCSeLxYvOGAmUIm2v5jcOYqkBodKrDQ2FGKmoCGB9xt5MIZ8+hr
BjGNEslRoV2ggz1SjWAv6KwvGD3zkRKW56/4pXkKrUHSYBJSP4Yuh4+P4eXAKe4n
E2Vfzcmswf8OW9yUYQcbgu24W9ShTSGjQ6ADlplaIB/6y6Ezgp1Jiqhtjl6QCY+I
Pm0yQTGR1dDmF+mmTMWkqZ2saOObyz3lw2mRPEAvoR0MZU4ngYWVmTCDZogNwgAm
pOPQ/kcGBb2G5+9BbPO8ZkLQVMvtUg/3oAikG03PCAh+7GEI48FWjYOkvGy71VhC
R6OvAr25OF4XENQYjzl0SQ87wXy6zgLy19V9c3PhtSdaiUvFA1znmiXP+niTsZYh
fUKAxV2VBYozuv63hx6re071+ffSgMI576mtkF21vu7QUC8Nrw1Ge7f31/zxbFbj
YAuumDhHc2ef83ZH+wYE9LQi57ACvtJ5jBx3WyQQGFefBTizuJyjUO0+qBx+X5d/
Yjf21mOIX3M0M4nnNRnrl4U15D16wMpChzAeed95tNqOIw1tpoEFN+5xIVdqiZPX
ZdAiRPOsPrYNpM9dw6cmKfYr3O4RODnWU5H1ThLn3t8CKhoHEuazeeu8ouOaCo1g
RTW+86MLy3jzx9QAkaYBhYFAYuCtUduyoWX7cYPSJnpzc2+WjMdYn0fpHDHCPeCv
9yBenmE2exRXYbuoCFDET8NIRkZpvc61jYtSnfeVlw7bBYiIGq2XcPpiMLco7f98
2CUiI7poSg5A+qkQyCuHI+9Ffv3h0YYfoqg2rQvEABW2nDZeR37io1rswwn/lfbx
Oki+AYWiq2jnT8Kre08sT7Du8ofv1BMARt4bwR6uUsDcqltkJ9upZEMEH/FMGEjg
uExjVO9udv4bojUAvKodzbEPrsdImwKkRkw22ROxrVj+vaUvmkRGfwtHD8non8Jr
InSpyaOn1dmojkz7prATCwi/Cnm8dzDcKaEuOP6SfbTujTxznTLCqs/ys4GBKlRh
czkT8IO/y8eN7h4eBBs6+6H1EWy1vCQbwwEfRKNgW7DyCP1i5V222FqXN5WJ0erj
0UZB1dEH6ytN2D1ot2uIw6ew0ekeJMZe3WDR297fu1wP85sXi5Dyke81eyUemYKh
rDnKDN6wFMI24OJGh6kWQBq8tNyAbBDh0EqEOfS+nD458qwcSkeqYsHyuw1lmJqu
QnR+tuqWjd9Xh8s8A4QzfXD8abuiAT9U3K/sBAbyLed5CBZl5FcVkV0GQBJ+P1fn
O/pnmfhQadMso99xpSWnu4OmLFJk3phNV2mDX4BFstKkdXuClUH8pnncj4u0d4NK
g/1Sh4a3IF/No0aFM2Fy9KV433L3t7mALlWmOb382e/lSfg45J6cTZl4oBu9Dhyv
xMBZUcJ0p9GdmuG7KHaH49/DLOnBZFoAfjwWrExF+G+XaFoSmaAInh5BQQ8kB4PL
z6gmDleVTGsFVVKmpOHbk729TDBaRJZYYQorF8SKYMvmmOLzGWQoyUownKDEptKz
xbLVBnvFME6UcQuNey/G2jsgXxumPr9HDCEWMADeI1hskwsZ+M5hCWpBJxhvKdsi
JEfGWB9QpZqN2cXzTlOR8eOjIcB5GDV0G/ZMqk946KPo/Z9ULIWDQKrFAbMlGMG5
xGKLv5ibRxyjVGg0NX/kl1ZUmJ564yqkM9VRb0G4qMAJ+5jFpnPAsI0TskjyMnew
F3knktZ/wAAZjG8kulq6CnIDeEwE0Jpk8PeEcNEWVlTCdU+n0wWucQbbDuWnlmHO
mqaLaPh03YYn0T7/hveUbzex08uigDK23ShMBK/rhUFayXYC1TGaZEBAbs7Ykjco
iOCIg7vETqKDBWqmX8vtaVuaGm8ETxayVQd6AfdUM2VWQe+LCibtJOV/4oeyHoLZ
sa6HDKtbsWf5cjutR8Pk0KwM27skZclrMeBsDiD0jmaEe+wqwJ6y8qXVcUUUYm6y
W8XCY3r+1ad4ZZniDX8xoebi4goM2MXkj1iinQkufjrz2q+mqvwbDCalTzFY3O54
wjpIZcNbbo8Jqnvh2L9j+A8iLZ+FbQkofFHpQhG6PC1OTA0cvi1hXx3G54wBoT51
RFhiWMA3XlWLdC+KyJvPaAMp9+a8pFqS+XH4r7xIF3agSDBBAmnLYUdKIa4CYsPF
FV+Vxvy02M8vjcPWMiSA2SXOLLtNyNmabEIqoHsa7AU7FzKWvVVBNpEQCuHVgSLs
qpXZNIUWMSapNqw+oEsvhImA86O1pwGs3zajX7eJ1wDMHJ/u7OYZHB9x8qz0l+NQ
N6RmX0VJ7/QdYacgB+7bo0SNg0jS/NEBGECNHS6DB3Ne/kXK22dN5LW+kPjIcypw
9pu4G4VGKPiO2SE2AbYLolxLKxuOneXt5Mi1q4/RNmYarZ6Cvk13jZKlibQ7opA/
sJjPr/grnIKDSMRFTYvRt180nXK+Id/6tqPjaRcw1DVCKzBlCiKk6JN60AMtIcSH
EKqBbfLEGWEB9X9u3WYd8fauNnTOqbTuiHtkA1mOqGe8uk6vlNCk/Iy0cA3xY/NH
SnUV6dSDF9UaHuwNls/weM1KsvDIT6gYOaRAc3CNnu6vuLEXQjKXKahbkxkox5ir
s4upeqG3dh/IXdLnvY3/X5dVnuk7wo39hXT77v1Ve+jqwsnv9sxA1ys9pBfCSeMw
woC3ptpL152XkOHL7IeQqP2Fa/ydgnUdVeKf8TVwViC0lMa+5efZIW0IZOUbYGzw
L0zO/9PvWjmrQLpLCgC6JFfBsa8HdSUtZ+l1mVApb8gmliNtOy9FltOZXKOCP6Ju
GEyDLWwYKgITib62oj6yAVvW7kZG3eU8KdF2RiZZ4I1mk/b2x6eRAlio/J8noxd5
oVad+4yY7ESgznaMm7YFC+caDxFKn5yh/hJkRU2vqDXJCHfL5bAEMDOZBhYPKKPI
zVl+kJ7xTgCjewPMC0Fs7+sO2fQuT9VhchkTQ1NLclPt0J4RMBtxn4lD1E8/9tf9
MMOIceaKTeL0gXB+kwip5xXUfJdzEpuSfWsY6lgrdnj6uq093ecL8fJJXx3Gf9us
go/FSlGD8V928ltrozjuECSfLlJssN2B5DnEGoc1CceUzirZ0XrrJIFl8BK4GljH
RHXQ0Pm1lgIN1Vtz2/H4Y+Xn/lg94pHg17xaOb64GtbzUa3h5yB8hzstptqfs238
sjES3v2ePl2HZxm/Y0P/zd6NJDoPRmpQaXeHmLXb9RyMtIEv7rd6fCdm5c+Lkjjn
Kd+QEGICGOP/Y91p6PpABxIeYMvgYlMk69NH9fjG5U9MxAT9TUbV4Z09CX47AO0q
uUgCgxf2oMcHaH1ghgt8JehqS+LRbRFi2bnhDpEivreLLhetyANSXZhKTPdlBz0W
Xi3ICy+1hsNR5kPvqZLmGipHeOiVGaEt8JsLldYh+4v1DYSU+CNuZl2eK8Pm46jE
+i/dBUoW0ARhMOIKV9fR1muHF0YgnTfuMg7QdbytFYiIfgJH4rrK5gsyed0bAvIj
Ktf7Md5E8Rkhy805+Pcsk4JgDUSzoRiOEpshpyq7Xu1j3jXXI6xWnCWFhzE5qOfF
YmHEyUG9qkVeHni9EFliPCZaKrEgp4eiYH0Zn9wxMI18ymTKU0o7ITq5FbL6/cO8
5vfoZ01ukiYgLRZTk5cgUrXuznQI2ZGun2MyE4NLdhXDJGSCJkMfurGHzCmAxv7J
Gx+Mi+RDSbO4g84S1cOBPqFPwoL7lQWLARxCDGQ4celRlsr/mKMG4zFRu5he0Hyk
UNZP8mQxwH6ZAt/Gy1MW8Dd6PKBnA0d5wcJwZfH7uEGT+w2CtuZCq/E9AvcCmt2G
Ujp+UyNfk9/Gj3aLAwWwLcn1T7rKuyiLWQzhNmSoL0jJVACbBBYo+3DFzblCHnX5
O109rPY+t4c/C1gliGbbrfsHOzBe7ivMdeU2BUpP94p9O7laChK1YORvwB1t6wEc
eOG/E5ILGNdy+erjSWl7vQPZHP0moGhuceYCqaEFgyQMc1iq7Y69c/LHyMSklkb3
XrZe1dfzZFw4lPfiGHydgwRZfCLFLLEogomFyfoeGggwREmLxkXqtjYcMtnCD3OG
efpGJxIU2GjbZgtaeZETNxYNC4c0P+TGBSAFN+r9pPAi9hiBc2Hdargm4dJGW3Bx
C1+wfJpdEEah8jHsDs8kBQSuuBxJ6MJRWUIaG6ElSL8/aBpsuRY0JmXNiipsDOGO
ni+o2YXQOafWtcJe3B1Ixne49ZVMmOYTccTOU7ic/+URhRxRzDteyzSX/vkFA3BX
lttP+WeABRKF90C3YV0GlKqLMfg9B30TfZAuKa5eG4wWZgYS5yUZaaxMpu/teHQ5
y5gFek1HhEt4KkvVAXpEuGLc7S3QY0SLUmJas9XVmBjLBAdK4ZWxk+KAYfAeqK8J
zT6SmQHo4MeZexU+QZLLjqEpm+yU35dmRZCNQU2a/+Tev4TbpiwrDjNrG1WStaR9
9PKgI6fSkVegOjUc+wf+ilO6ePfQxGTo4/CZW8dWlutH6RvGqBHebDfUL94pPGKw
SqiSJgf4Mq/u2yGRZjTUMAvZVYOwrHw1hzLFOb4iVYCPUCYkVahR37UD1pf89gkE
Yk0jiFqag18T0HZLn31Qgiy0z5tjpBpamwrZTHex8ORBUZLd2oySCxmGjgEEaDhC
7wGhXm2ZvkWTjrhLwSYDvdhvWA/FBAmfILB0p1a2r+qlRHM51G+CiaiZ41vhvjgG
vFhtvODOKa3jIIKWvQNxQIrJM9dbLAFCveIb4sRr5ZuW/in2iiH/G1mJj8MGEDb+
A6H1reXWNmo+nV0RQDDjvlzpX/IksI3UDYoHdzQc7xp9tugRr+NdCnZz+u4H9hCU
jsw3WnCOCZ37pms78k8VXfY9ran9UfQVwcWFryLjKuOz0hUhxm8RXfe8i6DpMPgi
eRuMSvRo+Jk7z7Ytff47FUQJpUkiw51anmjO3ZOXKfkohNFvcsMIQvGWYk2PUQ09
cE6LeBJw6sjXwhjxn8AJrrcWdvpYyhDlY/o4z/jryjn/WGXs/heuvC87LJjL5ciY
TnOmKSrGt98gKyZFijUTO2hlPucA9UzWM7iCFkU5xIAALBJYRQKs02sjL3YaZSIe
qFuk+zpTQKXlubzclHz2qA2omjNfzk2PcYBRuXIBXC0htmfJkTc1wGoiXZUFOZNb
3UIljw/XxtK3LLcIzXr98P0zVlhe7G3l41FANXEX0KwK9H1slU+nQsWn8VrB49co
JQSMuOL2JIKMnapt7Zmz8Y7KAbBpHcsP3qv7V7I7m42a8CitJldtsGZxyt57DZci
3BvR8iEvfIXxvhqrvUMsj+Y2Fm3a+eclv+gxmC2fUJX7YAQpvarCBgsxVRtY5xLx
U5Npp/qcCDCfIemBU3XG9FEETisFa1DK3YY/Hy0qwCsWHsnh6WmK8BdvvYoc6c8j
PUSV0lkx2hJHtjgXzR+A8ytesiNAZvuNUXN4MBWf+IbKpnz40OuOOEzNH5JiBnGv
l2J2hQ9Yoo9dpQ9xrcsXGnlYFK0uurVZR7Q62StP7h4Yu/92IFV+2znaRxIQbsNr
1xIYTBtF99WGEk3CvxJQdH297AeP432udLNlxrWITZ5s51IuUAPnWOM2XCWjIi9y
/xH+q53cjof9ki7Bz8xMvF3Nm9sx2ScluNKC+6n85kcORenupxitFgg6RndTtv5d
GhWfo5RK70VccOgriieWCNNr1JdlP0bWukLbEz0BNASChXtPvkFsxnG4MmbS+DqJ
llGl9L5E3BrqptPYh+qZNoGVZ+EuACBIhJJKG8/FadkPvXEEeOgG98aGmFcCAII5
9K4PHWLPU9NOXlKq5OKYAxaF/61ILg0nWEsnHDOCIpNQewhzflhiSjjmDQQ3GAg9
4uMMVFEONZ4XJ6gqS2EhBOBw6wvCiYk04F3PKcQzAyzx63qu/Xe70lBzkbM4wtGG
pqEH0h5MYqFLSeUyjQMkTft2Fdvc9ELu38H+WX1pZut1XYbvSvQ9Rm6Lbe2bYDfS
5h/q9m5lLPbWFXjzZ2Zm+CGNh50yGzaC025ipx569JhqMpF5hXBOsWN1JUIu5Yfx
+P9jt5b2f7g1MjTvXu7Rv8fqRt5wI9WXtuJGau21tQEBEdl3L/QFwQEX2PH6joLr
uUB8uPAuFTWY/BOJl8iNh1F2+IpPvGALRAEOJXs5Bah3GqutluIdC5LZnubOEb92
Ys++9QC0yIXL5QeaKvHMUzaS3U40abyemFno+puRB4RqIbI13/N4tVLpJ8mQhmij
pog3jGG4MBauIjvgbw6EBpNQw5VcwqtBql8Ey9hxzPxy6EtUyLIAFdr4PLRlkHxi
O3kcz3wLFsSDVcJjcGuygIEH5eyl0kRf9WppurWcYPiWU2FXA4xD7nAxKfOTnahF
Fh81Zq/IahWFqa/SzSrQ/ID60mmwpPjbx6YuzYInouuqgTESCrt4JmDqhnQZawJA
0Qx58xi8yzJ6a2utQpJM62BcAqj8MP5qyGct6qQf5tG22wgqILPgREFONB/UHAdp
2QwdRgjGo+Tq8bjU6USRaArNFl5tCeD+THH2Op/4DmDM2ed+NomjdtR5U1YC3+BY
oyXueteFwpiMAmYC3Sl8fRVJBcnV+ZYjazrvpJrXKTlq9hpi010AUYx/cdTDTnY0
0NIKzQbaHPzt0iYaLME6MphljlFfgophAnoefhvpfT2Zksy7zvm/vk5sKAG/GTV+
I/Ad8RewPGBFg1MIJqsh4Xe4Cvky+N+FzEMZqO8aqShwkuhUjbwxUwV6iYQC3fEX
rXfRvdovRyfqxUGgFJM1D1bBUbJveL0PqC1tvyJIBLtPyjCv+knzKo0p0MzfV6N5
d8uStBC8s4xFZeRrlwefALfi2rmItWcqOzlRB84qXhaL66eAdCnJEaahF9r/dLu4
GkxXDlUZ/VxxLiIBNVGOeW91POhnWJ+Klkj0WjB9lBNwv0dRVgIH+7bYVdmdiL0Y
3tGtR37mQfBQwSVbBUi/rNa4Txc23qJwYtzMXnHw0sYlhToFUPoGO7I4KQxxvaWy
QND+KYxuKPqR2FYdke4KIZagESVKdWbzeEpZ9osBLu9TyJEdWartTLGg9ga3iIlD
ScP5Gg8qDFwRMOCgisR2PqjhGSTL6rV8okQZn6atywelsrc8rCyUiJFHcydwG4/9
8CZN76hhWaa4TBW+XoHXgQqu/ccUiTO6Grvux1mOZgQGIJOv2wZJABh4Je1+xL1f
x8C+GSMTiCDvwDOXbYePG3lsuFvgyQZTEBH8TSUPXZ7RnsM42X+AIaw8xaqagTpm
CcW/IdgjbzyHopICBpOOwsaB6avcsqRHMMoCoHGu5YONyi2mbS7YAEzALRp7TC2Q
Kyoi/QgWcPeFTk43EaIUI/BX62vaI7XGij8iCxb7Jlxe6k7O2e06FjmGpcFyXEQG
EunZ2j94aERxTelD1g7ySnuivViijFsNdlVCI+0Ikq/y1WyZ7rTpdgoAfgyPK994
1qSqaivQBk0fAGV6qmfRep+xhCn5UI7Nv/TeirJROvc6GQ7Qn+J5jqcSKZM8bHcs
BqIp5Xud0COuOKxk/UbEBJh3nlTNfSsRzdmWqkJMeHvfF215XG/7TRvngygw0uHz
eYRPk4T20cdNdqWIJ/oA3twCh0HiV6tyr6BjcOfH4bhnPyFNpDwwjr88SDkG+6mI
f2r18f+xid0alEVxX0HokKyqWjrX5/gqhsnRFcXm0/YxRMeX0Vjd1uNpn8BOoBft
cCQHffRaBPsTOmY27jYcV/dAzi+3NnLq6MdYx0KDKO7TV8SUy7dRyPcgn1+on7YJ
kVslLPAmusdltGA40r/xLoanxVOxyMs2r6LklcvTrcZeknI4BxBsX54BnehSCqo9
2IIatkhgm+JFK0ZM/OE7Tk7kvPWf29f3ZE8bpAzWp1E8MjMHBMrRNdaavoOAyJCM
t7Zh/c6x9N0qmC+XZ1yeWPCFTvH3WBX9v4A5CrnHlcNOdeeqCnA1RmVTNFynxIPg
oLHxPP8STN3iICNq1VUDS0mfBMXFlfM3ugRCA/7PaRNPwEZXaLbl1jKroV+lIozR
fjpgfQ6K1J+hEnRNO30jgsvuJql7prJxJCXo8DtJd3p3r/LfDaaGNeGY7gaBITkX
Dx55q4g9sq4yzjz3r8vBNUV79MWTY9Fw2+DoljJ10qt0DNk/wy2s9aTb9OS1Y+cy
sWC6VxzE/mxWmCQ8VdlutLxasxaizES+2FXq9Yuvztt6wc5pUGJED6jX/Mt/IgkY
sk2dDI//iYA1R0El7Od3Pk2Ury5z+9jlC86hgJX7Cg7r5ILTSeRhdSzFeq/9ZBUC
QzHdjDv2lp056Mkt9oKQHdVPNEpMz4kZAdiV4BTTcjMaZhjtrV4Up/iAJvPHDfBZ
XgDX85m+Tw93H/Hw0CQh8/UesHpPCcm88Sr/Wh0n2s4iZPspJL2WkT55qPIpoJVz
xI0O9SyKLtH0V6SW5Rh+vcQNULNHD62see1aTYGfBVpVxyBMfa/0nC13UmmfV72E
vgRmNAXYLZqJld3DLzZNa2EL/2/oBaP8PEPgVmtW4hRwGUYdttvMc26N6TYzYmp4
JedyO+E+H3ufnQfGLWLAHXzw1JQbfzHiYNeMUh/KBa6geLf0d6F++Pt2i16TT0Sa
ZYt8/k1mfyD/cmEIJZwCZaew4isFWC+Q81b1to8lPnG3543OEV1DTeg6fjVyAAKN
waZKcqevXGYBFSwBKRRtA3TndD/1y6AV9Zay6DGvfzTQgEXeXjwHHd1XWvjKALXQ
2A0K/LbId92RWC6CnYA8Eiao6tH/oPlSE6wFeoRCVR4dsjPZRJds8ASHvGvdbo90
ZaHWhB+bOFJFWBX76wX2X15cB40mdv3L/WgQ8CNKLTZpLrqaMu+QYP3jYdpxWEbW
wdRZ107oeDNg/w6dhhSqAV1FW03TWpYR0//I1GeIKLzO+uD+se10/j/uFe8UzB+I
W2Hj7LAh3e+IgB4oGEVxEp+g9JG8/7p+0U5Zm7A13QYyM1PiEjZlfBPQt/cI3jYv
083/Tgb8vA+EY6RUajZR11Q6qmZpDv/WdW0vdwBKhOiGiKwadHKyvfKGyhRomkTm
/MyAYpIircNaUI6FhNfHjbqt+qtoy8Bz5HRi8U70vih1aHIDARz8tQSiFUHZWSq/
xmpqDlHAwkcABQpjZq0KV8J19lICbBNxn1lKTpaOHDYPR0KF3JNic0LsCWz+9733
ftYG2Fa/g7MS1wpztnO/Rv//FTLlaQ8wrzv7YYSgBzo+/Pn711r86q9LZ0c5ksZr
yXjU+xXaWQSu67MDwbtBZN7VuRz2KQudzKIPqC8626Nr++fDYQ78/E3kJJ2orQI3
az5sZOhoZI8l5Uqjn53uo1yG7eiRIvIjjbC5jTB3ZFy8pn1/Z29Z2co4eJCXUlqS
g7c3SJZogXEKXsndsZ8mVdXhaBx1W0rAKc7PclJM1fJ7fPcS9xrbXYE2fdMAGgQh
etqdVVAOEQyAq2FWERSEAmmzL/3z++DB6LbHkLLGTHooapeOOL2yViteyULkPJD3
sFuiZn+Rju9OhMM/KuobH+sslQph3VLsJP/jstuxmKDrGbglB6WWb7MK1CJvZbr/
MKvlB0KAZy0lVJguY4zNOt0vWagGBoUBpnJ5eU1tG2r3cQUZVyzX88rNPwGSAnhX
G6krhjg4f89hBbKRGQIq84K++IT2SLD3xcXOHQhyiT+JHy5gre24FjJXRwpXOG1g
r3swB4/CVp3HDx7c/JfozbCqNdOMBhkGMWDPgiDOy9yq3t6IOZ9lIz8Pb0fkApXB
8gUSZ9aEZ4ME5ofVXrP8j+SrBkiam9Hp3b+U3eRJvbVl2g88x6l/NFuyJ2MeXoXh
XTkK6rqKU8ZBlsgE02nKGqXEC18S4l5GhgMa3jFMZju75qvHBGdW0vjcbmQqQUYU
7NGR2an9SzqNTlyodd9Yf8P8tPhYpyV4RMCRhxC9nV4/sRGT6Mgd+BBafhbCvY2g
IZO08YdPM4N4ORvBcgUgJ1XXA3MwgW5Pbh9J3OHIS9t4w5vsNCovfjI8XI3PAw8s
SZoDjYUnFrty8jwIoAwqUxoL7OK9Ro3/IeG19WcdJ1n37FpzK9tMwyeUNJ8e2fXb
UIxvswYiWpoE+/0iQxtF4wpniyr2BXxxBf2+4uEwIf060mj1aJFJqKOWQe3WE62Z
hrcSWq4cSE6fbrSj6GzU9foyHNBz7CyPzi2pzUQ5A/KC7xmkuZV3XeTqa/C7r9EP
1iHE36UEEstYBaXh+e0zD0qoizFkIkX1Tbozq+4HPYIasPVSObnT3ttqPgnkzxgC
AmsBx1bqWEM194zg043F/xqjL5uTkBkjRnG49xcS4lczbHe24RcRHXbmZqRdBeVo
Pf8H5TUHkeS+sdtbNDjh/3AKRRNHR5Z294wWtqQmSiBgwUMAiowdSX2JNG8/NS3A
EpBkIai4rpnIf/gTs0BV5ozhnvtnb5+qkdjlG7DOVCdssIChjBvPSQGS84O1Xllo
4Nt32Jj3wwq21VCQt3tBLJ3apbgzPu39c997FcmY8Hkl0WSwxa1UyXjEHiDGQab8
CY0Yi93LMEYaUyZD55boH4p5ZyEawTBIbhuD+Av/0L8Pv45DKjJyjHtWNXJbZ5C6
VdJMWoffRECgFH2Vj0Ds7+gzYT0xr4YaLwMhCQuBf99WHiq+CuaTvs0VfqAXkdBh
GYX4agqJBscSsKkx37Qf1+q4thhy/5tPWGYNoR9rP5MIUVCbcQpHZTVFTDF+DIc/
UMXS+636V+ER9XxaybuGken+t2OQU8o/kzU1HOCpzPw9PIDUtWbwdfbt62pn7JU3
Yrywj6DZx+2j4XwgYKg2jny+ExuUYaEjibZ4yTeu1WjqcqirEx6xXzL77vnYl+WB
hBkslQptqwGAqMXBC/vO/Ap3bDKLLPYEe9detV+z1FpJk+8DNXPzoFsmR6L9ls3S
FjiIQWJF6j+h2YeoW0DSYMSoYIcTx6Inqn2WowOcm6S1yuF553sj59iYPVzyL8DN
HvHw/8Orn7Cj+HE+Q9PdsDcEfaYo1HwlF6gRcChTkBPYR9xhafGwmr7ZMa35toIl
ARhP/uyBYyRdb68/EPYxJL/wD+LriQ5ywHMbU6FYHWtIThlDcDVAX/MMvli3Ewgh
8Xg4pO5Hg7AQzZHyzC0TEYqlPo1HmiojZvnLe3qgD65g5ydnh80AKmWyuuxTY52Z
sqYELxl9bx479OU0v80HhzGYc/SJXutZk1KniO1E8J8YQNJgKoimUij0IEPdH0DC
NzRI+rwoT7cArjMR/SSfMrHubBL9N4A8RkjAccQ9jPEmKwvpH+/YUXYnQNlMAINc
+Y5UGmSbDmYLPeQzBPsfvQK+818i8uG6Eqlg1Rc2+/qJakPs1OVg9CQsd30OlbHd
gsAZvY9vCYBZoFCq2NUMamh0HoSEI3hvIlXKv3mg8TuiIgTA+KEy3Sa5So2nMrJi
mTy336d1wDwkKzwx35G8YNc1Q92nIfAxWkeRX48CHDZ9MIp/3Pm7ZSF+nyR9HOiW
i62b4laYhlWx1pNagSyjSaTyEZER+lk7aD7mtF7by9yuO9BF1X21ajxUR5fu/KIi
pRTY/dyfrlrucjNu8qH7pcrNojVs4nYGeoHWCO2wD5C8/fhvgnSb228C3A1X09vw
rsWg/xmDWo/6KmGbVKZ8+ufCy/3XeMq86+gc+CdX/ekxFPz9Loz+Qw5V9B7DVF2l
KojoLQi0SsBjg7CCq57cuduA2lwgxnhOHWFfTCorCRKMzN/ZC4PUWuKcJ5WYkj3f
O9imF0/CoFBA3PnoqssvgMEjA691v5mjbkHe23D+s12lr6LMl1qCcMPvD0T6vXls
+PCXstE2unLZk6Y12ETHJqIqLJ/sxcOJ0+UMGLJqZeJtQSN/Sb+73LZ2AJX/EX4E
9D5gQC4yB6aot4jeMpb4DO3F51Kik/VxaXLBj4WtzL7F6XmHjDEtBR70cSgWhVNp
riTmUh+rK6BDi9rKvSifmbZOVvA3oQZLBmgL5qrgY6yNmfdc5NloGTouj1LVT51g
8++OLE9y2sblVCjyYXHPQG5waNa+XTJQeYlk5yCwKwQU5Gmwhw/1b+XTGCAE7bkr
K0/Pf6HV9+v1pjTZi5NXhcR4yQZmjLSi0ruYeu+i2v8ES2AATr3PfXkgp/PaSCh4
EcIfJQ3kWwydTqseihFfaJIZXcu3FjZanV5t4WH6WX0REp1oZqu69jHL/18XpTSE
x7cySPDRda6YmXaspM8Ll4T/JYU8DxmYOlYCiaVBXqlEq3rsLj1DHF++VAUrX3Qt
yMzAWaDPK3t1ilRbZ9gAzRtNsAKk6DTRtKmwRqHe/8ZFsPd1wq6FAPKMrPKNex94
jwT88/lX72iP8KisPjNBIrC6i5C4BPwHI3GoopnYMhPXZ+3nGPsbE8bLl2MehcAm
tG4yCXInACsaj9bob1YzfiEa/8oRSMq1nyoBsmicxwoO9ZoDYYeHgLpWf27Kj57R
QB5n3r1qwESGTxaVaizRH8xNWf2XEECJ/PZJNibMIKJOTFpX5Zeo/h0/PWqvvhji
xOUUWm90gXa+o3oK9BO74OktTcz+S02PvUkwoK1iUzJ7mCl1LrrW1rF/C9aYBjYY
TUdvj9d5HCjEvXPt1w74oeeIju+iUKfSv7DzJOLVCKRawIuVIt3mHAyheS30Jedh
kOjjqH2yGh059x5/3NCNsSkxhGr12EC7O0AjcGKzD5F26/fmjBLr0agFd2adn1P4
QmQLtskAF4p9C2LtQS/i50PxlDr3GhgUQreJBGybHA/4NKMat6QBUuMN/jgc5glM
ZS6kMPXxh8D6t5DgLbOqMD8GpOY33TkOeHxW8BqLiormYOgz/VtyfuIQJA8yELIe
V/Y2EUk7UqyIA/cpL47SG/E4sVCKRE5ciT2wrQu8yi7r2iGZlIJhLvPXOAoBds7/
00h1Mc8pnxyQjrstO/NRHY30AoCz5n++SWQdoD+ly/51QwNE1LeUR1vXfkNxCX1Z
Io2npHKb7Hspl7i78ukQ1E0/YsV23r9R2AB/8HGCDXRjaUgfdKe/4B+24OkcK7Ij
IhH6VPt8EEj1nl4Z8zBBrQK7ea9/cLtgNHywBlmitT3jpliWJQzAiwNzxY1Bn/eq
37xIiE+U46L4wTbubexJxIw0AwXQfYusIpeIUTpUR9cRlnt9RqQLzNjnyj1o9KPR
2V8kFhbieHAX0b6+uVyycROzN6ECf/EbqB3ARm0J8fXm5AXyOJ0sVbmFnNEHgIzc
YZJjt/tEl86YtIw6SA/2Jhi0kek9uL/VxOg46dlZLnAQ42m5m+QxYAPe/yltg4Jj
4ZungGAu/aKK8+rmZpAPhlRi8ILTnujxtMX304ako2Wcia+Bf1OLVBOK3AeoLdH/
JCqlpZQkCADlP4GMHR8UoGw6KaeUr+63/kePo7S+uHFaVHo19wjnpalkEUHUISM5
aNunnvbju+xEGNkYdaw3zWVdoJpJPkWhUc3Jb3MB4DRBaXKeDO8IhL/kAvHd6Qla
akwc7hLD9PU5X46X8wlLxJYT7VzvO3pA40Czwslzfyzh9pjqSYWdkixlE50seOt1
ClpvhlrOU0lc3whX6+LShCk5QA2h04DDvseeYSqmflGmYnx1o3ptNQB9RwjnGi9Q
jvEELcx5UFEepJ4kIs6A5xpRQwyrviSN9xvSFwenxFB8AWdWjvlFuvWD9Dl7vRkl
EmurA93usGFcvB4rmZVfKyoyt9MYRJKcJ0sY7v6KK4EInt58BdLYbrP/073w+EgX
XXoRpAFU9PDd+6r+UcWVZHsnlFMDmg/6skzng8KAQ7yzTOtpzI/DfKec55AjO/Ao
3kM3FUmGgqVzbSxtEhKCffCzQUxs/sfTVfDvIeoOswZwxbKfQzZeHW8Y2zeQkZUn
3mfwZI8JrYf5HOPo06ml+hyUpi9ynHJ3cwYJBy7Nkg2IdC/Drre02aJ731qRd/pt
Gw4e0FhCc+Eq/2T6EBxPGZqdMNjvv0zxAcneM1kO3Dv3aB0TaGCSJ9Zp1BBHhahl
GOAOC1LTNGVfbf3l1DL1laCBgDa2gp7RQkK8irrmOcFKu8VVVN5doeRki/sxynfU
/cfkvkEoY73VgsYm+DWgayk3l7QJrKVv0gqHkbWgxpAyYiC4dRwsv56bwn0QumhG
yLPUZ0+Tn8dS+jt3PLMMWRDjK0t95EptFZ8EL3hVlqhgVxQChGUws/9OdUS5RUau
N97ubED5kX1YavU3g1O4PiR0Mj/ts2aUb+YHrT8Xe0SHlsj5qwxLKCSl68AIWddC
VEYS1E1w3XiRdsRyayRWxQsQ8BKz/a5+7M6l5VjeFXwIi4dzn+mwc63HezSY9VUu
qOugu2sMsIDv9X+6eu1Ge+Igwc6Ezc4gY+Ag/iKlE284OERnZs+zIgKvm6t35s3W
xZIEhxxkE7nlwK2jQVhEd+Dld2G1n5tyFwV4KtGO9Chl6a/JV2eF02w2M5iSxRiW
tD9qgAQ+WJNN4jUuussaA3BoDEKmrO23AyE5U+/65Nt7NwpBVyxITDrOspFiuMg6
CcsLSxvWVqnWOgZ6yTQ1lX1zlufGTDgcwZ1G0qEP8nAJsRJYXaxtwxFGKLjo/9bK
7LljgRK7WwP2PLzhPSQzwl/1n+gaI6KNoeZZho9sOcerGbD+7aCQkVBRm722QiOI
hn2P3k1KYwIuClW0ZHqvG6nt6zctiR4yyEAHqAz+tvL0Ji/zQDYAF+ofFu3v4N0J
bJNx/jjiqwLHTOF+07bfOsoeRIicU1XgytRn2/u62d6nP4U59ZCigOw+FdhjBEa9
QoeurYltTVNMVG4kMl4WQmITdmuAr0qzqr28aoAg0sIYdHhEd4AaZ0jfq1+7St9o
n/HPZ/p4wVavcbYp08B4hh+4LdtBC7gzbAZnsSAqMntyWHKH6NpQW4XR/X/JDBWd
EwijswgmjfaeQ3G12Ke2RGMKi94uUB/awqDmhXY2GKYqgClrw3g2cuOPHgk4sP6I
aNpv5Mw1X06lv6r4+qyReaDsvayCgP2hR8LFWIKXRR9BzBr7GBDU/G2us2T9eCc5
VLzU1y1vvnQyn7nMxPEIDCLdHC5t08qpKcs6Jcxu0/EAMRpW6eFpxIXnsiU73062
KPblA5uth7BpVXz8NMx6uNfbWwC4wugWOfJhQot6n9Giq/XIvjL2lcfGl0Oq04vW
YsFlmQE8A8Qz1DfC3aL/7NfWMM+jAlONHvt8iNeNPbMOMRDRtWWTiT+7/jNoGN/4
vWSI8Bi12APo30YNKXSCL0FLk3Ky+cKQzihRbBRpC7JXgf/aV188ei+5iS+hAEiM
lQNinaaOOwpZ5Dcy6PnHdjxeMscYePFSEN+mkvhQYfZC4il07y5ZwVNfvyu5woBB
Kmij+8G3VoAXzZG779CUuQUkHNh+1nL0bIB/tzZhiiPC9kRyGGms6m1cGtvhet0z
275/RotRyLB/OhnJCpB8KR1HSFoWbmTs5Lpuzpyg1wEtr1r/XulJPOw1P+cnMWj+
MdOePqCZXvWBHNOn2krMIPW1gJxaqtyJIp0d3GYkQkUExH/08NMv85oNuElvt/bu
o8qgRdNb7fKRBOaOXFAd+7wXDjFA93QlQWBEokEJVS4RyZKvGKSJIzgNNJb+rH34
pRUv/mebv1Clp0rYtgTPA9yJjZ78aq03d21iO/iWGZQmuF4HwAW8IIrQHIe2oAwb
kSKB4nXmLW2057K5bI/Z29LuB7+GzSIqVFGf5AO67DKhxZVRWei5ZQPbj/dyW6F3
QgXGvrZd/e3cyhN8twNUflnA/Q/2jxD3ZEmJkqYknu1KvqwLsQ4MTTWyTU248enG
G2PeQi4RDGM/vUjoWKxGFczQLXOYBlLKJmWVMpvyX4PoXGFOu3OhzYYetG68ctCX
iF+uwVmXJhrROtlamBkKOk5oZD+XHIlqo0VRWPhGrv1bCsPWInTWoM9toF8b8/vY
6ShB3tdopHegi7HcCtontM/mZ2Ieso+RjaVZ2PLH1W6LYCT4pKtjMiyHQ2U3i+ku
UnMCDWvKASyDqNVU3F/R2b0VkeVb69wxItEWsuzdfCqfkCeVDa97EDaop8u68zC3
YC9IKLfVduXOJ8lqvHp9NGVwnUZx1KkEnpBR6h8FWxY+1qln8CbXOcIpzlmX2UQm
f4EmlKiHPWhpynHSOIYV7reYwHQoeLmuMFhHrw+hR1EW6mKywG1id7n5VodVypw5
BBgUixGMY5W0oingapMFYCiNTo3zYUx5o21Wt6Llm9/FlenN3V7Kg0Mqp6vhY0fM
t/Wc8RmStiUNvDXbXE/3qncZin0JSRTEDpB5TJSD85eOSxq6dCZNH/rSAOzJAxqU
5jvduslKgrKsRyd6W69h0OWz6CaLZJ5OHzxxzDZytvT3oDPCTC/Jl/N/QxNG5hVx
obeBDxAZN77Rjc5m/3UJ8F5rDCnnWExzd49iE4P1kioQuSotZim3br6nyKS5Ds2N
Mk3hR42w/yFzbyuUBeegYMY7THcti3bmOtJQfwAobw2RC4KbdwqdtAmRaEG+9YUV
FrnQHzpefDHelL0pzGcCcEEECv7avtFzc1G9/NLF+t/S1asPSG40g72o5L4LbLrv
pAqmW/RL19DWmRE491xdtHLuznKpH6EoESP63M1p2fJ46Z65ykB/+GI3VQBb2Xzo
dnLC2CzZDvmyPdNUctzSTP7y5SKgFKbY9b6llWLl4u6xAqDfEPIrYTzfCeTBJy5R
eEtdFTPNApaGe8oo3R6M4S2MWuKzmDWtWuk2iElk7F2DpsTQZl6oiwxby03KKoKT
pqO/25TQTu0DnukrJ9mdciVRyT28qJE9GGU+b2ECA4KVh1jGBNJLFQUdAGwDq0af
gJRySpglogfrOxZeIrH5ZUCj/jYWzuG2zTnLhQK9gqPjjqgU5ezC7TrrqcX4NxBR
IzzktxRAzOEvETNpgF9fPz/x406clIqfRWvgNxxUAGD+8wDlc2LGyLlWd29Rlyun
MDLnVzdVAhHeC27xxKh90Gafc8zF54xRfeM8jfUmgf6kzGHvn+90S+hC8Yj/0BhF
fLGxfrN9GV533sKqzF1b9Dd48kIdnFzn785HkA3/TpWRnuN8G8794eF+enEfVj03
0Xo2cOZ3PMPLZgz2KlRUUTeHDHeQmxEsKzvPkIKR2tYBrGPXS36EhMxjKwadJQJg
+L0lP8tX5dh3Qw4Brx586g3Xxq+Nad8aDJWan1A9F4cYIvzmA91M/LdsyQK5mxEd
0HdcnAbqFl+TsjuxESWy9bqjXSc8+fFUOmXZU8PfSXM0fBkO/C4qCAavMoWPJ62s
/iRqfipT89cpQXICQpAPI8yTSQiqDmgMA34zxjG56kAiR/S1HorsHA/pMj8Jindr
nTowOiwtFjn39IYb/m3trs8RxBYlo0I+GtLKD32jmWVZRCKNIJqAZUoZ/LrzGwS2
Jdv/N58Ajmuls3hL6t+j8/MKRHen0Bl6BzqqCNAnRTSf0hg1dnsonia24rXnRR0h
6jE4HcLoZvFk/m0BODVsfkB8pd/+L0C1+KKDoSLqh4Bt0wJW8ecmCJoS99tykmQW
BZnzu9Y7+riJ6Wk1RpIMy6vRk4zOn8BWLzZs/mPBqEcXH++csrilGU+Eai/KE43Q
dh3U4kIScNaiDFKtMbJD95lVo8SplWEXoPKF5hj8veIhyJizgg8+8sS0WfnaWaoF
yLahRVOy0m5AlTHgVNiCG0YjDY3RssBQlnOwLAksCduNzGQXAPBdWtJrf4129J+n
OwO5QDFtZZQK7WY5skv/NVl23DOM6VW2W9E1of0D6CVzYqXSmaZPYO33SW7iChqH
0Iiyp+/7B3fSZDLTtW0DuGMSmKivyLE13EY6ktLb5/E7KOCGHQP/EwNcmDYXyfLP
SPCCkGpdt57N2Ay9uc35n4l/OSG/rzWmYFXceMmIDHX34PyKufvQBc0VPDw+8kUE
k3pxia7FKo/cgqfrYMwXzz01Y4qmyGpIx0yXWhL+PHgzjzy1cpI1FlJaZZjiPwlN
hg7f3+VihAndMtGOMcMDiCcUp6cvGJ2dEddvgUShwmKxREWjaTTuODkR9vTAjrbr
bi6hTDCxZ7wrTQfpkcjFFks33OOmtHoSeXnF1UDTn1ijVS8Jhc55ALOim/M/z7sx
xhBH4c5Wk/e9bg+duTLKVAQhKN5yFhmUA4koRlnDR5wITwekXRJE8vxgpsk8f3Xm
LtNrc9f16KB7DCjfQAV8ZUsf2AtRUdgw4IFDj5mvMX5sm7uFeT2ADDBCHIJgZyHl
BNrzyBsQ92gHTCtQ2rohmI6yDnWgOOia7UorhHdNykLvmpJX3Hw+vF1qI/8u+Lcu
b0jdyaVrNOfdw1IzNlpCUPzLkyXFRJLriUnuHKGUbmXFuX6JICWjStPh1bTBkEt8
5CcIPZLdHXOA3vgjbDX+6cTks3VNFi5x0p3bE5P9EtOANA4LHjFZj4YSLHmrdkuT
BogEwDCXQCTKX6Qy2Uj9YSbn0O4vwmbzNd2fY++B++qHN2wG+kWEwrRd8KDFj0jD
d+2NJQChMDLmYAHAY/kqRt5hsyNyEHgKJL5YskqAsLXCu9C9NI5yf7hQbE0WnOr0
5OY7MgZjxgT4ZulO9nnJ7OaA5vqv88BMM5Npc6dYf/vLsHlbXvnn3LP3GJnHN+aV
VvH1Z0v4qbYcNaU9qVTLRa4wJh9WULhUESKTUKh0cXeQ78RPRsWUUhjrL4cgPy54
gVOhQJ36dV+qCHMkhDes47Hj6nnnCuq4vuNho22cNkyv88FGDfVG+IOQKk4UvMt6
qOa1wLNHRuSVPP1rzT2tiqZg89X7PKdxgk2PwxSgN5xzsMQp4SAcrQVuexyfBXsg
IYvlD1hG66GcKy7Y6ZqYXSU6d0kY41L1K2PFjxIyxFUvS/d1cZ88Tzs1FOSj/9s3
9qTBBt03jXWromGxkYkH+poR0d4RTSqLXl3PBXwSmF+1tcncExUX4qnXj2MSTUiL
V2qj4r93OhYeHIiZ70qQeIRCb4vwqZwvKczClu+xfxWxTtXj1tEOhz+tojIl1Oda
NlsKHEvHZN0n7plDtVA/MTC0PtUfuiUMfh4y9a2M0Bnm9izDE56TxL030pL+QsQ/
Lk0lpy+DAR+jAcmjtFnxdalNRr5tB1Gl7CryqStO+CNNImF9UYdN42hM52GS49g2
NmnaBU4HADd/dctzTe/G/9H/M+KNCGH5n8hjqRxDNqnPxIhg3eE4dM8BqV/P4Xue
UlVNv8GhEwe6PWoOo6rneqAFZ+W74AaOPR/TS5OfGBw+jw5SwQHwgWM4z9PQt8kg
QXv8rXa84vTwyBTknxqioWtKrUSslIED3lKEH/3tnWnNwNTYqjfNXtYwSVQwXfgg
QsQhYZMCsQwykQuiStL9BPwYE9ZHJPrlzvP0zGe7YOF0lEC9wh3u6MfCUjDOH854
aUZd1bQJFqQZmgyASxniLgUPL+L9yLkma/ai0/gdtKbvNWoU0l3tlNhInFKbrLz/
eN+rFDzcqngTA7qZbCYXqcSD1ZNTJaQCfUtPjhws/AmNLA2fh5GRpN1lcZ3UaY+a
UP1beJaJuIf8AvmV+TapbHO1F4vlYUNG/BNOv3ZKY8sjTiSgMB8C5GLKcoZU4LwA
QkRsSRBBygSuU5q1reNIkS6BvSfdy1iQXxhF5sqGpvLuSbGAthR2SUIQCbB0x0N4
Xvg+HIUzn8tLLF3JfLHv3UtQn7KJFskrOM9Ey6yQ2pIWyuxJQvVIPzCsA4d3eRfH
gM/3WptjtD0S7Mi3+SQEXSyapuNGtH54ZVxlZqgMOHj/7iWOb/jnY2/ruZXxgqdo
rO6BTs9YikZGylgH5U+MPJ6loHy4gMvrrV1jXCq4UJbXETYgFAbxuZF8iS73mYym
a/cJ6/pQkS+YzGoqUkKowAe5TpGvdtclSSRZln28LLIIXNmVO+0rYCFM8Vdm4vQ/
FybuWwyAhlC1q9+p1xEp1XHEwmmPq75y7Sch2F7u8gbjcI0P9AXcW9co2iqV2WDi
AMNmE5KSU6pG5n61VntUaNyuBc2iWuanl4t78PdCorC/9EIkffpIr/berlEAqm/y
DFcCTxOuuCd2UFTV4N3+xB4pzPlwJIJiftqQvm0TQ7wAaryaaszybHLd1+posCbV
RW0vcxdlsbBlxrZ+OFRQiT6ABVh98T3UTpuME6LUwqY4JKoSXM2jfNeqbJicWJz9
ybtCQggRDoQT8YwdSYd793ag/J2HDiCEvQg4LZxE2bHfbJzeKedco3FC12TdBKTh
EhocvaLkn20ZyEHH/3zzVhMv8EDqoKskshhYOgiOeeHrxyYM/AFDsUUIDXe1Cr7s
zDPLvvN9gV7Zte0Zeb0uM4gapidDzh0CjyhU7cfVMPPZiCPr8txXecyvgPnrbJdD
cm1Uue5ocvfz9Bhr6GB7YE7U9hzR6GzOTvmpCTYKja8nx+0TtV6YtFpZmEd7nJ4i
/+Zmuu2LRYuQHskDOSlv9L1bgkFqs/0QznYnQwivDW4WM0ci7D1Vg8xyrI3txM+i
wzdwFPO7C+231sPcSI+ZKN6cBVfrfygJYWdLYZwXym9tKsgk1v/YJYirvNVCyKus
yXe7bYfx88uG/rcRsyX5/TuwLIpy1C9ku9qFZjF3Kf6EZxxrYkMKd0H7xBMCY4lS
LnNxuKVfDXyPE6dEXwyqMVOHmBlXY4IlOzihTSys0daUzUFaczDyuvgzis3zdZRF
m39cJNMI03S/ciBOQ75eFn46Q0gUwpV0Bcc002SopUMS3wppqZtLffBQVZZvRAKF
R/wLS4bo2bWiVzX9Ldwa2Vls10FcT059Xj89GtVM7TbpAqpg5IvrFf/uSTfipVZd
3CP5TYF1uNsTW5Gb/mAiUqo38oju5wxgzYhAj47th3OG9EK7bkrfKtVhQjDFLR90
FxNX2ePrbAWfpvM9l7L4ZOrivCq96sVJw/CAmfyQM1bWJNVNF7xB0YTpnp89btNC
P78UT4hCUOeR/QDABr5BUs9lX0thmUcad6pk8ERsRxFljrrVsbvb562d6h3tNT12
+cy40//mUWzO5+VZ66twAgRa+RkAyDf3bAjW6xFiLvdWWEwq2fsDoaXnPVXVunNo
iciKmlu52Oyi4diJxWhVmNpPf4E/Ota10c7wUA3Ats18Iw669ttcBNXQcGMJES+w
DRLNtIXouoiNqXZaMB52hh1Y7andVdxTJk9XdcSzm/fbfRYpWfR7l/BidEu2xZ5s
3Av2F3v8qDSPnhsoQiLXFh4WJWOyrwCRqCJHOoTyuygPagpZ86qVfBIAx1QDFcg2
Z712RUZWWDEkwg6z79fQtFZ6+e3EE+RDTMlJT9IaEv2jbD8SX/8UMXYoCHNA3u1k
zcQjtsrP3mriv8IAXElWqaJhpP33rbCBN+NNvmL/3ys2uMnWbuwKxbiB55nykHyo
a5/i/OsKRjy3AKvjixKJbe89mWY3syebD8i9KgIRuKuluvfa4JUMHXLq4DPmUcM7
ooAC3TZhWc9Eegi9XLZRX5l6BWWRil+LZ27a+ts1516G1urKATomatrQsgYGFoNe
BW2s/bKLbQFed8T91e5Zli+6kOS2MgedoFbJPXXgg8qIFNv7Cz5htsKweeCJvB2i
iDZOBCRe9TYt3HsfT1ra52kRLh5eAslMQul4iZuebhuAH4D51qSF5se19XEUmXfI
XM9a3rpUxQwWUXa7bi+Dt3Q3pNHf3QOUWY6IFq3NB796AShdGiE0LPjAYYgRgO2x
tWlO59E3Y0crRZFPDQAUDC8JMMT24+HnM4romz4aY0IQZ1qQP8VxsqmXXmvmQ5pS
YcIBFH5qN3+mlctKyxVrPTuHc1IRhTH8YkVQdQMi+9yipqmf7F/Uwg9jSkY5/oVS
4ynei1SMvPcna/E4zGVKDRxPfTxai5ZobycIlh9Tq5x8+KXOZyPR6q208I8MUGA4
OZOLIEsJCtMkwiN/RvCsS/Edr3S6vQ68vkj7lVUtaBbjKoKlw1C0c/hvDEvswdm9
Irkge3DZxrAqV388ynDymlR/bG6HU10g0ARaNKMDy7lKghlsC1rcUWQUBvs06BTs
oCF9MdCjph6MPPDafvJ8v3HVlvWyf9WxJXuxE3xDvYXT2pIS+1S9TNqQGcBywI8i
JNPSPyRVO67BywdXN7L8MejXwvaT+/tJaTpv2sQWr9u9G7zdbu1H1WrEq/RhnSEC
cOZ0JvjMxQslhhuAK8m7ka1Ca5BOgtZl6hf4NJFQASHgQXvL5oRX0SUm4jPDB6f+
27vrAJUS56R0ikx0KEy9y5zZzvRAMXEBFnf6fN5y5VK1USNNHVFf0L4LftMLdpvR
MVHFwLnD5GRDDRnDqk7Wvz+YSNEMwWGgvfwBlr885tKBbXL5M5OCQ/Bhvn6CQX5i
/bv73mndyxz94EbK9s3T+qRQP2YlkEUVKXoT97Jn7OItwKf8UAQeBYH26K6MM7O9
++kVO2NwmnQa+cLsMm1b4wt+e4JAnGIyM7isYAXBu6yaq0jEW8/qkBkWFc3UEmlV
sZLu0NQ5KWV8SZDTYxt39R6rOfGuAqZa3m36D4xZFyydR1KGYa05yJtFwXuuctIK
K6md88mhLldXa51D5BwHMevXwe20PdPQ+FFFaEH1dORYoSVeaF1yWDN36roFFNEl
s/ZrVEUYaQkXEZ9GLSsAJwYuOP3B4C2D6uMHLeC4OA5MxqWoeyRkU5nShTAaKxTc
RzIhkS0X/MkVWAxRMWEMDR0zhRMWQiZCIHAZUARZYLbJYr68l5E2jRr8B/daXdOu
gtu9zfvJNhF7l/ejoahTj9JtlcHI8hpdogF4ZgmpnF7MFr+3dRzaajgNtROqWU9l
qKHpInbquuiH7x9onu+Nc+j9Dt4d50XZtkY4PVFvtbzhs9d2KQTGehIbchkDSP42
NUaPLOil7x+TwNJa/2PXjYNscOK9Xa0eORvJ0tUXP6xKzA5pBTJWhcf2nbXT4TzG
FCyRrzwCdfx57m13UGhGCKi8DnkIP8bMH/3Z3qXSG6G396G9h5bO41Facj7DE2K/
VsI5scT3TmMGiXSbbjGrWJ+UMFzNRSuLq79wkiXLQpgXTlVOeRRJMNU3pVl08qTJ
iqJTGjv3gxC28TdTB5W4Z8q1qVFLaXIHM/67WTOo8ySsHS7r8+B+CGtArGUrD/qV
VlD45gYmFeK5g0uHu7Tcdm+cxGbTMPWmMzzq0uJ/itffiFufVjN6GvI56Cn6Odlx
zaBWmMcb7UVUeOEnMuew5FeRNbLzKl29MqUrjQUsQGM9xnUYLF0xs6sbkxlq2O8E
GJGPdHKsA8HF9Sqou/RxzDzMWInb8ku6SfHIEFDU3AMTMX51YPmGE5kEVXHCxv0G
l09YPNa7JyFXc7TNnXj9O7KZgEkezxHCG7Pmqr0yXeG1rPE3FQmIr9QwMN9S581z
AIXbW6YR3xbsRGeKhme4PKik28zwDut10NsRPoe4HfgAJZtz141irRal8xK06F1L
k49B3vF2TfUfoIlrU3CpXeggtdBOYtBFjqgo3zufdNZtrs0c84i9K42oOIGZwqlN
OdNGZpU7vDk4EUWiMOhTrWTAszPie4MIqtcnccTYYDlie0w4U35mqluK+YusunvF
eFu/m2llEF1cE97z1MDq7H1uS/cL6cDmN4Rw9UD6kJgRUpmrQ0j89Pa+rvPpAlOA
7teQDkA6DIB9rqcLPOFBqfrbaPutNy4HDie0TzzjeXoMd/VfDbLSLt88FwoJD9hz
oUk/NjBYOXKnDRUP606imC9sh2Z5uCiS94ohOg0iuOhIW3efJsOcfFjKPG/BatbH
OmZV6WOR8Kdc0OYJ26+mqtvUJV9a6LorxMcgAnTrvGvGHx+1QcqyTJms/uxp6tZN
/SwdICRszBYgGN05d5en8nfU5rDBSrjy4L9lUSyFvLz//EXCy8R2KuZ9lKPFbgal
lMIy5FKlcbAdijOgmrdGiOtYW4e1Z2H6GHQEJNQFPvIsSH8QXKLaFJoB/Jke0lJG
5zwkMTpsFANqza1+lV95F5qK23z8fDKZdCzLDGfacHR1Z1LjaGfi1KdXEaeMMErq
EZtCp3ptj7BIoOvoRiM1CbQM+fvqzyM6ctLo12mtz199o/nllG/IZuGcd6/blY7V
UO4FvwbvqBMEApkFXs2YoGCQjcAfnOA27ORJPE3UdCT3ZosSdaM2xTarJrOhoUAG
qwmdGFaP6f9H6pDOUiW5QWpBfjlN9zyDwZc61IKj5xtjC1aF4W6Xy4rFVO8BGjc0
JBgTkI8WgYS0Pue678j5lBZ0jA7F/JL0KRwXhlnc7RQ6m3ZUomY5pPjMuAteMrw2
BMjcZLMrNkVHEs0XcJN0pLLHMLIX8hlHjEwRyLiKeoWT5ciD15ENqHZ8bx8tpeft
+NZHjy3qJ8VAwAcAKZb5fR6L46gEITSAkUrjoHCnX1fiZA4qVkw2yXY0i7JPs7OQ
VU2VyLBKga5RZAwInzDqJQZMga9KpH1vFDz6kEC+AHdjRCzooXi60g5ZmhrKVxoW
r6GWOA7sNmFcBTo3QmG/oZiGv0xARaJGfuuKRJYWQ1X12b5ZFR0XZTrFtdAir412
ozbQ2iPWyz0pGY3LvE1x8LGe1y5ucQsz94jB3JJQ3p0s5F7vfqMOp/qjS37iQZOH
5US2upYtr4v7U01bfm3AXUetrwlSBNMrnZu/LusxRRMtVuIOri4KfniIZOZTHTL/
mdpY0GsZL7KLZHw+B6D8KccLTm7C4/YZLhDIIsx7Q8ILOIhyC7k5EA8NhClXT1YS
aDj324xsGpxtJ5JxVVuE/3Hvt2AVgGZ2UFK1oswOzU2dnu/KxlyobIDxl7QdLjIF
UgDaEJb6f+ZsPOIjMySNpK05esvWaEXMT0gAlyIXTU3AR37dyrB37M9ft5l+PBlt
5nG1H6FzlhuQ8K6mHG9aFe9jFBQTbpmpKs33gzAfmtsy/MO78we3YN8XTdX1U4W8
O5abvBDiFP0SY1Y8wjyib1T/aS4Wyuw9yuxCXNiZWu0OI9Z/TG0jjD6cPb4vFEAO
hnJUy5+fgNPykIg8lfEtifZ9cAxL1hwLn/sc57f7mSI8ecKR5QVsEYypVw1qGWRX
Lu7CtH+6kikC5+Cmsf+6gOOQbyMwmsg4cSyDbkQXS6low/effB32XmhevhpcnCCY
8iiO603hibED3bXwoP6b6XLmnh0rX3jsb6f0Nwdekwhy1dtsC56qV+U+CEuoxaBx
vSsUDoCYNJ54hOmkiSMKDRF07BLsQeahqbwdLG+NP+uh1uN/w6bMMXMfAgGgcc0U
78DxlJdnZoeORAjBs2OCGmx0cSXBzXroUo3ng1je3ukZwp8xbnVIy1crsZs9QWHL
N8LrxIxuPcpiyYSwMgsoBvKYbTsZRyghG2wj76raKVpcnLWx3hz1Zlcf2o6gXBYg
tGRXeMiv+FycbZZGLMcpD9v57C3FKRD83DdHPhllLGzCLYgWLoDs7/9rgPEm8bZf
Ikzi4/4WE2UYEqjWWPmPaf32ZZ3K4IgVjoyHCwWkz5AdfiCesJ31qj8FZFyc9Lwb
ePbpsjUUE24Yqpe8gCP5mUUvtiA73Ut4KDzVLlkNfhAuu82keQmV9UMZgkXw8JgQ
8wGIXRPeBUqhh/lIFYVHBDD7oC/mS5ijzuE84kn+bPiQf19P72zLpvnHPMi9Tv6P
QKMNejYdSpT6RSLhX2DYxf3lX0fsZ3jw7uqRB9i2GrzFvZMHe2/NP5Wx0EvFhATg
O30JYdu+d8dY1XUlE8Vw9oX69nMAPemNtT7Fko8spEGNGEq7J8bsAl/tJBWLrwLu
MM0DNAK4qfoXQgfrUI/P5U73KxgM9a1wXpDy53StwOfsNiD3GJeNdxFXa0xLASfB
hfn7YN1CUzzrjhVJckPBkDwEGYGtaWsYdxN6AlHGsWaXwmrAHY/4Iam8tRJ8eYi9
Uz8XnUTxvtA3dBd6fIbv1TaA+hQSIzlszOUqD94TT5pCH2bussCnAElBNTBrva9S
jh7++AC5P3dMOsUxlgJ/QUbY8KZkzoUcGN6uN4VjpkEf1A84xSxlWHbPaitV8ThV
tK2ne9TWaQkUZkiOqO/Vc7w3D/tNs5NZvHZfBdLIov87TJYMOD3bXDlwebc1Ozvs
Sgy1ypsjp5gl8TGe21BTk14q7yOhhTTBiTbxauIQs4r2X4nU5tsJ1v4t9ymqQ3H9
4wGTWf3eAEiXzJJVPRov9RtNs0Eo/fvgk1FsEZXKk1laHj4pF//p8Pl9QFAm5O2L
vC9g3m+ZVwYHAA8oGKmUAm6IV7aaEF/fBb/fc9gjejrzLB+kiz7NBeu0G9tCk+A9
7GpJgH/SFLwkkDd0++ttiuLKLaW6ZSyDFFyAaI5ThoBAxmYC0BF52UzzXvC5uL9s
ocwCgyUQ64/98FsGpxXHVw2f0q7gXWg0sxvRYGevW+ksy8QpCRqWEOmPCJBlUM/B
Pn+WzRWaAUu4MN9r1CUirRiWdgBZTcP7LYNCjw39IP/vRt/03DMYCYlWS666EMVV
MRpaVmnoGzoPsFs4Bhm4OdDr338ccVMgeWZPFtwkDQVaFQtOOJjHBvhG0DaRk5j+
SSZ5jhphRmcpfv6Ea7im3jRaYs/sbNedZ+Eq14JAfpTdSL+t1pflKlpovEwHE8UU
KKchcj0iQpQ1w6r2vzRCKb5NZaPhKdMwZiR+rXsF5/X/cGwDjKonl91H5A/N6F+0
+2lnRPSsm/KO0X25ZP3NL5/PzfD9TdhPZdv18jZXOO0zzdSHWz1PJlESIEpHAS3O
U+xpvEX6IGFEe+FPBqxE6Eu4dlly/dV9CBrCRlILgBQHklr19e/3sUSMc9E9BDNC
Xs4+Nn1bTenDILEEK6jIAAtLUqwRAUDfHAJ/k9NYlsQ6BTbyDHGnkDv+D1fklvg5
Eh2nw84sF/BphlpG+kQLIw7vq22O3lkHb5plx3ZjYvbqVtMXukzcgclzmL/G1Qoz
+WWLHNXvoxImjj6F7+LPxNljun5cpDueEflLvsupGiI/YiYQh4OJfh2MjZ9nuSpj
J21fTV2vXCjFsPeW0ZKPD0PQkXKZOAYzaLc6PwUxj9Vqzcrppd4Y849bzR84kxFt
VS/UTEpx58h17fNOmcww2eX7anpM4MAZ6PRI55QgngqYoKERyS9nKtppmiDSdNOf
jrphxNpe1j9jJ3rUKr7zeRQq8oSuFeMxH+5GUS4JOsuFNURHr6/SUZksZKEd5kTc
n467bkrU0XmxMV2W6trBv0eOdh6l8REOaC2s234+Mtwr42AKsrPz+On4B2pWyQv9
ppopRKkwrgwVtGeZiqp/cOSs/8rHqM68zyHeUcxlgJDl4vo/TJ/D7/4IivTEMbTa
6q59s70Ljw25cirALc3GAYVLQFS3wiNQMDjkxjwuvfis+/tDAEAYBnlhXx1SBFUJ
ZCSfub5ZtG+e+Cv9hQ8qqbXNTEDCjurUU3KytaVBRUDO/vPDVuTEnhzjAcTRByxY
EAuqhmp+9rKToquLiL0NA7LRvnhOgJA+UWytjASlqQA/1WulCHAVL1Ws2H9qL/Y+
lALd0SLSGALTzS2B6H8HJc0zMFOUvQde2hx78gymEks3b3EEl96G2prxtUhs3eDB
kzl6zIbIfu17TmfDXq1NScFVtoXpOd23V4x2wilwQkQZvSFmtDKr/g3Sk8BX+byn
eas1u3MNx5ebZH2OxaSx8QWXucP1NgnWixz6F5oZ5ZvndiGTzwKfc5gwPMBQQcKD
rxi0Ivh3eMoCOH6GHhwy3bZQ5Xx5s9EIRmsV3wexwkBlMDJ3F2qqf4/CGUhLxtm6
/8kzWDMXQRzJK2P5Ly23DkzsTecBmdd72KJzvHdh0DXmo2HUGN/Bq6v2C69H61KW
/FyeqP/8TKbt4VboipPEDEu2PWc15J8dYaxI2q1CYeVQ7obwVUt6vZZhl3UCEsQa
PAA21iawarKp94/UOynyQenz9CEq84fMNE9NqiAaaQCmG2mM0JNjwwvTQN1h0hgm
ZNwPZVouyTUhnIrYeX/JuMCMYRW/cgRsErnLvDCgqyN+Z8WGnbufcWIZyn51B6yD
tY71tgWpQDmu6ZRfVS2uN5e0GN+ZpPG4YUc4uUxwUdFs1BJgi5ThSLr14NDqd9he
zcXWi3C6Y7+l2sLqaoMBRgmZfT8lxLn5RzArV4xxObguyjmQ6IOzjbYWCI18hfwc
sUDgspuVxFjEyVfI860EDEYuRwAZbMv39lngc5rR3lbL6mzyvDjHEdp928uZXnn6
tBDke8m+48nOB0x+7CIlXmml8qjyWsWZeTtUmmUrFKralj+TTvl1CuCedY2nx2pO
sKI6ODNAKtf1JVZbphP528ylqy0+RNmOZFrFX1UQpYyLG70C/b+RtTMqdX6hMqyj
DakHTmBqnm2LvEtHtm/boilGSL7kWw2fTNGL2/XO/XobTghvgm743ta5O+ACSG0y
r+rcbfoHSnsGigKI2w3OVdk4TWztAkImFFG4c34R0FGAFfpEFfK8//N1RVjIa1AT
yT6npyMHKbVfTpncmI0YhW27w1ZhLNpBxdrIX8LQSCXcDn6cAaZCEcXSWnWqPpqP
A+zmzbBnDdksiATfgvwTaS8pCn4McNGooTC0fRn5GPfmCWRxm6BNGAoAaG25JkUt
HM5zhcUOC648YsRgw43r56PVUAxXLy1iBa1k1naPRK+gqL+KsQcwMoMPx54DmT3a
ABWdhtzUg3OLtY9e6FLtqyskVInMKOilKmxwNqv1KZ5ra1cozkLd7XOzwXMQjk5c
qlarGi8w7pgUvQMCgEaIyiXufECaxfkGhNTNJWg0SIk+HTq3Mq4Bks5wO2Mv8qZC
lmvZbv+2riMMt55kmOdINGDNzajeazQgPIFe9Gl8If7TnxtOqsFbQHnl0mKLiUtd
QNIOn5R3jJ0bQ7XFHAdXzMLSAgAt+jyfS9ziKVNfPZtblYR8jzz9WB0E5hZUFSQL
j2cEeKFWFAeZgE45Bc/wwK3a8bHXStXLXOFAaeO1wrJ0jG5neGOC5UcbaVVml3yO
DQZKrfSMSmHKCsFbthG6gLELNgyYQQ0sjGr3EEoKs+SWDaWghe2Pz2PaFAww4ucz
/ocZ7oy+6MUrFPPXEWbnIWVwsCFHhtfJtnLOx9th1TNkjSddnM63RZqSLMsoUtSI
a8F540nzWihqYSGQsXkBmyv7nVAjSBDdMB0xMIlVv+jKo2pKKEQXqr1XiXtgtrTM
fVOrQaPecdoDEc6whJ6Ef/TIKaQlLEY0DRMf2hjtsaO1jiv9l30dZAn55F5GzgGf
f+hweN7fS+tbZ7ZesvTDcHBtpRb4ypnSA0aBAVa26on8jtK0fjqFliuejj3M73Tk
C5VGC1RGCUrq+Gs5b8W85xJkzh+MqIbUTjisO9CiXEmaFzrbYyWe9NHA97nxUd5b
x4pMxpJOboORtVtO4+0RBHvi6r9w1NwFnHx0iZOD3NsbpY2lrUf4yC6bjTeqvd37
Gw1t5cmLxqJusgEakPgFIDA7HFKGQNxfTE59WfRmj0gsp1EE7xj9XENS/NBg2ozc
KjyQtSDCA3m4/pvVKb3uLcYK4HqHjaNvF5xQQKZvW8hjSjIDTAFwCLbfgjEoMsm0
5iFzLXkNsctsf4OdQORxNO13V28dcy1zhGezS9gaaYp/R1xGvf3WzwcXh5O7QcJx
iR7Q4adnCOR9ILdLcBc16qRtiI0dZ7uL6DZURE5lE32YK4ID9/iYAd5+QByb2RAy
BlL+Wm574e/MPOX8/IzR8/55C4kXCroVlHQagbYRIWRcob6HwNSKJPOAR8LTFrXU
Aa7hnSEEOwwYzBzDVEiyUVxblbWdszVQRblfwxdWeHg9udH3ENsrelY3ugrh1gi7
KBFqhnuKbgpaU9MBZwp7XkuXUSn+gGjHV9xpDofQz29ZIR0ovUR7EU61x6UUZ7Oh
GCJ1ZDiJlsGlkkF/sgGrLvxMhL66oe6qM6QREnXyuhFdtEmAyO58VjPUkYz35ZRP
D2mTl/+Qu1pyrwBk5Nyy6PmxM0S4relweS1v358x1hevvJTv3h0XztLSME/GEJSF
QpamhDzagZW/OGbXmD/zvlYwlqrUnIBUpnn0DY6faVkXcZPxwMzXfaxY6AN3YR2g
nwJH7npfmypUY6xKgnehXVCX6xAy2QWpM/6L9I5cfj5KvkgRzW9UGfhQEcbxmUa9
faEkVW0SlzztQ8SG2tY46iWPqZfQ/04EX7HDWX3PqofPGzzlLGwLPwxchHmZMHEW
4BVGgsLKndPr/BOU+haEXCJAPyFKm+3C6nGF2rWbZXkbEojaTB+jy8kYAwVrRg8f
cqRXsUr6l1VAmnpNoCVQJirC43WfuRGtwpnmgGAGPaDeWLTaeyhuwtxZGTwnGhba
kFdAjQjOhJZR99fqZjFXowIMlH0KVStb1Lxap1Rj28tYBl7xDSiFVT/4lpW662DK
30pYvZG6iKv4caVaJSyv5Zpx2bHkKGjZRtUpEQXz7TXRm4hQzPmusmJDp2I6zIFD
VIRRrNU3lvs0ewFxvUnFo87Nmfxd26y++JrstI79n05ajL4lYcbUZw+d5uQ2Ot2C
yujOcZRswBB4me93OXefwYfGy2mPZlV3qZ6ZEKhvCOCbCU/a2bl9rvGsp+2qPosU
v5n+15GZudZhwN8edWB2VljVhpckjiSKXcezLzeXC2CFTaINyEl//As96tqLesP+
PqK+WcgsD2Cz5xz45l7SfV+xnBmkEYv6AVVI6uZaemSilYkVIMW8zZjPr8SWJAzx
uCkGx79pwFjaMWhLTb1n2B9BPGarr3dNcDKsIrw0wI8EAJoKM95P9VNBPF/RQ4eC
H3kFOmYM5kzB5xgmCHXrvAxA8tp63q9N9/ti5DFCH+yrKi9PtWS1QH+e/atNSRzv
XzRFTpaUn9yS2PMWCFJ1GGiiVVJQPv+mrODGnXxBs2oqZBdRCHnezhoKHrPAsiUV
VO6Z+2LhxLSoh89ulmj9hCdWb4r8nNiyhO2TwlCcdw1fJp3mu8JLk2KDz+RaHQaw
xdyQ52FWr+cusGv+q6EcHPXxOqZlmWrYQ6NoiTB5OwFs4/SycJsZjuh5Ituphb3G
IUNoG6UAc1Cidw62uCy+sE6YvuUHia2fr7/fzqrClihVLsDGtCYQ6PBLPOdG7XZo
0kwbjjGoaCmsY9VJ7kCbysgEK5YOCb1/VxGxY8K1ln9AUkBWRhiXPWrOqFIYm4S9
4ujAh4ihYyn5HUX4cZhy3gn52olJA8+cYtYXUNohuyH/fRA1D4Zx+dVSxAkOodSF
PUrqtSnntIMJUqNup0Inn4IrvhIPt14YfEXrld2KKL/QeHefY7inSaQ38t56qUcl
Ao5iVgYPLmDH5tw2B4xZVXwVrbFedfTZBjLObENXhJfwL+MdE9SIMqd+cTAHQhMS
xX/ymC9rvobB9eCJnS3afIcOgnu7bLeRkGQp4e992ame1Qj4dMhfHjv3jhd2Xjem
fGQ5MTvJgESwnodglY6scI6ysBGrJg8czooIEHvhvPkVdEa2v9beyatHm6hxjIRs
gyitluq3hHD/iQH4Bvf0hIBKsMyZ5C3RW6SvZrH8lX3V6h05nOsUDSYJUkm7OUgk
YKve1+GnhyEQ3jliBLtvtsHiVR3WCuj3HzIbuluqafIoffW92lmW9wJRhTS03ZaK
4aFzC4i5LvSTA2Wl0S9FCvbQalYJyoxVt2FfZGzvtEQSmLMzFHyB0603XQ2HZju9
QSQIO8X82eFqT8rJXkILa/3w0L6CcI7689Leg1jMHn1VsmkF6jpkQI/cmYZJye3l
OosvH3Ml12Ebtt25TnTmRx4wyR8S+kFh6gXbkLOOncVcPgxRGNMnGncUuJSJrJXU
cqNoSBpUjOSqKKHkZEa2bu0dQjX9cA3tD5Rh+L00JNPZOT8HuQz97ocNn82lCnF5
9DSGqVrlFaxOJPYU80EJ8d2yaMEQbNtIulFNW5IR3pE/l8oMcF32PhCPcvFzyyxK
CV5ybY9kdv1tzmQ6lvf2IDE4W3fFmhA8khRo62GGylIdr6QqawWk2BAOSZ+bceKk
ULGh0tCoVfTDi1Lq4SGwQ+eBMN3tWX7wapqumXMipaFbuQGwS/TKABJtUJ3lEXO1
FX8UAqmGHQeEEnTctyL13RXvlPzsANmWp7N17VMIbTO73KVd13bOpuegVlHCBaQS
7tk4aZUC4vgAMvwzU1aWMNcBjcMtUT7mzNpL58LjKQGPP5AM4aQqgK4WLwzPOva5
AVJ+Uo5Maa56ogAkfDLpDsvd6eixJ1UdZyD1o9u6AxqRjWh/p/3wON8in5VM/z+C
ncGV3cp9mKepuLcIbPq38bVY3731SR6dByc0M4KUlm21E1V7Wqt+2bs1Byr0dCrw
lMHqPRlowStXWlT+8X1uYGTMeLFWSoaWCTE4Lp6nHiGSzoH+kHmpzDOhHo44fDPd
NILQbEJRMlOM6BYcLZcapgbQROJRXKZYF/y5vCGJ4ug11EgBoOlWoIACNBwPP+6y
maDAynAO1mTQVhfY2H78fhiJaoX6SgMQAQ0+VOIqurJ7er2rlQ0r7LeCGYAog6q7
+OSJZnmtW4mJxAdEaOVldq39Kjrw/MBkEbu1ZYhR9iniBmqO31WARgCqxMw1prmq
gAlBIzHtykaUDyQMz0zKRCSNZBP6OF7PrNfOMySLxSZpZJSK0goFTeg2DyDcHEOe
AAs1Agp45d93W7w/7bboSHQciAiB9z6InZrOj1x66G+el/9Nucv9lDjJV2ghjIpY
GD9Tv+0+1z1NbEWcrqh5KMSvokMvG85ngjnMwOg8QCUA5Tk28FtX0FG34V9qT3/3
UwEb+C5gF6JVaF1f+hKxuDpp4lIT+sEBaNThS52C9KPuNthIbqQW//E7pHWBCOkd
FM7lWtDUAIYJFEcZhm7LG2rQjRU+Cc/vXJYpnmbSD91iTgFKJHWAvJ5mZ5ZCii3T
BtUnDLucikdPQrJV/loZV1XAHjwZF/l1V03TsFNfmW4g6Ob0tUaIXB1dkJHD1wlP
9NLaqA4cKqIs7oQou+npCm57hrKSe+/IGiDfOqO8pCN9PsTegABJG+jL4mnsxsh3
39iPjor0ECNU0O5lIVs6nr2e3ONFEPKtX6B9LHQy5BNlPXEY76Wk+ZmHDx36sXyf
e9oRGGqsotHDmYO8CJNyjWq54Vak58ZX3+/t7MKXrRnDfxeUp/PX7rirk4Mz9It5
G1+SMPIbLPkXRhzJ1uTjCilOM/x3/8C44Dvn78FOJ9Ja1BBesSY636uX2N0pWH8u
JJzHEfOwUSgbbBSa2KAhzvZgXCZa8YGbgVHfcoFaJtnMJVyw+LmX2K5KNFvUA9G+
UQdsv4wQTcmyi/bV0ASLPqy7xeFUTkNjphXQoSIUb1dPZUM+2aRy5fkhvBNh0gM2
BDsCv4bUnFYTwW6mPlgMZiczAm/DSlpzoLc6xBFMlNAOJs4IeikcRHOXxkUkRSmp
5DngXmD5hMKymLRp02gLYEybhjuODPhO2XkhC3cOmXrspbEFaCxANqhYMeKs5KDH
EnTTvKgWTZnNXnm6MHBYMrNbTft6OYHDTO1PevCWZMs9C7657Q90UIwbIwuI6dKU
XpIuBW7wnjAk1WY/4iHVypZb39FBC00enpY/i5i2FTNvGf2hWQK3BXC+SZUVvHXH
F8YOZTd2AO98rMCxZUDqeIPemJypbMb7NfQzp7LMdrLdEVSPAo//NFGaZPK10w9J
KXZBIMBWYCMy/xXIRGMbY2Hx94u6x+qx217tbLko0SkSI1GNMOi30tezjWcgI2FW
c+bR36CyvqhCl9PpQxQMAoCXiA/8MqeBCeOTOqo+3jTZ7bHy8s5C6eJ7oHLO/KLW
pt6TYwidO4+5g9NNeVNYZEepP++47X9ZnG97xohJXLvqnmVmHMPj+H8V3dcxsm0T
fNORRxuP43j3m6F4Ik0r6vvlG2o8CTew7FQIrmY8nmz1gPPnrF4WaiiBgfk8nZDj
rE6GfBdLA7WhHvqNfBUbmmPfRalNgod8JV1QG9TwXknuNq3jDKICcmGl2T+7bANN
MTKL2y+q75lMamKaqbYEWjt6xS14kHMh1sqE500UpxZ7vWMnw9LohlekIqYlGn2b
nVIxcYzCCgeGS+D+ksoAizvA6je1vhD5mtODSfn6ie4V49RlSp70y/or8Iv4AisR
BXVGnYStUW9YonAbFg5ViEgWZIk6piStRvXuFjUtldoP/gXHC8fwi5gvyubLyzgg
BPDfRuSgtXLIWa2RYR+4Y+IML0kHeqGR4mYQ/YXj0kVQPkS5cRPTjtKpJtbHttV/
fg1RtsSnYhWS7PRsq9V1q8lSS//n5ey2G5qwJwdxZn/R5Cak5SPDoVvrQQevX+ro
b2q/VRRV5y/8bzsyvhz4CXIHZIRC+TF0+gFooFwDeGVOrnLZWMYEqumR1l0YGx1n
kmPi9k+1lO4RhKdpf6c7dbCULF7VMD+qJFloMXmKSG77y/F8BmGXYxnZJw2sBHZJ
1NO/unJbAy6dJdVcWh1Q/1MmxxEAYafyjSXaht5QkSEOWAuwkPlwzvTz4SWokEx/
QP0MiyB9bfjufLrbAvvVGz5cJpI35/AnlVWtZ12Pc0mplB688fhEyOSERNFtYXxM
r542YVafYUAYawoAacpPN0ZGTYiiHgLD1khwy6WW5qK1PM5lAv2VdqtXJv7z7B24
Hwm5MBaNSb5/RdODxkgwSlaOsNDmJWZDDIkjGfg/NuPkYzw/T3RIfq78Xij9hXPX
kNkaWMh2WhM94leg5OIDIpDqKRq0ew24gXovPtq6J6TNOmXC2YOsM3AZHeNmahwZ
gUodBA83DoVTF4UoB7V31PTPOAiofnnd5wxj/8UXPpZriB7bjLWmoK/pUI6FgTT/
LckD+G6Opg29YQ7eN20AqvKBvrS3DeoBBKS+KnJ5wPrP3HhwDpDZqyuTunXbf5Wt
ySI32xU9yW5mUZ9X+cpP+hkkKH+nHBXvzmDjS+WVwiBTSO77u6lrx2etAaEtAye4
6YEwHbYzEP0CTnEEACT6n4FHlJ8eBfvA2ZU8UuFXntAlz3uqOfSk7/KicnbW1uCC
Gfqt8stdJBWvchbUMQtgMd5B3YyVE3Czt9erwzpkdjVhOJuRjVHb60B0k96d9X6c
ziVCzJAQ3GJ9gG3fEL22e5iNv1je2RHi+I23TWDHPbG6bo1KSrTtc0dle3qqLrmU
rZCAFhCYtq1BrQRwwQ0hetz74UfQ8tJ4LxY4u98vsJHx9SLAuyBLmijoGkxL7zIT
0+AC54he63Ow7+i+nDh245MkBy1AUU861nwBcaO1qz+fDOusmGJUbTF6GuPwEBkZ
N+bkfIDRQ3EwrhwRQ3L/Q24T/R9ouruAjLHDB00S5GabMRfiaa3fm4mSHpVnKxiq
gZQE49KrTIZ6OA5QRP3K52tAsL6vefHc+I6qYH//cHHy1nW0ms0F4scjN5IMbXIE
zZS7iTCL/SCD/877vgAMpDyoT2B2ozpGs2qR6f3E7hZ3bS+s90CtuAMZ4ucH6E0x
SGkGGdi16kawVs/7gl1lMXBvwi0SHbCTTmCYKTxfdnaH7bb7llhMj5ShLpCYZyPp
PX40+k1BH9QVFMkBDz9lnGrtkjEevPRsJXC6bQNf8/pzuOJzwhTDR2w+poa7d3Av
gXPEHnZjlQUtZvIfT8gJJcLuW6BTqLl6TivJDyccmuBBBkFFXlan5iIIS8bkIweh
PA8Mqxw+vk95/V6JYpsDXH/M5ARmFrGk7i1LTpg3/vdQ978yfrxamz7TgzwmOTHF
S+Apqu0zt6zyPMy6h3v3MP6otQ7PWuOxIywgX3b4QlrASp+979ibao2J5Ty67K9Y
rtW+QuSpJG8R5vaNNZ+1M1uaUud3WrZzFt5BYNRrb0gHjFCPPObopY/g1i5VtLWG
Y/DEkOZQDlEe2jtE+SmuRaxsPSuu4G3a+Bj+oiGLbhFMIhsGekHfZCw7NGwQ6jL0
8EWu64UBbbHQlE73A7PPFqHp+XK/7ZJTnCiXk4OMiAstE3JZ3ug0O3961GKH46ef
keO37wpkcUc00qB1H0gzFj1HTvNclcWjEs9MndyE0iSqg88na2AJn8/TVzQiLY8Y
C6dxgNw2OAnPS2z/8N+M7Omv+A4Kl54let5KMGCR5m7z3evbtTsGn7tUpgR4cRqA
2Ts3QtAIignXgi+RQyiu1JIJF69XO+38v5Esvgc8vT7oX4NbDOddGmVXBJurzz+M
c8FdwWWDpmRmNb28F0eL/2vqS8MCwMrj2gIP+rxQx/JyVhBEj2u52lgZbtdJCqx8
9lfeVE5QqhD8jIxEgLBT19yk6u3+3i40fTPbUJ7vGm9RDL5ty5Z1JaGEaR+Efg9u
VYv72hgZwwQnxBV4Tuf9EQEp+sqL/gKCjJSZ5QqmUhKmbL9bcJbgYqV0xilBAKRp
8XMrsPCTznNsTdH/sFgp3L9dHowkiUz1uA7G2CTN6rRkfZcVa205DUHWTxFIT92Y
xItktRfOsrAsWNQSUxKatQYZ4Cvb1bZajvrA7ccFzXNvA0xFQIl2rP9h1cDgC+ux
iydGNWU0RZ4koq282nVlGp57pTCrQAsR0ZLz3zXDqIcNff8td/roFAXWLn1Yb1Ei
qGD4sK+WW1rB3e4TkxnhHjCWYBWkMAoXMRPILdybAPPL+7CrkljMp4z9gv+RMane
7gEYhIllTNHnEkemXUYnpnshfs0xoXt2azyEAo7EPf67poB0zDncJSgKDNx1SYeK
PcLbThNAIqLnvAFjK7++y3BGdATa3zZUzOk9GqK5qgD0o3+OX3vUafLX7BkHNuQ9
GXyfUvEopcIzO5vA/9oY810vm6OcPRN36QHkTJrImpUvUup3FD4fo9vn/9D/3dic
OmHHKh1rTf9n7V9CJom4b0XGdXtVK90c/Juk+TmVVIAIIEcL2RvmFjwg2m4+JTGM
SSF6UZwO5CSSaT9Cgrd6j6x/YLd/AUr3zPndRwDMKJfL7VAX6OkkZ4SuaDgXU7gY
OGB/lHK92np2aRtLEaBhZNyiGGXH/YSbqPPnHC+wC35ixmU1bscomR/MqsdLEgld
HPPOB07ABL/fqOrkwErRxXRFnu+bheKQUb5HZ9gKSqWHvIO376Hs3DoATEPjw3lw
tqYlrxYkZ1JsQdLC7o9b2dG5hpUlGLigrAzZYownGBOpFIChjkBWQ+en2x47fVBA
pv1TlbzRmRyay7DelW5Wc4/BWAmmwYDm+//6yP0T9Skgoy9Ck/RsdieUXy8g6xuc
taX2N6rx599kO7a3KFh6enymo3hde+YwrvvPIh68AcHuomjaf28vR0Wdzp05yzpl
mniqwNEYrYYriSDWD6Jbj14HLKzc6K2dyhDiJmMkejEiJEROh9gBgukyzuBzS8T4
8THekIqM8TQH/fd8uJwTn4JljZ6p1tOnzTjtKhloYMea4Jg/I9X5h/1exvKDuCDr
4rHL+AOpnKeUUy4X9zlUW5RHJRWB+iHrriwDOWzcxs05gfCPJiyMgZHv5d/KDYgr
r2XUml1tcLnj4VcoeSlv81hW1Z6gndDgMq6DMF0GzWM6XiwE0OpXF2h3LLAk9FBT
FtugxSH8wdvc6ku01llF/6c5uAlWyQxoDSuCeZ3s50Ba4UJZ/DXBqkzsPs2esvuD
+WhnczkAlhHI3vSClzaVrBaBhZ7QP6q3WdBKm8AHGyE9a6JDllSR35MJZqrZPJy4
UJ/JtL4N6kvDSYwFmoTUqgMDJNKcye8KqYCRXfszWfO5KdTPZrjr9McslAbu+F63
dFgMSkRtZGNuPNuPoDiGo4VKe6jv3Zg3yAMCS/roi0RCJSAWzTQcAl3LeNyx097P
lAe9f26awemcQy8Nbuu8c9B3HFLJXAg5areLweC5Rvu2aWy1bHkYcTwOmZKrGd5y
eAlqoorHviBhcAVatBcb/NRUHzQk/WsXxba3L7aOs4UUAwbo9QilVoWZkXMC1LGk
LYlU77+2vK+/MLjyt/ZyOnvoaX5AXSxHZCt1U7dtI/GkUhQB9nQSlx+IbCnHfB//
cmuD97vaaOo6m+LCodzwaXZc9Pon+IVVzipQvnaM1debh5BaVzMqRMKUG1OmW6WD
JaiggvE1fdpyRYR0wd4c52SzZVRtHKnKhOx+exWQV5O1ZyzteOY43Wg5NKJhr/9G
qctAz9Ih1SFPKttMxdmfppe5wJf7XJ6ZusGD/6Dn0tqHnEKMnU7FaEZ+F9ObfRAx
tPzOraCQtomicyVKAMAqvIeLDGWL9wXJs4FFI1A9BNIT/6bv/W2P6L3xfwrQwDWS
E7lxQvtbtZ0dr4BX6DuOLqZ3tZWrBDf0NQJZRKA9PRFoHBVq2x6lxVeLeoXowJQI
MYU8wd4S1mqB6YhcHcWhxC7wpeMI0+R1waR05BjBm52fAsbilkShdLNj8mxTuRvU
qbUGAtmWyjlQytoi6nQ6xcqhdFoA55vgZDntiTw6n1V6q3h4+GVqaWXRVWYqqYRs
OxUpQve0oB0okbL2uEvCBF0w66x73X6qpF55/sLErxLy9TF0RZbRIFMJpGxNVAO4
FPOfy5JrSYNXpeRU5D8E4JoBSbYZeasQzvAidWqsgHopzEKVry+/SpKgQ8Mnfhce
APjj9jQVe3vT4aDLrMjTkmdS44NFlcSw136fOiLSc7x4SsubveMcGPwKZGCcDoEZ
57NPLqItWfyPdtDHNzeuD3QG58mtdtQ3RAzoWuxx12hJBIBugPqnWiZi31oZH7di
CRR04WUsF7+lEmB/dBJlrGvpIdy1ogpPHNEpbdB/cPxZMYkP/iZoj98/bZRdMrJe
YY5LR0HfT+axCqjuvKvu7EbeNrEPc/neEjwVXFk5Dn4pkLi1vapcoZ2ZqogxnuGs
biXyX4OsKOhm2I6dw7bGsv7JW6Sc++/yGi7gkbrtqDF8t+N8DkWh7nbX3OmFHwOC
bpVv5cS4SwDMCXpg6ZFB7VCpWO5voPCreB0PpxGRnkxisvF64QbFjVaz1A1BPwzy
BXSJ9yEnkVx7KgDI0Gc/zFOBvdDENtudGLcDOIkhft7HQaT6WZLCxhb6NL0DVY+J
TXph4ETzbgBaWdT37Bx2UT4T2lMj8ebAK2MMSamOIpMFOX1naZfKLEIU+cT0yCzG
5ZNRkax46x0rQpgWlVDa3cQXiPJEAykpe2xLzINFSCItgwOkGyQlUDQWNx1eiABB
btY7A929YJfbInP5PbyPQsvDM+sK3egeDEyF1t8rDmSoap5wew6c1bXGNl1/sW2V
t2mngVqEJF4CgxBSJoPiRpbWvOe9C2RWeYJFhOCYkTT/rm+3rT0Up4SYL5s9QUGx
szhvU/BAs5vkH3aYBX1DVtQfZzg1N139KdJIM3JA/ds1OFgIvOwl6OHc794BTzoJ
FF9AnnjQ1KraWkOVzYi5duaHg0BsHokD//MbTqp66C4y1Rh78KmixffB2Pj4G/aO
YyOFeAZxXmFAac53e2/QrAypsLEJK8mFfRtUwphzTUXm9jDZrZt7O3g7Mhe2shZf
PeX58AB8v8lcnJkUTDsnCw239c/pDUCqi9maSAdtWcZNQyAjeskBeMD+k77LkgBr
EL7GZf2DY4/QLJHWz9toFH3dkIkL9PQPs2US7reZ/tmaKPdjjIqWukroMp/AIdqe
7/vJFQs+bMMqwagrHEl5bY8GiGWN20C7XJhdGi3JV8HG2Oqev4ycjLhgTDz5Gw9Z
UsgqEiO56M+6lgDwBWpYte34SZQ3NyykdR+2NTFXnL0BtHZrCgQP5J5dawefRmWn
hGHtV2+EzfknYhXNYhNfxny4DKgXoqrxPfj2Xx+sCWAG+pOqUT2UtUyJK7Snhu2i
1IJ9t1sW7eklRxOVg6EdinLj8GVzVp32MuhtBuwpP3FP/+7YJqNQeH134dKf0rV6
S1a8Yz+/wbhmKpD8tDJEIFCP9dygutAtkBkDB8AFE+EZp6HXgMHdfdt9C32ClMow
/EObqv1Lm11qKHZ/isPK3K39lZB8v44SG7n00tIAlIDAePNh94piUiUNCtVHAaCI
b5WRR4GhjvGBQf2AQc1Lbb6Fb9m0gf66uHcK0aLSu5/44KJWTcd6oWL+PIF8pzrA
oiCTMbNu9HbcKYyFJ2XajHPV79BgU+MuSUIlUgC8gRg9HYrTAKSm2T3uRollaGoo
5sGDAOEHZZKRFWOqIAnAxh54SPFkPrGhzCLDaalla2tFxbQunM16Vke7LBCfaxAu
M1XztvTh+D7EqINWBffw9vshqteg/np3qbANTZ1npYpeUk/fDOcOmnl9oOsXAwOi
iulYjvkVQhg9tRDmuky5ASFLhffNmSQkXWjm0d3DNWI7CnO7xxuE97xO+caEWHA2
u513rV6Jd4W6VLeo+wrOuqMeZ7VfMXvGB68MfJusTPwTg9epmOLkAz6Mv/A89lWf
1lNd8w3hAc27zZmqPR4qHzjPUQeVoDU1v/VXY/IiY4Mh8yWQbYPrIvpYa4BEBDM/
iLqh0dqCIlxyzZ6/YBkAl24gDKXBkmnSdfNFNAZwuKfCa2LB7OYmR1M1GQbmmevD
VG9s1a1LYB5YWvQLYdGxvY+hSdUBrKLTmI/whsuyWP7pXLXlNtbpiSuBfdCM0bEw
F5tMYezMln0DDroL1j2m/XjhySHVyOJX67d2XAIavmZnHuR8Zju53bqneNK86NSo
WLYELnH9fceg9gDloJXK2giXS3viwdcEvhGMLKz6l04S5yIuLSUn8wbk/Ab+/cf1
qU0rMtXhO2pC44kka3g59cTBWWQVmaIngJ6QoZajDka1p+sk5rsewpTKHhXo08Z6
MeZT35oopxkH5l4ifv7/7Gja9ucrmij4Fa7XVnxhGWeBLhZAij0iV5tqvxQPCjns
50an8aJEydfGHzyNrJvKbdneg8NI3OadFJqXYNRk4z3dnZVgL881mYGjrzdssn6+
U3t2/TWD0tXiSM2SeS8pnge9buc7xnwfA+T8wmftTDYt41zZxSccOLSCoPFQZh2v
Ym9WYbrHyPu6aCXQjvKRVdVZM94rM2R7KpLQuCHAm945zObE72UeUeCNvWcGPf67
jrMqc4kijtQPBzGbq+290JYhpIqHhz7Se/jRFx04YqsBVsr0WizwmmM6xAVwWbwu
fYSlajtTKBKL7l8RX3/B2p8iLXUMdKaALmgedDYgx9blSvWrskt/qYYgtqedxJN7
QfJadjYSzvtVkljtKOXK6rVoN37/XHm1/Pq6i0b4g0Aw9eLHi3EaIqD4nFvyMte8
/+anG9b4wrkM2Zu6TZzV4390duY9A9frUWZViE7VX4VXhiXtoN4JVVUaaaFzCABP
urVEPXQ+Ut+hefTI8YgsezTGcehDs5fE8b+AwjgjNcW4T2JUeEfhdIO3ADW6H460
G22I6gkzFis64vcR8wdyTsqZOrIvax2JAEstTL51U+CkqPBztronAZgS4JZ6wIQe
aIL1O+Ho5A2q1aqR8mBatCKlFNc0dL3qrrXGd7EGAW95zVlmWhArdGYVOSbq7Y+R
e+Wta5FQV6NH0O9VF4uPU8DBmvMpvvWMVW+jE0tiVW6b4iE1qzZfL8NmNLx0L8FQ
bhMtunWUIxyJ96T70ou0+0qM6erIEFs32ZpkOfW9NLuHdbeD1FPnt9b9e4iPuCxq
OSgZV+FI3MxvcMt/dC46luMCfJa2gndFlQ7jStFsKLiHLTCTLf/1zPRA3QZu0Yuv
/O5gOu3ou6MiChw3m17PXronTTlbQqnmLRyG9dwWeprmllTdHujSMyn3wUswLosN
K4ih7whCnj/M1YNhGY+wg3HweA3FJ0fW1hoK76XtUpTtY+kgV2TLfb0oOS/fnM8y
qila2AH2qYj/KZqshYYR3NIY0xSGUH1CoOOGBzttTzsDaweFIdK5asBHlei/3idG
eqecmQdoGDwESpPpCMJtp7BVgYCjbvWVyGOug1V5uODBhhootHDeaRsvTHLyJdGP
m38DLN/UeE7hse2NxdVkBuG3HwNU6wO3w8S5iUsQwncfVAGsCC/ITgAwfopga++c
LF2+dLdaRQmcTNoFobWwXzAvDwhCLavrn0pgEPHE6eLgWlySbxioC5Aja0l7R1VZ
PssBnk8PEigtTn/sJRNCWdV8QZ95eGgQ21XsQl9ITZLr8HUpjfUotHW28Sndu60S
o2VKdnPwk1+57+uMyDmiInYAFQPAWv64+7tGv+Neag1DUbpJjnsitX+83hDB5IX+
vdSPVsChiHCZiJiHhuSEN5PJFNt5AGcVRo6SpI8SM/lPMZjNo0NmUA3SqHtgOk14
0jHBTAr/vpFDx0YI3C9termii/DA7fxhHk16kq0tRA3PJK3L2YRyBmhcooZoUx8R
F/KNzq3o8jAImvmtqaSD1HPovaquevOFMzCoHPlfCy8I1h5QzyB4Iyl0Vpq1Dh0/
Sk+iTQDGS7a/rIzFr/itHL1UE40QYk3Z+RxAcnnePaaNYbzbGdZstvPeYwpGNATF
DuvfUyCfCnl2HOiqe2Q+d9Zkv1g+q1iZDzza7D4jnzdIQxPkD8MNWe0u0uZa595W
3I4vNF6PXRHDtrFf3h9kPd8cJxpCsDxbh4kTOa46Rubq8Z8Zhqi28psnyEAQJolA
3VpZjX2oqE60wa0LkFjDybrDZSIrfNIjRyPElx2bpk29PEYthkyyFXcpY3OZUc/U
PcijquxUcksu/hU4nFK/6hjH7gJLQ0NWC07AbUikuHRfpO1slOC+PC5mmu5j++d2
BMOpBRLOSZVkyRgtjETaJtibW0Qak7QHDHq5Z2Sn8OxUjt93iqwsUS92eMOJ7sS8
gw5MS1ToYG0QaS4fGvwsNfBQwQobHZlAjYkyPRXc0Hh5BEXjOv3HCCx6wRdrnTtx
MzCIeCMXXekubY0NO7xnrWyXBPW4jEWP+OcNjz73VXr5JDje3UAumHZbYn3H9VGB
WsHmy+dqbGjh0m88LAZQ1ZWScHka8NGVxlJCXjGFuknDAKWnCs36tfQ1NfbVtfHI
V+KM3XcsrWBfC/5mhfieylXZ7qxyb2Oi+4Q8pZJfREgm/V6qWEbRPhDhOgISmqf0
3oAYP7whLUR8kXytTRwcQo7ADDpimBsvA8M7U4y7uiPC5dRHjscyI4WxAjpfeS2v
rGxYWo2JrWS2XLNnWzFuK28YU59hmqn9ehap6XZnHxXytnnoVdfbqRODsMR6FZk9
uD2amuA3pfbmN4dXqYoWMst0x0qnUSm81Nsk/1ZZxr610Kr+bFtNWDDDrMusj48K
nZjTa83J2yS4j5KVZH+m1N5RxtoBpY34pLTHZLCMRMOvl4HTPOqB3M0kP73/m+zv
OmnXePMo6lYC5aaWPCfNqhQDT6s1lQF7r8BKMRWEWu6RcMRoQJbCV5dTbwpHzv+O
zqyf62OQhBzPO8TgOxvSkCf00BlsMDvnUm36LUJIHsTJvJhqUIGBq/sWLccPCw+U
C5NiDbVmw1rSZHLuJLisqU7g4r5DtNozo+u2uiZt3LqrCDhP8qUtqTcLNZFChBpG
VMo06mySHObeXsaO4+StRbbMC1U96OxR1P6RqG57bQmdIIQv29qvZgDzT1GLLRH5
Jwvfb+xM03FVYEig5aAO8Zdr97VqSojdnV3+mm/64LzRdcwWl+OBdjriSCkCxvY0
15enbusRKjfsn/8iF8Ns+soC5nfmPk1VxoAL7y3X+o/mMrTwU+3QRsY8OaeRPzA/
liY8wvmsatcDXHWSKN3ly2YsC0Y/htbfPDNR2UjpdanF1p3F6oPBHCLgQGwwd7TG
aPpJuW2pdVBpZMv0I/a9dqpVbepPSkKEfzF3FX71Awb+XW+2lFxCMJqVJTp+18lu
/nLcxw3T8TxrqbyEcokUdGft1t24ATc2qoL7VgGtp0jpYMzMd+kGcFSsf6IuZZNJ
3t/4PqPvSHfTfg+eCZji8aNnh4KJL3crAytVgyX2yP0frjUBCfMC8hBAxLnYWr4H
a9OvJ2wlSFi6NwRhXwetX35BCWvXvBdzyMeNarfcLSruCwj4KtUWlkgTXuV8rXSl
aNagI8upviJr4rieNMnFA208dT66H9vdgbjw/BybHvIg/HTLfX1hztb30eh9DTQY
y++iQT/S+YOhim+C7VsPa7EwBnjz8RJw7QRr2drBDXQLVItfrceVRq5ztWscP2mQ
XxfGtK+ToSmwEzrTl584Xkt6FadpkrHZ9avRCmWnLgI2FOBJfS5st1mHXK5DqFM5
MCXmbUDBpMBDy5P6WZaVohp8hMqkyjIY+VzYjVAa6Ti7elG3ca1rSHnaVBG4m0Gv
klDIYsQmoGZ3pbUD7pXcOUBsiczz3xgywg1KnVXdslNOOtuOwUvRH0cmDcK09ZQE
pw9ZIjTvHPFijC+O1jmzUBxnRjNQr60PwzZo+ZI7ah2EdbMRbtGOrEGEAnWWyheR
uQWT7/pPmbqBdu2K5sDeoiZM2QhvN2N8+oliGugccFoE1zcCYm+tObQ0gRl+vcTy
gMDzMPSO6Yy76k74UHofu68OEMwtgX7BF9EU1syNBmlY5Gsz27JyBl/D35fdaSx7
4vu03Upw7qwIWlvYsl5cGzxoLD1vRzZopWTPfU6DPzrkchA3tltxSw2VDcuhifEh
2Kyapgxtiy81AyoURZRz/Vy+X6QG37OX9MCc6bMWV5a1qDlxSBi0PfN2IrngkbUN
Oj+FKxHBdDTFbq4B1yc/atS8500z6VZTQKzm6FA0YxdvDN3AIk1P+O7liXvXwqDz
tZ7N8OFbxNIts7BegFcIulcwlEa8CKjX8ffF84iKiEx/tJ+cjigwt/2eVAjNaTZo
VDgeoan8FRjRW8I7E89hhSOkJz7c3CySAyFzpxy4c6dyCYXPIUtY7cBTNZCU7/c6
Rv0PNh0H/bHm+b0OB6ak+s61+83TStLidEjLPhJfQVmAw644WU1kNGCDVTFLhLkq
GcAdv1xGdcVM7DeJRRc+LZlZRIBqRZ1EOkMmbX6EviRukxaWBXAdPBbrrBsZ94w3
uv4Bmy/mrMIJh0/bd8x1kaO3FRlLB/6gQ8ZN6wC0fMWr/lzRsXypqM29AUFNIMLh
CzuosSKhx5J5cadepXeowYvc43hiu30GczvtHb3GXX/Q3hCSULTooJEVZHIhNMIs
zkrhmJnNHKmWLhuVal3VvBjmLpbuIjof47Wy+phJSad3X/yn+oJGhrSW0Lz+Q60U
xACMxG1AAVLyEMT4Y/3YolI2nOf15sHYiRSeTssFQC664rTyTZlAd5/mesZetWwA
9qlCCxVd9pwrbtYgiiXkF4MCQY3X0kv5ZOo5xvZq0ML0wSBrsQbgqXIn6nv+2yE4
TR0E5y6P1Vh8xXC/rkUv8+MdGEiCMIRO2qqbmKEnLySW+/lPLhUAqWHACM9xvarV
8gG6Xr0CtRJwUY5sVNZJtyk3kGu8TYzmy5H3EuzuTgu8k3zL5EmUQX/7ag/0wx1t
OdZPMgw0zxEpO5+nl3kY32kzfZsnWC52OvzfsoGXKOgxPVmKbu6bQH6hhdGUSOaG
gHuK0pNZtQ1jySUYiIvHUdDOKTPd4vE1nNVsVae2WsNFFHqNnfLcz8ZUEpAhNIaG
pYW6fCRxuLaHR+9bIFDaTnNFrZtfAMF6pBiqqLRZEpQWCbrlF/yiyhUto5P0zUJI
lyYIFvfmHmg3coRK0EenwIk+vz4sSYxqvkl9n3G/F+ia7PWe0Cm464G3DUtLBhUL
ogt9F0hn0oKwkezrR5btFFqHJc8ezp7JBlmnmCTGgGz7eJi5Et33+EKDNWomU/6C
YVFgP4Et4QEtm0A1exHnkLY2dxars5HpBx5rFmwo4CvMuXgirJLx3hn7d0hEtrrw
k86PeZivf7uScKcnrV9OfioWTk1UKG56Sm+6GZNp8Hkn3YaNr+3p78tVlKgZzk4O
Zo167LZqn3zGs++d8DWQy6c4ERnut2ZV7Lg6JQbr8k0wCyHeYxLG2xBfqIKDyW/2
ic/vWf1rwPqQCUSpNB+u6BG/jsyoNbhzfYPEZAyq3D2PyzeuCtHVwQIGRj6rANsa
9sG4QXAyQt1NifDfNMBmK5H4LBaV1nMhOrEAPo7uJW/Z3VWzOn0z19Iowqr9MERq
YpohGTGB54Vu/rBJajV0uOT8i4FeCAkruPvmJ140O2rl09SIg/zY6GYplc4A+XgH
Oa20gFQiXsiFF1B+jr31pg2xFsuLHhuEQ9iw6QTNNILR1SKQEdmnvOUCGB/LhhzG
RqnYo7XGaWt1TD4Fhnk+5Mo6WWoKGCYvRYEWarnJspB8DYOHY0QeXE2ZesQANYko
gE2iu3BbfV0zMzNm/4vCQqoGHU/PZx44Su0WDw5F+dY/NA4sBZpj2OMJ8nNtTLbs
B0iwdJ3Fbz0xKgpZHVb9md0vIIxN6y3g/N/FxQnNK092Q5gKJA4s2TDQ/ep8jXt+
5ZJ4r/hMn3fQ2o8WE8XbxdlY6Tuhz0c5wHnyLDGzytw6L5pP/ABzBSKToOJtLGnc
48VTr5yOQNjjSdtDd6z0Ba5bqCGidCO/LHpxz91n3JMIVdreLuAIL/aRSj5wx1MN
VvuRlljMH+01wqO3BNIXbEgHiMmGroRfBuTnx9txR78G2/n9XnT8YR2p0+WDcxrF
l4CBXoS465Hc1XANCZL7NR2QX845Z3coQ8WDSYP/xKLpf+gURqLvKnJ2MlRMsTLu
/r2HP9wrPjpZLmua4cs9ziBwJGUD3TKLI1RkBs2LofKY49uxAQ3JvDNqTFup7Gl3
fHVRRpsXjG6TUyqLSEZgPH9t306AmBiL8SgJm9a95y/dla68gjGqhRjYLsBEMRqy
wuCT6MWZ8zdp1ws1zpSL55PpDiQzz/g70tIxZzGCQJ/Vc1Rm2a9eG7TNj6QtSl5k
qFdNjJxtI2lT17b3ZdWShSecz959XSLfzPhlk1iomINhFYJe/pPyH0o779PCS5zj
j44ivlLG00S9FiZtJ6ykFGInqBvFByUnwQ0RilFWaP9RNKtOhLr1YMaYmI3PgP3A
NyTkO2/fZOYvq4HWyOqxEVv0nTeql8pXY2fDE80u2NHPrrkN+OOWjOS3J9BsXwUk
BMc3r79ByD1cBuci5Zmhpc1/otLcxYbk1mOR/N3alc/WJc3Uc12np1UKWAyLVWnr
/u2+5v6weLlZ2ateJBP1JWqrollUFY8Bslm36qJZVsoQ7oe2Z6SPzoOAb3gxTLVD
ZUEigTFXSdMIg7CUn0o2Lki+oc2CjBk4CLqMZHNdlNH69PXmXAtefQ1+yVlinDX/
vZnxsFbQ9N6T+cktI4CJFWxUELONpHwAF7ppCg9VmVscBDfp8kmDgqezT5P8mq1S
ZwitNhjPMfInkXqZwB/6O7zLtHivJZM/SJ9rPvDf+vvva6BhsgUXhP1OcacJ0Qsh
G0NgYMOZnzYebH9FzK7MnH2/SQ99Bra4W3xrTLp8nQs4xRtzC57qztZtITGuNF7l
Ht4xoS/fFuhk8k+zsQMdq8/x4d9l/CiEdjDjhW5vPRSLk6sn+PTVPNEd/FUeskAp
zxrCkRtwve7p2vm0L/deRyzTHXPx59niVj5a58TvyugNRwy5k/Lf5uXd+dMVUUNw
T6xlA++A1aUiojLZOjEsk63BA3un8n9OPjbIHUpo72WHHcyblVBf78X2m+6BUPPW
+KlFhnT2RJOSjtLRBY9WMBHQTSf8R/cI/OEf5NxvwwSZUPNcUrcV20Iy1czCl3mT
kI6OLhTFZPABJW0dw5TbtySb/2Imqn0UzIN2iupIqmaHLA+BDFBF0kzBXW+g9Y9x
KaRQpfNHl9IlxKVAMFnbGF9df3GyGcIyfjguLAARafuoVvG7ZueCLLgxEjmJWjgi
bRhQow6nS0SeUuXDLeKLQ2n1YKAu0kFugwxSZyWdEiK2bri8WB1ObvE1/xcBU6Dq
KvPtvITtrqWHXl4YFT5QXmH3FTWLPZyVBK0pmy+XqHxjh7LQAkQBfqPqUgyDoEpF
E9iICUKLODGaB/qLys8ue3JB09BXZRq+rj+WBHe6Uccye9TC00r0tx7geQwCrQBE
UsEkudguGKn8re6K+qE/1jGetFZmSUoOB6gtXnopRAEJ2TYf3kVjVZrwxkMlfOVp
s5KFZx1KVOkvCr6oIh70mRhoZi1KzC64nC1Jb7P3rRNcGmn0raIeKJESwUEx5fBO
6Jkf/DYy1PAAH0pzzrILisoEItXQOpnRJHczRwOJ+mPj79bbrtKqgVM2YdK27i0C
wxd5j6R1KA+IVGuuGzGmiE2Hpa8tihYGYU9vJBWRGKmtwVps3cbVpXVzuZ/MePdG
EEPllketmlhOqiH4M1698NDpxnUglPGCAnvxCftfbjAzAG2Dxr+orUSGsow8lBc8
nRgd0QbZnoHVNRpU1gpIX8b/gs7zazM+YT/ZG73DEouB1HKm4Lf4Gd2eFytKidgr
w1I8DsfE+yvPB3faAttGwBBMqFvcpdLu/L+eKBqvhPhMKpByApTScGGvpC/KXqNH
xjAbjO0I15o8isf67AoyiIKxOB+m6Zux17oO2XS2b/QdGgCuJvBNcIa46Z2QwsSB
B88jGK5GZGBslCZZcPUneF6JdZKw3fkNoO9Auk+1VKIQYter0P7ui92EdHnIvYwk
O1Gw9K99Kllb/E92TkOyBV6LZ15dmFvUh4YpblMtquoerqQPwPyhsKuyv+0JMBnX
kVblHQ+IAXL3Su9qT9b0OFofkmvQGkEbwfQc/SAehLw1VX+SGAc0XhFvSTzz8diK
F2sDT84Qix0f3cMmLWU2Kl5luI53hhnTwhUIwxeh7PZfWIRNL99ThSI0W+dKagQq
0ZjXTKLNe//V1K3tAGt9pw7ry34C44WEQPUpZb4HjxlxrwvTuEC3B7WdoxYAhmpB
iZu+zv7+P8PRMcQo8qyIwtePJ9l6G1n0y7uoZNjRs9GYCt+wPrRnlOMEgsdPyTPK
sqiITX3F7EZOdsr1v8m9aGiBU0RgBfEN9NmO8Mq+bFkPdeaFbBqB1NmWXdjQohcY
BoCBiGMx8nLjGujbhm+4mwRuSSghPb+33VIcOhMn09Kb5cARyk0JbeplH5fmh7gm
UDw+EUmZCY0aIfL7Bk2stkh3SQeHcoXLxw1zVdUCQ9D4NojE6f9PfEd+E+RKnst6
vYYHn2GPuD+Olcyt191fdy+noZSGdMSQwARe0FQq0bYM1075xlmXjn33mGVUpCs5
ceo28d7GRtzM1LUvNdzUtUQMcxGLnoN8dmKFOiwYUmHRkaxDoK3tonQXUr1266g6
tpjSU9VGDU3OdPDdIZCmX6VYGMyCtle+RGmUzOQ2PpbtY1JvvpnN+hPbZnwBzWLP
c+PstjHT+0KuRzDcks8Z/mSbeC4eb4PzBmddSQtComrLnYV3ytnQX1Xe4Tv4nI1d
kI34PLDuCDm2cvVDdXw9xLu2xkgjyKRO26X+3yl43qwhsbrrQ0WNp8CKJ6Dljpg+
mJWEtanPlGyC7AnrTxgwBkv5JsH7g6/7YO+mKxJZmzFLPxAh/tJoh2AYOi1CuddI
hsG70dainBHtGftb2ZiIDR8Lkzw6k7XysecNmQZPAD1Rh9bun5wgGke0LDeVEk86
aPCFovZw+w8ajSe20dYL+C/AJu1/jVTzXMdfCBdu9CST0UqR2+FeCh2GlArChuOv
EatwkV6sCsu/mjq4xG53hjQROHXtwVBxA2RywJXsvAsP/9fKdFtViT6vSGnkatqp
zv+aTI7j62Bpb3+1blbjqd2YTeN7k0wqEgqcUupohFH9WR3QaDGYLW6ykHyxArxe
nkI66wj9V9J3MCfRy8MdbELKOwDQ+NVf7j85KvwuO/Ans0VrEe6Nf4zQ0RdE6gxl
SqT0tXRtHZssDXBPURvoBkZpSVUUS0LxQwLPCXC9zuko/vihuQI+O1dlLm0jOjij
SRBBXQ05arq2MqoKYpQ2u5LdL+YKJZrDRMRFk1ln8gplqwr8IvG39qnjZp2FUlZD
N6GoXsZOEV1bgLxIvGrl9GYhNDP7xl3hhR3nHoSH0U/sS9p5dUrYWNu1vTccvDC6
jn69NT5kVqXEIroWHCkC2Q/SVR4YSodU7m1vv1VVaZpMcJpyk+0Y1g4oEn804a2b
DMMtsJbPf6uWdeVGGJYLRu/bS9TWPNjdJ8YLb01ycxY9coJauSTKh+e1+w/LewQ4
YqTXaP8bHcJeadR9fHYEZw075RT0rfH9mi2gt5Im4jj6Ce3tPPkAI+fN2fN/kbP9
te52E7Zw/MpvM4dEyiUVTHRYjd2m08tnFm5ksfBWoK8S189HTnoawf1e6ERFx+RJ
7Jzy0tid90aRR5yj1qLXog3emfGf0dlFblpkGR6yhuKwv6YcNcqdqirl+K+ErJol
pnEH5oaOKxM9mWMWmH6oC2Y7W7p0LQmxcgPGhTvLw/GuMPtdEnQY/pMnBOf6o23L
XYlzXmtZ109WWBYo7/UmFu2Ub2bdqIF+UwTr6hJn1u77Kqk4UcqA/lpl88Ygci3m
zVEIzrRKjVgi/4VhgiyJ2gabS8Ceual6OrFVxBjPzsCGb3x8NtY4kMRuV7CD0aFE
TcsjVEqiEGWmxsTnBjt56k7XNlqWU/oesy/r7VnVMA+5JIO0Xl5XCjiSZY5Erd+S
g5SQ0eooyMPjwniVp/k4d5jJPt0mOTdLpjq3M2ryZr8YRxTTQRhZirQhVJmGTmMi
KmJadI3TP5zE4ubhI8bz2D4Oi5s+mE8yWt3vaJeoKUtonkebs9QSSnEfRxV03sSW
H1574oXapD4rhvGJu+XSBFn0ZAesdkoPkKQ8Z8eZqtMZ0W6m+Cbv25tef3WE/usz
KMovDub0p1CiKvfgdQ0D1ovQj7yRgudyQuE9bhVVrtn+mjucxP0wAVvnlQdrSUXr
M8R1GIJajqvbE0Du1/8ojECpcxC0s6Le8+t5LO1N64ac2IUPda7ro7UeNTROq6P2
ol1p4xnm3WdJx6uCBGctv6oBpf+t1g1MN4vpB6+X68cVPrsF7XuxleFbj3sTbU1q
Sr7erwe5hiWPZYBt7lDWXQ9ucELAibjkiy8e/jEhIxQmxHLFvaUeyvKJz7RYrcSq
jJFc2IFt2dpPt+6lK9zwaGlNHkcqqVtvw72J0DEJrxkecz52oQaBn6aWprE5Smk/
j8Pq5UB5EaRyhBTPCl3h340blJbWwVbXqpudB5SG2seN0Pm6olm7RZowJOtMG8uC
LknuYIC4iBNklXeQaDY8KCQm3h5mV6HHO1oPAaYJnwMlArVjZd7xTRcvpK3FQ503
Aj5KgUEktfPByIwMz6I0mM41cW8Xmd+y9I83RfeOabRdObhphzl+RFK7FJnp9toi
C//LrtJCf5goTr7JRUZrMlNue6zXHt6Y9NUQtiv1zRRTHzejLjSxtNVJI3Eu+iGK
dVqiLasVwLQQ1ISum8mePMCdKO8TZqkuPXZfekFRt4CjnpRB975oBgn8zYm/oJdc
1RR+bE6xbZTxLS76wvsthIT1egU7saE7dlXz9UgxhF2pUAzW6snUSlf+MGPpIW/t
eiTO9fAsgLdGQqxuVz77mRsLjkExcKYbwH38Hv7LnKIx6bLlnh2iBBhDy8PlJmyi
kHh05hFBSBRuTlmH9Ul/QBGgpdQAeBdBbvINm2XWpCCjaOETL7pBbt7ligUTqWL+
Onul67ZrKroE8GvKFB1FBfgc5aVHG/aC1YTfJfsPthC3fe4I47dBdkm/qo7+mALd
ATLnP5JhhME1ycbYF2v9iszSrYFS9bM5DEkBGdRCiFk0ZLq5t8wvqO2f7enk2TOT
AcjFFzf3ng17dkuuW1OaMmeJ+kaLl2uBFapxGg4bQk0swu1KX8FAw94rwTrRIuUP
z0T/qhWMa4mfHS3OyrvhWJH3Dv9rIIjPK2zikQvJhOb5UVd33nP8dQhO12eoKTWg
s9CZdV+kKSL/B54KJOHqE+ix7XJxwFwiL1elWj9b9jzBG+477Nq2u5KCAeknVk3x
5fCppgX5G+JNDT28+TmJdwOhFpz2PoZVb4bL1WqM2FuHe3Y/5pSP7aeQdslXGmQG
cAE9hIiplnmAFttgGPYkJnZ965A9zCgoGHoDTvdZYXLWkfZnu624Swb/0EnZw9ye
mpONKSHGho+onVZRlY6OGqtpTmMps7suHvaPJujuvhLJcmxwkAvi3teuGI3XQXZN
XfLolEPfnVHZ4743VE/kTcbeNqbmme7SPgvj9TAhxVqV8mfaBJqpCkjNVs5NAitr
YItgS5RpJD3+/nRFNIHUxFBh644X8BUFC8Y4GXgKRhGasRUf7c7cJcNj+CJ3cFKc
D9ZprPWx325h0wj8T/eI178nk8sxYBeiF6AD00fb15ejbq124o4j7O3FXChnRpmX
8cbhdCVcNeRpqSH7LHafd9XNgiJQW+Q34W7f6FyCQCnmRC/NoYv11O0BnnS8Z/qs
pzbYhtKA5NXi33c3AtIzJ38iVvIebmiV4lQiG5/lzNSIriyibEo4GYiEkyZeycyl
SlSKioq63Bg8PeWugULfeDp15hg0bSFiGI0tLNoFqOlpMh0z+c1cP1O+00J7nlY4
RCZ9KTD75bRbuQikhE7vjsrnDxEbfXsAtR0F5oN29qUqy/CSYd0c4dyZr9nftvWd
d0iMQuS/p+9lfPU+zqCbfKcL9PUpB7eIbDKnQBDS1Y3k2awcQqST2wSKEq97JuJC
iL9sk64wo+zN2g/zIDHRgt5yI/nswzk2NDVf4NLAgOZX+uxQifJoHuy+eK7oy0Gk
o2fOXhL/3+m0acGeE0+S3BRF8FwFT/1aGur5aAP+C6R4oayodBYoBWfND5hYg3Z/
uqo3grvtkPmAgFEaxIWkn4w9FEq3pF57U4b2oT0v06A/iNr2EbYdcya2v8r5dc92
dVbYiXp4wig5Je35d9aPzL9krdsfnsrQ8fYDEiY/Ee0N+SWYOlkdevrIqQX0oYv+
4cPMZhcXxZRknPpWT8Wv/iUq0AOQYGo69U0AbJ2zPcnH6R5E5qQdP6DOceQ3GXRV
PzdmjchtBOazP1CGDTP7Kve0KjNUJ6Be/B6ffLPBMvvF/5oFrBBxNrm2sAOzt8FX
OC36iujkAPupC0bCDGrhlrppdrEPx+x1FQotvXzYIjcud0X6TpfYSa1PRfe78qTF
5K0KK5RV+2AUDUkFWZmZ5ZFjUBNf8FNtiSXVzYVgTXCVMzx2OLjAsUsqkb+sa7L+
IPPlNFCoyFSTdFgXLvxPc9mB3MJoBr/N6fHybpowMenFuatxwB1OTqzYUGWnmbW8
4gYWLCrcFaPEl6uPfjZezBqFJ5cQquxq26t5D+sCnR1ermofuStIWzx9uSbwi/Nm
DADvNHNQR4J50iY4lkDUtAwb5md1dMbPv1A4lx/5zuyGYbqgYCu5DgaBdmnM4zhV
ZC1iz5TZo6rH1e7v/vCTG4IROSOFUO8y6+0i1Lb5J0VgioAp0VXkibe6+JfZaOLX
fLM//SA4xh8xFvF7re78Ckule2w4rxI5h7A1szcLeZwz9mhQ00onidW8VDy4v+cN
VwTdMmfcZxhNct+jEe3htsr/YBFZiHg7lV5DTwDOCImWPBpJ5H/08wH+Eyvt/GN8
IrbzryMGlg9yvlvBK8HCsLt+0QBIC531JIKno6qmUaVO3ze9Vkrki25oP8fwv101
6dginUPquOnUHtFeS1roJTh0l8RQJOpgpdRsqWIfCdcupYA9Th2fzH31NDWQ5fTz
kgo9ebxXVl80j/Vd/eEJcTND8rM2TEuTBheS4QM+3E0GwCT0tnbockZINADNqrjb
RufyXe7UR5wlUOajtvSQWvZNCzB5Gda+/Q09OTSPzxoQTt92CzMU+hpYqzK/tm5O
RvkhD4W31cdGzIiJpCaDCM+8vY4ywLsf7K7cKya/9Cp0X7uw+9sjpZ4rvYK/4itV
2uMlK1Sploe76+sqXhTUTBf6qirat5bg8SemcQHmbmAx3/hHPVthlxB05w6cOHl8
KAsPgdIuyQxy+kFWNwOL40s32ZG+QVL0OuNa6oN1cE8p/5zHLBZLyFt/2KhnMQEV
CEiAD/N5unanoHu9LcEYT570pg1gf5jinnbRD2xUEUv7GlYVfRQYqVnbB6xZOLTk
ZRrpatdsq5E9aRt90PWyqfgsXRDc+xm3Ah37ncstr3EnlZgy9XQVtHHMlfLPBo6H
PehqTo4nojydXDN7InLLMr87k3udYYtneKnR0ak3Tm7NngqClU7bRCzhygQ+StP4
7j+tIByMaK0a2eAgQhWi3s38JGe5LnSiw9irgkg4k9yox5TOafdUNcpL1svm/Unp
diSLxwRk0f6w9rHQyi0oGb25b8wGH4EKRLH22ijiuvYNtMLLXFeBWAfEblX0KwhM
cRai6AP8QRW7AfiyXQbebT7dtrcnHmuEnYSgN36wNX3KkZm4P7vIxciwpuln2And
ZVXxtEmHlpHmvrGet+Bvw1Hl0Q/gUibYZwMjexaO22pKw1bFvFhq6I6fcqvLiDv1
LJmmKNxKPqyLw2Il8IVMTKxw36dhSkk/XS6+A7MY7WwIewrRawALFdxOyCa2h+ex
HD/SU7Pgi70rdGY406itxNks5fYsNWEL/wLVCqgw68R2ImBmJ3gDa2FC0CuKb91v
lmG+UndR71Yg2LXoqyczfWnTCLRjHThqpIB4AO5TBMr1E/YQaLey4rSo+ofD7JIc
/IUgF9vWEgnWDE/aB+lDNVplL5D3O5j9WXJKBoutAE/52Ukt0LxTRlkyZZPqbdHK
0labRZ+cZbdai7+/7UyPcmfE8ISzICPG+yzYk7fJgitO353puvlc4bCBqkcNGBY7
nBg+rf6pLaSLatuxrQFXVbUqlAcwe780CMZWPtlwjQfxQdCmm1aPjwISv/X0o8H8
1aebVcn1N1lqdUgwHXr5zL33N6IFex9aXgoQn0h8nbQQl5te4cLsruWYz0fsuTkZ
BsLVsUuzKx74KImEqICjmnk9milfHR4xhGEqD9UTbJjbYv+m7Zdrzzb+O7MBuWqV
attnwfw+SOBOGSp4iPA+SlIMLmKp3+trFJqhSD/lpbtewYkcJFwD102E2m34gAIO
oe7HyQ8GjU3BrmlO/34gh+iJ8Ar51a+OI0qj7kEUXus8JLMzHhI/a0LZxnS/gs03
2At3DlN0pMyrWghX+f5d1hNYz4caSIC6yJhQkIJTPykLGsLkJKVanXKMT4d/ctPa
RfquDP2gOAXC2yKiX/MxruiXTFpqCH22vud7UQ0TDiA+u4H3eD8vYZVyGm/LDOfQ
U6BFf/ICUGGGPheTo6yGc7utWpwUIhbvngdXhqilR6+ZiDxNRMK3VLAGRc2r+i+M
PRn8/p2Rnzd2B7rxGhG6q9HwfwPRaEVpItA+OEGUzmXphIx/JZFyXcp9TRPK67tk
5YSKpRIjtqighVymufTUhu7Hmz5rXMJw6m0W5HJ+l8FBy6EuV0lQuez3o0Iz+25K
8XsClRI8PyeTSY4DduyAoEsO71DLskq9bZc8mC5czb6JuGSvulSYYR11jOOPw/lw
m3nZEbjI765ozwVZ6jJb4QcxzJwLvmGLorJZNxWdw5sEIV076OHZJ5yDW7P6M7lu
2d8V0CtU07oEuoMcbW9V+jRiLqi/bNjiz4EShH5u/0R+1hl41Ioy7XUBePoPzSta
oUID/s+mRfQe3WgWjEbxa4gIRtO8zowJhC/AAWyYaU9QszICBdjtHFGL2fStvqAF
h0EGQDSblz4yK635T2KudQ6JVc5gS8jqe/6+HLRarxap1Lo1ldvE3qtpUQRo2bf4
oLLQdcLmbfaFnP72it7RjA8MWcQ4/GqAqXIdHIm2nbnVFFxl/fjxYYhamIRJNuqo
wa3ynZeX9toZlChzwktlxtWtu1PHERM/GVZK7V8DSyMiXQsB/shewFLs2A7y0nvF
XAMNjVd8WymWQ0EHre2S+Dg4gvdd6ugizVJrluqXrR6Q+1hiJDDY1NsDIB7fgNFn
w6UJIf9xzKYOlTdidc0SQyTngrsbVsi4Q5LC/i8AysdQN+NC7M9jNi1O2L5i2tQw
CCbZcj6jo2uhvyVfkPeQUIBgV1wapYaOzbluGPubE8YzqqbmyuC6aWYUyBv6Pxl3
ew+68JI2IzvQ83FFoRBhasXKRo6kpYxet53a0oWegVg9AT3qXupdVu8xjL5xYUG3
8dauwO08tpXy0J4KEQvrZnttpWCKuME85eDUHc2JlIzAfHhiNq0lyNmFMAsdWRjo
G850LhOoVQKcNm3RIjFsSw63mJRzR5ud1WyYLxZJLelS6/hv7+76A0srf5O55xdw
OAcRZFvn7lrrQWS8hHu1BRWkhFs8SByt4S9dlubFrEqtOCytnI65lBNaIDoF5xoj
0/UsbDwBhzdiKCBnrM4whTxA+4YI0OouDcShS4ZuIufVZb84GZ/twVgb2hkbplSW
x9tiSfS5K9X7zCtvMEdMdSp7cXFcd65ZEm3Kz99OOo/pjL76iphaD8A4o4459j9T
ZkqqrxR81mV9GgnHNxMmN4wymypIfmIZ5TFQUWbMIBEklAcx0zgjlcF7QGNwPbmg
9Wf2Tnk6Nyqp8dM+rHdtlMzhbWHY84d77l57AvR/Tb8pyWNDlIUCccTEKpTceyq8
6cTszuOZFL8cWz6eHYIo4V5tgbpIWDd0wIHjbYcao8rnHkKooQGfJmpfWQGDUAHO
aJ/vmcsMSfO/fcpnvveXKUvarub2kJOQopsthBcPk+EBF3UtwQh7CoHpBbVN854u
zPz7ldTAKwprbwfscMJEmmFLoffopTGYUOY90q/eO3DXtKX28d4h5wV7h9YY8k6b
Denx1K4vML6UtqaKU9yNBLkFLAS0xZNhvOvGf+0wxYOCEDK1hdfHKUq8NjSqe/Wh
WjuGvN6Jwk0wlepb7r6kKZrngT3rpDOL8B9wa2wMLZTCn2IbVMde0V8xC5J/I2s4
o8TcJdJkL1nFp7MjunW72OWrNPlffbl+pwDpjSXBU817t12B8OLHDfI+5lNOkoAO
lCGY2nJUZNIxTEL8xAy3EU4D7GY28Flb0jOgsjz4GgykMGK25L/8cIPqn9/pAV4B
niHqBLAJ6HC0e4DFPEAfqJNMB/0+ZXqXL/Lh6i3/aBz1fPj5/ys+p+2LaqrxyV2z
CnUxKq8ezjalYn2lY2vEZkwXGa0vyjTtMLqFYieJuXfbpsg3G8OPfAg9etUJLzl/
KRgxwm9MW0eDKawrBTj6Ce1PoFQFtMrDHSpTw0cRerzbCHKMZRmmC+KT1MOC16A3
TInG/qgdYopZvO3kzP1Dwl+PMexv1LPmuh/6wMrd3DvTRDs7x9jLBN44aGgBJ2iJ
ofYqgMrmvFKDgvbXPTeUnL+hg/KSKbK4uVLbTnie7GWN5iIIc1Uw+4DHtX/40l4T
qzWWxdZW6gdm3Ef6TjCIUt1phG27AorW4DKA+85U6zpCQqUy1npMjcHwue5cCjPT
46Jgu1j3c3TNtNgj8od0vg9WlK6oZFAU2ULysLrKG2xwp2b9lMcF78Mw58hAY+yo
VxDX++iX+wGMO2w7BqRP2x6WqJeRusebHYSEcbNGahVPH/nSu0pOjXMvk4iilLMV
s+WqUxQtsmGX00aFzbTYxTaZ9ip3m2XRXUTnf79hrr9HgoIoqHCC17XpCcDx7G/j
FFpVMOzKhhdhmHx4Mof2LzoULF1vlNg4Jc21Psso7Fz3Ny1qH6IRGZgFqPa5Wno6
oaKzQ44yZ18hBk6gK+rpChZztVZFOleXH+fQF6Ovrob9zuN0bO0MSRNGoM/FDo5T
BL7JHBV1NMTBPXASIJwKln3+dB2sejfHJToSSEY8SNExgKF0r9g0vS3E8Mt+SQR8
oAe9cZPiMp6nvERgRDtdKQIUk8XOwgB/FKStOfqorFUw5Tpj96dttE8EiVgTu9/Y
z5ceHqJdIPB21hm2vi/mTBKzs/YGKlfiuPIFrygX61npZoetg8H6POJoKrWnZwD4
eaA6odUQdqnBCw73bUmVyHDIXYsiDXJJxZhMyZzFRmbC9vWFOx5s1dn+3wJ2ExQW
80clw8GwMSj5Evf5aekf6aNLXurjKNoXwMasObzRnCvy9Ymt2zwktFJ9cRylcEbg
pK8OsziNytFcB9l2uW9CLwWsWdPSrZwBAgGZ01FYYcgwR/QNsOG1aKHUKmPLz6l7
f0Xy5vX9yLyLYOaJA25r5t0AoL2rTuqb8OsGnjSbBmR9BVaYRwWY0mdaKqFpkySv
42je3Xs+HNnIsQCWx6Sj0WfwzPe5QnyxF1hVURmnSuq6VH814sMbm/IxjqWAm3OH
nO9fKdQh8XGuWTLGQjinKfWHv8gr9ZOQHdAVJZaGGNKuvSbkw9jlifLlwMdICQNQ
x04NQz8aB0gNZKlMD5R43B97SABEMInFMTTKgeMvlD+xUw0V/Qvb8/kJzf4nqhsa
0o4l/3omExjuu+D0/XO3n1JWCEqC3k67fym7vO6nTlKaM4NHm3vugH81smW6hDhI
Snq2Q0lYG1Jh1G7rQtAxMsOIvDYwipt2/Ofj9u9clut1h2eJxlaJr8DLWNBktMZi
LNKuGu+JzxWAhmMJgvvtivqUKgSD7xehZ8BPEPTprudj3KaFqQa/lEWYqv1Rnb4m
ESRYn6KFIQhjcmtmp7wosgVLAeG5inAddex/2IxnPld/jPOOPLt9wedptrTD5+tK
N6QevwbNuKWY5v2qttA380K00FbqBFD+mDImK30PNpJRmpenXTHOexxmWzGNLe5u
PZ5SzdWHrEGslgHKMpqpA2sl8NW4GZtjCXsrhiigjqPIBGrqRzLDrat+t6bo9Gdx
rdMgBQ9Fr9q0FA1UYV90RJESkXDXvUnQCEoCI+R5cd60BtpZkJUr1aJjYby3RqfX
64kej6uQZh/JlTPiyc7pwW2d0teZu33BeqBsmhr9EOVvnK/JaSHrAIqUMp8lRfqu
h/c17pwKAw3KNrCC8bKLA1Jay66YIkHIwTVi3uwSZ/iAasWtcpyTWfJpXSa90Ay1
ikvx2ObcqL7BAolptcsjHPh9xzlTOlRsaPhmnd96OekFPFOzpS4JnPgjgErjuL5H
1aunO9UABSA8E6l1plyNH3YT2PbNJsdKCBlZC5Css4EPGP/jbJQJnfWJbMFJbsX4
vAyzJCmzbKAcoYMTfdvZDIelVqn49DtAuBdqkUTNWeEyioVF35Z81p/mPE6FDqYv
U6cfN0Ip3s9QgqPxGKv+kpFh4PGM6NTMmWgtD9V9tAl8CaHg4rjVfSTzuhqOWhju
6RxXsv65ox5n7gy5oqSHH4NNIGXdkShzxuuT5FUZR3SJvbWnU/PGbLV3aaNva94L
c9NvEsayb7thD6ZxbeMS8PICs2p18D8ykhjAzDzXU507IHTg2v8T/7Mm+Pbi7rTl
GdEeQsX6CS9t7dFR7fL3Di0mS47UIRseOU0e/bW/faXOk3skUjWObuSt9ZhJCt2w
nt2BFHb/XVCq5azEVJGNsSq4p+TTpJccgapSIYk6wsIBwMaRRQI8rZml0LnPWBGq
EqauTi2XVVAnq5r/LzrxJcgRdMjCZ4aRkU68PT8aeWNU0is4RdOIO55IbiA4T6sh
PpFBt3HlAt2ZlaGkH1sJxVlk2BhdkiCWq8u4mU/vNuvkXuYeK6zsn6JP2be7f207
AQBYIc0aGGoHautHN3r0Wj4FIw/+On/I7NO7d1W7r/IFUAy6gkHmIldgfWCvpune
xoEM4zEPfoOMfZCBjeDSyHpXSE0MyBNoPIaTO4eiSRGk6VoN03uB14QSo4MNUW6w
q7Qw4iMtyuqzrh8C0YP9o1y68M5XsHF/MBUcOOlbAvuR4C1Lf3bsMpLqtTGaRYIp
7JQjf3HR7fED1E06mC2wwciz4ku/O/aqme9yrbOzjr+IoEXwpi/i78CE7Cab9vkW
O265j1FA+E+IttA1RpDuDPs+46VZ3jGJJsoIElTj8bo+SOtS/wEMWRMORy54yS0T
gtiDNLVWXExLa16QkG796IHva66xEIBIW8nXuvUvPHyToSvsel/thIPwmQ7xT/E/
1RBkumjA7MI2BJg+6LP3rrSDuV5Mas83FqWknB5i78KmksMPgUovLeit4leXdBBc
vhO2Bh6f+arCmsZix/QXNzbNKZGEg/jEHAcC42SGZzhrnQIddSILPtOUwtHsiklC
vcbTqaYdFZ9AzTRIRElyFhw4x5U7WncdgR6d5q14YklNxeSLrldeAwJA1XLjQ+jt
9kkkGoswCjwTMYDYVMehBbJEOj4PRqwtd4V8/XzrQ3JA8QkVBvUnbwA2SOx66/Ze
ioPMaUW6/CbgqWC9Gtn0Mnl2inVMmmHZUU52GIbDZw1g2wlV70ldkcDLhZn5Hk6i
g0TAyIwFwoADSyz+0t1XHpE6w0HZuRnAgILzoJ87KBfJATUIy19qmPh+2lNxayLu
kHMlFmCgowjgbRo2++FTLnEOET5JPCp7fCAbDJb7FfTzneLK0wtEV9WRGaSDB+Yt
xYsYQqDowtHoRdm2FVuorJ/X5vFFcFiG7DcZIWpIDgLRAjMpOFOLPO7Ul/vcP8H+
GWA8gClldd7D0BIp50sNd1c94EwqzdEpce+w5+/maa5Yyu4z8kBpQGhFg7NwRMuy
/bUUdTOscatV/nRdh0X6FqoQwXEujvGWBH44Tb1iKVgiOQa4tUFI5VmvYRwJI3oe
TC3rHstYtDSvEVts/yjdh4hI1BhtN8YOrJ4568cu0WONVG9xdOZyygMVlebaMY7h
szI5DIC/l7dAixbJOJSx9lN1l503aGub7T4ozDxxzVCzumSfSv//Ku5/6JGRC9kw
jP0gqZj8kxyvb3lsToPYdQ1INACBRC/lqtVJVdOFzjdJkudOgDMghwoAFNLesjyZ
O7iUgXBmzubU/2JGt049PFi8f6HHe9S850eqiOc+wvb+EuB6jZyB6XUiXqtIRw6M
FJzN9p8eis1e8nTSBikCVeIDAoWSlT9/UylQVc8TJon5ZObpf9X7qeYpV+fDSAbq
YToxxQNahM3up0bZtvlDk3UGv0taqajIk2lrerb1c+bY0jrWmmibv92gggsbRS2l
LHjldpskhLY8BszgUmCDYdKiwc9MPTONdK+OSWkvlF9FsJyMDfg5MT0XV0a5pM7A
Za1/UXdjJgpzCO0dREuuONJN3j2mfDLr/cAVHGcTI3sbzCPSCQwn2PHbK38bWVq2
7wlyzNowHxu0jcaxb0G6SBLTK3/UTqlY0gtferSgU3uqY9ZXL8KL0TZS55SRrQBc
XtB7pWMR6EKXrh6pOhVX7s57+86Vd4xYFscDvTed4nAQIXlLwm/tgeSE5iG3gI4Y
sHx5eeKgsSSAedkVeWsYV/M97hyLNB619Wh7FlFoBCUsSQHrY0UZLMHb66kBpDmi
W18m7QZICpOnPWJoDn97Qn3TYgB5MHKeM1AND8GI86J5ws+ql1DE3W4ZHIXleqfI
N4qAUDRRAX+yXRyM643buLtZmoux5GznvbC45FGfjs2tgHP9SKbeb3fmfHmp553u
7IF6q4DmHolflw8iWNohI0MDRwUdb5qh/djBvpUgrDUL3tRKopI/Jk8ISaJCdnmW
XyvnjhQANsYLU9VXjlh8NZ8ieYltwwMdIwHWuIKPlevPxM2zGPDQK4f6ssstniLx
G8A59915mcHBqbV2ZUvxZGeq7g0Q60bI0Y6VqumjAslU02cRq3ys/Ar1OagxA74X
gU5lxN4JEdDgbaAZoUJRbzPFubbd1HcLbTilK/SP7BH6wTLmNZe6XhIX7XQmzRd+
sIf3B7NCgbGdqLiVbQsDmThkEKqHL0Qejda1pmUIAqgEzQt9epoyWjwn6xtkO1Eb
fREEJrPn2rOYQwfiNdRE+XSzgDPRbpjkghFCDjV1t1mcnzyeJcl26YZctFsa0i+g
r/Auv5GctKoKkEcJGogxzpRCBugJb5SDjU/Msp508jXQCJmqugItXkuSFaTZEdZH
TZJiA/IPbFsNYZKjDyEb7h1a0qt8fomiB5PwZeofJkHvNDGB4qLP88LT9MrNuosB
NqedMbjBAE4+Ow9fhHn3o76AsTHzKtoF+bB7qPSaz+Ya1oTF4GIn/gJq0slFqJxV
uLPl24Tejcb/JapFY/59x9jPjJHoDd8ATqu+0eJ1dWHVI8LsXW6tsQHBJi3UFtNJ
XuXP+gLutRCf6kjm4QVqQOC1kHOSrpqQSk/LkiS/4b/lr5Z8SwIuuTTlj5E3IQL+
3LXO9MgyO5N++j0K4U1VebY/jcpOzmLE49Lx/2NnN94CTvDKWAKYo1jTY/UwWLFS
vhrlHHvky7Kx52JIN6KbJvnw3nsBBydswsMOAGqRcxbwOLfFpC/PiO1K6i5/yOVL
An9sNvUhXyRR9MnsWEUjux847Hnnmj3Y2ERxtdJI328FmSxToPPiD+/8m4LqIuba
N0lQQLxhx/U1/FZvtAGcuXkjAKGhMmDGotdox5EL9WIaY6t2B5aryiW6bft8XT4x
2AA+HzJZ5qCLSYMeGn63FKw7zPBxePp+BIPFacNrfAg6KgdSXv5yzyBI+8miQMor
ZTg/FS6aMzuqM284RTdSFPcUNhtFffb7JGgoCgeCz1xXvdM8Lx0vODLAV3ugsTUY
UBbQ5KnY8iqCeWhkCauyCVG/JQe4z82Q++U5wLwk8SdOU/wDFFmolcaD8mBjVOu9
r/637HJBauUvTUi4k2EWIUQTwvqdGgvPQNI1aCUWV6kFmA2sR9V3mgEUkqeX6vFK
1TMQbR+ZpJXe0jAqswSup6Ft3TcEbZJzUdGPpYX4alXUaYNbbmCNPLVU9Guu6+sd
4fNMtPNBsiCpBhmImLARLY+9SaKXQ0hC0HR1uLpeA++iJNGj+/YkO6oXClnQIK4b
4UO66tu3icxV6IQaX+N/11dAKhBnr/8ZSU/W/Mqw3cIzCiXvJty+jOkDtU1zSmlQ
XpdGDjvoJBzFc19Xu40GV7kbcGmxKiEHHncOgQMXRezOfamtlD55c48AKKdc8x44
/9f/PqopY/B96R7iKGgdL2Nt2DgaXzPbelEG1nMsFQ2I4PVZnKdeulVXwKyTYuw8
c16ydnf5Y3IUnscZ5r5hfDjHxtwpSm5RC8JdpNpBTZ667T1bVDGJHIQy64gMnGuB
nv8FTXdqtT3Je27qw/BQ2HxXBMeQDplTbbdou5qEbZ4cN2L7+neoBC3HKetJ0Z10
PwWvjrNiiv7zKgVkXEvpftnjKsQuDxDGxMWikAFf9YJAKl0aMzkNkaWz3WFVYOEF
DTQ+j6XpMb21n+tXX/jbUMIz0Z6PTia1YwAWWMYHt+qejCzxBB6Y/sbS33fDHe7X
XA9c1vl5lWe2+09wVFl2fMAMT7FGdQzf/QcCKL0toUpNOp0AUPyMAUJOHkNoTuXY
107dc2an1v+LUKu1IC7Y6fH6HE/HctcSO29rcNi7KUItnh23TJ1NKhkwuplLrqa8
m+AErExKo49x22L0dRsvnM6KC3MElktVi8xF7RulQJf1oCibMBDRTEPIc8/vagOH
pn3nZGZFW5zWbL57T8r/nvNVSSvCCUIS1nUpccw4NRYv1B9lO25fVQsqg/xk59BI
veYwDZ0daRREH4n+rxU0uDeZTDxt/CYk3OqpxQ9famf1X5ornsKi5P2oMQqQwEdT
HYk9HPBL6WTZ4Yo0+zeSMRUmp1jY6jAQKipngyhDx6WEeYGmiFvQcwti9Zw3d1fU
Gwc4AIQPyRjnwoudexjWfXwvFVR3XyfhnZYkQaKR8nVkR3G1ZDLfEHR2X0TUq21+
WG6cRXjU/8VXxc/YpcufICnZhkC+HDV37KHiggTP8ieQexg7JwgemjjgIkSLzf1R
n+nFPMcpfSN2AQtN1d3YGvaGvv5Ch9F6H28txL14x7j8XYamtlzt3FG3BMd6axS8
qlAjj9P5hLbJH5NU9k9d/G/azQR36C+0rqfaN5lfSIJdeId6neX6AqQEERywEOPr
M4fXuGglI0EasZTJDH76mUkZDwCFvYrJ+RNQLuhvZUp8Mmsj0AAC2dYnyZpgkaiQ
0OHpk2+b11PW0kcRvwex0OqILyxbf94903ZGhTMDIQJz12y9hA77ue/WTfvqQHnP
b4hrFwrVpinfS36oTq70LYAme9/LgF4WlIbdtNUM32auY4BIyvmeFGu4LM5LDArY
dgLbGciqh63f9orIO/lHa9GuughtL6hPMp8lP6/nnZxu5BHpZib3KekXFNxWH+eD
uP9A2J/wXBvEfbmaWWL9ARMrjSPrjODjK+IiGPxYiSPck0zQ7khjcxyIEo/GI8/V
31Hvcr22hB5SyNHdPoJ9nHBgP9Fc52ynyiQacBiDOWf348Yfs0z3PzYEjYKj/JsD
nHbTqVeg9uDGBWT+Ij9AqXSDWv/Kyt23rsMmFWJJrdlYmV+mRtMPslhTdyLFGzTM
ESZl9RfGzMDpT79CZGuc1o8RDrXXNvrCMtP5kS+hzA6XOTE9hdLrWBXB1eGusD+B
HjQ857eojdGud6T3I3/EXoOmn27iolTvhOU5ylh+2Wx6tgOqe6hPzuzKly0gGvhZ
WIuetbi/+70i2Nr/WsLqIWxvP7ajBZvOPSYeYt2cOjYxov6G3grCxUBIJASdLNsX
8Da8+C/1fLaTUoAA887KEixO8Q2SqcFk57jViOV0mfQSiymTauXZwpP9L8mcq5e4
zgPhQcushLUeeDLJhAdstom+M+bTxf1TvKuAy3mTlN5zl6uhr4s14LxgkbmB/SCe
IPQjKPYqiZ3PpwcYVyIDGm92i1Qyui6hi1QE0KytOM+yfxt+6zox4gkqMnYlGnFW
Q6Jkz72OeZBCFEXPNOjVeKN+NdQdy/hZEzmFoNYerpRLG3zIa5tZqPSHE2y0zw2o
3nbhO61h5xh3xoXE7PqTJ8OndmDXZfJ2wFrRLch2lfwm6A0GLXht3Fg4m6R3+4nF
uE9BuOw3AZxrP6pQiK8nJLj4SrnyMXNUDVKt8qV6UDlR1p2p/mIF0X/7QAGE1Acu
kVeEefR8fvKk9CNuAWKQzhNvB9K/E256EJzxJ1qtgSpD0Endm83CLdSh16zv1kHj
LsAO66+UaBn8WwUjlNz76GK+7aeKIaGipXUt5Hk19tn8Q2TAj0w42jIDyxAscl72
FA1bq884coSYMqzLzxeILGU0MTzmIYpG39GdLE3m7lq14hAdmUngOoaIYpgSe5LT
ZJ6oWoDP6vQny3rCks8JEECvD2jiF49K+D6KG1Cljqb71+zUeW4RFLOVf7rGkshB
//t4US7sOWLf303OduIVv4KIZ7xBzHlvfEUwA0HpNNut6rTSFWqebAoltz+db6T5
J1VEkhfqZ4olBmCJNHaqOy2pRoAmFlmJUCGNaJVKdY96jEKlhpO9cLLkv5WQmaUQ
CHaRnk/VBHM2HXaeMuIHhFaTGsvHQzh5573OkyD81URBrffuLRaUI3L4y3wpSIcf
UKaPvp3JmC0aiNHxykFjEkX/iVSg1i6HjIqHl20PdSG8M0nLHnRIpfeZKNH8NXwt
Bkx4vrQmCTI4tGpnAsgpQ0SwTmTtCKVgJ6gtIW9Au0q4f/vMpqPm0bzhX8OvIGKa
V29cPh22z5aZKD1SLNHKHG/aFzy3sse1fRWvE6WfYnA2CoCIj2c7Y2+dgIHSsehM
mS+a1hIcUfvrcW0S20ot/qWixAAJxwNM8RQKccCK2bBWg0jNDd0bQwilRi23Y9Ob
1Rpnb4cowVL+iZwSBXLcTGeC9jM5il2dtIFmaBWrZte46wI9N2OK5AeY6pwG8ot8
hLV/cEE+5+ujLlu95fc4jItGJsHsqts7kqgXARopSMub1szzBYC8tJfGkmE5HJHF
XMgyxb4wBpsny4QCD75r8Fv7bBKKIB4m/E+bTfYHQgXwGTAl1KPcRKWjF46JLIl2
x9NQYpXuJRB+tfC2KUMFgDhLUmuOm+UBIDhyuexm1UpauHb+V83aqS/zDXK5jgbb
0uEOgnIBoHPMN2QtgfDa6xkT9DSAQSTvu/0KSJiNWHPmAXURz1iJX+0aYmTNwI/p
RGyPj+9B7FtVyHRxlPthykCAxoJqCUIv/CwKPurdWazryaU94v9l8uXTKdwdmv6H
L7XO56t+gs8ISk0IlYLMI+eICaWqZaBSIxB3lZS2btzPjbrIH8jXn02yyTFKBJUR
pKdGVJd+wA6GC2uOG9RYkNJek572r8NnUv76452hAxv+Yu6jihYXe8BlhycOGG7T
yy/a/hXpGi/lyppVKDTbVEqHS4CLLOcjO+p7+AmctSMQ+m/EX9kJPJpn8zqpfEL5
AvvCKX7/oaV7oAkAxdznFiB/vilsXrOjueiat1SjYHLY0/ki3XAVQXnyU6515278
vTj0LJvfPddwGxZkb98Y5EpgqpysIj7HR2HbQjK/T/4m5XSyclAr8f7MlbrXnfbU
aRQdvrPZ/65Hv64BfqMnI5ImH9ntEVqWmFzGPHSlw3fSC9W/H1k6Lmu34UQFDSKb
02h7oyKB9VuqOT53paiiDFc/iCfiqbIozhroRqwoJ981wx8I3loXt5H4kD2iNarR
28MK4csERw8shr7pcgwmadg3nMp3w2TrqerypgUzHuo6VPy9V0cr1x2KlNHwJl80
Uy+JYBCnkbCiiscS7O8Or1bCHU8GLQ++6jhzqdFBac9sPW0FW+geA7+d2RhMoiZT
wpc7nmLUM/mlr11v9uvZrihQ278teGLCLNbo+P+oWEWf7sD5PRUERRbF4b8B+K76
opHLQTX0oAGY7BkNdk0gCrKx8tx3qNsUEzq8JDhUn5pgGPda5aqPLTJ9dGicdlAv
5hdsalCtqVHhxGA1Eo/XgcwFgZRh7DEu7IMH9oAtYu3v+mllDjT6fsb6wyfi15zo
14TiCNRruQUNJl6YmJLTddzA3aMwBkQVykDiszNRpz39b4igJS2bBJjC8jGX0gio
bBu+HK7nFk0hBkro9NW9aLsfnq5Kq/djUcXcx/o4szocmjsb0wgaiTEae2Or+FLA
+x61C8hG/Ca8ZRQuSxR/4k6rXpqkMSpdySd/AxeTLaax+WJYVg882cUV17EAIP8e
a6ZphRXAZFgOPcNGpjCFDaE977npv1FBbYAqNeNigFoXsZakeZhbS9Vb9bR6TMVL
Bloz7Qd0r/duBclQ8ogj5b96Bpf9C3mIMiFXxETXpg0noHPtJdpYVrIeh0j5T0mT
E00nt4iAizvMlTCJa0v4k44q5kpyv5ckh+joaYYYMxpx0vB+LOmDWlR8dL2oRBcn
VKR6ywBYo2tfZUFpejXTfWvlwzVDzG33n27lXjdyZE95Ti2xE7vaIv1mW+ahgfWF
xeOtjBtyHhkLggZ+UPhNX8mruy2LJXToeadwhyEAxyLY+B0cM+SaGfnvmgymVV8O
8yknpVd/0jv+SgIF+yeY1EkaFmkaSNgOLt3n/5akqhe16kTSpfCiXFxICZJzHjSM
EGyTCbp7hntCHESsMCPDL1v95jk4/oFL2Eux5N06cZuGCtIAeuUjiyzGr9FS7/qO
9XxH3FosEe2B9h+V66LAQjhx79ajLvfIa5dNOwqX8Arft5i3/CStjLnVQi1cdXVd
v4Cw/QJcStgDnB4u3QdShVhihRW9ypuKpYktSH50QU7/4keOb1kLHv/qrA9upEk/
q/eCd6Ma2Js6UiZJqgfXl9Jc345YuPxpSGf7tM66COMOrNydga6lst+wU5O7eLtT
0uuFowgkv9byMSektf61/n+6JyzIVsU8anlLeK+yjJqLY9wUxHRdlwN26fHmPgrm
2GJtxJQZu/gQ0jmERtTTWL3uP/GrMDGstpqGxy3AybMRLFsRVqx9DN7vLJVnDMEk
YqxSzd500z67OvyyYmjf2xRhpYt0ho2Bwogbl/kW/B8MEn4pH7tTXpfD7C0aWrZZ
sdqhvHWKYk7kdQwTsnSRS8Coa8KTap0Ks7WXrw8CWc+wXHVRJ1L3Uw9bZBcc6/NP
e51O+A/rsqL7HrcctjsGUH1KLPD3/xG1Aip1nK7zLdDeAqp4hV1zR9IrZsIjn2po
PdVQbNULYZmUqHsJ8EM3yoE+USReP4qTBpXEl+M81ecjoYgNW45Qn/mcxmHzPBJs
t8W8XxCrcAogmyWox4VYp/CKsHEh1Mzx/oOiBap8kOlLnHRxHg5cbxaHwhQmTwvt
vfRHBLyzJ0O3MQajLn5PBSazKnY1ScSRR7PSmqvUz0RyvrvAy4fG8YfZoaehLKKg
3OuWzmi3tJ0aK0Wt4B7IJ3tp+HhlxUA3n2ydWOleXJRpb8xzBllHp1CmFnmhItgi
5f1OJ3f/m7RzhsWheZPPC7zVUIqokQNfsEiSw8mXUUvibs8uUHpY7Ut48s3X5nKN
gWFGM/E7FRLRjqO7puauC6+HE10rIhItcV8tw5DQSVBYPYQr7wUe4wlVSBnJadJO
kEUkrCiijcpWv4H67FtEoQ7yFx1jGUv/ctTA9vNDAz9fJUBzO7J+g78ju43lAOtP
8i0YUZ9ba/rPhiNafi6wUphy3LDJXH3eqIHIgM3Iu6FMcLdkTX5vE8AwydQ8vCv8
xW4Lavtci+weNXnYpU770XUTTpvPgLsCICaQcurhto9ZCj72vbH08EdULhPnQcj7
pLQous2Y6XKxEIjPaEywHNJGHdPprhuhxxjGC3FqhQh2AGvQKVxM6kITSEy2lt78
f2mSFCpVKgOrwz1kAIuJXchOgiUaz8XJOaeatXxvlyPmz9VZalHwloaWEHAYbAjf
L0XhMMIxr0wHbNN/OnCzaZv24Ahkazkwa0tS4XQuvaJ4zNtMB+//Ov2rrGZyry0U
ltwyyS3Fe2YBsIAd9AGpICS0ypa1QUx0r7jInBAMfrliyMUetJZhr+IMwbkotxW8
A8zlxYiCgTYNelaGiZjUtSfLxv1yNxVaZSLgsBb7O/TMcFlmOfYAciQYVcQn8KbA
+PJ/62YinT4gK0rYIjFFdoSrvGfKfCres+cnZXBSENpC0S92ijQ0hLktcu3KxedX
Rbwq2g0YRpP23WnyC1uSknZh9MoKcpfavMsGCMWO34pyoM7gXd0n/uwUpgOe7fT/
jyBfX5z41B3XUzRXiB6QxgYwBMrjcPGONUnnCEh9i00XsB2OTLS0SjE16MCWjn40
5batBPBzipB1oa59laYqSx/cY/iwEDC/OzC3UNUfzD/bpCrzYNp8gpWF8b23wJSD
YY/b5PEWe3NzxMJllfZCi1RdkoaNJeBZtMFFTZhUI72sWC+Gbm4NtpgzE2Pw3Gz7
XezrxsTPyWr+UDjd7CNPy9XzXfGKiRGwo+T14AlSxZpIBLWh4gvmNyIUM6lWoVlF
5nEiL2pr/FnulpAnbI5kWH0A07B6bpTHiW1efrd3v4s5OjL4jQmESVRv+Ur0i3wH
WnU1InR2PbWGapyJ62nHficHOxinhcnMcbIsWtzGwQnSKT3zlHmqzVNL0Gv6Ltli
5ynN6RjrScvjhVafVNIysMKFBd+5I3q38amFkrx135NMuyu47uem0XnPS98PIYkb
3mJ41ZWdlHo6HWlrqVXYmLCGDdOUmwxoYrSy4RUnzl4DjQ0Ecr0wPOSLFnXmvtKG
HyCW5TSF4SuHtLeTrUqmKwKPMj2edKd3KShgWLtYMlYDbD3IcX0AfhieWI/5XKnA
n1FqYMsmBbflBo4Zt7tRPj1AyivEu+V+GJHvsskrY4iKKH6ldl/bVoIFycTo8UMx
+MlQs0Bpo11z8LXpPbIKaery1HKy6JXDlAUrCs7ixrYB5N3cjOaZEcUKZzVTRA4z
MxzLgsSwAC503WxvG8uoEUv+zV32Gyb2yZf5RXzsxKl3f58q2pPTEZF3taBTKsvq
nRU0ZrX54NnsVvgif5S0OQWHw+6PRrbXB5Hdy0LLrlWaFrfyVVGFQA9D6brwOuS8
JfLeOsyKd9qtgHNmyBcItLKjZxUHlTx9NrCWhikxB/YL9RPzhPOxzE6wdVqZKEwp
nzaLnShvxBlm9inJBA8yv/K4x7AsKEDEVxtQpYL7Yw1pZBlSg5nGWeSduEY8p9Wl
X7OS+52HA9+XMMom2T8R+ztDQzySPpnYIDlsG+eFLNYm7D21OwLX5Ez/biZSCAgB
uFs56zF5W+vy05Q9ncgE1LObi7vyRRw+ttf8EENC7kTu8iZhkQl+FoUSYVqqckKC
R+1TtoqkTiMRTaWKrXbmDuRsyWIpsAg0hKB9Mo1fOIpyCab6LGJKHkRkG16mgtBo
MJcV3NowtwezIGiwW8U64O5vajSYzrSMN9SImtzA1oybb82C3cThze5n4jJji1JN
+sAQ8hTfRFVS6p+35Xc53CKMO2LJXFEx5B/O2IqXCI/+Um0JJydO40cQAVVVHZwW
McmXy/+IOc0PU81leunOXq89AnLfJStyxXmbFSYcJBqeA+TnyqjwreZb6pJnFcYh
etDkmOI+QDqruAM5pE2+Km60kePvlEsffJBskXWwFH2RhlX1Yiy0CNzSk4A9FON1
WCzbbF6+Ei0Z9n+hBU6Y50EiUZN8szLM3ptl7oJcFCcvlOVLXxOmvsfOaVgW3OgC
8OChffLVeH6Slka5oeC/l8Rt5aPXwLOXl2X++Lr8F3IEPk7ewolmPObBpmMaOdY+
5wljEiR2uhdF1xtnrVlLftKJIUduah/2WL5anybeZPr71UvRpabgYQOsX/H8D4k9
r4qxsdf//Mvx2C+Nm9nfVSVp3bH0tA15vyaamLv4qO8yMccFro1jwJegSehWpvIi
gKYd62V0XylYrToEtO63L3GzqrsIpbDJvr+ed/6JlurqIzCruHcQAzJJ4chRRl0G
7ZA/4OQkwrq9AoCdA+RVco+qu+b2s0UPshjr+Mtc2Hsd2smTSXKLZuXfKq2QTw9L
V+9IlNsMyNJ5Q1OiTDbfChQep/JUgrAGXmS3Dz5GtK9v1sq8j0x9IDUMAkc5H1Dm
M/yfcIsMr/paq0FPs+BsNb39LEsVSTjBkApN3UJ7Y73CH08i+RRAD326yvXAPmLz
30ETP84jQsJtWouIWfwIH7oxYmNGuCZ+aE+8iGNNTWfw+n+md/cGEOnvrQHTDuY/
/nyGhxLt23rLyyYTbmTWseox9XIDzZGxCFRjgbMXrYj4swjNcwwU6xbpp4q+e7y9
JKYBkPHWTbHm62zWyHY9I3kZ6TwLrCJ8csoc/IQQgLlJgXPkE2ZxZJIMXgu3Qq7X
7HH4sNpPdHxndYTiBLpdDtdNIsTS9NTg47iGfkFQgPMWebsDecfALj+CvzqTNz8n
P3o4pcuPsF1d1kJlR4sDGs73/UqNf1Bkam/DqFmTkyJTmGaC3iegF8OXxgEsgsY9
QOHeCkhS7qgUN1mzY/o7Awux2LOYrvpF5VBxroojJXXnBIV1cEY2gkAbP6fLHHno
hocswToyabScbDB1kjnY75ceh/zDdtfulYqO10LP3/o++aSJItetlFCgt/S+B8Iv
r0fRSsCgXXCn6VZei1T6qQpyq946IzK6HvPxGdYFTylSIkOUwSETqqdqvGRazV08
UCV3Amf4CQKh5Yn4gkdZOAYdQcodFNryGT2D3ZwImL5U9vCv+y7UY/B4NzdkOdpr
lKXCRpXrjzJTRS4zSC330/Fg7Bmjs5IGmnA1TLuphObHJAiYfPxxMWobT65tdw1J
c0jfzjPymbtAGP8sr0DOx7BKuxXfOn342qF0VhzDWJv6qjiMyJ7/g38yhpAGDJzY
VUtG5yhgvrQx4Ax4dAVD2EXYRAXGeaxTyrXh1TEzVKy8t2b8rUgDq8Rh+3yc3eHd
Fn/i3+ZSDX0Jy1l+Rm+gAWaNRDqompvgtUmCSZTjsxtx83/ELtz7Q2ncYZIQe0qp
HsHnk9Cn3xnKnk5RiA8Lg4cpJ12hkrDJ+NVowdQZ4U7ypU9qVmbvM+FyTV3iB917
A9Fhllpfc1aj2HDVtbeJPm60ztNYgAZN4I+VRUlfdeDgYhnjLoBmaPk1WN7PQWrQ
jKMGoBI675dspRQVK51U1VA+ZxSTU2tkbw+S2jEf6aC8fC5ia5nbfs7zwBk3vvdi
WW1OsV7NqmV8TrXerTjy9M+UoErfVgtUg/TxGy9XtGuuhEvhUSPHHD2NtovISn5+
rCqbZi5M/Z7PenjTJ3HtVWOXYq0IaIlZwcG3KvWX/3bOWs1FHe5/8sNAkE82UKXL
jwkEGrqUfRD/J1YqlipmiZqiRmQ4Yr5rtTGCfkkbmD74s6gGIzHYnQmPrGLPtTPB
A2j5XvLhSvO/4MI41osarHKO8f540kxTf0LlBm6RDueGUkpU0aW+Zoi4yF8+E+DN
n4sRJLVsqqCRlK6+ivh5RM1d39lyjpkhct+EBnOcJh+DJ2ZRAv2UV7qWqM7iaH82
G4FVRYCB7n0VkZVGrML/h4Pn8k/LsjKC8VSlxqUN3KDKAfJaCeTEPhwOkvD+X4L5
EcZ4E1pjJbAWR/IU7k/L4yf1umGciWgpJ480rawXWd45H0hq672sUAgsiObRon60
7VjH+4iKKy2VS9+6vCjpWjIo133o64BPxfF4xed4PUWV5zbBo+YxmP75T5WxFTX2
QMu17o53DVqL+0bgBdwYevAFCvfSITYiU9mrQcemqGGsoaE+Y/RFezJ1psffEx3b
MO0iyNcElxk4H9UoH5sU4iydn8cyLc9qFRekUpzQuuo4rR3gZdyexJ3ilogAK29n
Xbdy4lIu8eVXPwZjVIyp5fAbrnB8BklQ4yS2MZYXq8OIbTD5+xGKIBLqqgc4Ol+u
qWK7rqrhIKbiltZmD/dflfhKgwtm5GFxqO74T5//H5QZ1+5NKtMZ7N3ylF0wxufn
eKGALM5ED/IaQgLFEyfVt5E43jWuHyeiDxwN/pSDf4BIIsSvQbp3eFagY9aoglg3
X2HPJhFO34d+OAckJy2ncCRU1qIav7XDBRrw/RAGP7IE2G3eJjMsyJMnB7/jpB9Q
JrIG/3vHCYCH14mO+FOVktuzwKE9vZ+JPmYY+nfz0WWeniYSDln6WdPQlk3rqF29
gU4g5N1GlY4EwJq17YKx0LCSyB+toKpTQrxm32vl9mdpLtqDq4pOnvX1IPsbrE5T
Hk/xqrZx5+hZjK2i/5Wz4DM6ivvTBbFKbPMGMRqa2ztwgqpiQhduUJHYmOZEuXZW
H1Gpemow0U45ED+kFGhZDhRRFjU04grubclkFfx4t1EspFRNDJo9Q9xPj/hVfRzY
/L9MnAFmPdsn+DJgunqFb/MErl63YYpYkktsXnAgXg3oTvxo/9oAaOgZ65qPTtEi
mM2RLoTzKhaGAnL5+PbmzZW/9+tFhdq5zLICynX00EcSZNhDkwlWSEWwtmk0nHdZ
Tv2AKsFAzwrIlBlIvPNr3DHd84FQUWX5WfDVJYM807ih7OMtAp89Q/rZme0cCkJT
2YHp4vV8kwuKPv3w8x1RCWWlsG2fv6r/3D5mxEljgd2nJjFsBatjZVw+elUsAxGS
x0IBFFY7M4qB/Tv1cxEUUrf9Ft8CAT83OUs0K+T1lVdMsdXs72rQjjVTWu+QFGpO
eWKgbSfRLGlidHtlfQ4+VTmAmSDWJmWuSJ8oCSxgypUn40OigjOxq72pXKg+YAsZ
j9rTRHpRO8/8WtKGSSUyEpL8z+r9qAIytp2oIpa3JBK/3aSxyk835V44deB2NhPv
58tv74OKUgQd+K+gICNuECtDkPdIFhHlpA1qjc2qwidDnyke3UeVjRXbdkhhOYFO
pNnRL9Wv8ByMAKINEP/3ytBVU3oqKeRtjykbwCieh5MaNrQWc+afVuGyvzb2+3gY
cix1rII2zywKt2pkUT2pfoE9jKgMZJ95hsABR5QYkWWvn4SLj0+oWgO8+8nCtOx3
qCz8QJ2Qb6TY5zLMeaHtzrYpUG8obX+533sQev0X72HmknMx/RvuLTEii2py2VvP
wx4tFxQohPnNi++zmZLx5I/lo2ARyofKaorawYFQ3uAu03IT6UJy67BCfE1mvhJQ
q5lzz/zTbUYN19JSSObab/qYvASEmLXK87LnnBPDdNwsZ5PB1OEIo9LGQ2dA9rtA
JaGzdImoZ41tBz2qQN52o6ZeVED/d+zt6N5M5+QBPqhdJaU1E/D/h21XPOR7VajK
u0Wsvyls1lTXrLclQK5R2cj9V9C1cADL+3HLBNv85Uiwm8FhsL2+0RGE6Bi3CrYr
5gqn2tmc2j8Cp9zu2fneNq/ITvSWEbzTILOr3+X24wwd/Eolzf7J5PHs8r3P7LE7
LfHM2QDpTm9o3Lx6FLsuPabsnkbHuAGRW/lb6gBKoOZVnmnnTjWdmowaSoRYnpfJ
tNqoAOArd75TIvBwl+TuYZkYhHPjBseR9RrKe76SeD7E/2b001ZGyGZZc4a6uKHk
y5jG5jHYNWAPa0Fxi+PZ/DdJ5fxIb0MLntkJG1TKfuwYi4QdRv42x3YUyBLYoPr0
P7mN8nI4hA/jDFjPdS7X4yA9wU/cgR0i3efRA20JIAa3wvbvYzuuv/xuAai1Um17
Wf+NCDp/8cfWDOpuief3CWdeL1Ma7Bsh+9GHGyazC6mfe4pCb9pcVRyekCqlMYRD
8euxrwYo+pKpMc7VWGUuyXvRnAv8u5NnFGsKvvhRa/V//6RDEHQfH1fmR+ssM1h0
BrVLA6LW9n/hRGyzjLEULZFSd4hOVGsFQi+83fKORnTSr99XbimSocVeCAcircec
jAZEfXkE2CoV6fVqapSQrDXsFK4W1OWB31//DOzKVz8Gjou3Z7JWJ0kfPJDikgaN
Jap30zusJwrhT7dkjvRh/KNlYVxBxgVL1jjnD5nzRN0zi1CQCBK4FpG+5cwaUYit
8VtXwSl+aMI5bimXDEswhTnnCJhbE6n8HDWFbnqNVHGf6+yTH+ofs8IHzqHAkNoY
GD/NDxcVZ5FFUsxlT+I0hTJJreYCQmNmUK1h9oWJKwjEs/HgoAUWngGQIEPm01wb
9E/JsfHE0oTAhPsmx+kOaxhxTCsmpLzIL1cfkCaXT5l6ZEqKp+dIQGCiPaQT+r4O
QvelN2RXtMmdkiZSnmPryAHhrXSR8yeFhgowG3IW1IdH28LbWVt3BzJTZ8lxpW3I
AYqfCxL03U/4FoxfT8Fy94sR7LXkFis5S9gNoI29QdlfuPPZ0gY9N2uP3a3Lkmlr
+HCRBuo5ipzDrnVhIuFV06Uv5YkeFxJK9ujkRq+2jNrQgW1ha2RTuG6L6eSGpOv1
Mv+q1aEYfU9/CYxv8h1f4ySsBTzVcK/GigAcjLmO1F2hZngAbERf2y5+v4AssYda
Eg5M31zkctHpKeodDGGMGXGVH8THM69jowPSTnbj5ANO11BjSFYMusGy0xvSWNpJ
h8Hzznl8aQx8gmepEwS7mMJKugzuRktxyw8yO33qrfHYIaH98rYkW/wdWWsNAcdM
Sei6UyzFuiW1v54oo1M2OstptIC4VnDGRL0ivQbjr0rrGApfDAS5svtKM/YsxKxJ
Kur77z8zwBco8laZEFnmVFUZOH18IX2CQ1/EOafVrpMO44pJ9OtTee3uM7KVfhjL
Lfbdy20sUF7iTCzu90ZBqGj2gxq5Byzk8hb6zeHxMb7QM6GVQKrbhK7ohpF/teQ5
bQCmJ7TOdyzw/BVm7s09Z6k0KuTWlVFoYZa2Aysl/URBzI1IMjdsu5GqFBdFk8Mv
SAc2vcM3Iz3JTtVgw7kzUUlN18r0Js8naHdpyPZk6A8Yz8PG5D1ZqJdB+eFgtxo8
ugaqxKa1Cjq4nG3MpVRY3fPpnnuDNbaprZUKLCeuwiYjnkI+NbfgyJw1/06c/Po9
KCME48EcGj5UXM2UEhB/i7iKieEtN5P0WP0fcUoNkSTQ1180zD3rXCTVpFjWij0p
/a9DD2DqDOot8w/3yrj1enEAm2ubzMw6ecWfe2c99rpjEv+8GTbrVLolHfwTRZJd
A1hZ5GEi2C+JwhS73ETA0QovtGJl3SSGmS2kOmSi6FHT5qlaZULwChq0M2LTfY6G
e56RzsOtzM1iBUKZFyopS7myxEcW2uaPdJhyB5fYkTy2WVHZXLN4EVLvErqsb6ZU
HXAoLhn0AthPJgsTZ78d5B/1/WYn5Okz8FKzYe9ir4lEHWPEz8BE+08UIjvCuLjL
JGg4DTrFH6DWNKm+hqOepjurl2/gPs1fPL39CFSprqxjQPZZLQsv0MpeWnXee8RT
+o6hShLCCnXb8pzrQDeWOK1AYqNVgnuX6flPa7tOyPhVuO+PtvQoJ+bmakZg8AXg
5nAPDR79VKLS3brD2NPn+wt8YRMLaJaq1b+5PSAwjhnNl5Y0sD8n9ZF6YBh64Ezj
+L0m8u8JxnSit6aFUjp0i+zw1LFnCLGGxm6eOzMHxXd/gCe4vCRFVf/dXtepQihD
njtPiWkf4DKMq6vnjpSEqa6PJ+bqJdm6UzUuZzEYxdkSm9Vdd7OIRvl2yRUz+U2P
mSY7JONbUSwJq0hDpKAzMx9sX3Py5MayUPSfcFAI0/P4WxpI48KN5HjIV95COI6V
coVvfb8cuMddvtBydaI6G5NlJQTlhoPjdO1XKESgfPMbibBbylCOURGbu+z+dkSF
4ne1LM2a0jOLQox8OZLWa5TSbJFeC3WDMxcDDVYUD1nj3ahoz2CNQZ8MQKgtu+mq
IygkX8EIQUH9KEm3yuSrTkc+AzonXMQ79MNzqpBZ8I9UbDxvfx6GlZvzWQ0av3ZK
pyjJjZx+49xo126PlrNBKM9ddlXVuRlRFTouMEA1/clSUZXignN9veQQbHxM8Zof
F4d8sT930UdRzzF1Go2AWKTQTSvXvuEoFcUtniGNHgRSx1VI/GBJi4LNWmxKP5De
mUcARZceFOkOt2uMCW/IHe8HA0bNeoJN7wnCc3YJ8b26kyQw++HjxNzIgexafVbQ
0abcf1USCvyaX/r3Tng8mpxd3PUtaRr0GidfSOdEAkghoASvC/Ool30PHo5471U4
oaSYlKfp0K4jzw0Lypu/exGI/t6Bu0T1LpUZckvrvVl+astihq2Do8TsQDzmAAtY
2F9gfbIUP5DVjM3eXNZIyVUbRtACNfCcKW27M2SgqS3igxBaMOGQwQLt9+0PYF4X
5W9zIojqIlTb3Yl/MqdSkyP/6GhpyaVVgXN4Ojjo/mxFUwmrTgXbX9WbgPxi7aTq
1yewRxOB79zkYfpXuKdudZuo6QVqOudIAMUM4gfhGs/wNmoro2RacKnlzL3FRxyE
2t9axTbtHWHUvxkxzZOsi7KsQsw7V03b5xpoBXg3yxjCTYIEEtYMSU4TYh0iGyLh
4bEk8bRBJc079jGgkzUyOg8RPwisbO0AazG69WoJ7OOPYwj+CtTaGHuWqa/B+vCa
tn3sej0YvPn6QKJJ1q0OTMDHGkK2U8RJrZJn+4tiACT84Dvb237ulZCVran687FY
wIG8S0qmWbGdEIU6Uoul8oER3Uozjc2nIQp8u49U3f24y4UFxVOOZJSuoaw+GvmT
/Dittni2gG6pUniGEKLNVo+kmAufr3MLHg7OOHTNaaJq4+2Sj0+nQLkwyRFGbYfX
FX0mq2UZNppP7nhGQiQNvwiksIkuSS2GAyDiW964L1AESIrWGqxtny96g9qfQYMH
lQq8JPxckhNyetFvc/N1RzVzGsN1sHGOAsp66cU9FsZGHpaWxg1u12VnhjSoCi/R
GRuJt3f85YrDQeYAalArgVmdpMicunmqRah9vvLnjTDi4RCHLRf3RXY6HmpYCazl
Jd2AX7D79rlyeHe5/Exyml/jmWds98bkXWtMEGoIXmSLbi2IJgBLXd3RXqLn8Zce
67ae5V0MX/88B7K1EKhDhgTKFoHNuXeHyN7kTiLIfaY9ljTO4R7S+cqrjIBzbcFE
Tnq4KH3tVYskZgghOo2D3N7qtgnkYTIWi/TsEs7ODIOPVGmM848xg000jEWcnFpa
j7RhtcwbRaGTk0PO1Ia6jyIXyQ0x1q10nh3/f4HSOHtpiax+7gZrINNr+UPDa9uq
6qr3JSQR6V6h304ic0JiYAslPGd8q99sS6pcGkQ8PPIp9AVI1Pt5EXiGA/Vtrh4z
1q0OtAQiOHDTqa7pLjhzNJ/L9HgOcBuHdoKP0qLuicWju2P9bFZmo6AX/fG81PHX
8hym21GDxiaVZEiRbyrdk5yuzeE623XOULQFXdoUCZq5LEkHZWh7XMhrYO+xRGLW
NqHJSiPRIdkXp/NnER2/FzqvYda5AlPVBiDLhtl4veDZXNNZdZPiVqAqE9fco3H2
ZhpcXy8Z3EDltGLq8Ba4jTplxbkCgvfFTBVrvAgqZ1RUHnnT2bo0DGgQs9OEUgcS
lengw2zhMGnqjZYO3Yg+rtWuLQYY/mTXo4/EzvhTfiyMigdWy55wtNwHd8qE9QnU
E1aWrnL8G1cCUW7sMXIwbmuNkh9MUDtj6aCPvx8GYz8FLXsAusO5M3GHzt4CsiBV
J7AQOVXO/+ut1bvjWmpEky6XK6rL+e8ET9oGUq8TXdACDU+AtC8cFl6twbRNPmH/
nQ83h8QTJMg2sc/avkrlHfR9fpj8A2zzNnuFHj8sWmL5EIBVmO5QfqBNu04QpRW0
hdD1iQxPhbdfgdUnsOedu5zsgJefL9A28oDIE0y8h+xSDI/KA4rCNxhQMt2sya9a
rQyx/Qt18bMyHSuMz1NtuZY/x4ePDSGrUkU7zCAUht5u5Fo12K0NwZ7FQ47J2i/J
pULcaxZUWqeRgXKnJbPae+LzL+uIOyDjVAr1HSp/c/vyEm6EUY2m8FkiJPFuWmmi
ASbCqQq92G4IrLQKCjiDXWg5DPDIP6zd0S5V89L5jCSjf8ZuLGznlU94bX+DfEL6
wz8dKOAGTxoTlW8opUw8pHLpsj2Mq114rFJSOPYnsU41lLq5yT+VbENB0XyZ/fxp
VTukAqWlcf4PG7PRXFPV90DRO1iSjqr5RG/Ua8REqhQxBnRTuRcxQFi0YK9kHAz6
2xxM/tJaWjJFrkQquvxS+6Ps5+6s1OAYCk3EIIg8ZmliefGFNjXWLF6fyVrYFfnr
lB5Qz/BZ0AXGqhof4Ra9WDkR1RZwrlTJyt7JW+IfBJstwgs0jB3wJKp8+uDL23wd
n2QWPY3dMuky5fILRr2YWbmYhU6TY+pZU5LyphF0XsGf7tQ1FbxAByfQ8By4ML4o
52WylcLAUS95g+G7otGijrn6IzDz0sjmn3/4joXJ/fJMGs/yB6Y7rn7+RG0OChSr
rjLHi08BvMV35VYTxb0NBvifkgB6KxiAant26xoRiFiALoVs/U6Ag9LH8RFBymVq
ryWJBMJ+ueiVjXqGfDhLkGgRBCHIprdfxdjA8TzynNSehDASTxlskmJIUYN3typT
TVysYymrpo4hysKK4MmAmwMNovFViOAlipCCyks+QPKFg6joQrnpeEn+gABnSLXJ
m8DkTOseqxAoqJSuJ4z6mgdZ25Wi1/FZqzu8HLnF/UXI6NHUMbt6lShkbdNaek3C
N35s3C8ePHVnqskI0H30ql+zr+PXOjHuAIGZ8ayt5Kd0oApRHdBv6n6N91bdRkMV
qymaU8yf9W4L6z+RnyyL+/UMmTHYVgetjhE2oH1oS7wZ8ZEiW71bFuRNR7pZqQ5e
db/ZNoWzoTB6uGfmKmD6lQJ0Ar5u2ts2hES6nYf8Noso6GuVPtrY/uBaX3D/kfWM
6X4X8UtzWZyQUE+E3kU0UvXDU1sXpmVQBKTtvdsYa//UDKTCb+nhLZCzeHL7V5+d
Nvvd94nY9M0GK0PJfmYmi9WC7+Wl0QL2GgFtL7ojfG9x1E3LVdpN48tjwzB/0p6K
HNrsQUBbZgJHLaJrGbWiap3qSVHWuS5HzGoyDm08F7YLI/yZH0dGn6cIWxild42Q
1FB92U1age+TLyxgCfzaSMW8rHzm9FOA9kvgRClsVbHKHPY+vRYW8ccnffek2NPP
X8//O9W0d1J1scL4G50ZnyRBE4Iahc87yl9qVPyv81AoLq18uhIiGaRT4tydOr7C
MlZFLzcB9PQUfv6s7NjCbnmWCyoWsehaxLrqPZhvu7MI9jqKFk7Nvbhc9YqqrMEi
D9F/8Fg7cvnyIHmzzU2TnmPjWrNaBXZOx33EtPYZoRIALVE/nM3fQO7X5oayDfQg
QccjVQP43ffoNVHT3dVqzqKNp/yNhSMfSuuaCxCi93x5YBiX6ium52dNDUSYP3Dp
Z72DxCjNFkZym3QvvKQbqw00EQXHFYBVFi7a/8rWzhHV9dwmNux85eNbs+ueWbbb
HgYQwyLSJn2XywJQhNo1D9hy/E9CQiIEC5v2O9g/GAvb5dgsVR0R3m9unfSbxLy+
nFIIL3Ail7O4W3TZevMuzeNI0Eh0oOIkXlvR8SP53Plml1/VPg1wxHzb8NdUiKIq
Vtwg4kiG+IGZUBjsUl8JBrYo2kCNgQX3aZoQ4AO971ZIdFHiv6CXJhHaIrPxzXDL
Kgd5eLXzKIqWM/1f5f5yzIyBXuk5PAJcZ4zkSGEo+BTmd0WlzJ+EGRDUZxMdJlM4
/cFHZRJ1yKDBEBeFp0LPFfaMMRr7itEbP+z3MWswUw6wmgd6g2+zaEfZunMD0ji/
81DyXnyVsyKhcbj9iKYvke+ZPXrIOKNYQ0nKIDjGh0EPBRPu/GaoEcQBzwIUdjuK
6GfFshZvXgqiAqLJ5+fp3VzuTLKyzMCI8TI7jnXKApsHcG1lFwIa3gHOYJO3Z2j0
UkaOlimfD8BP/7nqK2Ir5D+NlkJsBzqkvwzEsbDLMm9h1Vb52bFxiE5PIWvzprMj
jmNLuqkUL4Xsp8t/xOC6IFcnFi7siCgJe3rh9qMV2nG5PGQRBC3m8Pmz45WA6Zyx
XHJ4eiEllQ5owfLXBncdC2/v0KBnnFFpcyYoucysI0F9DiSg+hkL7PZWr+Ie1/s5
9uFCOjiIw1clw6a4aVS/kuM7I9qq60dKk8ASoUj1BQS5yolau4MJxBTRKhpedQUz
MPH3yJGIO9eJWVKdKZ2s2y1GUpoLGEIpeXfuPOUvn4weC8DQY4zjfOuoQPtGjBsh
Ly9TYQg4AdeYMCFkyHKCPzG3ZcHnQ+N7bw1jl3hB8I7sfcm5uOnfcOqERKPFh1/I
6PuGW6+SdOUlu/l+n4oOFbaR9uHoD3zn3+ONYCV2bwRVXd482FLTz8xbLfRxZGyr
jQwfmPVGWwpipYRqASeZs832CjP0aZ5NMH8diYq0+9vIIGIAAqOciN6tSHc5ea1i
kAO5AWMXdF1uv0HowjKyBaJbxfQgiWDpkgItDvE/LT+2pX+JkKE2Aa2m8+/33Kt2
ItaJ/FaEasoPW2Np7bsnPjSnsVHdIexWDkNqqP4iBWZTLt3AujB193GHFomqW1+b
wwLcbbTC1PBaw3ExxzUIrikJmPEtFAe8XtUXnghjQfP8Q8szptfm1oVShpE8Yf4P
2ziIikAYAVMViOLdXQzV55imt0sLNw1tKOtpQcyPPfDhZwxUXw4FSFNSy7ZlZY/8
RLPSBeZEIFMfvWgkYoGM0CUdlJ1BJY2Bu5jdlmPAaIgG8xK5i7JXZF1esqmvYOK+
FPZDuhAvOY2qWOl5pao18aXFx3C6M/WoufyVyhwj4pNB9SvkXOmne0ePxVZKHk69
/KUgoiq+FI5aK9nZRJ6gBsDSIDXlo4zLrnGMAFncQYCSMUmEC2ZZzSqcbc2Hzis8
2DnC/4cXIZgAzfvM5OjpsrE4RG68k9jE3FJcCCeOV5ixsv0yU7nQ5vWsPINilg1e
j3oabxJweoSizk0UZNFKGT+ZqVp1RGY9ajnIQjocovtqb2nesBnmPKYkDjd/46ZU
9IPnp632qXyRnRWvn9NRNSzW9JfBcCcaxWkOaWRaAuGKOcjUQLOKyuH2O6FuFj5V
szUNwZDBmoB/Az3SLAFfh1+QyCJBqXWC8oT9lsxheICd0PMZRr4dPSBgI6hBWAtG
OsorVULmgkBDta+7ippsTDaZZpPk2P8FCgo2BB0JfvN7sT2rpVU3N7cin1mEzDG0
99e/ZIDvhhsHyQsq0noRcshiuZBgbjWCoANXxj1Iw6M4bhUrazOf5fqc1G58b0BA
0PO6H+Qb5vlPD4JE6RvfnvSTejBus+xAr1XKNfSHE1MhqgRt8CEKRiHLm50ypUjI
C7A8QLexE6W/O//MsXmWIJ946zewoiIOZXnvCvtjELE5WLP1Y0cqcSxK1Lzg6hTZ
lbaZGvTf0jEElBgud9zaQXjT9IpTbakeHYEUH8ETRv2t/Iufw+fvROCIUOgmPeAZ
pMRFrg5p5jU4y/DKg/unh3z7Ti9YlRvTVp2W+edCqtJmEEIHmq25SIm368d3sxbP
4EhfBxxTd5YFR9ayRfn2VqkCCUuGpJ8khh1RFGdeCpWQbRirbjXdWIj3kw1Jo0u6
KkwSGlgznWegfaxaH3Bz1Iv8y/YjrRLY3S7kpMknZ3mGCVemiNxyclBxEgTbuqfs
lxtyj94nnxK9qgdoDOwqzV1dECCdO0w0Omshkgg3+z1wqna/qT4NQQIoL4Nt+x7J
uUzUXSVIg1bBPaFfh8aWQCf4gubuGm2fXZh5pqjvCcjQKtrQuPcu7zSIvqjQpuDj
Rrc8D4ehqyGKdgEY1FktMNyKY7GAqZdgaJkZofycKrzaxiiDdWVvrZeEWZiKwoeh
M1vNRNUWQbbe1hrZ0hhhFoSA9ltT+GSsr90oZVeOC728gr8QBYNIKoZZ5L3xUyNB
SKpsophtleEtRcSHFWFwKY1hJvHSPfPSUOEamRoOwMqKcpKNx9jKL5aEbcgm1c1D
eMBUzAvYfhr38o6iRaBKMElpakRmyqERLVc/fdTpvFXiTln/8d3oHEDuOoxepBwT
jcUv9pSeBAcSzvmzbF03zHTFs68QRjgJVYWV+kPPEepseuYGddVKMvdBfJqKtQIJ
vRWHcv3SATFvMGSBt0L0QTFIveKQCR4qoi/uxulIqaZxrSeiTcR7WUyCvIbLr9oP
8XVrIB/fbnl0NpUFHT9K2hauSQrp1yqoWKrcM8gZXrrHwDDSZxp+500tEu7d5RpK
WYPgYSxJmYMn0kDTh/AeLg9Ldj4Fzvc6XlgtfE664/eEA++RGf9g+Gv22uE6+dQn
092kCu78vC9xMv2l67GaQkqMqsDIBFH5FzIVVGh6XASZDLROXKM3ZyMNCob37V8/
Zm2dqVdXePA1wyef8zut92aE1TD/8gmfmw6lp64y4+zK0aDdOx7d8Vxx1QjGCHOO
dtL3GuCU5znnH9M+qznKQ0gxvH+Ewzq1fQk1MfcZL9thnEteD0XTqG68dPQtJVZD
GD9JL2K29gjeEpDFu2/O0I1dLgLojbxGzYAS9g/F7CSYOprEtZHt0DGihWrh+AmE
evT9w71mpxMyl04ePo7XLWNcglwd4s2C3z48W7p4soBbr8O4vUMPpeGTt1mYZQp3
8cUfUi+Yx9aS6DByQ7Y9On1oPe+ytk1vVdOeakCyQNHMFi4YYblm5lTQOY7rt5my
euMBhx3bKn2zNRDI2d51ZNFY/rWOG4c7wV8CMrqwUC6AryIZDXeLV1dC83FqsI2N
X8Kvi+P8a3PnR8H/vK2pgYLc0g8uHX+BHCu+eJRrN/HE7p4lqX4LJM1qf2f7pLfW
/82Dk3P4CJRZ3YpL3Oj8GzVYlB/k3e8NK0nOAOsrq598og03HVDUxgSkSgPbhGkC
cJ8pM8Es3JrfW4heJt4Oq551deSwmLbQbaSX1pvq//wKz+X70JUyF5ioOJY4s1H4
5WnIoPNFqwTFplnUv2hKXliinf0m73N23z2nFOSdCxGtknFzXmv0vm6uDNDL8hPy
nAjW98N3/BfR65i/c8+MhBP4ma+UVu2OFDKyDxEcBHuSw/IKcrDEkhSv2Dj5GyFs
QOMhu419IUkiGQtVMYOZKOC9oDEiush2/7i5IH1fAKtMMlu6BGzmQvkvl8J9H50W
2IQY0nQyT+mc5YVEOMuTtOal3HLIqZaRySkAt/XwhKkFXVE2OgZ0DpRtgtnmfWnv
2KVADi6yG74Uj5/9HC241YE6N/ldrts5awQ5ehsou1Nxica4pfyUKxlCJaRk5CNN
O0bx/jRBP2kz/KcvpHfd3U5aiBRe+qGQcz/D8sanksB6b8JvLKfkYEXc/zdtOo8D
lGjdZKuZt3qvxoahhH/+W6PScCgxZuKK1mjVR+CJE0OMwAjD8qw9tU0EWbZkkZDG
ugLtSlDMJC4M/Szi9OyoOPYVvDpaLfZ18EYaz9igqB6AbnkVsdmmNcgImCl/hQgP
4BV+D8Wcdz+k3rCJO7jI7s8/vQAc9PdXwUDTKHkFjs2TBHwGV5G+f76tqnY+KQJe
N5OucJIqlhsDuAURzDjs7raP9EnQEV7uLTrdIBI7UHzNX481bNTOlRd2ywXFevVu
5zBWHwdV8mEhBVSlyJ2Hl26WMbjgfLVZ6E01qgwvGGeRbduc322xpr7VQIofmTZU
J2MsjDowXFW7oqAB48oLbQKO+QcvzUKRFf6LgBGnJ+KOCp2moSS03e4r1AKL+7fs
9N1MrVf98x+K+pReTr0TCd94YIehWvs9NcHxP6MVffqz9yXqNDgCdNMU/FkyHRKP
Ji3PTk/8SkJllt7wX0WQRA6V1acQU18JOcf3IWObRpY8VbdJD4mpoiKFOTNZOVxx
bCu1puq1mKWi95eaVb97DhAvY09812GzLQXzvuPBQNFHqlAijujt3LMNrzTns4vR
rz2KbjkKByhZCFpKGP6LJoNsSsMYeBKqokchcicks4lb/EjQVmXYmaQSGcv7IcES
qvDbv/uPjuNQCVbLsfMG97yG8drQ2gIzFfl/nnVIRxMrhqiPuXN2ubDGHkFSYq3p
CVuJEmOGd/glZ6Hh60E17Icp5SbwuhNLnmMmdxRLzkfsrkp71iYlMBQjQaUlMxQU
6jN9g7bMo9NjgHqhT1FhOu1LN2N+ecCiUa8CNmlz9Xo3EugdGcxTC+5TuH9Xb4Il
r4gyap3Ohhho09fkh1SuoS2TKDfgt3Edt44t4n0YoyfeVxxGaTccF+ct6RR3rY5Y
Gi+hnCc+KjTVkKUVhIsQIsy45jdXxFZuou+/Ls+78SwWwj3O4A8tphT+a/XFJHzg
2KPu2/QbU9w7B+VfBw8fhbEnqj2s6me8uhf/6O7du5VGAqYH4rnjgI4ZsHC2EC+z
tTtUvuvAy2NiAxAbFzTjaZ1lJZ0LjoMo95BIbk7bkQlonZb4FDdTeRMViV6cO2SV
EQryUjNIb+wW7R4pj5FjsojfEO2AHI198/PklYDfPGQ2K/yFH0l0zKBHl2F6YaWM
7mupNglBdmqg5QdWHe5vQQfGI6AvgnvoK2XxjMY8pnbSTV7KEZZ/uBNmtnZBFQ1Z
ZI/XuMTde4qpP72TG5084XwIrpNVf1O5ZaQEOu3ExAQ2P8WqUPzE2MQlcv7ztWcm
N9wEQE+GrlMj3y7lO7jQJX5awdoltABdXz2B25EFqR6O2j/VRnSGwmylWjZSxmOB
3RGo2NfUeQbg0gpEZASuwoZvyIkwlq6GiGmuOmkiPWi17EHZ318lgVb9l4EgdjU+
tGYjwXL6XCZXZ16vRPrPBfGI/Lds/cCINiUqW13MiGlWtvdXkBwLAn8GOyQwtMtl
LAzZx1TYPL1I58Jku+q+qoXyUS0NsM9w8buB/vfMNi6YIcR//a3MiQh6jLWax0L5
fI2L5fhVvyYIWFhI61D0tXAiE2R3SFYR3Jx3sbbQv16RNTjHiFBYdiyAkI1aa4PR
yAT+TayrRf1EVZF8VeXEAiL/84tJMmZNFNPzU5xKklrsOU9aCz7vdgZvwC3YLURG
Wd0NUQTAaeT3eOUnyNssc0dOLTHwGVu4QjEebi7Jpn9Dm/kL6CTsWa5AL3YztTGH
s4vxhPrdGtYGlUQVpw2oEtAvk9XeMSfoaVr8uozxWET7p4/sSj05e6GGcLKOorPH
oerLAPsS5LtQxsyiQPEoMzDr1SjtS2fmI5hBunV8h13yYAK8Rx519iGX7Xe8X+50
SOqUq5fGjDY0aGCZXs2vlzpVAnQ2RMjSCaQ22Rze8RMKgEbEsXi1nZL8RTrPh1/m
q+dZUFXkbZ1to1ZszVhvleQvhlgf/7X/2kgUmbkOUU6QWcIfBKje0IKMq/S8kxfj
0IWVDIcHY5U+gZAYvAYfRg8UF30tXgU9lQ/mY3fXH44nY70M/bxK3OZdyqTeJlkb
MzI1mtaNorikRu/1rnbXIEIJEJytDX1i8zp/YxME72SJXst80Tpi1/jlt9hFlL7R
BOWaqd2Jzf4eZY0dwBWFGqkW7UoNhVR6CDRXjoKV+5yyz3s05Hi8IwIEfi30HflC
xdrC8c9FNJTIuE9I1mQQ/ZUWfBP8RY393VxlWpJICIisvyH58oDBADy5K7U5FY17
TKe0WTCpAX0pIft6YNrVxNr6w7ZNr9b3JHg8c99i4MHCO2BuePe3bVyhrGZzkh3w
hzcXMlrM9gTQbbWePfGSnloGVSemCHYE0/9p+Xx576vB1lylYyaDuueGtIT7NfkH
+BvJVkwl34LIXgmAMTC3P6IAUA0MDO8oRCs3ayBb0fATN4eHlMjbuK4c/7L6lUYa
p7RLmtEn0y7XIMU2bAANwkqktZJ7iuOenjOgmuvwRe5zDhnKtmhvtzgXGt0pgaDT
3IywrJ6FnUljuoSLFYeLhkvLOE2pMbsbOQZ3c1lSauZdAhf5nVDl1sPnjn7fu6Io
QcSqCP3BQcoRPRCq57npavHqQHxoAMkjudPdFEiAcLEQHvIcih0IpmXgIZolLfA9
kCEn3xLYV2YAHsixgRp+9qpD59F3GJJ9Eave8qBnocG6ec/PaPuCbQnfoWgMArvg
8Nxl1ue4HadTg8OB6ORrBh7LdJTMLQxm3eSWX2jZOFFVCxNjBJf6fAiEELjz4hl8
Ee2klAzFSzAJSIUEraTU+szBAhSMEB8XCzRBZ3swntufyiwg/nTY9hPJtxjGi1JY
UvxqB+Iyxrc8BAHoMBo3IUoZbzzCLyr4muD9+CheHMG4GZdkXoPyVCI6CTR7zk/b
OxoqWNHtro5JB3lGBnadbjqbxBM3UBHiF9mrtSKc2pxUVHF4HfiSLWFXC1Lo99u0
/pt0IDXPfx1jutYJ1hLpx2gdIrxzHNSFYVsFbt166jY66ZEDmYcFqGduR5plWiyF
Jt6324PQjV/dJ9xUNPSuIZ+NVvNPB+sMqwJNRMIOEN0T9t3zecv5uYwJWe/nqL0N
SY0iobnfcLs6yIWQPw3u/ok4mbElhWytWKguvva2Ng5Q2Q2v1tpcCtTa49mdyEoW
xT07cYY6vxGdTInDyxD7vu0J4deTNEy6FB8GTcWbv1fUYsQi2XqRSUt8HYhzwl5c
4DQoyvVkNMJI3mxGwZ7+hK0u8i4s+LFG0St9U17uI1fr8G92YBk/ZrSjmWFjtBjy
1SeG4V2Dm/QaCjGXngZ2FtA/o5j+JwD0MHL1rZAMGKEhFs866PPfMlgeoZtRyM+x
hoNJ+SyjpQlSiX9KmwYCvF0TxWz3Dwa68zg/Tdqq3G5ckRxlBkVjVY4YlJaVUHwQ
Ii4xrHfMKHofkYobyuuV5mkH8wfBwyvxh3EfpO9+M69IOvdu6//m6U/IIa/9HEGU
WrxhXb7/znaEHRJDvIkesXeIfJWOXHTNr6y5hr8RLz/nk5gsKAq94DT1URPxL+pK
YborpYi4cCDfnuer1oLIQD3lDBs3f0e7P7ev9tjia44P2UCwNNqvwC+jC8J2lxsG
NyaFHz44DqW6tGriG91/MnfOKY6vkf8IKxjpcoVFLlRer4Ut7uiV5Zc5zPOGFVml
2TlbAqdKPgkRbbbeQMf/+Z2jXwFU+k7AkL43/4ftl1D74VjwDqUPyEZHDZgpb71X
XSEghmlfDdXfxO+TnEZ7Mp1vsTzWEAGyoxD8FQ5xdEVAgjNHZbMpf8gOe4hbyMOh
I/Qhl0yMeaMDTJvuPAP8GvsL80gp5UAbO3TReqKBV/q7E78DXuAk+MlxIx7JBsFy
txlZg39Iw3i6VEwYu6mkI8c2V4JSbBq8bb9gqnVjPYvADiQbGnXzaKvG+D9HCHxM
urUjbd3TrK+WkdUQmOmgI0/eX3Qfvlk6MwKE+qwV4ZX8WeWMPzZBMGFzbeUf+Mkd
YSBOng5heT0n+T3ylHugkq12flFzF37R19Y7cqHadmoY+xqPClLqwoDi7cd8MOpi
wamelz6hqBXGnTX+s9QpD2Qz8xcRNShr+Yq+y67tGP/eo6WIgq6WPYbJKiuNzYYw
bcUJxqaushblI3yL5UiyYkwro435DDoYJGqZsKRETenklrBv7Ve0mU3mwl6IkuVb
/oJ/hJe91yorHztDbFrFX1/LIBY8BpUq66T3mn+sSMGHuZ035fXu0hN4yuRltVaJ
fTLc9LEuJSKmBZ/fNJhLT0CJrGiGxNDIx713Y1u+vKWabPjNnwzRhU1YHXW09WoG
FZ2rOla29uFfBvqcpoUu5SsFdZy87jIMD6UXj2W4/mFnppi6Cl4pE1KyW27QIIgd
k4NuxmfuCMsrJfTwo2k8obkXTZfHtnTd/KeqI/kt+RODPopOQqyOXu7I0XZY1aJv
pZU7EExMQTN6HISDon+0fm31uzqu6HF1Uo5A7S0l3y7+KLH/K5DwUHQByCReOFeO
56EgIEgKRCSYPXaemjF+Tj9nOqoo2V2SstC101w4cJhl8KJJfw3muady4EJAQ74m
lpHdfYnsO2AcrEATvC8jbonmxFHCWn1PirnpbBthi+Qs6YfuC5hiYQ2Nry+oJ9+C
ZDAYjrgSQA6FLbvqIB2tb4orjeVOOVd+Yl0vGB9PkQhY7EcxT6utDFx9YhE0TryV
fLZbPKQsgncNpLlpifzFk3uxShe8WuiK8ZMM1UnOnLn+ZHwfiSwc3hv2QsddNrLF
vNUF1hB4cQhC860FzZsMSZNcph40frsfj6wFJ9hWOZEmc3TVetwpFPUZYPCSFbYT
FMvfUGk1Av73goaS5VeV3qoE1bs+up1ifUghNx+6yA2sEjvfLOM1qL8J4NQmov9/
T5eeHwDiBDW11htHdGF0MlXx0vh6cQnOpKnytU5DZSPPoEvbpgCWfTh+Y0IZJg/x
C+icEehRniMsmf87biKErFCngI0Pnp33JzEKNUb0Ai6WkPjhb0SWKJmibBelqOZN
r13M31KzOB/nwrTWmEHGarwTsW2DEuxbct1LqQFEdiVSKdeMiz31xEmcDL9aAbRr
bHE62+7JBt6L+Luil/dRNv84bFebPljalg7TiAUEr45OD7yX+ienZIm6tE3mgoY+
93CmXTwh43v0p+OfA2fimqYMFuyaW8AAZvOjMd5eCO57KHfho0kulilPoqV1Ez5N
FnZtuaonc48wVkIWZ78+bgi4rS6dZmOlahPIG5Fble+9mJzcnhpD4UeeK1x8Imst
MCIgcQkfdQtv4vZTiojyUwmLEu08CccdOTGLZZIyGKH1S28uReunG3MghhyHCF03
+ZlG1XSq7Y+ASWrysG3WVlv/Wxy4zHCjL6YmE6mIlGUoCTwnmoRKSulp+CGOAyiG
GBaY7Eh1/szSJcb0LUEOcmNR6bTqiOS3PqBxy6haUFA5hSetnG5hHeMye4IBN38u
qdxx8eRMSG/fPh2Q14zK+SLPjMYdjoHiA0lLp1yZP8mY+41XuGQH9HKz7fU+f5kB
EDXe/MEBWIhNsaS1DE6dvjV17KIVkVk6hKdYCvkZufFd2Jhfkor1vlswms0FysLX
7aIkFvvCO6jM8R4aCU/sp1XJk9mdNelIQ5qZTtR63M717TWdFVG33/2hj44D1ct5
4XnS0cSkCBiZkxySYEpa0yxXBKUHWVfjoOHW82xCAFNH+a9eBAzziistPBWF1ofl
rQFMxr0SJSpez/zDr87NE0oHoVrWbbEQAVRTVp1eVQLauU7EHzWqM8EBEKmZKdhI
Tbw2P1dx37FGHvBB8WxhV6e23Ftp/+c46Z+HExf3w/u2H3wC+xE57bkqJkPYbvNl
agxSMl1wBoiFj2Dlgz7jdf78nQ983WXMvHoCB4MxxUqWiav623UgcouAFtM6n9zI
9/FJCNE2upaF7JC76dbfBGXl1/rGCmQ4f8Q/UXeYI7LM59/PtVeRo/11F66N+iev
ZGybub+i1Jzz3+6mS0Nzrj1UKEXRsQjcYWc8ug9bMuFaBXUn/J1ML+Rnni3zyqvC
HXYAPmugfXVDdoTYiDlf5NeCQpKZ/rSN024SO7NZfmso384o9TPVAYcr3mpW5qOy
nJK4f3kcstc4tQEGH3YPGm9paIgUffaEdRWcBaM3J/FucseFFcshnFEIyMDg+PP6
A1EcWwYHro89InqlKItnQo7YzqkOBZSTmpYOmX2QuoBhfsjcZ5jRJOFWDUQbmIHH
GXWi/UAOuAcDXZr+p2tA8HFYO1hMNtMThCA764Qz8rBKZ6xNNl8g54UL7kx5O74x
7TfwLTR5LLAI5xYaXMVza7VmTuGkLDQEXcwRlQ5CqA9BxaHIoD0i+sYdPCWECdPI
/SiWM68fJ/vVlvZ8/a7UG6q+gq/CO36mFrB1MGE2f9Zl+rdshoLeaatMltQzuBjB
qHTeK09+i5yZODm0ui0q31n05oN/aC1h56sd+nGdP/31+jpKVBUDOG7pAdRq258w
4OfgHGPb0dhVWI8BStjlnyTGOHSQcRL85/Owei5s7blU9+Zk2iYrDmfiS2DQKZHz
x0oIsnBkBKGGzuKMlxAbjnGDP34MzIx5K4p2AAC1D1YG9aPN5+CK72+i3pV5pcQh
L0UQT12yHcoauxbNBhOHWnSTqB94b0dV+ZwkR0yCkcAZ280eKFoFNwl0t3+jCsnT
UA5Igem6k2KK3g6BhOy/Dh09yqUi+oZXBWkDiOrEywa3BWsZu1bs682ys9oQ2p5p
xzv+15qo1lLl/V6ujgiOBhFI9MZ9E9xMPU1bWRMDfAiiOd7vCT3IqK+qgTHfYg1U
EPO1VCr41UHP9Q9SWklSjExyQ2IlorP/cKJGXhMIDzK4pPsFpkLU0ZX/+twkKb27
kjU5VVftonsgWE1zdvhtY/6KddFZ97dxMjmAR71pV3v82JhYNIpJxKfcL8XttXlp
ewlMPiN4CkX8BqpseobAiBHO/zLZ0E28gvImG+kHHL7BAMpXRyqvl/RMbaeoNQyO
SUrITCraSBzf3PlqPyADdbzCO5hsTc2FIPcKIsxDiqw3EPswWkeq9ASl57JBOsFG
qvmT3OXbHTP+sU3eaw0BxuLvS1HbItuhfySVPsBWbHnltpwp0g3OkN4jMRSb4qm2
50P/WXmlfOopMnSTOIIIbY4qmSRgs/SvAZNKCMTljefbW5AAUUddOQQLZhmhk5b0
6nyYvFilbXoMMAjijuutLZGyd0n0LcbQ2bDvbqI2mtXgnRjm//uTN/oFbbFWRQv/
aoq5rpxTiD8PmrFIUIlI9ErC+ELkw2REHZnTRI8AVFUzbs+0DIBvGsyMq0AkTDg0
doZcxv2b6hl8NTckYEVL6+UKl3rZWAUvEK1d2xsrIoDIuNK+/MLcDoI9PZ5IK6jn
lzHrQaMLujp+j3UJh6AWQQIEva+U3wpZVAtyvuPlAnLMzrJacTYb/quHnfE0lVuv
kcISEhWoejm8925kBKf6dFBSLriP3GZgLll2+gMQEoRN1GfaKbFLHV5nyZKoaIWv
kO80EGg2LzcZ1q+DZEkh6pGOgU87YWhG2Ez88dMakaJbHE7C5G5wdFDf2K45+IJ9
EtCm6EK0cnfLiyrvCTyRGVwfBlmXdxeSC8+lxSosTUNpvLTD/RkIOIyThy1zGksV
sHdv5oC3K0alkUi+KOwXSns+DjgklVv4dVkENxl88gI/2yj5IXaKgOtF7jOktp1p
w2syAtUlZybKmwL196XxwQoXaUk1K7OHt9TeKP+MTiwAEjlGJDcxB721IHqTm1Hs
ge85jRGgL4Q/k7iO30eKoCV9bgU3JMWNqs8InrWrkj7CRLHOPI3Rt2t+b2g8xD7j
Qzsj1HV+sxAmj5jDLtRuNO3/lJ7NMuW1Xv8KXXblBQK+xxns+/22/TnUDhVXwvf1
5MyOOWc7YE8bqpeNE+IOu9f1vGekEx3Oamhyk5oV+eADKe9BQywN5Ty6RwaRVE8O
MGN9cFzIIZg0IMWA5xlUE6y0HwlhpqWojOiSOaGrSncTjG9r2Lco28bSquA5JfS5
XYnjeQXfL7VFnmLtdRg/JzA8P00HCkq8h/xqyim+msTvgNvKIBMRI7fXatL1hwFz
VAK6HQDjXhPLJlf3X8Y+Ov85cnyydUYJKEw/680V0vVY6lcU7aAfc9oo1CTP4kvS
l3xF9s7Lwex4H76NRpou3zBjLvtAfyXRpUOXYblBWz7eSGbpCe8BhkkLD3roXUQv
wozGRLumx6IMNgdasvsoZXUCKWVlheVHH25AlR5NLwLMFI85jRu+4tS+dpAFNfyC
Jp+XQvEfuf1JLwL7Bxho3+izLhN4r1rSSWMj0XjBfpCar6/bT+7c9CVetIVI6dUQ
EMavNxoJ3YDi3mhuH7//isHID0nUJZ1uBWgGEPS2PLYT6sCeDzYPOw4mAsOf73G9
L38YxtkAIYj+fHh6ectzenMZoGI0MEb8KzeIiVfmGbMqDziTGQFbpvUYOkt+cy+e
pM4nT+mEsjPonekp/gtgpYRAvxETuttxucxQFcz3axu4j4ECb+PJVyQa44JHRYk3
wWf9kRLfHuQeoWsqCkCzMncfF5gEXCz3MuVifsmq1Piw5JGCzcWlRpDSTMpDeLnX
kI/aglk+oDHh/lK4EReovhfkWehKiGfkv+6iL/y1+755X86q9ucDgFFm5qZxXvNl
WfyaO4dFoPRrJ1eLcVgM4VRKxYjMidFhsBHbTr2HuxQFC85mAn4uCphjmNh6gPJD
UPtHzPriXGchIfGZfOZUuCHZJtEvAK5NTTRYrAnA5koIlN1x5kh65tAETx63WMlS
KJH9vxHRj/zKbkSSG77enw3jAyEtR4/FHHq8jur5iAmKvq3fRohmQW8XGD7O3sIc
Q0tXGevCTHG+OQ91jl2t1PlcZvzCA2Q42oXkhBts7/bTke234e4KW0CjwhcIbe1g
xOKWJd69Nm1WZSelk+GGhCmxdkyj8BcFiCWyIdgvvo0IFrpfgEBNOCfXMpOqkEED
VkCbfjmKVAbzBoAUyv6dVpZ/IhIOB8gDUGTNGIkSKj2FcLgWdMZnHbOkLB7bLu4F
tRjl0rO6DbpxaZeltkTCPtwo/B72AyuT7HSpFiIoKzeW4ovwP9GVgvI9b2XiHQDX
ur8eBBBhUKLfLwTuYiInwJ9b2lGUGL6wIch7wmeUuB9zzWC7/nQCEjTD+xARkXrD
y2Su5xokbMF9NvzMippoCW1BdygJ8D5t1lBTwHxauCEqNQTvfiiNSUe5F86Q+Y/S
XOlKZjMAIUUwls2mIG+UE5jN0NvjKI90yKvyD+Odd63rQNXJxYssXSlxAUItsPKb
CaL6H7rLH7QtTNBoyXJWzv8OH5WUQlSxhw6ZjeHwoJT0NAPMGWn52cZgWA3q0KBi
i1DAKWiud4XQtdtHKC56KmJBx71aOiQrFVyITL0ZW4H3tBMsRXDa1D9o3qPYE2Nf
Wo3XL3w77mSK6tTYjbhsPZo+J7w9PIo6AcIYdxV7uNmlo4/P26h87F8b2M355Gkc
KLyV8+sbb7JuzLXld8jBt+04SK3yQdgS6WGCgj6wiPNILBoNSMZrJQxuL1ZjScHg
Hc5SAqqJit/IOWw3wb7DP/BPI5apUs6YhXVU+eu5yPbCh2EDzrW9XcHoHUTk/Qxp
n0p8XRQ/kVc2DMCUc0fK3esCE/WrdgvbcaB9WraEzW5jS3Vq0L4Pi91DaSR3eNJh
zeQh6qgEc/OfmYz1giRyxt5Dt0uT4EZ8r0+0gLJ5OIb3gU1xe6v4JJWFkf7Zo2/g
DY3Kw6mmLySKubw7dIW6yEW+O0s7I6ezvzrI5R5u+YuEHWvyqdc6dW6RVKWe4IUQ
thxQDpspe66uZh5M9q0t2rnG6IuWSlZAyiFEKapiwYBabGxwQu0NZZw79GJHFdg8
a0FshkqGWQg2YPG6YNo6mj+kC5JcjR3LpJIHu7P7p6U4kApnR91artauOZFHJIW7
yn0+1rG0dgqg3xcmnTfJ/arXVku2zKkb/HKMhutja3ezxdTdJx1CZ0Ve/Pa45JyM
gC4lWINi5jr/NPvWd24zwCM7BwCK4Qo92uKv10vuJ+TnQVxz8jB1r5ErEqWDA4iz
kbYbRQe51v9hCdyFUAqK5bx7zT6Ziqfd+Trf9F/Q16lmRJRYV30gmfJkL496QSkq
d/2+TqNsaRBBD2aJP9mI2Q91HGamvKzAp4c+4DSkdGCjDt9CLiBaNzDUI/0CyS5f
eC46mF0MXr/Z94SEfZoT4OAGxSB5MN3fVevk6zgKe2m+XHe9fxqA58EcoiIoTxq3
Jo6M8SGtEh06dZMLali7L8BiVgr5IFGQjUp1iFzM0T+9GezX+tkXaaLRKM2wg0qq
P6tPcqM3uY+hjV4dytT/DnG9jY108qqB3kbcpZ8ugbG4uucC63UriG5e9A9eYG+o
3okbvUHbgkYHOhkyigmqUYRl0ODTfFnH5nXUQxkH3OV9eLTKVD8F62fFbp9KzB/n
yeTnkvVColKLZwqwHkq4A/OP+zBefKn+niBBW9g6r1kzN2fMQ2CF/q2OA0nEXAZk
S68yvIawVTdCZ/XH9XQz5xc2ydIDvTSa+Yj7fr7NouaAB6bX4qFWCluAu8kbI7so
Fa5lgN4jtrENoQsSkefcD5PCefE8h5Q+HRw1irz3BaUycQXwvPCvKFTPUylIQaXF
m2Yzk1DbCnvkw8rtK/1pd/bzYMbXWbpo5t8k8x5s0h+6z9YwYtKP03eaF+Ic/vK8
hJW9mA0rg3EXyBSRNbCc07BhfiUmBSVJd8FPLJcNdBrVnok1okN/+EDu/YVL1YD5
VcGRtBSXjJEkiNGGEu0xP0F5hl5yhpI2Eu1gGXw/U69D7MzqLy9DaVVSfDyKINca
3N7g7KzQCAY9qTK+eCBowoU8aorS54UGQ4TYYpKongQliRIYaIHF18e+tU/V8v5n
wVnsUFJan/GXSRQycExJKAUylCh5o53n28Gz1C9bbJn8qEXWrv+4sqkJesUq0kJO
HBv0EOUiekqCtRQX7qbP6QoIFQx7GYnjy4dYWhLK0rwwiZztMPoXUiSPIb+JprwE
6UfqcZqlFWn7PeSQY+kNf1P2DlEX1K1NP9lXaBiIYLfG+6bJdom1Wbt5GUt57eaU
LjYiG80cNbbklYhTEXU4CJDJOVpoQdbYtlH51q7lxAzXiXMe+TpV+nZxS/oSta5U
jy2RkyQbZRc4iVV68TPmfEG9FI1j5cjcaJb1B6iBPqPv4bPJSl8OIyDi1mImXkpK
8BpcagyOQTBwcu2Vt9vDSLKbFG/r5sl8VxzKc4mnzx+VV82qg8SOc4p70cgZknzr
dOL86Arl7OtUhyZO7cX70FII7ixMxcl6iC5mZBOjlfCOF1Uy+eoiRRFDXJlKEADY
CIHhRw/TrhyXNS0B5oDFtF6SLFPD5pGAgdvrb2CxJZRDQPAzmCL3Rfdc1bm5DfFK
DGEbpmI8/7VTgzV2HtgJiLWDBKBe9bBr782FN0eAZ5pd9Ygz+FI4VrBanL9byWof
I2+LNFPPGJzSTn5ReivsmEozOew7g3y+kBwwt3ezjn/85zONYZYh8TWSK/MSowcg
bfyivy036MfnhGa33eSD1ldC+6jeu38BUtVg/7FnOAV16OLnEgBmjO5FiIZzooCg
xFdCwikZ5wWBSFDLD9WoHGPAGeilbJu0jGbBi8Uj2AD4EodDx+F0CN9XwurDZAla
tmHxSY+NL6ytZEGpAI+wUDV7mnH7YCcZKmHfbDpLQdjbg2pCvrqqoXLod6ah6XwC
2UisRzF5w0BcRkDBDg8q1Vrs5Bq2fLyDZ9Cmhol/QcPb//iZfYDs7YGfnuqWbiys
1B3DTLWo7Bmc9sgCI7mbh1Ra7qNI7hKVD0/SzTzBxai64ou14uK8ULAqzRpMu18Q
bQ7grBUEHeiKHIhrWvfTyi9lB1xJ30TEJTvbaPBgesMCsQhb6aKbSCCEW4gbKUV9
4wZ1RYmLzqj/eWqbSpIGbCk8adVf02tJonW43vFDEPqsqAAW+zzCiA8r5+JJKeBd
xVNo79u3kzYneXelliOdPzjbyIxmVyS5kVQiXu7ZOkySX6jVRK3oXrC1yX9tL/AZ
4dJ5WXbwJgduR9tMx5C/xoEWA+Ljb0AnRipRwPYcE4WlcOaZ3MI2Zfiwnx8f58Ui
GfXyecUh8gYZ2DAqGdx6jtNrW8DzyamPOfDCtC+po2KSRWHvd6cjpaO/D96NI/SI
drOlBZnBIUTnGCfs4Qc+MCKY+SZCdO23zSciTbZ618FkzAw3C9Jwoh5rLKUiyS9Z
BQKBeGg2ipFaqzGUzamAqpUp8lpSNZixTkOACnPkg/dRfWEO47K8jS5CL+PM5e+9
5vYo2U3eaByrvWBHyvCyMb35cUBWVfJferqmn2FCU7YIvgZ2hSsloS626/Wr8RtJ
ZyrBgAOVXjy2ChoHswK5RwKcpwoljf6Xfq29X0Cr50VEWS5mxGatk7YGHCev3poA
8qNsxv/MRU+dZHXycfNSULap8QczkobF1xp+VZrkCW5KI+K6EUL4NJodOMRwxBLK
aEaNr/TxZo2sbqA2Fm+wijUFUBYFvF1kAFTC7xUf/W+H0/+a2h5XhL9/27V8uRHM
Mrm+Gzl9kavIwZpgIgYfs9k5w/kp7t5lqpQlOSpna9DfQeX2hXtmRA4DA0y3BYTK
LLFocHxC7pSALpKV6tLmRkwXHtMlc7CuAJGroXExfH2OC5SEKYGIN+Qa1RjkjP8e
axRuaAvFkfZt2XeROJZN1fA82xXJL4uWTYW7h93zpTTiKO0F5IdBrHVcT2RoIkkc
S941zIJ1Ch6B5FRQ4uJGj6lpyK2BE6xaFWuDppA1cmycHWkYnMCEOQhBHhNP72Yx
6VesXNvO/9OUMHYIf25y1qRtoNI5IWbSP8b86r/tBYf9xTD8i5meSOHFxygma8FY
5LccpZoJ/SmHLs2e7spgYDQ02wZ1PS4/pOq9LSU3S/B5BXVpZKTFthMvDFQPdHGf
zPqwSn2E0qGdx6CJP4FH0CfNLtDPDjW3R/Lx3AdIL5U7vp/mnUp09ZEiXef7LsSF
8m2oLA5IhHm5JmmX6gJxoqJqDpTiVnNV0CKN61eRuo9RWlesHOmRXyKWyWKYHzuJ
fH2SR+jsrGgVA98/U42KZiOVS5YoE6x/ta0N86h205R17R7GJEFjNQB/hyU3e7yH
oNfQXci8fB8xhwCXAG9WHS+Ts+jIj1Za0fYcwJBUxNLFkxlWvRUSrqRkDGsxPuOf
6DXG7OG1X5ka0Ek78zQTP9TjQgr8kLomFwcTe7rJU4n+UmrhhGHGTjfUaP1Lhn0i
fM2Y9ABa4LQ6GkqyPpQlHZt6RtUinsCgrp42LMA2TS/1R0l08lutTu8F4YyK2LQG
tnMBhpQ/Y6rkpBJnzFtk0YsOT4z5Fwfevo/C++pLA/icpULEWt0xxHPxMgG+vvxP
HKEjygCoFKiS77ktXmWnJGfFRIO36oPE+jze9LjD5EMMN9z2v84V/bc1vbk7s0eT
1Ww+qMWDovLsGyYaeOSHkxnfTuiRz23ffflh08l08Z+2Jsbpz6m3lAf9JJ4FINU8
zIlL6dJbFOEVnq283N2WpxTZBCtX2xrqhC/ZyV1J3iakCi6EwSEil/N6YzelUWvW
XK1aS/zfUvADkyCUwIFX5uWEsDLP9EaW5nvlaGywkG05olPyEYY1s4TMVhEHqW8p
37m7HhhxiZnwx+GpDNpeyGykXDuuXI+KbYPmyyLuN6gMVNT0bXKBjyb9mbT05SqZ
2/oVmE7+zS2ok/XKFp4Ppr/6yO1W00b8gDy2/28NGy7u+ih+f3u1nlarfa7Fp3rH
MDQXReSgi/Xb2BQ73c5YHsBHFtMKgK5Wj4Z/TmtFbLepRvwQg88sbjqTj9RRxY2V
2lZkkgqGU9Ji+BNclbYlKBJeC08fPcRI4fIz1FAypwSnsitiKHcGMoMCJh3u72BU
vhi/l2wKBg0XS3qirXOG6t6xzjoTQgWVzbKoC8wLL9dZem5GV7j0cxV4078uad08
ur/81hEBFvVs2LlwXhU2AJwpo/RG7juTTg84HCQ0Jeu/0WxMZiheK9jinj/VuMpN
yLq4m/lzei5x8ixXb+2qo4zsr3g1X3j1WxK7Y6u1WtoWeaJfbOXLCf7VPSq++iNq
gYZMLOsz/p+P9vcfyp8f/eRbYnKKnFX3/SFjUJaGOB9YbBLAhcvkroFqIeXDI/uO
SZpYNEKhA1HbJ3KgqzqioBK1IXltuRDjceaUWzr9QzH8LQm50Bu4xFjfl8PnUegc
Qk5B//jd2xKT1ddZ+Rz5WLygGyZLodRo0Am/qiMGek6sxS7my3y2AwR1PfBOb9pl
XONoa4i2XBzsIulXQGCyLANmlSee6FWwW97TTWRJrVOh6Fp6KD3dZP793m0JiSZ6
P8Aj7dcadxcySddeud7C931zQksv8Lq7BVi/5qsAHnblWfMaqdXU9bPDQCXs+imM
Kh1R7iJqOW1D+F1Dkdb5Lefr5/8dm6PdcPVmhAjssuZ5NBFzYDBi6sdX/FXmBdQS
LMtQp5PMLvPCv9hOHYlDHlRFDbLuLdK4c2LNhd/+CfBpLlqeQ+TeibveW1OZcsVl
FPZ1ASBfKaxqKK5iIU6ioY8eXWMlpwWW5ICb+wsI1LsJxHtgY8BZHqXQ+it7Dsp4
TtPDX68wXQjSva2f+Toz7/0I9aOYpS+WJ+0eOZB5QrCTstWCk810Jv62oUInwr/H
dRsfe9WEBOPAh2T/d+lgga0eHyBv3KltYij0oqWOJgdkYYBw5nRdxNu+M+rmkEdM
qYorXwUmrWEhiY2CRUqUAhvMlA1nkgrC0fU5slIn4GH1iXm7VMKWJBvPv/EPxpmo
Rn4qexU7jEN4jXexj5JJyOy7KEwHxw2tvnHFd684c9+6yyEG3rgxvp6kXXjYqSkR
8QgbhfRXs6bymhYJhR6m4YpnnMpx2JRYSITPoHwSnuS5ZOoQpqAVWAwmSmkEXjkZ
so3UN21t5zExLz8Fy5DTbczLlog6eElJSYtJG7ZNZa1yfotY+SoomjiZoXGFLn6Y
CwkYviCovflqzxVi4vrZVsb/aGhM8reskog1ircgWMk2qV5K7DfLcngPjF0xDJZi
vx/hJQ6jMMdWEjOvjDF258VoAl+Nd+uLBMCI8pWl8VHuu5C4XVnhLgDhvUA3zXjW
evT3QmWxwBvX/m5lJOuycCfoCs8XSefIyyvyW/mqO2CqAH/J/Por5ji9rXjfjGgU
+F9l9E9Y8JhZv/dtJ8u2uTtW7UZ97UcqEBvw1Y1o1W4f6qsPbkmurJ4wd2V6gJU6
OhgUuf0cQ/4Lbkt6NiVBQtY14QOZrth7F4pIpu6CiekIeXPL/W7eKMsqoNoD9SyV
Xma3YbzfhvmFJriiTuzeQQzVT90erRKSPqD5YHYG22HJuHciVtkoNzilCWOindWl
t2oL2Ri94D04K5bd+P9QYfYGq9TeedLSIz1hHYsRBnuYm9RqArQerftRFLLbvyMc
2XRT5mb9I/cFieive7ctc7YfkhqFuTwJUmPeSy3Usd2eY985clNm5QAWh3/h/d0+
0e9TENUyAKQbuzrpJZaEQEMi/Xu8senIoplbdUUou+vnaCRgw/GcJqg8Z15J9nlI
QN8Fu2Qht4sOxLoWn342sDzTMK29OkcZPp727sA/bkojj+vxN4RIz09ODZl0bQQV
Gsswm1WJFLKu7V36H3HPUgwFf/IrZW7rRtFbI7iNfPAQKJnbSfjWKLY4U3LL6EmI
zQvEhWLVJWSTxM4OuGc8MG4TaYL4Iln96ll1dlcV9G59koQwoKyWl2gPOD2JKLKU
SZoCcOSrhAH5RHKkfkKZdsBO0NKSkYauOjiMv7AQ8ylk/soS6r7xvKoi9J4XdUeO
vCb50TUItO1kHUBZnlfzS4LRNK1PZd9lvYlqJwLpoP6CX6J9nWpUkfmj6ilG5uW9
TkV3FWxWS9QQObk1sxreLpbusDT3H0Z3CBecKzP9mMv9hF7+VXf57ARPvSl+GGDT
J1tNeNAfRQbv5FeS4CR+A1pZVhSe9nFN4zjD3momKpzHs1UYYPwB2ntJuWmJIWJN
G52krP/nmAJi4bCN48iEib4qKP4K97T6JIvKz0ssLP50qINvSp3ag1vCtQuIJQuw
CvKwdMj3TAS+UR2DI6zk1RPXvn3dE2KQ1iXqIRLu79PmyjDJym8bN9QYt6KI/gPV
ZsogxZuwij9VCD6BjgScsNdOi0u0GbALO6ATVoSzBjP6O2WDeSp2+WNkBAaak0uj
9qd0u2To5dtbvDy4Gg2kmrm9IW1OLXMcuemfGyupFC9GxPE+9ryyKrnpoH5cv5D7
KB8mNdt9y/OYhBACCjNKybLuMbO1m6IelKKjxevXt+/8/vd8Z/ieDVw7zw3U2guO
0ScFf3/8haNThSsoWjF+ogv/u8hyVXLAJsE3hSSOOuAiaA+DYIVJgv6YLEWWicXU
AfDew5O5glTiVX64v46u8uO/irozJQmbFLAK/5u86AOP5ODjIToaPv65726vRAcD
UQMu/1u7RUwy1x+TEQqMxYYidp0RJKKWc8PQvJJfJEuf1HtYUitJnwNq+AobW4b1
hDzQSWtFjQgF0DFLCumK1JYxG+d1fSus8ryOjOjh3ilAOCsLioSE3FZgBruuD1Oj
XSGT5gbmpSMrCNo7frL0sz+ZcY+ERHE7NnLw7bhqT8m7XahlJ6oxOUl39Ge47mAd
ykERcEMGqIUy8BueQuigDV4McDkKXcwzcgxwmmeqg+Ea2vxQAeScfNhEjNMv/O0I
UHrDVi4uhO7cC63/2YOh4F+UM76KGvRw76q4jAUCcs8NV91uO4W1JmrzC8OYOmmH
D7rcF74pKpUxtakEvxM3Gi53gIO3ZwH6B+fy3xYfzjkw9TNDZwX1NeSLXWqNzSY0
IKjVS55/g8r8zKMMOQ3ozvQJb3UwyzFXXGbZDbT54OFYLPxoU5mpNZe6nS99v+gG
yFubC74AOda3B5OGy3R0JgEfyqZI0WQ9cl+8Su3Wz9Hd2LRx6Ylu3pPDNzcdES+Y
R/h8wZ0fyiYn88S82h3mmhN4JFGBJ70trcI5yNDhaJx4LTHZLQql9MSYWGNzy10R
fGap6AXxsLUMfTeWdXu+WCd4xCC+xHC9BCLp01Cz/kMjqDA3N/8To+fuajDO97Td
zmXVyMrTpsULLjI1+HfpQOCgkNG4H+yP/LRtaySYMRo9CQIUyysFDkdCOOgHgoww
O0cIuxgl61o/bo6jQG76L+gqWjE2zjTzWaWtoV0MI+MnNpZfn6XJGObxswbR695S
hxcEjBJF4K6QjonxGPo2IyBC+MdOyzwKDyX51bj68FkAlVmzFPDtKinjz65p8XT3
O50uOL8T34mIrqULOXo2boqZBAVUQFRrbr47s1gyBFP2E/E26uh7QvBsrZ/P9e5p
rqiP5gV7XAjrLk8O/m/tv6UYC6WqEC9sDQAnqtMOjHOSLOq5u8iv/+k5MrehQxCW
Fl6+0H/ZIMfb8lBTIZ3LY4vcZ/bno5k5KI7QQ4oWOqnW9nXwc5CmoL96vaOakZCX
ggU7nOXqyuDIDU+Du8NQtdH+a81SiZcB7zo3Pv++evMfMTLS4/YRp/YVYQTsQG9L
IpH2I2F7PlZ14jrCQq4D1wOOel4Y8hHqY9gID6JFIIlT3Y/y5bNuCDCCdFK6l8F5
g+DczNkjb29RbFX+9ewPrMhxagS4gWUNpgQbuT5+LiYf9TDo7xTIIVJZ04ASEthB
xjKrW0D5w867N32RqLFt/GAe/PUqFdwLsAd8rkYC2V/YQt2ng4EDqOvBccAk6P8k
K/Tmv6mUvJbT25rPqHaR6PpvJ9E1kCrdUsRa2R+seIHieJbtMErNWzsOlnx2KdVF
iS9HuJrA5VJfC406nWmegDQppw9Zm8LSrkjXn379+OkUyDDS0qmY6RKZQAeKWtfR
Z2Sgx+qINr0Yjz1FmLFx19iesTkpAgOYbe9/ZKzrNl8H+sSkpbvUbIZTti/xRLTg
0uYC+ASn1dX4Jxa9iAiO4HczVOi9TrdbtrPRJpNdvMut4K0jDnJBMcmXHJmw29yX
IjReev8DnApZPliOxfmuI4he0TPfaPHZt2S0I+Bv3Z5LNAiVoPj5afmZD5L3+ybi
MgDdZ9BDbHsMMuSv8FbGNjAv1jDJ2DQRUtsPY5kGAjjyatzme3wuSMBTwmbA97Aq
AEv7RwZkb1olUCOScH3pQgV92UuE6XSW/a7+EA7sdmT80TW17gCtrTcVCrREeYH0
W1oulmBKa2SothlIHIWjiOIs8+W+9+C9r4MTa9KKNpz3WdG6gRpQrkUaPGuIRUDD
AXqvJhAEQ/wW2KKrlSEnoC0MyCGOnUdnTZvY6gA+ryBz9gLRmhMQXFjYuXeC1CVw
Fcvnnfklo7N1glbWqfMzaZw6NQBPiZPuTtbRlmR0zA7iPpKfPPk1aTjuSCZGTjjE
djPx0BTEHviwd2iaqEPgwPKBzpZ8zwGkX+xzA0/42DDmV5YahQQhPISI/jwE6R1f
TghpW7wXCxsn76MQlx37nTBEz7Zrew2iQ+vPhbIxYCAtmzYpwNunvfToHA3Sh985
+Ul7evnfNhBqdWWNiDQe8pFcDgL6bd+PvoRpEk58jlDFdOaQch9NB1nmOFOk/xth
87j1HPxOjcOqtOGZ7+d1jD2KkksfoLFrEPPmaN0JPmVFeUt5LKo52UyiNlvuKL3x
+b1tYf3tLmCZY2qg9lTolFHEYaOaFEBOBWodE0v1nCVXkt4RyNVIEPcBN0hKhsD3
H+S8Vo3pemx9nCXhHpW6UOjWUQeP3QUQTc/XsSHXZwuuG9OBJjbU6n5LN0SytxlQ
oqCxlNyZGAS7ECJIuS1+FzoFi/vNecMVbfPw8dWAHsYfhzPtTC3Q6ppeThHFNzsC
iolWpQWgM+H7p4J7dtRegGwi7MR+iatqnN6MKfywUKKnF3qVCE9Q7uCjMLLvdK1Y
lEo/ooHgKkf7oHlAcv9hlSZYti0tty1tUXrujzIGycBIDYIb3KpYNKU6cQXXPDxx
Ml/I6CoAgY/39YjPC/WbWSvGFrxu1SUW7fqdbL2WWLiWJZm80ZrnNxtT+i7Nkj5S
YeB1bFjSjEvHq/FEhB+pQmLKxWLcRe6MBjfVjh8uhrL9QFGo7sYzDuN/7iNctOHJ
eeau85F+aoSu5uz+gZ/yXR2GRbGh7UXpdfctBUiBJb+k0xVghCh6cADMls0V+1FG
d0OgQU5UyIDlub9ww+8X1a/TjL+tnsh5SlzvRMBMVN+zB5x4XdHijpX6+wFzoVGH
duXzhkebkPfM1xDk9qaBTTMQtPmOnI6hjG7TwKR2+8/bkKCCGSeMDCy7d2erRWH5
os/3m/u+IJ/4ELy+01QFWu4WtbIcKgyaLQbg9pjojnwiDMOF7ItJLmtMA7zK9uZS
qvFNe6BcGQ24dqoFQaUMrzgYF31yHMZdKpMWbNHzPJk/fJ8bIi5DRPTqAsOnoiIa
TlsM7gZFD6w76L5bjOUz7sluT15vWXhg98h4mIoJN8MUFYReSyXXL6t/UbGqXomC
a/PI+ilPAtRf4uvLULHkyTneuRF8160y3Ndxt4tTBA/jjnXWJ4caGIuyVpjwz5Db
aTJGAc2yO7o6odXpm2Vj5m/EL6Hqdl5yy6INBgHYsfg0HoQOvoCj/t59TwOEk4uf
jRMC8YJ5QwEseND9WbfwcWUURVjUv0J0j8PT+e9oUgfKE8ZjWV8S/B0zlu/7i0x1
kSc+Nsp+/rz8Oq2v0R4oDR06Xde5vsP8YQhhgUMzWmebvhCVCjqdFBXkqs/FVTe5
2F9VpHMTW9vPelVTB6iyJrdZuzosQQohXf6TNLdKz//IRp59lDUZhy0Vq33nayfQ
rEBbgNraeomWQ1tBWZsBykO7MHRAOXWAXG5cJUPz3GQmxAzYhiOFfK8f0X5g9a+k
gObCogOceDvaB0wiGE/3jo5EZVdCL0KbIaycu06w6V2mHu5/Hgni0vdo42AE0Oam
fisW9pr/MafjhwcKVOCiHTbz0InFYRu4G3vzV6axW6o2LiKSIV+QHfIRjEYyMiAC
FobntJfubRqKaFBoaxPWU6gCGVcMNBGVAT0rAyKMQH4Eni4bzvGQe5llwMR8WJqB
5LnKsO/yhRk5s4r8bip5DKO/2ACgTlGhqZ9jvZyNxdG+BCKJoqv6CWbdWxa5WI/R
7ZKqaK999OHyIJXnMlgx+CCsrUJ/59iY3cMpNBwmyd789/i9je6XEhdhe2D0OGgE
4tDJjVAtQznCdfgTnHE2SQx/BMSd0Sno0msDPnvRfvbWIkXeAkaPOgqAV0PDs6e8
fheuhng0U053livn77AZDORtHzYq0gcCTldKBcqWuk0Jc6JBl1Rq8+gi5ALAUtBu
mNk7PBRsSkFtXpCthOnQ2M4pd4gIPmxW2Dhkp2ANmw02Bn4NmPkm6RtmMSs3n4XM
v/B4niIDEObr9zrshL9B6RygP/rAnboysNT3419bcdP7+hUFAUFbJp46h+e0pezW
47fukOF5N4JbKQYL5+b1eg2Qdaz1P8BWqi0oALmO/iKPeYe3sEtdhCiJkzewD8rK
4ZIQrb7NpbSGMxVYDfwzyZbnvdR+TJiVQY2j1EVarpDbed+pO3YXP+uxA/labnBx
80iWvbMe+JNnMqcxwWG1D3VSLArazuuWGI2alB1JT0O9Wh+freELa+W2Va18R0DR
iL87xRjtJuuCNuUgHF4fuz0Axdle4igeGdne5IwjLY7NAH/GxIEfGKZxZCaEpd18
TpjzcfebHpCaJsqFiMZTr8mHDul1t40fQYwRjIf02HBXThiSh5j3p427JQ3UFDXm
ZFY/hn0Vpke6555PdPohP6omuI16dCAo3hgpgHkoptNxVgW230IXekcJFn5d6Kmr
s8qsPBzfU7Iu5oc3RCTTYJaDQZuKoSfkljqslbDqucxUbNqGn2b1GYQeBmFeh02S
Z5cg+fTvafHR3wtO0l6cwwkoyVok/yUcDxTmfamqoy6R6m+KeX7jx9mj+kqiIiW2
wiP2kxR7alGwLrBrtZSlYmVIvdoon8YI/qjRY4jolRBKfEUjcm9xe+nikBq9MbGQ
1yRWKr7UmeQ8JOvEbb5lBg7Z43Y4SqXK1+gNF435LoQguJhiK9iEFXWafWD3SknX
Bp+NA9ohBS/l0/DC7K7ub8Xb+EYa9XiAeT66AEhMiJ0wZfCgKgOkYP2WSdl5KEq/
SxOUh03iYh6vvtxstIhoPdjVRX0/AEctXEMXThIOqjRyQ/mE/50p9W1aCq1flmL2
3G7lZhH6YsZ0WG8BOyrx4EzHH0q6VL3GRlOMtIj/YO18dFRK1vtDQcFIUPZnhVj8
5avyMBKaC1lV9apA+AyChiEGbngYewQfMBgQPQG+fOxILQnx5Sa1Qh/bBJP66zRF
9IY2+qDQ3x8UhcCCHXuBbhcd4A4i8g8Hk7r+xk7GXcpoolJfP8nS1PkfWIRjNQXP
Yuvru8o52IXjVDD5ZgXX+SyTnXteNHSSsvmALsMK+pJ/DQyn3zumByqcaPLebBMW
YKNJEu9HG3O0DKn801HzXpM8FWv9g6kcWnPGcC1r9ibUbmT3OYkpsJaZcvPCVEGS
J6d3zNogcgKW1fTX5UhhZPkWjlxRy2rvn1rd+tB77u6GZ5LzeZUB6BTtTa1THnTB
aML3juzFqA5FrKg2wThqeg3z3UwA9l+LphBRxnZCBVU7i/FJJ//jXuSWFXqB/ipe
0yCCSz9vKQS5vpRhHimO0wXL0pm7EBzbP3Dqjtsdu1yHS3v6S056CpXCXYkWpb0H
V3oREmSZ2s6XoulbOzt/tD6JDJ3kHtQNL5sWFhvdxS8MKt9DWcH1KYqJIlx7GyBR
WLWolh43ZDilo/wucyeHR3wJfvt76IHXjkS0yCLApz74CSWFY62sI2CBrnQvV8zi
mytRe2Ss6r3MwevUHzdqoURXBB8ea+PaOootYtSrsV4irvVGHrcHd6GzQs8WNTqK
fiKUpJynuTx+GzWYiXRlsldxtEIwzkB6iPEo8nIi7Y0AgX/LumQctT88Mz8oUt28
i5lq6hyY7lssQsVIUQmtN5TgHT/U6ZuWOcw+KsMG5wVip8MamUULjpvG7P0ncyzG
0kftlbo5D94aufDAC754xrO0kqptozXc85YmqvzjrT1JEAMnWQxKwYZR5/6iq0Kf
XUa/XKhJ9p+dix9pGU8ZjPMdxOYbxyLDM8HUabwdShnJ9rcpeHtHK9Yzhh/Zjpgg
psNjgKkRizYzUHA74P0klE76QZck8Z1kYDFQpnvHwP+c5E6BfNwXAoSZkVesiCd5
Z+IuXFzwaf0QQUvtFCQbtW+wFRT5slrhSnJCf6TwM5ThHuuvWB4kLV6mQ98VNFoV
FExalJsM3fZqH6VtYvhyghLrqg9fveKalWajs6WflKFbNkQPBPCR8Kwn0bZkqjXU
nj+SHZzyFyxygp36uqRzLrOiX+L4+Pux83DqQ8O2t+5BEoZYgdEdmAkRbVJdNWOG
xtMw5mfJHtgwEDSnzr2wJYYNLHMbOTVOnNQ4Avm4BLEyUs97RzGQU9xsHX9hcuPH
rGWUppZ6QxPZPQSnCGISihJndZMbRM/fYdE3NR3IHsU+ldiWM0mmU9ndwUr71lIM
zZ8QDqWJ58MpPEnSuujd7KKbI85X2iAfURXE4CYKLvf8JAYeS8T++DGkf4cPYglI
prqLzt7zh82+7C7hnk5OerDo2H6V5/ovJ3EfmSay6GBseVu2eN9VfXlLfblU16eB
O67B3cVhR1H1t29LqVZGs1n2YYqDK22eJQ30cNbHq9JX6AMb4qA93Z0ZjJNL++pJ
V0f1TqJLCF98tAmUhlqM44p1oZ9z0m/4xdXlJhLV25N7oDCR7beKAnhFr1k5XHDj
sbDcoaQK4hePCiFh+sAj4iY4S8SgOVwc+uNVwcr+eMjERWFx/NEASMasVZZzq3ed
6sQ7Pd18AZJgnYOApbx3AeoBiNUbIM1CVs31dV3uzpv1y0IWOjSMafnXbfzJbIiX
J2EOdk72Er7oXOz5WnTbxQyb9eYhQZDuzeJWINL9uB8ec/LHRqr7KB+fo4w0DB6q
K1h5dHRb8eJvcqVa95krFENZDdmJuE59WFH9ULQq4DhfHoEhymybwdhpMdeLRQHe
gZny8YBPKGTVDqQDuzA1lK6jKb4QMtstfnTbMxVZSSv55kycPmRynLx77wKIWQor
aGMjAXoi3tiWNekZfIkKz5WBC+p2LXU5+Y0b1enNzo20uUn758hPuiMqmVuwVFhV
j6n6soyZ3+oOO7dNLoTA9dDXPT4B7P5/j6AZHpkhziXbtspGpRUJSE7MQPPpE/3H
agcA1opE+pfPJulXSr1bbGIsRoXoP5cw60RpP2xragkJfoENoxp/kIy74tJD4fY1
Vt/bun8GAXmQBUtvHI16ZITpR7z+/MHEhWNBf2QGZWYiM72lp4wLFMh3ulZVSQNk
1g75reJTSYB+X9Dncj4eY8+fUrTVozKeNZZQ5nl+ex/UrKnuUZJLlk5lPjIYjDKv
Xv2LW+GlI92pxuRyjNNAgfTapfYxWrubMyUThSm5SxLxU0k9cLxVuJZdxH1hAwA6
SnZOwJ4dW1DFcOKKtfHsSrdZqqqITj8WnwDzV//aFib4I98gM6rXaF6m3GM3ZAZh
xNIrODz1Krqjiy0pbvLkm1pIGdhEYJ2BJbEHkvV/5uCGfpdQkQat9UBzDgzE1a7a
VoW7HDFKSLF8TLLv7BxwKQHAJhKvr5sCk/D2LnwBGyKBEVACxfSmZzRWy90yGGml
iIimld68ov3Bm6UzRKbiIKds1LTDdlwecwGCaufLiD/XFXagzY2snvelkdSbpobG
1Xrf8dBGZooDIHAAKTLnfd/ponXMqdRHNL0NNlOk2RDzVjNNugXYBGiBiPJGGyEL
rTMUYwySu2oxhnDb28hi9sy5B0KhdDfOHx/FIsBIu2Mio35QMDYNnKQw4oZl3TgA
1YtH8ERYCYjArTBkb8aebVRn+Mvt9OxZ93v0EjVvhnukCGqXO5RnsLXwM3O54Txu
2FSrNJqxZ750C2V8q/ujl8owVx8JdA4S7Kx3IYMa8iJOW3rHd/eEF3ZgpaPaZ5vn
kbv91r8DjiEpT/uUklO1sDDYitDxo/p6kqAxZ9LbbYifUns6XrmUnsgPvLqbUiaH
FcCFl2PmtKtLVoZYGDaYgzzBGHCUcas1fFO4R9dH0yGfgHHfz/ZMt1JoJL/mEz/G
w+kMzddqAtkU52r8xw4nW06HTjMEv91+k/c3hcA9rIc3vrjrS6DVVrGqu+9x1Rx9
3MJFBbIGAMy0i2zGPj0HUF4uMqq+qZvNiERjHfhHG4j9Juyy9dTE5LQrvlbcbzw/
05akKBxJIp8G0C3oZbUIilGkozyh6Sp8Q3mzG8M/m20hZzGjxo72CEcqEODrLVM6
U7Nx/BXonYBMbyCcKxMAMgX3U1K5sJfi46vmWr8nBPcA/FTR6BX7603XoYVJo4Nv
cJJRw3Nk1RAwtzGPRN9WAfTUcu0inMjTm3wLk8+bbCnvRjgees6F749DcYDbHtzH
Nof+QoeD72xkW+fasRXnQ60R7CO4cDeboWfrSJgm6WGL8qPOZ2zIL9SLd5EyBL2a
Dqaj6RjHAdfUs3PN9chtr+nobGTwAMCEZNF6fPpMr4N01vRGaH23jadUAcmYlUKw
6gv29PsEyMYQMHg1vzS7d+yWXNtlnL4IB/NN25lkk3+k//RfZTM2TD61wb/UIOw3
PLgsf0icAsn6t42C8w7Aeflv0SOHVVbyLWLsqDHzFrLlAGEWBAllmlflwdSEn1Kj
+JUHSRIkC2db4SklI9w7aQ5e+U2pUCTghzKLh3bG/UlrOlAy0R0rjOT8u8IMf/rr
I3ww4vHkwOW9e/vVKl2zgyNQPpnGFChuqLy8oJVb50S/zDdOhl3ge49bv/5aDcMn
xkuejmd1h/KuNn6nAE/lUoisUNdzsLNEi4kepHgdjeQ9blBujX0diVpaya/uxUwN
GdCFKAhbDevLbO5GO4EUBgHSO1EL75Rj0E52gLerKMiXEzDcYOOWTzDoqHw3zKxh
lNFg77wEYeK5FOSQdznRhKUzMtaUXpYcaT3V+O1mb6F4fS3klcT2b/lv1GttrvWO
0kll5lirU5F9bcAwWwsSv5KCey9qWwrPGKgqn1Z+zbKe3ulVrqvLn7CkNg7060/b
xnE4zVQ/nX8gFiZNgiOY4jVCSIvCGUSTM6a/vwCSTO7Uoos0wkBbzD3tcptclqON
uRKOixZASy0BD6JfeXG35Wfq0NUHZlqmmWNKGGCdP0sdgObWVgAQYMt4W2CtWGa2
rHa0aRRhda53ipKABiHJGU0a0JOPViGah7trs8uGQKMzLSbE5rAuU4PEtwqQBURA
Q1VEsulTwZ/3+lSB08bNxjQbu57cttenHJ0HFtrVK5SKVIc0r1t+MTEQ77C/Jff+
RcurzbaHk1cFfz5KxTFXLfqTh3D+MbFVpieJr1OSHc7bIDkFs80Gran7KSdjH0xP
uKIQE600+qCk+Xj00eDi5bU4Nk/Cn/wT9oNDA83hv7IjcI0xlLsfKldicOWQXhsk
cSm20TD5+8/xLmrRyqJY884V7comVTV91zD/QsdJRSkTDgWPryhriugGKTbnRbwE
KKxNaVqXgEegjzMc76bNqeFjCHBi2hgWmK2lRSte7zpOe00mweY9fSzfCpMSCn4l
vyh+QB6j9XDz82MT3WOuq3e6a2fsp+NR0zBiI8Dnb855IKc3AEWjOjmWBPauA9si
smgNBI6rSWBwyd7ncEeToPjIDzyfuV47uvVx5NppywqF0bDhqCNFSlIX9Ez90xOO
dT5GrgiNCMJF5yn0PD3xGT7ZcQJzQk9PcQXnRC42gjWwzxZELup3ZqoEAj2se8Qs
/bJeO9tMTtJO9jltW5Ku4Em9+wvIVD6+VuzYnwp6rfdA0vRWebwuq5wcWnJqADIV
teC+/TIjk/ZlvWYgsLI3VeY55vxogqAs/JHx9bArHgS7paP96lW1DH1uX0Y+vC9b
jmveb5keOvbd1Xbg68/v4HT/p6ecLjZnVeObIlWUYQAEd7QrLEHHWRoi23EbWcr3
EyAauIMin2Z6UdH40FZr/1jkd2Oavob2RCFCVxIPjiVQaL/VoenrkOBh8jUU4U4e
jA8mRcuuvKmZborfT28F23za3rJ9oCVuL9++om6Ql/hNdNwvjyMdRzOCf2HOcbr7
fyEIkyUMwUW3vTSeBkTfAcLN/HyKZrOpqDdyE3uD7p/EXQJRvD1AST1BhWyU4d6/
+55PaCQXb0R5LwXDmcrZMZ7lHnTGmUNkok09RAfi95nsnNdy+s+dsZDxZrakdqYV
ON0sGhES5/9q3xuClZWvJpdmX2ruwK5VBCt1JAhEwnPbqyfFG1uA0tKfNc6hXGjL
BTS1gWfyupjSEjfIGd0+DU1NIrV3ONp80vaF+VYCKB5uBDbYdLozpw/rx7t/gkHG
crgW/wXIvTUp26v86Zu2sTqhqcUqZtmkZERpqT8MvWEtkqa48dqWp0ys+shef9aJ
/fh4tZgcNVQLzHUdychzjQ4/jSDdZPt96htiB/ZJpCyHN0PkyKjbI2Y+20vZ4Wjx
Zm/Cd5rONf2EDqSdX0PHeA+AHYCiSuLpgaN/Tw36WG/6Mo15LOUB+hrcfim5sSYY
krnVLxQNttCfKwT3UmGJOTMC+amAGN2e9Y9BwJ5mwixq/ctJO+AeaL3fhVmLte3N
5+pnxxKS+CGvCtvf2ZH7Y8la7HIKnLc9W0AbGIlu8ZjFGLTpFgr8q4y40RQh8peo
fHssnOtfhpch50tbipjtYDeSt93eTWjcSbpSKKHnRfHROmp1lKPAYluWmdaWUrh7
do6rCbvnVHYuzExojYuiys6YR1COagzV3W193Zy0aRUemG1uPXJGz4cGwyLM08DM
K1qxYeGcti7D5VNlzkqJwLVwP95Wg8hcHkF3svySvO9GbGmO88SG6aRNPlsckunD
hQ1gDm45DJVcohPFi61C58IxtwceYTcgX72J/XwtuUoAj7nxgpuVVt91BoDfXqK8
1FzNTYQ6Oo36R8l9FAZBvTLYlghFaI19sp0E83NaryBmQGTCwwIDmXwA844JHyyg
j+wVVXN1UMetaSFkgV7Y68zG2bVbvrfjEQ1dNzbmIFdUni5aiPJqtKdLNZsh79GA
MENiTpG+yYs/+cNIZou0uI2Hq67jJ3He5GPYgn89bCrEP1brtsuv5GQDG/QBZ3D9
vj2R5wWGztRfwbf5D9RaolVkmtYB+zjdzrC2sxkdw6R9I0pg8b2FlHbkBIaJHY2Y
oWbBYQ32rMSKGjpY/25sqlhBa6JkFESOcjuHqGKMZsMdrdoihv6DwYPKBfVRQEYV
tc+AQBnroPS+gVyn11LXNcbdmOErTLW5RDLR42pIpHlrNRu0WN9u+lsGBJElKBVq
YBNi4WVuG7R3WnpbssYcHEMcHYn8jUZFJxBPRiFAtCUa3MfT9u0j97tnW3gkiUrR
w+Fddyhi4ZeJ0IS3fw86nV6xb9J4HcMS8pJIZn+udr5XYVsERQLjDlWQ9Ms61KYe
VxhguXrdHkm41RsUkMcV0FFu2gM4r1haKrhAtrzxTM53lA/iy3+c6+snhw8mz5cR
/PdeQBfah5Y6nmlk6YpqVlhHvzQCeTGUZChqjSY18rFlRK+KdMvNcZ5LkrYw6FhL
CDpNO/gb6XADiDG5cHr5ocnT0H48mLejamvEOxSA5o0sMnWzA7+fMuYm9rKZj23q
Pc1Gxe+onbDR4LHyDXWjj0cTwm1u1dbRfzU9JMWTHlwQOogoIPWPEoT/eDmU6MkC
/NJ9BRiOxjQCqov/vwgG9Zq/N8DqhzWvkh339YwsrjJZ4AI2dBn24g4pVnbA8cY/
OaRzIsmvGsjNfSWgoCZUKdgtHUDL+dYbKLiCf9i2qfkctu6IqsPrV2pf1y96lU5I
v3veEd0XX+iMeubehK2TRHnMsUowB88tdsbutxBwB7ZjXuOV3XhOvqU1YmcPOyep
66JxzDXJF6tFjp3PSTzVz67+YqapXqDvm3izPfqFn5iP53DgiAKkB5kL4SjWgXgC
2XuAc/DvrYhzQU+vWHCAYrtkzLjjf8lPg28qtP1C0ebxR7fAAM6Uz38BnxtIllQj
LWCpEtmLlgONpWM5Tu4gejxfX7j0IMwNq3TY8Rfxcjb77+rdVLmDJXQOzTNiaWxk
LwyC8vQ8BFHhmT4uR4MqKmWtqueY6YF5t/8lL3Vnkwup0R6w+knweDT58ofAwAeM
eFXUam0E4b71bioKKBxjPjce3Rgrf/Ak7mCnc3SSSMw55H9dRdhkl0+fKOVKMDQG
Lv2HO+6MfNd+WTBFHx+0xtgPbNKI2JgeYIioHG75TkllS5I5I69LXogi2Zi98ZVH
bY73/oXyu4THSYouco+MI4r1lfRFTWgJWPKthb3ol6pW4C+diQKqmu3Bb66lACjm
hW8CZg5uVaQfGhWh6XjUQwj9jqpL2+9B8CL9PkqSNMLpU/f6zzuuLy//3BBnj6TR
WlPhm7RrZZyuwR0hDnntC9QpIlSI3EPs8Nb5Jz0WUra4OFmjoo58+AITg4ZNZPde
+Kniax6Q7JKFRvd9KgFp6Ocse3/uPe2cXsd8cnOtz8FM1yGP+ZSefcL3uJ9EKqCb
zDWINwAvtPm4BHP3k41EuhWPowkJ//NabWdWDUt2cRXksDjghWlnB4a1o1pemgSP
Gb5NpZ9pPrDHeFfHFhtmYGsZKFZUi/KA5fZHnCaW1ZUjBvn4TfxRc8CvSKIFoARL
KkQs3/AxKlYSR6wM9g+PWa8RKRMALrTS6l6/ly1NPzuhV9qagR/IFpxc41RBuY9A
FhKs3lrIbdwCGPR5+TkTnDkHoEcrBwbnekZNnDcoMxoWZ54DwTUmZeicfexTNS79
LWihXX1jQf6XR7XMY/6XSYGDt964rT1zX/MRUcYYjdGy0TTiiLR70Xi8DHDGkq6a
AKxCOv9Mr1LYOkrdIIHPUQa3RHBHQUonNETTfggIMs/8JYEtPB9PDqexLkRMVjLI
bZrhqHu2R2wreJmm79WUI3KYMc5ozI1QD0Vw2sPX/Php9ITxRMJNu+wmdal6RiZA
iiO23/scndaeW57wghs4JJJS1ApyfZ72BfTUXLn2eZkwbEbChAHw3R6ODi1aTlrX
L2rofgRSzansEHSD8OvwDlrIIJPNLGjermyY/zlPhq6W57Vif4aWQ1Ca19dhgSZV
cPq6mP3Js+ESEW4iNjxL69o+SnhYPL4LZS301cMsprl20Uih2cY/tcskKlsz7QAQ
Imgk6SokDVdabrJiS5R9MgUpv/gNaNkOpBuxdxA3SIt7fXqTJGdTWHITBENwbENi
r1IcorIYxnVvbEbM7dG/a6NEeNQ2BeNFTLvLY2Tjk/jzhQXwVCcD80tQ0JkAxokM
BnwK64Y5tXvSfgjYMK5fnmosLv8mIPcn6rqiQw66QVAKeL/tZAu3iiPamfoH2Tic
H5cnkoaZb0GNLVDPIxmzKFuznA1Ew3wf06IsYNO6LzlscSaUEhA6+BPoJa7M5iDC
76caTrq14uQN/V7lt5bVKK45Ko11Uev6+CmVZkMV2tn1hwBE8bp+nq8nepIg+Ytl
HSZcTqfmdq9rX8pvjjoj8DWLEjxZVpipGZRY+P6l+x9E+s09asfsbTHLHSAEykFx
mJykPLIDekMfaTcSScBRJ2Id+S6PgtjFLPVJi2L/cA8MzUgPbz1OisuhSltGkD+f
P5dmgtO5pTdOhAhxFIcjIKN8D5S18D7f4pbs7FDLpZ9QXHTOTo5bts35Dk2pyB4D
jcE/IP39E/erhuWUQey6VmZ0kvITc3yQAZWYYn98GfcytL98ZSOxLLZ/jPh7Hbzm
q8fjs/Pb2wPr0rLymfly+H1m0AaAcHsNKT+B0NEbY5mhvKvE/Fx1QJgcEquE0ipm
/v0fbuykzHrRbJspvnZLwQyhR8TD0SjNPYMtJ7f/PkoYgMzwOtxeVQdkz00lOLNg
qS+QFGE7ZYJ5CAotQ5M2csfisDytuCTVmulYKDRlyjtLIsEw6PEvWaVJdWcgU+Q5
gVzPxHo4OW7FfivWE1eIg1eC0BY1nryMfMPwQn8WdnabP1fNcyFWqdDstB56VtXc
I1kqEbGnFiRSKo4qmtHBcT3HsbILIcJJGk2YMAxaHB6wfNuonPynz6YWmacSYRF4
ba03wndKGHfId0pDAzdY7IHA32LQMFbaDpsyubkkVJGR/ylu8XP7123jw6BlZtyw
U0XczZgvztgGScgZZQEUtgQHYyybTFU5gS3zjxK6J95Zd/BePQkzLlnfX9eSrHMm
PQT1Xelt3UCTATSW0TYn0wY/JRfRg1jM77HZd1FvN13cv1wfttVkzWYYEo/DMI4e
9VJgU2joiECevrJ8QCSbvkJn+UkKVtXYSYUT5kXRuiIKZPKrjlmKFRmJRxEryUME
DIo4Htc8y7OaGcX5oonOZy5fLUDs2gRJC7VJ28KdzP455qLeI+1zWzQhN/8xVpIB
ohWFATJWD0pRYLiy1qKVuPTEqhIk51SlaGmMNn5mtIN9hEClBlPpP/i2fWou7eV3
2vBunkavhDPqXt6foBDX0bs4vBnsvW9dh+1PrVxJx9P4Gq34175Hp4GtXRD1utX/
zFD4YjeXzNzGX0Y9v5KN92Bq3T4fkq2x019TPcJVo2tkh2O+ul/zmhwPLzX0/Vzm
edqDMkh9jRUf66sHigNqj57uVHlLJp5mhHD2ZtWUwk8CE7TqRk17OMUgd3PfgDWE
DLs3Y08r0jYFnm1vJrrYapqAqXrKhn52njGggdhPKmdF28PFh33vrrf0J3H+VEy7
MNZ/iGxWddVQv9BqqMVjth/PTaXdxyXdSYaNulw5kQCxXpsqRMw4A2xTMw8MqCw7
i4/GZZaHIW+Lcgb9yuokC9oe3qe2KsJkZW+pN7QSn2tAWx2kDquV9U7RwHuZc2Ud
oyP3cJ5BAbObD4859jg1VIM8PRcsXCGNL68wQJXFVUjjDnzFgRWAvHli3xUB9jwA
nHclxmZsXGbJK2YNiDl0FDOX5/fjtIBWTuH9pHQ1lpgsawPwcMoT25qEJPxtXSld
0vRa8XP7uGOQGxziUlKD9T28nmQzgca3BySllsx8mFZ2DywdADRdEmEn+Tc+l0TX
yYJ0TzM8uz8HVM/BdfHdKIakBXMywhOPpdzkA4Nj6QMztsrmAf/5i0OC+MeH6csG
Ul4Vp81GljuPIPwJoFWi/V/14HnCawKbvIzyfmzMSLEkZS0Bt53ZHj/roOMlgUEG
5pjyee8CxtfWc8l6OcZB/3JuAVnbF2ymF+jNkU/0UXKHceRlf3tlPJ3bVcWgJ8PA
SJ9Kpa/paTyPqT80SwiTWelcUnWSPHIiWTZ6td/V0UmmCankT84Tj9nuqWaf1hgO
MjA2Msn6GTaZyp/jbjgR96YwQZWRiOAHTugy8XwtiG+n5v/WsbEyJS+ukD9HORjp
LPcc3uBOj8mxwT7/O7w6uhweqXx0zFjmLbqWiV0jYIa1+k9heGxw4ciu7yUJ542W
7s97TL0LhKcDVeLKvrxEPreL5FhsDdoYjU7TuleTm1uZQoWCKDNXns0rk2MGb6E+
tGVtJfHn9di+aNbdqZ36/f8oxCN7h6YGZmR/7dFeYcZnKtbAtrR4eIUi+guYieKa
9/WlJos8rwIVHrxI8EwGBo7u3NfJkSdeEsFfg16Zp8JrcIZHBcE4vPDzl7b4yz4H
8+AVL7WF3x9MPYvqWWjQ8vspLwSLsC1smYjXUeK8MLQ6b4ubdflTJhy+OB0Mftpn
xkU+nu2eOaatZA7OCs+PDEtthpNMkiih2R5+qFBWAfQDjov5s+rnraMR3FL8kZfc
z3IqhWbST4RbP+l8zugrvyaruoKRX1C+MrJNdB/klDlss471gTaewSBGSLfmcTyl
iJBkCB5uZfYmJK595WqgLJY1dU8cSmxSz3Fu9VTer8iwKIUYl3GqIgzoPMLX/DJc
PT5SWQK+HzZpJH84MOXCc1SBjzGgXmnWhthD7sHsZ91ILcwhGFHCDCzM6VWiLxRK
dYcLXkt2eTFVrYdMFEus30nJutr+C9QCCYRwTLko15EH9Y+ilxxMKrOQf108rLiH
h2ldvhOSJwtSkbG7zY6kECpA3IMvDb2bePHl8tU5FwGUqtIRDnr6xGUKMB6DrI4w
z4Xrog8f3NDdwHyZW1f9GxCiPJHT/0WPMsEToknKq8MYMlKM0aGmOc32ULMkfMEC
qawFo+asjw9fS0060lcz7DnGuIdtYr7yPc/4EKpe+4L8+PX6NnYsR9vbU6KjNK2F
A3ccc4kWABh4wqZqlDLNldgAlxMICf8D5b0OrsrTIHSVLELVE2o7tzgScbCGgQWm
1flUdzp/D7V/Y2TnnTVYsFBajxF3vMQwXjYp4oRQlbOJSadPT5mm0xphrcXi2k30
QHhrjauvbUWBOjOmnVPN67CHAaqe9YU4bIs2W2icnh3m5JuiBFDJahDNkfnQR2r1
3TFKr8/Nw/0Qh1hzcG1hvzVE/iK4RnVNEFiJ6v3Op29n+6SremdfLGEQc21Li2Yo
kqw144a9/k9FOw/SWrwo+y2BsMHMTo1czkaPFg4kIYZCsyU8NifNz66JKXVvR5Aj
8Sx1HQOe6izDls5fXoVH9l6+vcP77YpMJgrHrrsaSX54zO+rN1+Mie9KKiyAMcub
QCke8jem71Y6KENBKyVQKChVZEsR4FS31mpBJ1lD4xgmNpuVXuN4L5bVnC+O+Zvc
u6gHEPtOAsxAthoVjgJTfLRflkDeYSLCY/W5vNBSIDSr0cTh8XEKVR2D+hT+dRm1
6igyIvsaFfEwGK0d48fU/XMJKDV7xUgTfmFDMslc2Ntf0q6i0tfyVOR+L8050Vw3
XQFlUZslGSzEMDxP/QM4vB5j15jeUsChDQfFFWuBKhsM6ZqQhss8Vbaj+dpYqOM+
vIOLmBUEu7+p3RCwgVmjBEsbVf+jhk92KiRSO8LrYxH+yaNx4H4aA+X4B5HJxcNI
mEVXJ/ArQrBkmVkqdEfV4k75q5QkoYBg6ymU77e5gKGwLtj5JE6Qi4zN08OtprEb
y703juTUoWqhGtRd55m4xpF1i3cMKmT6U8fIyP7q+AFTxLvO+9cCC6o6vSPVR+XP
7iB/x1RcN2TB0oN+q3A82TRWxsAB8UMX1VaQ6h8WyP/JX9YDwzjFYamVMyMU6icM
B9/gP5yfgXQjqNlu4nU6C/Zsa/pUTI7SMH7ex54m+ddtlg2F467oa6mfzaCT0+ET
2SgI2J1nGU7WwmiCxSHRoTiB9sBx8TUJ29oaQ5cECLKU6oFguv0vhC1YcuPbfZ6r
cF6QRXc+0BhSlNKn9SfAboyd0ZQ8u3FaLSVgBdtRBWNZ/41k/7nmP72oxILkkWV7
Kf5S5wWCy8bDQlnjIVXzrIEjgnZp8XPj+NrpFOzNyU9y2N+iAAHe3a+j8ADcR2ue
JmME4Po1n+EXgr5jSACDnm3R9CACZEmDE5sl0mCq9ask4xPP84c3Ryl92IOgxFZ0
VbtjA3bi4Aof5UWBc80oVs1/nBW4/Y1sPETeL6joZ2ydEBcT3RIPlPXmG3Fi9Ii3
SYe0jiWx50WNKyqtFss5VTEr1bB9kcEHkt5ygh88hegNIWxe+drHMNxzgZJODv8Q
JlFzR+VuPmEiiMoArOZVhdBiGpAxT6eZhQwahM5CAe3F94nPE+XG3Cgi8MoRJbWs
mZ8LThIdH9iAP6qxnNEidYyZV1eJSFv64skeFbTmeZuIFYh82oLrp9zW8mEySstM
KKc6vQz/z9MFFNWGb00dNoUiqfPyyzLenxWKGGYZdXeGT7cgXRvmoWqhx0J/PoUj
3GLm7z4AU7gOm1J04kuIIqWvzsimwsQlLmgquDglm7iwaSxls5TDbmpovOF3AKCs
BMgTMOJV3lpHtsER7MCaG+LS8Zyaqhs6SHMor3HnYqBrZz3rqCG50xoc+JzHUdwG
+KkL3JJzl7AHHWzl/0zUHb0Mcc3PGWFsujQ9qwOcNGrZI3coJVKlJyzs+8/SGLn6
jY56FiWy46A9YSTfgOc+EencBW6Nms+W6BX8s0/xTK+uMn153VpYKQuPGe9DF92p
XFtcEQgQ9sqlCV80DEYTYDuH+BAS5GsZz79geVw8Xb4V4k7SVY0D2GmzqGdAomrk
XVI/PGjAppOGfS3BAxOOh2MTdzAV6DBa1fJ/rl8Avb0OBfNmYyOD31FPpYO+cVLQ
fcQFw1ffTjRRwxuhUhDE7C8YDe8JaNVoL0CcWQTuXmghiLsupkdd5nCd1Vu8civy
Z07XnQ9xG49IxTt+NSSh9dSyiYsERMwihLavvhXr8JRSrfJm0J/IF/h5PJ0NZ6hd
gTK8oX0KLMHYfNMU3LFVIRHZu0GzL5bz7NM4oioVK9afIkmfnhwyMiFgLjoyriac
IbjA2B2MliKsNiDxYGARvH83crBskW/P3Yd3H0Fy0lUKpLBW/UWmrX55BYZ36+D+
6y6C944RSBBhF0nOy+OjnMhpDvkJhU96tANwjDZKbRxM7eMc0CSRnjPM4nd8eDR1
/CXRjdkKwGZJQBG4NHcVBmSzPPxcxkywunwpfdXCN2j6DzWwIApyn1nIhZg4t867
dtjKlMoFNbv2YgqT8S5irlaH2yrhjkrxvGcjm6qqx/+PE+wYszijxQ2bqG4JzhBY
c7Nu9ylWdEbzR3W6flivP59OVsAu57myh/54ilypOBxiuzH09OwPHNwu4jpBlbUh
ulTxtw6rfQxKRuZXhPQBRy0HWy2l6pAA9tNkastuwBzD5WzG4sjlLcqimL0KgWRG
MvZmovGpQXvha1JrNHfGPqP25uL8UXDcKs+tSJAdJWYPZhRNSUktX5xyepH2coXD
1px6AIDLSTdx+YgPZHtLOMVIFAPh02p6411EWGYCYVQ2jI2XeYIsgZWv+kLVtqm5
eFWg2h9WE601FYSbvYD2BKu/dA74dq8XQagUAoaqowZ4qB0H7h5MgPk1tFJ+FVCg
ekeSUkbuMyv9EvdKdICRvW4lwqatcq5IJaorZOlq5LY/ysvcIC/YoTFAQitCdzDN
0mSeJW76l3AtzM04K+S5RyPhdx7zdEwKGChwqIcCuwCCGYIe0DGT5tmDav8Ak9EN
iHtSTlD7+hkR24yMgjYRxV/KuTWgZmYQQLv4sgYoilFuUrlLv+LRpZy9p7ijRfwm
IadRltsJymOwiY0r00YRX/oueSCXqQnfC3BZwzyWvl427lhpy0DgYgVaycos+6Nd
pLld2+dAyJPI2d/6oWbXQfSXNwoG0dJSWPc//PZII3UHhNwnL8MCjimRtA74mjS9
+w2JBORAUHyuKlpcz8r++pAlAlvDGwFFyTaCov/kpLA0ancHZSAlrFxhD3ZrgYZt
Ju+VX2WjxAyhQ2hXfbdV3RfeKMmGZ/ccMdUBMvfxKun6VtXsnJp5VdBgim1jexVV
Y/VgE2UWBLS0fnNRvESCkKEHwdPUzWseJRs6ShyVSAWDDllMeAkhG9pN00wgr0rZ
txCMTXTojzZHn8mhslF1edNzI/Q8eHIEYSLD5AKvmNVNY9TImlepsNT4cBJDaJy1
9DwhroVWSKZ5OLZB820kVFjAgaPqxoR79X3CXADICM0z+YPkSFRD74/uZgcmjOmi
gFdobqidEoWdLWwqvbQ6aVcnjyZvt1AaFUEVekcGAMPGDEyoossMzG4SwJQE3AmC
NYeNqBw4jByY7qfZcrXrDppJsCJiXpND76yrjPgUdeoxrRPA/cSOIyPjgScZoQt1
eSmfzn58B94c5vg25IeR9n7x4/O0CJCYRKmbayK56DxUrzpG1T5W361eaU85RNzV
Zn5y8WqzHqzE41kZ9VQn4NfFn8F3V3xPCOBxikJm19M6lTvnyoeYC77jFPVHpC6O
nZYoiK5dUakh21F35gnkfhtZV4FoiZNstDIfueiLPpT6jUlzdV03wxzs1K6AmQOS
ztuyWkB5F7HbobCXPoz1We8gBIzEMFCaKgsOyn9zlHQJiBN4GRSiod/Yl71RR9hg
jRVaFvNAsC+KfoXbpv2AlRAYyBfQaQDCpLQdwV5hmvB9xsTucFCQOO+M3gWRox1h
pY2BAFodNzhrUa9jYk0XObSQVxfpw38kCPNA9Cx5XpA8udNwQRlOfRTMjR2Awrd9
LuweSPi0FihKhXKpY+PGHvjNEyD/P7SMxD+DSgREc/7ninNXC2tcK9cUzt+vjhhu
aTLJpgHc9JmnNb0Y7MtQza9QN/rUls4JfUbXMBlc4UBUkRF68d9n3wc9EhDcKtzt
Z4ZFjOHq/05n8X1COwLrYH/nQg+MkUQCiHSpbFwkoFjoLTZAjzNwXEX2In+8g6Bs
/W1fb8dBoJp1aqtRh2KgpABOn5lo+utVaHVrJe4GxEfB/cMhO90g/meeLQgqsQqZ
wwoek9TN8JQDpGkMab9pfU9ug/EbA1XnSTnFdX4zr4NV3NCOyzRq3Z7LM+hsWSJf
6kBRoeVdchjhvc85EwKN3ki97n3QrzkFWHXhDMSiHjhfnxeG8OVsgQd7Y4WioCox
hTPY3lr8nD1dAItA3bZ+JpFPAgbi0toxFsI8JMfB0UPxOZ4cI27u5wLe3ts/kxXG
6CXdEuhgAO8FB6OPieyNLUCWth2mZ5RvH5eiwMj8iKqiUcKxhbB1TpfY6kC6CwfH
w0ZgX2V2v3HFp8fv7yMLXlDEX0G56P6EZ2PDHOyGJh8v9Pqn+VsDeGFXk9vFD0ji
f2HiT8kOtI25hfDxSCAMJ1VhSC/eF+dI0BmXMl4dfbxNuqwF/5FEZaI5KJNbljMU
TSkBnnU2jGmu0vmkYAkypUEkB8Ac9ZYeOGw52Nc+YecpyInOxWkLgpTtRMhs048C
W5qff2F4xJGPTh0zgqq/Un69pm4WWhk9GU92pFJeoTEC3R8fO46KJQGd74xP28wa
cg8dPzeANzuJztbOLLRZTASaPDkZ6ZAt/PCkiQpYrjoH8+mPHvbjRdjabVnLSnfU
+KjdlCNlcMsWfruLVV8X/8Sfi0wIOb75099HtOVijhm1TYFKK3rnwj9zyr6VuIif
rix5+xKpMe+p+x7XfRDjxTsvuGFHU854F4a43mtrbidce8rp56T1/x5n44K981rg
M4m2oxxC5isguMKqfgxFVmoFussHTIr1NKO3kJWQsg3tAM7teTiT3e1KyBYpkztc
Oi48oi3gGoK+ExN+11ne/ACkkFmRG3RvRRDMwZ0R0N9BiHyq05k/LZ2QgoPEg2Ct
UMrHzCFbjaw0lb0ehPPD0aJdezRObyxvoLVCoymYiOfwAff7zGQsHkYRt5OeuMhe
VEDvoU1+b4dpA0LWRJQ17zu1qM2V/eOnP+ZcBPw/Mz1llKpMDhkC4993POGYgegH
pPCMWrOPKwL3FBFu6HL0S2QA1feEhs4gT17eJHcqN3ZRiYooTWJvjHbueh3vb1fG
qQS6JURXWufc2DgYaQCVkbytA98HPL0JCgjD2zyLEbMIiboAelYy179zGthDn3pi
mm/eisAEelyda5SIbJ8sXqma2nVYmlMPkOjU7uQfozm1j8IXa4ibbGk25fKxWlgt
v9WLzdEtDbJSzNzmago/1tMfPcdqT//HQtsH7Qe3TBRlyhOaap288Fz5Iw3LSY03
GqNgjq/3Ni7ol1R/4xfprPMo305O1mlfa05XnAT9Ib9nlMCyUczU1ERTU+A/zHrv
QqD/sJYl/Kz07zYsdem/0ZJmeYihhzc/t9izUo3GXiayHtsPwV2tTKnzOvIh6ex3
dlq3ABZIBzryHKkuoEa/HrTbnJvy5J+4gt1r5XBd4BYBvEFPfUGAj6T6KODY96zk
dLZzdtkcfaxENNuXAqN7yuAYMfo+nAX+PlHyTt+i7LO3hwxT9+7ZH4KFJsGclNnM
nqS3YRbJsIR9aU83Ilb8YDo6bChXfeYzbRZVTrsHxgU0Z7aG3DV3+VEcVZEtsp8X
KiKxqpBFqWtW/VLvR4aExJ5FzVCTPFBE1sXuTJ5Cg5c0ACYbJP6PWTcSUb4/BCp3
FIPlDbXA5q2nVh5JLc7QLqN10RZYd+aRrkUZUnD4MvRd673qPrAoLiFx3aQoFCAg
IDMKoPnrrFDC/Id0m+862kUdpCK9Pei+gRRzS3AqhndpGsX79yupU0pKx6q7O0hI
uEHn8KY3ErRTu2BWZIQKdQModt+uzkSN8nvLsYD9lw1UWPaD5QDL0m868iFljFiM
IOHLGx0paXxEnsxfMSgyPj/rWGod6dmGiDzjT/tOi383TqAlBF1NDHdj4OjObhBC
Nbl9XHmwPbWDadEH3i6iJ3f427hvDYYegqemMltMNJC2LgtN50m4hWqQEms9kxqy
NqBcraEswq62avJ+CR1ZcnYeXD9M/3FgPfHPy/6WpH//I+jqExyVebJSbrngp38I
e8VyxAZC9nG24bSWwsbvlare0yCECctScP9KDpyALaCm5Kt/qIwqiT7/2NJXrwAQ
wfN8Nc8hCQmmlZcDbKhi7Q7j6mrIAU+2Gbb/U4DpfbaP+INjZVMdQN9oWX3P6nc/
B3oRxsRdCrZK23hJjlWoS2XZVD6fBTAGdE0PyNqGDvGgapjnm/+zyFA8OSluh09t
6IpWrBR2HGEmcAIvxI5i1yQ0n8G91Xn18rzecdPuoe4leaFOWKBZYvOniU05QhpX
23wGCkQ7aSIXlWtGisLZgDN5OxK0YEdDXGeh9bfpyXbf4FeS0Mzb4TDpE7ARKMFP
cjdyak1fMSublnZicw2RIEoJ267zOvXkUsy3QkJeGmIchSJZ0OfRCVlp/7t33RjF
fF4GesAL2NnAevxdG03MPFuS7PJ83g83ParKrxofCZaW7bcJMhUdA4T6WUrhPMCQ
719LmAF8DsRlcnILDnAP/VcnfZ84eXCYXNlKuV5LoHtUz2SaheZDWRr+uq0EE847
FBd/FSrUrX1nPWJEzhpCbb1Y8lBITlRcgoW4zns9U3UoX8U/Op55aJqD0IAS3bES
Xd7W9kszNLnoyo41j4TUzoKXQ3q883Xa+GItDRH9Z6nGZ5n4E4bqD7DyEASPAzut
cD38eu5neG2amyOCoaJr8ugjCtsJMfTV9EoNb5EA3jq6fc6d5JQCPCu7d7wa+Wvm
5DQhJuvuiyqKjpWUmQywHmI2NYasC8STmOH9qzekGRZMGRU1DuoujmD9AyNXyZsh
IVT3Bkk01BS63bRvP9Xp+ElbXEjmlCcaZPGXhNejrwAhl7UePQLkci7Z/Ay9THPy
5P+jIBmJfCHkiu3oKzUUUboO63ismC88zau+3GBht51ypvm7eKUr7cGoJ/VLtpmE
T0LHifw1xKfqdwEaJ3TUup9jqK05oIe+CDeVv4qIlsXmA8hWyR7kIwR1dUKmiHGl
ejX3+Kfa+rrRGpKhGbaljoayAcS4fuTUbC+NGG8+kwE6p9lV2MiGaD/9pbleoG7B
1Smj+1t0d53ZAC7oggD7TsMVqpa0+6HSOTnlwyROtMvpvaeC70s7gJyCE4t4dI4w
8z2SdDQMtEwOzs7n+aDKLdVjlWMwtzJiSUAqyNV+sa0kA0+9TvD2AbDNHfnejhta
pXcgEgz355jy7rnKAD6atuv3TlXb3IreYJVEqAUh5SmMYidAQb92PB9F64K0DVkh
a4vayPigYzCf4eAqY6DWkAa1YYUoOa5aj9SlKBmqCaU2Z7XyAhuELt5guVMn3Ghc
S246lfRa5yNaL8HtPzu7H+0BE39qAirkfrbBkwrRomhlztIJ90W/08IMVE2Ni+0P
JP1jOhm6LI6RhcbiBVyyqJZYgRfVABSqsZ5fJr11rj1jdyvqjg+VHW537wRDWbOK
TWg97sZagNZIXhUhmwIKxiASkQTjvi0m9tTWS9Mk9o4XTp/u23YjpBoJmP1h9n8u
FiuupcPZiGbFCvvaAque0xbctIAfM/MTaEusHANfOB/IwiSyZMIWBFnwtd8DPkkr
q3YRFcCTtxxBmfatsT7MBcz5WGSpGasYB9qz5gaY+vQiBLB2Aq1anc4hp7sZh2p7
KlKVPwPijPQf5qDuj6XRn8t9N+R9jBpQ2xY1vmQJEhbDrLjkEwuX4BpkoHEYtjUe
uWh06xTZS7AXCnfISuMDk5rghghxF6O6vQwn2WpLp+kIf/u38fUGQQRH8mk7ZRXr
mor+HWx7MjFNFH6HFqDVswwHAZ8asmMRDB0VSXdVFVYg5mkgwe9aIejXOjdwT3RK
oHd2Jd++ItJ2dh9zLuDnmVGnOXJfU5CgrePcvsX9IzBuYxTCXDMW3xITtWNlMrFU
aX5/oXpSnQvfYfSQufGMuyajB9pNvyHooPlFlAm1S5GxvQHbCy6f9HWKiqh3+KHw
PC6cp/WYnrkJyAV9ub2akQkZxYT2S+MTLp3LMPKlndEcTyyO0WQTqKlKfnBYZZZX
dGp17m6nehOCfGQrl8r8e7HS5vpZuQ6aBv+OS6y7Z044ZwSTpEE17UHMyIJqq0T1
KA0MVs6fXahXt62m0PfxTCcPLECXNfu1TgpwQYEv8/batWIt8o2WGW7jfLpQreSU
9YPtLqLBO3bBnx3FwFxupLruvItFGpTNmb3tOGC/pJacASo4Lr75Rz/n2EGz9X6J
iZcjqP/t0O4xvqziHKWD2Uoz2VlGig64MiKna6SMu6ptvIMpMSQAam3jcDph7kAY
sn9eybfqJMKDSYLSh4TQCqkkuGVRIjZB9+k7VuHsQhCQBu8S+vAU5t5XRh0jdP3n
286ifMV8BxMPODImmngRWvA+SXfSOopEYQrz1hwZUsKK3vpD2KVM5/gkLsnyG1DG
XgArmVjxu/Mqt3ncMcK52/0ZxR4p4eEL/UGWNqblYh1ZjYmp6uy/MDNjfsE6O5xh
opi+GBvuvA3rA9+67jFbHDfG/+JOtAG9hMdTalpmJdBUUAIsEp4vpCRnlQNFKMyo
wJY2YXOWFSX3yrXhwT3VL7tIZ5C6M/QVzkUyWTIXTHVqSNU4A0AWqWdGRI9mRBO8
wwA6FUpVT5z5quzXqSllTvMDvfHY12mNPbblLcXbjG/czwGmGJRxBXKrgdXCUeMv
T3dhGJBWW251Z/LRlpSDG4uzqnMvDlXckszXrTrTqLn7ctHb3cqnuKsVo6EjTe8I
NDJzAEVObazLMzfboS+y7LA6fuYDPqaz0Golxul/Q9XKJtjAgfNjh4Mu/ePOpieP
b1gZ86EDUyAJxT3Gqdjke3t9nVccQZAoxS4QQWf6wJiy4GlRS9KWCYkQ5U9WZCgM
IRY2qeZF0TWabvCuC3Und6I0y5+T4OG3W7wZqU/28+olS4pV+z15SBi49nWcSkLx
bqjwTeeOCe1uhlpWIAMU06zLP9rHXONxb01uYGkJVat6sg3xCUJCcm6MmLsDrlzm
1PKqfpBhMAX1iCFAbsvYrB5UWitqYuDVP2Onl5xxzJGK8sX/ARl5m6qA5d0V1StT
bUa04mEZFvR2cfuJNECr+n0w2Di7vLCEOdCe2O0lTm41G8n/2JJDRCWhmx/1cElZ
1C/cqo8rixRRbXC8KU/mGc0R0vzv87rc/N//GrY2j9hWCW3OkbH9iu7T8IVttoi9
Gg3LScK2O3aF1ikii3QOZz2iQjTi9sGcAY5DlJDJtTwsrOa2hafAk/5dMSwL7UVg
L565Wa19GfxAEpHrC487olovmxZAL7jWQQMAX8Flh21XTFYJoq62qf/zkgYEX+3Z
ghoZT2hPfJIDR5MGuA+5Q0LZBP2n5TBq+1Yt5EQKa+QL1hjjoWfeg5niY6RguZLn
hOrap8R5NmJoyuW7kPOWCXm//ewnyKMVSUiWb4ARY5VCi6xw9qUHBQ66X187XmN1
LYUGDm68mPaH5PC1Nv4FfLCQ+lZso9/85LjPZa4IXzRkhgJtOnsLKYrFJbv61JN7
PNzQHX1Iwy5xGZBaU9gzTuYo1d1NijLZr97nJ6oD2bm0TfQm/wdQSC4TmgnltEWS
ZY+a5/jh9tHHZl+S4Xt57U7bkaxhIJbuV7PHbGRM+lKQf83vwmNrv51KP/+HQlg+
FEEouRfxavinOrFSI2rdNXlHRmDBxDcf+mFIMviw7IZ6gj6DC6QpWVH1AtcG/Oy5
AMMZRVrCV0qbYoTDmngpfcnbzav9dEmv+n1JVsCTzPCg5WS4m0sjKcmDyC1SDp0L
zktb/c+JbiMH7a+N+3Ug8vps2Zn83/DBMQKZyQV+C6Y271lIX6fPSIXPooIuo5bX
YnkKKWVixEguGOxyzv0fxGBBpcFDtjqdMsYkVQWZ3TpFR4u1gi6bdBVhiJxCC/jb
C+laExq/dGpiHvzbLG5H8Jx1yPLV0Pm02IcjETJubEF2hj/n+fkCcGzdRugfHt+x
uyo6P24XYsnuk4aCq3+CX73kGeRZAowheQk/gfyyFv3Z/07xrABQL2yZCooQz0mG
Dyqlj6Zxw/SCTze8K/K6mHHQLkywKMgHV0VvOtoQXqD0rBjP+L9H9XFrzW22ClIG
ETawI5dXZ04f/OBV/TtGCIMgntdvBsxz3p+2g4JW7MoW0IGDd+WU8Gniu6DjNGq7
C0GqtBsWmGb++l/bMRJyBEtwJ/+R9xdFSRdz/GQt3BvF9hxB64GDVn2JbxbpXOja
ohWcZbdRnvry1T6SiIJIrdnjwsmSfsNGQFvH0qNTWDTYqbYdyJ6P2bCIMkwXTKec
phJg4qTWziQRW28USBywOQrpO/rwvqX4RW36EVmfevx/7VcQhBRQwq8VgwswdmVE
EJu4ZJx+vRX4XX2IcNvjz+SjwTxd8Da14j/AC5XBhbIJnXKmEvnot23V+4SP+4Tx
HhMOLDpGpX7dkyJp0pZxL2RN5PDTRUn/w8l7V5w1yVwhpqbk4BSqpo7HjaRvtu5r
7tPiVhS4Q+51n63M4KhHBTFNSsEeVvNSl3ETa3e3PKK8QMGqCDvKSDMl19FWxJ+S
uLLHDhLRhthmvnuKJB0zTi2oRCR4XqIxYCoGOaIMZ9Joey8J84OHADVwC2b0M8aw
Eg79dOXjOoj3nv4XdCZhTTllAuSfUjiE019wkivZAkFwCohHElsXk/QNamAx3zEg
jZsA6YmbI1enrthsThZqZX29j170MUX3JXcHlfc4C9XD10fGy2BOTG6m+p4jaRJb
+HdXA8AR60aLl7jAIliPLwbaSIpGWbMW3CFn0i2xAR3pQp1s1mruNzF4nKTtZpdt
nB2zW8/KNfvBtHRrq85tEPx3KDWpsiqbmfEP0kbS4SSF19vQoBY/4OZkPmcJanZM
f051B1tIFz+lYYZJupXjFc4HnbCjMM9Ew+5IUFLRrNQ7ZHx7P/sWSa67cw8OuNYw
D914EQpXu0ZX2qX5w/9/hNqaIT0cscgA/nA7Y3ou7O8a03VWZCAFkXl626+5fF5M
zXC//TOOASZIRJT/AVY9uBMQ6ZcQqs+PhzSLniEsGxJ2FAi83L9t2sLukXmptFLh
ayb0jcSjsYSM3eP3YcTlxGb/opO8DwcWaU7X0QTL+0XzGPXn0gWMRbZi4sm43RPE
39GB3ChZ7mDgPtVPokhbDZweAG9zQJt10myA84yHHNyi4Kw85BImCZ8qWFNxqJsw
54ZotMJH3WUMRw+gmKrX6aAeIDQCBxIwMMq3sgY0ApCd/aErGclb4IVM4KoiLprW
dEnDLsmx0s1Bk6ByBER3295t9o8f4PsmkmkfNwHZ3M39bEIqH565EYuRMHMFjyEF
uHT4Nqwt/Cxt40fRoCwC0JgQoADQfvDHp00Blh/8ReRnFNiK0qbAZ1bVynahlyOo
AuGMS/NAmcTaQeja65HWoVD/CGRJU0+uDka/EwkAgIrYYGAMRCVfuI1aaVkudczJ
qBuzIL7q0bMYyZWgfZy+OR/NrqdTZbH+K6eIFbID1XY9XmwFT31XWweXt0xhyxmv
l3VSm3pj40iln/3gXzl+BwevOu0IsusARQ47ZVbEah96RbRzisz5+t7/HU9YOoKy
endJvCIHJhOsEDZXmew32P9Vlr48LKdiR3IWdNg8Tg4UPxba2yvchIu5mbJnhhff
XjCSTXBg8KBpgPGt3NgPLZ/iRscXTBt3IJQdc8cZRhBhoXeqObG8PinqxA0XvaNd
Dz7lESjlxIFnCdMn8NrBae6IGaI4rn0ExtxG5V9C7VBqbP1feOpDuwrXvjn4+vJD
b47UPMWODSHKBw8W+8cG3VNmxJB0+XqQysc83lk/lBdFcU2cwijXAd3k/NTLplv+
eBMNgcjOn7NNg08jlEAbMaglqe8u00ErkzkDRr9f5cW7PzOFWM1EfOWOh7cb7Mm7
EEOIeRRPFOt1HBdx0rpt960uiftCo//TPdEZFK9NeI9xyLswDsxPOB8gs4mvAwln
vcwnm5DILMHg1QXuas+UCSFXVj7ODHR8JSWj1GnymMJGbAekoFHovg8vgh8Nkw1o
zkx+Tj9tmSqfFjZzmdW/BHYBFUH+l9CPuZUNIX6Oc+9A0WcXOJ5q8w7+5Cg63F+x
IdwKZt9eWCZwyo3b1qD+eG/BAdpopZ0SL8SvC08Fw2FGPS7Enf/pR457Oc5M3yNv
m2KFZFpwC6Z+/lhMPYQTA59E4+4x+pUnUDYun3lXOQQ24uB/KY4ul111HucHM2Ty
uUYsUr3l0wOfALZS8E6oVwnE5LHT48uPi9ncaK3KLFMX3ko6phicwNpyo8hSOVwx
C1y/645maAfahSvo0ReUAbQ5vobvcJx5WcM3yvEelUVLft7VYNZqvx2zOkKtmZ0u
GlHHak8oc2aWJmPLttT/Na0V0G5dHeaiyKhgjILd3doBihJ45lYMRrnLrj0P8jTw
ygR6LDNV5+mHQm4ud0X3R8iariAvTHFYfzZODiX+6z8oa4l8QTmHVCdXLRXE5UNk
iEe5nGPsrLUPNT8pMdBIcOOXazUuLO7eQX7pe6BzJkEj7lfD86fl8IqpXMuS+h6r
DYzclE2UzSSYxOKHkx/p9F7v1Lel8qlSjO/FMToYNKQEFuhNPIWdxxnj1RlodulZ
KJk+mPCoLFbMhURDlU7wm9VTuzrapsYOwZUqzvc8ExHYXj90itThlEUYyJN7u9Ym
1zsK6rJ5yhz7rhD/hT9F+Z2vaSVmH20/vIsz8W62N8CdhJY8jhB86DZWlZiv1XyN
Y8A0bMycY9zKGzP9rqZTIwMh8GuKREE3P9yuO7WP/c1lK2iGhpWH/rksN8ERD6cz
K4amrVx+HG41IFum4wzXO1oFoMInF21Su5oGVK8VhpKB8EWNebHYcTOq4oxgz4Pt
hgBXIPJx6regBZkMfyxEfGrS6J1rSfc4l24PYmp08BYwiFU85a2jfv5dIxOEcSye
qs1cvv95dH4oNVgdkblpqIKnL8Fkn88PUF1d17y/OTkCPqB+rp1DWKjOZTsOVA97
2cuXNi2DPFt8kuKZFb9JbxqcBCzGN9FKBvpCo2En5FlgCSpwvtsNcUOevwlp4MvS
sP40afWHmUfouVhM2aq7OjLWoG2AM7swU+8gAJTl6gi57297/VKnwPwoMXY8G0tF
sMVehQq+u4QQcg+StkPz3Yyy3CIH+Xzj5QQpnkIAriy+UPq8Ws4nDI4jgU27kBVz
n3SEvRrXRzfruMf50Nb5aeLaklz8zkjpUUJDYp/5GbBptH5yBqZxWN3LSIr9Mwx/
/TecdloSHnjC7AYX/8GSQQtZesplAnUeQP8uFM5TplTIVxHxdKUvaK9HQ1floEYi
JSlQ+yCRykk3q5ZbPaSIPGD0bsU+5Y04F3IeiKlUlFpmKd9SkURcedrCMlsUrH5P
Dmjo19K4c20vvGa8tUpa8iqfnRfW5pab41Norf90QncXDlGzrugnQf928ylOrdgH
A9XK5vPPvlPx5tA4jR+8cPbMCKrllg2Ek9govxEpCN6zuf9VXIBhnI0zYPMVNRTy
eaFv2L6+yb4aMnoD2H37e97uJauL0FeyP5y7MBQUf8APhbzaDmQokTMjZsWKWioQ
ZD3l4BcEQTgf9Co/8FVCjbz336IAz509ldw2KVMbxHOQuzPiN21IPX/tJmrMdPg7
kNLrIkcJMpg9l5AFF+gHm9yR9H71UHfR+LFr+qBmXkNzi7QjYAYNPp3XCq3O9eXk
bLrW/WSZzVdxvZRJvnxcY7iZ5v8GKN+/md4FOaLEfDI67BcteYQDKonyIWepxHfJ
cxhjhrsr0KLoq6Wx2bY+Noxj67AnR42tApd4neu7VMI0daHLVv5d8NuXyPUB8jpy
4EZuNl4QIYgC58PI38wXoku0EyY5DnLB0O3DvvrcMCe0Doa3ciE9z5P6Od3pH2xK
vM6PihxOnZyErIzNwoCSF8ji6IDFeDyvvGUpZ1g8g0RdDmOZ+3wS/Sv7MqHsA9lI
n4C1XS7CmXfZEReRxOpZM3AB/Pv9TvqnZnoNvE0uUBmYP3BNsDgzf5KlZ1WZ6DZS
dYA3TIVkozoDfpgoohnfqzUpELrofno6hdgpMg5AGU/sTOEEkzJas5/BcC3KNcrv
a5IqIJfPm50mcU+PZgId3QC7k/25SQxBf2ymoXdnOno99cA9gn65hnyNzCuF3A+U
u/aMMwgdkVYWgPRSDYXtUeqjyj8doKcFv7wAMhR88R57490PaSK6yK+Ki4hvf3AU
E2NJ/uTg4Xncf8FevuJLt3C/7diraj2kj/4iZgAAXhuZtJvEKMnvA3q29yeChqgG
IVRai9RGjTKDlbYcN6p62+DolzdYB9UXiv7cAX5yjvaUIvDAMDRLGmtI3zGUtknt
O2Ld+SCy0mpgHzRc/oWyopSROSbutRuCILz5BGDhAHnTFLM5a2KnBcmMfsXph/qq
/czy0D2lwMSPfVXDqY+f013vQj9IUSCPmARhvoKZhkQkJcMh3SXmlMewhDH4oIMz
wEMI1j/2J+CpvDb49XEwIRtyqQkv6hZKhdEdI4QivnN5dCqMlbfP2Vm2qBvloAXr
pzWMN6KvRIJYmFLNwQOhId/p6Pg8nykmYdm5GAABbEVMIMSRjYicHEyQ7Wip1xW+
dqchM9DJqaYNxdZuIAchJ1HwtIP+A9qwJHv/xA3kskd4Ej5Tvnout9MEW+ghb1Qo
0qm+01fmeR/vt9m0cdJjZkzK8B76Udiza0x36wX4R7tlM1NF96hRsxA7oHIiqKC9
ZYClrlJU7cBoPm7YxMoevzFc1EMIlQLezpXEc6yDjS5hGzXcSoqgF5s7/dIcKD+H
T0QUrTRQe8zLO1C/uj24DvLYtU5ix7Ydk8QO37UodslH83k9i+I4jkXv68Zs0VFI
FUHGzmmLcnbGSCvrxacKyFeD9k+kPn1GUYx4U7o0y3ToOlKNAcAvNIDpRQvwR6BC
+X6bnaoGo8KtFHGjlBr6w2+aH13P9mcuT1WJFMGrbKO5dc+R5huEKKQjANdrpO+i
kjw/003Rwx4gv+LxoJHQrzrXizURZ+cI2k0hVZQVGXb15fMy/uMZJz8t8C2AKyIq
cs6aUiYH42VXnNaWFHg/lUn6UYMSwyYZ/SKtrwEpbCkePyLgqNwVRjUC0CvSVKXT
fy623osde6sjbWCgxBIP/T2MDvD3j49nCiwl6GP63cbZhlxnJ9fdhpAW8NsSXbHd
mUSMbP5YKaVM58ycB3LFO9ynThBeP1vO2yQC99jEdAzOZF7nt3t5N8FJmf6kAC7d
0E/LI30lmFkiekk2V8/t5Fn8uBHjOJnbHuMeR0v9+pD2qWZlp9NIlDmE/9pAMaXz
Q9GzKdXMcK1VxhMwTgO51dJ0S5J1vL0EC2hhyyUioFbYYxUxcBF6ky2faqAwEanS
1+8SwrBNrk3Zsa6jkUbz23gRRA3MEkOkErKlEIlZy+xJamOEkAOwci9/JPJX9PXm
LWbhGmy0Feo/E1yJkX4XHRITSlxHOC1BPj/BPNZVg720GNBkG0vhYD+8LonubhTT
663B86cytloK062ppBBb+TYryGaHCWsaTVucpN3aOEcHjNpV5sFJ5NNBidwp7XYK
Vex81apjp5/RcSfL0Ynw/xLcm/brXZ2VvJIhX9+FhIIIXPWudaXMe+nuxjUz2BWa
zNZD60rEfvmpBz8dvUWgnbcLt77kNX/rxzR1wBu17PZZ/50C1MoHIFaV3bAzYAW1
GuZhUAsmodKCWQu+OPocEjOOoNgobW6wpMF7gZ1I+rhqNeTZyqW/vv7UH8z+d4DE
RacZAqpYqcBK0n7z/nGUcbD+vMkQPlLMQAo7sn8zo4iSp9YJuXrnHJWsWGujFAcc
aXfuDwghl1zDo54nebDySNJG9jN9xspYf7FWJ7KOYcgwWa7WGHQEjqgiTB+yiw12
avjby68ZuFliPc8lbJUyquDJo5JQZCSGHiA30OlWo+c1oHbxKPJjdnTWe8b0SXXS
PHe3xzM7eEbGgTemPIgSdHidG5poYcda3nw8dK1ZZX/+79vf7+kWmzMLbszMBkGG
hLwKkxRSBv8SvKrlbl+weebr0ct/PWH6eIbFYa63ZqJGsb9h7mG+HFGd2a9hrkXT
Z8E9toLB2qQTC8xdGB3ZgyyzCdAyj3/K1BoR5RnTXM5OI+D8Gux78sI+yLItUywm
Q23dZhFHZAvkkk+aBNqWw1FMrqRIlxSHdUpvOLS+34yUEZbceQQIdlk366qU3/fr
9WglruleLyNCqcA/w798TsHWGTgdha/dJkhBuRiafTscd4K54AnBg8YngJ3LFdWK
JHTKP6Y6QTG1ysoKA7odXabav2QXhV0vfdQ5lZkmehr+s2QXquqHRRKU+biuDDmp
l7ySLeHU0Gn43+Wb1M0QYTmoQ3YNJDedmmkGFHj43wlCsVHMGi5vPbs7YspfK+hF
psUHnDKSKMEHWh+XntP2w9zGESTVtuWZNVgowDZ8Ul1PUBG2b713mLUZg9JWXUU8
Zf078yyNVmgRCjio6oe3eBWTbwDZNe7ZZqCRrCEkUOiGuSSEIOg8RR0Xmk4+ZCkl
QaHEs2F1ijubDWygQo4EOE0l28Zemo227fm/iOB0Rv0g9C0kfE0gDogsrdQQC1Zf
ID705mSTmxipJ1L7MKGGnaLU858MVECPQQ3lsJ34dQgURAYUTrrRZt54AjSYXgRv
lT4Rm/ThzocDM7LT3eBH9ddsQQqy8BrsBBFirh9kquyQ/nLhzVnlbXN2PtO7KOZ/
neAz8+AvyI9fbSM6czXGpeN0O7hi//cpDOyD8bLi5SCyB8ACKOTY1a9yGJxtvM3/
iyO4NFhBz2xouEKWZqQ7L9gR8ZV5HW7jawJ+iULYkjVwXm3odLKtSYWLMh7bMYU7
LTEYt4898lmNUOp8l3UjTaY54zCGXuZJFgaXW1Fl4Yleyg8hvaYyTKEf5aiWCbx8
OPO68sQUXWRcZCsbvjTPnj1Z5GZCqFRMcJRhcBouN0Y3HfrTKZLsTIBs0K9GkJLj
Cyox3uSZH7NaF7CTVNHyOKSI15jn9L0H19OBR59IGSkfv1WLImE2VLuckGIaC9rX
2SQyJG+Y1OdFpFWf+3IhNmUKiuCj6UphdmEUlf/Gwht+hn6iEPZuQBcIrRvIdS1F
Rk9zqmV0MhOkAmLUg/H26vx7nplG1nZ66ITIOWJCH8xrgGwl/qH74fFWoDErQ5JP
gik4IvCH8XuB5IuhS6DC0uZiIG9rvvnQKxVpFsZpT0Q1JjCK1dJlxIh6vy8Q0ris
4hubAEo+UxkVt8xnkB+6hWmxsO/GZuZ9Dbm9yno5sMQ2XMhp20o2nvo4xbsaI+s0
iDmXE+Mb6WJUc0bMGiuBiE6x5R9GUdta6i4w4SLU7BjeJpI6RMy8tEkFxP9Jq9nZ
cK9zxrbf4wlRhfmTWLva/QjVzAXiR3wUaTQ0BVlm5/5kMEHXZtJCGk0p2Gv0uUeh
zqDvID0uWQ1G4Md9AK/yZybbHVNHL/O7iKhI24vRfE4C5IXeK6vuoOZEKgk8+fNK
eE7liOzG/2qBokkQC5quYEnaGMlZVyOERIVki3Nm9slxT73ahm2cugN/pysZn/6r
yR7Jg2ecN1nXpv9yi1XNa+lHeWzCXIn42RvOaQPOqdVHVNGJlSbWM1UyJ3pAccVu
bPa2G4KXORRkF90QOFRoP0o1AR9192FVHFrIKve+jm0pypbojOFxQw7LUoyaexeV
9gGuqqUs8gvJOJow32euKjmKvXReATxNkZPdaVC9cY+oIGDDZC2pz4Bs3505w4NY
h/OE83heuiZYHc3/vWQOwtK/RC/Nl5zzNVFBBUk5CMTUhwGh1niCYht4fVho1Hl5
FXYbDJCHRfxQvf+r/eLZzxKWAp29dmFFBAC1+7/d8Yu3rwB5M+mC85HQXkwR7kyX
YhN2ynspjzolrs6oF2PzSZvkKWL6ZFL40BGl/G4z02a5HapBXf00tLX1iyHT9q0B
5cVPDRkkNapUiTpVgVMKBdPgiKL7RkJnUXnO9thNgXSeJH/6pCLtHBaWOaG/rMjy
CiHDTYmdqdv0y9GU3r4BcFmt0yxZFBDPpRi1TXhSdd+8zD93ysQ1+Br0Phw9WghI
Vum0Eou6Im7cD48k3olwdS0btwN5585itZK1O9YAXKlo0EF7+kcPaaYJ1ffIY2+I
oglCGj2DPWRrAC270t/K1ZZrn68al73ffC9LYM5Y9I3gUmGlgtLT8GD7pQu970n3
xV3nK9+XwRfYTfeIlzjUjWX7Sn528NcQPLk4S63Q5uq0DZaCcO/E2ravfWD19FIy
ZOZTQicpa2EKgiXj6ZLbI/6vMWJMwM/3MW1OvvZKckWUH9yOWQjuI+6hWeZWEhG1
UUABqVmxayuRPdv5JPEK7ffUJqlpaTGhcFYNe9EekSYTaNc7+rBrPCLHJ1fbWtmL
0u2/9zWcrwj9fy/dJMFbpUblYeBxBmCWFMV+SyeFt5+MFEVAsNIoesm41YRHiKSA
6yOIWICn+wQSWxE6divD6MeGl1QTiwJ7A8qyyvr3s47qkOH/NruE9S6V4h2+il+e
P2owb6rzvvTPlRz9Nk5gIgah1So2HGKO2KtWm6jT43/ogPKEEwkfxH/UZ7cIYxBD
hssZgLRfXa3rX+D6+NiHFo0tbhQCuzMU2hPkqrHZY9dacnpjx4PsvHn+74vqXQeB
EjLbLMDOmIXdr7LjJIJIQEe/q1FK2OUQCyNrz/lS9o92QPX3mBiRzyX9UU9TMc2c
SP7p5MtaJXWtysiNJNTa1nq7/7Ta89Zv8dyyE8pD+UAabOdqHvWMAKxCddHXGbUm
JSohgGF4zGjygIJ8J1GzyV+wuedzdzmu4HqqJ7ucQVGOt0jDwEfX0R4XcLp4xVm3
UCQSYBvvcDdVJO9MZn9wBuK5sj4ALSC63LEMRxJF9d3yedSR+YuJ6EoWclIbVULy
7hF+Bm8ZmuSOHmx47TUeZhoXeZvYx9hy7RB1mM2wvAV0t2lkdBpR9aKtZfkEhzov
rX0w2RpEOl0IWG9tdP933MabdJGUqVN6VntgL+NwXLdjxvYH6e+PVPuflNbtLT4n
85MlPB1jM206mfNEbD1aBGGn1AB800TZqf6kNmw4likjTvJ5xhjbdLiP8geFHNbd
3nKzIuMVswfy/OWNb1FRop7Ji2aE4NGByd4Il6Dsx7nx8FCnUqh8QfhI6048IflD
WtFBOvR1PX5dY9IZCtlcFNqVZGAxweZ6keqfcLXJWeXPdZQgyxeStHGNlGv4e5iR
qC/6lwMUHudCHX20V5py53yECKWwivhdaKF8L6KKW3Ny0K1b1U1BToWPW5gZC65o
mKiswV4VMAXxFKy6jgVUQhJxD9E0i1TuwVDdsZ8y2WykZlP4UnjdZaTXUXVCo35y
cLJYw/E8REheJ5yJdMck+vrltRjAVZEFIiUacU6lnlMKxSPGGOvdpcR1G+HnHuW9
eqkuQBgck4Uyo4/2M1IJHWEGB0wqLmuQ3YiNws5SxaE3wKG4dOgVMHcQoadmyeFV
KXPtEuBbwf89u7ldyDYW72mrE4EdpBOc8MbswrYDkScI2d74Ep1Ej6V/Ez5JFIPt
T1sRuH4IiAROXc2k0lsiY4BxqVF5//VTsRc0JLez9DhI1AhtG8ODTskACjOBg535
Qicn0SADj9pgUMwnlYRYj0/haUPOoVTqDX0mIhuR2ObNMTcqY+bYfhW64o/MI+8z
sxgivte5ZFvXBNOi5QyfUqbs3Ki8ZEGio36kSBZfVf1DPJB6umWkiRe6d/ki5xLg
TM5ZmxY6OOyMpeDsyLR1G4UU19HG1ER7KPNrJDrg4DxZU51V6iMK0TVPBeIKvZ2J
TZWlW9em6+W4PcGZjH4V0LkxRFsnybbTUG28+NDkImwh9INd5zCrRpjhNyjUPvPN
wx3RP8Box3GvbRNxA+HGBbXfgEtb1CLbp1ydvD/M1ZjoJXx96TLOA5m3ucB3eB0z
kNbSe0NG9RsESpx1B8W9M1T1gvpPBTDYn8mFgPUiCwiaEa1hmgiyts2577d6Wxwz
DgmteHFrUTTb/ZUFmBLeG4T4sxWKPEZU3CTSpkIWhZXjyMzpW/vrDPudVo4mupJ0
Xt0rrlIAmsFMbTDorlamoC9Pt8UGTnQeU5hoOQgRU7zGfDXcjKAXlQISmL9+DVuJ
g7XXtSRXn1EVunoUdA9IHq8Nah4VQnA+mUQyFSuPqfY/Ri4zYTIQN95AvUdm4lfi
3xZrr2M9l6eU6xzlnY3QLTWO6V4Mr8W1gC+AsKVxbJQyQdvvflwaeW8+aCqmln4t
CasepcheQoxQCLMB+MLkqkZ6FHtusX66L4oJf+clvQzUQh2yZ6BTi4wNgPCsnW2Z
uJLVXm6Ahyax5n3Gh0+Ix1GTQ5l+sG7TtVTRMZvb5JOIUBQX6OhVcDj1hU15LQ+h
OEHsJ0dE/C3fqlzMQdE9PVx21SS2JkB+eLn6YUfcrfWnPwVaSCF6z3Arggwt2DOB
epydj9r/OoLo113IVm32htOl5eoXs6wk839u7LWav40/MsaJHCuPjwIlVcDnzwrk
nnlK7DwOzlkOwrBI3z9zbMUN78NA1pKHf/R8ssEWJzxjJKbmWxaZ7ZgaM5uRLr1y
63pLccbC63jkd2Ea7RJGNRif4CtEL8qME7deHh+pvgPH+bDSvF/NO9C2Bqzw/AyU
7f7NUFdEFKusnDStP3LJXH1+dOaFPrrZIW8oPjh+x4Q+hjfj3baVpHVbeNFsHPce
8xxdW8yhWLDGgBfvBV/lrJyuZMKXmX2hdD/WdeAHTlMTxJrD2+Ju/pU8Y85gd6hL
kkCtgWlUcHMIKFiYKmy7JR0ZQBs3OcEgKChrcRLo+uTNlfRcq7eywYGsonMAxzzR
uwwxXD7nMgj8xr4x0Af3+KDx2ty/IopO6CrEOePICcIF1xZMiJjcpO2ntzY3OXVf
hv8mvyF5bk6VddN/pepUrZrSgjXMes/JISJyV520TIm3SQaSK4XEGqTVheSMpVEK
dv/uBch94OBDjZbYGBcaWdTWE2efZA909IqDh6vEU5kLpI60IQZBrZ8ywvrLcNjq
9LLB8iWfWtVTLLK4BD6IPpKHR/xUjEabtelVKlRsgu2nO1ilYC20tgsl07Sgv5Nl
FoTchkpkWE6eAf8U5ShfPJvHULA+R3yMAgQwd2SanBJcZ4L45uWvhhjKZIZ6v0tT
NIXlNy6GdGaT+7G+pb4yHDcfo5R1OCQ13UpIiaflZrcWS1PhivDyUDIUoyZsSlvN
wFyrE14ggRHeWkDBTDMlt6g2k7AUYm/Mz3+xeQN8AYHqhxOSYcEc/uxYsmCYkYD8
HjeWFwB5TrCqLKZYtYgA1tiJAE9Qcn1aDVcI9ndXoqZuYO+0Bu0farvXNxzAH1HM
OGqoXlZElenPCOoZrXXkiLGpNLeqNQDKGB7wHKsfTbtSMTPZZRvabKgLoqhjuB3m
TR+SCLk7jWGUlzU3dTBVldgxbXi0YFO8e3JM50xBrB80bB71qEyRyhaU0QtLTXLU
wjZn2ZYoSg2F6V6mi/GF2gWzLxNVxi1EuAgSRoCyRFrp+X/cL02MCvvV87603wFt
ztL0RTGAUM2gwbhTJhDXNBACHebDmJLAZfHcwJwMzFQEsh/NAwnxgJ4SYjiXFAtI
1gd9U0aOMIvBpoEqDi2+6idamLgdgE+JIbca6P1X39AqQBl8kfFNsQQlR1wqNV6p
zG9c+OJe7qqpur+lgqtx4nO0F7iZsCkWaR1tIurSwCUK+wCO+ab6tR2Wwh+aGvDC
QMF20HotvAf/g2y99tk/6kX6YoBOt7Fvkw3huomabl+OjIIXQY0D2xOIU9dhwljr
WpobXm3l81EaaRlLLsq0JDWKJnE+CdiACN5vovPWkjjxXLVum/sY16bzOxyHgeF7
eAMM74E5CuH+Fz5plg12s8VKgaRo5+DpB7uJDlMDhSnfcM/FkwfZUDBtg7G8Vg8O
Po8OUbHwgaZspxVW7sdWoGnpEw7CePEx5/4zNCAVaO3C5H2sVESEOH/nK+DgwboK
R6CT5fUdWBskabtp3RmYsLnQv6CCp8JjiWcVw3slsiu8q5IleLBBCNjUC408t5D2
uEiu1zuNL9z/no8k1FTiJmmaM1LHAFawxzWIFbqkWZc4RoJj2kQd+D2eOa9oytO9
RSn9BSPoPWjSvnsW0FI3xcCHxM4cCXq5YUh+0SNa3b240iCc2LXdLbC0DdMxXOhb
ZI+1gAr2HCmF55Sq4ajz8/KePQSLDGv/VrZC7tCHW5Ztcm43++Hq4jZIF93TjUyt
0llzrDJ/DwbNL1CY5SN3D015ZktXBnM2SriXQkg9NtcOK3sdm/axn1gHBvfcbj74
ZKxaOfzlEitadalfer99dA8iYMFe89lMq7JYhn82SzkRn6uLv5vgXh7mrRfiJ4wm
cgyt3uL69ACNKmhfz0rDEEEx+8XTT2Jnj+SIFE1jz+IiobMRODfC1SKZaSIrZcVN
XbpNN9cwbwxpIGcICz5xyXCKhHcWInC8DpjqxSqX07xAvbkParGEhJZ8pC4hKJHn
g5seyOjvQ/xIMwqBxoFK8snxs2DizCz4zJehTuZfdvrJcDjXLtBgNaXW+cLsGUKd
FyIF08oBJD3rqbenxO2RA7rWPOuy0h+fAfNktwzX4uy0oj8TqtqOSBCUWa7GqySE
TWxKZhtq1zqvYTP0U1C1T95ybkXVFi1TYEfcC+WJ0fEd9UQq50qaLi9CU8jNVSVe
k39yqOlkm13LO2NMvad0ysnRDAgBhMgmlnvADaL/LwHafHwIr9BCcGBg05w3j6ii
4vi6Przqik0uEltVssutAHiO2Pu7lgtCLq3cWptTqEM/Bi9wP7IHXc9mYzuFdc/s
LuIL5vO8M0EmZU249qdNL5JsBlf1lw9SzcZgSXWqEMb6j4X2CnAe2x/Kljc12AJw
t+oZLyw7yd8aHbTw2DaRQXgf6PN8cmDwINS7PMpetBIQ1gnTznkaQZZDTiVigZhN
QTXw2IZlOfw0GV2iKuV2hCRFEYCBbvvUCLMkYaz8VY5KDYST0nw3vdGuQgzrH7ox
msBG3wa1AZDW0Il2J08Gt5894c0eul6hLGDLToK96xTb8LSkR9mdu6BfQEW316/g
xq5B0s0uDRcOg6l4hX0yADGM8pJmUQI5F0pjDS8pfNJmKnIdQULtieras3WFdo3u
dPfA2l+O+dRIQR2eSNLPccGxGLKu+zfjRXonmknsF3GhGIh3oJlW+VqPz/uoFD4l
nT0Wh2ppDtDE6m14Kw5MMHOPMoSmzR4nsO1gEhaqOrqPu9vzKhDZqqU4lWrMWTOw
Vd/u+1xsKazZlBa422l/zg43Jizh+3ElrRhzh2Uydf/fIb6Q+m4Ktl4OAc8XLlI9
/9NL/ZqexHemHpFvp2coGDShtYl29JLihfCopNGyJUQIsI6CfQRXsJCjDfKaTqlN
tMRzBHImja9iAiKMfJAio4+GXvWy8pPM1bTIP6WbE+8o/CeBFGcGDPkoWLh+hPIk
SljLagaZ5CCTNu9l8gZ2j3YBDdSzVHmJa1uJLYdfYJuO2/zgNO9oyraMXyUkJ8xu
LNaHp80yBjqcbEprSiCeVGeaVNjfWZRxGi8eljbkB551NQzVuMt0k0oQSc18Uplb
bDkoBSWOKU3vvA42dQdLOFH5FXsGjYZZsFNsJ3ac2+QP1balrhm6q8NQTmjlLLXT
kHhcb1dCH2pWsnKmJ3saY9tbb8MpqCLaQrIZu33/0vIlthC4l1GmAc46jzVowWbm
e51jJuQ58d8do7qXwrJDJMlyLHW6fdISo/jMiERdJM26r3LbvS4/3NfJI0Aj040D
1YjFcY7tPl96xW4bmw9dVYIIyLhwnvYcFHd1J/YX3M0A8s3tQo4O7InGazAuF88u
k/e1cdsxBT4zJcb8NMWTirOY17iYpAHEzzNQg3agzmdTJLtugTltIUddES2JhOiY
FAALvBvP1d280q4aufOahf1gnJCgvPkjHkncnO2BbPbhGrXAtezrH1LiveNJ/C/n
tqXMVE1BXgr4ptHvHQnpY4l5vNp0QLqS0CCkROKuT/H7utJITJZtDt7TmFe7RYdv
XNq8xdIgsHs8ygWN0MpkGUu27etc3vn/jK1Y2IDpChwrxbW7mSJqpl7oXiwcxsyr
DVv12+28rktO5JiYlLoS6T+GUANAGeWm9SDGM2SlY+i5XmICX5FExYSAgayY9Ns6
nVVPfrvWREUIrAau0PqG4kqXj4U/SZc/2DFCvNlWnETg8kmAo6P6VOcNMOHOkLmC
QDOoGjRQ8twBSnbbDH74XU22xnifypOXRcTgjPf5zJekxogYdH2Z/9aGH9WU8HKG
rtMS6gPC3UcDZiqLB+NVN5vUyJE+GYiLi69n7T87cj1mxJ8RFYO109NwEkn9fM2P
hwOazHWe4Q8tGIOp7WNfJUfC5klYQq01sX40LWL9Il/0YP/lDg9GKIAgitZ6oBVp
lq7WiifshUgSqsSgesyLXPk7yyfnhj0kwB9f2tjrPtrcQq8OhLAsPsCEVEskO55e
cXns0SKxUzSnc9MOgF9+2qfNcrw12R8lnglsFVqg0pM8KyNQUx0UactVh9GaXD80
zjNkJyvHJiONSFIvOR1mu10g9IRMhUznW4Wgx7eWixNM8Z0KLV5MCL25bLOKKWgg
LMAMYdfdiI3D9DMrMrXQEd6otI8j1l2UZw7qlDRG135DfLtDFKb++T8SYaLCTE4l
/b/3jC3zMNqgbMf+gODdkMQKUo42itqGuyJkgBIZCQkMM4w3eQUHEP786JKJKeip
HE3V2AJyN2vvHjks0oann4CsZrxMH3TLvA+RzXj5EyZLw7xuQg0QMPPZ1wyYaCdw
hJyg4a5ciG0ktByZn2iJ9b86g35UKwNKcMNc2BmobAly53KLc7l+FljwG1vtt+3u
46+2/2MhKuxaYiE2ZYM34N0ohWdaok6j5Ukhg5giTrDFkbxImEKIjYdRMCP1dZ5b
Jy8m8LGV3NEj78ucgXWp881cpsPotriUvVdYF3Su63IKKnMwM6hu+e1YlcNormkf
9CH79fK3hY96XPO3yRISZpZFXGpFQHm0mPgEGcp+S/LdsOubz+2rRRhUPrM9M1ZE
9gnT0BVyPjQv4/4nnawYCj+LpDCyl2GJhdcH/AiVkWnKGt8nnou/oN44bJVcN+fS
UwQ5n8EMXDzmzDuJBRnfbK3NfW6OzFhg3DzdLbIPAZIKI6R7kWUWwVEaYt7CSHT4
rsRU2YROCBL/T4os5Yod0wWNfHjPmS2LJKu3sIh4DQq7hwVOvD/Q4wfceCM0GkEa
4PB/0R74SpfI3OKDjWA8c6nd21rHp7m09himD+K2Drzm8qjV8+UM5FZesW+urKmw
dmgQwPJ8yplR4rItkuE9lxR1C13PsgRnq5mxNaT3xvTJxpOgrHGhCx1YpxSZIiFr
ZyEYAiTksl9uo51+xklAHUqZojpHzYs7Q2Jp0ucaDcB/q0BtBsZ4b2rEX1+93DGi
74fzvz7Wc1wpNhke6JghcA+9lplHmKe+U5TFjBRDz+FlBkjRLwwoi9Nf2K2qZP/D
POnhRA4xfozWgJuO3IHyuVljCyE+yWzY7Z1RiAoIYEFyhjHa+sSHY2Yok+PJ42RU
GNeoZo/JSlgDgH5U56r9RITkOnk0/Om0JfNkuLp9xxaXesfyPHj8frjb3EZkRYa9
1UWwFDFHkJfPltuebcsaKLDFfaFP1gFikBp7tEqMLFi8jKm6oIU9mu2nREG2c8Ds
6f866eL7ObIiMdjqR34DSFQaXwp6RqA/68Q9MfVfVqh2WcS0P/DxPvLU8pYBdADz
UKrFGf+19HSBW8Ewt5sF6LAzjtPF7FZaqzhs3zmiNb/HRZgRc9tj7cRXWa3yPE5P
UkkMrHcysL3D5+wD2jPGaX6z1yyuj6789O4CoAguMzONNBCSjENK+vgbrL1UPm5H
0Ig3wOPnlkpDuba+Btnc1GPUYcNwBfdIuB/+mRrBAa55+v6shg1jgGA5ErnSH236
AChlp27SCVsuEQoGcgOC32IrZ+3ClpYF+mC/Zx4xIOeLvgUsl2li2HkT6n0rDImQ
I47tAUkcecHYzqfFE5I34WRJWBqnn2y+MIPLbs2ziy1BGxMe73VrIPptJaO5pVSU
UesQ+KRqDLsiuFz5StwyqMfs3N0E3zu+swzNIRsfBedTUvMSnxyVcgEmlRqYHPBZ
QGlMWyisf2q0oERIgGSeiRuKNVYzsd2Fh6mU1Gs/juJ2gGaAE0EMoP40xeQIxZuZ
sUbOkvPwxmUtKg6R/J1QkIqAdrdsTIt3BongnwpDEub7caR+XaxZpnmRWiAs/kzg
zTLj0AbIE1PMcxm2oH5tE0yIvk3+RwsSxUaVSZfejJ/ocYtu2lnE4pcp5qIl6Gyp
+F0SEiE7JHnXrrS3O3fnoo+DoGG9JuAOwgRKOMGHm+vbvV8hZB/w9/AA86brIl0v
io1+zKlxn9PXRcFe58LjxEuia7gp2wtxV7/oKqArg8Z8x/vOnH54GFwNRFjf9oG6
Vzosq+2+ab+2fB79+nn+kUI6jXhg+QwfjMylL3UACYrxAQAkzRyNOcerJ6xAfhKd
+fdCnTfvmkRXm6T3RuHcQuk0BypbdqEYN87Y9W+UCCuoWeFXt3SaSkhwHAsNZp7d
3lsoEdTKMFj+qHnjKb+mZ33lcMcK6OgZgOnAoFqObzchJzoG2kdxCwPV6DOhK6+b
c2rg6Q1H8HgoOvN+kjSEpxQNHrklodBMc/DAZvUg9GndbtBE127OmjUZ3QkZxqzn
aEZ4/f47uY435MP2kMo9klSYu98ZYvZCf7j/ZaFMXIRC8kvkVXNwh8JLXliE1n1H
mq5gn0s3CoRooWeaKXKN0Vhiyj9qw0xESVVxTOViMU15u+W2jF2wQCGVzFRAkY/d
Ip0HHs6vG548A4iKH1Wys5DUyF6fUujVtkGl9b8YwGGZY/7o1xuuADF9ONSZ8Goj
lFp2wneJIOf1tQcXcaiu0Cy+S4IBHUz9aRptLJGLjIwsx0mt3aw6yAERYNRhpN6W
uOQzBbIwarAT5xOSs8DijdTskruLYmlDBkiUf/mKgiMyyrGF0NOwUECl4xO1wjk2
zJBr+rI6q9YFvYglRg/zSlhmyJV3kFpnhNo5i/KqzBTc8cywJgaJyDpVlFbR00ME
QqOvQ4YJG5flteEaXJLeI525i9H7l0iCYnBFxHwLW8DV2q5/bsLhdj4CIh6Bj0cA
+RRLtzvqN9djA2lb7sXOzC0WbZITMlg8Y4fMKR8GctKuvFOGuh2bcypQXjDmei+z
XCw5JJp82hoZIchKytPH0qJ+zhXpbOS67M6ThAZp53ERB8m1xoS7zQaXTfnEkuAD
UVMH9pvrD7NXh+J9BV/Ieat0R9v1HDczrWxZixNgqjsdmb+c1i8wxJl+27v7nu9N
Dkb0MThIqbVoqPY5sbznzREJ+EP9PJHtTHweCQRPS0KXYzHkasULqM/lZCvusXsF
atbAPc7kgo2vJ8r4ZRU6Q3pR5Dvj/srAGVL7Sm6W1zXZZhcPHO6U4YvkTSefRo10
AFU1ZBxgQ2Ir6oaiunhTvz/OG26eq6AsN4muRLPxviYymQqrn2nBOzb9oRHi08bp
/5lPQXczXllGz2RStRiSi0eRUKL0/PtAcD41ysn92guI4LzJgC9CDaol+CTOydBG
+J/zH4gzfePEe4OvGFfhHOewAbYmqmW274IMZe//Tr1+lxFCzrk7CpAFD++dF719
iLKNrVLhA08wf+SjFHZa6wpfL5FrYJdtTDtNiWdQSFwfTG1Oq6VW9aRI4yNbfu9t
UvfLzOW4gxqixaDJqr44jgQ76qWx8FCiGI/f5s5iIErJkhbLtlB0XgnZC3s6xjLl
GiVGYHZ5JF8U8Uxmyxn50lLJyK/vaUp9OnNa2BXOSjIF4PNkhC+IGVAfcqkWqhs3
E7SoMLZdFRWkuNu3RmPuT70/XfXD+/EmeugbCOYhqc4PlLZXOZHHm5wKq+Y0OLwV
S80zOgTyKiVrQNjFlfRqgtjJ+QVz6ls/fXKIlXLPLoHRi4qe9m/9C3WDaEyvhM9i
6L9lpcOQDM04V1jMnva0FKdqDawcXbMWeXRJK6CmNp2NUZ3BR0GleG8R7oGD4D7Y
hXVMhO5k+/UDMpd8CQoiScsnHm3eK1/1A4k8tnQl6Up9pmcoB9DfJC/0pTiVIHzA
Cg/GvcN3ykS9s4nmRuFqPwc9pSMh8HKOjEEOG7EYbdKMss8vDPlCdh+Tu7lXHq3Q
4+u0jX/AW0XM4Eb6jrzD20AsQRHIWKSB6DNKemFxiuhPgAqD1benRAzAGYiBHYIs
8TVydN2ukycbCP8TviGmVQ0UaUC6sWskSgh5BA0xveEv+78JIZ+Nc9Xac2m38i8q
zDfEipp+MR5HQEvu6HhkbsXchXHzxhrK8BtUrMsMILx+HjoCrWiXu8np1CDmWUV0
H2lm6KoNZ18gsOCBbLb9rEl7aYdD2FLDTz+auOtAuGkDUS/a4I7oKo2TGr9/MrDe
H9T9TsNBFo5nxWjLAoUatBughrfeOLwZ02dlgE1Do03lghfDRym0QpYQXl0Avpy9
UtzHBiFheYVsbFNq5LOCvIeSNgYp7QqnuiNDO7cr3oTi6laTO1rofI2JQehbjfH2
TZOu4H8jJr6f1gi380zrimWgg20gCexhovWTwb9l0JNzrDsuXrTNBSOVRPi/fP3H
j7Ls0hGmz/0JQAWIWbSWZarGXbuHJQZbkyFnuXRrp9n3cAWatpLvp+cF98WAGt0l
1ZCD0yz9CwvX3MV87XS939K71+lPK01Cij7sQPNfzEJEacZobay5CeaK9uPDP1My
cmUfGMGfh8YUduJPb2mK5GiWkMsw17764qrkO78BTXR3vKaqeH5NHFhtQXTj7odp
y+YrLmdJB9Nnm+59idNShOKTwfEOsDCPmsEmAf16jOXg03v0C254vMbNu2D2kyrx
Ax7gNrHvznou1hw8MO9G2/tieWZGpH9BEDEKE3iP+XmT40dsmT33iu2FdRjK3yR2
IstvPF117A0gqeyJ7wc7J2u0q+SntIvurmiyw7glxWxGztdFquHJ4Aqn1Nh68gyy
1p5CAq4ibkRPakd0gsoxOxcrG8+CoNTwUvC/yG636De5hVE/pZr5IScVtrBud73V
BOnJPYy54OGoy1piILqvu+rMKvj8VzIaOPFd1M/gQuVNZMOJY9RNcStx20feqP3Y
/jDuyHXmvGqEDQEOVmr6C6Z5o9cn0rXpchHrGp2i8pBIHaKy/aezENdPIcskuaYO
l7Ch778ISfEy2Bh7QNX0XN0hyXgo6CbMViWUFuwAfFe1NA8N7LK737kUF8FVSSvq
g1mvsFA4Ubq+lfhu2VkRzkwMCK8jbKFXXYyV0koJV2fRj7BG5JBiqoGByWOVHwYe
XRUGpmyOycAUhy3OqsmBcIB5CwPtSuN2nKqVwp9ISQhMYnp+JyptRo9zKvXugMW4
5WGUC/t1chwUE8Z3WW2C+67oxpq0nBXqryRkQKcbZKHlLtl7Vkv2jwbV/bpUHCHc
qxSSVBBnXY6/Q6MQv43DXLzdwQfszj9f4pYO/pSHADWX01+TpSIXlbWU/4bmHHpt
tydlEfTc2gXwH7RTQ4Ewihlmr3mwNGZgxTZZaJKqwVxa//Z7QBJmjDJp8x/29Rue
AC5ZTQJW0dnBqJClgL3BmKVKphQwLdDGVo/vMBLAXwFRMIj3G04PLqvkNj9IAsmk
qmPST4T+XFWTOXCo8gj7zs6aCB2ltiFdIaQPtf56q0bjSifGtJVSVSIS77EvnsR/
JiqWOzEcRBazU1EWUVF/ci1HVTtVIHQKA/uDB6diEe9QQ83qi6Jm4C2KZd2E/zsf
3B3aDGnIuRseKNO528uBqpvnfRWligSpJZ9d8bD/wvqNy8fKoVmTnnnIcvHOTNvM
DeVSOPF9zE0RP/Au6+FSLiouS5kLAi59oucMytDnRFuCHnKUaTpxnVWHfT8t5QUI
7P2dwaeVWTwxzu2+13032Vs+Eq8cX765JC1OgHOhJvR7uC1a+ly0xBkuAH97fR0o
zsUelfneiRDH/3GFiVCFspjcxiR2cJ52WXrbNqDWMkeE/jNMNzDnLyZYDnJ/AyLv
votQT3Gh0qbqwEJqRiVo+6AS1+D/oR9QgrOnOZiSy08CDVBWXSBsJT490Hvd6voF
3hq5QzACbFXNlCDJy0+7XSK3KfvdcjqKwPwYYMr36bH/pFQk51d7p+3SGP2UXSAD
D1CtsjMrb+GgmZJPYCm74TmqilGhFy6fxJfaRLfYoiqe3GjNOuTetjLW1Xa5ND3i
Pd3XN/tStO1y6xGKEp5r2jD9pncH4E7x0yuUa26/biG9/iRW7MylwRLkkZKqNm9F
CuRcOApN5wYOE9fsQRDMCHSO6rrDqRJUjnYf1Ka7nNGkyC4F6jK9vHQX0RprNneI
5+PbS6Y51/jQxtDo1XmTxAtUMEgkgAoJOcvigXr9Q0RSKQiRS62OTtQE9+0HJeJF
uxr1tIOmWikyJbNj/FH0gX63AcEcKR1nQ20hYNXzNIddT9iZdPXJxGC2zz+OyOUc
iUo2zb9fbbflRI22aLxBO5viZ7nTRINeo1q6IFe11uagTZy/ThFJQa9kcrcp8Kdv
A0T6T5fXima5UusEescGQ5t+968IDbryu6xxDsfZzL5WP07R+pKQXauiosdvwy1n
rxWy/vmIqI+Jsj6D0cAbp8dOzHxfgzGdTcwD1aweySjPcrm17fzihe54j/HoH+dc
OZKDzg8NDhSXLeUB7lMIE6WaAqQt1KVbtK5sktdGp1fjburcI3yCtJSoT3PQ4oPI
wTDkXq4BPIFlbQsyRAsPzo+WZagMYILQWqMUrmtKfQXsWvYt7kY51dfFIpFiexk+
SE2A6TQDoZrc5vCrsT5N9J13l9fxGRnrEbR6IRhJCx4UoaIctk33na9KxUC9TCJT
lBU0pkgBB36PuRrj+Ar9Jafo7t7miCokTMimZmAcfBk1/gklmHVMw6WCJIUOMNAz
Ixs+AwUIDi7U9r42lJk+kW0eMBpDtR4S0CVypX3nNn+8OjDugxnVPmta7FnRmgzR
iitkJ1Ibfqdkq3VjVixsnXDzrhwyN7pXfItAGgZdsv6P1ovMboKF2sQ9xOnq7yXS
Am+FUIHok7lGBJqgszBlhbCRm+5wUwVRnDsqfRyEHdF2SjiPx5Iz77xyuQ/3cnEH
7aZBqDcB3XsqptiKZkRlgjrk1eI8Hy8AE+DNwzZwHxf9VGTzw0rUZTt8oVesBUom
sAtpphL081sW20+4oX5XMFVhX5GViCtPNipPN2xGaFL8owhtIaKUYp+F/+1V7jRH
xD5WNO1KVDBa/54xoE9r4hP+vJDlDJBhrjRcMsAV/O8fOowu/LwfmfdE/XEcoJai
T/pyxHO5OyjO3XeNz/T3aogaqb4HhT7jVdHes3ux5dEVQEv6UttUuyTkkVi9eRCn
N1lmNRuYN2d7MS9/TzS3emKw4OEoXHVyivC0vvSeWa2A0joEd7zOfdYl3Qchl1ME
GDE7vHRGrGVH7kdZHng6lSzybMdaLkM+U60H8FgV7lDAsrMLsvVPWi4oD/963VUx
WHMWJTgEJlDQuxeMni1HDQ0/pbzK1802Lz0EYwtUmH1fMdSJrZ8oXgjv8zsQ0glz
OK0gzELeXYD9y/06WoigRzpZYw2CdmujU2h0uEIY67J3O76WZ0Svpgf+OCP/6/zH
YrLB6xSkPahbxOqkTZfEiR+FDoALDZ9TrFp4fa/C+qDkqncz6gQJLIEXRMe0OplC
e5C/IvX4c5mSSyEDbkN2E+3YjkXSYfQkhojI7WTiS/s5Fi9j3wX2zGFv0qlXeegy
te9YFo/LaUTfvtj9hwTDoUQbEwa/sVtBlifg6wY7S3DOrPlgFmmueGAW1ntOarCm
25AUdmYfr//87iyG67JqcmgADPUpbNH8wvi15z8vP1QJgIH9CVPZnVoVxgNrydg9
1VvYuUH1RtRLgEhkoV3c/iYrMymStjS3sz06I2mUzXJyf000/EG5sPdY/ctt1Pfn
h+hJAKACZty67PiQLjC3dRTND9tUjUwgIy/mZDM4TDjILGNkytpbrym/i5f5uqbr
R+QSd0iGm2iGheBuPIG6+JFmRumren+doYD4xjaVGq/NNk+HttXjuF12/rpvuByW
Uswck+na3ItPZ9CjoRkcaTPuDs4UPAzk/UwrKgjLVzXXxawKgc4y5VBNApph3EzY
gUdqQnmlQzbcGLn8YZCXacybGVNz8DSgcl14np2iATw4Rgi+nxp6xRh5MQI3jKFz
w01v6tjHu9KCVobyCUTOT9wIfQku95zIVr71DBy/8FNlwNW0SqGXdZ/IsaxgJ01p
HaLOe1QDAT9lqFbKgfMl5jGT59fkfxDpr3o5g7rFPzi+x+WHKjVqhFf/SnzQXBB+
gqr5qiCtL+e7QO4JcNI1lbWm3JW1DLQGjPfFZJIYSdbyKH+AD0gTI1mn/PuG3J8o
CfC8votrvfJYOpCFjdJCXXzySWFhxIsWP5LZTzwknuBeApIL1hxF+EeLbno8ae3Q
FSAUx0tALrwW51EQ/bAPIvrC8aV3rosBtl/T4jtZTfN9mL7225mouvof7xc49oB8
IKnIsPx/4msBQRouw+KHsEOgiQqQumzOcL0L/iMxeM4M9Rpr71hEUdbghm9P1bEt
sASKn4f73oQ6HQyBRpk9WPl0jigUZBIkHuVl3mSoRu2TOKyoTwILSTIfApcoqzxB
9njLFTVuVEd9Zkj6gyjIowb1Z0qgaMeqWkxfsYFfM1k4EjW/XSxBskNrlDXVfDIX
+G5oxD6i/RqXNOKfVPwzMBa2kTvvIk/yOWPuR4Jdd8tuM9jgSsmhSULWKs1jHwnw
up8oIthcxrTkk7iqxP8nZV3sMYa5aeEy2Qg7BMhFQ7HxLtdcBHG10zOygRTakKf5
bbyv550vCkH+m9AO9mOev/o8xoPCVZeuBMvGWowurDxoGwvcfmZf6XPEOho6CYfa
K1ayhWaWr2ov9mP7vj8Zblhxh72WxKxy/gxV5shgMicmZznTbCIe2fXyoW+R0JPF
M/GQzIkHxVYvjwrKXnc9ZrFBKOVzyKwcMDRu6KLR2WCCfmkzcAKXkgg3KB2qhUka
ozXY+0QGqLyR5bL8ojCq6vdjFvlrA2oRI7NE2feFTqaGy1/aV/ypUKb2FUEO09Ci
huqiNyth9sXV7k/Nwf3b5SOulEhIrKplP0z7djmKAdLdeGG/Gw998/ArSXokFoDV
RNCHNTMtqHLQzM5DJFGRi6XDZrUWahdRwXu6TPhM9eHrjPxPaPU+Vr6BNGgq4IYM
7vjHT58kGX+IgIs17EGliiqU4NMFMbPL4h1rGa3LSBbkEOK6o/93nHRipnCQWSF4
1097h1hWAeWwWgt9VP5GlwD2VfxRrW2VE3sBXJV1UfyekhGxPQ8nQoxGoIh6Pbd+
tMKp95dN1J9eEUbcY7pIGHV/fggPR252znS4+w7B7Wt0BlyQ8nfAXFfz8Nen+y2x
C5oWqZSsSMbODPHnMfkfYgm5x403hX+KCNgf4icxQL8QiOO3YvkItLxfOAU6Vq7p
/G3wAU/+vYrF/whRZRGRr6MEk5nZBvfokGqIPmwrjmTD1z8UsD6xH1QMUayEtNrX
cCf99do258+9oy4TP+aSqZuNMPs3X0xqe4TDsaevxHg5OTHaTUaQ1SyE3vDvyP+z
hvYKV60uUF5r0qeceZ655fMJlNw0Rw0Kazew0nhl25eUKM00oia6zFmHpybgdk+W
zWbNZkl3jmoHsdZNk0gWhxrQMBdYwZRxOD1jNFOj7UrJsnI8nyuJpRMsjG9yiQnO
jKE9sw/aNlvncWWbKmQF8+OxlqQyPAMEjouXd0emD4X19g/8dpK3ijG55uWvHGaI
cDGXLOS/L5wFJKwn8ynaDrBegBfDt5jDRNWFXUFzKxJkfNspfv3lohPQKhle8y97
2ysd9F//Tek95SAps/UayNZrV+jR8k7LK52rbCsfWRCEH/mVcADMdTdbxTZztTgd
nTmPpea2VGvOVtNyC94elAURzqz/Z9oKwCBqs7BXyoup+Mf3Ppij1FlVZ09MPcbY
PPdufRGmfrx4G41bjbhyM6rJhSealkhALWS0K8LnMTd+uHe+gaCjLKdg7RiLg3Mg
6tA++5XgQGGdN+YlvtEF962v5vs07UfOPHNBgMiuDM3gARgbspANHOSPLpwA4JD8
TPIcEnGJYyLED9NS376Bi8EWEWSV9Iz4rW/p7ZQzAdeB00bP84GJ4C0MQZ0zw4oM
DVZql+r1hCAfQGzeZpEFuE2vBgsaDmHaWGGqr5BJmyshVF6i6OhJtOKunwjYPLj8
y8kvg8YMhHEoAAGDBplbZAEfcLjAou1xUJt4ZzZ7/MzuNtjaFncCBKDUCfbR8hEz
4J+BMmYtCFVowUZIovZH1DLRKgfIPNLE/GLU78gNdzKwC5hV5SNwPSYEl3JUq67T
0sx0yc2HvxqBn2N4UBAO3ZwwTGKlzLL137Mj/oooeUjSjazGP7V09T537yRPjeqO
jij9iY7BJ7t0L6WwSErW+edISSfNmV3WiQ5Z37XIGJgTGg/2alIsbBeTspC5EmgP
Iirj3/QS8kNqXYunWPo5TPUXHtm1WKORsopGX37tWoBhY/WdF8Y1nrN7IjJMBHmZ
ckWRPJ4nLB364HVcH3KnXxXsT6rq4l9aFmVteuX6icvgn1AUU/PF2NIIHLRtxMXx
tw/B+Wf9403oZ2mEUR504j4eYkPVZ11GtdJb1A3r4WuoAxIrstPFIMNGfnbDOCBg
NpVQv8ERFH2dUltplTyezWzloTx2nhVGNOx7+sq2RrdyxchlqQQbb95PjlTpGqIj
+Fg5i/Wlmhd3D9vcjjuj9x/3Mxn5pL0fpbJu+6MuMycaF1ASMOu5vTf5uxWF3H73
AFgTLIuriqqI04eDbCys2MviUkRsXJUatmJ6rIFwa556H7np6GI8ikb1+krZ+dRM
Uu4q5D45F5tvOEPv4kpGgziJmWRmlIn6zdYDax+lg48eH/eihKmg62TegrIzAHZc
tCGr/Ont8coDnr8EEvQk1cBk7zkwE+sZZ1atDzI1DPGugTXoK+OW0smVLji0f3/P
8jrQqcZ8LisWTN4zPqH9DnHs8Jl89MjfxPMz6WWremfI4LDfU99baTm6AoaprUfA
Mtk8uMqvqbJCmzgiYiyxgKAxs3xey6HQUYPaQvzCTsT46iT6/NBlXzKW2f+0nekr
7wFRhBuifmYxF07BvF84S89C6nzlEGEGLjWAEFyQ+54gISY0lRBoGI7HclTRsVLH
1I/btM8c3kmgm27Dpd4VfQrJwS82YxpC2LXsTNcVsII22ej+suvo9O4vExtjxB0W
NwrDdb6QgoJ/yg3qA0syr2K4brHS2m16CHTJvjNtl4BDJVv89aUd+iQUJCoEdosT
0seCoyjnTrAfpXxCMEKjwBPup7m5f23zMMFIAGxvixTpRxi+IP/76/wvAWd6bUiC
+Kv1fqcpaMNOCI2sqqsScZcp370oXOacvBuV5wJYR2c1lG9rCnYhmG1HmbvgnnEC
EvMtZ3lrsnObQ0o7J35iVVQuuSMRpPcYr/iDLV0BST6JxItmiXbg0mCnGGfyGE4/
i8ktS0KGLXoVzQ+RNzi07N+A4+2ZR3qXJCDvdgbAu4vTvaHhX/WDwrh/M5XJ6a8J
JrqofeskZ2nzBd8svPJ+5cX2RIs288mpUksBKETSUD6CKbPrMjPl26gdFaBKOH9s
5ZWK1ANrACOXbYBKbSXi9+LRwmmsYIHB5EMOXVzVfwk96yITvMjUbM1uB1QtPJua
u9o+OpBGuwH5pIv09dFisJCLkT72OHqOejZi6qMEKThKa5iHWayis8VCtatsAgCN
h7N8DCGBKdabyBEI/bDdtCn/6F+Q4N8h7dNoYdvBNqIcyMY7zPgwyzBtx0ZXu6Va
bkEo8QImHrjOwjQ5+ygUrFW1hwxii3qqxlQbvN3DG+nqfcHb1jscB4WTIG4+x/lb
G3Z9s8BnelSZN7+u2WqsikzEwSstnXpWkrfaN5lPeQR0mOCfAqhJJjX3L3AaJYBR
5uBo4ICyXFTkLO+9nwy+DzttOJqmpIgKtfq1eZe2IJBYENQKuS7yd+MBdmNOqoZO
OSTXfWseLo/736LeCrmJzMS9RCvz7RkQnSiwF12fwRjMo3Lc78JdCEOpvPzA+MlC
VKzY3FrO8K7Q02aO4Wcoh9h0S2IRFgGjeXWPqdU82BX9AOI9pvrzJEEyC+ANwicz
2qJB4B3KfXisplzdt28gfyH4f47hqMwnYv8G9nsekCyNukGnn1big/0Kxrv0V53L
G3KzFhYt+Mnht5nSywjznrTImfThOBnLcc1coa94szc9mJqkMoRGRxcjiiYL0PHh
hUyMupOyAEymwl88LwRmwLD6AISoHWeQUB9UZqPpt7WmNNtjNP9vJU95qU6NFnA3
KrX1uGeq+tzZkbQTv4x0OmscREMqJFKQ/z4t2wErNaM1P20c6lKQRvE5xf5SUg4R
oS6JZoNsnZ6MraUoHq2AzYmFPHu/wohj4wm4K/SAIgSpoDmXHaYaa7QoAMbwSi/q
zTLvqLPviXWjb32Vv4eBjcpHSjToFHkoeTbkgRyu2U0nDExrkWja6IkEiDZuduiN
jcjWDrF1uoYWXms7QNOt4DtgrLG5kDt7ZZ7Ah6tQdU8wwiieUTPsuUsV9grTPq3D
vK9rjvKBJnfKMAoWm0VsOBpRFo6u0ybOEzXKf8csL5dXtip8ChFKrcDvQrP4sIc4
1DjLlTZbkE2x8/oVc/Vp2ea5WN/Hwr1ygBFbcfbNxImkIAeT2NQHzCVHasB2fOZ0
04+u0vPDETATlPAU9BwMl1o9xDc6Qe+K9DrmReG1pNQFrC17tLIBwM0mSU2g+o5X
fH8rtNd/001taTTVWZHPTJal6JwfSB0uvVG4u272Cu6K4B58pDfV+fE9sMcCB6vf
KX3ycqor7nufhYg24Iw3/X6c6A8uVJUg3fzSgrP4Sd/5q1/p92pzQb6763NKOc2t
aBEi5GeEHRpp95k1PD1Q7oM2r1e74FjG3sTjVIfT00bpa4JEHuOas4tZz+8qqtiJ
XRSi2ghrzT7EbO+r4AziruXtKgwZeg3BNDKEjdvEh1bEW/XZ8nsgyOpqUE4jppzE
avWXnYs29Fc8frJugBm2KuDmq8ih18IN0NN+SOjqzqy1ohuNNmZszFTbyqEDir/s
rvq6WZ+7sDVTvZf+cxdSkNzsiBlUFJZGa1xtFYpPLNsKwD1zBNPabspDz+ah5hbq
QLaTZ/4pX4oMX83Ov/tVdI+UP0tRG0p01NpahRHnZz0iN9kFD9uwd8cBSq4saWOP
56uNEMpyNMiIzUWzaEEB3Moapkkd6raThuW6O0i+v1v1SGaTZfBamwfl/qwVpgQc
t3oTyaB2lrA7CRyuFQhhrlbBnEYWGlbJj/zTjRzwPB8+cp662O+52MU/hATIH4Ld
DLlYgpyBcrEInfYoAm7cyVn67Nahna/quespEBp45hYSPT1CWYos0lYSm8LOpGtW
tV2iA/boW5DZlZWywfLVR2sJVKGfnNsjWYtUHKPfKOLzMsSbJTjtExBVNuNBbYIt
Gz39tmapLrNwr9y9LEXZwAX5rpzmFdNJsVq5EV6BzbVCRp2L1L6VDOkQAtjSO1dQ
M5LXb5Q+WngHNEUVCLoOzJlGFiH6wwvLOW7MUzp6/LajxweCja7dEdBx3q4xAMty
ftcr/6yx5Pp05xwkV4/mA+biu9OSmhcdNk9njvuRMshz6V6kYKd1UvY+45II433W
zN+ujzEpsTPFG0d4Z1wRxjPPm1vXpXmkFphhZvOPkZRJSUxxphuVGJ+Igg8RNsPC
xpOYzC+J2O7h/ZkxSkAeDdvsrSTm1FPraWz1/noPtIug9adri6Pg8AFcn/0SfO1I
37ANXwlOuXR1j7+W2sm13J5l2+ojmg+BRrXfeXYxPHTO7/eHmm+4XONv3ryYzia2
E4EzR/9FcV0y8KR0TOd6ibe3OS6bXKTDDCh0PD5wONx2+aZqSMuMPNPSfRC3/qYT
KKdVCHgxwSFIheZvF9Im1o9CeFKZPDeUD+8pOyzY/Yk3OtIF6EjxtztQURpbqugy
EpjBWtM+4AOXmjsELxGauvfrPipf74e+TdJW3Qt5wKumOv7AQZuch6mW/GMlpTp7
1UvQqAhYQazKxWQk7H4JCRuehidV9gMgIuz3LClb3atmNJW8IzgZ24TeRmvmdvV8
i0jqWj76k5LJYg3onrtrghbZPBxVFnaGh98tE3vMyhBtU5Au3s0EAPNqMWiBvEPc
WYPolzEunDPfHkqUgyCfKpR9/rTfmTtN5n3Q/PsAvTYOJUXBKi9DMi24O8z7Amwf
GPQVLsilbxvkh+WHo9d3e48AXgWf10mvYNcK+x+gMOTkTAHZzKiKS8+9GcxgIyne
FoB8mu4Ob6SPL7UCpj4FzsBl8QvJtBWJkTotzZWjgppAdofV6AH1cLRNcFSK8S3L
fPhlW7hA/B9W9zSE76WQknXSo3wNFi6NdhSa6qklTAfTKQ7XzO91Ea7n2RCyoGG9
iLFO4IGFGJOykWkf7PYngfU/Bgftt1tYX9sAbfgip9ktbBZlGWf2F3HvRU4z9lp2
zo38EAAMOJKrem9DJnzZRE1zIMXX3wVALYL14PoftgHagHyisbXjvjZt4Gq4IOfu
Ml//bT0AL+gl4/4qz3Utscd9BUN7HiJ3BXarmvcFvCyuEOW7zMV2E5UAXQ+K0NGp
05G1mTuNDE79GsL76YdREupFAgfuVP27acD+XUt8jYLHXyhbqrsYMVqXD5sfZHjx
zLSwxZbHYilX8RIicGvmIElBzXj3IFOw88jat9wog8dPoHXEzuYMHQ9TsHgFueBB
ef1LbISshIpbDQozMK8YT72hIyFeGxKO2t/WqNZygty22rwrwcthBZK6JbZ4/wpc
mWKdS0dUqVyE1puuy/GXDtgh7JqRMPt4UTrzuYa9lLTKwz+yEwOvaRShRawVTyTM
2L2jBSA1O9tm1CcEsnrIkn71ZkWpW1P09weOaYj8U19laVq/KkJMiuWUxKr4anjF
kdd5d+qEt0uEb3rbhBzK6VWY/pO3jMPTeVn/n5LeuoAl4UPdWwVKTXWAlsJ3dNSn
De6PPG6po/Yu27zWgj6+kmabxoalUDmAl5EsWnki4fSv5uCJWRptng+2GPUrIjjE
nLTFUhWYTbvr6aLm6kNZ2QtXC+M8CFbnB4UAFbPalbjKQyl8fbgJOYfamoZCtWYc
GN0MrS3RIzdbz5Co3TVCfXuIluvGb/IejGxB63iilImidDA6tCxfAEYU/5JnQDEb
mQsfB6piYxtE9G+miL9z5z55kSexqf42kfRzsYHwvG5hN835FiF7vylSmnzfi3M+
n16WswiRnBytv7RwdlxA+AIFR/OrjU7B1VifmwUtl8EpZo1wNRM1MrCqjKFgi7yg
79r+bUe1YmHAx1/N9FH490W0oCy8l6ia0vsQ263Yw+E7CC88DNlrkXx0YtONdW3c
geyfmAraiDhKB7a3U/y0Xlb5dhN+iZvSj4IvVJduum7VLNY73lWkZQ7Hr1EEBuN8
GrDS2wOsN3nOovt3ZgI9tc/bFE+Cbke4UH/kHrVKlx9IyPRfF2VT6vpFeuiQbIrO
Fi9JYWuMf2+N9ktBItBYZzk7T6n2O+TDaFr9jW8wQEoaz2VSMfIY3qfCv/lsCITE
hsIUtmqUNM5LSwGqf2kNR4yFOk1KMxBrQttnS+J/pjfUr95V0zXOhyraNbFcpeQv
vmSiDSBN7BPgbPPmHq0JEfU2laq946W/k4XbMaayfTLHkc20OtHAo2J6EOSGCFfB
IzQfHxSqcSRw0fwlY0yTBKzxzVgQTU1C1iUSSuLIIds+Y1Qkc0+8v6Y6/bM5Mauw
GIxuut9LWnwaiLxHXfJ1anQrduMXQuRNm8CR7W70Hr+4X0ny1wswgYJZS7zW1Udx
S9PvBn7wPXRNpadVbrmi1pQrkiFJn3Lyux/dQk6OLy3uQtzGGZBIBYmaLlWsCs77
H8sXur69+Zw+WeQXPsTUV6Y26KyjF6NpJku7JLUWjAR6XSn0fABG7ljLQ7CBfR31
yPMCrj7cdHgZ7H5tcsSopLOQb3iHNACc+bIeFHP0PURX4VBVFa45hnTkIs04Mm0z
Jy/yb1HUlpGynt/9djMZ4B+AgN0u0KNBGPXT6/dJ6ZtuWTKDiBSuVeyzZFpsBS74
WC+xv5mtm1xgfWvktQ/VXqa2SiPs0KS/Q7utMvMH9DAIhuhdfgUg2xB4+bDzzzZ7
uZgyNC4VaTFIS4K+JSyF06NGsNVYC1hg491hQwfQEtJcFan/5Mjj6ZUNYsolq95k
xMzFeNBRK8M0fs9nPFug6cYJLLZpqop/ansNjzgQZE8mQql5Pk0aqNHxO3TIOZgY
1cu1y9oN3vFb5IASz+fKn0X7Z9NiT6TPmvWqwhZ+tAIUY/hvbBDZuOOoZHCrw/02
gywAog3wJLSjlOFl8cUtM4XGCywaTsA+ObA1aueelkZuHprxlndTwtc/Aeg1v8G3
7Yqvn450QaKVHvUbZR/Ucl0u/2mE+A02pCkpEl6N8WBgeUAdJ709RB6ea1P8KDpK
PvevmFBRlS8SvOo6T+P0JPKPD4FPmU33xvoyh/8Zx6VVsegA8PqQf9dUwFOsCqst
kL9r835xfh8gC4AaJGr7qetC3VLoRboqp8onDvO/82pJVMc8tmsWIW48SBBqal5X
n9xPPHxlt3AcBaFzi7AdqdJTJCpYNeX1c1pD1bTDYd77Zth25+s7NVInShodXTnT
nR2HP8E7dewFWRxjLVNtoNETCU1aaq++odeKLpbS/cR2NE0W/+rRkpAWa4jUGvb2
acQZYHPKr2ryVHXuSVgiAAu04WbqMUVGqTxb6ThogwSrT3Ox2sSRv1Cln8K5KtTw
t9EQu8ryO7dYgmuBY+a1+X66X7eUvZ3kPhVCDmhhqyUwTc/l032FgCF1qvoVLSmV
ijPXMk3X7km5x8zDcPM6T61D1P7TEud6OXx1/uMYU6iT60fNH60bb+gKMBKf5W07
7POCUfZM+Ov4yJhVjEv7q0SuTdSj9/jfzDtc4GXdOhkshNju0AMvYAdms7vk5j5P
GOLaplB/RTgIOaStbwN18tceXgjffKkHQdwAD/YnxsB0IhAa3ywTkKV7iNcz1X73
DDmvsSooCBT6bBE18NMAPDiUkdangx/T6+dBM+fuj352NflOIyFSbVdRxixpYQ/2
z26X1vWQDUNPbm+n6tpPaf9uhxNNbciZRhgmu2+gtSG47xTF3i9f11NDvolzKzR8
t8Vo9GI26a6eBc6LRGyR2/l3016ftaHU5O9+3ygeGedxTJpFSRgRlmb0uvUtF7ba
cL62Y1HbJ7bmQ1vBMjoPlMSEnEYEoRLblSH+PC9Uh1yt5sz9oTJ2lSkKzdfjdAsT
6vbGfUtyeUI3Tp2sukcldw/7e8CtzKXYyOlbIALGYyOyokMBVhPu3iANVbcSSPGg
P3vN2dttv854RyLasjtwEY82059bST7K/xaujFUxWGRWqKtNbUwVZy/QBDah9twf
3lKJtaxmFkJG+O64JpSFlq1OrpkrFEi4jRqOGJux9QJ1m0z1ag2BCFL4P4ooKh9N
40yjAhEn8yckNPozI58XecF5LpVLHAEufdjVEa84edaEJdVvwdYfVGmsdAktImc2
mc1mBLHzxKUC5EQMnVGrXMHKNbrM+st9G0FLSSUNLYZ3IjiYlt4gIL/u6MidPvTz
n8btP2HL3r1T0CPkJ76wn0ZCrLMGc5FO/N42kdm33ab1tpjDCiW98PBEr4offnvP
6jwVJfnHc+0G5/uClcY3T1OvGU2CmwNQDV4/1SxgvPIjOnzYVbDFd4ZPcPDc/05c
p5M47X8BTB/hGt+HZx4vLEbBF7rjQHknPc1kWrNZ8O37R2B8+KNc7oruHJByVT/1
aVb4PMv8BBz0akBW8u5YmC0hfycMArhO784GKnTwPgo+L7AzbJg4wc3SUlKvmEhc
JpBg+XalJoqMLDEot7igKp2qYrVQNCtqSuXWVFMVMmIi4OZ2Q16RzjYRVk0qLZu7
+rsta3oLoHQZYof0LyqrkStjA0v23GqjwKMYj32h9LLvkvenpqNSI3GsYIsxAbOR
k9U85Aj6cEWPkdRog4q8erD6S91HRzS5L8l9xr1tyyEhT1ywLkwA4jN8zOwFNCRg
or2/veK7FJ7vgPwh7UV1i96k+I/fwoUEuL/KJPseMqpnlWGbqYkThgqv1DiesxIa
QycG7+kcdvbWE8uEq7S0zkLYt5Ccu8VXOYk2uPFJYbAwzfHsSD6F23LbZVi25KeA
lflQH1tD+1tQguFRnEjgsw6X1+/uG2vb7QLDcrqw1o2KKv5yPq3VKyYck0ErRrdv
X6GgwkxS+LxnxAaeUrRwMdZdDNm/VzryOtc80laFrPsqjAGiJpUZmICjpO96K7wz
TKJuTRuQ0TBXa1E4kBh6CMClWGt9la5LzSTpXdmu+leeA08pOKJLZpn8DRhkc6AE
+wysaj3zKaApa9EWdxP/k6ZUr+kOoMMOoIsaiZCDNI8ayPNmXsTis0ENyjyT1Olf
cKNPdz3nWoNdaT3bRL8kCh4YwM6uxZXueVvyt+9chq8r4AGZf9xHOxOZxJIloczH
RJXNM1HGdBiM99Ryz3r91hpGfpXkoIv8suD46O/MW3jNBECd2yzbwq55j/vwI5pt
R2igEuP8DhVKFMxsTbwGF8ZjvL1EQ73YABlZzLcM66Hwk6juDXjsyAGZYZvZsiz8
85Qqn4JoD5vWhPdW+L7q2k/ahdGU9zdTyYTnGvSMiHg62T5w+I7TO2RW/r5y4eZR
c0jZ/eqQ1CYbbjCOl/XnyGggsy5FemDu08eIbFecgNV67gHRxY9XytE5liOUqCsO
NkDnP7AcSgy6uOo2LBjUdZak/5WNHSLfO/dItXnxgsL99ilbbml3J4SutPWPT/CZ
6UlFWQx9sh3VjggoaxLDdTSbf5RU2AnpW6mcGm7H1ewF8VgT2b0aMiHhQ0Ct5Ewk
7RrreC6yI3HklltnweC4izzcK1Mvdu/8apguQLBPX5YJV6VfrIVYfhkrzCGtgWZr
LmEt2ax/FiAAR/BYuCCrpcEW+NDb5wk4/J6GSfNzA2KV9pUD7yUBySQgCsfn4PUP
j/VBtMq/CcWhJ02Zh4mbvueVPvJOo7GkD3Z8qntkmBBDtD2lzLF9cp8n7luGd4vo
h5CJch6Vcv4R6zoGTsS2e3YdCZEfvrLLkkXoL8iF8cYxjK1DyzabctMR5EBWSEYx
d2k3R3vgpPCsQr6nlTurB2HB91RKoTvWwGMF9Y8h7OixYaSIT1ScQVy7sEdGJv7k
SqxIUB0nTw8n9j2uJiR8nr1WP5wACm5nF3JuO/qEQRYAz2gXqGp3KpbE5Qi5Td/K
lSPEqaVFzreBTateFOZwm2t4sye3BCxGw8mAZVU3yw71ve6/qvxzb6TcLT8kDfn8
HoWb1XpLuuiJxrJEyFndQte5wdllx8UeXt7n/wzMmKBZR0h7WUE04lV8YYWBk5XC
6fwSZZbkVDH1nyonjlth0339OKlh/hZ47sxAdt6Gc0lx1rqytW9psQK6XXiWVWBn
u8Wae/e2OKtvCVrYWZ1DJVT1NDIxNuhN6LLa3AaMwJJsR4Ke0hPZeRF9QqvidQCm
epuXBTWp5KZsRwBpn61bLALkIpXYJmTWSuX4v7564xFAZP6Pk7641BsZciWsZYyS
JlkDrHHCDjW4V2WThZTMAwVSkOLKszoIqXrkNmDfJpk+U0rSUKhieTI2KSVrC5Vk
jLmy3dFLHlhCVl45nw+mCVSExs+FH2UltdH0l0J4y5ZDhIC0ZAKkft7Y4CZf/RnY
d6PheDyWgEuDtiZjBcV4C8l4P/YrHcHOFkLFQeDdmeJvXF+pL9seSJCVDdmI0Ok1
n69g5oLEUIUDqXbR+C4FvkDPqhTihUGaMnES7y9gjlZFxo0dVRqD9Is2yO0nuxS+
ql9Jqan+3c3djt0SLFEspKsv/Ry2ahCQRzz1mPkpOD5/ZEf5c3IqYSVFPiYPR5ls
j1BwWqPE7JLJiU0tGrO9e65Zh1KeUmUyJN7YXx9XRBenBbOfPuR3c7NopXwhei2Q
Wt7y6J10qffUZsJ2ZfoGEJWyBv2PBPTycaMVwdVBS2850QnD4tzIasgPLev0lkd9
9D2yHxzAdJ2vyhKhRDiNFUKfCzhjsDpzymqnAN8YLMC4PtJHeWiRVq2+G5nJhPHb
d28J8X4vcF81NrFypm5Haiaf1eVAmNTpwHgM8Et2UJdyB+iVS8a2nftv34d9QD9b
BZzijpJB6mbvt9SE8hbut6ZwUxYQ0wXsrosE9XH6oCr3LVsaUQIHXtma5zp5V2Ex
t8X2Yd0/k6AROLO8vBfNH9x21lcc6m3hldsFqTShzAc24l2wQzT1XDLDMPVcdwRn
Qgnim+g5E7gHIrsjITdOk5s2ufNYtk4RroRmJxEHx9jc1gNfjevi4xOtuGs0akg/
0uT0Z1PsXEKprBT16ZgUr4+C6JqEyg8TrGh9xA6WX0nPOEjRD3UTkcagnM4ZjSbW
pInE9Wu292TLfLKmarQA/AKmJCiS+7rk5sV/lBWuVPy/yeLx5WqDYNgAxth+RsZ9
JgtAawhnSG1j4wO9j+WADc4085tlQvIl8Zq5NgennFakuVbtz1v4ltgl6hI597Bi
qXSoEz/s85nyIVzm85cAPGgHscMTps0jLOHH1TPp03EtlhbBhe1RoRCGWMJAka5S
ZJuZxPfAGxy+0cdxFcv3L2FxDJX3mx4qijt/JjswR1WmbTH0B6NWrR9L+SuJbVCf
Q0GWhPiO0+gz1R80SQzht7tncJYN1V5DG37jj6EDmBz7cBiG8gIMcMjEhKmJUfzj
qg0xeiAu8kPWB4tzz8vCa5c1wfUIOpNMpzaY7TWbiRGXKWgKHnNoJGGBHd8Mmdb5
p6y+IqmPa/QboC4Qw//ANpRYT09ITME8c+OmaJorgr5u/t/HXFif3iG60gp/SgZT
MwAwZF6nt+jRiqD/WaHzPhrzdQPHzLG7zqiuFJa9t77H7fG7otLXOCGhHMrsReGF
jDIxbtxIpPOSKPtTCQNRIa3avCQjFThGrw3ddQjrALxRhOORCPayIcLnA6x1Ov2B
5r9qeqwUF94irVkCEBnCldL1NzEQC8jRu7dk4dUnoSCEM0bI/X05uMPTlKOlqCJe
l10w8Hb0jnDmYblz8yv80FUtjCrCEZBowkBL2wS5M0ZL5X8NW17e4uzV4MKnzAnZ
wYcCQp2d4yApwRtbHr4FLIWqpYbBU0/a/PLaVjB2k0C+ABaU1xatSBAe0JcxLWJc
pPEGNrYpvSZiRkZc55r3RaeLkP0Iw0crj9c0H4OzHOOXfLeZ04HPLJ/FUy3AdrcR
VlFEjvhDpCXKGLbu4bfH9myukhg6cE4otqfV/BO4Sr3iNZyqQPISvW2oscSSaYWk
DvK9qc7Z9CkH8N09R56Yz5sYiteKaNrCCvnwyQ7mahlxUV3uvsXCt6XFBGtOAU+Z
fGkAV1Ebtkc22nelNiFdEGl5GD4zf5UqzizTK+efvxHAcxfCip0zk9oQUdrY+MFX
qRMNZPS3aCJsS74wvtdUya6YW89jO7EjFcUQJnBVhaQUXdnCmxAjjbxRW5jO4j/q
0w9lZUKGfPcl7ZL9lWQ2Iq0w+W5CACjOdKsJbaEyUuLLlGsFccX0r5PxuMFeZYIB
1IYwTJuPB5x5boR97wLEJX1koakqK7aN0DjPok534wIvcMEe1hB+YKXeiwYvhmmR
TuAMrPc1Jq8foKF4cT9Qtm5xaBjug7imCxRwikTVrQ19In/3ZvIoFNHzW4xI2nVs
0YlcA3oUl8jF8S9+STBXg3cXyldx7U05xVAYxVSDa7oAN6Bk6zPrEp/Niq6GNyy2
Kb0GWjted0LI/zXFv2ZiCzGfxl7Na0g+xPmB6aFqxgSLwfD32cQGmj7Hbilgy8Lt
GiMzBqLKrT364c8fO4yh/5euetHIS0kDcWUkboe23jN2IDe3/FQtHDnl69HmJhPt
cuYrueFHPPOKRlUC1wcwxX8MnlAL+KczCHpbAHemuzO2n5OXGFtGQDkNSpWKwAy1
SRlsm5bRHPqj0jD84vuU0kpR3+0Aa0H76p+soaYVCLv2QtdLuVRVhL3N0VWLJFdw
pir9/QiGNYCeBr6wdBZASN871C+FPA80auPLGD+KPTYx2Nnp+3nARYZu10BmsYaI
o/6JwQ+QWb6IUhX7wPCPbAHtAppRAlD8vWRBNF/Tac+AQVCY57pvV1dGEYY3EqNk
xw2gXB6TJ6kUxiFhLczqzxyIV3Iezxe2y+d5oEIb74Ge20WNu3L7TUntWDVkqaqZ
hs4aWDbku6hmTbtjz9xjjhrTSFvs3SMjqf+owAgLuJTPm2R5tI5evSft0MdyMUgo
KmK0lCxXQMDzr4Y60qZqc2jwByNknXktLkHGcNZBBOMBd4/wdgOxALgfDqdESyET
KTVow94uqajB1Kl6fphRcoz70WepsEA7d1JOZEQBB+3RG1jIHpS/8BwOIeKtP7NQ
AIctP/lEsUUXS+sTWxywKysEUUf2RnEZiUETWStlP3BW93ZR13JcnbJIORzhE0hX
IS5p6zmDQCGr/gvjeHmClAw+7nwyDxEiZnhFXpIStmaPQ3cCGupsIx3tEZcOLXaq
HTGDkvLuSD5/6dEfObjywGThy1a0yc3JZHZHRYrxBmMTYqTbcP5N7xWIRboADXzS
oZ//BBPp8PIzHFD9OEUGBmHi2bB7buiN85n1cZvbCUfyuQ6hS6YlMS7QEwPr/reC
rSYrYppuEr0xsmCxjQKlCHsar8csRw3NFNmGCzU2uRdfVujZZl1VXRwbFePTrNjl
rMSP576Ri9ntpOCRV1ICrlu0TFHpXIWeRnHdkzDAqP+JE77k3Kkha7933rf9n26B
d7h8O8mbXtgNbtUoaMhy6LqQPb64PiU4idHwbbSbfC5Lwv8U0vNpA4pw8Nu9/3BD
Id46PZj0OHs9ZCgCx8aD2TO/5STFXZo5Rqj9OPZZTmJQUfxJzM4m4VVVNdMtCI8r
7OwmK7fX3VciXxPYgvI9/JqQqDGHpp2x5Z60x1LsTQhnDwH1XoMxpCEuhQxbZdRW
e7i4D+lkNrXk7FJFODBPnWCK+l5XZXfjspGipBfH0liLHceHCrMz9skfs9JW0mAG
w4b7NDnc3rEIxLWYR6BErMw+7Y5CGL5/qYxiYuEc5qo0gOm0skOCNba6W1fy+7f4
qzwDjL+M31zhv5SwJ090NFDDH74zkKuwXCBugGcCxTFDs8DB6g5zh//J+IV/1l2B
6FGXHPOk36nTu18aAlg9NbVkkAds/tIBaNq6v4eMH8oTbQlY5aXUUoAtY+7XobJ8
LUa1gdVcSgdeQIJ+geEMECyJoxwygzUboJk3sns1hrKkrbIB/EKW5Dgka2EaqlJ7
KbwWgn6kRyb2Zd+xjYdN9YbBk+ndRQ4zXhimHGkrYII6HTc0eIqlGfBlysakbaEZ
KpRPmwBlZ70P2xkkLXNFDbGiufNjxx/7/Cidpwbjf3UjEBmn1Rrqy4JIygKpFg5U
NVIrBir1dS3xrE584iNQCLQq6Xs9Q87GBBOwWYBy0ceFQyT0cUvYvCrEjm8VS/Pl
rNxCWei3O82rWaeGotjjRwtPLqlK2nmXJZ10eVDLj5b8610ADG/5Uk+xqurOYa+W
LWI8OfZTKN/EDF3FPGYDWPDYAzy1RHGjp7Sl4TEaZ9xKza4ei48jCINB9Zmv6OHn
BFWooUxVgMntlyDzam/iE8K0858H5sWHSBjoOgGB92UXbnl07PWZLgyUjm11+yZQ
rghjztxcJYYxdJZ/WQHhNQehKGtuEOT1NyCzAsUovPtDIH/ShMMH1kjkKDFYJBIe
TE6wnavBrlgJpqQrXqvQ35Rm+sSmWUl74Qt4Amv6J5o/t7xN9P/D6ke7ZPQjaiX6
zH2oHvFYMhUJRyIjtf9C8gc/mv1fTzgWDt2/JAGxxuiThmVQYp+Yi5Rdj4dAf0rR
G1ut1zMYJHPModGxmvZfa9wdgNyNGYRtc/RD/keeSMNqnZjAqIsR2wucsp59nAah
esSx/Z0latnX8aOaA4qHLJ451gkMQk1Q8b0OtuFuIpM1IXS+9FGeDBQf/IOtmzX5
JgGe3EB/pltns0/0WA30GtqJdgr8J7R0EHukoCWVXX2BlIADKEYbEMNv03ub5ijE
brUXZ8MMVogDN3j/n2x1l1vq3f9pOmk75gNPalw79YgL7CjWNbWxx5U3ID8/mT3Y
qkiDW3wp7GaOpU16uoheea5JvPv6FyKo965mk32q2ZKpBP7coXeKj5h8Xo+Uvn6b
CZjyj5HzC5QYFmGC+1iqp0x4laXfbl9azEe5wB9WhSKd/zPv41eP1nNUlamvyJyK
rl2Uq/Stbf7HqLmLurBh16l6D3mqzEJyjaSejc/INDuCz9sS//LlgFeTtBegWuC+
Ur4Kn0gVVUSpQ6QWg7Fss8p7N2+E0YNtSyV5SrM6ZJ3UG40qOk7AqtoC//SxQ1g9
ThMemkkEDogDMuYu2JVPbLoNkSoJIlKPIP1d8ofHgpxlHfx6D1KiRZ+XsUesXBKF
H+AtRgWSBpUsBQJTnDqoILuiXpMokx2/Ph2HbHCv9LKR2yXpxUDAP4X9WDx1BeC2
oS8uiPjTWk5iFPqA7dgaYLhB8aBOjfV8yl2Ys2SORddLwP7jyXzFC6A/Jtpu4AlZ
f4q34XbdIrfnRi2HoFXQ9W7iR4m9mo+3AwWjAST0uDaoDWXORYP25jLrAOu5PVKe
tsNTcbbdrXCbjCN1r9AkVHN73jPM0ixZAUh2mJGxbIp3ewv3PNscujNeCG2MUYvA
WmBYYrfBwY2VlsmeGI8L76qJz67dJujeDGodvFvG16Sk+ZHLpoYC09smNDotWFaH
EZnVA7YBnqRAzEnpUehJA7zCeyaPvnf+zokUJDBKf+TpxTKVWTBua9LRYFj4Feo/
lw+rpgrNrVuqt5CSKBbETkAM2y5ksXqzk0ziFVZCVETuT7pu8Luq3XWzFkOTpElJ
KksTqARD2HBf62fI7h/PD0HubyxRQdaWfRW6ePvSWtBlvcFuj61+sBg7fHjfeVeb
461NeVYvVdUaECZy4bg8NdlWu6YGYv/64H5SlAVcbpmXS2EyfircUoQ6Nff/gPdD
1LLabP1XJDfTTe1+uQKg4/Wf+ilbFymnw5slqNCyS9XnSD6EPH7Rx036Ko4eSFeO
oQIt9Hly1RWnlKyNDuecrxTmHgtmHmbsj3LvyUuGDTBk7bLVD9pqoRQlSSpIYCv/
x0gBmKwr5GYyiaAWmsc6LtK2UPDbXwlf3s1SprmPVBGbkyUNsmgJ/3nlWzXp+yOF
lCs90vNcgfCW2e4xMj3DSB18B7aiv7KeD3gqRnYp1avzoInx0wtpx4ODWKqYGd1G
R4Gzq5J9xUvYOTcO6eVXo/s9U9C3STBeg9lcG6wjMKMF7d/WTASLg31UlmWGloeu
HF3xTFnvzJLnj/J5a/id4N3RFbbCUWRQHmQ0e4tYL03zQtIVRaQV4lWpvImniX2k
oS9WxeMBUVWJTOUonrZTph0mHbtIlIxdRb92OAMJlYoOE3KiR7pGJZcbFGNQ3cur
vtIyWIIjw5VXsPvrHw/FPmHgRmLwem4qxQs/XZlhcLjqvlwfwdOfMEqMXunrz1Xo
Zc1g5cffKW5PUBD+zXCpze0NDiegWZWxVsARX4QqumOjIzuHExvrzqvBZeNMC3+q
ZfjtDbMSq44IIMg2NEpG7eoNs9uq9sGuel5WI3HMk6qEBgXVEeS2fi4v8hErZrWB
QFsRlCDLPPLLjY951SzjN1A+RAkTcpjENipRoEUohqXhAMy30Xy6Xt0Q2Y1EDtRp
YYRnH8U0/CdmMV+vBpiWeNAdPx5iqBcXXYChn0nGQE25c6N+iJgK5ZwhGayCEVin
6X3fIhrsf/X9P+DZ4sohimkyz8WOSJHhEl/d1DOq7HLSQEkedo2DPunMO+0y96kK
K+FyVgrIGqltD5RvAPfa1ESI0SVSw8+g/Xb/4Dht1VUWbTRPlwlHJMEsfOxztgPU
bkOgGOl/SXkyvOjxiRGSTuoXIKleGU3e9nmRc6q9ZyjNTcmAzMwS10t7pvjcJ2WK
+j/8nOI6XsaoPYOXRKqn60Bwo36EsRdfAzSxLyfB0dmU328be2z0jBrUCtRNvZpz
1ky1CZ2Cak6W9/s6bzmK1D89bNDAy8j1QM6TJoVBwAD4dhCg6TotyHkEkOQs7dsq
n7yDyhv16tPrT6EC5c5xZKX2MxlFEsWNwwggyJZzGAiWl9SBUrOSTmYuH8TMNuS3
oDlTcYhw+Wzl7R28dJQXP7ENvGVuLIeTKJLGtC1CfHyRjlurPxBqBCyaP1qAwA2s
3bpUhpFlNbDZVrctQKohJRxpRkAabBNpUluQ8gonxksM4MUb8Qtd3HoJA+DlpFSl
zq+A6jz74nt0IfsUmA6gBCaupVZ3Z47PCbPwHyrj896m6H+zEV4mAjGLyKse9iDK
wvaGKvtUM+kadpw2M/QolHQAm+8Ad/wm6VJnXQ95EcvD9hjeqdCdsx51u1z9rmma
YXywv09B053A3uqi7GfBsOTSQPwjeKz3X3Ublk8ZVq3qmAqdXUE09TdzV7ewkq5n
/hLRUJFZ0vemUrg4PUfC6lANqXDtyQ9PAAeFZJMub++Xng4xO3iAfl3hCYmFsZl0
yXb6PLXuv1GdYdjQSvBejuN5t7dAQu5uFrSqjuIgGL/FkHKnhpBIi7BVfPRnwbHb
Qrma7pq6ObVNNmuXc1P7aE8uBKEsveneU4R3WM6te8erE07Bz8QR67QBY80PzXfi
hX6D1rQYEqo5PXuuiwKECn181OaIphYs4fbGkT1veJVTUlLx5dL5v4VH0IlP58L2
W8++rTKQmmI5ALIb+tgzl8o/YiKs6uJLJ7+Bbawtv19Ui4FtzdbG3OnxwYlfGTAc
Yb3Euxqvb6ILfJH+F8OhFazzLqUwdKxsltsHTuWruGF0p0prvCZR4/2M8hsTMkb6
sN+h/9QfF2KhqrKS0ORd/mrC3Gsq1hOrzcs2wuKQKUTH1+2zmW++Q2I7+MwyKzG2
iDHz7jnhVEkxiIjnMBazrEWZS/H20xfEyV28ea55uk/Ht78M3fTDiXzemfMffq7d
WnGGwmYJtRaD+m8mw0i/iawRSkXfEGG64hGiQWpwYp/0whTUxl0bRVT7xF3r/fRB
KdJNdNYKchWYnc1DtS7D3X+So3P35bYvH9j9C6uWHElhoYYBif3kp+jHasnUPyJv
hjOWvxQ222DfYifzHNAd3syBpLdMANo4LtmXAG4sEUf/5gzv+WyiQCZpB++zF41V
ztVtcC3joLtZiS1nT0mFpToTIAsgDpzJ5kCC2ekmQ8MU0LudH+j7iOSgcjeDIysR
JKoSaOnwjBpSJ8WtFPvbwE1VO3X1gYWViumuqsJVvyc4MOqbobp8kWQEVttQMBCl
PR+FJuM4HfF7zkDC/4W3715MK3Qroo4JDyIYEA/jbwsjMmDxUwyaOjAiIQKUQgIY
OKsmNek/+qdFuMStnVdYrXtyb8NDIV/y6vsPZZApW46gGt1LXNFExR1Fj8TG4a3s
0GcpiZAbYckJSMo6pzR0OQOav9aAYzyljRzzbySupoa4wcraZMCoCn5PxUzEDzLY
6qRUMikVE2O4p56u2iTElmPURPAuj6hRViN82v+p91Xbeb+Daqpkz3kqvnP8N/0S
uR6PRs+/VT8cZGuFznu0cRPtwn6yH3F/Bijz2+w5W/ltGIMs4EpRfeN+wrsThaxi
PrClMDYG10/kYyDD9UWaUfVU704wmPQrYbwHQKHo4yzfbrpJkAopxkeSN/K7TVH/
zdv8LrW6YViZ6dnacvDDrtAREUjiYGybnNb+Kji0sSkRfLRscdgy17bEkfCwUJbs
Sj6kQ365PpI6HanDg+1plyb6TvDEwPdbRU56yL0DRIxLWj8OGFd7eW7WUzWMQR/P
Ntti9LFxfBYJbEhKeouFb1LsOCdt1BtiZxKwScb3hVo1LFdYzz5Vj+qBo7v0glgJ
zYLVXQx5cTKDJ7Z1cNzhAJl62OUtz6rfnHo12MxxCEaEaqlNI+8cX0+PKxgoM9Ct
Tug/EizL6/5SmEfQNXgzCjEILZEX9Tr6qH+qXZ20c2GMX5UAwGb9EsHNjdPASuzO
UP/9UUW5DrQ/w1f+1+dDDCTF+CU2jiWkIwyemkcnmGvmPGRgHYC6OZezxNOrCKfS
Z+5qm6bDlEk9a72gbTA9HcxrsFZMe63O5Tmm/aFwODDM2EO88CgZO2C6BUzND0T5
3A4BKbPQ+jpp4pq4mBNWbANphyq3fYR5GQsXVIQ0UAeaBFaejLqkCjWh3qEaSJ+V
NxUz2ip8qaIzSzOheWulbT+46odP8qIySsqcxGuzLH2NvIeq5asWnVdm/de/jfh0
qmVxVxzQ/41B2TUPFLviNbPXux84jj3Q15UaNxAFDTJgx1TTRknZKyiFVOag+BS/
mbRo0rPBiP2zgm2MTn7r5vw2QheXfLN05uXOXWpUR06wBuNBN8wZboqtqTJRdLHG
CdlEktH12GNeH+zIdTEbSHfklRt5DxTXXRuCLtZbamdqe17Yq2LGM63LMy5fz3Xl
r5sLpfBq/YKBGKNWxxPGhzdRt61GbrrJIX59Go1wv2117+mZICcKMFaSS+Wc7PmT
tgbZJQxHn+YTOKUSeEWgbVxexqoRBOFBgbSLAkS4XxnJmI+eBW49lUlvF8DIjYBw
cm9Z5wreGUlTHHWKw468X91itwjf010YMLoT/k1unfmzt+4RGvD4suHomYBoR0QD
zqk4Z3Zb6BTZO/5If18RZxRd1lmSADrEnL08gA1E3Ee27SacpXh8NJu3cT0GuORc
POfwvAQKHZo11xHp7hYoIQWRLU+aKwuvsElkvuA50OtjnpPxOL4DR2o1buK3q6ak
ic2CtbzSvNXbGGJpfY1b8ScwHkgGDeW/MoDp/YbPPlQbU2m6G8+2aVAyEPS/xZii
q1WgYesSck6At+8o6cui3fU6WYfyePz5KiOpqiSyHB/bPAFaVKSl3IoO2JlCFhN0
kj02XU9RPwQiKFStyDQV2lXVyJSF3sC79rrd4Deff/UKUUmMd3D9mISCqBVTud/E
DupTSJcT0Ct9WA6H2DmXLRXAvi1qfIZMsvBN/8pjgcrugq0NDO6jHyjS5OtSDbRz
Uq+gwUYC36wZQ/P2X21FN4rh+76ot2cPwLUzkJOuE5ZfMYyQ3FBp0WGmiFcnfMkE
QfWUOqqaXDiRUpj+s/+HnIHbK5LLcwAkMCPXWXdwcLMw+6oZj7lllwHEiMeucsFt
RHZlke0OjP+DoV/cr30DBDPLfO9K+9czuzObls5O5m4/3pe/vMgr1wUgUVseeNpO
sSOh99WB6OXmjipqZdvGJ1gkXMHf2NXHQlQ3uj+AZE1BVvBZDqjHLDAPM2PSZT+1
D9qzIitgcXFnpoXNwKyst+FcQM7+j2IR3T66+xuVzYp1dUj4Y2QVvamTwDVKWD5M
DtbLklEZo/iWAIpvmbsBLfq3RXgEySAHhQMDWaiuU0+enBuRQ/VrdK9ybWf4/fcC
Od4uObngRyafXjQzIozLMqft4D19Yq1iu1RIrcQOw/9Gn6Rbd8NKJODY9V9oeb9t
k7EkjSLF3WEC5779dVtYrR1lCCc+ab+XlIUy3Dg1qBUyGK1B2tC/mIHszKqy7FYn
p/PydOHRRtyBcpvdC03saUAOVj4Vyh0gg3B9C+vSvK8UR/MgAS157abPm8FZbPPT
TM527dpAZGyTAt7GBFSt2SUofxCDzaHcHNC25EwSSq7gcV699BgG3I92Q3+wdT+Q
6ea9cyo8wuVrI7f2GX7zT0TOZr6hOC8jj3H9DyFdarV4aQNqnkdKzlHnXDhSojX/
eqSoNM9pC45tjZcxtEy/2Z6ldHzwUcRnHzPCdqEj0Y58SajxtwDNg2C4OyZml51X
pG8jI0vi9qKhec1oY1smerAe7yUGTeKP0x3+fiUhbWVx6owuvaxkwaEAvnwETHBH
RjE5ZNYUEPUntcT7e8AmS0tGa9ybgBrNwveYzbT3yWgC0fVEoKRu3Mub67gNubuE
3JnZndqhBGpd6Q5NC3k1mNcKtZPRu18Ayij+XcgsuWHvmTsvjp4eRuOSbDglU7CH
CHUDdaQzIvoWrzuNndvpDzLqlsrbOGrq+WZxghxZ1ffcIbf2AZaCz7ST9rYhHucO
CKJjHq0ZGkoG3oXO4LjCd+k1B5gyw+o3BBcYx2uV9ea1N2w4w7ieVt5m3SDcE95J
1Hyoa4H7rFNZtlnpZDy2ULul0uwd9M/iPibI6rWPOlFFb+VE/9ts0LhX5oY8BOS/
Me29zeNasSe53qE/FDoGhlaqGsq+Hqur1yMZlgQskcHhskNNvkfEiH06PfwjOXlV
yiMsvL3iGNuriMnxnlezNQOQSCnNKp587ZN1gG8XTMgWxRddHeTGgVujCD3Op4fw
Af/6J+VJEjwa9ILsAzm8AgIPXE9hdRCcCU2X7oYTj1/M/z8svfXb9T/lfPAJuRUW
9WNtpOmeh+RA8+Gfmk6Hq4I0zg9+oNhSuj1U/CeXKqG1gpN2nHlv63ex9/e3XG3j
2BSEzwgN65kbHEyFTYK6EPLJYdKcTgSJAzuqQIKDHpnA81y1QhWs5H/14k4n2MXp
aZCmS+qats8yKGaYBd1vamLfI1/XmwecMp0d0DeQagChleiUCcBW2SJQKuyM/WKs
+tNRMk3Hp48YTm5deBo7z8y37O17dWhliAMfSJIbFZDzMuftHFANBJRm5+ZkuqzI
xhf5oAZnzlhNeEwNlGdW6SDvsqt9SNSHFRBo5S/XgzWoYMsgtuUCb1gEGLN8vMjF
rrgxpHij3Nk97n3dG8UWc9+EkLigv4SKyD4aB1jCRS3Ec0IM0yQdvY2gkJvN8+Kx
oD+L0b0S8QroFczdbgld9xaGBb44z/G3xSimgHEhV6ro4J+AC7ifyNsLopRbYlOf
DicSkHOjt/g++vl2ErMzdRGHU1rArIMv2a6XxAUoPjSOzDYXFC/pR60Sg3M1R5wr
lpRYoMPGnSUHgIJsM1wsGivFSSz3RZlbdLM3eDOfJa0k9bLXDlimnGJKvwwY/bvF
gHQtpaigVBgKOzq7aEvWUASThVTkNV3L4jLixkITJ4xtmiciYbTXrEsYoyN53GLx
tf8FUlPDFP3MAZcRvfVV+3vPnFvCokaRDB/cKc8lZDweljmZbfOvFwbrAPbSW78S
Z8TGZpa9IkUH1HoF7rnLXUM+7w+au4kefFVGlfGw+SAaRlXjGOEF/VCgNzGJciij
GBeCuHebARd3OkK20zkX180C/u8pPppwXBgxqAbaGnxTzdn0jCS68MDRrbE0Apb0
DeBODUiDzMQKq+m03h2ORImEwNU8v0LfmMmyE7lolz99BAnMVo9HRtN6RSN5Ga01
HQ/c+nAq+R9/nUT+ZmEGIM8VSlphcOXk+Iqqw2JqqClhhF5GyCvw1txLnzLTPstS
neYPtJnospazYH56lqovvyUelGmHr3cGsiI8rUWPnkvVeDIA+PV2NGPhmbie43dg
NpQCg8eGAra/F1TmJOO17zASu81TIXLGUbUwGWbt1V0hPWcV1lF7AIq5owCPPQOK
72fj8We4x567buEyukRF/Ck0U139QKmPPOMOEfBHEuzMc7pKXoBUNVwjka67zNWn
uaBQk3y2V0b6LLvfO6pwWmcI3pKbDx76mCKE1snjfNfW5yveKSwoyutbwHm6On+m
24TyTlBoHIGKE+RkoqCdN/eCujH/StXt2HpQ7K97idFuJXnufcfwQdUWH0zDqcAU
h0sAZs6pK8A0trjpVe/ALwWO42kJR4ywQcYwXdv0AQisjrL1XOW4416tAYdr+lgE
27J0OYsocozHEjX+Aj2oVgvzWIlpy0rTrGEKBtRwrDoYoBJo/++sRhn1gam/shmh
voN5rwJM7OtsUg/50RQYgLyH2xhjOHBQP2wK1BstWMn2cduQCPHppSYFMEdULxnp
oHxNYhL1n/KQuSA390z3EDLshOPBsEb+KgCdMVTypldZk1lF1igjwI6ZCTe2y7/q
ob4ZMuZDnh4ziflE0EGstEy8LQ3PA9rLZ386dOLXlGnGTg4Y1lTqVieDEV0Shwkq
PAPWQQWMkXIE+PDlHfUxOGc9z21cHz+dZs9KWqxMo5L/pR2B2P7uEqxgabnpVnJm
R+Kjut6wnpcrnUyu/z0aSa6TWZROElzadwJtxznhqgkEhOHWhLac/TGaX0OPWsgp
T6aWTA2FQ892uHzJdxAyAt89cXdmOjuud+l/9nGgmnrfxYFkp2ndWoj7NhWWrWO9
EWy/8J/nMOOWebKDT+XDDeNW0cwt7jkhSqXy9Dn2jo0l2WCLakYrsVvz5RUrH4Bt
hoabUmaLiGPiQsyf+IRxuPk68jYP/cIpR76Jvim2/2CGbl7EmLoBp7HIk5KQCvNQ
ikRlKXxZXzLoA8jLM2ZgIFFZJeRDlsGAvJAwmRFTYJrnmcGzefArjJO9wFuY4dQo
fnWREX0jQyZyz4LNE8NYe7HrBm8302Qgb9K9ExSdrzhtgHpwWlNMU5cg61SNNt7q
1lm11NBKTxB+MhDRE9oaJiJULQaOk1Ev92ubeSE2MA5CkPDlVRVHlaZmv4DE85Uc
qUOQZlMk+7cXVMZlLk0fQRfd3xwlNTlXMSIarhjR2YY4PGi6d3D5bUMmlYKAQHdR
3EGaDt85FxfkjNmOBM5ZshZ3QWtsGzwd6ireZgeGhBocnMgj5XA4Grwf5+yFIPxY
Ftw3KqJk1gfi7KtzOnGVi7h2Rbmi/GGTb6owdevB+Px59dYHkB+1cAXQiDFgeh4W
nAyhHbxaN53Q0QHPO8+KpdkVd1W7KW6KeaXwGKqv9rxd3kzCRZqK5zgJc42iucHE
jXa+0IcOsWd09b/QBDiAkDNuSixn3UlcVHe85SC6IvMgZpHo95agdzUu6SRk7U/e
yZxuM0jHMgPwbLGUz4e0vlMGlYiouEbOYZ2K2qBBwuC9OVZz8pYio9QN/ED4RlSh
G6Rie+mATAepVYqx5kWGPU8DBI7BHR4TNSNXqbmTmRwBid+ZZSX7kzyqE3YttDyz
qXAdusZkgwsXZWFWZFLoxSSX3H8SqDeRINpnB2NuurPbp6sLxdFH936KXC16qapG
ObhptdfPpwB7hXjJZ5NsaOfGBYd4CCFtvG7I0bfo27t5S1xarW9r7SukAn/kKL+e
LrBNh6YEi5jL2J+DNd1a1FA77mUl/0SuhiKYh/79qvqXh1n6rtBXtqQfJkIO+kU3
rJEHHqaxiN6p/YMHFt4iJ/yM7LInLdScMnxu1bp6yitOujhFxTRgQ9ENlbG8DFuK
uaOSKX92QVrVUQCqFKfPTcbezj5KIio4R2qWVTmMpt1JTh1HhOZiFnChy5kbSR4v
E54RnU9t1SHfHliIYT8FyN8mYqp+JG/bzER184E3iK9LBMK1Flzj9VWW/TAVMZPi
5PlWTikqzWrAtsnwfWf8uDpRQyk+Y3phkNHWPXzHLhVO0f2JJvkJLzw7ec3Xxa5x
r6/wnEH+mFFLBpHa6qG4scAlfU+U0q3Ix49+xRJQF/q1kJz3twTl1onHsM8KvI5p
nvl7x86zOnVDPDCRTEk0bfg1fZMy4maJi7BOwxcQ/+V1EBHtOIiksCNCt+nS4cjm
Vw4t5Y0z9T/RSWmt6BuAGOf/XSOt7S4cZaIJdpvdPizZf8A2mWFcMkPXlnTf5Uo1
OojqYB1aUFZ/zYEqKanufRi11Mu39KwXmCFIOKNcAapFHPqMAhmy53h4M6DVNJd7
hcQNqz46hckqKWxRg8buNIhUTvx3hZEO8fjWNqqNRaNC5fFvpkkZBVR0hnbtoH53
Jng1VQj0OwU5YkQtw7x44nrTf4NuyLdBalMCRVlEFSxrEHKPuVcnpth64/KwUS8K
Dfk0sg5hnNVz6tIrrKg4Ep6yOzWDViD48LCV0VslLXWIwCjAQ33K56BRXPZsyCj1
EpwWVaiwWIeVU/I2InXjDj8mSeL6Rq3Z+dx+Az7mjjaoAoEmPaGH8KGwIkKjv2rU
rFr98/0hPFqNfNm/WSbkLPz4nMPlCopL6SGtUYhmX6FTv+Tq7aeAtYE8llLSMBAM
/H/nhhljYptooCx95O/42/lUXWBWvbDPVFQKi9jHXPr0nMab1IAKWtjsValeTp0/
CQmE9ZQkABWVgeIuZ/run2jng+r3R9gZhBAscJUjHjDx5bUFheKv/LhqdzGtjluY
Nn1Hq/9BniFUU+DhCGcgILuEJQtzcVJEum4G4Q9vGje43fLLA2EMe3F3uof0DoVh
Ag0ca2Qqv1/uNKUpMsYtlRHwLNeyM/vZZxzXPCQTGwQ4sPl1p9OJKstP+lX57RG3
Zgide44ELprXLK2dz2olRpR3yE3weiIIEapb0GhUOLvZ2IF7mWyDiZWvQB37CLDU
1YE0XbpQNVC0MzJtuB7Fj1AhVMd3Ki8wntBHrC4XzUuLn+Hlo+9jxytTgox9zEK8
ddy5BbvahHj2FmW1aOspKIlACHpZ1xiWtiqT/kI8+pTv7mW6lUyfaM4L+fsVUOsT
ljL2ElpA7ME6uv7dCU16Vyuwbpj+AHDTGA6Xq/oOUgLppy/q0O2hhJszWafDMvlz
Y5ARvtgthuVWm3jsfgYXWwUozzRTK8BJLRHQcERjF+VncwFJTklfsF7YKuKBjOfV
bD+QcpPkbjMwQBXYLQETWJiuchH/sA5cC2l9dX/4LWmUggktU4LW0j8A+H24hmDi
T93AR5F9knKwPb6pv3w1dvJUMK+kbM1+I30DelgEPf4XeEnKSJ5sMz2jNhqCChJ+
XVWNbb11lyxsdpzwCTUJMmU/rgJLBKzvNATGxQlKhLisPshcMgvj9TzR73Z5uEJA
fLhbT5E5VrfmnNVam4o4KvtjAzq5p+ERsdFMw+YDiL2CzSQnaE+BPSjfS4YFkdyq
eSsC7edREumfapxLoe9DwxrKISp5piXtWoQemNpPmQUogMLSrkZ6RiFY/ccEUIEa
90fBjCJ4OzW6lsUEyXlSUCIvvZUTe1LwAapGhyJHUEylbDuwcE+1o2ml7CUmToya
dqUx59HLZLm4EYpkRVseNPIAqUYfVwqKlo+KLeZdbor3OeY0aEnN8KoajDeerA+Q
bocrjPHQ83obtyJgBnE+wxSCh4VPT6Ykn2cDTbMqLZ3J85nbADkxfaaZgs+VpF0R
qddNjc8w1nrvRz936tVXY1UVFt6vW6s0oiD0SGNPjgp/IhQ4QklWsJzz4inbw6Eo
HFxJxSamEGhJXhtb0bWQFd2ikiUCaGHCxYWHTYPUnH2GxiVSdBsUJxk7YyptKJ/X
0YF47848g/UQGe/RPmCRZOc4BT2/d2/ddkEuUwcNZdG5+6ep00vZbJPY9p63Nqq0
axQTePfjQnros/rouwm81ohDa2kRjjIG9N85EQlSNfT11HJyqY5lg6XG9gnzpbrB
1iWRoYxdt2rdy9EJf2UnLDOtV/or8U6/qzS3V/AdrUUTOuL2z9hmPGXkWbP9iW4B
KywgmoWiacSkmauafQjgnxlNATVrRbvM/1jQz7he6+i4+8PjWBemp5YlAkJgWowV
uukByEfrLZJBPfi1UiHDLXiwGKWvz0e/VQKGbn/zggqcjxRWb1VhQ8UvCWPaj/uu
oWRipGWjgUWw4aUTiDidjnB1PX3oZ4UdU5TmHLppNkKuHVfoX67ToLAZ1rrsOrjh
fB8OZ/juZQ3XulAR4pY7cPco0n7qK9D0y8QHYnFkfiuyMxZSW1Pn82E7GuLb3FrO
D4VV/hnPmOWZ6UMfY593mb4Y2KBmHVAh46YErhdrZzRaoPVnyi8p8Loh4n/ZZk+R
j4sYFmR8iN3kBv4BH12El8Y26fa4vp94GOtBS//jwiDFebc3FkYDNikhBE4myXF3
Ipc7aZE8OmijdiB00iueAFB9fB1P/gln4tlKI7HkeRUY6aiq8ZZTNTqwy48ofz8R
7quPEa6SbOihWj/c83asg7zOi99b+sOA3DHT+Z0NIhPqnrKZ30sSuZhJGHkBgac0
pzc7iAHhampcyFsRifBEHzo3C5F2LmF5Md5714lSwDIVtPJkVKnE1ormx6O6vw+D
l8+o+VBAacX3CLQGauNfnFvPcGFtUIahjXbCD3LuML55M36ogt6DxGo9pIs/naY+
GX7XMn75cqd9EUNcUDxRUW38bPOkW2mcJW/HZU8N9l1YM2y7UkTw/WVNO3vWk7wm
79NgXBTGJe/z6O+e2GqFmOTIfOIQMh1RUTm5tOEhmJXGrWaJdEYjnoYCWb8PTOY2
XA9o6JbLdJR4LddamkBki8m3p5pFTNCrywrHDa+Fc/9PMRyD1GT8iN7eIJBbIKp2
tAqkgPgxaK/OTjsyrsSr8N8UozOHpAwe7arCR0OqLb7h2wcU70e9I/ItYsYfevXW
f5S7/bSR2j+Pv0uxh69BqIH85qec8tAGHE4RT50LHOK+9qguk+D7FlebeCpYfC0g
scmnYri6o6s573MfiI0rpJYITLep0pjaKIJK11GMNmpZgAmroQ7CX6RXzRnthwWL
SSxUhx5zGLGziNa8GAZRSqveJL6lNAqFComRv5vc9NIhxHUd+kWgpJzfkaBrzcaS
nmXTh88UNAFBE37ip49/zOWzNJFIbmJhoAZ+u2GFfUMuw5ri6uhGmSErj6LU7W2V
FYkc70TvII12g1N09s1WoSUCjATSnWpKL4db2y5nLXuBEYZLaAC2SMX1jVVGPr2X
ZItjC+nkZ1FtroLvT3ocIyvhMl/6r/7V8rJFp2AJlVRw8gHs1dk1gVMgEKS8Q6Q4
LBHgtZxJtL6dfXrBs8z6si0cRplOYO+hjmhQyZeFnLvrdcYQ8ousXjbm5UUXmjMz
wWjR8iK79JsprzMxFWTGRDV1zVr0dnrY2ijHEhR0/30AETOCsZdluSHIMY5gGEv7
ut4Tz5K9V8o2p6IhO2gVwTQIldQOFGYs9sP9A3wmSclXza2FqzEmgxTqLW80/DQN
GIFd1w5vyP0HF0eDoqxjZgF1KLwjAkBjsNJW4W8s3cTxjuIh7JrEXN8I4g9Qt5+U
3OB8jupdIUTI05xQt7bONj16QQnc9VH7LGCIfOP2q8hYi5kK+B6dKjCPKKuBHHlM
kZzX5qWbvEM8sAaYFkxL/jGnBP/coZWjDniW6xUQNn4UYM9j+FEPfE9BqHRWJYdS
CxuX59sxUFRK5ABaMLeqY7uqsxZUPTguXOf7zOZlLslVnUk/sgqi76OfuA5KjieB
tME1b19Lo72wPJM095UZMqFEJinNOqQlRYl7V8nZApY489d1Ku10VR6y2ulY4Hdj
yANzKChK5qFXrL1eOHC7pS4AHllAQ2qgXqa5szYyDaqBhVGHZi3ho4M+Af3MylsP
F7OBr5NT0S0HTfIkmL+DRVVJjYsbfc/jZuzOqVJSHot4jz/QN0nc8MyNBOTaPu6Z
BxvbazrUvV+PpdOaRKbcRm2BRN5pX5Oyn8XyT4z2Znf+6ZhIxf/GbtcK4WiYNEJZ
hKBwC67bs1Zem9r2sUYgHjf/2hEoXsEBcAUVCiG3v2ZB5pQJ18jFWlP2LFuRClg1
IvaltVNCMbHqHcIOPEgPrQsCM4F+MJ0I7v7WhJ9WYwZ+3UvUupWTne7fu9iaLKwy
RURxKJT08fCd5UWYhkuFMJbwbW7Qg8uwLgDFAjIcSXPdCBpB0Z7GWt/74Q6bQRfL
JnnZWL+70/KiJiX+ALK/yna59mbxT+vDQ4lJ4rjImnm4YyTpl4Y9OD1+6z2HizWI
DrVnB8GswDYIaQVKjAdQk1XrYZxC3aRW8qDBwynrq6DMjSkup9NEztiLxFSt5lJQ
QEzW0zsZpm1HaNkCLMWwJp/bXQNCwiBmAP2zH5x25UU5+243xNdH8J6f9wzd6Wjs
gqRtSNUSGBMJ33VguiGCllJwVWKqByagSUljSngDGBmCqzzj4tmhza6gwgqGUU1n
1/1UyQ1RW43Rpt5jCGj5RzCs+3gVWNDIcNmxiPu4AbV94WaF7Bmr2ZN/7UU7RH/0
/skA+NWS15pt/wOiYe2ZjfAIpb/LNjumnvEZ9FJhTozv9y64m5Y0uoeWEbqRHDIq
BBIOrNgKat6JVshg+RNaVFVRGoZB4iDWa4bFO4rhiZA9etSLCkmmQbr5gQ3F3H4T
EPLU2UkEm9A3p4SEsNeAcJvpGjqYM+yfb7TFqBMQlZNyZK9eYq/Ezdvbafz/IptP
4IL5E25LOAgp3CeYbemOZRv3k8MH+zUYCim+1nLueTSnDzUNmi36Lg0liAyQx/a5
AzxD1WiFEDwm9dc64vVzZ5D6+RNNITuxJBGcFBurZ/K2oML60+IXQK2Huk85O9f1
8bxrD7lyYCeaBravaB86D3gyKl7EYo6aoxJJilh+Y0UXA8fc1s62c+HEOxwnhNWr
28ScCYg0Jt63Ov4KQLVAB1fAewdqAmMwlKQwcJkBN1jqhp10d73alvhaUCNKaYNC
CaXcS1ezmy2aHwbNjz7v9wz4GXm4cE4wlieFdaqY3mJWQWQmOlaEuW5BwiouoSz+
DSdo6EzkKLlhSDaKE32nIbjf0S9s7Ij2yrM5qWKyvFxW1EWwV8JoosigPWzPpam2
w7cf3j8Nr0m7OXMHfuSPIo0pJ2eh6/AajJGwSkukxIP9fzp68zmBWjjupDO/o6b8
whd+gTAMOoVBHiLQ+hgkk/d4/J3q+gE16YXbIJrdM+yTkd4tbZ/EbDu0HyKOadj/
CFHUz+Ub4bQPFwNmgBt4hmLO+dgDdZu1jOs6Lna4wtk/kjiSZZfPF6ZDh4Tc4JL7
zaVbe/mmcmZNZ44rl3X9m69DCqdWbTvzK46IN7zUAyFbViZN0Dl7H1nMP+E7J5Fv
ZurD4LNTXFlAzyPl1Tw7v/1ss2Bs7Q7IZcDvLWGUPCtoshZB8hXQXxxKqdbqZI6k
vx/oDUs0OXOtoJaWpsvrIJShumnVVwHPJLFSDSkml7hXv2guapbIjRKePOVGBnzR
2SLuKF3Qe7cX+YmzcDdRBXwgs+0R9nh3uVtseErV1sRqQbTRwDv6GGn4xmeP6COV
pmt2f1riWfdt8fubMRnk3Oq3/lieo8Q+GiRjlhurhZRVLcsweN2frPsZBGm6P0aj
7bNNjWxan7CLj4uDDbiIOFoLrdt4OzRbBOhZb7jBTvP/f9T4N85Y2vrnoWP2BCqG
7laiYKD0cUTLD32LPcPtdqKjWyD7papl3LHpskh9aH8omd22ODgJaERP9VA333e2
CQQRBjuJBCLGrElYtS05amkJ4A2fqdBqVpXOIVgfIwyRJsk8HkbzAsk70f3SP2TZ
N7PqLnpfZlfHHYY4qPrfTStc9mQ69Z4ovBWeD/FwDon1l3HJoubSvdg4Tp+YDNam
EcH3WWDSaF2eeuXQ/A5bqfBUGY6G5BZ3KvQO46ArXF5wnq6GANGz8QYN6R284i62
QNn5nPyQNPmz0pJ5YU3EetgWY/YoNTqL8Wv7RhhbB7goLQfMUP322DG4qTRUTrYI
oeTBbiUP5talG8XOU4Mu/uWE8yo6aLehVa8OjOupPfqotGCb1KpjrYCYGhu2LHQm
K0bioagoQAAw0Om2nnYnl2aEqr5Jo/jlBmXlKkgDxDgBZNlph7iQiyaxmrah5RsE
seu5+/8G7tnryBNFcqVJkmpvwDs1dAZyIsFNthsZGiU/6Kb3ry28kUuoN4XrmFGl
O7scOtLOF9z2a7LM2hAnrHwwzcXmnYIud3BlZ5zAughJLutHquklPrlNckjlYQWr
3olL6c0u0hgk9S5BLODePBsKYi5y9Jw/JHbad58rWH2jXxVulyAwTS2iKe9mCsuX
CfronNrCGRIzZvqRH0g9YhlGSW68EpqSiw4jC5D/ndqrJWg0u1W/k5mVEVtDDdBR
L1814ldnDp2hmuuugGYalKWFo3Yq4G60SuDI+DNbZbXeuIY6hW9wIgzE7g+aoUAE
ZmX/8JE3iNH7lSvalg5x1l+bVL7MR3Mf8JufcTjetk3JVoITYw6Vb7p4M85IXrel
+n7HKIy0g2jvW/xY5plmK9nu2tisu7LxDvqe2MmYB1NWULGlyw3xUCxL4O5Isw7E
fQCPNCXXrsx/4K4L5cte1Y6wT3y5mPR2rolOPMMWplepSKujrlcEWREUR40BycV1
H3iCIxq4Yj+VFLjjpnm1Nr7OtEhL3wWEVSI4pXobKAiFve9JJUHCEMmo2bwgDFU4
oCFjSqphpOv9TCGJBW4Nr8Ppi1sopIFhT9ZxM+4XemLw13KoCuGO8CZZgnzDS5+G
BR+prSR63uwzMjif+AzR7GmuiyAepXe0xqvn+XFD4fTFw7J0XeBlXmTdlr3Wil8Y
Ogg8BOThOICpDO2o9O0ZVOP5V6v0v2k9Z+w1+S0xPnOjAr5jMkLg+pQQKj2IjBfu
AItBtQpdTVPvHwU4zVMOIHxwSbd8UWl8vrEo0H9eZl6phQfI9TGXYmyZKVn12+Fe
rwrmrqS2hXR1NXw1vWIVOt2rRm3L+FrergZAklx43rwNzsBQC8/8B8Ktj/o1tnyQ
8YaSqA9a0nvEWoCuav9P7Mi9Bn/b2zEh3H6RxpheKhT7o8hY5k9XqKoeO4Y7gLV6
dnvt7o8u/gLqA775ugCztZ4hF0Hh0hgaCTK/I/ryye6zZPDpr/0/fO5JT1A+liMA
PXiwmprLTFWuQfjf+iiBOcb4bzniVonHgUwO3SqLHKkvn+0tGCZwPhmc/q5/JF9Z
CjTA13qUE8vIqgGx/6+v1ZZWpKbxATiB909gwJdJzHy7dXb/YlrH2nfH8X78MavF
oUBu7lPq13ncCzemxT+0R60LWPYoZKqhO7nDtAEaLonB7zQXG1tpLhPdQrmqlG4L
9t2G5p4WgnPcCuEff9NOT/DgpG9SfX2FMZqySUgi2JFpokMlPeuBZvzmASO1Ptbf
fxj8Icykjv8qn0zpCdJmZnsTx0rD2gL5F2hKar0xq0SEXES1YAmm9aYHenTmu8Oc
snrjbTdfjLkTwgQZCEzofVxKIS+p1SLcIRQzm/gXzO74JgVo44jZjK59EdSsfcLM
uvSOlNjHxTysNhRSEiVB2kdhgtrWtTlhodo3y2wsVC0rtTrJ2iPKTLDOW9L3pP1G
TCYykembI1MFo+HlgHJGrDGc0QZqf94oESTa22EfAIvyGjbb1KI9Af+p+DPgrTxi
sPICi2SShUGwXHjM4Y+lciFoF9PjEbbkpXtE8NztSuebFnBWy8zt5V9fOpbpo+7d
OzcYCgWasRTI47oQF+x/CpSTsMRJ7QDbVnXUHIItiVUiDd4Z33HFNH+54pI0rFNE
64cTVlagj7xyXrp5MlPLt/UEZjR0+15o3gwuNVtT3IBTUHInCurm4XWS+WdosHXv
uKe1MFrhXN3xiZEKBzujQ6HmailJJsQ90/AKiWeZ0Zcen8vpoa8Jfn2SZnKoEIHC
yUjFWNaCl/doK+7A8NKiBPdP+dvQFnJvO5q2/XMd4NZMziH+elrq++vysyh8u6K4
XLCGroHRla7pHX0V7URHQBSghYncjn35lQUpcCTMtx3jxgaf+NkmbrkwgZcnvKTB
vNrQdA3z+qVV9CQ2Vc74ng2bga0QC1uVAVUeQ46YhroRAZGWWAGJ05wpMqAKrleW
9CCGaDR//vv7VM5bFD9KZHzLTJJAUsGQAapZCwtl2ZXpmQvofdHIoXABomVTdlUQ
R3FY8UPMVf0IiP/5EtO4tNxR+KuL5Sj7Mn3hh3OO3NgtAPx0xCFdC4I/0jmjOD3S
HnowK1ewh3zpkA7FTRZ9YaXhpY+xCYM0esSAuR9wHEctMvzpDABfM3OEbwcH5i/k
DkEzexHJEVe0032w+vYEezuIBA1gGQG6pEmoBcXkwvqXxhwmim5byD3xi3ssGj8W
sAXSoaftVBbkdRM1KoB07cz6f0vuU3SmVUuJUaGPQFaaP637HgwNGUk3vVc50fuf
I8/qw3iw3OD/E2E2AdGtqYgYTqJO7gabkTmwc+F9DL00kkPAcheI1v/QSUni82C3
/P7rnK2yeyeb9HBiX343kKeX9rydx+mbvm6SlRl3cXkpmr5AqCgs4hDAZ3QuCOqA
A5QwIoUEH8pmb3hlJNaaIDpA+vOGqJLLjcUT4GRCj2hMpaig6jeBT5CcpPC+IOUQ
T9P7toKaA5fFt9hu+k6NUJ/wyjnxy+cENRTTuKWwWkyAfG9kyyK4IG/xhCHwTvjR
KHNUYaMW6lHwLEbv2+ivly85Jm2/9O9YDWulhgOJROAO+328nP1ekw5CzvYun7ak
FU+GgfRI6H5smNjpweUtI9OgCXfFs5RhZoLRMtTggKlm5jtBMEms3tWngyIw9HLw
0cdnIM8C+8xTqCo5rTfrTH3/4PPe3IVdol83tlEAW1WlSEIo62HhGwfw0eLoLNHz
WveTxlzvnW+W7lhRKKB8OPHkXTULRve6JrX0s4VjDzRhA20OH1kXPS/4NL7xakCH
K2ewIodjbrLlZOT5L1lUXFtNTgEfEveck3aN3heYi96xf9Jve0UqijwNaT8i0Ses
RpVIk9jIie8BzgoDZukboRESs++0GAkDLZ0+LFGrBTU2qH/MGGSwE7b3Yke4ahyX
uh8oWmggPVBogDn6I8+0RA9VvCiKhbST3aaxaixwV2nnlj/IoLhjBghZHdOSdcVC
Chm7qD/OvC4shsuByH9kRRw2XIBPe9lKbTnPiOAeU+quJknZ9J1jHJCz5NEguM7O
n7taFRM25R76lXy6DVYzqBOj2FCHQHhr7gQI4BO1bpWXx08/fFG+M0ckfrUJTkMC
lTI5HhdvgWxpHfNLw0TwwcbVrh8tAC3ZTyF1a4H0gO4sTGkKlcPS9cVnpMizGTsG
04SsssIOucQacbBQWuets4WuSo7iqEu7F9Y3bWmIuS7w+1fOloaq4GeCu9LNs+6c
6Ofs3bzGqleLbQeWWd1ELgvsCxalmmhEPpo6A/7xYOvD7FgpNgDqJgvHX4920uSn
C9pHkTetaefdim0iqfYIzzVg/I65FvjcD9MXb/hAK2cPppzNf45bySyDvp4vhfOX
FU5hmkonZP2gb45rj06/GBiwH/cF1QASQ9Amc4czNQFsHEWwVrf4joON1fByvfJB
tmCucdaVJZEMy0dW/BBRZuey67iGcSUsmu/eEzZu/a5/u53nm+HiCYoG261RyD83
YI/RoJ1O8JC6pOY1BY/fiZaWOgDWWSaRbpTyFvvOpkfMwVhaZuvmKRTu0TRrlzqH
ox4GbWIq5MHU8XNbKvNTv5q6PRnKf872hMJfr4fBdEwoEAoLFX448at1398vgfUL
UfDy65KA2/XjQIB3nPGU6TOrBSnTaWmLnVaIW9WJLyrgnXG2iOENuF6LhxIbzsYY
IQbQNjevz2nPVwad/hM+Ig1dCaftsS2wEVTmY+uF6f5Cpby+IZvCzUMWe71DcIHE
RVS2hzNZLU1NtfrUqfXHPk40mjeudENHBIkFImXJHiSdpyyUlKP02ej6ZwjILPFX
JDgGBnvMk/MH+j0R31JJX8ZCOx9foNVwc2fmp5OzzAXeM0JQfvbbOKNOZq6+Eshj
HnWmZg5EWre15dQhnh1xiiy/emxSMWpTPxS24drjl1Y18arkALmF4NAPlrh/IN6H
W4tfnGlutWv/D8nQiW/JShHxja8aXja6OhzQ9Z6cayCDx9hqANI2OS/vWyPrlPi3
q7581xBRCfyTctZVMxBv80emCJoLwbW+rMerH/92G0qhMFf1UILJQRMeqAENC6aI
bPFttxFtG/t+pW7yDxbevKETidsbq7Pb9UYFUI56z44ZN521yq0baydOciAlE/lB
+vvIkP8O2J0OSwgPcDiZULWzeOaW4RJxsGjZkRtmIOJCt5KaEELHIp0+Wsxs9ELe
9RT0Ri16RlK3J2IknQySbkgSPZorXDH0XRf7ijk1NUitRAFTG4cKVTHq899U72kT
5DbmslJy6dc8HJDP4kMq9Ulq4IK2IcKRM7nnJsOH/DND1W0NypR/ZEYonhHTIVpJ
9sjxHdepKwaV/rqWDz1v23n9K+ijplS4JEhL2xb9CxIRtuYQOd0Obaf3sCBEbDIv
clObk4vK3hOtszlxSJPiHzdYhrFbWNOrSAitQQXvCZ1cITxAnD3Qco/7mwGM0G/h
Zuttio6TMvP/woKITDF5sIEoGwyS+CKDs+47bCdz6M3xPabDOWIsYAIZYnwWZllY
wG28wbsrUeVc7086blbb5WDiRIK/rgcwW1emEwoWOYd1ojYO5O6nUyHA2eYdvHRP
EaJmFTTa6lPMWFytQS4Sw7v3qWLGFHj8LxG+JVRRPIltDbrR4tu/5Bz8lTUKr7sw
y4V6f+MEQe0FW0rF9QlyhgnTytpWK626FFXkNfEXmQXZVwHfUInDWhCgf92kJmOY
sYDb2CZeeJMmXz8zU072p6FqzrNRTJYMNhqL4hlb2xdM+lk2zUJ2OX9EY311nd5K
Te9YxvIZLjc+LMkDjC4n81adoEwQtNfViu4zV3NnJGgUUfUqBTWQnw7EAOprRupa
eaJW+sjg0iGcxUiNb+yjZBRdt+EtvOtp5x3HpS/V3mH+3Mi8Q7n2+6/yiHGndZMM
Es5UEefNjkdZEI4VcKfqhXivZ0SUCkGCIs2yNEkfG7SuQjSJEi/m6seZcLfz1Bt6
Jf9aEbFdUkzj/19CMe1cg5UXw3uRKbDLum8kChwpw48NUz+iU+w12NHMX4YiXBSn
NqNWr4DAK3l1+VK806vwZkKkWLksUnEn10LDNa031RMBl0FPT8TUptcNCY74sPIR
A+rnirOjZvG5gBh5AZrb742VQYJ1khwEazHhNQfKw16xDtjJxRzIknxGca5tjGpY
oTcyG0iEhKzgv6r8n17Xq1lCLcDZlHJRyLz8e9wqyIVXZ7RelUhQqc7gtJ3gAHOq
waFtG54uB5nrTcfxcvWWHy7lB/JwKDX7UPCzYH1l2w2VL+B9gs9O5r7yKbp4YA6w
Pj1d2uXPzlGgy4omUGJ4m1WQskTc5eNXaI+/9zhMmzSj0lSj97uC1SfZoOdwD1Ct
xIwNVBdbGdZJ5XPe+jogV12QPrCbPvMK5D0n/7YgRbv9rsjxm74f1pPQv7l8pSKT
teVo6ZyR/mduy5Mk6Jb5NrF47gnu0S0EN/iUtbkMeXu2rwQ1kk9MWtFghlqQQLn5
9nFabUFEtR8tHZNy0fLJihp4zAcUXDYwmiU989hPGC9jEEMUXS+GkWsaVvJ1UP8V
5/uGdx6q7OxYdP08OZ0owAPjhRBPP9s6ouLIzpnQs/7sl9kTKLFR40GWyO5M9fVy
gYs2jVd9akEFZdglu54dfhi2PF0y6c71/+25qAjxVOY0k7Ff7p4CA2ulGFXMC52p
H7Nckc8alheIiB4QUvZgrRRxRc1Ntjt88f/34HJvE9zFV5F3OhZ8fXjMpbDQwNz4
NsDQTDAtQuTSfsD+UvPRAB+aC2vfiJX7nAv9Y9+X5FC1ufnAS5AxzxJ4SaNIA1zs
LlPnqAKk3b4mAnm+1aX/vgyo8UJSOtQfWBF3pJiVUcpoA8YhX4UWYxEo5274dfWZ
GC7+kLNta+j+pobeQKXUzE9jSpI9zRw3buWELFGrHuuIQx3lwqEbN/NiY6c9s4vS
bgC3pCgBNr4IUZlvUkrUFzIP0d3coglymjpzYRxAzOVA+amzBzu5qToQhlA4+n40
nZUB6UE6cDCrebhEGQ96KMD40JM45KK9tiII+oRYX+K+o2Pwip9zFQIKspjDztrH
kL+ppQbWvCo7UW8lC16h6sEjXj6X461d5Xtq2wscCwbfparizOe18eoXvTNc89Fg
Tw6bZDStYp7hDgJOz+X8h2S46XMeR/sSqCB7LFkP7jVdZAODaE78ef4d4cwvghQq
qf4/CkCl9WYmdMmO+5VIHR4a9rNSTygdKd/YqtZX+oaEdNIvjN4CdSsUMYDj4flR
P1ypB422Um6G3wtdupNo5xlfwIpBe7x74+uqYiHXxUIGWNVeqBRzruyzjpNsYJ0I
CwCQHgGtqSz6KlBTXayaXmysmfqDaMjYt5BfW5yH10+UOyj2zXrbK1ISNOCZ7XTr
3bV8rHjt2NHNvhoeIXGtyC1rHqSwJnfotwLc+AeroAgzcUOirOgOOBN9y/AmYdQr
QxupY/XhiOne5IxgWq8QFxjDuQqTX1QGQCif7/97X4DTsfrJsNYc/3cO0GMMxWSA
PUerL+hJAdpLHrUcYH1ka/GDGKp3zpzSB3cT15/qZzwGGSApdlnPJQj9FJm4FPgB
uXdU+gAHPFeLIefZzovlLIbH9RxJQdzm3zANZ4weCX2RGeoEaVZvtZFYFogOi/7h
Ztaulcp1GkPSY6qPw2op0si2hSZOIiJndV3euk1EwlY17FtIRsTwq7E4GWth5lt6
e+1tb/oabnBFg4ETIRq+1XmGAAy4QF0MqpNQKe3IbyIgPSafU/VosXMKPuR1frR8
PwnfjQFjw/a5GOD74kPMta3M+S7XnDO1B+ap1af/Gb/bjxOi7SiISO/SA+i6VOHP
yNepcttTSBJBp9C4sVraWtgoc+9pIf8wCXker55JVbbf88yUeOiAJlGpxfArZ2Q6
NOP5nYoswuR8dUrQVA01zxbXqwWfF3+zXpYFrwFxPYs16EF/EZBUOsn7UDc7RD9G
4jIos6GVQKycJry65IZZjDzH5fopPQe6sPz0qJeHMCsLGqXDOHt//8PKkn/jlCDN
Zyd1itVkKOb9LJQQZFrL/qHhdhv9XWeFQ2XA1tHq74bCiBpWKNUn76sBH+XoXGUa
tI9ClcjfWce5qY1uPNWstBHbrO8TLQH7n9C5xWe+pkQj8WCR6uarut8ki7M9g7+k
qPDRt4g6ngBzGdWTxscTI1HjfRMZeE1rUQz2TTCXZ3Bas7Co2FhC4XW9SOFhk8ml
tFjQc1iURJ0O5yD1z8zMsazoL0ZuHeJIS98Qax8DAb15Diz5mlQ1BqXay4/eJrJj
3KADs5jykjlIo4KDS8YkRokeGS9Be2JHgxnDCVrBKjlelC9GuFquMgv8elI2nXcY
A3BAO8KcNxqSvX6bxzvYHmR8JruqVNj+agdMz2uYS1BuceYBgXo5Y24iPHtf1fEi
VUJ6QcpdfSPvmpIvGs+LWc+wg9isckNYc4hL/F7lP5Xlnd93uT0qbh3gNFmetes2
uz5kE8YL9RLaH/Kvd9XX3fi1cYeq5MmfbitkVDzynRUtjkph2onfQLb2vvs9f38i
zbtMYYbtC3T7LMm/YV4TS7eTGF7Xf1fBxtbwKcqLtnd8ayPynepfkKFHBHauIlLj
bv/Ctp4D4jQEXOeyOOpzAH8xPDUKjLmmY5BIn3CzrQ9TwctwaV4YDEIQRuvMx263
FyP9s5oiTq2ttn/jL85BozY9NuzU+AbSNKWCWNuWu1BiczvNn9OuxqIDgecfYgpz
z1NXpNVXvlRo1mqcmNEeLJi+8Dc1ExRW65a+/uOlRWKrO09wYxVd5cfJy95XSq+o
OAcx6RQiCqXnlKcPczX/0A0i3wynsUn5/sYy2JIhbx0e4ao7D++c1PZklYMv/Dzd
+ZjWd/zNX9+RoxB0d8eeWk4U8H/yo6Jk6rZRF7lDQkV+d1sc/LoNgUuK/hRTappe
P30YwO/SUwDBGpCzUmdWJhxrex33GQghAWq5f5eIgLonbEu2vgaGHWp14d/1TToY
8PAqtlHiBJ1MAEbeZaAsWimNobDVvVcH+X1VwtWerIiiCRFvPOasuZJmyLjY3lpz
0vzJwXnYgWsRUId82Ya2YZegYGmNW2TmRBui11I1pdn/deEE8uZQ1eYxcXlptu+I
kZPrlUXZbJ+1eKWz8LARMn24d6laangYOxDGTfz0MkBR3H3jCOuYY354NeSa3e3C
12CgKM9jVmiAYpeeT95zhvwVSA9Edtkg4uDWYWFz3ddxISpiox9aaCtkH+B47jCB
tDdSdagSceRobfn0SMM8Tbwll8tFi+mDTaDgZrwqhHfI7a1iKsKn02arJUFrjBIz
hgqXgl//1MAqRye1DllxOETwIZ9ZoKdI0C7TxqOkSrT8Ns14U2BpB+hYyOryXdXV
TRb8EMkTiyKtV4vKUaOLR65vOPJommBVWU7zmsBJNc0HkD59MD1DZFD97lf1fOO4
n8ayQBWTRTgy21vr7LTk5cOy0BKAOgTY7xAFEpBbNItFYFWWApV7QcQJlT22Hd3B
X0ZWgPRSRsnf2XKo9Be6yAEt0Kbw452aMgrfIfY2e8ptYS+Hi1hx1kawpydQIbPb
fMsQpqR64L5se23bo+hHRUdPKh4PidZjNRjFcnRIeg06EvbZOhDhXjCU9jm7bYhK
6xLETdnovfQcfhJsQXY66Z6ZswrXIp6+Xeq2DNh48cbeORlR0rqx+Dlh3BDXt2Up
Bcy5FxH3RlAAAeiJMS5hva9vv9es5M7m1NHsPkrjnoGH4P4mYckqeFASK61zJqVs
XubsEckwMe2pyvHo2EdE4zgNezBs4xzACKDAuNmU+h7+AfYHFrur3y5Lligc23TC
0vMoegAamCvlFvt7Cc8Z3XcqZ4M436Kq1JhIvYyPjn+x4zYfyATucxVaxxLoHB4q
nXVumwFa/y353qj83w309Z0lH74UIR3TvJKCNd/rJ4QBavIveKS1QyvmYngf39E6
CTgIQbiJkpypIJ3KWlNnVgFl8pUlcyRkW1tB5f0wbPc+nIvpqTVU/4FcVS0bjs6X
LeAXNCXxVAfdtZr6KLcZYfMwdqKZNwTrxqf3Hh349akQNkTcc4M9DJVkFO+s27Fn
DF+doMtM4sJwMwX4ALCWqNa2Oybdz6RbSm1/z/bJSxBj/QuPZTEoIXvdiWHTtcIW
86mNAENmTmng0lZvmq0alHe1PW+9tq/AG6JZP+Tnt1ATYSI5ZDEph58vMwcbiApj
R0PrXdA4BNW6ClO9t/+JIsaINMD2TrMPccBsfIlnZBKFr/3eo8sJjhBNbyNeOto/
GucE0QRp/QJ2jDoUq0R8dLYjJyb46BqBMr2qGHsI16MUN0hMkbYdylohg1a6QlQi
OF+SXJsHBPCY0sEOyYVU0CAyIlX85xcWvzwR441mVbBZfFgUFnEkxUWhTVKBkJZH
VUqIAlGK/cj/HUoe7tH/l0OkP8GsU9GWFycZYXtVpOar3Q79XB6su6HlGJjTZ7ay
Kuy/rcAja4gQUHpw29AHBBXeHyUP14AAVursC2BUyFQwO5IJawBnODrnFMTEV9jD
LLI0ZGxAgpmzJob55OG2oBt84GTbUX2LC8HUtCT8UJn+Z3DFj8LKC6peaIE5mezd
YsDVYHmysDJXdPMVu88UT0AYY3xNe/PZ+LGFFbSFaLSMq5q8OzpmCJLonPvcz8Rb
mByFgOH1hFL/5jkuVo0swFuqEwOCkoQ2UnlT3XJOV2aowsiy5kxhQU9NTwxIHzVA
TQ7VPslHVjsd1SusyhFGsKNyvO7zh8tfgjmF9nm60EnIE5alfgAy2sa39dxijhsG
AHHFhdqdstkWrEarbR/YDgOuaRAn9C/UnmHGqdd8SsMoWdbYbwhBO4B3s0b6zsw8
ID9wmDiKn/tVPJiVPadE6HjAzvTzdgZVrvadT0nY07ul39vNgqo2I5hcKZ6jSWUU
+yQigf4l06A96e3kUAoOAwWCIFdxmAprcq2sCW1XHbF/ye0lbklNFVht4+n5IROT
IkvtJzonEG54SVk/yzcsMd9wpadzFdpeu7pMm0ISeinzOLkD37EwHBvB7tiF8QCT
+AuEGpVUeBFfgx2r5djZCInrZTW471GBDiwM6vE4UqpFXCQnlZoia6EbEaZ0d4Vp
ZtJfaBQEK4oOG/oBXkH7bli96ShKpxVaGKvEiXtL5BAEo9RpHZ+7lZMUnsm9gdKO
swEo4T5ierLg4QIVn59R05EuTjMQSYqE6J69ehnhfpwdTjr7dtrb5NVjngYD9HKK
3DbBZDMgkTS9GSIbj19Dqn6GttX8W9fSdLZcVtrRFBun7Lkk9R1RyngU55cT7F4V
tTBoE4XqCLgnuaRi9/d3FXtm/IgDjIi8ZEz85yLiWXACYlShuLHkODH2gZzZqLsX
dfzuQeHiCcOlpv8NsgyLprV1jY/iU/cqVoB9E0YZ/yzR08pzB5rn+mzy4zlMutEM
KlmhLrzcB2dm1XdC3RFz3IUS/XKGSlWa9Y9pQAsLG0PMp1hBjpu8fSGXt8tGF4l6
Is69P3abpczKq6WL8Fmtsp8dqO/T5hoIeI7NWpfqCyQBiinF3zmJ+zqwLQB3YzNv
W3mHKX7JWMRXHqSx1jh+UPwCpQaQFIsqnV+sy6JHWtZCml6w13NaICCMRw5yAF2N
QnyFtUBMorQj0gC6beTqoXkp2+aX1POu2hCh04QmKktijnfLg2fko4Gx41as7Cz+
vm+Fi2hBAl8woQCNjxFjT1B1QKKu7UPx0c5/8NtzE02NcaCJXY17Fz3Yjl4bhqta
ktXvSzzNxBjqj0149JWQnTwR2JDYmkTX3QiOEE2yWgwoRpbDXZ9DHOk6luAYjBWo
vYppLGt2DuRWftQz4rLDhDdn8Ghiy1tkwqyvfK8NfNurI4fK/a9O8vmiRsBoT2QR
OnM+izG2tQBauGgbGgasDWqqCRNnPclDAMrnrcSGJj+4r4jYLuqoa85CgFDvM9ts
vrcLQdzf3z8GW4IlAxRfeUMWJxcU1HtoEOOGE53qFKtNJQADkLmtGi2jBYTEtE9t
/Qgit+hAwwg/4/x6ykvoXUtwDlxiaIWmpbjMKBKqH1tzRbvlbJfdqG755+UvK1oT
j0j32xoiKkUrby+FfRlfX2XD6Xp3BvdU3FBDNWVBJtBrMIvcqDyi6Btfisq3ubgh
dpeGUKJqfIi1MGPQP2dUMGcWo3SiPtI8Wc88MAj4ha+NC0seRcoUiCYS3DPx6bQh
PKDdfmojPRdgdpTW2OhQ9vGk1WBpjdbDaJdyIpgXvCAnXmi7bwV9xO/ekVvaRJmC
QzyCS5XktT4YjNT+b6+V/9C75E3QvvM4xZnQLQJjTGqDnI+ciCY+C8ITf3PLETtc
NKo2BIwg1WWD8cogVfnUM6KoaW1Ehpoe6mxkGj29C8v1P4SE889W4DPnih5z990t
H7pTWHPkZb6Vi0wVgOaYQEc7rT4ztaonhQd0lVIhfuqd20vha0EUtVMOHkBIwAsm
2j8yT9yCZ4FMhrJikOc3m/lUTzKQaMaIpP8PRyzxC4zuMDkpoKtT8pZ9Gr1iOu5T
GzrGTXzcgLR4VZjp2nklRSFq4XaZUAj19j/mxDRdwbKyVv65Gb32LjPUd1zSqrd5
fcuCPDKMguCPqhCEg1aNvHoXasN/Fvi53gPzeoajWLi0/X98V27KgRfTKcvswPEJ
jo8Kfnq9RAONumqFbBwjOMz59ZBgGRJgNmdhlutDkU7qmIn3N9vIva8wkxC0h8Qa
pYKkpLdGWE/BsEMA4+p3mf0FyD7XECJ0Y1NUVG37qc0bs31Ac994mDWJE28rVEUl
+VsFmtOVNZyW/7Ex2P9YqaGfHER9CPsn+7s558x81Aqg4lOkpifLlOCNSDjYEJHs
KzQ4CumkuNuYleY13JRh83OsSPGxTQbhsspqI5b9Mixo2tjtLbyZc1yQl5ORBOd1
9+UhToC43GhYHYRJFGpJh2VyXZ0T+Z1JIV/57gQvomXZFUvUSdYXp8bU6HaGp+7U
uWHn0GRsfna52y7LtK678SBDC7K+0eamcDmEw3UMZGk6ScUhVz1wnklw9Z3fCYop
1BYqJuMPcGSszynNlIulbtEMNwqJIwiQ7epvbI94JFoy5n6ymA43e9/mRzq8u6xa
LC7WnXxSn1CW/BVEwQ64gL4gajDkA/IpxzGFSfY/1WI815c1hascspswaBj1cMl5
aprgwHbBwFEt80ngKgW7ksH1QKRrSUWPEjzy8lORQfConH/Txk5c86+SQDwJKOf1
bJZ7MMhbTfG2QnVmUViaTUV+ZGZhHU+33Hatbxxyv35HLVnY6bazs09pZ3pNvd3L
fNgqbGf8e2141OZ0xQd9Ssl+ndOTPiNxJpW9h4/ulv5NOFzX/4OMudAawpul/2op
QNq0GvtZqeK/xSMENMxBVJ0JfspV6hMe8zD5F3b76X5lzukl/zB2RQs2eCQQonse
iS/147XIHF8s7HALuNr05YBuqizUHGi2yDUs3On1Q//EDjr8lrymqoC/MmxOUJIA
8q/4dK/L4HFhqcKohmNf9AbeBP0Wjcvq3qptpGSKB5/ZfvVix7/AUpdKPzVeZGuU
2QutnDDNhXyL+0h7PTh1WaI8C/3HWI+O6arDmGllhW/HfJ93IkNv1lWwu7rJUdou
vM/vN7hEid4uaPbpxHAvkRCK5V14ifg1Gi+GOaHrQuoXyHvNsEdVhjAJ0feyhLWB
o4/0rQmQD1jB+G9sPHSFfZDZ84hXxRTC2PL5P9vP6A97Mu4Vn0R5Y9AnzFKmZJc6
28vA/sknWOgdfhvBXihocZR8h3ei62gjkLlGhat/dbxaZnfDgLRqDe4VioakAUGs
FgqqIM9O0x9xVUQaW+EgiFRVS9wXaTPW446jUDzffoRL/3Tj1UZoP3FWVOJnLL3J
NaoYhlCxZl+VFgKdYSzD3yqo0i3YAZzsLFCwWt7cq+NCH3vmM5BAEF6T/YvJejOU
POLTMfhoFguUZUCgz60EX/TSb+DwjS2746Ct4BZcbZAVkOQtzhLIBe4YOEjcdzCF
AqVOzBK0WRpo/UY51VgoIydh76U5sj9u82q0F0TamrgsxmDoNHMod/SYQUDRNX7f
LL4ydSH78+jygCwITLipeez7Va2i/VcbsUAtcpuorfWjmif+OfPyB7LZezsklTcP
tYA4u6dEo3/WEBUdR9vajFohfG541ehi3H0KV/VGJGnQuBVS4RUOvb5POcK+lHSV
LSRKs8hdcv7YIotLdif/lQciLho3LRf5M4oCImbnLLq/pq86FfTA4uWK9GBFn0OB
WZmciccy3pZzSGno31QCkoSKATJLDaqkWdomSuNJ4ZQ3o3Jg9WBG6nWWzxmaTkch
BCVU8PbPV5kNEL6zHZgHBmsYg1iEDtdPMgig4NL7hoBlpvh0lNIITD/CzGa+yFot
gaMXA9WVI4E54FvNKkw75BXf9wJjoRQNhMJUb1WEIDlQOg6hd91e5dueVKJEl4K9
SoXPwhgEcDvero+jtGoqcdHIp5I2teQC0B0Nt3jzVtHMUL+w3nd27djTdmlXx+YI
Zcs5dg7MtFng3yYT35llWlLbDMmrcib89W7JQjwXLI+UfllBwf3CFbi3qHUlRxZo
Yx0Rwd/bxzS54ABnOgpNzodGpLla4P2srpBw7VbnxYSX/FbWClS2Z8MdxeW2Sp3Y
aQMnHKF6OzFEfJOc9AGjHcBdRM1WqrYjMK8Q9vomPzs/9Q4I0xOJbb2Hp6AYjgiS
jKfli5xt/kIsmGttJbP5t/RhGQ+xOFnrnOG0KMnEz2LPikjuValLyWAEaJnM5sAu
Z3uQVR8i4+Cxmg00GyhXfZE4d/A8zb8ptcYDbMJuNJjeOaCAQebnOjt8YvjKM9xE
2VnIkyyhGFDaaPc5vyva1dki7+ltnDWTC1ZfHn30jVdmCADd7emqNODF808CVIbz
PMhWGfBNAT5oPQwX6Viv92iPSRJtkrm9MZD0nmeBWXw2jgnTh434kRCDmjO7Gdht
08na9uOXETWwSZOl2wCnP30bB6yrljTUVlL1fGCfhcDssNJt3iooVlRdRsfLbqv7
gkWpMKWYpgmRE+0IPrbFsb/XZIXeXnIgHkNmJSHkwbFHGJHV5GEeCIe8CJd6YkiW
qRYH40jprl8Nz/Id56y4s15z/fxcoM3xeHXFugVGBRMJLsrLoRwDNUxezfiFdbxQ
ouneilyZ/vuR70tSXlQUcqEyMp9XEkevkRE7u6pqik308p3nE/xIPL93xHnOUgmh
0gqzRrLfTQYOvdEf6P9jsYxi8eTXWevnt1KY+ABViqSCPCcQTws4xx+pRI+DUpmD
O8Ygl/7ja8c20CkdZiPK6esNjWwGGgpGI9YVIWID3VhVdWPuj+FsTvFouitp0+Sw
f06UZsapXk+MBHsBR2lEusfsEu3A6j94iq+pSz3IOPHpFVMGES4vAfwd+tgiTlcU
VvJwwWRd/gMOfwHgHh7z/n6Loca77/a1Xy7mdk71TryvdZ76JOQcbTXNoG+irv8x
KsRZL5/St8IIquoiQoPapkagILUVpG7x9bxIBXhZNZ46T3P9QJ+VPTCeUr8esN97
8gXUHAYml6FC6pK0SHjbaH/vO4yEYuupbCMQi/zmiqPbkSyUnAs3ProLaCv59ASV
QcCO4CIVMF7O0Ekgpwd1xUAMpvcFltF8/6HqIo6DILx2BdFR8DHb33H+TotkPsTy
FfpvHCHikXT0lJxxTTryzcT5ydhqunCdCAeJDBkATLGpok9gBsK1cv/iP6eEOnxS
hFIBQdGCf0FfDreGe28g69krmeZYeoncgj/Hv08VtFvx7nluTa47JYM9FUf2Nh2l
D3RRBlp/G4ZP4voIOh/D37Gnq1KMy65irjIb8Y/km62rQx0hwGmPLnuGQTTtKisU
U7IeH5i36extP/oX6DnH2BlLypl0APP+bjEwMG0wanR0WzIkdck1WENqk3evhoST
8goI3RLGolmlRnDmg+JhNBgI2PFxy5ZwtoB65jgjeCjAUQtpYoAjbuKX6K6epM25
hvPUu/MXxgwg+/IoDSeJizUkDKRFNPxeDagdwUXUsuW8UGux/HqGEIOMJBPs9jqF
vizoVXRe9ZEAkQF1RiW7wEv2gYhajg49lZEyIJlA6jVIUzd6e5eNEorLN5Fx7a1U
KbXzhQhNq0+lBHectcyWqzWZmBLSaQ983J+/dHtwWdA4ccoMLbU1zjAatRFK9Yj6
9N+cgKShjHVoGLDot2rnmexLZDZtZD5PSVYi8y0ozBTqN7Zk7Mdq5yPuRZuvA5oN
m1CkOGq4dcn232lK9ZExI3jHkTkaNma2DMdmr1EMPR6LB8riP++Gsw3dbsdgzgqC
SPSZbPXoa5G9Bk4M0URC24faKfAEVhEm9XxY1yrc+6TZWHB2LU6uKpNHy6hCeiK3
S6f5A2jKqN6WtTlQO42ehNf9IkkkHkORCHFQtNEOGBp0U8bQxPL1pNxJBBt13FIo
2LGAr0//g/0VLz8hExrJSaregJQHWoS9ezg5ga2eL9tiztZ8JrQAogCE6r/4lSrl
Lbu459EhZtl96MPEw9E1IbEfdWD50uT6jQa5ZTQ4V5UV/4/LwdT8x8CO0aOdmbYY
HaTRP4qoLGzkOCLJkHbUqfzudMtMVPAJxg16BISa1gistWTjkJyoYdh/SQPhbMWO
6M9rFHMiB+peHGkO5dEzrQiD6Ymsi1ZLfZIV8z6/BC0RRZ1jMK320RhFbLYAuoXs
MngR4oSwfNU7i06EPD+lxX8LGBT+d91PNWF0kYpB32aop1xwwA3zzB0PYFamhO4z
p5xaaYLB+3CXv2gUNaSuboBp2dYT/Yw4osShmsZVAw0iLdPwo3Pok/L0PoHlii32
DgzulZsV+9wnmV2n2F6/gkkGVKix658cWa7U+/WnBBMje/CpzoiWPe3Sg1uJBJzg
sYe8qXfYH2qcjbwH712Do5pI7Tz2CaenzObouw3ACtu3hJlZMgTP8EIis7tPoWel
9nPgpmOxoVRKDqjIQKxTbdEbOKpKYkC48MRi8812tlgffZLIlO2yiDx1ErErGFPP
FOjIa5Xm02WBNJ5DS7B6HvpqsvVTPOLwUroVZC2YhQx2lavgGKgKz3Ig7W9YT+JM
lCwPJPWXiIVDS/fMO3xIuBrxQjnz2FHp9oPa3vyeh4ah52iGleModbtM67iS4ucK
uErz2VXjnvS/TuPOHOVHA6geOGcCDDxJaOCRasUNdwnTXPmIrTKaenK5xivedWsc
ZkBddIvy2EnsvQ/JI1wtPqaihN62HZ1d6UbXu05ekq5yjCM9zfAvYip2AYvkYNEt
DMNOTYcK9qa26dXjDP2Iidjn+q62f8rhT8ubiwdNKIDBxMu551nIHrTEsVIgysiV
aEIwfFVz4egaP3gG53cDRh+tHJsFF0NdTE1ZTqVJDUhipxqEyn4JC8jsCfZT/Ny2
vT6tXmRPjIxz+I4n9w72tpRlo24O2p9xb9oJUbps4X3MnVF1meeCfzon6oxvHowc
BrdP55ZNB4YdTZMvhJD2I6Fhx8G09pTi5ekBMYeLXgUC0VtKyZ5dGLhyQoILfjA3
Q5vmxykP4u6p43aGOHQCjKlU9l86V2ArNvn8Qt144Kz2VBswd+JZu9q/UQsm974B
GiOlLrMEvu0gHS89I8IXVZfIJH1PdkPUU0Zudg0JAB8/0NTP7aKI9DLtEZJQ22Md
5cHn5nazCMe8k3zVxhzwyZiDRqW2J2R4kvXVkYLPTXSyH+KT1wslw1j6/XN8+Dw4
OnaIuc3zSo93Kyp9ziMFCu3d98ANVq1SssfRkab4OlEhfiwcvGBHawTehlzmqTv+
NhWZgsblc0cLhBBhgfRbIRja0o2yZ8OsY1DAD+gXmH1RPp1AWHJYLf2qob1u7XM0
FScRiheYDw/jCdrS81O7xbA8QQhfpQVp0aJBypdFNdRCXLZ94ir9reTz5oqcY/J/
cQYIXXMmgajb4VDxSkvT2wo1yXZEQLxYwF9YXf0ueHm8/Ck8Hu8rL0Rj1HCfxJqQ
lkIT8r99I/REmfGjSqP3yzbiEtplURDLISWZOCWAhoHbs4xq5y8jj3ZRbBZc4ZtY
wSGSfrWC2TsRO4vnPrHpVX4jjh343+Snp4HK0AvKSw/e8tY/ofSsDFuhwEdrjfZQ
0iKS/e2QFL9QDhSwavQwR4FjwzI9Cb1hDKVgRTIEUZcKQ+CH99rqUdCaUXF/Af2d
TsV3jmr5vFpN1DBmKfnGMUt9SCzDExvxNioyfBQlAyM2K9q26/M790SYWMrKGylw
/gSWRdYewRlXizEOHN1/vvw6ypNI6J4w3pi0KVuGAeIcRvf8bzXq0eVx5P2vagrr
/cgXvJOpCN96byoaRgount0YfIogeXWU7ZcZgkdgzrmY6y31n3MQgmGUYD2LxuMG
6z9/DXtVgz6ipEUxiehYaq+zOp9mXWNj6IKz782NnnwElEJBMg5yiRS7Ze6rW5lc
IXjK0FuPdfas2WoZtWOndd5VgmsRJUaybnYgLam/ZJKSlgmVJd2LSD8nYbOz0qfw
g/2SFGHNMOyT0TESHbZ/s5A/MSD0lXy7lYrC5RDXtW7Qg7HCQUZV3W1dFOjEZMVT
ELxeblHHFl2gb91CT8uOSSu9FO61b5z1wlPyY/6bpQY4V5FL5TzE3m8iD2xAEPBo
YqOA1GlmGces2aFnnKU6IaYOm85EoeKWzAP3k27/pqCoAqqwNcISrYxg9ou35DfT
F1NnqclWGqXFmrZ2s921zd5big4u9Rnr+aWswllKv9KQum2SsPRZ4ywUCpQE8ma0
Mi7aBnf7hCPAK5ufeBbbpbc81lm2y6GYvv7dscKJADQtNSa4CkEB22vHDKptUxKb
oHLOBOoOhuNkRNgxdgHXye4Z34unFOKYT6Ri18Ln9h/sBYz1/duxcqR38paxMEHM
ZKd87LVsYBjAE6Enx31kmocETRLtiFEFcmBQeKExUOuv7ugBL0W+ZSM7rmdNBAzW
g4PXMN80zLeCIDRRttDQE3h5fd7G0DaN00KjGDIe1WuzZAl2YXPgsSDmgF1GaQQw
BRsm4+GbM9CTQqqyKod5796GdvA2/7b0xDz+Skbwf02FIBdRGWrayG/EAZe8XpIl
OmYVWCbDTrT3hgle9bhasDoJEYPsvT8+WkpzI56dW0MLXvEkgtKdPhXFgxKID6K3
/3rj0BSbHlhY95BEs2ad9YlHjzZccGw7NpGPjStBAaR48bleM9t5ZCDJcV7tggZC
hqukLyB1juArpzsc2J5hjVPoIf6+Aak/K9eFaoj2q+AQE8We2gAyrcxoCLt5piid
3r+fqmHmxb/WpJ53ULesSbLLnLXiFqdjPhbOwL7EUWl704ztVEFmtjPlPZSqdjwa
CkuNOo1SWyhXPhRK+Ap0L2ZBhOqLJFplnt0Z3p76GuDh9cyHh2+fMG5yaSPhKBAh
2QIwhVqoIZfsrOUHh3UD6l99gaR3ytVyc9mlLqwMaWBNFGIvlXOelXGiIZkF5eLH
uMzQNe8Ic2UwmrM2nNhwxUdtXN9D2/2Bi+FFIyiT6XUwktTZ23xyaPy+ivXxrTYf
57sQjFLf4A4s6r0zJD+61YibyM4y29XFFsKetzr9bsEpOxqRsigg2ngWlbI3Ajw1
CU1QZami49R/dSs32J88cJbk4sfC0mMCC/g5+385iCROD6NQ6lXfjEPlMOnMbO0v
4+e9XNNV370pGHDPaHY2eUvxGNQPUnBQgi0XKPzzfIcpiujsjOthYkX/ROLmvsyR
4UhOJ+F019j4qYMgNMKMqswur6XnD5SVRxA+dISkQAJ1oiFs3ZMBtI5JsrO2ljo1
tvnwKgKOkiy3byt1FHtqWHiGOeZUZyq0hXeNDY0t0sC6kpBls8fNEQWnAZLH9Vgw
9vhOFj5nt53FuTZAKXzI6WxeD92nDr/qJ6r40ydzD6htTyV8dt0sMOCAhDaBt/fE
lGIUnk82ckptSTMmcrtaboENa2K1k40d74KcOQAtHfKQuPhmUKOJi6MHpWm9Cr+E
3nP1h0jclWHnJwdYg2g7nhYPzY/7uNT4hP8zwHLxdls01a/RxQVhSvg7IW98gYFQ
E/NUJWKSg7/C1iXgERpkPxwiToWH/PjpnKZvruZEyCgN7rWRxeDiTkn1jidwfuqn
3dGzYWNgdm7+NkyI4Ixg4K6SKR6semlAlJImVz5slFq9PcXCQfbQCFz2Mz9BB+1d
S3BCiFk9HH+ZGczQALGoAHxdYEidAeVIZ6Eu4aFgbKA0UM3CBMLw8O9FJzw7NBpr
iJJaZeKv14p5Kd3yPWFYYOClLFQJ7HJV37StqgOegXCtzTQuUUhA2Fw6OqIa/Xmm
jTdbIHz0PZ6/GVROM/XD/LzHuSY0xji7UA5rjuJyeFseU1RQG9MrDMTHXTFntVI0
nS9s/Oupe5wKg4kN5YW1jT0kPQ7g5cEbyRktniydCUXT33zWHZQcmjzRSRv2SS1D
ufzeo9UE6dKJTWQVJXLfof5jT/PU920AdcCGDLpgNsYaUz6iS5gp7Bq2s5J78+3J
dUq/TtAzjEZLZYFXbDehEzJ2jjDbxryHoGKVXV49Rae89EC4K/lngBSOcyr89FLl
DwLx99ZgEKilWLcqQhzgWsK93lri1XovKprEkBqeAr4GpJRYGAWqtClhFhibTFkl
Smfjjrbdhx3ZyoBM89WWIwMSH2/ABpFuWAnd0tnuFvsoM8SJB0eqnsSO90ezo0ux
EYkQvUTzN4jfXhhuFQMeGv0liZUbs6Av3V9j49ye+QXu8PrfPgWzzs8V0P2OMAgs
abTXyqdIUW9BGiO7V1y8tPxO4YiSRba/yKNk7W4CXSLdsomkiq1UczHazjKCMVJL
p9NY2N4VUE0lWFmOiqlvs4VkYNtHgiv/ythI4sqlWa9CPMISQTisPiHnlNZ8oqNC
FFwV6GhzzxMag8F9xG6kkD4UBPfqkk3Fs1/PKIIrBvzmsKE2Zzf8vTocrCS+kdYb
6Fyoj6EEQtJAzPXAoQ0e6b0n6ZjULyek+RvmZ38xL0PrUfDDIy517+IEw/VYH0Rs
VjWD1SFBkvBiC3cqiqat/R4pl7g2oMk2MDbXgpsrZnMS8fwJBI/m1v5rAN0M7XdY
h7Tt33oLRSfr/grXW+Oe95qjkm2gB4cUbmCZngmHPafz0X485yX96/Wkn/fk5ocR
EcTDJfTbxKlVG8qc1VU5mMcCemC0aGq6g8LKC+UOZTVvLPeCXednZ+hggHKmQ/i0
vV8eSYZWtijz4ns0VUnGKhbuoO1PRSAkFe0JMcb9OykdW5dyTz1bGkuALGycgA3r
dUDwcPGZTy+kt7Vl4Xa7nRSyZ/ZqB1T/mAXDpk8Les0mmohxiF9YfKkcMzuPlY6m
hjnL6lWMXJavZEUrlPlJ5WfEaT6MqugkIwxYLLLtr2SK7tohXCkOmiYxlyTIwcpq
yp2gLrhxoGR415TjGF7IW9XWlqgAEY45AS41whR+aghiitvRxNuSlcCJ3ElLFwT/
7bDmPhHetHaBooYwTEVRHmEH8mAw7Ef2Gv0h4FU0bgnGbI6ag76Y1S+mJfgNZ3OK
Kc/AX2phmU8UzNRHvIATGcskL4VkmRHPSngSuMlWD0TtDJnLrAGfZhbFMv7zW2nj
bRCctc2f3YkP/Ish4osgo8WpPTKaSoDeRSLYzzIFm8wqNiFPcMB7i0wEGeMGaHcb
0SliUcXZoOAMCFEJXcQsp3s8WXq5AMeQK5YveyWBOinzmP2L8d64OR22ScnchZw8
a9JcL73TBbfSXt8BEzB+7Idf1nAbIqdvPBpcnGIMEWv55LlUoXw/97KYrnk5MpNH
xzxPU+OyzC0Knp1tfwdw1yhy6s+0rPE7+ybaxNuBNhPlYkM79+acMoZEQhmcnKCH
bkWms6HA0YDteZ2XENsPHQAMJ2oWBKKCt2AGK5D3FH5f8UIm+cK876pd7lSUs4Vg
QRTvXauyzMGH0mz1hQ37pZ//+StKNr7QKX/2mTfV3tPtZzKhfKsXNZIF4aXV6XqD
Y9cyQg5Erh/y8K+ozROkey0peJUm6kfbSi3D3TlfUpqHxoUwf+G/qw1mPVIuC+n5
PYjfXWKgeL+M99DXmoy1t4KJvB2JQDYhi2VE7J7FIfgs9j16LDrDAHhKvINf1ARw
YfukkPMz3GcUK2obActfrAVwJ7kPhf4yPDNO4sCOSSzH3OPwz2wdhRpHw+iApv8s
smoH53i/Zbton0jUgVWBalhLlx5+qbqff0vuvfbRZk7zOjFqlv940MDMtWyb4xC2
O/LmIR3PRJPsWlaCEFaGELFzmLDDMPqc4IOCJl4OxS0NVfbHLwaDoFsdx4PuYvUs
UbBzA0NaXVrG1dTB+EjCECC2Pz6s34dKXFizMji1Sof3qu21zoNM4X4kkSUlxcQF
/mq6F/JXvVYiF1FOr7x4k/r3uhtaMrfhjby+sfCm5ZMKMKEd1fBB9xmlpTuj+WwS
2fbw/b8wft2XncrgHNA8xH0HncIBmfxM0tRLhsuc641oe8rCCH9hEVbs33VRuskV
9tKw35/W3Sb7qfFf3OAFKZz8t6uXIf8OQWapVMq5W9CJ3lrIySlHh6sUtYV8wt7r
mj5zbh4WsxfOFVAl7yi1G4ZtoeQw7031UaZYXGQlu1LgZSs0fvHoGGPzvLGmI63v
A5p/L5jdZDLMNwif9PbMTFoL+cp+oPNwNDmuHoivvtAuFInVtMD1RUB5+2cHd4Aw
3riTNcFi7ZLwxuMydE3MLvTnEhi69vpJNvhXJR/La/00oJW0m/wW/m7WCGqc0WPU
JdU73HHaKgtF51l7as0knZ/FdIhuKgEovaNnREeHLy+WClTROa1uxkumxLI3Omk7
7aC2ct6vOpBCOCJZjpgB6uTHGvZsV/hdS51nJlo4cUSoSeDtNVGoWGH1AryS7qCu
b2/FQ42qXcHQlJ3+9a7vaLe+8CbI9ktNv0610EzlhZbIbmGij/pqVNk7s2tkLno6
RQFyIHYaO6Rrfth/JJ+ZVOjaGEvKs4HcDAUJuFWUXt96LK+Zvdcm0IeApWtZ8n+L
HlDoIC4VJ71Q6sUI/aCp8LjsVEdcMlNF8n9DzM+PtVkK36zpka2AvXMCNtVO27Sx
bU4h1YKroEr3gDUTEnsNlOZtPof+ccAhy1S2U0kIm07dkvE4zqExv+3Fa60EuntU
9+Y7U1DPI98Xly8M8rhJRY2xxQ/HmXMvLzUCDsm0HVi4s7xVZtL50FCxj0NWly21
NExP0H1NJqaVuhrwPH0af6Zu4yfBnumZrOdPdUfPR7jASCv+1QZB3H6fFKs9nSWI
NLAFw+FnQ/wGFb/V5GbWi8JJQXuOwM358BtahW4rECvYPL50+w18G4oD9HBj8EKP
OTy2Hjg1mv7YzmAxPTW7ghbPxxVkLCCiqf5EY9bfby8wzTEOwTTmu4wO1d345xSF
aZ0mzfWtoytep5lzeB8pfBix89mxNoimsYCNkDqBmLOdFWeNe+a6C3eroTP/KDIL
atRGvzeW3mP0RJtF9sN9nP9ohexGwZCy0YZqs11sYZN20CzrEtjeSGsUwYsIN+5v
WtDbsW7oPjyEbnaQ8sf5rfvtsf628qIqQhUdo6nCn9P2onwkD5MK+10nYT8M9EQY
b4x5cBI/pUnh2cQWE1zEk/qu8A4Z72ZanM7udub9CspKTOIlbNHkDVnnYiIQ8UZG
j0/3fFC8TM94Xg0CAWqt3eNBap4nYh1aNqcJVfjnSrktDqdLPfJXfCcw92F+F1ny
Bp4EqJk41Kj5PH9ry4Gjuy2xyhaHdEALOl0pqn3w85V8eZ2GTOMipXwRn9t+jyuT
PDXdAfwkoMb7m5oTOWKR+twqXWxupM20wRvLQsC26cEcMNpV9iEYMCQLBhZK/RrN
zoeQzjdmQl9hNbST2XgDNFWS3kA8L1waP111RDhBbYsaYeuIaznNuGNNZpUYfohz
jTKvJtoaTN/hLlo5sSEwnLaaTVMAPHDVMHfpBYOMW/89hEXOABlfldSCRR0Rd86y
pYWqhAwovW2BIHqii+v194FB7xtbhKKx76/c65IPPhwF48MmdCMerM8NuwL+cDsE
m+CGqHHH9PVvYuB5r2xOOYFDmOJi+47JQt9piwu7QDmrNWsTMzPTg5y0vJtJ02E0
Zur2oZkZ9Np2EVOfSEn9q0n2xXx8hEracfLGFj2cqr1UE+ZYKRniLCr75fKZiV1S
o9ubaY3X6XBuZQYsuCb1HYkJ8Zivf4aB5A8HLWEGGdp8ksyXDDgGXYEBGkIZ5Ul8
OcKj7C+pUhONJsaefQyxQmg9ghm2+DnSacSrwNUp5zeHWjQ7i1bJVDLtSOgtMqEi
eb83M1NzDwYsoPAiYkBy+jR0T/HfgeAnrt02uyiabhvhSO3aFzZ5gykiG5eyM72a
9DxaI8Fj09PvDimU7VCOgExYPgz5BRDiO+FNbaf0t6soEaE1nCKPzyf8cUWB2+rQ
lxuHFw0vb14+L0wcfnlHqZEBlWCtiePI0hVeMAgWlgSTBLZ8za4kOQ9JkI5/1/P5
a8uk3OIw6mcFnTnbFxEDIv5VirNUjq+j//qxmgZTDtKtm+LsLWbZeUNYsTHcullD
2GAROPJVdIsxx1CQBpj7DknBbktUdvYq+Ft6Y5Vi3+8sUm2Ga/4lYsVfMfsfO36i
Rt8cPnwi079yD9GxgSlqeDM0n6U1DMFY6230g//gcQftbnZpcUBUFfylzMXSA3lN
TxTHB+R9xIXRC68Jwvts3YnYmYe+XFnDKSgkxiHrr77i96vL20z0kZlohH6u+Lom
Hmf2hd62FgRZfgIho6RNp7R3bLtzXPEnGA46IUOIW5zUo5B/BRJ2rRC0xnp94pEC
crOKPJxSa5cC4GqLGzVf7nAZUIVZ4Fz/uWwdMu0HnUfs6oljxNqx6loGGpKkuOLs
S57tmNMcmEc0Nd/htTq0cRUxoPSrYrVPCCFczmGFBDPE9lmpKUJCyzeU2lmeCpQe
xd73Uu9GeZsbHJA4cUTe0IgiipUmTv4VrWeGHKjmqA+ej8+etGHC8xW1D3UxrzV7
+DfOFZfuwpK/hgn9cryou8YSV3YWhXRIwSRX+5ZK2z7E4WZPxKWIZ25rQwsZeMWy
nlYiFyShY73FfGkfzRVEf/pEQYPEhIXefEianqoFL++TKACwf1vX7sSBfWzGjgXE
+K1MXYhWGpnTatcHHVnpsSNTtjVghHSekFZ6Cn3XlRCwIX5/cHm6BqzoPaE+45Ue
zO9AmKL6ddrt7Y9EFiMar3cy89iGbO25Nw5mSgey6aqmvW33iLeM7RjbFNOg3dJg
OxvKxMK2SMcDS2UPhcrWJrw8nReAXjmNbQ2Wv1RTyr8vhj4K8ojelOuBl7BlbnU2
XQdjJJ8mUZXCVgDQc4T+nWSCAyYGZyg+i7IsQaKirE4VXQmFZcP+W8dQTMGywYvU
cpqVpu5K+PtEpp6cCG3YVrni6POcLJ81MPVZAUlh1C4VKfhV3XYGYHQGAxONbqVR
M/6oUQzdXaQpzCu7KCWYjBKkxqfjudrS4u3vmQYdpLGD+qFYyGhfiMPYJRKr0MCV
TJUp+tWguslyH5gxYClfTUO9KlQyQjfldl4G1RBDZSB/xbRzIuPHRw/W7eBfoFD/
yzxjF28aG8E2dwTZa7u7Ot6JGguOpcgZAgyKFGYaJXNe/i4e9UNkbCzgAkzq+dwi
P2AefNqEfUmWB7qxpLXtectaLKtc/cB0KRY83aho1QRf/O4tHsQQPbw1ZN4bZNNz
6ORomxlKhHG2ry36AoIAJnLjPVwRN8UY31gMGvEt3vkQFXP4B5SwDPcieTP0885H
FWcmwMAe/WMbkJUJ8PpPkzUQRVD1PJqyl7gsdIsmTKKW1nKhd/ObyXXg6splWNhn
S2nsSc1UeVkp4qB4CIopChe3eHuz+jxP+kazemRZTItqGhCW/jujjwuEYvb9d1/Y
PcWp8ttKMI0Vt2vWX/wZQyXvpFq2zCKxTa9Tt8fvoCod6+64jRfPq7oSELCD2v70
Dmf6sWnkFcjHP+sBOwK70fsJDHYmYtA5tpFSlaDSC6zvhBNW+mL+7pG9scWBFkzb
SifJgmhRY0j7fkMU7f3FfknBfiRQwlWcnn8XzU+wM+L9aJx1kmMdyimY/XCM7h9V
eC3LqKLLbeU+o926lxbMvPr7Ds6EHcbmcJMdfYlqjog5zwnc8EEfreayVloMtfVm
WnWie8stK+xvxdhmc7g987jl1x0uzi+6GR9T64QbQA7jkstoHpttODO4bCquBHhe
x5RyIsn0HQ2StTKu4j+a1/W+iWlE+VNOPjuyWnlXvwzAYkoDj/YElSIZBYAIRzIo
0tFLT5EXGSVx95XNYa0U50D8Stjwg8GZrqfjK4AE+5XPFjwKflfWetg28YvPEUrO
HkDOEGVikwIlOWpPqGem346RzvBncBfKioEuDVhglIn9jkYXx3UY2nFcXhUIHsb2
j1OQZYiIIUZQXYPZgGs7kwL6wUVdOoQSNqJafjW4fzAJ+2rEK/MK2BxNhWOurPz0
CC/28tGnRtpn/lWvBSGKHVAAGWFzXKsjRkLe0eLkYlk5VEjZIY5DjV9XTjDB4zCg
hd05jGQzvK0TvipXE5+t2LhwFQqvkOkX74JnZj2maUTvcks2scpINNynEUn2Y3xZ
kIG3pJn6I3uTxjvCR7e3Erj8jhpHuT3q9dk4zSkaHn8eO/Z8LaYJDB6Mwuq8yUXX
CPCs7Xc9qWchKq5ZNY3c4VVRV9cMNA0YrsEZRh9q0yIH8OqfoCvJI4Mrmi1xXCIK
CpaN0GDTK31PhpBNeWgpu4Wj/2oF2gsE1uAjWK/GUdNT+uA/fCU1/EHsfcd6U3D5
LLlc5/JYlZGNrhsmii6a0O954AXmoC2kAws5sJsfahBnaZRj0wGdjqota5B27b/1
9j9Di3bVb56oW2Qa0fpLe52LI9qeJyIr9uGafJaBsxht5SA9CO6Ke6gtGhRIyypD
llVjXglbDBeSPCdnfB9ORhj4Od12z+8vAREbvuZFo6i2O3pJqSGO2WF6b+3hHky2
nWSF2V1qoNNmfVC55uPoAUdgKDkmUyTuM3w1kyEW5hEgv9Z0FMcizWsMz57LFoBY
FpkKeXuvPChcVsRTSVQVy5Qgh34vXfkY95SXcfO16ld9k6DxNh0ZJddIatwE5biM
9z9+YMqH1ExrhE2n1tgq3L2uGYF3zQy4jH7GxKJAnmnuKj/MdSbp2rEkK+ZMIPZF
L106IQRZCiNvanFAkBpR4H7SadlewQ39LLYGSqm2iyCN3u/QpX+6ZyfZo09ps0c2
kXLO1pUbUWxOJj1Vp2vAY3srT8x7XXE22g9TmBGKPidclXW4DCTdb8hxPakEvL4/
wd7HJIfUhWakFt11vwDqIaQbzG55aLvf+V8qStQh8Zejho+vSDTWt8VfVYpeVG/H
YEP9GIQ0vdO6ZepR9IhAePKkv9okkAIqtRRHsxoy32ElfC+NUd2z+JPpXrgtwVDm
m83ktCxoH1m3ZZfofJp1rxLBvaVNg8RiAAWLZ3zHjSGx5Jl9+xnrBHsA3sb1+Hj0
mZYmfNl1bfLYxYd6DT3svNgHRbJbE9DyW8e9Nk01BNq1O97UR6j2P+OiXmBPEuFK
nZQuQaiqmWwN5d87nhrJaSkHqMZtCDcA6Z7G4fmV/bqy1EfCKGuEbwZk3qf7bilz
aawFcEnEkMw/eisyHlK4SkHdjlxogDufAmJtrjv87tn/3o/ceZM5Tnt5rn+S5OlG
jTGEP11kpBPCcugP43hnhsnCfdeEmj+r6mea1ssCinuvaWTft18HgXH/5UMc4YXu
WrZJI+Dcx7NA5zyi5RPIzFuRk2/w8SIro3c7fn0NJBt1LL5poHUuSfkGt7pDtZqT
3XyUZKCBQBJ0ZoEhnQyFXkYxRsbbtdRfebA6nKhkr4/fRpPxYfopqrtsD5kwE9Of
WgHDefHwv88zpMSQTD076AFJUMeaUHwN5W7NU4XnHLsjhq2wjWssW7tktGxoMNsF
D18ssvfJ1IUvwa3demf/vt6XDHjmrE8bu00kSs14662o+QrE7hiE3MWBHb9dkDJ7
0XVqib5gPhYUZYeoTNlpZqZYBuGGjRPDV5t1oj5JEGYoI9i5Deo2mpre9dL0wMJP
z9AGK7XiY4MQjgscD9O82YsgDsotQUe7XuK8nO2XHYshJabhU/BVfQTLVKc3ptHs
uDR83XF1H52GEqMROR5vu1B30SAPjtYKgtCwZiJP8NmbgMKe3Pyn3ucbOIMnmQx6
HSrWWHkK2oEczJT1JihuirBQESbI/03nY0RKbWY63Lke2Rv54E6lKRM4h0vt+fOs
m4Hfg+Wnke9XY6Bo9v2E4ud+RuajAgdMOOR2qPozsJh2svPfkwK7evF4fX/U6v74
aJD8XeXZlskVVzEGfT+i94XUkFmZrB1ByyXD01pSfGvLP0Hj383Z4fbJLgR1hlrs
r4ARNlUBMAOHjg5zd8sMReJzHnhbpXpIWfxx2Kvbf4TlknJuK9yLVcFsz21jMVBz
1jhlBFWwI3dd1OO+bq/+i6wUm4yEJsDh8FXiwm+6MTN71DwLcJcrqJMsQoVKnh4L
h9TXYRc1rzfW340UI0Y4Rgm8ZJ6U3DsdEct5UkqiRQykj22UUXU1e/aVCVDcIEjj
+DUbZFQmyZGIOpBLHzUMWdLoAwRpjJs0q6RppK2vLcYBpVK8J///qGvb76fOUQ/Q
sUoPJW/P04X4ebTx1YSgS8ZdWRpNkwJ6aSZ5tL2AUwdICr6xKETsLEBF0lFJXR3u
aiO0GOAA3Tyh3z3X7MebsUBgSCydFzNdu6GIrhJoM14Sv4w5hOP3zLU8S4VbeGTJ
cczZJ/wn9p5Z/K5tFNCeJdZZg/SnUqb95m13dw9JNauTrNeCLz6Xw6qmre0Pt9vG
KdVxyDN6BLwDpn8FN3ZOeyDmQdkICfzirDAK8Qhyvz+RBmQfy2rA8u3HOJRhqdDt
6sAqMDNbxtBEK9M7TP+XbEyu3GBDA4jqvBuS0X26/71CsyHyp4TW8NhWn20HW/xH
1dEB60GF9dhV4puJUwfg9sQEa6Cud6RLkilFoefg10VQ8BK1ESFr2nGT3vW/6IhT
lxVQZuh2eUJS1eIiDQhPzKmvs7whn0uGgTazG5ou9V0muh6T28fypnmBE0CWu6+K
O3Vel4/r6RnPCwHD6t5SzvYvtxzSPOx9Lk69YvDXRBF0/jHvwyaToHrYD3ny5Opx
webnGBkGSxs+HFNnvWLtlY3wk6fjRdsAFtDE9cDxJ6+48NJpN8lW57uNLZujdIa8
//ZyU1Hf6zVbj5rjKCAp5ilEuEUTfEhT5cIKiCkeSBXy+nMWUN/xVlV3NT2mIBAf
gbrpeC7Euux1iwoDJfLNFtxe3SEkfzaPdGhZP6Y7Sy2VohC7gEbKEkBy92ncz2xT
S6WPf45vRVMIDw7AWJCVJ+wpchFYwjyFLzOuoJyB8hCMl8+npKyLJm82LLWmkoSL
6Eu/Z1nKJUBCvXDbGSqcfkugDSCqCc8ZyKd2hVKrVcAaqRFoA3mByQP7ajZSnyAl
m3ZViLj6xXqPiUdcLvbk3tNdcMjMLTniDJ47GD/YMfSVkG/YdOkclvLN2GiUUKdW
cpIs2WrRk32Tv2lxIhX9ljIXmw340y8fZlnRolc2JQo4USZtRrXavYd2sN+ZfCxH
LAdbW6qxLY4+oVVUT+JmcPZAz0iBvjUfL1etfRqWs/mymHD9JMS0f3coDuHg9yno
ZHbzFXMVt9/K6QBxA6nL/GKwFLS4CCajMQ+2rYYJQD/va/7UDD8w6Rdgy8AATdcl
UZ0zzQJSc5uLzyQiysGSWH+5tAkb1PaMwFp8aGdvL7XpculClQrwXT0HSKcfg2yY
O8M6+L+MDrHBWx/QgoYKjEz94uS/aHskmho4HBVoNDeRzjFT7lQgWUFMDlIdjDZf
5Y5ka4fWe3iSwI1ikexVDNTsTJGwkfZAQqgXeTMOmW3WqaN8wQRLkLaHDHfp62qM
8vvACczZ0nnjHcp8rTaJneQcHlTkNbYM2tmlNrxMSd2qH+PJrrEyymv06I4KLa6Y
JcS/KpUC4YRIBsvHx0+rF/IpixuqnJ6lh6y5D1yyiJ8H+sOkG3MDLWxcuZgGCKZ1
QyZgMeuV8pF9ydpmF2KbgOgk0dcYQ1js7uMTI/KXYjrJRVBvvGf6O4Uuon9P6i4F
V+r4oI35Gm8tTHF0xRNwb4CQFVLTyNsFRLScrKE6LjWzNgf0Qh0kxAMsVvmrsZze
K5VkIoOQa0D2IEftaPSC5EiZMyB/x1yCWvPr0wxnGpaB8hQi6TjWCIRG0RnDER7i
kUKpME2R1Zv/jYS5DDR3ZQgxDmZrBkvsdD/Bc37D7+rhcYnYcn2jWtEWb1MaJp9m
snqPzvu93jBD21B203TPfQQNKnzevzn31o7rUttKzoK4R+skuEjLhpGpjIy9P8XP
uG5m7a113ms+gdGhn6F+99ApucaVLy2s2JIlN4gAPrlbDPi//PDCFMbDVaNtWj36
HcktRA1eGqpgYa5Ft9h4+f6Z8Ya0sxoTtkToq/mgMEaunovVvgwLLOSVIQ5CRFv7
wswoGJRmmYKN/keJZnHrLO0dVmd5ATleYxygaF5y9vkT1cP1YbEBd8Xh3L3C9wiO
p2DjoYwb88Ox72wGVg4fvmpsQoC3z60wT/vCGiEuOWbcWJbbQUZb2u97eCXt9jJV
ZSxb6Bu1wH+Kq4GCRV4BXZUwISURoMxOzSZ+tCahmGbJa/6KPxH7m/H3vg3+gnfe
eVjOb7cnuPELLvjPnwLQuq1r3vdqewv3PmyED/LI2i80flyyycS3v1ThHYQ3ed0+
+z3GWmtBebtMWPAqkaCmZKt/1ooQaicou7pY4hM9dIniUDiQ288sL+K1BstwvR6T
ADvXFCykmQzHzTpMfbmKJHVEaT/QzZq+v5rQbksTtF/SDMbXvCNpfNC+ygMqdzEv
RnwfYd1YmgtZuahs4PQZp6CndT+GERjzzspyrx1YM1WBWYIzBvzf4CcFMwRlroj8
Akz52I9wSe8ARkDhinZmxL5rpbyRTwudPzCPRNWZie+YdAgJLGCSsjIq5uChIowb
rANuwX0GwulJ7qoeOa12O6yXyKSHgLUvfOXRfQEn+LFI9LNRqQORVDQhnvF4sDns
PzHbP/milz7PSjOyempA3U7BSS2bm41G2gobWCJ2G7zuwFqUrRJ4bwvy17Jpiu9V
NHXbb0BAtvPY3FUsimqgZRRGRuqTQtjk/+iW9sNA0AjbKItVD19PJohqgh7JM5IZ
IAay9tciCH0/gWyBeshxaoDySl1OmwmuVlmppD0TKySXJ4bhTRbPFyTwYZdAxETW
zg68q1qelrh8Y6+ERZztlr2B52pi6jp3NiGd0UhTuSPsXyQNNLz5rFZpby8ehR1S
Q2so3OeJ3jT2alyfStGRzlAPqwnPzwX5Ms9Gr5hAHp66UBsYd1VL5TbbBf2cdCbY
/TSW/4giaqfOBf1VgXiSL31H4f2KrfL+pH/QgsrMCH6drkl1cL5B5feij+F4Dd8R
SQCHAHqGn8L/IwSpGcbZIHUXt+99Mz2pSg0AXiyjurArfrCvMGfkJQPzRxaK+Wcc
HSbIcbATeH/hkhA3W8L2VSWDNXTOJrNuMFL/ZJQZnMeqkgVii6EQEJuD/Uo5WnhM
yGIO7CL1g7Frjfac7d3dYwtG1rSB9NXaa9lvb2eoJNvIPoj1KrDSDp7z7uDOA7ad
wZzVEUKIlSZZ51ZHtPKPojFuaIKIqIVgH32emMKc44T0zfWdV2806srbYH/J3lmW
3e36ItNiiduR0v8IP9MW/pbn1tnTaYCVHkm52tt3GR4vGxRZxievPWe5IFqO/u2f
AgOitjHao1a9AC+GOuIrmSJi9AfYccwQmtxQp2MrLyC9kxsYTMnn4UtL25MiBRMM
IiH8qFOjdVMgvx4Uiy7ZdPVeIBa8m5Wi3DxDqh2DZvL2lK0KwlMvkMc468R0yMna
/HfjFNJ+MOciWyAbQODFpq+mNRnSbXBa/JBJfCxHBHnPYVTVIeLhafopCR1cuztH
mg69qlVsmQ8mygVnskHw1dZKDF+EmQyx5LprfavPtLvVjz72RGb+sSPog1ta37Sr
HKohi1+SZx1zQzXdCVxwYG8+o6KQbc7ZidwRQ7Ot93OeREquPZMMMUTyDs5akSTn
cXxgTK9wru3kMY7Gz5KQPBpsjGlXCR6YmWXKM9BQ/mHWYwdsB3m6ivH5OKIxdTeJ
b3AjgusLqekQk7N6Tch4znsthg5zUj2tXkEYyuI89DF62TezQRIvGsN+H98YUx24
SwXsiKLbEOnowEJaVXvqdONisvxV0i3VLOeiV9pz/rJ6ETBR9uS7HFn8hfXHWCio
u2Eieg8ezE60nlILwdpeiRBZFJtIWsAJ7wZXKntjS/maL9JIBSCYx6xkcslEKsTw
eYSU4VlF9aLsX8MVTnxQmBv0/8pfrcXAGKHCIjafxsR5L564JxxrEvRxYus57kUt
Yaqiq5WmlAzus3Ql8ZLF5buRTcqi3sy2UGLOLBHnP/DtNv9+9iEphyR+r941IXDV
Uckib3ufluR7hWLgR7uHzJpgRynurRmi7diyK5N/Agoti+Wg6RtHyJxT8EjDJlk1
LIPBpu9iZfNTtgK3UN0tk2RKhyQRHf6yq8sBeQL4HgvpyOUQhDuN3rECQTStOmn6
6U51tyw02odhorCQ+S/L8ExsHfOYC5hkIKGBJxw83OFaD9MwaZT+fn2jNUT3mmz9
/gryS9SWjEE0AQYnabJ++MwmfugxMkF78Q+b03Ahpm1dGpwj0uFfw51qvo8AA/2J
P9t+JtZCHNtWlWw48csFAf1/oah+ru8lm7iII8FDv+jyuz6VfoQSOuNOy8OXaatA
rPb8losLjtTDoimPnNpB0lk0SfzZs5DT/XDfCGvHaOmPncomsEB+GHYIpXL6hq0e
2EvOjMP7fx/vZR4vp5dipvllIwwMeUGKCs2Lm0wSlDMRrxo6dQMD5fyimmGoqme9
cg6l0hb8NHiB0y5iSafRijy8MDj+mJFH3RgCbj1aazgOLof+9oxVBsmNdo4/OFo4
GUtGDSMe9jP5b7x2ARJ93LWTipr2i2FtGW0nc/Kc7C1m4n5SAWiVZStQv9WzTe8N
cyNk/fYecCsJMiC3/p04kMBsaUpiIasiUKWt2LSR/44IRmWHQPlrSjFxJ94NgxU4
JjuCJ+sjFQ08PPBXG9/DDbhuLIm0MBgFa4YFYofoSqs7sZZZXWD4gP37iiGXXwtQ
Mcs160m4nKovIc2asZxBHC1CLP18nzeNomSZNACvmb4ODKJoSh+DycyMBZUi4EX7
2ogMwMiiU9da3qxtyslnnfArg3QoKjsFQjekq6ymBO02Xg03LFW7HIq1qdfL+laF
vlJE2xr2X27xrNCeFawdM6qtUWlWkYyW06eVeOHjU8DjhWg19gEj3xw8XxrH0jpC
lf1oZTCrRWGsDsvBfd4Wa0Mi4NdRZMq1Pn4LI6+1pNF+pGfF5ktBTOhjO39f61XX
5QuNfFugs+dxlJsXEsSrKFhgPhhTTH6CwhcWORC/7fdB9trYPEb7Q+nSbPJDKqpC
lXsL/8AoTNYHu+xXY6Ck5fMIs5cZwbITR8B24Quljlk28EpFdM+tNJAf0EbBNkm7
rHqNoNjF1SgrY6UkUSM1n9ncour8JAfkE29yJy4CmzeR4FSm5oVifYVJJlJoSoyP
hNj5keVCQlCavpnjeG48lEbY3NZKWzMg2FlYiIGGDGQBjMCU0jUgnhkNjOTYd+jx
qu3yVEV9NlLgFnUaEk2wvxIxnqPgSfcl1vDOYrncgxaiXEAnBdOLw2Xvcl4FglEv
Mm/jL7BrV1welaqAEwKi66W2E0ST4g+V/xmRZVdkXJEUdmzEydw0Qn5tmnBCt/eu
8YVJJD1l4x6RHKNc4xwWty48SOZGeHkgSwo9vNdnPPvGolXXCn1akC9vlMXwwxvV
ICl0OoOFJZfleoRF7QyqhXBRjcWGctlsVsQTKaMy7eA+to2N2G86MJPZVC+1pYqZ
vwmP2h+RK4umu4hDQFoFQ+f3muaTClHb8nVbJ+lvPFbSpPw4Bg/axlEH/JF1iJT7
QVGCh+yCMDwS4K5/O6R01n3o1IA/TrapVoJHeV/PMIINwNrWZWPm2X/RQPXBhEef
XPLh/QcX9LuHZewpIH79YmRvC60CEN3fHoHGRh1/277NkSM8pAIfEF1IgSm23Z0g
hmyf0DyeH5cqdkIexkZtNXNysP19OPiz2F76r193AG+uoQtrkYcb1mcfgz6IEcWV
kOFcxHwGbf2GlWyPlufJ25dW/+5jHl9Hid1Ntbet6NLtlhfQKqhRq8uAkLJdxPyG
nvrF4/9y+D34tCLFmhAXbpK5zv0F/dw/jTQQvFZs7/N/L9vm+gDqiYaxUFA2x4k1
OKwoG6jDIDbFjQE91VAntrQS9CRL4IJ4Ijl/OnAOwuiB9B9N7oh0s9VLxwKJgw6g
VAKXDyWR2kDMTb2+7dAP/HL6X45b1XSGCjf6KHHWM0LofR0qMcYyTK+VeMw8ZUE/
tt62jzU6I6Awq1eS9K3c4IXNk461DQZHoLUUe//jWe9YjGWl/s1HU49vLVjEHvgl
UwkMSJ/Z1+ZBeoqRolehxH85SvQJ/wpTLtkEdR6tsWFou48n7igU8qPw9TFjDbaV
DIaXE37xbz8VVWcH98YFRkLuwDm2lIL20gYNXu5X5CJQqY+qYUkPrBMBYumgqmYi
ha4P9LUGl2gsb9AfrhvaKzlrhLj8x9nGO4QqgxiXxptTnTP9fSmUhUILB/FZsT3v
TNvRLBQxIMsQDVtp8X8m1t9e1flrGsG/9d1ijdVJnapygsXrK5ltB0mqx8+yj/H4
T5X1wtFpE66OHlCkoyF9TomWcGzAg/2s7Dp7Ub29Y5ZN28J0Wfg6fB8OrkgXTCjU
1myGygpyFsK3pmoyNw+wGnvDs4bV+kpuCWDrS4n9U6iTOQMWXg0jRbK7U18vwUCU
Gk8n+oxldAOjlRPLqEjWnktXuLgJms70mZlX4aB53YcwHrcaL9tmGVqbfvpLETnY
GBdqyA002wkW+cwly/vCG4Iki0sOKOY89OwuFb7Q0YQ+FVz1/YopZA/2sv6G5AtZ
rD3XS3so3hj6Lm/pw0DW2A0VOk5KFrQHitgjvoBKBsBtt04g5pZX61SMbYXC/jZz
UpjFwl7i50JufDBmmM4z+HL08iOw/dYMpvR3yMnFlTj1maL3u+Jcpu4LZcsrEKks
QU6hN2X90xT+dbeiQYvdIYYuKUylMNTe13NgdTMRjX7UR+UuE6JLMntGc3XF5WiF
uQfNy1HwiNdw9Su8LrXibkRZvuHj6ETrx8DFYmxtF9IKfQLBdnIBz2BvMF6+iFOb
eP5msjj9Wh1yvpwSE/NK0HaX3RP3vJeKJPZ7xRlLaW6UJwuMKV2PLiacd+SwIbSX
0PgAzCt/OGBh7XiJRkZorYgmlPbbz9BdjbIjlb3pyrtHG4f6BTKmxvmPvqcJoQ0A
Gs+hB6NPnMvd2qMXk8qS3FFrdwEdDe0hIAsme3lB1iQtlL5WW9cUv4Mwc/kEx5pR
sbr19mnqRDD6VanpmweaP7aHHgXrVvy4dfPnLsqqgxzF9Om699uSVVWg5+GoScgu
PU3Rpu6WgSLb4L7G4FkIjnFzMd9tifES/9rvbggl8rMF50C/59uWSBmHmgrkrFft
9E9o+IF5VrCfBWaJY1MrkcVvN1LtzsDyQy2XMnrVsHoIknvkJInihQ71FMYct9sw
lLAXO4242ee6PhB4uotcbzv1ucWM4w/ovIg6pep3PThpSvHmDrx8/3qvXcZ/+Jvr
17jjoWJ/zdCipQ2lOuz7pji+y0iQSp69yZZC3MX5ED9aDpG24bEoAagzhfrprjVc
zkwi8lPBekvHPcFD7LYBOVvnZZF1bmcxG6BrBgQyAkAC+6ZOhuNE8pIHSKt9hK86
IL+YMdCM948uERxCEXeLh3Z9h3EOcyFAQtFUhEPA5jaSyVCE6v0ETq3hlm/k+i1w
8kvCMXZ8XvOfzAwb9J4oYsvrHQk7HuyuwzEYW/9BW7rjW4m4Iad8V9x7Wwq0GwuN
sm60amHoWaA0TXzU4WvSYWAY9zRsTdqnL6/iZ5bomBtvThxhoL58HI9P2a+U0xZw
M5f3CVPj+Sg4rAdAok7FFVz4fBWP7776Nq8cw6pp77Ivji0kwiE4BNYgMjFCzTVD
fkthjfzxkk459NsY3fiPfZB52V3KEq7ENaRMNcmV7qKvDOcAr2Kw0gEHrr44Hn3U
YD92hSymA9TyWDypmHDYJTjDbvrf1A1QuE2qDhSGNwk0/3v72GMJ8srcZTL3bpwe
JOETNReWiN2NF97ldBf68zEngRT0pUnsCEmwZJk2zYBbrRhqlzgB0Xbs0J1lQ5e3
2RyreP4JHXC5uiS3l3Um/+cCTXoSwTh0NfGpZbgvy/kTd7jZzjqNsoucC+6Mjbhn
zjAd1F3vX3vAD6JocLyBPpIfrDjxDPEvglNHgWEbHgtGlBCKGP54wDTuwdaky5c2
lNVKowxYOlZjWHTyKpdNtVK0CZKIwd7jsuYghR/khVyAzV8qb21KAG9hc47CGdbW
68/4RqO4/TkYHm/xRc9NifmwdoJleORRsGDg0GLUqHEl9tDpvvbnG0+XJto9GsFD
S1mPH3U/V7RtDtLTEZlOBK7ryUluyD1OXyTMbkmL51CVOgXISn1AILLGEyHBp1zS
y0E2l+mmWyxRwvXHsVwc68LXJYKQgSpi5UnIsfWGAPkjZYs+LoDRgyqO1Ah5oXXG
mhLKBiDJy+G0zajbYE+oLe67UQPk085bPLEUTY9twSVvtwE541rvy72Bn1m9pauy
rIjuEFNnfjFKtef9RUIBjDl6c59PdnQBZb1+0rNrugoSBw3IFNgbWgdd5e9PC9nj
nrvgB2UxnmB9mUSRUVpcrWawRtgc1S6TeapwAl0Rds9pmtNKV28y71KswdVjEyLl
I6LpFHwijINVa/VOoT8tdOr2xhAmqXNyTjDhepeNkbdEIqO6gz1/IMEWVrugzN8H
Jx8jAxRDtOEdCJ3VZg3cz4ZFDIYxeH81sxE2Tuoo68abvmDYtitkJI8aeBARH5jD
kr8EliuAl/gi+qwQ0bbrWkPp+c4vcS0KKa4NKxRGWQuzxIerhzmEQFdpzMG2mSuM
Iu5ycGJVhfp2q1RhqVxe3wuLhM8tE1S3MBfKCZgRFMgBsmMashEqiMsUSxYi5lM5
0pinS5Imzv63WV8VvnVyImXcyj875PMHG4kA2LmGE7w4tD9UWXeWIdiYFK3BLL3M
rmn+UV9QOaMSrcxEHKUv9YrPAixLdGEUCZujWYmRvdDeWq5eY58zuj7i0hTIIOyq
oV/4nbvJmIS0BdA6o8dDpv0uPlOkiVSO2L3Q2VbSe/vYKiX8YQM81iU8+XaoD+bv
u5SdHBSSDZK9vMq+lcbaI5dPoCQPtnpUv+yR+ab+Tg5+L4H8JnsrPamfFYtbsGvO
HPvhcBGPteTk78MB1nLJFUIWgt6767aQ6BQX/TxdqZjMiyJ+xS3G/GZg6Pew1sqL
KRnoSjqN4sp5DNnoMc+Gb9C+TOHZgVRnFdgT1CDKEzTP+uFKmSqT0PNZjNUuS6Kv
jW5AamKTE+7JhGR2W2Vug8LHJ2LApQZIDaxPYyQVDAIWFXGB8hMnmkpce1UF5bgr
fGGPcfdsx/eZcTvqGojia9wxgnWvg0zs6o1kXXChv1sK/PEnFZjfwhTgqTrTulXX
ZUb0UZY4wmvPnJBkLcG23XJYn+Slmuy5qKGhl9KAygEcCTLOIrloLHYosM4l2got
9umi+oiVsqUehwI3lK8ouV4SK8npCAY+MozLzFF7t5b9h9BdhtMPevtF7M38Unu0
Nk8ENGCOwcHbqjgIgWgQIe8zIsFFqOoS9jdWclVCrNNSIV1cIKvvEj1teXpzfjq2
GS6D6TrjOGp8BC7/e3o96rObZBs0/QWSjY+rGpy+BwF7/rB7v22uewkiAuQzcVlr
oaI2vyqfxzkLWP/hCtBjcny7qeJCrrEJ65qWiN7tGO8lzZodSma5iRRlHRfgtYVk
G3ce96j9X+yRlpBk/zp/IGqiqE4C9/3gEKX9qp1BjOd5x0xqnhGiys5OwRxp1rNi
r96oG7RUjy3LPmT3Tozs3VMeQ9ZZq/4AWj1bqsJoEpxLBQUhcpIO8snvIcTltn5Z
a79bmpi4NwRLLinyqrqK/lSDBEzp6pq7CouuA0J+5jFsheU+ScCaQ3zxdY4OEtq4
PTi1S7utgpcu0spw+su1kgt4dfCu33WvoINUiVuYZ1FPsomM+dZNjQaSUu9144eA
UC+ngo5wDV5Y3/oxp0klNMs+ZPz4aU4ceFW+L5RbOT4oHMWne4WtwmKjG/v7axad
Ona5PAoFuXGKmATDJj6bvJLKOyECSVEcV2x4B6BxEQPRalreIlhVgJ19ZjTYdsaD
u2WxlQ//DckRXMXPD2+xzmx5cSDufNmAaDPvD+4Mpn7QUqnMv8IOtAX6XpxdewhI
vCdq/Nz9gfYH6WQkreS+J3CQTBQc3yoQj3Zh+t2FNI2dNJd3Vhw5tH8pJ++6tn65
2DrBWZ3ruY63FQZAnRn/27bJb2KYiw/MhZXqzo7b187Y58lgM0lscs3aGCPgszUu
xX97PCM+mJ/fXQ/wcB6AjN2UaS8y3YEdMBgeFVffmyLxVH3ys9hhg5GZc2WhL9zj
C18wbHGOD/wbKS6DuVcNhLwfg4KxcOGS66Fmub6gJB81QJtS19Ddvz0UdAZRTEb/
CMcJxtTXkUXqxhN3U9AFe3RkKvm2ajodQJzRfNPjZKQmN2mWwA4nuJSPnUIVmQVa
4nSFjSnKfTN3v7iEDUypyuAbfjTgyTNaPxUgGTaP7y1BAnOlvz0U8Fbpy1xPD7/H
7sFnaFwRtyLrM3AQfI6FUj9B6qXtl4SB24ym1B7UAe3QrYC6T7F7gX6u/d0fHFkM
mhJtXp4c9DlI03mdEvyA0W1CkwsjDU0pyfI3gq0MyodL31rVz+sAjXr6r3QVDa0Y
nRY5y9vIeduOWXG0oBDXKV1rSwBuJ+ZHqg++2yNKmTN7fIQ/JXQCNjG3Biqs7w5L
83wNW0V5nkla0t8Z5eKpV8d2v51GXkn3C2KDPETG0npUvJb4oHKzvhVJmMrqjWqd
h0wlVzNhR8OAR9jsbgXTg5uzmGFr9W9uB9kyGglPiCxtT7kvwlKH5KqlNi84Razi
tbg9klWRlOHRyT5Mqv1lKa3GYfe3qSzfYkG2FuWa8rSooAyEbKxemQn8lHYwcz9o
T0b8VvrZ+j/L+mq4O7drmbHNh6VNSedGpB7C63mcNKLS0g5FcrOj1Q40kWkjADMd
tkUFPG/LhPn9tqpjNXD7mosDtQ7hzHpssw3/tRCyxsUhlEW+CV3nSbXsU2GtdYJJ
Y5IKwAulGM4x9c0wvdNtnvDX8dtNRRc4rJUKyTH5M4S9GVqaWiXHKkrdFsPm15Td
Owy5SdS+j+nDdJ532i+d7mPizzOHdCmV8fmVGhdULD12hTrphN+NwRlqXHaemcrg
8Efan16nvsLFLaJbWYCTKf8iaZxn5OHWaY5uP19UisY+TKKLfBeIaGCLjIAC11vH
xuS6IXGs3wYQqqn85PhQtk7LdvNO4sh6E8CUOdQVIooln9DSEY2/e8/dt5xVGoDO
COszP5lMrmul+WCODoxY0MFObrWxe4IkJDRPaegNvju7xdmP443VV2feH9+VGEk6
jksj1vYrRGSDk3IFJBvrGrEzFVn6L+FBZBXhke4lS2r/YpCJHNfOaFub93IJTc02
ZCXkPGgKsAA7TvJxQdHWC7NIeSvsOZ6ql5C+KAf3Ie836xnH+VmCGhs6frML0C9r
Fh3/v9qSOjNCUdTYw9s6TAFEj7BbjdOVgTEesIU0eNk/qR1VlSswsiFm6VKqPG3G
3tSPIgPKYlBqAss8zKNxHhlx7okzUgQAcJtsXJxPQ7Idylk3W2IhDXTsngBC2+xS
Wpd/LIY0RhxL7c6azxIlwghKJ52r6+eurU9kMO+UgYY8VkKW08rA/RZ/iKxPtM2h
PjW+Axcdh986N2MxIwVYlKM60FRVy2NFVQWtz1WC/xD3WYuz9ndYcZZBxYW+FBos
JrMkbEjNZSZ91IvZLG2Eyl3zPc8Y4TkPDAssby4Azya50N64J4wZ4RXM7F7MpFFB
562RML751ye0Ql2/bYRkFk7unA4kEul9w+TrBYYJ8A4kGOGIKgDiONBImT51nhtW
bmgW4AJgWEHCVHZL3W5hIKERBCR608XL4UgoIRtsypQrj8e34wKONNGhs9AnDpBR
PcsQ7kxIn77HROCXz52gD64JGGus1QKe44kl+9aw2Np2kdNfFQQFDW/rTztHEJFM
mpTUezJWktJYBLspVMjXm5LMRHqiCmiBFaGcvBvQFvRtEsAsVeZapk5n/87jLZDN
YVSZWaa/cBVrODb2nGGcI7kzXHHx5Bm5nQpIWxfbb4WSiJbzBKyVF3DFqcUPQ2+0
XLBmfpDuIOnU2gt+U4F0UaaLTD7iSI7FA2glC2df/0t9aUn/qKje5tuzsEmyMl9n
RV0oOqUCSjBRg3gdtSxn/qKpR5EF8alQli5KdCK3OAhGrxtU+2GAXG8mdKYvDgsW
U1xt1C4uXCS79xtQ/qMsa8qSYfSJXW8jL5aVCHV/L6KG9BQZ8Zg1nasSmCelFu9R
Rmrt4/qBEkuVUNy18f9MniIYGVe7sF4VpdewNdFbPZ6yCBaDhYpU7svnfWKk9Pav
oGNQttZ0ks2G8I4+h86IPpDWXN5t2JXu8IHgawq8OLQLHzw6WJQGSrLmhoLCsDMp
TlEI1e4yLsF6KzxMS8Bv0Q9X2gPJRTvtq6vcu3B69b6f86Mk8TYpS1lTOTwgRMYt
sc0gA9F6oT9EjVGjLIuV+PM2UuekE6+rikzLwVt1ByBXgGB+iUqpoFlFviSDnm/I
bsPKwJMqKSaebA7JWP1XPgLmj2Wvttc+hfEbFqy2xsmNRYDzugBCOxk8PfNry12R
jT/rWOu/N5lnmwk7qRvho3H//GV5ZDkRwhj3AE32Ng+3yB/ePyZNlbKJdoVeQutm
gO2h9YLzxvcJICgvqBEpViKPvW9zvlu153MEj6YFhWxdDt30Ri45hQzfcfSNvfd3
y8hYp7l/wXOG7ZaotDgKAC4vSJ09u290LnNFGI3mpRGuDiz4xVXuWVfJELSy6Fk/
kUBnZTukK1TsYziDb6q/HwJ2FvEeVelz/niPNvvgqC0EpQvkBDKQFcxE5v7ZgPB2
nAuRuNG5Mg7hQoBR2QC7vfesippfc8Fnv2gvd1V7d2ZzTslxMaeVDWDrY84rO4n2
kb5h4YMkxA8jgK+d8IO5u7o6EIlPb4KNkvWzoxR01PHf1iiy1mkRiynDEAT91H3c
vX9QibIqaLLZnk7Shlf3Xw7IQNp+Vvq/0ErRT1G6zgk9lonqCcAIAAx0PhS1iXO0
Hmt0mt6rDgKG1Hzz77OPL7m8FfGU1+f0J2tHiA9fPyTBRcjuHKjAjLEQWBlb1Pbj
o7NEmSo4/g4JUA1FW2is8aISILwnAT33CXRvFN5VDuecEu2bqHarNoVsCS1lvQP4
/dfoZUZ+fg9lhTDoKGnWZFGVq14rLOLswKk1kk8jrZ+nQZZm9BeTPrar5ykoVwBq
TJVFOTmBE+f9sQ5YYexYgpatEgN5eFkyrBC4qPmODpUgMubtT8nx3zNMKSu9DWs6
LPHpu4Qd0MVZUSoosWH+zJMOeqMGwHFDrDO0YzzJH1rjuJ/fP/PaCTum8PGHmXOz
H9HMYVbkRGUGkhibClbOL0RMxXtZb9D99rzg0ErpXISJfQ0wBKDjl334NsQSXgyA
pin88hWvqxp3BtDdFJJmpKLvglEel940WOcPqVLciI00lAm8WQVRLUz0h69HMr4L
oXWzG4rWOPDg+exwzLpHw14r7m3ODCzLhiFiBWl4BjNDT1kKY6LfC97FLLlqALfZ
60bnhX1oWIIFOPmDlzTypZ1F1Zj+MjjHE44SNAvqA3JDX7F0WFONhGDTGPG+2W8P
7AYueYUKKDovFw7tnuauQX/ksuRObaqSK3tiCN9tLufJTE019OgCHVf8FmKax0se
bolHwjE8vqUbzfMDCMDmXW5G96nGITT0DdZoF3nVBVNzi1e9VxJ9JP0yrxcJNCje
BAoE04gKzcKBGQ7bteVnq/e9PVYBsUDcFZoGYE+hzTYSC0rclEyjMnzT/LJ2pp14
g2JhpxHdNaGS7cJzm8JrpN/9EbbMBMvkxBCSTpDG1xbB+msRivPd8X8GbzjPJZtn
84peYVmcApsMHZ5i3j9vBbk/zX9lFKc4lK+qpIbKVGxV+iRJBodJ+nm6ZK/VJ/UV
3eDIMPd3ye9Gp8dL9uqfUiH3h9ry6Hl1R2CWoZSf+paRJsbabRkXjXvDco+01Ww9
rw+B3OHArErNPFUBt8RkP5PWC6qFUnHQWWPp1kEKBy8sjZBSFQwhn0dh5OV5qXPN
ebPFvEGnjnhl4UTi5NJjV2EcFoEfU+XAfyWGzRuntkjEOZS4O4dsdKNwxbNfvM7h
bZE7W9uDYlH9KuxsWoMOxym+869Ak1BrJ0/jrSUzIBWrEGAu6xNkWdjc4ZfrYI9W
hjmZRDPF7AjKqWFgmOeCLoNdJ8fopq1YOoizWjX8BJmln5509nj49Q0F7zqDeBvk
QBVVMeFMDMZvAJSqq3hQ56+dsGNtKvje2e7amg4VVgtnzUYl7pegzZJqaIVhX96q
nmUWhMMHGGNC8PF/dnvYCkpfhPIRJUL2+9juY7QbKZO/iaXL+csRYo4eckvMHS+4
27pLOSBf7uFnWBdnctKszO0YG5MBgwNlrTAgqJCEf8eMAFk2woDdoYIQfKShZ9go
PXBIor7D9lPPeJ2px2sHtlzveA8TO7x7sMl65QpaULDwXp8X+0lcSJIWt5XOgl2o
w1tOf1/NoyIRKUfd4/k1dpOP86e6oP/8043949xIyOjuKbnePx4cTBv22vAmpAfd
Hrx+4MxYMz+jHzlzssQhTUfx6PyC+5124D2DDrihwvIZCcs1fWA3NqAl5aks7Ooh
/Dy6BosDHsoISfPYmK10eFO93/lLgRclXMeh+EDw4lc9srdMZxBALCEdeolERMqq
vcCt2sFfUa+yy6WNglFgqIE6cj+a0hr1sjzZhLHYWu4WwgeCPcjGIJgjK6uJPG68
wK9+MoB3CgnKvMeYzDpir9H1GLIg68ASf2CkmgYZgMUXhzfkB4K5hvImUDKs7jh7
+j1fQi8E1GJE2NKxfcM4wERFcIwn46ptZTLVeSqCJdYdSjRLZAXU6oEoCSlVD+jK
y//Jd4KNomukXWB0U/Nlue2UeX0l/9WF5jH9WTOAXWySCYoma7oJC8oD5qNWshJZ
ajX1Zh4PwtOJD/7nwm6ATulnqV+/IjYIa0QPA+96cZM0zu69GnJG9n/wjIRvNRn6
q5upYmloKu7cHAfRjRoeQCTOzuW4Wuek2BcWbmMs1VhbozfIR3se5auW9RHdYf2P
FIRa3uJ0y96zEqQEAtGk7uO+sxZ69rKwsJaa56kk6QLvUAGTI7b+b3lTu4WAH3Dr
W+Y6OCkf9xqwjGFmnDBajET8B0/FJwX7tLzZEmFdrHgRgQUICy+WLE/Iy8ZIBsD0
bmaoGrT+9YyOM3VD7SVk8D1OLxDf1Y1mvjxWOogT6ixd5fkJmx4indnE1POFM/5f
tGPi0xrPjY1gW8a1tM3PSzrmaOAHYAboD7czAy81N78mGWrH41UyfGxqK/SCqZ94
goG0p0iKJG9aIIX4i3v5EuNDpGs3uksVYXXolRFBJFJ8y/vVX2xpLRLxzPqyo/VQ
8cEV37V1Gm3CF7gJD8xotuRsj3qq0v9UcFAFjLUjMBVbVluMKEiKiAj3bzyAC30F
GjE9HtjxgfcuF4hYgmQADvM/XbtBEjonRxtIehfHlcpYnlsPMJkjEml2awLTi+rs
j1uHwwCRB08bWvr7ziDbfKMz9tJh0oRwue23HeGoesMO/cvlZbkET78GY7W4HXSm
8hAIfifbB8VMPABDa3FR3B3qobGulnIqCaCF8ZrXAcH7IS/6xutJ2QdXEMOC3Jkq
ThPQpfx6u0CiiJ1S903q225DqxufkzEJ3NOpXfimAVzUm7Iqa84sPPBvF7gDdb5I
VuGxhO+SoEZ/xFmhQ/Bs5a0WERxD0lqGBPeZzBTn3k5klrdrnMGC0f2SXFnJppMO
N5Dfl5MhddZ+yW2WInX00WIgGt5FrevqWBXdWD97hYSo8MEQbT/QnJRtjUyjZlX9
/kpeUiP4ALYV4/cXqwGcDDjsRHSGb5tHQ33U+jZ3iFSagH4vqzjMPa+zGFzqEOLg
9I2unmnBHcQ1KoG5LJ1Ks4heoIeKMeH18hHfYTK77aE4t26BGDEamlsEejHMZK6Q
eIumt49YUtI3dxjBiuZK8ZVAF8QgrG2Nx3LsuEIxGKOCb7G56ZDJibr1uPWL0OGE
ypNnMew2lgoHxG+3HVyLytI9qyrFexc4Rldn9K504KcZiznQSIPyulMIk7C8MWdB
keqzm58bjoUb8mo16OVGWvTDZN9o5U/oK5C3wIVGE0k75OI+9G6CVevHV5TL87hH
h1xhqdVPn6PHJAFBfC7XqUQkXdBwczdZZtkvnBCTyt41HIAqNdHy8jZLHb8DmPJQ
d3hDKZXtWRRbY6d+z0oNTwxDbHaI00ssTTTVKgYSUIaLWxYjTCq4u8jUHgEPmIUc
HYT9xyLDU//dQEEnsAq95kq7gEZsgy0efyW9GBLoqbkqSdyLHSjlTOhAeH0MA22Z
t30NWglMfXlhTNG6SRTlYBOPlkRUlxCYSrXDMvM0AzhttmTox97HNEdUM5e036/h
+XpwcCkZIHJ2anMqjNANy17mej+0oxfVH+gFrGrINJ+1d7SSGqx/szDPk5BsS9rX
pwnm43rykbSmsjc6+8fE4YcYbMnlRfQk6x2EvssPZjfYeFWggiKdnocsMK3hdpWO
OdGBo8omhbxzkq7yLSgD10hxtGdoYQ2p+jVXNLVxcxd2TAoca+NXceMMT+5me5hJ
u+M0I4YXsXgI8cR8/LRWhgd+EFuCL6HAAOD68islpndd7mGk9Ge+y2XYke55tAa3
+f1+D0KH10W1aXRlLec7pE9OV3SVux4DxLeymtGZjgvXEFCqoiviLm0eiLKhluo0
C797J2zbIA9CaNDr/qjI3IDoLYpKhBOdCOcJSEeTlyzSSjaUrtfr3lBY0MJM8pnk
xlWD+xQyQ/X74LJsTu/TxYUqnG5Cc/YI2p/YBOPZE8Ex+OGnZ9nDpEO/9/dqgTNB
Um48swh8KycfEvr/JEXVs7eAvs3Y8YjIjB3aXheBvU+f4oXsb5HgT8tjhN75vqBY
FHPivHso9osbKtoOJIkJZONIdCzwfeR+7Oun/GXORqKRSQp8X0Zddi2QeXMpM03f
2sYlOi/9/q9G6eeX5eKhgd/NhxgHMnGbIpCnPe4thwAhvu9rwrbh+pZM6WyS40hy
ZLfg0KJlMQ/lpiUqVfYKOGns79lZB/B5E0W379QaeVu5lD3keqa5gwEwAyS7qGis
E19I9ToeXh/utNrd2EkS7y8yBlPkhZFyfa+wgGQxy805qiGsSDJqO88ut6I/VX0g
/QeUhPQ44sXvznLVCeR13Gj4I3PIMdanhaW6u4/N1WY95vcvPZXpVH/GO6Xscc+X
s9TeuKcT0b/OlOBXcoj/LIAkz/J6MTfc8TBtXYW07z+kiuECaxTUeHV0QOOlJ6G5
Y+Gbx2IR+zGMNjTPLZVJTGAEHGZElrTHCFJ5LnbpvBHQEM5j2Pzk70l8nHGbZ9m0
Xv3q58yokyxwz6gb1PAm+/uptBw+BJlfGbIjFM+qxDrIc+9RV+y/EsskyJyEASDC
RTOEI1CVoKaXi4WWjx2yVGYpgor4JoU/CEHC74xTdDkHhAdg/R2NbGoDjo01XV3N
Pg0pntFlBhnzv1gwAZ4s9TYQEaw5xZUTJ+cdBtfICrc9LWmgjAnfxmAPcdMIi+W1
qxpedJGTOhMNyjKzFvBAR8Y/tYZ8uTS8Wb6H8mhJMnXpdLBDJUfhmem4Z1ED5ymh
VVINWwHOUz5q3IZ+ccLqYe6X5uXs+hzixOYqNNbsaxr6Ugzx+2+GRDSACpjirLhj
fLojKuMPY1S+4yjrI2wmy+dmGJXgxEeQD4AOtl4ul05bks69Q3MUqZLkAWLn6xXe
+dRWNO2/xEECzdFhvA/QVQtJb2D0xM5EeIdjnCwuxzSyzOeReclt1tSg7T7e3EXA
xl1/bFWs0+HgF3kkfHTP9M3tMlrsTACA4YTW5Ve7FDE2uZIYzBDmf3riB/5yp5Em
R1o+/UhzdpeQXW8dgIJxn4FIHsiZJ+SAkh0a4rzcvUJOc/hhgW4t3uzO7rOFf8tw
3Rs3WkKoGXuEAFqwPN774nE8IZBqkMq9Gle10PgAZFqVFDbCchddsiLNd0PO1AGS
PZj6G+diD1KAeUzHz1uy33ZaWVbqksoLljyLfCOZMNrN1fPvU7vJ51+L8VBpKOxt
83LUMQV0d29Ig7JRmjsdPDHBTW5ve9BgtLHOl4tsmJvomEbYHDpDDZBbZh4Q1eRg
0yfDv6iKl3ihwKjsksUnMIzL6RTTzYacsvaX1ZqYt/kp04w2RAeiOfgOOVRHBDOU
SLba25VdPHj3SCCkwJlAMQa4q0oVVvM0PIulUbO0bOK/G02d2bbotmxCoHgrZtBH
okM2EW8y+f8y9L8Qibm99rVkl6hMWG1jFvmSsuk1GVdPxChEuAMwjLd0PpRQoKAR
iUuoP5895LYRZKu+BCgCgqZ1Ht8RLvutPSbT7OaxW+6XbDXOJyomvpm6yHTg00na
+XjjmYJB6ErKB8gRdHO90eytZr5OMaAuR67FbColV5eWYVL4U21L0J80ZxkzPS3e
uzQyI0/TjJndFGM/Soz4vYgjJY0Vyfg6YOZVGKZwpe5QuFzLxCJdIrhDLcbHo+Un
TotJr+T4LXq9avj5GSukVyr3uLQYKbpfoECwzMSsCFA4UKUru1aZBDWDOqvPtD9o
qDDpgtMKA+psJmtkIUXpnphiwnL9sL9eOuUWuErb5pG/YXI1ZcJKs8zmIv74FRa1
gpKARjrf9bzd0Gq4rbPS/hRG92zJ67GiylZoTtd6gLtcrqJuer5wvWs0ohHziKgh
LZCE4zDoWgwTNh90jUern4jAZs55lJ3gnTi3f9MTJxS+w1ltIzXD0VodkqpL6GjZ
kv2o5A9LHvj0IeRCpiopL98ZkfyAWzxIIp/u5HB9Rr1xGKLYEhaL6YM4LeJfB1jJ
ttVYMde1Wt/cWgq5f2QjqMavkOxzK0Pve821xaLdSW5HfkMQI4Xz4tOmtLp7ZHUq
kC7RAAiXxYUNNYipgCZt2T5T3boDC42Rg5NcX3ZCfQaYaKzBe3yMOTxiJvQs0mqS
TM6EKMuQx3fd9H0e3+HlmAO+fnqSoESHYFWy2KW/4bF2nGiqFvcCf5AFYVhHUpkI
HTQIlClNyQXUzAjLk+vqX/8GkbZl+LFipzIAFbN22uapRhNE5iBhnxJsG3u99eOo
SZ9B1bSmudTDbyvkUhFhjCr8RzPlFfYL7/nl3RCYDEOS5COG6SgIbVf+IjKQRRDv
6vcdLDbNLRgt7N/4DtBqdInHbO7kYLVzMs0hCTTphuSYEWyZBcMTvpG3vk9dDtkG
F+I3HaGl2H6q+JLhEBG8HKEvuSP0Vc1vCytRaDzVbx2MV2PP0lt5itku2lHo3mCs
0n5zFjyndLIBX1W2N88beugMfg0QIEU7/RwR20Ck4RrcRVQMXUSVbEf5PPquj0o7
tmFMVFzmIATXMOPm19VKp2vAwXyPvNtgUSlMRjHcy16wdp2ALGUA1PJ/5UtQex+w
5LYRSYv4pkKxFzta/2fV8AHyIoG5kHAWQn6g40uzJW9zxlvvhQbzMdsdBV9yTaxI
WmqC1zNfETXrV+xEGjK0eld9uEgcyyI1s3vLESpfE9DDtiFCTz18yiaEYV26hbJZ
HYYjyFyRRAcZ8u2Sii5Sxryb5kXr1M7jo/B/y9bIpvlemXPAHGcWKImfI8hSeche
PZDd2TrLR14xtnMKuRPbnOFagFGDepHOGIcSQ7xsuZb6+w5DCOfHPWVGy+yKv2Jr
sPI/xDCECRzt/x4VLVLiaNb6CizXcZNq1gHxQVp79tINGdNf15Jt16DZu1a0GEw8
/z6HZlohJuFDK4LbBrGKAFCU2uEKFMstVUhssv7GGEJ7kUFtbA71k7FiZJilRj7q
S7A8NGueyyT2bCN71MGh7HeBrSGmbrjhvDxTc6i/f0R2AW1V6HpnxWlu+nyk5PzC
luHOb/IbwsxQb5MgEVvsijJq9i4WEtjLvhT9ckNc5Y6Qg5STCjdPAcNTRYs7A9Qa
fmjp1Hr5B02t8nfc1JF+0Fz/Ljg+EbZDTFowic+/G6W3x5wHqRV1DOs9KOWPJJkf
kttmA430l6OfAV/fW3epU4C90KM+DTNhPox+o+ssNghg4Hhw2X1ki4fMlzM8cXfT
WS5y2+fOjHnngwF4gc+SVGRfmgEejSTDXGKT/QvCgKm9MdAlAoSHdM5ktZKLN1dD
6DElB8Hc3Mj1GIbi+5fvwakLoCsjZQnaQEl1SJy94WYBnX4E2bQBdwGRT8EM0IWW
ig70k0ni2WCnrqCOSBBweSNBp6CFNH7J2qwdt7Wc1JdqsVHu5nI0tWkbWGldgCnZ
BcCAfClxEmGiR3upnKLhS+JK7Uh1HxGkDH0XwdooVbpJiZZES9vc2jMb2tfkVeJ8
R9HfPvcQu6R7PZUbIvkZ6GRqAy8/xK5/cEKW1x2WM7ez+Gl7Mr5s3MWvSX77iYUt
fXlx01EC8YMagfqHJAeCejEQClXQdTHZH+dzwrF/VxlmErKTMwvmqhec8oovazty
PKi8DQZuoCh0r3+n7lbZPxOo/IogLCf0jYWvTuSxsl7ijQGthYmWvMxP+ZYAYHwS
4ox32E5DlbKmiyu/Tk8s4VO2hv030C/3Xi/2XaVH5w6x7Bb9dUpcPA+UJvm9ZwvI
8IX+nbYlFINIs3jCYdAUfRAiaIqAir7BlZnL/XoQuMjvV+E0zylH864haFYyT5RN
JopC5DnU2WxaOi7TbVI9Q2Vcxys9afEgvxYx4VebAZWsZO5FIMH5J3GUl2g4uqEt
ufeaLDcHY42ZkdtTo2pLDbKRMAucevsV6LWltpW37jzbv+r7eWuktBVfxI044cMK
IAmX5L/WLM8plU2BGEloFttASWX+FN6zrARSnP2L9UiDnQG/ulR5BVCwyrh8kR/y
y1ihUquiwR23QT+mY89t3AI77FBvUksHYAVOmjPF73TSDlfr7Kw3SrK7gQidhY9p
LPhKn+31uG6w08BQJaj6iWSEZ+BD7LezKeye54aLEaqXFBDu47gOm9I28dVhMed5
+85wVykyCdF68F2riVglxal/7yDRKqSo0KRo+rdIDF8zH/j/5zElQMLM9viynF7O
WR/BMbRcKuparFasRswCKRsORdo/dSOzg050h4MU6FufXbVeTniMMqs5c8x+hlrx
M+94iM3HJzGBPgqpuDTkBCYW4GW6j7LA6YyaIy6c3tJk0Hho5H1fAFi6BAtD46Xu
08ivwXFCQpI4QWm7C4C02cUEPtp6x8Nw1ese3sIMcOHa7gwAc+757VbFZnIcUF1U
H5Q5LOIP5iL5EgqNjm53kWUclIGbqT8p9pdC8MxAyTXH3yGS05+K0nVMyUuJxzr7
yARSewlYBHJX2IEXYNrEbQbbzYZZXVI0qEOQmCWPUz85kHKFnXIUEYEcatcu5j/i
yx3kiJe7cV+opy5KLYUUp6jimOq49IJAcmDMRoux9OEzyyHwnA3caduY/azMkVEA
Jes2zmi90iCtI7YriXDPMFeyhQ6GugxjlQMk4zCuHcu3CEiNiqYt1/dmfQxc+zyt
P8cKG8pumYfEd+2chsIiyqHAE7in881c6TgD0NwwCorXrpoFJus7j/HiG5uB5G9G
N3Hk81FzJXppRH+PRAXmBYsqJMriOWzV7xbsnE4RTCd7/v1Y3eFu36h2rCmhlswj
lYQJCYIvAIMOWwDbFIFdpWu8r65rmjgirFZ9v3mp8dBlR5TEuf9lc0iloLRXZYOt
fJD4bV0KKtxM+EacYmvCGTWripHFnoXgu8EUr955TDmcb3NnL+RS++usCs3Fuigx
vHL90hsRyAV070vfulaW9FV0MOvOSFJosItkApHTbHjL/lyWMFV2JkblVySJL9xT
kNy1nn4YR1n5x5V8XcHDXyrUZY4A9vAg76/DH1EKAvAk3AqV+uuZOuY9gmrq5Cia
0vZT3XNV7A6J/xTcxMff6UMWFocSi/EJDLOAV4rYa80yKBz9j5NapqtlFHeYZ3u7
Q02TqeWMMw24p69XUF6Q+Za11WVjfPM4/dj9IyIFZygp5LIIUe3rQ0FyVPGKOdNa
UbrA4a5eoqfl4XxME/4YoFXH372Ns+2iVWaIsVwqsBphsxll6gTXTvKHHl2Xb1GB
+88fmB8/mVX/Ktb7XWJ6wNV9FQBX1Uy3a+q3giWFTLIM0FnRrP6Ox2tptLtjOJ3z
z1UncpZZtEGCFdO5Yb+t3zzTELS2nULako/yG7eZOp9eVlU7stzwd/qrYyftaL50
IrNcd2X4Qs1VZesPYG912BUlZd7xsgtLwmHiggb+UvHjBIgc6+m/QBMXWuvKWiY2
y1mWa4COiuJnK/mqgQKZNvSt63IrHr3cpLxIkV3+DHBzP1xMQkOSDcSY3ggnf2S3
MBN0MpVMTW54fNE9gKE3THxm4tsTNAbI0fArZdL5bBi4xIJNaQTvmagP9zcc8aIu
d4qLCy6vX98hEhgJ+6rk7YK78NPJHdorPeqM23XJ3bCc0CDxSzns05uE4PMOy5zI
Pd+EXHkBADGjl+DO+9fzaSaz+3eNlhxXtEeJnzWInlsM92JRs1xqmJHMhJs8NIxK
IZrhbhRYTH4gr4vPDUbrC1U/1WH1yFhWUO+qZTrJCIT9GmMRRUjW76PRpw0JpZBH
Are/FkR8CfocuPmrqNLDVwMPtf3E8VjdfIQuBwflXBhRZQIsN35mspxiELtJ18yP
E+Eu+SEw17cB05jrBM7BMNoMsT/dRIRf8trM7hVGqiM+rPkgGvfEsNwMlwEd1XZ+
mklXFb/MU/BTjGTW/5ExKgyjI7d9/4VS0prFJ4Rt2avtfaWxfj64o9uhji4YjQ3e
YT5lHp2qouRFW/0i+UMceNjVu3T8EU56W/BO9VchdqXFaTxJtNEgJ6m2GpJ+2JKq
cUL53ah0PjvQvYDGnY412WE+bCcWsNQvt1r6YNQew/5psXOI9nXelMPhmER8nCvY
RFR+xIhMLC7XHz9EADspAZ1dBw5nxtOYThACIaoQhiNlPPF/8OEavcCdthfu5zYl
JXczDQ8mX0/Rz89Ouhc/Vic7RvTGyliNWcjhrgmnjA/VIN477SBU8q+moY7Zcwq9
0d6yJcTtLb8PFqmj98ngFOSHSBpw+RUBIMvdDHQ0DVCeYnMWeuW2+xQ/njfbfACa
8u+YGrNfynSzr0Mia7n5q1TgAgRrCYiQed5tLXAnnjRTQ56KV4n0t+sk+WkfEPKi
S7xp8ft2dSIc/2UJ9DYo/l+z/UdVpgxlQ3F3su8vzTWi/yuvG17HEkXI+Y9dxQcr
OOCI6145cZfMkvkAIfYj4wSNePl43qy2cgjAaVoLlnarT+OpLd/ZhJqfQPDtxWXT
w4f/qYy9MGV6PM+JNbW4uE7tFGNP1YYZJrXUf19MFExiXtwq0JCkGqa3YyfYFSmK
IObHHK7qzmZWM5Bo/657xsqJCWqRhXNYrAezXiZIPhlnK9riCCY4oBAP9JLVS9hu
fnoPsfvGb8AgXiL8Vg8mpSj0zyktvYBXKOUWC9XjtOYZ5CTTVSY+YrWprIRlRqdv
PdxnmDL1pN0nGDaj03Ag92XoxfsrARXbItPTebWDT00np9bRq0xTLf54vVFyghZ0
KcBGRj4xnS+saDnOuP/D+UI8ScKgnAokmkcWIDvpGd97ct4wA2Q/y5BBC456RWur
kwomJ6bE1pzN8xaIlHKO/+RASBddZj5FFUFYSJctiIr6U2n1o952iZYmiy6aWOdg
AmOEjSjre6w1beQ680jpDOgdJeqRKwiz22p1mEVy48Qtyt8fLTQsAMYfOHHqeL3n
DfEHqqmCtxlLLcOSxF/EXgot0cqB3GkEPwhIxT9j07uSji3IXdCMSXBQ3+uf/hqT
/nmbYAJBZb/QhBGa1auuyjp2lcTjp6WD0Cr8yQKruzhWB50OcuY4X6KmpNunTzk8
05B7FsvJiW9IXhyIW+P7miHgELavSGBUj8cOJU9lCPRNow8UHGaeREmSA44SSXQc
1inZgwtGFpIfZCjwwcqRTLewe9a2UJ7GtoiUw8y5rKyKLrgk3sSYThwg9Z8k4Hyj
lq2vxUqYKuCa+nQuNLvK2odR5YrWo1mUrav2/9ZAK0U5slpvbYzl0QL2U9nmlP2/
4DqI4RVjJf/7OE+UbSrUJUOAZ6djNOwBthNfyXyMabch/PF4FcUxX30ASYlKhfWq
V7Vy0OKdOy1oUUlIN5+A4MOCEGArYcKtlfijZmnJ4iIr343/a+VB/EuPZvh4web9
lvci+SxyhJ/DuJxW8sAdxzYK4zz38xnxdCs9PxMjnDwuPgsummTfqe5YVthtk9Oo
ifUrnV5wMwA2clhq8X7KPsY/rm2e9gEOgP1pnAMLPjbyM+EsbQ3NDMuyYjE1XkBy
LWXOM03EEg4qqVNVVfB7sJma8ZHOStYuvLm7+yzWX6OkUh65A+AnyGz0kvIcSsqC
eY5+1aTfpcFmxyIm70OMN2lWRb67SsjwFNGGgd0KqWXGEdUve4cMIqFKsLmrVMEF
QGC28wEq2QpGE4Pg4seqh1QsbsisFMO0rwJ+TNKFTPWt/yLURT/mhsK39sPYyicp
tg2aCQ6us6/tzauxgzBpy5KoJswwrFOVvyHzxwrqivNyfQ7dZ2U/2lq8g8lf40ki
bk7pSwXEcaLTcW53qggmjXVmOKZDXoqIcSegaEmawgrhsJxkmFDO3XW916RPlsq/
rvq+nFfKtC/KOdwuA3isc/KbePcj5AotvD4perpGdS0OFWN0WW0VMnSqRKFKq30S
XjkajrFW7iT5mGW7nsVh+SGhgOQmP1YG52JSxIrwxPKXIU7K2TIakaTHfROmON0L
wcCjzO6t5U4FPaGZwzrswGv7g8I6hzhJ46fF3bDPfLl5cGUlnExCqSbcs4msB1A7
Dn598UR0aLy2O3TYHubBrAXd29PZEgfBkFdSd1XalB/ElEYXWQejse4IKjIxRk6n
gU31TuMAf3dqn+hBLgCdTZ+fIGCUhHU82qwVH6AzwYI5edW2WGsUR0ORZO3QkvRo
p4k9XofD92GdJiPcJSQMMyZCNIiQCCT9H56+i8qRWdprzibmH8Bnw2B0/dw6nVQ3
cwWdw/ckEWQb04fpWvwDnKRbjGOD/iMJaULfbrRyjhxoZGgUP3KQ2ZVGAb0Lxbo+
wT8ucjJALox6rfgG2lCj0MtAZM8UmZqMWEejH5N2opd2d36PAhtNhJM6J9U+OJyf
PTM0EZhzDUv9LifYEqY/Vi+8xBFls9o+hfqZ2RDeojj/lZLh+99dfOfOaV2p55U6
02+/L0RqWFIY3L0cKbwrMYFRbrcbyLJ8jfSXBqi2XG+twHOGMhhK8Kr1gOh6dUJ2
kv2TC+ZsuM3eEYTSm4+tLlrO7F9HwttomiEttEgNMtqBo0szHDztq/a/PXpQjBbb
C0b0N1EyW4lmA2XbdkJOdNVGzzXEQkmTVQ7ThWyIy65UwV883y7EIX6MvEp2ixib
NoiMYRuifPKlj1c/gy3kQ3BvEQVeHro6LGa/z7aWBEQDmEB62GeJU6DNKauJNt61
OpLyLf9942yX3G5WP2hT8Vs/VDbHgqIVdjSPy8hh2vGdrPueVfwGKiYlBQIVhMLe
fIbcMUroXQLf8pxdvDLb9CbWWHtwdhRRMARXElNGSztCiY9mrFO/qkmPyyIQ66W5
BSisPN8KiiMBRokneGJRTAkpYSnBzvhaZ8LAQsGjpCdYPJEqdhfH+hX94wj07Di1
Qa47esT27WW9Z0+RDj0/b1tI2dkl8iJEna+YLV1QX0k8WN4TIf+kkzCWZTe4AAno
U+hTovvEdosZ2I+e+4M+HI9ScWZrhlI4c4MkHOVb1D4hzVMluj66+eiaHHT6sW+X
hjW3y9XeWOOkuz1d5TcOoLFGaaGq1H9JZZ3drYxDkx+WsNNpBAZG51kGPlWRVMDd
6EYcoiVuSzpzrDpcL4n0xCthLsVYALjeWlQLQ4pNkWe7Da0VPzIolL6Bzu/Had4l
jHdeGhhetlQokP2r/VCHmTFYHrwJ1iI3R6m/Y+uQCDbZoROv1t8WYvc3Ra6Yrt2F
Wfg5N0ObIFYnX+1qf62Vi9+POBaRRQkMMalcLY/Mdg+IGCR3jPKhN+idzoHxSD55
jSudmigT76kvhGhMbQCNVF4gbQmD1WIyQaEQK+VN6e00TYUchzHKRGUn2tswSDKn
yMwwcwzuJiB5oW9vee9lBXr43TvEBICJioxlEhUHDgyzAMbKqw2SDxexj2wMdvAz
mNdJl1dPzTZunhHcpgqSSK4DWWCSq7E/HV3Aw8F/qAPX0u3uAmEpnnR9LPYz7eFF
tJzU4m6b9RHFletYtw+I8om8TaNHOyjr2x6uIFmje316DS7FA2LWD9R0pDMPVrzS
dL0HK2lXrf5EPS3RJedusnPauLA1uoIdtWtoDTrCT5lT1uqSrc49H4UcCacn0Wy0
0hKKZj2o8BH5JPu2VbTgW0NNOi8Dyb2rCyR+RFhr3lOGPBJubrj7r71PRl+46gia
pauEQIhaamvF/fG6fGDOS+z7D2juVD7alKgeEnpyIBDZ0KkHHNNWVEHB0+yeVw1Y
hNrwJDWkuCUnbLCgeImUdhNq4O4D7mnjO/y65h1qedxj+1eO9/pnr6Xz1WMfNdRb
uOeemkR39Tu1vbTpdCCHZEwVbMnWUElQEk6AjXJ5ZwovCfR/PKl7+QOdzkvI4CVF
m3YwJtItfzStmOrXkdZjirbTMsD821tSJKbxqwgGzMvZa8EsUCX/geFvl0zstEEP
nXIyVw0X8qFus34LTU8lb5/o75+cNBg50AKoLONrYJ2wGHmjgtXcCIN2wiuqg48i
FUzFnsXh+LBjVUWq/zn2RNkLCJGz2/c3fykpTNVbkhbI2b8umYYBEGnbLkt4efiI
nSaBjgPRRkD6CIv1PynhLUbqRm3scebayPuQU6ecN86L7KjNzFE/XWKwpSRUAdh8
CJMPHyCHIGBMz01UpteLHvBPbM6FSfXFO7O9hyFok90mrAnAM8IwlPhQRGqu3Giu
lb93siDYjwDLPx9PAdql2NWPnKYR3lD0/whSA2O/4B9iE1RXQDQ0fFzaMqueqCNO
GSfhprK51gepGY8kAq2NwVcvZrUDlqWUP7jQlK2lpaFXqTHl1F4VlTGUznxAPtwH
8CVatHvoMb2Y3nvKzgf84aUpM6YAv1BM+7in+97PlTQGVMgRRMeENS4cXyEjWEr/
gK89KtnPnQw7+skHRxUgTPQsmGEWpNwY+3RN+O1RXomO6Br4g76fLLLax5/Qq/sp
XqU/mz0GmoaxjFg/poySYS0Oukhj1IMthnPBPqrSgxwDxeWOIelomKAwLsU/rWyQ
ZB7gJp3aT1cN1YNlqn11aFIEPzApjHt95+yBVP0mLo2Ld28ndJ4lVJmY0SqeIWj/
S8U4S2R4DlcbXMIpgZloots+o2x7uyqRFQK4nMzC1snVSjz22XL7Q7dBz52YZRQQ
Pfzbi++iOiUPgWXTMs9lgGgFFYJ5hJzPy2ooedNr1dZVKX3WPX4UHOtej5OGK6Qj
GmFx7roSA2eOVkBzap6jGXTTpeTut8fv3zI8wUaBnLdDCmpF4U9hOzrHIokynT0o
89whCLrrg3TwvdzLDwV7yv4JLJ6OmsQEKChIAUHdfjooMpmIIj+1/rHMCHYFwr/q
7wd11+wG52NgxhZRZGvSQSeUHu57Y2r4tFk1DKAUpIkyz8BRquxFs62ja8sVjYvS
ctkM7SXpKRrcDJhNTMf7quSvflNvRRgv/I5d8IMOdxMNS4iIa7rSPNUQriu2KfPa
sa2jau7h8eF6vqgSUxLHcZNP0VPPrqmglMI96yCdQ6Qu6c6GhInbx/B+vAeis/hW
iLmCmq4TBU1nVQb4xPvK3F8T92wrJW6AE2cuq8TiqRUPZJxzeVe62EOsDALBVJ/T
nhyLySFWnwntrz/xH90T7x5NBSxvLgKl6LexlAQ2D7ri2HmNiO19oU4fb7WEdEk9
a4VOG43qNsuR5SM6uRcGrppQO2g86gWebFMzRpcSztsbAqwXWzsDpw/FRFOzN1LO
91jXmuZmk2lO+b2ILS3aXGoDYCUAk6zO1pMHaWomUIV2Kd2OVpDbugvKJuJxLb7w
F93saEIF9iD42TCJqKfJEK/ez/xq3agwKK66skaiklapEw/MFJezKXDYdIRvw3OC
XmgLFs3Djbga7oRAwskujRlzQP9hJ58DGqERyTd8hhBoVx6XTWaAXaocNr2xuD/j
EnlEO+cmaW4Lm828VYDFe5e5vS+w0jsf3ZrJoYt0owvYhI0gG+JmCFHNkP8ZdEAQ
PTKrXLw2BjLLoh/ZSa1zFKsxdWz02RrK3OnSwgLQJWU50ITVe0lipMzwesc/0VSQ
LT2nSm6Ng3LtybQCrZYTxuz+DS02/CXwvUQKBaLd7RoxQT1QI3FjpISKTBY7+oNT
7vPpSVaNAuch10pnhqeglLHWKC9Ycz3dMj2PLtxsRRZ26qAXp/HYXh2uWEkkKyS5
Vz5liOZzCJV7TmZFAWOBwqcyhO5EivnrdHCGgXwxhYAxqhd1rsQNNdgVR2g0OcZo
rQNmlhrFKbzijH+B9pMsNqm8KXgMUYZ+vz1PCSXivgrCdbCgkDK9pLcFPqQ/7YXo
Dy8SNUsrItt3o9K9jxCLPJNIHf3YYubnCoO8Oj08vYZr1VFUpCT6URRD/mhi/QNN
sFNm2nMrpVL2KG8G2QMFEx2gOcDgI1O3EPP/u4X2XAGU/RJzicdwM9mz44VWwPaQ
+/8+3OP3HU8M4FyBA3WmmYtzxkbIlr8V2IUj8tR5wA3S7G9rCqQ46l4qVueUwMNq
nX39iL+wEYjG9M5oq1X5YBUPDY7mxIXi8AR/82X0WgrqIw7KU/twG1xF7DmuX0M3
RSnb0CRSZdLLkwZi2Yl3JnD6EGBeAGh/RiRnF4gV8G8zlK4B7aJUPWoY2RJAMmx0
ruZYKKz8G51aeuyLh22Lrq9qE4XedMIYbJq+CGeb4QV1oisscw3Py3MAR+lrXOQi
5ckWcIDN5y/WfnA7HWXp2XaeX4pJxsGDCpaqYTbVJ1rIzOllFtxk+oUjrzhRHZ7W
rwqMWfFsZGyEisXN+OraJ+cZlr0o2GyKA22v74ITOi0mJ5FCSTM0ElXv4FCNME2T
f469TkSYY76q+2z2rb5pXMm1xK751HHan0wBNns22/b8AudvhFY5EOnHCsGPoKcO
VatakjIe7ccNmxWaqa8/7w/5MOY/QhedvBjzW3Dg8DVq8awXYcyvlR6lISFFL8hY
Sc4e3KbUwer2oFz25N/uLqyBxyfKyHyMMwzYpwJ8Xj6zXqCXqexZyeiks8wDPD36
sw542BEQxEq2IBVncQoJH/IeRm9I9Boa3+ER9YgBH+AcrN+MyH4MF5DwPqmYSGYT
niy1eqanZ+XzBavk9/mityIhRLkbXdMg9apUUbs9EndhGBuCSnkOHc5Dn1G66bHy
CMoQCiY6urCdKxH4i/3QsRAHhlGaLR70phi8SYcvaUANw0dYyLtDpE38dkmj3JMv
yf4bgkZ/zgxZn1MR+iiwrgR3NtTCtKc6HivpVG6ljZ1kwnWptrVb2YPzV3fjnZCh
3oglO1cB67OLwzAfV0A02r65P2W1C3owPytUePu4NkaVZylpMgy17/hRGWAHqWmq
NXver5d4MszcmCpdIXKTjvzeJRkkPG7QozfEZaUyjkcgA6eZH0ujqgE3yDpuXHar
snlXXQDO8YnzUcNjyQXj6Bjhc4lVp/JRmLSYmQ6DWRcpMX7ypi76OBWgmnwdGcM7
8QOCW5nw+H37tsgNXX+7czAELvCFaHYOoCBtDvQn+ZL6DfFxJKXh/xGLJUKHBUfx
P/IrI1Kg/s/PGsox6+F2K/IYEUpMe7MzH1DRx8f1o+DtHyLBnWsTunIwmFWFRqYY
2dBKOsna7AMVsNjJe1fWNaxODVV+wo3h07rLY948WIAz9bv0YQQgTOzTVxAVPSbJ
AfTQrS3V/wwKL9lqZOT3mCQisP+OHferewADIMfGQXqSFQrgG5c0S48ZlSFQHptI
GbqsEwI4VuUum+QyFXFmMU8yerCbJtReo80aD0I7YHa0X7xkK0Z2vsTVH2FGrgUu
XivcrUEYlaA53/J1ec3lO2auW45aUsnYv4hLKawJgV+uWdsUBWTzxVE8bqnTn+WQ
+803/9hZo/eHNIq5zkkiqk1sM4QH7mwtqzpoCtHP3L978hxOQbe8nnvGHkEOYuMy
SG3it4rSi3STSTQHPQCOvpY5FUnv5PdhHMefARYbw7aCQ2VaCh3fkAsUzKT21aqH
abvbfwjwpgoMTijViJilX1vcqQioGH6p5oMMEIXIJY/sXaEUteE75kHHkJyBLfzU
ttCBfeaEr6aeIrBzRWzg25uPSERB10fYm1RvS15MCs4sKwCeTUAeExBFry5XDgio
xRz3E3opr7Vs4gLDOwOthDVKbCEgEunRwb8CyKaUOwr+iyAj+UbPO8XoLK4ZIwoK
M0BaxEAcSTKKdxff6mvhSlxQmE3ddxQTTjXWmV9EcFkJhcuXSvOxgPH8nlzQT0/8
u9XV7ApmIiMKynFbN62if/ATmW51/67LjVl+jna7CWGHS7RDRlIb3CmNm3MyQ1iY
cVhejciSYdZHgIVaJn3jHpY/gPm/WfZNcteXYzOvRQ7UMy4xGhOfyG4Dtc1QtpNW
0Kt29ZrV+BTnWTaxUoJPIWfBNeBRhbVtTWqEK7GI1gsdjv+Y76VAWVfKY8V/fu8q
qXdo4KZwVUJqOhI4X9gXF6Yrks8LlqgCaqAlIFFzgAkSLDSHW+fpm+Cc4beMRYJf
CTSQmmMiVT4tJDk/eh4DVPjTubjoFPNu36zvlbRGrnMOSTwMCy2HNqPJj225i37u
b9uJ+44msdTUtsi10JMQeGGlEUYXns3psl1lGuDt3UI4lyGbT8o2v1l+yq9Bhiz7
OpDQfM1pMYHDsyMOfN1F6s6Uh2jBnEPzFgYJdl5JfebUIij0fiH+lHqvbX6V8MDZ
HRy8B7NClMJGXN1+Qm4dWuHVzm+320dYoBDz7lo+1EHb1b4p7/0tfkiAR9oNw2Nx
X44pLBnXR8GmOPNmdUhjF6FJQO7zPeLT0xZVR97Xv8OGEZ8vPmHN8gFciwExY0X0
MsQM5hLs3aPx+ypOJw6UkTP31Vf3WxCTQdPFLq8YU3iCj/OiendYALn91rgzrrjp
MSOqWqZecdwZsXFsyzGz0nOAzQtwCopAEk9wgTTZ7vhWGad0+TT2hklF5LlFa/Bc
5ioUIVEoI0IrwVLvnCpJDnjn284c/Trd98WCGfdQCz5+QstqNZGQ1pIcgjLcJJws
edCeMIZFOr2izWnKlR1hLleFBZmnbe+77prMabLo99GgiZqKhZO7OQhCSsGSonv6
VRpAvCRhSgMR02kfhGSqn+/Wi0nwsDSL9Rwp/XP5Zkse45AlBG+gz8+O/dmuyv6j
nLVbP/zUiDyG2pVsOXN6YOw2iIpJrIQCZ/1j085OpmkD2AnMBGyVQl8BNUdLLlSn
PzZFfaIyiEe3M2tlfhYWECGh6WLtb/uE1xWQ10pFz9LbvkEJpYnHEGgsqD+APpf4
0OirjR9yyBn0oxd6mJoLjvWbi8z+/+YlE1Mvuofgz0OWO+3QAcDQiJU20DHJuLUq
gMeTaNr4T9h5JDC0TsBx/YI6VmrKqh6u4a8ZZPsdKcLi5X7t2vwZE/I9npMO3oN5
yhXeWeBJA79R6qYYSs6rG7dBr9zSRVMlfAblLvSCe0mPt2h3672Ihl7H5knZf5TU
w9OOze7sTb5Z8oPTgGC8Wg2u7VXcmhOKKmduqaLN305IjSw73zJMQkb3onNu01xm
hO3jh9bQhnPKodBXYD7VDL5IQ5lLfDF0CnuTacHV4NR4ZcmdfGcZ/er/z9NPrpDd
roBj//1jWeNIm7yJvGckaRw1wFdmxTlHYCRr3pHyoBwMJiwzQCadsNaRm117IRuX
w45O3FnwXI+66klCMxVO3/71qXxf1Ue0ZB+hp5aRvnfMkBoudL5iu/FhOHwjUmKr
QkEAENNemOMz7WrXgjnv/nT0oo+gd7xHZdN9Bk7aah7jSxaRmhgykv3OmX8IXQQ1
61dMTgH5dE9ovVWSbnioiOxZvVVRG6iT8kxPPjAqS5HLoDanS8P1eUlnQBUR2+ba
rMzfc7f1vfAiLtlAdQmFfs5ckjwb0MlBfq/7Qrs2me1JVpkLGkQRW+BCyVOJMIYN
S7neUwvRaJyYd2snVFSCkjnaGtoHvzWLpc/i0o/cRiaMsxd6k4gtxX0kPhA+w6Fe
Z1WhwLkQyaOJakq3rm9lta5NgqtC3cc4RADtau7aZdSQ+oSsQyHqTum7lDHZ8xV9
lsG1odjTyUN3Nc9JRcfh0qWVkoszrdygQ5BT6oybj2H15SuCrc43gqOvmFexAza9
DtiJmtOr+nGoVmQbAdPb6Gmn6qUFWAXSp8XkaVLxiwy3CvdnxZCgx0/sVtRyhHiW
sGeIvRvY1eA2DJU4gJA4BAsGWoNhMpRkmYRsVkDmRuH6oppoi6miMlqlIvtJT74F
3jO7TpCuTbX9gSjubbHtzXluTa9DPfSpHzOIvmcU7yWljFf5etQdPvWhAgkWHzKZ
9rctt0IKf5SFoashqxVf5gHmLUtrbpS24bMGFKxm0jkWZTl2pX9g02tvMDFYTp3a
wpUV4/3TBK41md3TEym8FW7IxXM45RlNf1Up2LdR5DVeYVJ4qLhTnzi8rJ6zk7LS
2ZVuC0JpXxyYDyYD7fJo1ArziVQ/+VuIdbQMxbMM+wCsv0EdF2WgyhocOimUw16f
thpapGi6LdieDWrz/V3mZe7zwKwRHj2pUU9+pqNme0VYHv94QxgmeSYrhsKC3Ne5
F/hXvUp7BZQHyOAAYyrXAztJWB8neDpCnclvWta6sx/J3k8TVHJyKPUFMgEIPUuD
QimDPxr1Qw7ZWRPR+PUPxDxVAHhdVTO40KTjAotjd779UOXtYcfPu16Hh4q4F0mX
GLGzAv5cXjF1wcf3MgvzPAiiCGkvn/iYHIbHE7j522l+uyWhH4gMnfzFUuyHIXPK
TkwnaXqraX0ErStnL9cnHVt6mGkTpXfETTv360z7/bwUyxKoOhzwnwy87wGEvyfF
m94SEdsozClH+f/ktEGhnsw1msHPNUaSv3DMCUpxFOCwk4FgXW+CDFHXhm13w8BE
tN07GnS/m/tgF6sP5A29q82vmRfPKxD8h+ha1bFT73Ks8uTBn0Wvbj2RqIQyvXqc
eJ/2QHVZ3/5kmzuT3m0MxgOzb30EPNZjIZsOds4efB0MOT3Bkyxp8R3C61YWKwrK
MjC/4/TOuRZKtBjwMjntFfgF366ngWhMlLPt8UzcdmEo9tt/LUPfllT7yRTLANC4
Gouf6iCUohW2ty6i167Qa+LxXh2I+rzF3S/t3cC/neaUlq5MDbclh0N4iHDSX2jx
WgI6KdvVpIeGrh1hpUwf5PEWe3a914oZihUx9HWgRg6JKU7AAsUEznpVDDEdEM3d
CNLM4zEZ8ecO0GsWMKGlExtDGipnbR1EP+4SxaLoOiKrMIBfjhtyOD/7+3ew2Sfg
1am0yhgty5zYdBwC9BVXGy5WeiJSfszt65B+Qu9qsV9eS+qx63RftRK1VxZRrHKc
RZE7FuX1JwPv+ppT09xCKXNtZp5c1FXxOD9SP9i68ImrrdZhNNF/6bcJA4APl5CR
T5irYIezj0XLlLAY5l/uK0CiAYTgD4O9cVmNnoCRru09D82X11ZlV5g5kc6yMqwZ
riTBODp2STeQBfSsTMYkCiq6frioQ8ELb5Ig0eemQd9kqR423MVuWevmOp8MgFZ3
c9DYZ2sQxH9/AoU93IJLkG5yI4rfd8PDbyL54T/G1OYelafmnj6WZIgbFOviGgpA
dllRtsFK6xSSChwqJKmWO3hgLb4UAn4CgaQch7wPL/wIS9LCAK2kScY2tApkjDxg
fF0yVLxsxgjAWfmybE8naorRytZmbnBq3d+3JirrHhyUugxs28cHijmbERDa6BOb
0dFLeE32Iknvh6tk3gRlhSkmWKERxPWN7TXDndxDROw4hUhXNrxqzIXpr6/liQ98
YnEyXAND3Kr9wdVZKguqYkR2rZtUay3aGP1geFLWlnHu2MHLlr2MG4v/uqgP6ylc
wY8IbjzWvtkMP2BSflJ+vEQoWXmQGBUtCkgS3rn+gnulG3ECO5YqqvkMh5t7vkzJ
zPrS1JSt0Lb83pyBVmLlSbx3N5ocQMvzf5TAaxTFs7jayewbHFxzvceQ7d4AvHrv
hMxEVnLnHoY9V2LxEqIae/Zx2XfD2erV6SzBe62JQgTWsPS2XuubeFV7ChGGYSKm
LPHrHq1Z1lDbKKh6CP7Fx+NLBnSGbQvktsR7IXxrWPxultBZGZeaPGwxEEgmaoYG
0LUFYlIz26ukk6GUOX1Rk4+K1nNy/IwPxyEEPTm4djjImvs6DkM0FGQDr3YiPSrF
1WRL6uq3p9nKrsMg0Xu2PyGet1hP4W855Mvl9vyhdzmtGrONHHm0YCL9ybhCYdcd
BRJHIxaEdcr7I9SaGw6VxNYL1NeXSh4LPNxRSdVfQY+AcYAacxYDXdhsrqueQmBf
F0IIlhaN3l1npI+lXVp7+Gja15uqukRlvVXGq/WumCMJoBu01jBM3uFxX126tRmZ
fYYVQVmHqqsQmKeAkbmcFRN9vyCEy0J465GDjAfyfGqX6cH0MZFze02bdQ/5vUQ3
Ge2yz7tb8LFvImSyXArwONccTehBzwJmVh3KPHHuf2vwNLLbZYHwHDugzmghQoNO
EJPD58J3XyzzH5VmZqMTrenfFeBt8G+2IwmFa/lADVi74VA68fqPxIxeZ4ZE5/SE
ZB+PGHv4JdmR6ZsNJPajDtAjlgV/cswhrEYdYTZYsnK3wQISOhVy3wa/SkbMu1Il
+Yptv2HHknhBJqTMdyzLkYIw8UB5PQhOHilgnurTHNFwseo6kQ9acpABamoy9SQ0
4Doy9e3/Sf3Bk4+bFdFKgJ7VUzD6mDLEaJ6sdGkcQzwifSLP40qBSlbAnM9iPzo8
qZlgQPEr3qWtIJ5VmtXSzq6/pcPvcuzl/ajuaaFyPtE69BPtzj3wxzmzLUJ59SCG
sUo7D8XOq5r8GbJ2MjXRSCbMYUBS/7s1iuMt7wkaTLx5XqlfTMcVnZIoEqUfG2Z5
/Se0JFJguCo0yEq+ylQ//DJU7y9RN8QzRnzfW4X86SVxWhaqp3pLNizdxOoC1iQX
higjgq01SY6ggESL5HVHyWxUIAiJdCBlVEhdtZZFwZcWRQaV/jM42ex7fpj7G7sF
TjYK9/N6UzLSXuL3PEzJ5nLA3SSbWsiMx5bwBmcIBRdFlOHiUU/hnnBhxxefHlwq
Tu1OMDFIFv7UwCod5e2aHZ/+NuVkCFG4T86kIZ+Skn2pcL3uJq1kOL1QLem+Rh0m
02XpO19MPdpHkIrYdyUhDo9UW6S2G+kIOwbM39M78S8BwAT2imUrwBk5EW7xbO4a
5ytkmRi3k0E/Mh9Z8hhFgZO1zkKZz0qK9ii1qrB+wIPEETWcmLYRn7d1EzbJRy6W
BL6hRHe3BI/AdYoFJk5GKT9F6oc7nhhWv4YRITtqRD7Q3lusDINkwKuRgJSXo43I
Elf56BR0DI5upOBRqlIqx3vwBlJ91m1ynVrWgGVdoHf0zxf7A2rulQvb8x4sk5SR
MlZxM+SN2HunzX8tvF8zu1iBK3nDeEyRLtUnKzrOrpIr+tHv3MB7Jt8m+GibZbdT
TW5dHbSKY9gV+YrjrRlBW9RWJ8TG86pN2ez4GWIonVLzW7qyuakeKE+c0QrI5iSF
0h1pccs5HbSAl/iddlnTn0YeHVYblYO3RZcUYiT/NgZSY536rvB+FVxgpIFT8NpQ
Knqed/4+yCXCqAS8izNbqbW4LUPhQafs1sOG16S06Y3IVSTg5BYpmLtCf+bHqqnZ
QHmZFA7z15V9EcbgKexVQW4f0vje1SOcz8ZDD1FfGd9XlFsFHiOd8R9+0p5fFX+4
FQQ12JBTyYVDD9JbBicZ2WTNsCBFyyAxYzi/fz0Z1O25719/2xRAci7jmihQkUZj
pOW88b9dpW2qIbb87pPtzAXCYj9IpE7AK3r0HN5U94MOwtuusQdWaiogzyYf9IsF
D8mXNouE6fM9MWpZbgVIvYbZ/qlD6BLdMf5Z96X66dFqaqQhaOyrPCdSD7zEGgL6
fp5pPoeeZCXf4ToIsHXwPGmvTg4HrKfzmjRFT8sadQlEI5v1q9wny86HCED5oqiy
hABTImgcNBV3A2sQGmnRmRGdRZFgGwFZH5XC3y2wyh9n/xLHAwOd96+fPNxdC1L1
aQVG4y4ekIgTmExOcwdlQ3FW681rPkCVP2hfHzfIXbuWSHWr4MXw2Jrmff1Vv4ov
0mpLQH/D16l4oZo6JXhn5YidG7ZfpD+gu4WBdvtudaoiIp+9Voftapz8yjhMKkXj
x76AXSOO9Nwtpz9slcXMEVwv/tXjQnJyFcfA43Mlc1sIRsol1miL1RyOyGmniHjO
3V/9A/2tEaI13i/Z+ydlNH5TDlhavkVAnPAAcGw6S/+cLIkyQffhx5w9B/C0j6+m
9zyFfOnJwdnGGaB1rgSr3SngXpLow3ltA+pDxEWtEzJ4uSDr0aoAial/STbqwzJf
E5GKkO2R1KDKsyL17O6iG0gdPS5dcdDaJnYc9V0JY4tQZ+SxZ+CIRt/2dUiLBWg9
gSBJ9sTvh9H8rvC5neocUtgn6wI1AdES2cAoR42IRELC2kDkWFun+/bOXuv9dJSc
nM0uJxaPYKl+T8PSDeQItCaYrQlzTHg8PMPv79wSbtJQpqGxZbEGQCA6t4FtYUzo
4ZjVa94sndxilavhJJD57vo/Tnt1sOq+wAMR1Vqt2wocK496kI/uezb87t7gH5Ig
0F0wVtcowsq2Phe8RfnBr8xKaiL4L6H9waXW+pLf6Lo0HoSDyKJmQ1/LWIrOGPzA
S4G9+BGSK1hFH2SMlih5dK8MPmYdTyXNaehuqxUFdKd8lWJ/TCDrdkK5M636B40U
t3RAHhzmAxKebtRzyv9GzgrTEN1PZBteVhdntYJEBcnjZ5/R6GYlkIUAap7i61Ca
f1+KzmPerYKVd/9Iv/STifqt4w3ajd1GMDhDpUdzr5VkiNrow4v77FFWntRElZYY
KlDiiR3+xWK78W1bNizgPKO4O+QNQFn2ltqzXcLB8lqI1goFGPgSLV2N5IAB0KeZ
gwfFLKiBYQ9rdNCV5jDQOwvSNeFD25U3bvsQxK90/pw1HoLrTR4f2E3yJKzgKaSb
dadx3hCOK7jMhS+xHD1yqA+j8AZUoJyvsCX7Jaah9mjvvSn3uIC1JGu8p3SRq8IG
LQXeernmGTuvPYGyZKOEX1X64o+p9l89IuExNDGuWcn7rhPYIWWnKPG7QSiPkC9f
Sj9qp4WYA0KLtxo2/UYy7/OSXh4wyYXBciI+z5xHcmVWmosGcaWLsMNVWXAWTZoA
kGZb8Fh4LubtZ5PWBx66lHEZE4zndqB0Bapu4TRtYFDDsMyvL8vQytodQNo1In98
ahln6guVoCF6liJm3/Ulh7dxPx0PEY/4ossuzY/WlTn4BG53sIzg63EuEFjybDJ6
gHUd6VaLokX+hZI1mlC2eyab/SZLwaH9awdDfjvFBUj8BS+cecDgAkjy546XusqL
qeZFIHqr/HP5/7SYCjJiwIZn9IeOB7Cw5VAue5B65Ovu8iY02UWGUn0W0GRN7vQb
GKE6RZ/u1EpLSwr3TeSCPjEGWkrRaX2q81K2dcyHmfQ8SUCSFgSSzhxrK8TrVXoQ
2hD/qKx4QoWL6dbiHhyNXzcNd1NnoYn1OOP3LqnCp4eBAG5clCFaMIOSy3wTSYAq
WtzvdZJmfE7O9NRbqUh30fKY7N9gGuvINNEQP+SK3RXVyWsPrkbavtNR9hoGvPXh
WqvlNw/olPuj2v+23hjWk0+kCmOeSZhjmP9cUWCLwCl5luHQ0Pf1TkSn/Bq/gla3
sojGzyx6uZfYS1AwyYAVZnbIrQvyISf13vwaEwlJTNwhD+e2+CMBoaOGCPJO1qym
OUsChGEJ65G2NCZ+Je6vhNKhjln+OFOkwk9+Z6a7vMskB+0q/OAqN33Yz+x3ToMk
yUUaF+UA18+RXPT/LM3wuvEJP/vHpYhuO2JCKVM/zCqWyGmAwru9dV1S69T+8UrC
1E2rtYrO6RyTmziAdB0t+VZkK0oY4V9ZS4UeUysoPVqOBr6wi4lGu6VrJ3We1lBa
Dd5cuf3lvkcdvYtcytOajhhYcybAChAkP7dEpeemwRfsqEnj5/H9f/NuShHU5EM3
lvKd/sattYMZyZsW2As9p+lJPx6YQsPddgiBafLATTVQSgF2q5XKJ3z7z5bVKhlA
mqISaZogXpz6bX0TYP5GNyDS+T4PThzLz5J1Jkt0cSt34aOscF4Es3mKwqmKBYtu
0ygALWTkEOlQgk0hbO99d/NjB3QUYt+UMRpVJVGigWUTf95SbjN/QF61hNbsIbGR
gJ2kN8pka3VUrLUKkJ/GCcoxNzJSDSaaBSCdIA4jf5lc+VcHzFVjLpC4tD9jtXCa
iHdaIJSKRXLCFrafNcnEzjScfZVjvsBFptx2SzGpqNe57BAd7A7dKTlzcR0dQBOt
DOPX8m/jkQz/3HZxZi1VnjgBiVZnrr7d8OFuFGbIsVivx1r+MBD7IBsSxTzlz0oJ
tAMeT7/2Dyg9daamTR6xhaCocH2ObKiyMsow6uNu7YapQFq03e+lV5gnc2LcXaQ6
nCUlN60WxAWAtPpkTQnI3p1crf2fy9mrSB7sPOU+vx79e3s6hNslqGTGuGpccJFx
XLKNaM7HXQZk0FRclzlE8Rxshf1ILoWfnO81YNk24wIm6xZdZR7ap9JsSgNTG3Oq
nhFrY+pZdWNU6MdiGsjpEAHqF5SxL/GHgj8R4oSRw+8XE8t2li9kM0etvBumVK/x
bA0shRpin3NpYdHwQn3vO2l4uMjzgQG2yA6xRNTxwdr42vmatvnQ6QI92dIo4qGw
5vZmmH+BeJM/D4yrKs0x273ZKZFhs564T1AdiyZDy9w3emOhQhWHNart5DP4ElIO
HMWJzeCprL/qWw4hhmmN13qrNGik53DfRDGAxKawqBitFaf6wFtDVV42g6K6AGaz
zmhTz0zRrXB8OhESPnoQFPxjCRs2X592vVdKbuWN4KhQm/tJ52Te3XksbdiG/OAr
KoJFApCh5/J14ls4/yhSZViKN3awG1wg9+/sPVJjb6+nfDVbbZxZD016J2N6G37b
a7qRBaE7QEgZ8GMfHEZTle1UtE0+x/LgCESpmbIJTz2jivVfjq3tMQIkiPlTA08v
I1WfRC0kDcwNyy1j2HNzZp0aw91FqgolGDQ84kj13iZluHV6ujnTyBwFBGhVyrzb
hfeSPQaC4Tw8OTzv6SGVaXtwYdjyU+gy0GKYxc80MWaSJlw5Io0zYiLvay0NKD5h
mjBll7IjDFwjM44vrvrBQ4eBdew7+2UMu5+YElDFnBjd0Q6g67KKJwYUbab/Yl1V
nXwyaKrM87n3OZSLA4pRMBS0kU6nsuVrbroVHH90Vrca/RCJfnQS8UIarGvwNzK9
cwO8B7E+nl0aehL1vCP1QaIxMW/oC00ic9C6kK8T8RnZ8+YfK95CY63oK2OtvBhv
JlxcxaG1LGHXn7OlVds5PKq2gSu+M1222xjcnJ0w+JrSQgdNYPOJ/J70SAnAKKeC
mDVMYpdLcQXXvqr1Gx/9WzafMJbiBj6zFe1zcM0k4BUZQcKvy9NkfpvK0v9fYaZX
7vf+XI6VxufsOZX4747fG1NTH1l8Mzdhp8A2yFd/O8Hg9NVMnaz2E20CFRoKF4yL
zuI0xGK2dSZv8d3EdP3bL2rxg6GTkYtX6mU1mWGLQjcjKNIS664X50n4mnGZLVwq
BvEjwAwPmteG2rjT49+WlRRzlilakLOEGotUsy33xRlc5FR0z+0vW6Axwk3Npwa3
LDa6aAybz2HN5ABIlQAgcwEvDpauj7yx+u57XVjN8QSxCS+Ql4aQLlIpqRrhPn8s
7kGNUpOxbDqV73CXTK3rwX07/Ryzj5WUmRY0hlUBP+puBmy93PLrFbswPBmnSA0z
/wglhQjsH/uPyxXq13vBHLoK7z1TVYp1afrNnnJaYtrbtqy2ZThiJhef6oxjPobR
gv0u/sBBrm+rXrPd7zbME8iwoMXKo4gLCHC6Y7TSj5l0EQdWxkvdnE1uB6ZVTt2T
y3hAYUnmEs3Dg4mCW21AAHt85xvAYD/LHzRVoP5zFwV6EbTO1N2Wq+2ZSLr3G8zz
bdVd/sYr9uN4zzi2CLSq+ykf8t/6vOHK/FUhPeSMgL/3AWeIQhsQPYFk0VLvycY7
qUQTpsAzEGzBRTxynMiXKI8oTPw2PiSQCD2jOugoIZ5vbs+rUNH0Kt3ibg13dVlz
tTsXrwecW7MV6BxJCEAtRoKuWORhUYxczlOJZsv5NPFh5kfcYFQdNB5I1PrZMUaR
MxJhQmijpifwDhfNfg4Drdi3P9b5UMgFkQaMzOTGrC6z87Ge+iFAcMI6nhUKJqI1
XYZpwN1sZDJMiS/jq8PnSLW/EjGtgDlSA9iXwy75o/0EvSYBS6+C414nespMtjvn
klJ59S3F0VBLl61Ai/Vs7FOAJlqo9g+pdnqKnCevgmDpYWQG6nS8KBvSEVjhc78a
poWfINARGMjI3qmBul3KpwobBklHARzRIESk1JMBPajwt3wad6Rig2lCtFlXN6Al
D6ed1efce+vmRV4dzGHTX4sqWMsPH9xNedcu+hTbYpYxr5cackhyHoowBDMjjL3I
2Sem9w6nPJMhenv7X73UVWHRm2nALm9o6wy/rZj3abFNAU04ZEyRBeTrzsNCE8Gt
/Wn/8H+7M8hxxoXfYPOBTIbHYod5DSsCQ3zcCXacri4jFKCpgttUoaUPh9sXzgLw
1yVYRtTssyD3wOw7oXqDrEbRvrcpgKeyvqmf/NIqe21wnbjky+b+13+MasmW/PWR
JEjRtD0XGYPEgUiIVFLUlDc6Jz8tkvPJxT/kmgCMmKXCjPATfhPFpGvqvPCoa3VF
Z1Fw3IJ7sB2m2uQzDjHwljp7hAtji1iMO9W+QZONGUK0rwGdEV0HTcVMchFpwMtM
HfjRT2QpM7e4wQkR4m4T7kVRVB2K4PnV/TjUBI2AJJ8d7Fswud0y5sKPd/5wi4o6
gMYY/9z6BMXWBq13Gu4eyek7LfZgWELyhdAiYXdSTsNgqScB6bnJqzst1LDyZAmh
xhCTpd7VlR19oUk6rwCtOloY/nswiZTEzbriULPXabQEJayh67I7Sh+sURdUpTAB
idKCyTyHzg/+4S0vSxXZMX8cWlLMTDkktGX9KdShI20b/orjI+vojnNy3Dql1Tzw
RQhFLUejGfZ8PdkNglLX56J6HPIHR7e28B2jO/MFrOC0siq4SVMwXFYo3cF9DjVQ
4yVfu0+fPpCIJqNgZ9jBq+a+JKiFcyRdFoeauRtNe/n3U5YGYHvRAyTAL230rkD1
l0SJggfRh3mTUkwJIk9F2F3Q4VDb0veojd/YWvQt7aXGnCvc2Ni6srqIGthy1K0k
c1/rJOq/GO88QpBRbvb6mdkI72u21LGJ1dfRedZLEzX/cbf4QD2/UHvzYqHMJ/jK
VbP7FTtQydGa5L4NrggBBi63LlfxzIGJhxli01eDKKvwGMmZ9jplP0OUMKqCpm3s
cLDD5JWLg7tYB0LhjMLgpMp7n0Bv15k94Fqqb1J0aoipPgM+ExPCBJvruloztaZU
jKzqaO+1EljmXc4A3mkhxMZlAH/9oA/UJ9Rk2+S+N/T6XJqmbuUOwFOo6/nMyMcT
run+9bLXmh1z5du+sr3pEXhOxrvfUNeBkaAbd25ZIWdYFQFltJQSBux7RrX2xjRO
K+872gZu9d6bZ0SrlEZbsJd56Rvg/zoHyrgVI0R2clITa+16xNBsDryQQsQJsCWx
GEn/llU2tzT0SE8GN/IgWatqvZcrSwnBD3xcAvqksoopBv22f3TB+uBx1yl2THyE
KQ8ogZiVKquISy3r/WMx03EHKwkcFtTH01f7tLx8qv9xaAx8dpHcWIptu3E2yylr
f8ZSL/GkeWWJQnR7GuTAQ5D8Eh2xfJZWh8nmRa+pRAyqJ6bHFCn9uktpfjP0Qdyu
PhIwWlW0he3SaVKiMkoMeC5f3WQ2b/es9jXlHyHrTeIlSEG/Vqt8gEwLPuIDGfnP
+AMu/E73BNz5kPHRfjXpBLes3Ww/yKIXxXJek+9dwX82dgms/Thjs6GxuT5qQZSJ
Vr7n1+pAgbXcHk/v9kIDz7n/jSPsxRRd1BCvo4SLHTVVjhf4/ixa8HxvJ+fR93n/
4PHU75qVrd+3XHGw2NZTpKMdt9SyLwNVQY6uvwZ6FUnMXvQxmv3twsqG5DCAjZHH
3Kefw0T55pR5FWa9VeELH0dBjMBdMf0zZaO+EJwq6BcqrFtwh4JT4k6ECHRhAzlO
Iu0yBKhqyTGInml353Sfmr9fRu+1XkXH8ASXK27nANHckUbB4vAywI8kAYDQqVOI
jS1x28D13on+BCD6eonGXOlNdfjmQRM4Hs3SFp7YNor7GuAB87A4DrxQQJbGl/3C
NXUIhe1/35Us/Jys8vOb7WIwELzOqvjOCS7K1SBmR51PpwSLXcwSEV5pI9gMrJZl
juGBXBcTVtWBH9gAkUnXkRMQNHISOFh/TdnWQtKPUe23fqQ+v1FBl2O2rbq2qdLD
LNw8KpQvRJEviGba80VavVdqWidPS0XdFmN8Hhvl9t3s80qd2+riLv+SXUp1fUyb
V7eOwMlCYW/kN3o01APw1NiI+AH0uLDl6zVwWvl83gDTlSmI4e6gVQRkQ28kOA1S
27TIrVp7evwXfse1w6+0EHLvSCfa9YIT72RY4scjwcTfFzyC3X4R2Xp/uVVvoXUY
uoKqkPhV/CkT2q6SZqGEoCE6df2WutDc8MBCG19wfknYqaZ7kAo7hM85pePte4aC
gpXonnlAeiXaeRNzMTv62sGSY67Ep9g3+zgUubwzDlKdaszxrg4YdK5qWs91nawi
sHnL4iVkmTEfTsOsRkWY35aQlTDmJtJo4QRq6l9tEwoH3OsBWBcrOQbwHSL1fAlr
TVJ/N0cVDUfeeADreIZCZPj8VSrjYlUwdYcbJq4O5fLrFn4As8BUxvXj2MwAZegu
U5cD7/vuNq7WhMkQ1HQKSym3W69cNTyyIoHcW5Om90hunosV8JUs5yHa+Hlhna7t
uQSTUHJHm9ysrDnchY7iT3VC8fg1V97SJcgk9ONqxySVUhqHTZqBGlOQkKByOIxB
TugKhF47JUNppPW2YKwFP/yrIorG3UCtNqMTg+eI90RarXxM4j6VXzescYnTuCT9
v4j8zCYHIOUOZzj8bts5n+pe+taT5LGHLaEXDmnS+kEXBHlRc5rfdQugjEVCDyLw
Lo5t0zQNrmLSe247xKHsBZsqWkZDB0MTuVgFm7t0WRBeNJ8zFCbopMbgXP+9ZAEI
f1PSGq3tKFcTDtH9CURLAIfeONTBe7qNQhzPs6hE/PBLCHa1BPaf9sTj6fulP9SZ
sfeRP4JW4fhroJ9fN0pN5is3ntejCDqNa0cqHP8RgvG2NGUr8OJqfbZ83Y5vR5e8
+6L0ZiaYsR+w/wLclZJaz/kbxGZOhQ2opobUWOJSEfR6ZeSkSgs8Z+nBlOFvZjXc
H5lgpQ4r6r+hzRJhRcRCGwV9QG4jgCXH1GwPT8LaAEQKtRPenW32TLrJ50Pb3GL6
rxELM4z7hyp/IWVdRW5cZA6Staj3com6fn8UaawhFl3Bg/0ASVlbSz8cDVr+t49M
hgouGCItEdkkaKDOIM6jVSVQOBzmE/2Wt+C62R+n6xSmjkkcAnpHhNcLYQALlOuT
Cz2m3Vva+1kDRHr5E/E04VE1gaHire7Id8XctP6SqbE92ZSjkUWb+ekWqySPAMFH
VrF54mUgnjHkRQTwaVbuggz95hoC1G3rOdjg3ypD+p56DnKUCKniVWFqWF5Vn1zf
KoXBMixYZgV5wB/7ywlGvy3CIRnut/i/gd70qdFvQ+1qtaAroPcrXNzT2LUPOj0l
ocxazJu6givAB9vZL2nGPDgXg6hiFLm/9ar09FtSEIGzuj9oelqhrkiprMaYjmkP
CpnI6C5AvQTU0mjqL4w9fzuAiZzWuYk7+/EU4Mcd8j/mfUYvxy3dOdekKKF/Ceaz
645rzidcnmjNSNsTlm1RX0ighXeyc5vC/ekrEGqEpN6HFewgFg93/ZCrlXm1yB7I
5A0dfRUU9iYl9pMMtlBIuv65c0v7mYgNyMI/Hk+rvXszL271NY1Rzphugm1X0k/0
dKcan8gvleC1KB/ZJtWxq8lJD5jZM0CYV64B5YkLrH5smTvMamQ9hnIBtzKj8uif
jGcJOgZ+FjbWmiVnxaChYs5DjaddwiUox6WPcU2+z8J1msytME6uYL0VzIY3h5Mz
Ju6uCdAFFO4PRrbdY/VO/RsZHWSDukr4XdB5OlBqhKliLHQtt46MtpO5iLJ10Wt4
oBi4KFd5YLoUY7GBFmQq4UFqErb/KiN7r+By9rN0axkl55xzY8VB93wzOxD+1LKx
NDMnIHoc8jqmn99j5LHfBd3iKkQHJbbHl7qyZvlOk/Q1vabMnTJBOm4khucqY/Ar
XbSQ6lXpRGjETfqsfgEuI0bcxbctfFkeWktTBIePnYQsema4z0LL3JRvvcEPqyKP
QpBFm6fjdmApOFgph2dBASm3L4QsCUeQmBgHbuxTYUQK4iu7qAiH026FKIfJNi4G
nu7MQdyCl9Jt9N1LOweqMXrswt34gM6U5SusaZ47kGiFr9o+yR1vzff4R6WE7Vs+
Y04LheP//5QpiYOkTKbZPE6On4jyuFApe1ftc9xELXxz+GAli+jAWnBRdfp44FnA
M/bvIXTUKM4Fx79Bg9fYcZtlL9VddlaM5LmVtsS2MosMGK5zLBtTdQ/PdZN4HtGW
fOnGhsqDdi57nOJLeGySTok/+pmT8pd4nSqovk4yNWALIbdg5DqH7NZZ6DhPa3a9
d9k0Z+53o9GfIbdyG8GYj1iXrUwJWJIvKIzPxgf12oMe0HY4DqlWs03ic8AqfzfL
r2jGnEO6zOW/FL/X2u8YJt01W3XOfwBon3z3XlQGAV5knMayKR1QyGR3SzEM8Z43
vhv3roK5DMI55Ox+XIw0cw2neAvE2EQgSx97AqUR9JAQxjhvQD2FUpzhnpDzFBlN
I2VG4KYNt9BdnjEh81IiVWBXZ/Mhkp7CekLjDeVfARRpLu4Jv4ngsv3vMtzH4k/R
MUHpAP8OpRbTFlY2qaj9SgtYSQgt3TPq9ws97xyBRSxhDyscQSQF0kOOjHHfgGZ1
Fk5bqFFu33VYnbbTcBt7G+FhjGHqDQJzCXPelNRBoQdxQNNHNtrPq4+y1tHEJ2Co
8tpZDV5FCs+h7AsdI2QjbdPLvw8SB88VmceCyGDljwj05QYeq6jeIrEcr+GqQzTf
XJtTU+EY0en8x3MERabl6E76iCGSMpJd+oVGp5CD1p0/wnvrkt1+KTBxeCAKsLZe
lW4PIXGnyRjpgU3nwGrrD/7zpeEaUVTtuUgVyi6iHR+JBeJ17iL7pvsE9sG8MqOu
zjFSbIpWRZ/Dpx+bj/1qWbvM1unoViWkIPYMXjX10ERZw3xCQ1cMt81+ngCv2elA
IcVyrWzXw1Z73ApaWhXjygQBwqJ0u1uJ6ILgh2Yxj0N3FBhciIMrNVzc+bL60e1K
AtyTPPrRUa4iZ4UyQNkOPRtSKg4b3ZT8Gmte5Rvh9dAfaNcRwAqHDR9LTB8/tVic
F+Xi3i/KiGCLFdUfVo4hBGU7MB82TgIccb3iIAeO+pkIIBVvEIhgIUdiE9h306TR
INO3Z0xgNZxBrEIg0jjsjBCJMOgz5Sd7Y2NIuZpgDS21RgcvVi/mqykhMhNfCAkU
oXu7Ez+EjHt2UbHN1AZG4AbXEXaRkG6c5RaNipc8w4wPfoSaotB3aKOOsfp8XaO3
J+SevVGEYoDgvtvQpLQ3IeDhF6mQwgCsM6NUvHcRFJj1Ya9ZkHdX+ayMgYHG2GGh
ly4720zYpzAtmvnMn9HL0pentJ6sl1v1Pejizy9d/6BxVAs4rc0CNsoNXxc9CFrv
8jfTcXjVAeIYQ9WwiHPXQCpUJMM7tUPGyp81u6nNUcGMDCM+6aHn/HVNbqRDgz7z
FsF6HbjV7agyzLm9fvIl6a4tXY+Vx5QQeKgCJm2URATJ3QLOHK8qr9Sw2k/XWZBR
EUNNQz4vNcEanDrOQ8l/zycbfgtFVVuFSvLsq7kuuG/5m4N8bADuGvxCd8F3/ali
3q9NkXg65Ue6zqaaYEu0lVT/KN6NMk77WQX/JbgKNGfVYrTPNosblrERv2yqhh8h
f5Z19l7LvfrwdW2206CW6vNRa+5VsoihEiRsTtzzLvxZ+2qrVy9NnfjFlodwzwyF
yL8vXcqYs0uxv7H+lQbTe6kiP/hb6UTvrcCp3a+CKMnBEAb8Q+4tOOzoHQgFRsTN
/jl12Mk1iM8YCecaPHs6hmEbCA43holJNPVQR1ui73aMH0c6qDwpmm/atyqMTaqN
CkirZNoaKoBHYLzV4inb4Jh6xYO79K0ZeE4sRk6sU9PaUncxsTAmi6oBn0nxhx1c
V20bgWB2ByjYuFGIjFPPnaz6I/G4zaGxDYDbnZ0L5bl1mb1TncyFJEyw8KiojPD6
ZnrIXDof0ftlDsIbaM7VtzUeJMS/zparJYN0Qfqu2krNfv6AI85VrBd/Y1xtrqjo
9GZTH+cEE2uDX94n3b81rJJGhhy5R+8dXqS32EwYLJ/QRQM7DQk37b/BECWP3xpW
VqamVlkJ999hL0ySX7M3oTbqPy4flF7ELBxjf4sPR9KyQQtpGxKv+r9FOrMlSv6I
a7X5d4GEO8XNSg9fxOo7GJe5AarSBfOmAZ9GPAiAVL8wtMmZ9+0x2Y45oP254+Tp
IaHnK8BQ+doJrnO0cNil3MtMmPISdrqYeM536yBkwNNfCaBNZTqPAamNktizF9kQ
vMr3jmJ6AdU69HPRt5oA03Ez21Jlp3c1nJRdWPYpoUNuTkzKPdPGbOtw0Js6CoVo
Ro/RozmVYLTJTBBSC06/ZMHa5/hsOWvBqtemJXTSi0bDUsLPnJuxfoQr7ObU3Pla
yI0UGo8O0ToCSEhvfmJ8WNb/3qguTqRkQ2+YPpKbd5R0oCgkADP7a54z276JvlOE
C/xl3+sCXYDgTgjot6kRxDi/tdc+ERXO6YVROJQJsjZSlV/q6xsheU4wiEqI9eNK
Z5cinVCRmu52a+dufrup6G43nX34Zd9Gzb5FyXv1spOvH5KOHjRutk+2qGh2gKRh
I2p7SnWnys9J+TNUVmomh7AVYgo3wYgvcM/V3izd9HvLDwZCpk8psHZA/5GUhVqt
tOAypBPViz53kUUZtYpmz3BGeg7U1SHUB9MyS+yejF3vfzcf+IARtHI3ycTgscvv
x6x2swr9VKLDZDzU3AT08u24w1FmcCFOE1+4AMq1t55+gRJ6ZcQ49gZ0pc0eRq9t
kc/vSEK1bq8RRl95LZyC5ex3Q6jxUd4lXHJ8tgnzJwFrkkVz0yITgzaamnhfVHXh
Or8W8U3x6sHKid61H+612fS3hxLEK3azj1Jxynzr4wYaMGrQhAR8MPDm4XgK5l3N
f4AEbg/8SeHLuNlXtpI3rDVMHf5dksSiCt/1vEe441TCHjvM3YWAhaPFOkb5EGpn
GAqIj7KsCF7nKad9bXI8Hy6qOHSHORWVNlgRTP5I4uzmHgctfE287o/zbegph5sJ
/NH0wmJw+SyUqpChidANqtWEyrH6LEOZQRZ0slGFonKrEKqJ2Y9RKTkCzBdA12Bu
KY8Dwrh6y23VK7g91P0Lgmc59K3LN++0f/yW025tSRPMF7z8IDgw3WJpb+0mf+DR
Uncy2de2IMD2tKwuh2X0gYgAitT5U+9EnyHGPWqqhWNIyprvA3Xhz5RY6ld04ga+
RmAh30ejfMWYuCyXiPHz57sRpplQpdsWmgvQlbSu2UM74Te/Ufa8GcQtjMVdxQ61
3eq4zpC2y2fgEAVoXt1kcgPnvursMM9JW3LwS+x+D7xrJhMf7m8tBfWexfO1IVKR
SCL/gvWD/chApLRrWgHQKD4TGOEmrs0FLL5zKipjobKuNKFjeW5TRuJh5aqMr+RI
AOoj11m3U/tc5kS9e8ytRDk+bwk/hy85DVkfaEZiTdSXC7GBIoekYEJYhH8kpqDF
mtzZCPHpAGcs/DdWbT8WgccKaN0v04n7uKApUjmx1kG5tGJVBq6KdxXlGeqXXrUW
dJ7c4HL8q3TpoDWpo4ltItStYLnX3hULKX4aQEPi+nDFQ4z51s27QVnPA1yMhFll
oUPSIh8bYFpCfZb3xu8Njr4yrGIr+NFEzeD+m5vZQlnBbKKiaIgzXy/GotCHTCK0
3MSrmD9QEtvatXlaHSvXbSAwoPJeJHoesomtkg8WaSPKog3/sSbAZ79k80mSPjEM
s9mBkKJwt89Sp2sA5MdZxZJiY4rETAexacWCcm/duMT0Tud9X0v+XkKiPE7iyIeU
C9Ebm0X7aGvxie0RLvP+pNRgF8ar+u0h5oEN8n5ttDnHEa4aPOuIOmY0rLVQUMay
5oH50hZUYuI2wkGQ2UR8rdtpdd9qyFL2jFvwp/RgKYlD99yZGRSKUpFD3lLCkmrJ
AngFp+PABJ+WE367cOnZizwymgC3wQBD2PAMTR9c7OtROYaZXfvBKlV+cPLL7UWc
osWd7w2j357CF0a5fV2DtujZkejDkaTnlUMOttz24CDjVfgaCC1pSn6q/NFbfdFP
e3ZvgE3+0We7s0DmkssKfgM+qaKFB5YIJFQwnHDUlnyi8BHON3EiMLlgZSz/RAN4
7qSi+OxRJvPzNBXqGWOpNxHUEIZC/ww4AVqxl8YG+OI7ENldJzLrNnhroFbO/qRy
puE3F6M9HfJF++x69aJe29QJNzB4vcacxgETcTko8+AgVKVcwz8JgPx58lul4MVA
HOo+Zu2MwHHc6U4PMmAfEMgz6NBeLYx4ZvmzbUQ6/4oi/uDw/fkyToyvfD7Msu0n
VomIMXj36MfXShCbCDAO1U/pqxztpwEUPjgh3vmBb1Z7BU0uW7mBUXEsyyJf25Ub
zh16pMYl1oQ+28CDOcO6TMgH6+4yCWuSH8k7DkE/yy4FSdvmXpKbTYJeocIpK39s
nUDFlED0yEMNHpPMZXdo1OyQynxHV9+NpJ/T0/SVaf6w3LRQxk6WEzCsWzCxu00O
lnaVuqGUIDJx7zge+cssBjATOFcNBNwNI7Qc98Q2PEYbXBVQkr7QBoZMcrHCbyMw
2w8n0tvwLHulb1mUzBTgNq1D3XcdUe6cj/W50y1kieYJXU0iaC8sDEm+NwWhV3D3
WNLBEpGqiCquO0lp5yeOTYYSiYfvuQ9J2W6tAAUvyDaUnjNQz7CXBrQYctbYEqiF
3h4ctSMDdt92mp8f2dCIw9nWU8FkZnLt9igAi4iwemr339u8V5dZFEWF5gCa+O5m
PK2KUUZoRdsXlAbP3t92zpsWJgZaqg7vunzIvxHzio+k+bwvbKwEAcuONeN/eEHZ
8j4ikWDFV+xKS5gFLrUS9jLOCdInXQli4S7X7ZYf210w81k0kYH7H0BnDv+5kdVA
szMi+tWZQlYqfou5/Wnjjv9Hmw5I1KeO2xDLkZHwMsrEXxSqENAeqC69IbgoKGLS
8JaXDcGpu3Ziahyu/KhM9XBDE+wS81uTAuKs/OO1HuUEJonNin52QjoevvK1wHXy
2vmVmcxUYQftN258xWzBLB/yzs2/rjN7rCD3Ewyrem73V61TOvzI2/YWEsIZGJRx
qtcvqCHurXahMomDdeNU9HEQ7Woe4+JkVxwCmz/wtz4N3sWLs/XavunbqgC5NTDs
cFff2yzEQm3oa+UD50EHebKvTxhMArfws0Kzjh4wTPjrpycxVIJpC0zR/HTCQH1o
E6KMmOduV4/p3BSrlEN0Q+rrr8sQfiaqWQ2C2OeRpuo81CKjLXxtf4wnJBrpkeIq
AqNsnC4Qb5IKzoSPPrQ17dHl5cau+2OOtli6JGBH507zCfoomfKiCeeeeIPZQREX
u0W46tPCQnhtt6JIoA3O6SGCMiRvSWrOGfIBkCZ3Qg5gYZNwkdYjPjZNKN1DyT0s
UZJhbaJAJdDcBHVGR1zePnQzA5RKvkKUT4ZiWCxILtCCMdYizqA4Md8B0ie3apc0
bwGsw4WKq/3zXqvrwJf/63SgomtosrbnvY4ZuRVbnatapBNLtM6mGPJtR4LkZt/u
MSea1bGOR05QBpcetP9rx0XFSc/RaFI4Wv0ZsFYw2u8+IQTm8FYlcFghSUmvdi2G
jadmEI4jQvkCOoMHRNmJ8gZZIfYnp7hDXCDvXOxLZoMq9K/i0v8QlaffKJGTm7ra
lH1MVH4XSJF8xsv3O+6iUMwyLcyAMHLqY8ryAtisBnP9yEWZWjLqopaLYyTlmrrz
1WHSjE+ZIS1jd6OLROhmNOgPbjlk5K83MoN2IV5pJBQFwKto2u03Nl7ZoUnPf4eU
q+9No7JobQ/PDylXcPSQn9e4LbGSg9pcAgoZobXR8Ia8qQzloOtIT3H3c9ar/GD8
MekPwLNGezPQB29tIMY4G/Q7cD7KBFydcLSm249uSjV5Sw5TUhfAjSSnsc8sDVt0
NDmPB/NLQT/869jBKOlY2XxxKD38EjEU0jQQqatwXfIl4RTHsAtpntrl2CwhwxRR
q1AQNEOkO7LhTdw1AfVDmYTt1Rrf1nPUup1LlTJwGaWdn4PevPGg9b04mjywT487
+jXGRYJdCMH3gGjq1jEh0TzjD42nN+FYEYvJKie9Jc6a30dQMuWKv0tn5c126oNe
bDQYnUB+vKJhe14BuEiEc3kHTpLCwDqsVMcHnuLSRvbGmtBuurmkVrbSiuiZ/JJo
t3mRqzILrHGKmTA2ex+Yn7o+pR9PwOmCxlSmG56QYluQ6xewczdqVtSlFpEwCrkK
cDayegxUi/E8Qpm5TbFsPowh69e5tr9YDcpeBG2jwhuAp/e8421D4ON++4wChG58
a4HzOmcZf2frg7V6nc0psBNlDdwzbfFHuU0wXJBJ9rfeObnPPngxaPjsfDMOR/Kc
UdCsB7sTwtfpfvvAjQGfSwmGEu5lPhplZEhuhmFg0HTTlDOPMDi7ttMtsn8DKh96
dywzi8pVktM80t+fO5PbjtLtO11F6w8CcesIQ3OY+9tII4hX3aFNil6dIUcyjl6R
VAQJgzaQ6MC9ph1XSLl7NCuqqgh2FwNCtUDb1nSW1pH1zhYKGYs5jQPD/tYzA/XL
MPkloKLEsFNFwyjy8XJ6CAUeDzMe5NNhqnc1005JWLTfLFCd5UDBOLRTAQlLq5de
Opqf1MCfegyXx1l6k5Hj9IK9r9jXru2b5exryJ1vAwqPoiiEAE/4uXtM2IDFsun4
6aEfNZYGNu3w36hxwaApxahfQue8ZnPY88MsLMHutqYBpNu50GUuK6k4ZSSOR6h1
kOLe50Ex+4MVAIOCqGvMC47wJQBzCPg0tZ6L1ZrQh6J65Ngj+oxB+J4RsNcLFwLx
JBC7tRCSwEnpSNdXcy9YTv5XIS/rczaik7cceRttgqXBYOOrKffrpr+hG8sQgF/L
T0S5JHnCPf3be0kK+7V35GRGp92OHaVEQrX2TIYT5lIyCMqrRs7S4tM/04O0A/o2
fQpm1U+2wqPtVHR1sLcuKMcRZu4KlNSA/4f5mb9WL7kIRal+JgmswalOKn1XiG3u
IbO4QhFkyDMNtgyf0svdmQ55OmD+tGljm++dvsF7/UsPe8qUSXOLqfS0e1F1/XwG
rkJhhqb76iwcAmfXTbFfjGXRVMLJ/8HftGUssJqoUe0cdKU20e35e3lAPYZOVh/3
EpkxI5Isujb4MBpn4mXCMRUcfiosHhAM9CX/7FshsQSaHf1BtbGsvLCLXu2tl4Ik
7f9eU3jPwUk31yd7hgAHs51SxCrwEzuG2i2d/8F97RPX/lWvwAaLxSc4R3zEUPKf
nKGS7LkgeTJC11aJkc9nXg55XzhfI0apW2f0drjGxqZidWwWgFquLRxmthI9fli2
gnTVHP0MLxn4ls7Uw3cxzZtRNAZftLOYnhZYY3sM623tg1q/aKsowfi/li7nMiC1
+kQzb7kZF1V32mBnYRUdXT6/cHIRvqvIkISbFoRGFyfz/2F+WXRY7ze6ZiKLW7VM
6aSBkcLFI50r1cerQxDyTsWOyVEJbH6Ctlmw0XIl2gjxDJ8WDVqvoGCEesw7/7Mi
tzWnOuW2CsSTfsT3XHwt56gSMUTbg/sC/GdmgBGqa/FkY0bTQg/5ceA3X5bOtB01
OURsOYF9wqCiKZENwYMDvwtf1Nlm54P5trwzAHdYhsrrLPWQTpb5OyiYVU3A1j6y
dHOh87Jo+wUDLudYWAgUHbbfCq+MAGgCxuGa3vxr7vm6dPL7t7CUyzpmJDYouJfq
QdaRrC6G52VZfe8iDsRJzs9rVqMZMgyCE4usx61EIGscpuh9n6nzGLxdGWUXRps6
gwBbQcvR5qs0PKjjGKXMfSXweUfW/cC6+GzQg843v//kHNbfMwEL/JTFe7lj9H+v
VkNMXpNgjz9bQeIq553PhOR8uB5ZB9lDJrNnDoCpKUU+s5X+xpgwbxH8IvqTUIh2
+1jEBRs8etHpfWByrU4lz6iU5ydWIqqs3EfrSql2gJhG0vtH+HkgnC8xQVq/hNQY
1hxaBslPIoDtk7XuutG7Fv8fNCQTc1bRMvg5K+RJS10hBBbv5kLBkCSdijB8e99u
c5LefNaCjzJr072KgK8w5H6HlUqI7/nBYv8bdlKGvt2xqGjwMSsxVqtJXpR9KSte
/OEZ7SrR1qWoQ0H4IK4zJN5dHbix73VYWwOYkmb/67X9PnNxVrU3f8YJeu5NMlrR
o3HteIz3l1V+kEGP1HGOksGm+wP4lAZaQ7cbSr5J0X0xLA2U6TKCeRhlxU3nn1AU
rTjo70Ffx1+tNVzRzUmDFpyS+GXd4y9Sg2/OrIGBFRwbLjhfWHQVgrJu92uBHNgc
kp1ZVF434RysdgKnbVd0iCy73a0tjzx4/CjL5djBVshCR2oCLd1mT1/7BidQZH7+
APd/qKHn7o0v3pB67jan3F4IW1nPx2sy3Fci+KeZXjz9wX3o7M2jW1MjSgg2xKKM
ZXXVszy/cKy3MLjKZRgFnTqKE/B5/b6KfRgyVXWZd3g2u0R5k42MhCMQRfNx91xy
055EmdbVI9qMZTZvTJ4FrhS8Gl+y47iRw/o0958TkYBcw/0v1Gt1rEGaX7uBglb+
2tOvqvO1oOLlFWNlIgbR5HpbxiZzAEQ7idikr7W6gthnoplv3NSdwCHa14YUwq62
tjihrOzFWVaaAfBiU9FZDhWKwyuhBwO4HuYJQsNBZtV6ezivPm6leCzTmDCTzTXK
wHzFmmgxs86G+p5zigo0C+z4wEmo/3cn+ZUVka8qoL+NIcva/yFUII6BgTh6WacG
2hbYvdibOU7mUDYDnFUoyLxQG+qSNHc2urW+4Odfg+HWRB8dj2w+pX5U4M9JdEeg
nXTCY7aarTxepflert76CoOg55SP36stk8siXckJok0ZSjrAKJQeWOYWhaNxeT5D
p0HTL5IlrfCnQ+Ud01+3S8tH3VVNsesmQkenb84S4rL3N0boe9RjpVL6NkEwJCV+
dKoZ6N17xc2Xk+BE5Ae3qq7fRBBh+ts3v6lpU3zGv1myhCPTJ4K04za7phvpvOUS
vjvE2IFg/aRJjqmgcWXfVVuAuO5EK+WEuCTs/HgI45QAwge1VS+ykS9wG0t0nGUS
+ShyqvurEVaf2e0yQzVO1w1/AjeYTIk+Z3dXk75OIzLNq5PV5qJVJ7y9c26xOwvX
KwSmC3nUuP1wXsL9g6u3CI2EP3BPp1s0xElp9fe9KqX290eNOR8C7vy5H59jCwzK
bo6iHf3WE14NVCepAQ1AZ1ME0QLIX2iHQaE3XQsviIUUM5GW0zABITe0oqRCWAdn
rAq0Rc0SiHlEjbP7Xwgq3x/MwyzxlS1Y+d2dahGefhVt+SU9tK7FbC0/Tp0oWuV4
pmiv9qzYCo2kp3nEtKJgbPF7WjlQpZ86oufUD6MO2MnObcKJeDIr07mAZx361v50
hTyo8AudoWyyk6ZiBKS6RHo+lOVR2/oZsLENsCEXZeGgaE2Z31p6RevONHFQ+Qrl
qnkgO/pu1kH1ec9tJ78eciklwTHme5h7VRSh32LNhVGfp0W5/fEBAp0aa+dzP7dE
XO+/wHOhOxaBeDlNBeq5C+QH5ydK3vsqVZ3/7B8HIuC4Vzycf9DpWs/cf8JhFxLu
gMWE2jvvr8Ft2WqjW/fLrx/CZoTlR2zy+J8MQGnCVr47t5Smo2K1w2g6KOhSkNAe
TNdeaGnBekxXgTB5/IL8MxLn1Be1D6EhJKyV0UvONNznIDFrMSFrG5KC695XyehR
kh1Z299PdxcmAHvg03BCChmrsotHiyp1Xk1DTDIk72hDQRUQm36T3q+VldalVe35
1jx2UPIW+2mGsZx6BC/blZF47xqkwNJuixcSxtxWz+5Tjx7Gbbz2F0hQqOMVZ/qL
N0J5zqz5zE+b5csfMfAuRxbYKC7yqiXC+Cgmp5saIDjp8vF9qt6NWhAbuSGph1ZK
SnDcshn+pz0J7fMqW6J45Xq4EfBFMDG+PGzQqdKbjeeCOQ6pUuVn3RuaVybAHGsZ
yZneDdTC7BQmS83xTTXgJcgO6EmxBsabHXJmhBQoA3hnxan7i0z+5SP9/Sefgs0f
BBT0Ytg/iqqufvp1vkOKf7BethPtxNmdf1q7T1LptwGWhiA8E+MiO/SbK7f+b37y
NA5wew07Q0tAiOFwjfh57g7rEurLupx0rRbaHB8874nI8Do5Nv5jpsZFJFo9ibux
jEFKMb+6cr4pJZiQvKyzUaCh7z1ogn87h1YeLi0JsL3a/Bs57EVHBIR7cpAukV11
keZS2qMk5Z8gP6Pff7LouujbSIRC1P+oCXXfFQ+4GHrdJBgqR5LzYq4HFUZQprS7
tIHXfJG3D8Uyo21ql/GJm0KcDc/b4aKr+Y8nkF8Tpo+2VrHRMLCysaZ/6tPGn5Kx
NRhtsoJObvZeBEeiU+Xt/7Tl8BXfpSBcaemdSNkLvRqskYbKy9eFK7JZw3/EYUAx
nX3yIY5KYnZHNd+L6vkcCyz5gMZnhLUbjlvL6AgFJkRqxpK5O2fClE3MyvkKlvTX
OQWDznXq4B173EsZ8msqljvi596Lu1sqSv3cJm1cMICz35STokRurUqjL0/skqbj
utG8igvZ7OpOgqJ9jsDwhpGyeWflEV2Vj1BL7LFIz8/g0hbZw+46z1ZD+zSP8WBV
NzE3281/iWQVax4b1zcoBANJVHto1lvyMJNtQvZmFNA1NX+x7HbGfx0iGD9c8cRG
Zm5uAoeE+CgIQ25bZkGwHMwBEFsHOVBnZMsf6hHd/2VipC/7dXBQegIqsDt2kXn+
b/S2vh/6Jh8mgLLg83NSrk5Cn6uTmaPC5SIdOoy63Jy4iryECH4jYEiG2hC3k7H1
D5WR9FUrBiz1rCjt8PExDz+r1YxSdGHfrC4mKUjCbnQRUoDm2BwDo91dSeje1vgX
F8Dr+D7dxZ0LBHAOCZrmUNuqWG8Ih8+KgGZ2WO9FNcEqhoZ59MD2P2YmXjRdNFyx
AIIlJwek0UTkK2arkvDHxnFZVqBSkvwrU37U1BYswtS3J2mzXNoUGEY64t0NEQ2E
3m7b+QzarixhFYv8ATOO+pgy09m2CtfHRqzje7Z0gwOJwYn0eziGHXsZ1KDjj/li
Yi69wfE0HTAVs1Jd4gDcQWzLe069m7BNMXJ3MLK71eckrW8JDVOYhELg3EkKPp0z
3Fx+m/n/pK6mk2w0CCKlL1Xwid1nAr1NSpAxZBnHGzHMN9YV/SmSdQux62cYrSLA
F0c3FpogbfEz3tJmyAA8twDNnT3zjeYkBVGA4LUi5SZ1BzSqqtf34I0Y1y6DdKLG
CZibTTXKcENexRqCz4IgTe163iF9kjPCadrBTpRKEdsTCtDOA/L8Y0WicKGXXaCS
1iIlRlPV1d/GfQbvjXvQon9YVXkllR0Xz1X1U+zZnjMvCmbm4UfIFdmQwttmiM+O
KuaHe/P48Frj+U9Plsk+FmMiyoCKrZnq+sVibJ6RUDRq3M42nwvobX2gJcX2c7Nd
tqqFXfEHmFdgmNzjVDB29zQD7TRZKO/+jWHfInyhRrVbTv2HNAVZfSVqcm2Vpl18
oilhMQi1TPeipfqKDqVkfozXCvfW7PGX2C52PhPqCEYewCqRWBmYCaLnu5uwHAC9
mHVBYp3o3aTZxGaWxIhx0tPeQgwWfsRC6iRNnghEKScjmUXDoakuBK6yDqsPVQfn
XKWGMDjYFjf5DYUAjP5GCLFkAOGByOShC1RhxTGLg5LiAp+2V/tpi9azwl04u6Kl
MhDqxyGcqlBdFs01nanYHNUnTdasCP2lmkbeHA3VmsBkKGQvGXrykeRkkMMx7M+o
Ppkx+pctNxQUS6CIHYn90roICOgI6OVqWx77y/cSRkXTwuz/L7pjAJh+P0rnsulJ
0eT0q5u7DA8BpBwj3CqYhtlavnfNEzGLs/g/RbWxbEBhb8eXqtLUp6sFg03w8wjM
xUrIVG2b3b706ZE6YWn/MeUvq+zPzOCCrXVmTIjFYdoTDP8VOJ1rsGDjtFlhgrUl
tEGra4IHJB+MH0Ugr95qi+Hlb0rb9pv7rUmrpHsZsW+hgv2hRYOPUFuNt9k9icVg
BaDK7FhX0HkBBBL7YW2pPv5kTgG4ODR4l3Kuz56tlIo53ojD0LZRRMFn9FOXbdSm
f4rwBTZjagh3JKAAXg79l/vOQWVJGhKT+2t5gmzYoQXVUMbW3YiDSGP6h47Y+CgS
wtg5ZfZg0jLmJabs0n8o3T0s1xuXbgxjAwL3Do2V//S/xl9aG1aBKu97fOnH+19F
fPDI+wwyqGEKqdg8zeguzhW/u72PAMQDEqyFciEbHcced9lnoyO2X7UQq+NMbom0
IJ9x1qkL0bJv7Xi4TunUPK7bNb3M3wyYRZSsA364lBkthNDzNkDpchsGYvnchrL/
OeL3w+pIAjq5JBYlmTaAMwOs5azKrG0ePo8Nm/5/5GV5iGCVwixzQsvdoIx1oOlp
AJ1LStrDPFh6w/NWGviUf9To9lZfaI97tbHB3Nrn5X6CUAK8XgDsyyEDyZvbc+hI
MHQgQzXxBCqmzzCbHEtOkRVMrgxLzPtSAnVWHGZ+MTmBVpRY2q4kw/eCynnltjT3
Pcdx+nLppqpcJg9mDwqQB0IYBQwix5PHDHAn1L+r6xaphIEGUeisu5LtAwRIULM0
fLqnNPim4uQito+b2psVCXOE/c8fjrpWFbqPexN1bVL9MtH/o14JXV7uiLPtzUYA
xI9A3nnyUtF0qe8mtOAD4XC5qcmWnu6jddvkXTMTWpuQF8X4ar+fPFkD1j0dlQx/
DIE7bZWzSTcyr+uAq4Z64cDr+o/hReLthPHWJf1lhZaSh5qIbWDK/fFnzCTmf4DT
VMoUaPIaiALW68dRNMk3qxNW8oUFsm60o60QXRJz3I3sLesS6aQSvrLpVzUn8kPS
vCntFaKvJ9g3ekfGqXrTbb6R2O8Bjeznfw16nytv+Nb2+t59bYLoCbMHqJPovPNZ
wV/Qiiy0OlvvbFNkbpPDfhfgdFFHvwHt3gQZDmP0p+VwqkdI4WwWXu4vcKOBCdzV
+7fZLFWERMIy9eM5uaqQXxNy4zl1tSE1g2TO+gBo+9+pUrOqc/7yfX4wcVHhNKpj
GXsa5dLhu53W1xTNlEWk7wpORq7PT03Ot4e+846d6ZnYobJn+UvaDyUkTUVKvymR
9h02OkxhM/Pw0E5/ZapSSDGHTy01WP0YHCXai9o5uVtlhDdCVVQXOWzHXG+PJW29
/+lkPaC25HGZJYqKbtVzKH1lSsA/syENW6u25Jqi2XA9LneZxmnvwPi+Q78bXNiS
9QEkJF9YkUfSHg/3/5TjxsJJEbyiD8fn4vmxVMhWoK3nlCfi/Q/TgD0mfFEktkEC
nM8D2Cke9UxR4luDKBmQdbrNXKqSS7KpcypzkLsAhir8Ox0+B9fLvyrAkK9sLkd2
W1Ein+cYrWyBdv64IVLBzuQp96/bJLpZhkxwQcIDLCDKtMmss6QOquNCjkqY45L1
/nzhlKGYcrk4m7aPkUaHMSxVXf7cgSAgKNmuYpmqd/iV+mvSCZr4D6OtVpXwuymf
T7AP+wcdInMg6Er0PTAu9W+FjYYuEnHnLFI0Br0tZJARHYTeyNJq6eJhcUvz+YK3
OvvLnwGuo8AnQ1KSakggyHBgcfgdGWe4jZsbaD5qV4c8MxNrwRIKAa+l5rfBIkf+
5dIWZ1QuDduvDGgQr1nE0Rsau6Nr6X1xCg/rEZao+m2UYmO8lU2GXufEXATmGA/h
mAN0VfaYTQdt78GBY5sWjfZnbD7m5C2LbZajJJbqqxwvAukriHW1RleeY0NMxCPB
RiMUnxg0hIDejAskRwUA/lU7DGiU8YwqqDDRjcorl89xfZrLraG4dMptFIPMGTn2
SxJUlpaC/wneyOzp8yB/WQcMmOXaSUw+TRNi+JZ7AiN7zTgHbu+ZonrsNUQgHUcM
k992yUEy2Mb32yAvBgT2ZYLPgBfL9jb6JbjEaa9jjnNkwFRJkQ+KrAxZ5NuwVe1/
qLAijvek89U4Wb7dsyG+wzeJSmmAYHlnasi0XMJlVtYA4cRBScmqNk9eHwhSBuWO
Dp7bcGbVJCIiw8AVCMn2SpPnlFMmMIqSO7D3t5MTifiMnbfN2MTgFSSDTPqtenUX
lh7vbhRsNyg7S7KEMfs+7mof0M7Q24mvBor5q9+wFwf2F/bcLuyVXA0kUnnj5tYR
D5pGn9wLMZC4mr3jE7OgPLlvsKsvX3CgK2uxD+U1XIfSrySQ3UPbB1xYtlbFEKV/
hcBjQZiyTXzPtqGnr1ebTWTA75ju1qdreZQ4JAFZz8LmscWNwfwGiQLiu2nwhdpB
nGX6FDuICBJYsWH1k8JbUl6MLhG7qPDV5afZ+6/hNPbBLI+MkxTFWr78EzzV/ex8
+661I0Xft7n5WjRpEG0kstVF4lNssSJOtvIxnKLe5ThSn7zA4zxcvURNdXzdNFHr
iOh+oxB8scC3x/hg4GeRlXEgu6kxUENPm85uuGsO5ogA/BKpC8flvUSwLPnUqnyR
iiCPepVufsN3xGMsJrH/Tzpf4mvOkt4NPKkEEx/ZWlE+xFiO8+6KGRtxDotWzBBP
uQ2L0h5ifr1XdpAATHvSQI5iLdm0DmMNhmnJULENsgT41pwXYuikNxgnHXZf6uXE
+ZwdG1bumfh9uCR55Yvp3i0uUq80jsiokBWoKxqSRnHFTmSqHPesRmx6A2LR+FbM
wzQs9E1XSwT+yEYUBTymhdlFWp2EtPP/As4w2VHn5y1JzVhbEjUo4/r2HACgLkkM
zjZfG5PvMXSc/QBfRFXAt514cRLdgRXQaufP1EHKP9yF8eHnBez7iSoPK6fS9yEm
dOGnp/q+2aBz+9yv4zvFDpyo8T0Z4KrCoIC+cUph1nrf5rFjj1apXpnBEZQo2zlR
6Rc1JM/Xkv39lR8TEp70NP3mmT+eBHIFg2oZzHvVLyp5dIcSmTIkRScevzGqBAJa
3aVlLEztXk7khzWhPDHNtfBR4fvN2IRxt1Y9llheKAiB3HqJU3uKrPFOsFJNkbXs
tpzCk/9W+/NlpkCqQPdoKbyGITFSbThChAd34JO9AiGQWaDe13Z6Pi1oSG4xkCk1
Oh/SsQVdW7PfdQiAzGmrSQTjXOGTs/EwjW4b2cGHqP7aGrlY9nHlGClsYGuwnvS8
jvNdWlA5EV4us2d2nuOLAtpF31y7tLgZ1lxvPsMoylDXPGpSYtkuVmas0+JufEOe
UDrtUYYfT0YgQr2MJop8kBGHus3fhEpAs2JxAfRK7KdXj0sbF08h3oZhHQOIdevx
eC5S7kW+DWvgaICD/Qm7krXpyonfmnOOFe0FiiNhWrpra48GWg6gDkDnmEaxHOLZ
6g8nzsqd3XNLQAmyzD9nsuqI5AMusxrCjJuMIOTJU7MUJbTjtketcJDjPSTs6bVJ
TtYCyp0JNHXc3dHe3JYC068lW7+124X67VPHxgmH802Ivq3WBWan0v0nYe6YrDWN
epTjDuwDNZM3bZrIZAR9g0mKwHhWcx3q7+g5IyqXl6tAcjaZkIquMZnIKjZkJwhE
X5srxdqZ7ky520sQZOyhZmVJqTnQezNOCo8TTU2vv3ucAlUr+Tyk4C4QuIyp87r+
Q13Rqfy1DSmKYdpqAK6YHI5gs/jNaoY1D5R0k6icY6XlKhn0B6PhBwzEaRNzNkwq
mjM+lUxuUITdWfk4HhKWwkzYCGamhlIpAbfRcrZiBYOLT9Ayf7PHuf8MoZgdEPU/
KgjWkm/zOWxhoPBrjURwFR/S0z/PmZL+rb0MtuFxC+0Bdo7CWn/r7eJekNRbz0Pz
HugTdt4rAzUBpDuJjxNqKRIaUm/BKmMt2ULu+/sfhehPGkoKoH7A07If44lLEG97
5EmB/ydXXGh90iDavXO0O1JwuO5EEOwXjn20GFX/8gdV5y3WFqqBfPGNoCG5DMzq
bgFACnfjAwSUJMcjjRivRmvxvdLiLPajh9axmr+9BY8z1MXsy0NPxpLLJyNlQnX+
Sb3OYUWfxYJXObeF1xYUBNgl2BR7tK2rFuUtRRWMjVgATxLwZvV0kUCBlCjHJMh7
a9YTSyQmbl4brhVbEM4xAOrk2XgpARDqrqMbhYXk2PuNcutbzsh63wrrzXPLwpXQ
ZGMwULdeL//jvY0wNssllzu4Kdc9fNxNa3PQlrj0uFMuauqCbu36o+glInO6cDlc
Zt8mOlitjFdfGtnT5IpM/SBt7QFsA12IhLjdjcy5kmkh+962jejQvWsKxWRZ87kC
UsTYLF1IiSYKGjYYX4Iy65OLmJSKyMWq5esxsClIoZV4V7JaAfCrEIG/NbbkgdGr
qeqBXe+NyLE1G6jV14QQQRCkIu/BUbxLTxG4RIFzVTp3HSJuSnJzCbkWV9xbCGau
HGtkLO1ApOh1sJPnDeeD2C/HrazvfwKtBbzB5fmwmo4oOrdpu6OLjRAI8DCous3Z
YP92FpFvRqZ5+t3gVI8wGBDUUnB1Le3QgCHSM2PCUAiE/tgBwsPtXQHL+31TvVuZ
CKFTHIlWyzm3QadqLi3R//aTsZ6gH0QwsQo21yv+HAjhQ2YZHz4npQ7p/Pq/rKol
jIJYxCCM/1onzkFvPjPPJqaTVA42OyVEol32thZHbKEVlx2H8RbEBwLSx/vvPbyo
XDIqtv0cKWt0mo64vO/gJP9SEQ6DzAo2ksFXpPFADC8Xt2NhJeSpD90Vz1SrDMGw
oR0wA88A579kQn4HFyOGUPeOCsp36waVnmRzlv8B9escfmbT0qth66teHO9ckXV3
pZ9jYMn2qcJ9VWUm+8G6eEudbAQoZm5CugdahLMpWC/+00Z46dYcdFza7L+o9WaN
U6yEJ2WmAkuvxu4PPHWmlCoa7PyS6Yi0mPxiT2uxD7943TVgzKtiZIaBymFjIO2k
RFMEvhzXd0UkrZq4tajW54/ox/pVXZ9aiHY2BlhGjtTOH187KwmVV65tw0ejlUXL
jEB1k5sUkq8pW6i1cS501f08xr4OJTd9wzgCVd6/qOrV+tkEbDrosDVCqM0M303l
CSvlWTGl5aA5qCWjBeuuLTcdnBPW9U4dyr6xiF5MDCpFpjXji3V2BuWSVVie0P6D
XjuUrlfPLDOsTEWvccVt8K7bdmgggRrnqKNJ6PUlVB5G4JKf5GGA+S8fUxLcXrQo
k2yxPhls+ZpwQ+c39NdfFXQ1ZXoEJKgrjt1LCBY/VOvdY2wWW/KsmXIobKxNNzDb
78F9n30MoBaD7Bf1/o4m5xYm5P1FYAlfCOYBPCGZ1q/ZFbjY/RxPRLXwDIpglb8w
qoVxGc1PQ32+5l/HzgY4kaNy0AuuplNwBc8ScabUip++DvqHxEpgbOXmbhLP8Vh3
7i3SPzqK0xuNTRcCzyZaOichaAviXKD8VcHxsh3wr9OWK7PGlHJ7EKInjEsyJ3+t
r8WpO2OzREUWlg2tV3/XHTva8kTS+B3afT8RI3fnbxXJ6eQQyXRD3z7hjEWMsgUL
HwHpocpKUg6RPK1BXxvDpz/v7EO1uB60ErhFibO+0WUiJrGQzWSg4KbZsO1gzaPP
RzftHg4Z+J+MUScPrCflcctuNu/m+pemc0avOQ2Wv6F2qvxgqk4AaURN8hkRtJud
Ve12COAaPnEeF2jJFLbW98d3VfH9LCt+enLRIaWfZpc0Vr0VScKRVTmgcfyt3GPZ
llA/rHOsFsRoYkV9whjUUKvKiHh0UlTyU0DdJq2PcmUbBQamDMan02yFlx870y43
Tvny48yaJq1L3q64zwiZCEgI7ZXdU6ADsBH6jwXEHMFDFuMMUXqbOXWOSHzrd368
VIK05KfNAH03majWx7XTM8oNftEwejLTQttIbCK0JKcm/V/4Z+8SobMPDl0d9XeY
dq1OssV0FO6rA7Cn4sz8hS2YGsDH2mzGZ68wA3rOTEbjLTAbZq0pV5MXpyHgygGZ
cRx0Zw7n/QMgjKBoVu5PAUtwfYZFfrhpbkc6QAg2KwYTBcINsJLBckKG4OtbF5jI
X+Ah5l/NneQYHXMi2vMGpY8Jzy/4XngphUTY4cN4i9QhjDatWovog+cnHWmFeqfE
Zm46gYuEev/rdcBI+EDEZX8cHlYESdMFY/10GBblwW8fBDfc/LiyMxcvz2L7GEM8
/uzGtsKx/WiDlRSyHJls2o/gRIlYOlaLniGbQQksgJWTENy7RT0PevZSJcOLe2wG
mCjwvcugarZKTtdeNPqbullpK5oqJ+I4H8j+qqsPa+4T1AHBju+hjg3JomT+hPQJ
+aB/Od13Mfj2NltlZB7H0GlJVI2JIocW6h5tIBGmeEAS0zXAYuLMWO0AnVv0CIZH
PsZkFuetexgzNpyBhCnD/V/EpaNoZMiofTCTBqQTRi283zsiHUCFKhvRdOKBXuEB
KmFm1kdk53xU1wlmJt8fUN3yp2l6o/1upFW6Z80tXrjh7jUwfRSiLEPPJym2moum
QzGyzuPpgC2N3grb17PKp4bnuPfsWvMNVtaT33Hd5BEZywYFMViGwFeGy44wSwZX
WP+Hdxp0WOEfdUWm6HhSz/Xvz7F5t1IWnVzgmLg6g6JKPYMDWlwKQ7JBh0YzC37k
h3jB5T8MK4PKUmDXcA/4AC9k6nYkMBbNFABqUXCdmraSKCC6Slr7Qzl3V7f3Jhoe
LbsiEezGN5K+vkz93qcpAV1P6F5XiQujXDb317U/03k/wUpXlIVh8KbJIlJhBlQP
oWou5ljhxYHNMw/X0/kmsm0kynhDFY+dusUnTBWPfLOpet6OrTwL4ZKpoPgJIBlD
syFOIG++b4QfHYQ8YEBi7IQhPIHKqMzL30vlGeKtUpb/+VELRyDNLy3lJFJ2/1M/
uBgaSaDnHtId3ipZZWz9vSKZ2FAuq3tRAGL8Q5SFMH2ziayJNawmiBGS3OHQ4vtV
mjTg6UD4YELCTfKyQtuFWCDZYkQ9onSFP9WCs23zvBElYWmkXO0LSG0kLvzvHAmX
BhncMih4V8VlE5QwQqcIUdpu+4swhkJdCmnM6uyTa6rwNQiUIgTW1c4aNrLLaYIA
5EO7waanYiQVFMp324pHcP/BWWW2MMSG39XZbyRaJPm2172GGaBWkHjtDpDVQiFP
JU1gECyNwG0MvMOMMTqP1h7Idfww5qNgVWnozSFvyiBYIPFt3Lf0DFdLoTsEuxc0
7NRHB0KqJlpkQyKdDoluLndqe6AL6nkW5hpG4bUdECRZEYWU5JT+gFR1GeioOhvX
OyReMXvoAiLl2U4IBrBW2IpZWTaNc2ljMbuVerVS4CLnY3Eu7D+DKReBtPOKH58A
NMP5DkR4Cixe2VB2SSwg3eCD4LzJ2s6zlkFklQOfqbt+Wm9a5o+v29/H+MSjaBPG
B76uhCROjH7DKFpV4pWQrxsgWaJzt3b04psIXTtzjxCDNnQVberPfkybJhNedtBe
ZQPsXJRFjKBe/ILqwVSZ+hTQHjBQ43qU6neVh/mu2RngQn71kyV9FFknSl+1hInE
n/UfPhNTx/6OKemPDk+irp6Yp05sECX8sYaz+waLtQiAaxB3ItXdn/s9CrsEbpiY
rGNS6BuVMG88NPCfay+U1ki3X8N1NsMIKRXEYt5gjRHnWf+KH4pXzb3d0a3pW7+F
Gn7OmCeA9gGAAGXUM5aJTY/XIYzTwrz9MGAyTvZ/LJjcQ4F4aon+3ga6fQV1Dyc3
GBOEo1FUqh1ZdVv0Em8bepxo0WVnuAbJNNGBcJjqHkJpK/gcBZlzl5naqNEZ8AVZ
Ph5QabKM94/PoGsjjcDMblLdlb+RURfOha1F927YC3a85jlJNPISL7ul67YqFGmV
qrja7cf44pXftkBPOYYzl76Mzq8e490PK5HHURTWNMkO13nEUc5FaBtifHv51tKO
38Z6Xwd/vgvruO3lkLOer6XYWjQU+fK0fFC6n7aVu3pUHVBskjO3VXWju2J1iEzw
6wFdr8NmEi8xtF04F/FMmE2+s3zHPbNFFWkPbF0G+sY/Eok97yVElCrc77rc97xs
0DUE6VGDENcWoQc/ECpkIUIJZXAAQRcKu05X/CHrk9joFBURqpmUETA/qUy815jx
ao+RSTReBAOyFJEy4RjHVgWNTkd1Ekw0fMvE4FQlPTDAcWw5YRTMxz//TWrQtItm
FMPeCvpDh/hG25dEZZrTLGmZr+nMAFND1Q/xSqWwllTf2hoanKAJCiOmNk8gpmdV
UsSXC17ODs7nQmPDTLWHGk7rBaRwxQFd3YRQG0F8W/ykGxnm4TsCp+lPwmp6TmDg
zs5+gE0gRKCZ7LBu8CuqvRrcYe4+XVxKp1JzNUB/eWKQCtQG24z6ztNdPN6+DU9c
iSvFuJ0Xclxa5O7NdzR0KpPEhW7dspL06qHROWBji9vKk9l1d8QI/zpM0SIGr8RG
1n3WcPCNwp/W0o7YoYWtBaJjeWRwbFrIsJh15l4ZQPz/Z+Wp2uu3aUdMJd61GpNK
CjA0k2guRxeKGeCSotxGH11j+XgJ5Odl0A1+Sdq5qbV5+ke4gy/tot3Nuu3/Sy8m
eIino0oI4KQPJUkThbUjyQBL6BAFhIxWqpnna+mS6aXtKR2MyVonsbCUn164nmMj
cpsi+qwANxTQJtMai95IV7Yu2hjK7d01k/NtzdGGeNisaWXDL3xKldyinOXH2XaN
WmfEPbtH6tBd6wGPniPJ5u57JB6/zoFJR2QiS+rnjD3U9qLy0+inPBK0DkvZmOLa
0SKCk1KUTWVx7M7F9lFeVaAboHGXWjKz+zKaGbfpZGCA37+WUf6EHQ2sRPknMq7O
Mxg21qbP9SrIHl1nJBcjXKm+R5+g88U0PUIpvWiCwsWj2Emsh2R0wRvrrOBq77IN
fbeypeqM6mBnhuqcRMqWh9Rd45enlbxCzIBG16fYibu1qX3Ll0lVvb/wgxb8duDM
ZW+ls3Mz47hTP1O6r9h8UvFU3/RencaT5oPQ6K/JOc2G+5QGcVexAeYBhkYg6A/N
VqjhuBEwOPJdmhTXXKeWIVRspxxGYcXI7XX6s4yY/RXkqHxiQEtZtz6H879hxv32
XULgDxl8R6AzvosiR0xc+oqsW86pwa43jIabkuHsiq8rGu05LiJNKdNNNVHQveCV
P8/mwQLd2mb6FAzK1TqkaxZaO0jsKH6+amJJZsxdlEjyobcv8YKheeZ8sBg1SvI5
MdB5ATJUV1bfQ5Jsg1hQWkBqbk4qjBpKcmeB8lRV1fDLgOUkWc8QzaiUxyV4rAXS
nGc8Dg5qQb2UYc6yN7k+D6f09cgHC5m7FiHK/WfsjxhbV9b3xycMxtJ7240tHQTM
GkH5eu4WL9z1ueGtppFRmr01hYLxlcURSsPnBRv/zAcIyz9dt0gE/2llW1TW0gCY
j2fNakNgOnRcrD5oI/BczhTUjUgEDRgAMNo1b9BVWUL9mzPTJ5k6ZxK8JwxTmgh0
OjIWOiLIYX+Ec9/10q8ILVxnpvGQGpwHA4Vr82nL2+wCnH5kFKmjrNhKoMN+Cwky
6XGUoi1iXSWtMDdU+hEmj2lcEMcfUPxJoixFKPjY65sgP+3rlozjVFeaHSQET8yX
GbKe0x6lZNbG4YropI1XV9oixxcV7h5HGQDijrg23n1FJ5gdLJhW4yqWRSJDSjlN
eYj3pgt1Br0YN6EnHEiuQBJ4mDGxKkvmH7IQ7bKzqTMTKqGrLRBKrQZdznsC3Dt5
cCyy/pWxHEgmbDVjcu+dy7Er86Gnt38DHgPkWGmZE5UWrBjypqJlsPSaWv218K2W
0pe5lz4ipidra8D9KKqThFLOMKaIsQLHjIdqngDp7LJfIqNYgNDa+RCuZOPIdpJd
FQbC1B0UADB5Rlv3Qp4bi2g0ieHw1a1IEtmwpu5r9iROOoSgS05tUWp1RgcumYoF
48wijBJD5i3IMGhrBOegtLhnO+G8ayNfQu+m6Jsds2OfywkdbQge96Gj7sxizoIL
c0kMPUkvanZS1h/WbSgrUsJp/YsQ3v3QImsljnhYmBjlwyGyRgYuqD7TRBYdHVPN
WAvleOyRc3exB7Yk402Lwt2eYGS9PisuRXeRscjWDUDxS2vte+mIOuPpSdXqdOda
k4kSxSRt853tJ48wvSO9UqEcMoo3xVNxCzEyy4OrsZScsHIypCIirQsKdSfKB1G/
K67iBC0Nvz8IzWD9H0HWB8vmR3z6OHDho4X1WI279E9vci5Swm25AJzhN7cqGT6E
0C11+iA+x2ieblFsclU3Xj4BQTuVRrWm9DQxIiU0sPO/XOALKJhc3QErSq26beOc
dM59fMmwt9ohyJBW9PTe/HWNJ0k++IAKnQyHBe9lD8crRqj2yz/77nBtuZTsuna+
JsrToKXlmbBPdh+irZOL3woyfvQW6ckC0V7RSrfH3CUyWlPXV8g9AsC3kiXjOYkZ
f673M+47rSKwuQlHWQD4Hx19GX1K8qhks8dsswMBP4nVW6VW2OMbtRJhT5z4zPrJ
EDJ0TZ4xmsZSLdFohVd8mnwZDDYlVAC78CIU1ra+jVkY71AI6wsvEbaWMiz/5P+t
+PXB1haOahoBPJTZtMZyMnnuekf7Ne2Kv4ce7UIn3bDgLXKA76IOGVFOheQ+IkPj
08dsTImwOiQcYZalojXwHWR4ZoFKJvtQCaZZ5nD/nP/FzpXHwhr6MBXzLmRgbQz7
3MwPV2m4CTp1+W03JLMpIhj3SHdwfXDaf2X3qMbllKx2uqe7vIbV6zi+l6K62s8y
CCmoE7cAxiCZ6DMAlpZeQqhaPR4tKK5q/KVtSi1Se4KZ61IL6M1HqSZn2mmAxY6H
4SMnDK1P49UHWDwQiSxc0Yz8ayO8xvrbwgZgOpPJpxitC2aNMWIOPkyoZW6mWKYS
7KD/kzFh1ZTqgDYjKePNwh8t9cDkP1L4x2S9IfMp+Zez6q4DHpwxtKduwYFVTnpc
3Tf5mvahbGSaY8uuCysDdPjbyHhMEucOJIftblXcVO+SXISA7sl5OoysVEvDkqJC
ANn1BiErC15Gdt0afSgWoaccLqfPZJLleeTfeXZwVLCQgier90tDqF+sqt8YYIbR
9rHJF+DKI4He6N94v+daLQcSj6Cia2pwHjhIssVtlisfEun/Q0JELffdTu/u1wrw
I8ATjE88N1sWiECRp8VhWO0l/eyFenRtayC9ObNvtaKlmDjtD0XwOCtZWZwJTLag
H0ij1d/JD+X9k/QXtzRgFxUEbf+oLMr0s3Cwm1cyFvUrKlhmDFC85v2BH27TGM5l
oFxzJJpBGaD3Zst1S+BvA5GUt/YCoPRd2C597K6uCGWunNlyYw3pl7GpbomGsNwu
nmbevXmraMcLeGiftsO+DRuumllaQwzrsxuUKst6xU7QaupDg4HTLcEUXo74/28O
PTH9zMAIqtgh7IF2oflt0bmJkTCDLbMONnWlIrsHalOmIVYG/bZtHbvkZAj8HtlA
SQSorxp4e3MNrmMwraGRtFtJC0WBy4i3vh3ZgIpoFlGMgjbW2FlE90G3pp9c21eA
lyIbEKbm3Q3j46+K/S/c0TZkGqxKNbdox5y5dNYoSaFsSz9XWW7GhewViL+JvIoN
G1/8dDsxyMaj6WbPjkfy3G37bBH2HinHPDGela05zCHO1V7IThrphiJHVThNSQfJ
x/WEJdR8JSUfHNam7XbkukamdyjtZ6lY7FKR/a9cE1FmUPHab1ulteeCBvisTvTa
hD1eYnRdT8fFwWkLZnrBGroiqqrdO+CViUoAd09OsIDDFb3z/RMLTttUm56sl+s1
+Ins+P5X+9x7tyXAcv8LZZT+GOqSCEkmSj8JxWd9duN3nn0tTKE46qDLbOiwdAwn
r0Qapnd0qZIeXm1nqxh1+h2WtWUyKcc/G2t2mO/AUB/fZqEFOgTcuQTlkEGwshBm
T9FjLCPL/3m9iiAobWfSG2uTm/sT4lGfFo0aLXh+lbhbf9TXSG12FTY0TuRmh/yu
vjrVNLVk4OHqrH93t5fLcKOO4twGZ/rD7IG/pcllEZB+2+OeCFwzkddJfSkmHx4k
TypbVMzc28uzhKYu3hgfNOWSfeJ/FaIWYGharSniTdzlYPcxT06wFOxtyw5bK7O6
RtDiL+rS14PukxSiIAvwMCcDJBavtiszsAK7ufbE+46/lUdTRP6ETUm9JS0IDEe3
SrtSIrprtfY7cIfJj4YVeMZUteYw6Hx0QW5LfLZjhZGWkeQxhDECZqr8BU14HSb1
Q//gTLMPWzfh489FbU9dA3EJjR9UO9tGsG0pCTjhWWSQGri5FOkX60+kYnL9Yfp7
ufHn9GPcn+WkiyguVdHpdKz17TpxI75SpAawZRNMEj0RLIMkhjjHD60jLRrkzFHA
K+HXt6lCtwl6VG5klxmzxvxaekE5f9f1+udnYVjckw1AVPAXDoq9uuXwO/y6H90t
aUvxMTcm2DE4U31ZI+GiP98LqCbWJ08RBWf+jGplMJr4jHqAHb1rhPgl/q9oRpbR
hFCP/8DvxCXcdkTdq2rvwXhmQJhx+L0gk9wiqremCFeMgnaVdfALe7+1dOmGcFs0
16ryYqjKIoK1Ui18Q3AW3gr5PAD/tI6gsl0qyVZjBTDpyjwheq5zFMahF5bxVtOs
h1jpzn2dc89093yEIefToqc0K+v2ssd9T4Abl/8edZuI6kHfhLCAdBg5wbjkH68k
6QYlL8MdgFsvGe1sxxzXwdsnr6iS3bR4i8rfbaKnsB9TZUXgYb7/pkraMozvMF3K
H7qKb5wW+hPgby+seZrdmuKIXp/AKuYD0RRO5MYYURk+GSye8fC9zXAbb3RU1k1T
s8sryN6YgFVVNE37SaeBzoXbZCT90LHFBZENkAPuBH2IIOkLQxTGng3KyREeoRzn
gtp42/NQWNvrA29MGrgBMkVCgHdfV81BHdgylKnhAy60oZ41NtaiJf1RKSm+tq7o
eG/e1fVbv5BLtQOSDaCuwXGAa+iFPJZpWKBbbGBa76qiN0pRntxW/eN3JqAuuhJv
bf/KWJHvyaFhzQWYoehR0EvUN47xZtYbptxF9yGdbFIcgYjfI5l8n9ZUxejZVQLD
+Vpp6UKYT7oFzJoI13MtO6qcXXlLouRuwGItWp9cvfx6Sg1ojCF2lmOJFuxiarUJ
n/RmjoFQ6CAJwk3suMJ1OgnBC+gdIRgeOdI0dANZPUM1GSDZB7i2Lct0MjtGXmBV
7sF9EIEMSOh721pMDhlZzIEtU7pfE+gR2khTrYb8Q0yGwtC+0hdgLcWuueqceE1j
MTLgZ9VlJeCOWDNuM8fjbrVSFMKpHcj5YrBKJXDU2BkIlj+0RmfxyL2NU72GmOwD
3mB/oJ2mInvpPG+x21OwfSf8WXkZ8EAUSlsDznKPZ2BV0QGvGuaoJmHx2a66r07+
ucBLNoMrih34jSy50NQ95rcRry/hRfypPFWw6nexd4C6VoegxQiVeWuUCKGI+rLo
mmpp1V9PBDn7azWyblSYoCEXKTDu28RA02WKwYEBU9t6GVplzV2l5CArcDqIMz0v
u56WmbEPRf4ndHqjTDnVZpM/nxszpWyx6oRwxQY+vUZgDrHwtS1ALs7khGZP3+Sd
A5uLkHwRu9n6Lem7tBRH04fy1fVyiUK0id1WmxZ3SVJA/JsR5NgySOT4IJ986Wdz
xtyNDjkMTZm512CGRBL5SLJQI8UAJbJnw4+JXo4GDlMl0lw6dTjNtPY1Q4VxSSFd
F8ui8hZtitd5mDgWtAmJPoC6okF1B+cNWXUOZr3dt/iwid3QWlWILstjbxS8uuO4
8Q/z4zWN956VVRfx3QsKprskdaIvikHJa+k8JDFOzTt4G/aryEyig+nEZqnZ6eqO
va95qpjqhp/i5xXTUjbxbTLoyenvRF86Nwf1XqUu8P+mFJihufSswHE6IL4RpPA/
5eaZ5Ek/rgOnReQQhnKGRJljDjFxcjc+17Cfw7jGlQrzDt+EEGLKEkkoJsmSaqqi
Ibhk4c5KkD5mP3vBi7Dh5z6a9sIndLSHw+dJVk8KZJ/zT1dszLyULSfZQiRvkjOT
q1VVY2aSanc8d4W9pvBqFfY1nudqStb4pLstbE0cV4rG7RimwYQ1GRkf80hRysq6
6Yh4Hqo1DOU2IltpuyET3HaOai9Oai1FVQHzabdYUz8B8vLrY0UIxw/FNGkObC8C
3W2s3IhNkNxCbqOXbEGldyrfApeTAFU+Ccyyl9HKb3/EZhEJ5OZLxfpoRQYugpNJ
UckJipqCddoL835zopW6viFGwTTuSKkUPW8EMn0aMZIaQiaf13eyOYKCKyvBUzB/
WSpNFX+pLKMzxwwtRHeFEPNLifT0e/76d6mubTYtz69GEqKdq0A+RybVaQXkkv1+
Ube+etq0PEnD0fhvmOVuCQye2RHRglaGrcqmxpZLF7rnK+ni3H89DBzSYoNsnbP4
A+5P/KSWkFECpvg3vY3LEnrOWoHkdtgRSNxb1ZvAYlXDU2lMe4JJU6shY/2bxmUV
uoZ/Noxm0nU3/CErUesG0/CzeY8wmPMSK4r5s3wBvMOJGlfHKr742Od+ujkzHG9l
+eOaZCJPMWVscvO0DOXuYE0fR2DTqZiqKbB622PG70Tha+AQSnXRIXRUQljfvzMe
2c1fMsq2mM1vUd+mIjGxJW0HGCqGYkPi9m0cCzrH3TB1RA3X4PLT+avA9zMDA7r0
S/i0pF4BFE16NZD+OIN74pNPzEePvW9SUByBy5u692xo8ZXV+b8b3rRF33ravxpS
lOFSKi0dibtiJAL3EQ3/jAitHOoM5i+78DWXAcodoxhk+mNObOMlJlOFdpFPU6Jv
GASQ7PGWuGwx4LxoleMEoJwARDOCpkHtOTnLkibQzWhlMBHGdHTU8JFfg6w53hxw
v8xzzv3Hqt+HFB+j9X67qIT3whfzC9uzkEA6YOt0EGZxRpwQX9DcywshwzbnipDa
jkjc/HrpT4pT89C3k6VJxpywEm60x4RDHqDyFJ/n5iWdOfkU4cUEPF6x3PP0dQgj
l6NpMN2MtXTPRpB5wj/PF2IbI87BkMA2tE7J2g9oIMXJRvk7XV6AhSa2FIX++KZw
yJ1ltHxOZu3+Jol0YjYFkdVRbus+6w936BQATWLZm3zT3tyI7bSLydNbdVMV9UJ1
FahsPfFKHrbh12bi1PYK5azk6kMaNK6HF32pZaR/PZNJQoB1WhFhYzZYedZ3clkM
2EnVff6W4zCh/Nb7+RxVTUVXgbWOM4B3iplZvWQdiDkplxLRtP6O0lD7bl9e4ffD
WXcCzUjNEGhVvwt02gcRwwBm/lSUKaYhelPiodSu2R7LoAlgM7t1uZywWgzTetjQ
W5wZP+kI4VrS+TxhKuRPpQ69tMqNfCBoeScdwKy2ctJ/ID8nK+9026dkHgZvKqx5
iIXNqmrafRDd1KaSxl1Jtg5Z/to07/cff6GIk+TTpiZtIoy8YTMS0TNw3q/NqR41
XoO/SjPuQygIjfg1LH8YoElWSSRcz/3mI1YBZ5izPJPsvI57lheM7o0uuQ/7CMOd
DLb6DYD8zXg7nNorrLNfRFJWm+GS1VVdCxtoOeMzJqBhIrXtBBcbrp8QOsyknd8i
qItULHCPim1VBM2x7x1H99TSkpeANSBiIoNfvehXnbNf6MaXP+JMMyVf7HgTNwA8
8WV2eh1OTfvndEGAIVEAW8g9h9wBa3uir6npDoTc0XCKaXJorfIUXENi1QYdjU/H
WiMELU4iMoE8cVMnkWkKtch4dLhgOuV5DbkeGRcFYP/DkkEf/t6kzVhNgG3WR5++
8EIH4q1/xaTV4iMUNiqBfjdlvfnkiQMrRdEX8WIH5f0wLiSuRG5f/ayd5JhwH6+G
sqB1E/+sfzjeFGNKzMEaBLxgT6d9XCTo7kXX+LJ+JeVAQYdI/YqcqwKnJsYUhuO2
edGFuTBf6Fj5KKQbYas3TigjCnZi2Z4xeFfiO+sMJT6Jc+T8u7y1JnmGnHEEX6D1
3eYH9hcvfNKGGOK40akIuC9GaZMOtEZ+cWUxmdULzwunHlWDVkXpxzZrUrXq5CMI
ov4WJxKlZoAEL1ElV74cB82ZHyhu1znzRN4fStop0pY1P0O+DwjKAl6zucpuxx//
vpC6D9ArM/SUVJP80NzNngIH3XwnKx2Dyi5a+ZagJTlpt04s11eOVeZjB6HoyQrd
NxWEynj9JBnYAIo+ypIv+ydsWrCodQAyJcJSxkJ2hwWCQNUnREORT8mCFFsIRkVZ
zgv6uPb92GS84FdQVcxV6Qselqf18zAtPHsyrCZPKDcBj9l/Y2H5hLTplUcYS38h
zxAuU2UrzGrZYkEldysMORcYJIZMpvDIG0G4xboBP/NFjuSRMatZ+lkTYW08piw6
IDo769zAKUf/aJ2bIXUqQqrzvSKoSImh2+e4NDkzidgZ1AwP1nWum25VaMhhX0S5
Qk1ChG++WP3sdbRwck/IL0MY/MAudsTWnX6hMfL/XlhQV02yKPkRGfn8sHmqa2Ti
Uwkyz5PtEqckwoIKCmNlBf5LRpacbSsGdQgN0rlLebQIlj+viZ0L5eRRhTk04EJA
2cAF3+3RD0mQHLrG63XVNgMC4D6mJ2Q2CfsD/uWdSRc3gyo64xyubyF5VJv0VU6o
hVpZScz+50ghsgrO23OvfCb/5HsvTjwRYU0m5Ks3qIHNdASFSsy6PIP1UjmlPN0e
IgxJF45ha9P+kepq+1b7WpWP4fXt+6JuinWyXhRBsve7+WAioE6UaOgKBn5OlkRA
zAqDNe1inFl3HNIzIImDDRFOyLHE2HdCbyJjirhxxcK89LaSScnCXMEm6XlEP3Id
eSXKWshwTbdI6P3WDrouvWvtmQ3y1fXKU2cSy80cjC+DpNnL5kH/4ncqawRkWfoF
ygk5Waz3z8p4/o1shAi2wcIirBBPkHe7uXdEXiVW6Kf1ZNNi5gXZlXH0UpidWz3J
9NE0mSWYP/CT/4FoQHb0EAUujNw13QA1jxjKwQotwV7uZ/m9AH2EpliWHg5Qgmbz
YmR+wT8pVDQydtScblVZI+U/bt03TFkhbkryWF0TGWPsayDGsz93AG2btKZ+/CcG
jlrkMOCQ4H0D7sbE11RMCNoxMJ0hNa19NoBfZ7UQu+AI/02ipU/AJAELFA6mOVhl
QBXugFJVgJ4kVXp4fELOmi2jNm75PEu1EcxBdv88U5IlmcZ1qXHJHt1o1zO1h0JX
QB7e3o7Xc7cRDLJ1k6/HB4rUh4gElq20Nis8tV2ZJtYwu9mWQUFDGX/IYtStTznv
T0jEkkIvfOYqBNK/n+4mM911ZwEojP6if9L7y84hTOmKHqLt/xYWjtJ4HjQsFau7
ygg78K6tdg9YtK72SlBZZh9yc35BpOFdxuEUb1k4xGDwVRfIvdbvCnKj0OQrsqRJ
I/IR5Pfsd4b36Psmwpy1lreonSiC2Go9vET1g6l8U4M655QsGNZXlUnRa0guPQO5
XZazvwE/yDo4mmV7/TJ+JqyVvawBXzJTQi/gjDgS9aNwbyfrb/cnfSn+pvIqfVRR
xksCAN44c1VjyGKDO/NcTdnKpUgOuv9Yun9TpwiAFYWGJ0uxVShqZBp6q5wwEhEP
dD1a18KqOHl3YE72Fnv+IfhMnQItKfSMQIz7GaOGaMlWlq1aH7OPjF9/F1enJ8iF
3ZiiAOdlwp4uQMVYxAeReL2UPV+M+0jLBJIhMrHi0BslICPudo8gq9B1oXxO6HRb
KGDK/9Ubk+P2AZWFfCmw3stNCz8tlCYBcn5yOictVtzJRhLDfuME1qxSh36qi30N
EWIRMkP5W5k7AzW1lj3s8eCi8W5u2OuT4tOdigaijfLgwRpBuiYS76pMPciSjk1S
izhBCAmoviv5T98p5ER7HfzDvhi/8aABn/QRZKGkDqzsu7m7ui0omXwhehB8BjQi
ijPMS1/HHO2BRALy1wCxxnRmD1EFh/x3rkk/j1IlrqaQd1Vg68ssOkvaibhenJIB
E44GhAmZpbPeGKkBzGHLT+isuSFL+1yIzEHTUeBchb6zxxb0hAoiSIHLR5SugMp5
wghl7Oon/VlPA+xELxgnF+bIWnbh1dDz8+1746Dma1FrTBGgjt6b29vY1hyYwr/Z
n5FU/fPuTyM5GUEHIaqnobmXtra9Yfr3cSyRPkhlslsgf+XcvIjWktX2xhfDEAR1
wzgvwAdCIWiuKD+COSQQ+2BqpgD0hGtKrhINJXD0KU9+QYws/KV8MlzIiON6+O3l
/sdRvMzGvPhl8/ZxsqtIUpQ7jEW9VkNoclvK3paIL6zPyj+/XBTZeqyK3S9kcTeD
yFV3J9GnGrjuo9r8SL3RxRnN26qgl10L7d61iKgD5e43gkaVdAR65DNt+miqyCEP
960dlFeziUZFYghg22Vc7ZHYfOl9UZq8YowAoV77stLjkF1q44VQYTPhIyuxQGEE
UwH9YzvwE3ytTSnWpFBwlw8VC0aISZvVk42Dej7VleO2A0LTN8v53VJSkFRX5aJz
huiOi3Jxy9LDBtbZRB3lVpoKlKqB3Fqk7QOXeavqqFZ3sYyWVj1tVKypwnnT/z85
mq1JxJ3FsSBukdCc77Ba3ZI4P9jInmwDR+XZ8lcpu4gk+IFUKseef5zFeKSYsJxt
OOH3EOEKR51Oz9Gi0a6WbvY0TQ4iPbx7Mg3hNRJkgvF/IWc2fisqSdv1i2rEY5ip
UcfbCdwzrg3YrlimwGXvZfeswXOEAb3IWN1KFyd+B8ZmWq/CFy7ouu1/872EQFaO
aXY9N24/nYXllaQ7TGsnhI81ebTQCrPz2SixU58FMOEcu15g9HbjCzlGXeJ2qlSY
NVK/EIz+AKdSV+QFwiXdoZIQz18xGnuGJjLnSRmPwMJWvVtV/CIZTAyorTn3m4MX
WGhnJj2iz4agZB+2+kjauAe5LVh8FxHf7CcInkTxsQ17Zo3jH7zCF+/uO5GzrBYo
oFJ2zXFExRRlUpFsvHalvMEdB4kVcgoYEWfDaqHOZALQaeIa71W9JU9XV6Dxvks+
t48cR+25s9ufo2Vnk+vV7LIbAJC1sDHayyUxoXVGkznIwUZYKHsV4ASKcuACUkOm
+bjrm8s4K0SBLCMiTt0DUP/NzY0XdkN4TZcKgx81ARiyMWFg6Jc1zX4eDjRGKy/9
oSDsoUxaa6xOnr+Xpao1tOUR6QRpZHt7NStfvF7DXknTbeiK4BQW7T2HxDcEFT0h
tSLegH2ZPJ1KNTpoO2OxYT8RFy7Xm5oXoR7VzCeQ/Nzt/LVSS3+JvTK6ro0117fs
htFM2gEFH5x387z19K5h4QIBhAAULAyGfEGgSzNAaCo3GXmX7EtGUIitPqiITWMM
OIKe13KFmZN08/r4zR9yF3tE21ssmiT7KujJSMNSYoE+gGu3YLvxUq5PntZn4Alo
fS1MaPzHfJRdwERuzonbOfoio0y5VJg3ecfgSLXh5Aw15V6u5PqkJBJIBq9Unleq
YQ7rog792yQBo1RqlDTvZKQswaj3dEtMxH8gKuXHw9YfGjYnGrRv0LJ/pNpHXJFk
Eoz7FCJ7pUJX9QoXMP7gwYWoxIGRHijuaG/l/zWHoJshMNmdiw3ha81hspe2NKgY
1z3xsajGXaMMMi+TrA2ROY3gIR67acDq6uBWlmXwS+/SAT/eVIefvYe4Hc+xYa0x
00eNhMgwED05al0WlDm7kcoXK0yCFfuFnY9ROenAUNMYvaAyMlEJLHDPxVmaDqQM
p5o6tjAljVnXTRymXHoABeS4Q2NGjmcvnRHfpVYRKgwJAJ0k2Gk8CIyMIP94L9O2
06fz16A8umjdU2QcWnZf/2mNxGfwSdNR56tDFXsZkhkLSEbV3oC1k61eziRiiAPi
NriD8Eu1Z7iaNQyQRlOHeSRq5VYJQMozUis1qyF2fsoK/xAIVOwb6VaVsBKYph3Q
cG2h95EubQ1xjI9qr1O7nB78jrdius+U7WoaNM6eu/yzcAsBJoiYp8a42+1TlhO9
3sDoRD0NxUhiQt39Iuxjd7/7CFK0IzO7gFeqNIW/6MmyaN5oqez8PirQYGepquQC
78uNZGl1dzdy9PBh2M9oV6sWynQLFBskiCqcsHGmaW6Qs8N0QpEqGuw0SFqPRo91
D2ICXbT9ud9VnwD12m7S0klaZZcfXaODiuBS+6lQGZVZGTZdHfQIHYWf7AkzitlS
7l+cxZWRlwkG1YR9TLAopGP7jWBwlOch2iOe82p7jffDh6NMwVQEeUDjMKFztlDd
2/UoywDLLP2XWqzACZ03W3rmNNP15+Ee0dmdLSyxHC1GNg/zAVvCvi1k6x2fT3im
VtfUOP2zCIddwMfU/55YLKwtN0UpEO0B0rDykzXE7FP5R7Hej3n0PosGgFupk9bq
ls37hKjR9ziUaacxb96TEArGLZf+DshwjQYcVLWkleN/ctNgd+vhj3QPTsyirmQV
wXNyaieedvRnEG0pK6N1Of90DLj9UBniC4E9/CxCwTO5NWdgxzon9ddbFWjdQOkD
4PMXmNwmIR2tF3sGOsLp1cvbMYC5IOZn73AY+cyA/mWBMRUQ1p+VDrLY9Tvu1jHC
GkM6pwE62cIYiMTa3qNeehjtmuyFCYWQ4wix3i8YsSlsZ65D59pMPAVaCNFGtAvI
PfiNOCRxgrFfk/ztpx/hgpfpe0CuZS9fD8zXrt5IJoMp5TNGJ0uj6vA0r+6IEd8t
HkVHj/x3/NyZQ0nwSLchJK3y4bA2uhuGIaFDKYDXrORlIDtYRHDzHMwTvyY11jRs
aE8ed4nUvoucfUco5T4PqXf9VzkqVEOjEJhiSDtPz9+RpZxFOmnorI9oQC/PeijP
EXubj1406IiGt4unvZob7URZSoxUTUWAMEACW8lpdE9RCcSIAsHvZS55L2TkCV3j
DNT1IvOeDgG1qsH0f4Gn1yjdRoxGmIkN+1Rf6umj86Mymq++r1RkBUlY9EjkaTOk
W9z7yLCtvsNGE4i7F74Qa+YhvOBxYyErgpdIrrJT5pZtFryfwZ46go3MRhOn/PSC
DHjgN+CXNkkuYZOljYoDDxU510fnyquYXJN9q7i5T1h51Fz5NuzJooo2PlPb7diK
Dnt6d8Mxde+PGIaSnHNUQJDNeniXtaWLsAt1BtNtGuu2kZL1ZECMWb65ODTlckdM
MFMfFCBSxRJTd/0ZzjCppA/Xh6A9uFfx95IqmXit0lznE5bMWwseF0YE8nKVqNgK
AVNd8Sf2no76RARyg6/Gnyvzycfb7Q6KZOR9RZQA1mrEcWJPq0jBG6YzYXxT70ck
qlMf3fRq0HxG9gew8P/h5uI2Xieg6WH8KytvUc/NDI6KvYtpOqKAqRU3XJrQwXZB
Pdd2/gZqQr/Mq4McUmyIbZ4UD9UZsknj8e/uN+dPF1wgV5MwaUmS42qezOeJq/M9
6UB5FQkgFifg0sap3sUE+W77BTQKoqktQqsSGhiMNaz40hb3hGMR8S2+vs2jX8Zj
F03v8NUW+i4VibfBJIcOFznvHM3AyDBwQ8V+GQymNDtpI6w8IMDD6EEGsqshvAPd
4x8Rfs3xQMQWiMdD/nmKks5M6hcKpLITOgIx6y/S/rRVziys0ZQWms6rwU/qvjk0
qEa5pbvzEqp5bE2kC1gMhj3eJe23D961efm19LDCYKBz6EE51LTNPwx1N1XVacA9
h/cH/QyTTzLA5iPMCFt4yol5xS+LZsOqrZavQbb0+EE72mQzz0SlSH4Gf1FYLtJa
17kyRxpIIcEJGQNzHKU8S4vAp4+W+k4lE559bCRLzRyhY0U2fZ71WYzsHvkYcpV+
gCbyba1lUnPjufWF5HMorvUHWKguO3k3Yo4CzmqQt806Rgs8ky/qiXDt8y7Yu/E3
GHmOP+x1R5+T9ha64rNznerFPca2UX3BREkXe5kf2ZjsUbri68WIwNzoxfplSdQX
hQUgoWOW5mHGUv8Uteh2oVWlyf9H4PzuD47c6VBKYN67bZkEJsozNvl6DPYFkslj
szhcWJ1squTN6NXOYg6JrB0kuuWjmQ1XFjR2PqzoYrOu97V7gb8j+daaLQh6PiY4
eJGgTUVGqrLSHZ0yr5E9j8EcVReQgkI0T/FYWElP46pT7bmZBY37mV2ZeDwO4Eex
AiG28MVhLanbrJMStD4pAam+AdE6LjgW//Z5Dwif1SDK1LF1+YwegwzRN7d3g5f8
w9k7oAZFFGOn82B0s+f1j0D5ySOQF6zpaAr/L5dT6O5VMfVL/ZQtCoS/lRqlIJGA
n12zDIsSTOwpbxzLBhIpVGmHxkZh0unM9cbve33nNCPwGwplxRszP4F92tAc+7U/
dxvPbSxzcX2yglFQSfPK+lFsVQp+iWkDBMnOHEH9fbUQT6Yvobz15err4068dHui
3KCQ9NYDCE5UTrqFf1g2yGQlFfXEejF7Xck3P1xobdZznzvThJLtlg1SXxzJdO2P
SjKkPP/i6BFrXopEo8a661wiGV2y7XTOFz7hUEF6xSOkxhqOY3arStxpP8itwg3l
XearAtsnK3Qncibn3KW+k/EzUALHzZHwPtIMho9wm1kjM77UlOb1bLcEDSW1zvrs
JUyLPEI+DNs9iZZrm0OGGWfGmvbQ7B0/tPjpC9z7rVvE0XToTEyOA/1GlkJ8llGb
kBd13Ty4wUthoh3shKaL3DFvS7YWQjRB/8tEK4L4OX4iYGm+vu429CC8QhEe4pSl
a/nG+Jm3Syskvpyy4r9qxqwBo0DBMS3H8AgJdH3VpW5q3Uzl9woPRRy4FiKmFU+p
YD67lPvgSwRoU7vDS6JZtANKk8FbVNfJZP5sORU3dU+2pfz7rzdafmyB+zY9G4LN
gEdbZNyCi6ZqWfDh+sOm1t9fxvqVvePUUQpLz71Navk55B0/dGvGuNOB2CBMVHgO
edDej+862tUIZZ7jeo91r/7wcLMi7YFlB85kofcd8CdnDnyY3/XNIz2Hng0Em0SF
zG1dMLZbSF3BzD96njeLwibdtZEo9fXNE3IEjjd7MbtZP8ayTjeEEOv7BFyeWnnU
7+/WumYKUnMQKwZOgalL3JVCzt7eY8EE34JrmrzwnaW8C+U7KixJIEv6uG10fM90
AwJf/jTMoet3SYHbF9nR1/V64+Vm2oAp9XbdZdDYcpskWzn/fKcrREw0G4YcVX+y
Wo2QD/eUGt2UEKaCrcpyMYTM20UfMrWZGPpA3Pb9p96rOG7lUdKttdFbOwqpgEH8
mGM+T5QpmxD0IUbeMxj+N624F2ETZ0ViHWC26arErG7Z+k7AmZJsFJGp1/SKEMQS
laOIdHeo3+4L41q2pGDFRnnqLgFE/ujArESxrbBabInIQiT4PTF1GFi3siX4FaZm
8uq8NKAUFHHGsaYfHDFyJ3Tf3Aq2pG0upPqx1/CITHob0/a1MfPPRKTs1mZFEzYk
b9KyNd6hXPztczP43UU6f59kOSVGvh1khCLgwP3CIPmY/MixuxPxvQohUomnHlbz
xlv/AZhjBy6te4ijyqEkDbbd0QDzk84HJ/9WjUWQDVqbY2uzvkUwN/5zoCzkc7Rc
3cBlP+HW8rNUlwd1BK00zOXDWAftfCr8DzZK5E2s5+HJPRKyZ1WOTO/6bAmAEMtM
Ewwrd2Bj0LeldOfnOIdQBFways39NF/xCjeCrlgcpno6j56QjtPUmqNdhPIF/Zpr
TVJjQfdXIn55Cr76E/EFcuo5o2ckdKcmBZ1kCOrlO06/2oIiv5kTWFMn0oPoq+bo
45cqD6HdlGV9E+2ugeS7iKyuDx5fw/OGpTaomGYtzWcp+wJ8pDFLyKHPpLEQ1tq2
7lrMuK/79iFEz+4BkgvSI5PgGdWgX/zGRED6YRMWqL0mPzXlRHXZpjvghJtrsFFA
Xfxkj/1KDfeBnGBENTJTvAvVdYgb8LEpVWLMBHebIrQdqHMSa1mXvUMf1+zHfntK
dMN4AsJmG/Fzu9T9XIChlDdh2fyPcuQioRNwaSlGjkT3apfmclTeCJqXp/YM+hat
JKwZlAevUGiS7CBDFhAzw0kgJRsmbznA+A6WHLetEAWobhWb3L+Nip4CIOQfSoQI
yiJBXAtGvPGr41Nxm/ODv5RsxF/c12/VthW1PqsADKy3WIZ3Y6qjPAepD65MOyfX
6VZZdfovDF0nJ1j3KucAlGVSrLABwnQg3umvbDZ5jsxFibAlDl5wXZ3ckQr9cc21
IZXZDwXZ5bNJQQZal2GK6TX7mSQEw7AmBGtcOqZwuFn+2e5s1wNlyBszYkxmNt2w
9qePypa5grcPS9OL3d/Wtf29hcJO2sK1KVkj06oqmf50Qy84q5j//ptT23N92eiT
Lxu/Ogr4sqPLhIN6eHx9CAaJ4PyeQ4sOrmkOhzXhMN3V92OOilvHmqQENlGf4J/j
t/DEgsfVJMs1Z9xPAbGI6fXzTh1GVXY+N0K8RNOk5WFd8t/Uprma7kw17Pg1akJ4
4407iLroWiMYZKVFjDwpj7/jbkKafx+nYgyJoN13oSqogIc2XoqrX5jLKOg9OdE8
tKnu0ZyIOGfp4I+zuM9oDiag7gJ5uKw6MYP68Yv3igF/UUgmo3qP3Ho9sWHZq/O8
s3tsh3m+NisqSx4Lt6pvWytDC1d7Ri/2nIhTBcqVYXoueYamlOq/vXO7KBGef9gz
H3yZFLag4n0Hg0jiyA3DF7BtqD4QdbapiVLc+wX7TVArYCVCJ4rFxx3ufIA3kq7L
MiyXIeL+nRfU+PsEtMM8xggMS2DawuBnDhWMWZ1hT4cdzcLVUm18eqr6q4snNMJq
g4xf8F2S4i6JdpQzOpgsqj914MjXfhQzrMj0BdUuUq74vvSRMvvk716rmF5phU4q
ZTfOd8VDrByvKJw1xxg4+lBLBgewmOgtK3T1U+6dEDb9bu8iQ3F1clwaKxLMja17
V8Wfbn4iRYzmI77CMF22L4GyhvQpEv4OgNztvQRrA84fsR252nlUs+oUSFJztjqM
me147oRqgh2IIScch4SDipWzPT9Pz4RFON5U0HtXd1kPIqV+Q1k4sf8wKjjKurSd
SrYltROiNxwhPD2XwTBaYtfAoDaVBWRFj8x75dFzkPXM9sjDk5la1zpkiaegRr64
vdy1GBa2lc7e8Hm8yMEy9xX79J3GI53ZNYohn/hn3Qx0ybTriF8rSE0j6RmrMxVl
8EK4K/iymo4NPFTqMakTNIe69VZVZS/6NEV6zf6MR2HteuBSisRbkZ5D2BTyHad/
2nZRyrWskWjPYRwNdbBCOFhwNVIDh2rYJ+RGrLgTba/cHttJ/xbKuN+g1jflk+sy
o/Muok1IiUI7C/GsZV4gMz759d9eNahn0RUgtYvF+xbyDRDSbAor5APTTrTR4UmE
O/uEr756oNF+Kpmex31RzX18ZjeOY2h6fTRsbCHNrkdYh78z2lusBKjLATumk852
w9JFyhdbQxbdxtP/tI4TTEPCrR47jhABxoNnwwSR7DS/xearBRf/U/Z1qsm90Ry6
bslMT1AZUqYSJtqhlVDXeQvSgC6Oruf4bQI0/ajFPm34DOi7AUXCjQtO4Ht5Y5BL
ZX3sqm7rM4T6QQ2fUi+XIVrBc2YJuHkR6JeefJql6zhGhZppHR9oveqnZVsm5Y5o
MLadVBOmUqcTx2IEytD/ZdYedzeeZyXL503D8XEWP3/dFZ7gCmQS0zQZ9dzIV8Cq
+wqGexS/EbWGtbTfB+/RD/ZiH+tL612SxVsciJtojj360tXJO82osOYAEBOasTE1
NO3IpQt+q5TARIvzbiqhTpZfcW/yNMHP57n6MjYWBVy+0QI1CfRgitEWgyPyVBeI
69fc8KRNlQiqACXOuUIB3Y3cscy0OzQjN7EO9kEDdteVlS4e9aefxpzMaTl2Sodm
40yK77fsE7eszNGz6eCDhHx2sLzKKZyRf7w9GgXEngbe+LuFjTQIk0IZfbuSE+kb
YwDZDouY3lRZpKHUfzMag4OXIPwirnfteNZJ9jIWdUL34KoNJMIkdVbeIzCIRC3E
7MPquvaPf6LrgKv2CBGVDz7BdNgusWZCLJHoiP+PyPHb07Fxh7kS9ELm4v+RAmMZ
FYV6SfVtxyI6yxgXXCIEu7rPkEIs2i6fu5+bUt0ffzfQoF84NVuZL5uCoejnvscN
D8GwbT7/9vHM54OLaXbZcZ+sWSe3asLzLkabWnOk5C98HA5dNTGuqzHuXO7w8CXG
UgbEtdIfgtJhvvYkFpAzNwZiVmyONk94qxDLkTlP5nEapF+6kLC+GgtUzApFfjHg
r/csoqbENxbHh1UxpOGhDEZmeNUJweZ2e9FEhQmytfj5G/dMDQPPE2xyha9ovEWN
eXogS5jO8FOfP4Vvsbh4iiW/yHPS34MsCAogqr8xZLJgJn/z+dKPtuCMpLD6fWaL
DwVpbze2Bybrk7ylA3eHbRba/Sg25Zt4lt0UwsSnwhFazkS0Y9DaO50Wx386HZy3
bDHR9WOgQJ5YYxpRa+MrdKNpYk8+uDVV1EFU61SH33zre8FJfNv2isx/Zo3KWn03
5dT3ThMoczNYepwnr/JHZR2LCrsjcEYVP/CyzNCqL7toHYs7Us9EG4gcX9DDMmvl
Na26heab8rp20hYwuILjc+suO69CyFQ/NSfO5CreYe/3J9xZMka7w0/NM4oTS7O+
vOCXhfNS9UteU1Eqt4c9RLPWPubeYesZkaTv0YHDIzRNYZbEv3JcxbsB/XMcqkUc
2+NdETubVez4LBmgjWg5J5l2r2dw9JNhPDrf0EGNXUkujE4y09v/ACbicqQJlJgV
k68QOvPiNLbz+MbMmoRG0GUwCPgnYUqOHKQAi3yvDuz6E/GQCCwxwYdwoTgMAoLS
MDvZ3quQIj24/WBgLXBe+RlPEUBI05UjqFi9aB1RR/nTfRBtLtgyEmtCvJhxuO+Q
2ELMSG2Vld4BsfI2Cp6VaOFDW/fx68Fj/48+i5LQ+Rf76PigISp3UI9M7fXieeWL
OywcxWCa6Pj909w4Gg24E67LoviA2X6AoAdOpcHAaVTmhHVyCHJ1d0j8rbc5FJ2E
F9F4tsEoapDHxYmwDAdeAvvwwTrh/rvQNknQKRgueYDrLfYY1l5iH/te+48mg1mf
1f/JGiQpFUEaGFlRl6uRWM/jr4JJwAasiy7HHNAA5GroT4p/eB6Q8SheLhUyoS9V
wLg4Lw4PAX7IyanzZ/VdCvhgNStRS5rvU9DaUgzeRM22fePPrgx9wVPEuaEl8HMk
ASLTjBuxvE0DSSYuu9sS0CDBUZhXuvH73NflzcJNCClRsQnWzH9/YIUwjds0iatO
G7x3timmV5D08/ChHNxsD8sZ9Rqs/rrBVjTwR0NPAAipNMNtc4R5wCCJA1reqWyT
4KPad174MZjBuUVYWDcSmJm5hH5tBUG6QaRZv9QeKNtZSHU2M6TcIPqkVZ4NI/rM
CXcEmIh2TP1TaBlg7CGmxdUTe4ynq9eESydzX18HD5m8PHXizGttqU7//sEFgnRA
1UEySH9VSQU7G1WnWNskTQb2rrjhUxSqa4vD9IKLgwdMouO4zm1UpW5CjMm0jHUn
BTCJoX8vCJolnMYv0Z6bkMh6jEcNPvSReV/JU21CEQH1+QGXJhzk9Y5MCv/MuDb1
cskEaDFejsuudGO3phOIFt8wkFK0rfqyYuySJhXShmky0kTqhniGda9zFKiKffls
aQdJSWG595k/a+bwS+pWDEq6rakUI/vi4Lix8rtAtPVzha9Y2RInRFUr1IGgsFUB
wr4M9FFfFu8PDXJRqn0tfdHjT6emk/GEYDq/JlNDcIOX8SxFC5K9+Rd032E7AnNP
VO8SV7HYP0AeBUabei/QY6eNsxLje33qYbuu55GVddVBbnRpC+uoK7c+XMm0Fhyo
KsOgRAZFuSL/FfFjnryuH45IOYR9kkKUDsfnaxLhKd09gk+eefRRjlTz8NeZjs2R
HOj4Df4vw9pl1vcePGPDvQyZTzJoHZq5VsL5QxwVaVmOs8c0ufNzI0lecvMf1smB
X8RBkPKrW8O2r50qT0ZdzQMfhaWwXDOn+Guxa8nmTw8V22vm8dkZSuoZi/TjokCJ
dAc0blAtY/PqEJna3F4e4hKO95JzpmUOrZ8EQDtmh3fBwStKVpydA7ToWwfrrcB4
n9t0mCeshupMWDli1wZtlUHZ5+rohRePdryBwoVbJUIckYH7dbN5WmU1c4wayQpP
UVKvszPhA3XF8KPdbLtPKSjaGnS319gvo4AmoFxEalShNcmlqyB8Y7c7BvUtz9X1
ApzgqBuzx1cP5Vvzc2CIm8FmvFnc93RI4wu8N3k0JJvlTd+tMnJ3x+L38PEqEo/d
nv4boFec8DmlycdPvTLcnVD18VYsxUUb4qz6cj9lVGFonliIJV7lWURxKBn8McQI
gsc+LoO3Ea5Fpu6fIOjUCWnLoZYrmdkE7z+7anxdH/6U7OktEid22sm4zgYNbYt0
CWLLpkbDw5RkwJdlrTQCzR9W5Ny4TEbaXmYJ5vFxwGXwetTb2p+pePBNDi9SgPHV
huGhSEAgkNhH3IQqLeLqGtqgGG5IVFli2Ba0JlvrlhVPIfKIhgdw3W/qoXG8xDLL
4pHds+z9v7dlrskZJYmfLi4Uky3y1upRfZ8IwfVudIznoqvTz8QJ1KwgUXNaS7hR
9KyfioHvAQtXoc+WJyIc5DmePJbGKV/nITf4yWgkTBUAB14YwhR/yTjAsGmxE6YE
kC0W3SdeACiISx8Mb39x9cPk3qW3kepHUeDBGt8PovjWU92DjqfJzORA6veo3w1X
5wQp9afq6EYf6wKbQo5p0VmksQMN+dni5imnup20RU04ADGrLyC8DV5muzxBHRkB
XtyYvLl/Q+TxU4i6at6QRpfbdD+iixRSe3Ip5wJPPcJ6MqbQ+7bl9953h3Cw8d9f
3a98fuvhjmDgK9ve+IhF+LVtY2NA0EhulkrYTg2AsQ3eH0DWgAgpv3ngBwksKGQ2
654N0dZq9zTuGsUOsZ39MATVR/ZgHPenXYb9mYWngmWXaaROwrVLv5UljA4kzDzr
ygaOGTFtWoc2I42FLlFdS+FzKbnylpQNNbV2cS2VkrSJg2lBCxYmV/bNYXAroen2
yioE2HGhOO7fALyqy7kGm9eFHXhNb8AgMfHAmaCcIX222+mwZU3qHDEwkpo8COL6
a7MfsVfSEz4E7J8yUz/6sp9So1C5BOMGdPzjxBMFY7ZC8hGXSsS4ycg0QxQ+BRHd
tyw+qs+LR0K8wNGOuzjpMKMVY3kYRg5xSBLvZ6p6vSq3rnk4H40yMxUUnQaYT7h/
Skgew/VHR7llXOFeufsws2AzyERIjFDQVlxuLlA+3a5XAw9Q6qsdQFLTkQPBECY5
2aXnTvsTgnxN0RVabDQANW205IlgfpB6+GYTPk1R0+ZPNr7EQ5bvlfTlbP3dra9y
RLQH98ca9HrQWFsTRAcysQr/cWdcDos30H73NERocR6rYvlrKmTU2vt2hwDRlyxd
dfy7rGVPkvhjiuajS7vOqbF9XLcneAOcvrSwMSON7i1+J5/jNIoKPUbYF614xQQe
KK+H1aqfIWUCG8Pbx/TMqGSwMKRyKyjFpGsQgHjhtzDwhRSL2hJIQPhLv3Q2sRv4
gKl/AzB6oxShxo8CEjWF2P4OHelmRZTWPaiJvUkkFmc704LsLn/IhcE9XOKoUDG7
ou7aFLzfcLdQQjVL+l6Zqx0SqERieRJjbT5Ci+uRS0IcakJFvrbx8LiZ2d782evF
7dmqthTHqsEY1r4HlU6QTcko6bk+Ke5KHSnexV3qbNuwDSEFbKiEgZQ95TZo45um
S923p20Pw98QfYCJFRovrEF7MBwYnGh1A70konI/Mo/bkUO3YSrforSKSOG1pRw6
SHGXA+F7VkWOFYfWVt+8CZ61FYhEQtpJVLPuDo7yD1JgcSxZm+ZCulUdkYirt8AS
IptcdCB6zZyTI6xxkA7YwtunmbnlFLZ5+755mIjkh2NwKpz9mu5DaERsQCSNcHxa
EjEd+z/+dF5CgQ1msPTn9X8gnBCfO8fDjshkRzl494RfF3uYTUPHV7c+fwlbOhMu
pIBpf77VLa8zWGpEFXp7j56+6MfHOvd21rzzgLwmGVfK1lCgyfBm/ijA1YRPmC5k
vgC0YIpMUcsstH/JHPL6jm1U8QS1hKwV3JG6kF7xlxXkUhjj+PsiuLlgmtJYbsfT
m12HpuuiiMYqvZbgV/wvXgnQw6QLi+0pCybjUwCJJOStnaKmCj6tJiVEPGhvdEgf
fKHKXlxesefQW3kJLKTvh7hYF3kj2I0ruB8vg7oXVXFF/KVwsomNoeoMjHQHileG
LqoUHi6D+q8dzY1ZSh+dO6EKHA0YP21Wmslx19Qe7GYfUrVF+0zXtVpjcDJnZPlB
Bu9BuGfBhfi0Gl9l+cIpXLhdA+4zM2UYHn4XqPr/9dPXEjsh/rJ3nlIVJ6uxNi1P
i94DAWDsasVZdkz9xtNNmoLyqE93hcX6I+p1bC906KmdAF/wCkLkoTdKkDY0Y3Cb
aBs5OIiW7tx+iP5AGC2Ao2OCXg/SAdSneEaRewN+D6YAHHd2GGq5zK0CrRnmlNQs
Ax75i42neXsU25omNZbNSL/fpVtUYxAJa/5UHA2/6DY2gw1s4qTIIBTZiwx53qo+
1dMcy1gB37hYSqNkiucqs062o7L/u9B0RHnrkVCrjULJk6q/9+gdF+TEYcEqP5sm
Wi5tH/3Yf+sYYxJj4QEHFgCLY9OWodZQium5iCra8LoxOuTyNf+z+F7lYQs4q+QU
djNq0Gdsyqx/rJAh59H8AWkRvUmIrTAE0T0X8suiToJtJu2ZmWq1Q1CuOIPtZ2iD
EHiv5rUkYVQq1OGZQbdXtwUtMr+BJKa1wzy5oYodUVQlPGfepLY3DBYWd6eukcjZ
/+3g9EdOPWx3e3DjhiGnZERFWr4S247lqO6puKdhMkAWP0wqs3ikjWHOEDpehe0/
uTSchkwqCa9lCQx8WZMXPOHPIUU+nNY4tfslGquT5a8onhmUV+hGSYHk5dzN8Rm3
+bYY/bfO0rcSR++IPcEha3FAOTBE58paFCGqDPoj6qVjP+KzjTLkQLpJkkd6lV4L
EUhYpMIeG7aCVGEtkdXQ+VAfEvI30s833fdfuuKIPGLeYsPueFDSmqXAOxT6L1C6
jgyZHmS8UMEdkJTmn7i9zkqpImF7l5uI1DUBcIm+nUrvTh5hVtFHEuUfe2XS6zLY
cGxNI8NW+dpgUGxo8LhZlApLC0J9fkcDdWceqlatAoMtI8hRQH+JUoFaigXKGpGa
Aid2+5l7uQrK1s7ol47c06Gb+Ohpbt+RmGYvNlB39V8ENxQiIDr2dwNHEKSQ0yGn
AfO5YJU2EoAYuc4gCB6vRKTlXV3/VLHfgpr+M9dYiov3Ppcju69ofGiY1R8sJ6y4
uUG+oMnY1jKixDFInhuiQo5lfDlcAHgAW1VzQouTbwgc1nD3ZIM8onqoP523CKvu
mM24JPIoAV0NwSYYk+yV0SbMvXkeDcJMBi42/a5JKkSjrX8MEDU70hnF8d/KoUq3
V8BPibEiFPbrZdgk8+Zfkl0Zw+JSw8haHKgvz5hmpW4Lg/m3k53slLq470qZ8lRE
0phHM1zB9wDHU9iNC4kOadghU+ke2bOq3sWIMANvPbU6l7zF++zzR0iXmyKRMqGN
OHqa8GqJmlnB8qO6K2vDzhKXz9YBqhA30ZVMX4a8fGQhzU4cnrJeHkr4CN4ZiYty
aH+Wbp2oFJnQW1U8FTQQKi8vDUC3FVvtFPHy8KzBgJ6GSzJhm0nsSFy5nF7dIHca
WpPPcZ60uU7hoGrmqCOa6tEbPe+VtbPUhK0KsqNIarqcgLbewzDh/Q2Uk7ayDn5i
uuZnj33uAGoe29m0s06OJopAa7BzMpRHO3+Lj6Fg0+gfC7aSK8RHzY9bNztqhkal
RpIhcr0AIWm4SNiLWHh1m+ygdPAWPEteLXZD/8leTMVKB9OOkSuSg5/jIv/kzNuO
pRO2SyQFqxOmAxRoUR3Nyv2b2kXeoGWDRvVGiSZU0jJ/rnnZZEdpzuoqZe5E/ukK
Oqr3462J1CmKVJmxo20OaTfeXmkeSiIxBVAeGTgm0rwxtqg0Q8OReWTWGSD21f+0
mhPmJg+L6FPHRo4fOGfwszqi/s5kRz0fWnC+drLmy5Zj7o6vxdmCKPmfaYbDXj1l
Ki96O/lF+mO5eBDmPosKEWtL3ym6M7PX1VyeqAb1VqB3xyPX4nlCLl89704/tF1V
S0lxMWKMfsMXlF/ee37DbRUrNDBAKO8mHoGJsOVVc8YlRte/czJ0KzmODPMCMMcO
Rv/oF877PLSK5rEtXBR1gqVvE/c97QBzJJyVYgBc8vfC1J/MVEOkkV4q8E5DaLlp
ZPUeqe/wJ5AR3FfKA1iWZcX1eL5pPEiBF83THHwIp+VkaWQabP6Dr9kc3nmPBbwt
WS5xd544uQFUaZ/nWjveXHCI5Dy9P3aQwB7fZCG/5fB+aySypoe3Vdhqk79dvNKg
SBOR3fIrns1Fnkb7vz3IC7/HEXwdNIMWgpqS2j5Vuv7TNWc+CIJYh8NmiYOb3rbc
BbKn0UV2zsoxqNseh7G3vlKQOPE2d6+m2WszXz3nzqFqJ8cAwtEvV0Xc2OZgCiC8
4/Fuv+JlWZMOL1HFP3cleMe8lUlipH0mkVnDWD/y4xkEv047/uqPszg56Phk8+QP
b27ROxJz5R1VI/j0L0+OjEJT2AtGU8x7fRGBO+T7HglJf2H4ZZ3u4dFV1nmKk2hx
BKalujo0yaFOM5MZ/SuP52TMVsQP8/6lN5iNYG3t2StNI0CrrayXOBQegn30p7KG
JwLaFHlrivQ5udt5yANWG27bOIr3CxtyJDU91lvTq9XHDKIO59J1u/r8+X6In5I2
FLpFNOzDxErMRiN7Fm0skIFKUxO2QwL/asdIWmn7nq5TTNCM8fB8gkQojkpGDuLq
AuWYRkiZ9n5zZj2grtMqFlinUyEwRov7NdLWr1MHGt8jGialh7EodkzsyfAvB4dH
LYZCbcBF0Olf78CeRbweCQuHsHVC9LmE1xfqaF7+2++PlIfCZVhv3Oo6PJKDr3Eg
ywlTUqM26tYfLRJT31qJmZhWlPruBlX0hmFHbNT9bXo2dpL1ieDMmRTbDI5UiJfm
cpfIzVR7trRM0IhCuK4CkbeT5rjeo431XVWICgnxd6u8q6IIyJ3xurBKiS1mBAbJ
CuR0G1ovBz8+JeBL5/P9/JIePTJgGbpuejeWYmqefGhtjbwZ0yY83RW3Q0PBJmU8
HO8kHzuZGfXaCKCbcon3haSk5YA4WAFZQ71agD3aWF68M6Kyaey9yDko/4dB1XBk
WM5P7z57LiILu3XxobyFJ/nNYH67lLSuipElg0Rs8vcUwACc3bbg1F7YslLnlkvk
ozPanLNYTBpk/93bg6oujwerLhEsSs4TH0+wikYYDLufWf1J+0PqKJYwRYRwGXcQ
oRGxx73oLn/YMsAmj7uItTcC9I/T9/IQoja6S8rujp9u3qzHYTu7gOTmoDLAPS/a
s866aDDoCthY9Ifxql6SCPZ7p7QRsFWmYqdyvCtA93cdwYi3PGdkQVM5p9VqqeRl
BT/U11+34l3jGPnQ1+DCSjIiKMgRYYiKF4Jjm1Gq3V32c+vhHVBRQynow2ywYbkq
coNsS1wdVfg3hce4g192hLMlBN2Ib47FKGbTtg3KyHxfHZ2r/jcWFAiibQYYcjwH
uhB/dS8LLJt02kQToSzj0vVDz6+uGnwEKe31Ao2Pnx2Dmg7kB4zcxYkpjtnieu4a
GzCCeqUkTxLNIq8We3j7k+jkIMPDwJdrAisq0ZFWwO8ys+iPFXIZdDJRuyIXlO+D
ePKmrBanbLlEvOuZt9ZwjB57pHtYqvTO6dmakFvmc7G9aGgtM0H2+LMmXv/Z9eDH
qme2otoEK7ykCTosKJg7Xcb2N87R0gtt9kldCD959hgCp/9+t1/9Niw1lX0iD84J
OTTsbTGkLOwWmSOmgIaOVzAlCofg6tNLzwvyIthzbwuvOZcnTgnljPuNeEqt25hm
Ve7trOtR4UHtoO5GgqPy/dUEm8ApBXJXrpnZCTiB754hd1X68xyvvlkfTSHZ7PPT
oElGE21zvdsDTWGe0xcOIdnJZV4dH8Km38L2Jo4M1jPUYHmRpLI0WCqL0rqaj/cO
exDNW+sXMxzKB1gkYOK3pbFG9Hv7602FNi6NamBcnpb6U+wh8pylpumymh5O98su
fyLDGgcr5br5B+GUzmR6HXDvzjNMJ/3fzUptOt3jpcNc9kb0zrWzZJ/inNBAQDIu
leeNGmQlseA28gPoAFYNeM6YCtYy04GkO+H3eT76fW8+JiCtLUvrd0gAfCDRlCBn
+ZutXXDY43hJjqbXn/jlxkZwMW8j1538Q3d2wWdmHtIsIkHLbIu+So1eJc+87Icz
kGh7f5n57JT4x8SeYVCWV1GSaeucg5JdVgrliEr8x/w7p2HASYDLTIv2tcKQpZmp
5f/aPSBauMW8NsYQv4Sw9aymqhmiQFuujHf98nB5CzKArPIDsdfwMkbGYaaK1yEF
qF1Upx6WuC/LwNZeZm4dugshPTa7SOH58xi9sKzzoVUa6hkFlgPv4WCPRG73dmIi
eNFSKOm3VjEvbrEwdDxBZwfF8aAH/Ho+zEYHIpp91mbCFrQ+NA+03QCQyOl55VZV
1Hu7r2f+Oh1Tn/Qbjep1i2NovzqIz0ZayJ6vU7Dn+c2/LlZIi8CbbCIYXdzJEat/
Sd+7BReO261edCdiyVAaplBStVurJ+kfOQJIdIQEQKVBEBvp8lHkPHNECsA2d4Qb
rph+6jPRbmv6uMltd9GreWrJd89NKm6RSzHEQsAJKwodD7ATIm03nHGPfx0w3V5d
hyUtwMeTmv+sdJt6DOTRlLuZ5t7X+pXSVSeU7sy955FXVDKOtwV12c3gYO9ZPE2F
Tbj45bBzx93cW7pPKx5y1G7eP+43cvzhtH2b9KliEgZdeUG0GEqo3XH3YGffRUMo
hGDpZBOiq9SxJ+cvYeMLU97WZ9CDOlZqggJVNfkCjDNUlpFS6jeM7kiZPd6+aI/v
YCSHhNnkdnmwAyZwRaWF74A0gAHqyGgW5Cy6I+gByziqqr4RhCwa5G59hVysQ2y6
p15iYwdWR7EsDjGpNzijHf1ymSNC409XfFnDS8YCDGVVuSRjzmtbTBik2UOHTgy3
2//4eIuyO4dAjNFiW4C9KoupwSLZyFImVOJ4DXE1kKLvJF3MqbRn/Dk2EPmW+ORU
bEEjmhMi0wppEupV3bTDsfH/D13ljTGnslYjctEQa463R0etkSDp9uTap46b+MQB
GlEJxZFVXphIy49bmRWicDoitU703JYOGU/McdALCy1VyOf1TymPRJi7qwICRIgN
eyV+xavnToXnhttwauXr8aQ5txV9xpnKYvtfckVg9PnOQWXJGP2W6ZZDKmIqAM0K
xG7iTzrGsyTkScrAnNjIPZm+BkWEOcKR2GcSnxilGitSPbnQROVv9LYltEyvBdMU
ZA0bvP/3fFzBZODxL+9xzoxGtpaTSCpKQHUPHMh969jkCHWGLpuMtMlCd48vtViw
j2Fmv541Q4ERT2jcxkdXRUs+THoE/KPZZS/VZD/lSy/fmk5X8ZSc/H5IIZ75cIlD
mR+Q07GIfJOsj5f+8AZI37+GqAniVOC0BIJXL5HbWGIR1n5rN5/4+EcQF0KmBvBF
VreQGrp7JjvHXZxUb7pPIwXSm+b/IFbX9eCUvNx90KknrlifdisaqJRy+EvzRnms
MiUtaQ3R9nNW+iFfIHLjTqxZN5LDF2yvvjtOv3/POxvr6MWjjlDbY+TLCzl+vSr+
ror/iFmCZXION9KEM/3Ph5PZnz+prAP/CIYQ7fg/qcJRSpqCZWB8w/gDWuFqCCKY
sH/hfPZNYqAUEfPxsA5F7tM8BXTWLIM8pQffgUW/9uMAq/x/z5LzxMqQ5HeFjdgg
RaKt1c+6y79O2NNR3zFT3lN1wNeRNuDBSU51s94IeYXRZy/VNnbX2yvVhYgE6aYi
+QyaKtFCSWDpAjEeFBxERph+K2afvrfIk2oDuhi70sCBoS5huRG+kwxNe/GwcN7J
FF9Vfgy+lJjkX0aWmC6PSKSMwvNvHJZV6+YXoaef1oOGrGKYHBzGjadk6OYaUY1j
8RPApsdXpny5X9W55k2X9yRikShkmLONlVNw1DM6wrFJowTBB84HWPyT6Deuy/XB
g2RwPiaKjOEDiZi/FV8petH6vXs5JKAOE64pEurdEvNoQXA7BrAzezeOlW13IG1x
sdiBS3rtH8xuDGHqaHdDQ8xW5rf7bc/Xk9rvJqNxWuN6aVBTIi0+aAI94G/WJwW3
gjfZaANPWRJq9myFAoeMzgCgLnubWjYmvKojk6plLDtR5TILyJTbBAucw6gbHpDp
FijgGLMbF/zD06Xn+3mZaA3moKvhzyD9O2GEv6GHVQ6igjGLPHl3tXwfLKyKZBZb
i897UaqcrvKsqDxs2CpqSHBu+T5Nj0VRdjAU05sFyb0RTy6SUAI1CDCBr4KonD97
yEaSvRTedsKHDDqRDSlH6E3H7YZHmUwebZiZtZ8G7pWqvOU3wZx2HuCVUb54ar3W
gzzzs6sxhGuvxduhGcjwnnctZ1fOjDljpPYzRQjJ98eG9Eavy21W95orZ7FS4mn4
2w8wg6tAO5yIXepjqfEiRc9FtYiH4pOHkUwBhTcop35ovVjCASUnaUvYlqzSB+cq
J6cnLE7alJl24KDuoyoMD6WtF2F7LYUZJSuxEAgq9/jpRot/MZQ0hEnrOqYcKZlU
gZYXaThX6Mx6Ibv1coTBhjETCFVgBTgEnILxaZwdCxpsKS87pTQz5vn9hV+vpr5O
3nQuIjilF1tnv6m7ynUpbqrpgI8HOHmd8O3G5wCN3PcgnsH3OxjfOqD2UlL1Nqk+
jgSAzEGRM8qOkIvLsPlb/CNeusvs8BG3URVsCftSDQ4TgoZxfp/g+E9bXsnT2HpV
Y55wN4B3E4WcV916R4ZoeHOpXM+VczIS21l8yQkiHNppPNCcPGvQONpfSZci97jk
dsSSotyUeeCdr5XwXkhzGDQoHsYBoH28I+iX4nrbU6hJCnHWF9k8WMxbZfYmF2PM
RYz4WAmI44MoBkoUo+MmH+Bg0FD+eruFdbnMsDDhLqYvrl/PZy3lc3MN4QE6PXcs
PoJgqXlWWbR9zXjJB3xV/Z6ZbPiz28gd+Bce/LMbDTBqdY2C9/Zptifk+sro/2Uh
0QIX1R6DkD5ZbhalBufusP6EYH1mOjtkXQbWeptRNcIT1uL64Vd77il3tQXZ1sZ0
LBQlk6SPm13yaX2hsd3eJDOoMhyPkpkzUx02bBuqWMGKI3WzgTxWFPBf2gzBd54D
o8NRV2IBF+EgfBcr1PAI4oTpzEjt2jAeA0HlOJfTegy22OlzXn8HQOxUp/7+jMGD
BL1KwqxM+sxoVh3Up6oenzcXvMrLjerbHKXSNYs9jXCEMtQIm0JvlvRQ/ng0mCsE
rxF20k4vA9keZh5ZV/Ur5XcQnwM5BRdLOQ3SM2/o6boWqKu95mqBheDQJMg+ku0d
8RGftM1LISvdV1hFiAOgxAczMjjWcqqi3iioVmOZfYDhWywS0sOILwCD8uaGKHrS
e6Sh8YCUaP2T72AIdUdrEdpr0VwkKRq/RBt6xKvx4woWl6fe7NUphjWJs52lrEnv
f8Tyk1a17Zdt/fU3ZNb88jrXYyU0UX8nVejwCXY503SIUx/p1lcyfUGIGAQbF8Ec
yaduoY6xHPHxtrdFQI5EUhJpxfF/PL5Bxc1g689AwI9oKjfNFsOO2aV/k8EhALZ3
TrzgQ5q6/o3T6mCRtV34rwoXyYKOWlRtjJCe8lEgpWKkj87mGCoPskDHLcOOqQNB
ZKSd2Rnd42pePaZbN10w5i6rVijQU1ANHw7CO9Nf07fCDVD6rMsYX04rnIZmkFIi
EsMUEUvmBhJ7+UXveyYyTml/OI1xvSBDlf3BtbFR66BzIKrpnNaT/W6EmxPTDm8H
6HoUBiwjKSiaQ5iHNVXhrHmGp8uLbUCqm99jkeM+uUlA5kiLqLAAulA0LFIN0Yro
L584UBjkHqrNiyhoiyisKs0AYlvs+JJHF4YUaeSiVyhTyLvdEoGJDeSEDcNehJa9
9SnmycQr+7A+Ny8WF+Fo12WyG938XsBIjNvOONXUBxGW61vK+Ih20qijLi1J/xCt
0rE1UzWHySU9mLdZUIskxbxGaZZTAIg7szSQhlZEVMbnRUsXb7outWzLnc1UyZXV
Kuv5OSe8PaghzU9gesB2amfFbMx5wTiu5AgpoBnYGF3yEutzRPXa/oqK40udXbLv
EAPhxOpsA6It6HA8UfZuSGkRDEiS+sbWHrnGYhjsjpfwIQPMUVQbCLb+tDxby9Pa
6/3H8M1Ei8p6QsX0pJN/sq3SsD3PHY4W9QDI6IuX0AZ+Qd2DeRnfX/eRReAH3oj3
txyEsmOxcUrRo129lxnNqRr4KsGP96/36J1NOCSXRvzQ7NxZzwNfudrQcjx1HWfR
NxkR11Ss8B24dIzll3+CW0HBPyFyH3G6hxln8hhF1CYAIjHEGolnMoVIHRP2CqRs
1NUxMRjONYRVwabJRVqtm27TpXkkxWZ5GHjqFOrm8P6RRuT+dR8gHV6d6jOkJBJt
X5Ad3fg5OR6QZN7jk3aiLGhwjdhks50n2SnbIXixHmiA0U/aNUZzqnSqtEgUReJQ
OnqiTJyK2uZz7I7Phtt67c2OuFqo1mbawFlsI2nTMPWbT3XPgS0dhpvMe3lfboHK
Tmd6BYVzNC+nik9povHyTBErA9vXG7vvrPdfRFLcn5j0EZfp+JvVNsXmqK6+1GLZ
XBdFZeIt+A4ktffifTmDzclTdKgkf5q2VM2sQgrIKznC/1ua80JTpbu3S+RgJx0q
dinDRpokrqczUELBfqHcEaCU6a72gvomdoQYU2UaOB7R3ZPLmXcAUCi8S9NMbG8x
GMrrNQTyD9akCLHjGvOvU8OFqJzWrP8S47OpSQUH+93A7Ik3ejJ9lGXxioSNEGpZ
4Oxq0t+JcbmnmUfsrrnINtnRRw5KfQSd3ytfrLBFUBXpVpCPtPWgCXClFuQ5G/x+
1Ab9PQaDyb1ZL5V/UAADttClyj66R+gF6MyBfhvoCVTcQTA+8vZkvHjQK9yuI2Dy
cYPaL9HGXBXKG+C2K3+QucFx8kjtskJN9lEsA3GS+PZv7eFdeDGmHoOl0oG+2Coh
fU8f6nAiD+c6+dum6Yoqj2t9pMkHK8iKNQc9OPYU9NkWtFF3QaOZ3L2BnCHvzvGV
8+Wb9fXteIBbIP8yE1QjS9vuhrM6LQObEeQbl3/4DBd/qUjbf+i9BdAcgtqtIS/0
u542ZYQKX+Iy9zgiVgzZFo5KFOTd0l7Ghddp899w308/PH2oo6ArDTqqE9NdVEeb
8+NYPXGSOF6TxhR+rZH1W8Plm/+d2rs8JvAISmS9tBuRUDFi6LteVI0Z8KHdP6M2
hKV2vbJngnfDksWObBGkTOpHUmXg+wBWU6qG31BER3UV5YBYFx3CQ/3JvoK28Kja
oopUX8YHJiXW4CGQeDPmKcujw0D4Bbw8RGPNbyczu6eWWsW7Dmo9wI6+wJxVj1QP
couiMLZnCDrd1nOH7LryOYzo+2wvxMdnaBJGO3azJvzoKT5MwribguUi5ONzxoMS
VJ7TRh9hC+ttqMd89QCJPl7XUHJ+zsNppGCM8kTfXYAIOzzOJ6+7X36BMS7dXlvP
prS6UdSAEcnSi6hsV4IElUCiPk5pLxtf928ShgTcJjAFqg6GCtsInDe6hm2kXiKL
jvKmkt9mAE2jCL3OJzqb4WTSvhNuVFVnwhEDLB7VJfQx+7ST5ybClTj7H1Ps12tj
uD2M5ozXwDr/zrUI8S4rX7mDMfEh88PZIXwVwNINQc9Emef94rknaxkgShlC+FwU
FPAXy/UQD8EMbG4YTpQE6YB7BrCix61CKFOBbmb919YQswZkqJzL9EUmX/x+OnZ9
kc/9MDlMcYbgAfHQnaEAB9uqH4pEbX/A7jpw6rg0AbxbZ+9kklAJh4BQbEd5C6A4
R6oF6k9QkmKEGLQZtXmGGAdjMxNGp19Ohere1pAPATNoLhiTtZtcCO6zNpEp1IBT
VHxgnm+JoQOjJvjFPcxaE2UcROXYA15gVL3ovI+hj2zC45pFKsV+1iQ3pDHe6nnv
VTLLpPC8YFvDXb621/jFnOYSy3hFGPIUgC812kKEoRbx1Hw0r4Jid1Iln3kO5g+G
4brQMr6G3EwBsx6+cJJakydOA1Bm3gQdeQW1oUpSuLwqMK5RuWNVX2SO8CGCKwlK
HYWLzaS1o2xm3w4wz4KEKl3yc6rmlbdOyMwHFROC11AhVxKjVkbWJiH6WSwzmna6
x6mNcnVePk4VnmH90iaXp1pYSKjMYqe8Iu+QlkG5lrM6PeWxxcOaSQVfuw2UPTwU
Hg6n15nHTnOH9IbAp93mTqhrq3Arzw1BWNNltQd23WOlf1Juxv4MpTf53pBpIfGX
UwtmbcjMPuLw0ihL9V3Pcq8h5u3IPAvEleK21PiWE42WCrzXt5COoEYK/u84yPeS
IDYs52MeMsXKYUEWt6PFhT9ZSN216a3UJzdJO+XFTELSncFZsQKm5rUSTy28ce2J
geMVDcMouiHX5HyYfJD+CMixgCMQjNgXXnQibZGyMxDGh9+p/VUCv0uadW5jHljy
u1a5CY3pF1WYJr08eGd6CT4PFo9EFnFxRcu8h5PiNtBUOVAvbQ63gI8mKBhR0u/u
5Q6hZOqqbik/xVAW7dimAd+G+Q/8XF/VyswdCcvHAny/B6l19MyPVdyLPIjiwomQ
y/aw17IDJwIDIMUEUcfmLZASj5/qcOy/alptvON9AKJqEOQO4RXHA8kADDYumFaH
uPI5x/Quz+cnTeJZnTFcpRwOJZ6pEhlkZ1eE/xja/k+Jd1mP5GBnsGgHMzMhlDH/
p1Stm8ao+aS/WhKFQ+dC5HNNxOcyE11VvS8dZa10d1XKMlwf+U6vEcUxQX2J3BJ0
NFjMEiT/2TtTVA0Dtoc+QUFP44Fi9k/51JO6ovTYdK9enTqza5sjIqDsIt/pCWDV
rdGgHtjVKZsj6BQtzTZcK3oCrUUWboSNkX0hxWE6s06LJn2IJB1WFjGGCmTI48UI
/5X9iqwDNd8NApH6GQh9QYt4J0v20vuWM9788/LvQEihLryp1Dn/bG2MyYLW/JZx
AW0pvvN/Xxa6/cUdAyvvu3YdZSsrcfohZQnty5OGqxIXk38S0kSxnYWcoE/gxgqM
RSnG0qP+KbsqOguedGzi0botDM92bn7EMN9EQyMf4Sox9TR01EXWK6kjyw8nothu
RaWYCniCN/Je5euBSW1yG6HUAtJFAb5vkYzqCGNeQjIVxKR8xhvmbeS9aBrWmwqB
59k7L/TMEY3p4sFXs9B0AOdwx3rdvixGEOGMpPAaOTnt5MLFMy7ip85rFkWkJCl+
TrkLZUscWXQr85hFWNQLpPNfRnGrr8ymXFrbyojxlNYrtSK8PiOddK+y/Jfysm3r
yQCAP6Wii7a+IuGn/BJUyMWn5JepqEAzJn9xuyILQ/SvQ0quFWUsv5cPJL+J34VP
LNVFnejF5pifEcVOWczNXOHRrA1hVNeFG764ByOU9aq2Xf4OKdV8oH+s2fY1LBMc
sy1yO7KJ3fVM+NlnCQ8BIaa8c2mkXb4nrK3iTpa/Tt+R9RcyfhW/LC60CKh38SEy
Mro278qv/I7LYulxv1VMr5LXxNDdi69oaVfDlxb1PkIFJmAbaXiUw686orHgdIlx
BVigOmvdS2ccLqgdAC3js2cC863f6CekK3ZdfF6XwNGbEMmrXhem1z2g1eK0xlSy
sFaOB7NpPiwCj8DAYw46VwxXo5BnpAbHZTLUWuu8N70vGC2EMr/oqQJQ3V7R+KRj
g7WXmCuXUS7jE8Zpp/eMZ7CCcQ+SL2k5UKfHCjtgK3jbzU0nxn5mkUoha1mhNVIa
REJmINBD6DzV3iwE8H87KFopTLdRyOJdSP/TtfQYAPDdX71EhvHTy097XImbncFr
uGq/rgT4OqJhrYwFD7ReWb3/+P4oLBgxAkCgme/Mw8YbR6m702/x+y/m9Vnx6asm
TtvMkcWoZbVad33TUeH0lDf4nX/v/afUoRddTLQJGwyEnufLpBt9q8sxPkxkDsH7
NMwC9MSiXiBmvjkjv9eW57tykANOAji44sEMpgc9wdjA1fMQJtMb8qbOirCAa0yo
YhGCWVwgKpr965NKeq4ynke1c2v1FOF+SSo6c9E6oZ+9WUH56L7XMolW3zNNyg7s
LPC2ytzH+yXKN3eGj1u36ycSALRUR4AgL9BYuL6MjWeLr6xRMrs5K4/eVNeB/wvb
AlRCOErIxH2XOI5s9Ib2OTsEy9bSbtb0ad0jwYBm3WT4fE4EY1sG3w/az1CYvbWa
2S8JyhJrMfw5hKHIl3K7ocnXjJdficMOo+jqJjzWNRts3yRgc9LUqkLempfofHpQ
QXIIiAlvgaoR1qYADfrkyut1tA82WCoPMkn4kR8XrSwypw3u3lv8Ht72W7Yxw6HR
nHWVh5Xq63zvTuThMI8SiPNlPOlMZNKbrNr7jAFdtEQWsow2UANp1JPwnsRG6PMA
7p/HGY+3ycYBoK6HACmNnpI58m2aHmHlcIuZipLhgMLVbC5G3kxgBCJjKRgrCepY
CmU49zn4JhNQPl/aamJhuO4VAoZWQJcNPrPc+RFoBY7i/ZpiW8pzn83LynaTb+NE
oFRxCoHDYb5kSZfxkMj8ERoeA5JFxv+6kPGvqkWR0r2sq8bNTqW7+NMikhE9wR9B
EySMj3hIAUJ1qJpmM67rGnka1UEmwC1xvDzN05FAvHuXGumtYiXXr99d49mO2cBP
o0+TWa2NJt/J3NhJo3gL0IFoobjbLg5rRJLCMgLpEiz/3WfPEk28asU0SadP2zOn
N8z3NNQIggyhBZHUk+XYt0Sg189KqvkCgS2pISyD2z+kzX3YO573ukGgP5CkGQdR
OJY1kxvb4jnBXQ3GW76FSr/PRbB6CoA6FNX6I7pwpwKFPLMDvgjCazWHjl2LJOSF
RFcOPv3+GWxRelQT3/WBUmrSF3FvZ62Em8xIFEJwmvUe6KisclZzmS709D4mWD7s
61AgjKQmRsIOJuqfE5avKp0hQwac5skX+grG/1SXI3M8/kz7PII0r47gZNKCItxe
BXMSPIJUpgEzycHhrOu2slewemk7DOBIbvJ4gGTN45PxjgCihKHTB5g8bs/etxzH
ilP1hc5kh+iUes8JxU6iKXcvPQZABMNRA+cF8loO0HKahyDuo+h8Qw8AViMWyC/h
FfXCgKOEFrlIjEHXkOULel1uiUIT0CvnLC1qN3PycvB0nsF5zo3XXggUDOtwOhSZ
Q0UBUJ2AXcDYN/ReBzoJSSBM+pfY7Z8x84E/Oa0dsHTzjOXn4n9mr4tOq7nriWQN
JofhDbhZWLa3gAIwjXL8ID2yvq8CH8bczYm7ehdE2anWHyRvyE+unHebxZ1jTuS5
95BASWtE83YjSH2ngwJMY9MIJjFwLGgq2cRrEz3X6VND+LpWI8CskZwmBcPwgH2B
7lc1vzdxRMT9I1gd1lYQCqDz1axcOguxtfiVbPD2O3n27/7DMYw73yc7bDf3UvxG
iRBkA40elGS/1D4BTe6tvvqSd19aG19Ywh3D9+6g6NIY6HOykosCCWarIt2tgy2n
gUHdhYGhZIcd/Jbucwkuq7uz6c7rGjGyvWqyhwL3DutzRhfyq4oqcGeDOIu5j5HX
SziqOD7QwTt25yN5QgMvIZKD40p0p5thEBNh4heAQUFZMK7SCBTuHKwnSxs/0Es3
E/f2qZhUHgeKyu9oOxAlNDH7PidskSN7MC1HhN/ykNZDRkZtF4GfGQXROedDUR8A
Hj57g4uOdKSSKtyUxqwNk7GbcCNlmLBOS2YFlZHGWNRQ7RvUfqvQJKztHRdAnH6m
SRxKbBZmLOEzDWHbIODcJOmfpXQxkzgVOYzZE/dzaSQ/eyvOQ6gzlrL+sXwvn53L
jxxl2YEOeL2LNOEXPZw0QbpStGiJ+7I0mG3qJTqIp3tXCocqcdMeyM4cV5RlhltB
ctAo59fCNuyBu1oCmw6qXflHj0yGboT1s29eCSsGPvwtXiuYapcnBqQp7RYqdt1M
7J/iN2breIsiI74F2ulxyHJZib4P+2Gc1vPKw0wtdfU54SHokN+j5lO6x8rWcQzZ
eVUnhWvyDX3t2TBPR9gSvajNb3ySh5wl7aQ+K2ZLoFlxCDanZrjuCD16BKRW7Xre
Tm5B80aHDf9BoUz8eHryCidZscCodVODRVTAJQQnRod7xmNbqFhDyDeGiGlSW1L2
1qshoOe3aJp9qapLXWzwrq5R/fScjdKso0hU3DpZEhVxIpazJwUCgZCb2tZ/uB4j
CorlaWHtlFrEl2f+6Ba2x/Zwhg+ta7ySnxdKJnP9uUehARCMrZFe/MPOUm6fsGoi
8jpRfdzqzxbNGTsAZJ0pv0nPiHN4rWdH9nmHkyQk2kJQ9fZb4ZPq1Yi2hvD0MB9G
PCRTV58QFOarkOu8ZRxjtmX5H73JjvtuuJ0smJFhVBY7NIT9bHYEwQdLja4QTuB6
Q9GJEH3aeNv2hrElwVBQ4F5Sr/scxRZPXWV/UCDRoPfF5szXlWQthmIlgubssKOF
U/prSB63TS/D2/mbkgPVoFZ38cwp4diOVFFVjsulUg16Noyt9Gg3NXjwKWCNqUvf
6vuEGRA9yBxkf9VBMwJkvcPTpiYbomTIQplsZtTNNcB34JumDoQtsFb4z03GRcFP
+jlcj3rNkObJAFwhbB+h0yLkdkY69O9LKIf2O5dtV5/+P3IGVcPjsOYuW3J4haLq
IoXbMnGaL0sdx6BtC9/Y4XbL6k9APRiPT05mGFYi3B8X55ZyaEefnntblF5p8fkV
swVz+6iLP6jOLtGkGdHBQYb9F0KpoZEBIWtiZRgXrcXFH7WHI9Zssr2h1JEQb1KU
edkK9unI0VpnORH0mNyQZ6FxA5ng0bWgDV+ZwWA/+zTo6e3RaAYen+tEZzTXcSz6
KT2SeQB563SoT1KA+LhbjdGrGvyjRMoBqk/1CP3jsv1k2rtUIla2P84nzvAHo6d5
DjtYp8ModLzWypUZn8exgqdL6JKQDnt/A/u8TI9RfBZb+klKr0YJpw159YdoSx+V
FjAoabWpbcbv3Xc0xnW7ihDSqjvPFJn81U9+ymGmJLx0iVybicZky8v6eUQoYbNb
QlqQrIcxI5MiExruGRiCWSXkr9o9YMc40aS/ExUc0muj5Pwex8RK4z4MTedX44Oq
upbXWGdGb3sez2jzDy7/zdNQFx/gllcG7U9EWe1u6DjRnZjmddGO0u4jjT+ZmpgS
k27okN3V5Zgo+zDoiDWEaGdMEtBLkQu2A4II1cbR1TEj1ah+0Z3+4R2YAJ/X+QPf
xBVLG/Cxedara4J4wQ7UVBIrLVa6XyQ+pk6/A0mbIyw0elK3qFqOYCaLv2MiY27n
V1xMu2BP6QnqkO3C8NkB0KGkELX2a5Dluo0ZytftZ1G2NLSNVdaSt0FFGmoPUoCg
09KoFITSEYuiIJBOd+H+IWmok6MRW3pA8MbMDgWKcJ7qjYgZ+lYo1uXed5HvFMYS
IsTMKkRWcaZeGsZxSOoWNtLla3fAIReHz6OvNK62B6C7C98xpEJQ6JlJLj0TdQ3r
kNBmDxd+xv04d0D1qntun3UO2Y20OoUjmZ7JfiNgAF+5de4a92H8YEl63SxNEGfB
HVAVbaZnLblekOK46v558bkH7PWlgkr6LvzjXKreZ1w/UHkeo9sOQISF4kR2JzPd
EpZLrwoeE4e4oFGpPtNVO5owItoVadO5Q/rRyxsG9Z0qCLUn9CWfsYI09jRKwcmU
u5ZXplzoDn/jVGEONeCBOturifK/Mk5PJSLiisdcarf2dZbJ9+VnkIgoW3YCr2Hn
9qD4umd1gP3W/LuZR4Sx9/ZXQ/f1IyOzoBm1xAWaFKgpE5jkfOR19GVvX1twYSzR
y7SSv+HlI3FvumgJwytrZZanYluIrSY+x3HJ8D+tGnqhwG9rb30/9JKzez7YoaRP
4Hxoi6SJKrV4nN0CfG+Q7WLuZEcyRQNfMzEHTrOtB9EHL7RRFxjLR/nW3KGmAI06
36MeL//0mA3yctPAKdgB3vsm434b5cjWSAXg9a6VLLwK4NygDa3rAb3YNaW2uaU8
8BYyH6Dy8HzoroDeRLnNiqB5ovdPlqQHbg6is9BJv3CHl3baTanaJRhLVBeF37Pd
bs/CHNe3J3+BPpalxotlIGHQ7zB3Ferkg7hnzA7+jDqxioeJkUkuJwCebivMylsD
pAvjemIl/GAqazsRrDHzben5eMt+VgUkJVXo0D2alb3u1rsTg2WegcRAKK8opGGH
SqacexE1DuYIDPgmlwphaTgJsy2rRDyTTaM5WSKZr/V7ZxU2XzRA/BW39m8QDA+0
du4AfhXwNrQ2DXphBkKyPr3EVUBikLUylz/uSfp9XoMiPCdOdke0bcGYhd01lnH4
18VdXMwnwdrXzmIfAokH9rEiHizsJ41SS/jX+QPJq/7dX5pFWPnnWHIpIqLVRk2V
sfy4AJDl3uk6EQIMp0LHB5ZNwRE39ei5BALdnUP9stTCu3P5WLLu/HqPUrQ/ACY3
L067H6Y+8e7UwGKrYi7vuOAiuwHTBTbD9xYKY8uSehgmAwjRX2iZOqW4R/EEYAsz
PIJeXtwpwd/2qN9D+nKJTf4Dfv4etVVm0h8J8HT5GMwtiXKU5HPkaIfDIFqOv5It
Kcfm4G4E0qaC/aC1QoSSt/KRPXCdshJGAwFzzxXYPaFC8TEkDOocCTS4geHzcavN
PXpd7aKD3gz9VwJxPD2wSE6jky1ygcw55a5kdmJ0pSdoG1/oE6eNLASo4iyaIMGe
qyQeeg6XeR+NDoKVoJTLUqP8fy69IQrpBytalG/3lOyjwCRXFV8QAJTqo9UD1fZf
NUwzeEtC93Icosi/42Glk9xfYX0J/fSc5E6MuoyAM1OrfkOccHColTYGhCOZYMy+
K4k3FY0GGn92T+yAhf6rBKzgw2VyoA5Nl78TtgFt6XrSqzQn2yHWWPwhpmDy2yXC
RV/08J08hp4/swtr/OFiTZ5WCjY2/wwOL8syb9j0WOMLfDkQdT+Ej2WzbM3j93Xs
m0Hu6VSV7uYF0S/9gCeAY+Q3zzYG2AHilirgOvKbBrXVRBvkZR0dekeV4hzCBuCq
nfHpcQcPU4jjKVMKJPBLDFJ8KEsbWGmW+zz81KYz9WVM5/lA7vVaqwg6SrYcWnH6
zyWaE/tEWwJpRwe9nwLWI1ODDpAcIfP9I9UHPXxzkZzIsJDePkcdt2P4yTxJ4oRf
QIWXAn9QZjEmQfOAtkMNYFWbPd7afzwvUmVufXmX3Kzo/blEBjrLMS9zIpNR4XG5
hbX1X+QeeoXr6ZFlwCBfgSMjaxaJgfrrsrUSEHA+1MrlkZ6oKez93wrE65oEnODE
5Jr4viKG+l06kCh31RQ95zGLQVrwvTVGfzZ0KT7JjrueS917EWhaeYDvLSspPfHG
lUGUB9mdady5n4QZiA2CzeJwMIY8SZXL6WGxz6uI4YMJMRqktD+jHftZU1We9jWy
wBjQzqn1OmF8mnHJAYHXpxtG+5FblraHpb8fDeeurM6YtCgCxMWwagfRxrNycZzj
XgeQV6oqi8TW3WCmyvZoRJifoBldMHvgAc6Rdg3SilFezG8nuQ420sPL4X+LKbx5
HOX21OS/Y3gleti2CNVZx2FlkPfJqybwg+Kojj7Ogv/h1DWtCiTpfwxqOSQC5JRp
EbxEQnxQbV2WH1SagV+Qd5SW6BAAw/ALlV7STTp+OXEwwAibWJ28E6nxmA4AYfgZ
OvFo2X8G8Fr/IOaYoKNK6IjySXc1Bikpo1qW8Asss/0bHH7p51lqxh81FsuSpMxU
Lkq3VPLqzVfT88EZCi42TUl+KGy8mvWfqK6I7Pxd13iVjIT6U7EZUQ19d9WWgD0W
9dmJD/duv3BLx4+5GVJxpl6+/WJngkuIPHbP7ZMCJB73+hS41b2rxMqxQdnhyHEa
02CdZtI/VQEqgDMvTNuvWwLMO6bwl/uwQ++hXeS00D0EuuXjmUZ7T443G2xLiS0S
2o5AFNItzVYnol3iwqcDw8A9Mgvw83eOS2+ARAXkCvA2vp+uSJucYOjvt0QB9kID
TfJoFL+JE0oFSGCCqohjn0cryU7+KjnU/xL4mnEMelg0F/Ld3mkI6GGxW4gVENtf
2IUv5KVNxdyhEH8UT+eimOF03e/oc6s/GmcG9x2/JT9weJVjZWMOQRSblbkhd8dR
j7CJYN8yrbTT7sxwjQivpXCP42xtXUqXZEVUNV5pICfrJjTVkR1dx5MYbFkjE/iW
lueZZVjyUs5vZtubatiwQOPegaa4i1Ir/tOJAjTIl8DZSnKz3YSztqix1dI132MF
6x8h9KjAjLvITNCS2ymeq4KNnYApa9otdky+sflbBSN3e2COtbVzCTVGhOcMttvZ
TLh4CiUzomhLQn85p8sK0CH+ywZuhsFxKVimlKHoIHtK3gFFqGFyEsyDMQZJMZEq
Jqo8qk2Gkwg0EIyxVHKPgwBIhp782QsLJGWaghgdAaJJvqhveslF8rub7JeLeXhv
3HM7ZHc4nqKzZ4dj6RIP0+8YnIUSGC4VEZjnciueSdCmRrgWVXMQnmfO3Nvdvbie
fGitdY3XBYt8PeSypv4kk8A/YDZs+QPhyI322WX2W29/6hj05bi+1XHAHqDhKBpn
OZCx8d91B/zv5sWW2M1hW4j7e+DDWqBNhZVXkrd8snlNaW1WzKNS03AnGblaICyJ
6SDzlIiu5GOaY0w8o1zOjCw04pSUIrKLRm00t385IJ8nz0zQo3IuomDqTa5ofYm+
VAno+uEiIFPzKj4s1SSi+4TPbHkNCEAMSfpsL+5v6LSeGjXhvfaScGngZGZZFHvt
N9kbEpBLdwUeqZ1qXskSHe/Sa6RyQEDLSCkPfVFT6IO8s+v5taBP528jKoL/nAzb
jHK42z3kxdcrZDxIfT3DwACCACfG6Blua3+1iTCFIDauzALXMNmL94MftibgsWG5
Iqy/Y2oxA8RDKvoWj+4vpWaLGa2vKUhmCFJAi2rjC7RljP3G+gf1SjiIg7yIBFX7
Jh8RcYOboHiWOI2Vqdss7QPXVgZltQvKQr8TvUEzqs7o6HqlljHWChI03ElcV6iB
7muVOG+ab3qTdgqJaCX1i20Rkb0/12rN4mp4dYz+BkHQIb7dYP0UJdMeh4qIBuET
jUYnjLOpHLANbmHDYFf5PQDKIqF29BJay/c+8uBLvhQ5RJEb1I3ta7dkpShqcUUS
SDjJRxL+LMNCVrVfwISp2juYmTyAIG0QoRdBUllE/n4NysNbuHc+9D6V/Y6tSNyp
/cgCdh9dKKIKymlzj/Ee0qrPkVrJREJsU1VGSMnpQn+ehHp6YVCgY2gUmDzC61Pn
7TllyOD/SerRgXfaWE1rvqWGgnpnnVASm9kTnOnu6wLuI+onaE5ChH29AIRFYiKU
BeR06Rpij1FrvhG/pBnWrfMn+22DM+zp9bipUpTK8yUPy4DbGxPTcWeR/SUA4QZQ
PQEbtM04ofCwlfvs+8446nMq25M3CyapMY7xDeIQxRkTubnBP+V2xwuJuYEXlCZl
V04PdJt7Zb+bmZFzr8nAXm2Cl8Q0EX+PcQjGjXLn+y0sQWPJIswZLUuqAiKk9eoD
MoKQukUn7Pgehk+bcSzjapPURBJSSAsc616X/zVEbEtn4kcL7vYAvPYNMun2BfRz
19ZceWsIONVTl0OCJQgKdO9kwVmbn5QidEYnqAEobk6m+zo573gBUgryE9V9M6mj
KRyltk4Y+B43XKhKHD+Uy4A9xfHAeJ5wSLtqYapdKMZE+68uzITwFLOvkS+0OLSP
14ZHfPsT/hDeG6EHK1DcIv5qemzj0qq1q9ckuqvRgrDC2YGL9HxJtIuBiqvQVONp
HKiHdOzDQ7+0+7fxlZMtJY+XE+ffzNznu3PdMCyIZevHSDfI9WSsl6Xvw1f0mf8I
CatyD62ISTzkcFaXbJUvYx02tjC4vnR5xw2xeWzGeHQyJzWIAl8PMK9D5e/sb8mQ
qju8HEFXhlfREgcQDedzydksIh3JMD+NqzsBM4SOaqVVTmt3VpvnbAv4Div2hWKh
70IJaHqiOWtXj8mAIKB8Fh28JqAHbUdm7mN3qEoHd2hseGMaTB3wElHWMB5dGTiS
lOmJPa2hJgl9xXSLG42Gn6pXahk4GV13A+v8CWa63SRZVicEi5MEQbXa149QBCQR
mphs4+1yun3FdA4H5pVoa7VTpeYadlo96q0nPpKl8VtqmwjEhHxXXb7y+oyynJ4D
3b3G+GK7feXSnvYadtZYp+Bq2frlulV9UHwummHvd8Hf+dtiwcaJCOx1vPa/t6X3
KfYGmiVvdWz7ROb0dRQ6FyxtDC4dq4jlQRjaeZQwf9dBTg+4c5UD5G35A4nRvv3U
MXWMwMaOT0cSwxx7ymcvS+kewrKviCrRTtEMm4PJdLc3bomHE3yOs7C1/kyO9YKd
8PGRAqBbjGJTBSwWPftf+nWYt3zvIoYumS0e3bEgUV1NHlm9JAZVTXAtJ/tv3f6W
VennhDJHqdrArvK2hpXQb2TioelZnx/vNdb/d3itErZ9eYo4CwUbUcO2NOgy9q+L
9xbOvz+caPqZuoXX7e45DdPnq/tCQnsayGBV97mBxG3n2zrABSbt8u0YMW36s+mV
qMz5RjpIfdn7vtkgezN1qN9UunnzsnDUvlVIs5YUB6o0/3egTRAdOXCd8QpJFGo8
aU3GwXgQ9NSbFgiuHm98DpsUfjnyr4RGD5vy/VSa4o4kZ3F1Zd0QOLIviGQjLlHU
yCtqUMC9whIcNgaOvALSdcD5XPje3r5AQv5zfUmdaAcu0/rky6/RCMaofk7BOWMw
gmif1/+6y/BGW18anOlISJT5DizzyHT08f78obJd2NljjNX4okthf9aQ115QpfG/
rTfSfATjDZTss+qriaGggDLZHorWNSJQhrOoy2z0XjdvX4OcKUp5V3H2xq22fE4h
8DC+Z/2UvScSNDFGBv43uK46moFVhCa8bsMXm07wowTldwiBnTh14k0Lvk+o5C6U
tniGK8LFxLQ+o2NHnHCr6RReZ/z7VR4V6p4w3AA3K5sJ2ITlT336AUOFh++O5BNX
qj2QQZENVeLj8cNHrioTSyCJ/CC2bI9s/1EAbJxRkv+wcWhy+j+Jub8tyBa0+kp0
FyQTLEOwJJWk4TaOKsVGHJY/ucmQID9oEeeu1Mjar+3ludP241Mm7b+qYwcf3nFm
d+9+pdbo6KULXsXQOmaVscJQ0URoxnP0yIe3nRpHGauwjUWTzIYvzDWwoVVRM63z
lfAkEwPI5hZfcX7gCLSLWd045hx6eVOuH/LisMwLZdvqSCWq6eqCqDrrcNVXV90f
MXpneFtL701fvQ+UnAyRe2SVpo+4XRHxn12QEDZ4f3drNNF50vvrxQ1HHfrN27qf
MtgQLBdRG/bT3Iiq+jTqd//JrGHN7Ya3brVVmzNKufiofY1lByqr8lGwt7/Fr11w
aDN8B+9JZ4anlqftmpb5CPrTcJlU5pKGWG7NG8e9aCDdyyrReX4PMSNriTBgq23q
GMIAKDDvz24HT1HjVSCRYaK4Wnl1KPCDzJ1DWSRA3XLkAbMyZ1BhJKasHHbAHPUL
qBTQQjqFFRO4GclmcZuY/QF5uIvEcmdGiuPmSorvRaupe97+nmrijblaZNAMcF6G
NfkVwRFgiK+R6HUkiTqdYZhtNqd6/Z4A4iKdtuZbiAEYfAz/KEJY9mkSCiJwbOke
/pM3Xpo2fhk9sCALbpEzxBK01LFnjcB4zyI9anooi1/KDdh88S5wubz0jH78Ccbh
ZdwyKxjEDpWC3QwTZZxMX8K50UUe2pxu4b9Me7m9rWlmUGcnIvBQtbUqWLRtL/f6
qHyj6iL9Xb0GykUZdnImd12a+J5GNOoqT3jdQ5nzY23CtCJ0gg8cHUdTSFBOr3fe
0pn/vpAWKcQnTylTMYL6JL8QelbHyjY4kSFpYLHuimk1Zj4njzy1R7H8BqVaJU7m
eQIT7xOzbqR7jD8T5cfKf8GdEMBqisV62U0CZN4I8y6u8hmXVA3zrbd8xq+oG8qv
4Z7MbHmaszsLTSloggpqJbcGLJ3gL3HPXmm6/T5/p2Bm4EWDvy1pGB93ZRoCkl9t
/DiO5rdWKPE0cKK9el4Pb/aar9QbReMzEbJcYG8j+qrMwe1qBVce6CEL0fq3u1Un
FiQP7KRUxbxZXvH2SbHQJcT9AKcYqerG17ElnfHCCqf1YLxGQgm86jT1dcryBTMk
T8LAcnyUMUV2cVqSfviO4xE3aDzpR1wa/kr/e0kWewTH6ZYSZbz5Wj1ImDemcumu
dY1nI9T+9yoMpO2gHzkMyjmjdv9/pX/OeRQWi9bxK0Ly84rP7At66wGSLnkVS9Xh
1qZbmwauYz1eLv/x0A+TO3Fm6MweCw9IXWqhr3Q36AxElrL0sA/y06mfz1/w4IZO
NTz0nHDP/qq2APuukGZQQE7uAQn7BV0jZ3K7nVNxqOFXBwjg7tR/Js4NRD1SvQ37
N5K/Ib8CT/Sh3AgaOK3CjxWe97PEmNRFiSpLwec9pz/1fNik6fKVLCwXRg8KByVC
bUDDvGKHxNxFOWMNCPbS60sWiDCBSk/DQZdLn4IJmFrDM7IEPgkUJ0Dv+zkbLHpj
DaXfPRriqNWMwhEMVp83cfwu2nQJYwIzFs2YJv2Zd8+BlxQDqi1k3/zRekUPaoLd
7SSpNxRpsII51+qw8Jjej6Usbq9XBkACKSomFbnhEo17G1BICi5C7Zcbx0usb3aP
wj9YU9N5i5VKww5tV4Rjqp04qgbAE0oTPl+RSPyP+JqIAPfzr1L7wa6S5oE0qyHY
RCHlVNRQaWkqFwgEspr4Np0G2ESPRTAft6gJG1vxdrRJu64yE4cp8ZrfNyZsFtWX
ZSecgKDwwCl36QvjtllqlJ2j8h0RbCFa5CTMB3ABQPm2ntGKr4buTizRiHpDDA4k
+Nmpv+jnFs7VjUjCBnjTNm9LKGa7kwe2/TqZRlWWVTrSMZeTjgL09YLP1MN52p3C
HoDVq91DRhg4UPQ8f8Hmy6p/JDcSAooplVzt03NFnFZqcwJO1fYn1aafpslK7pU1
b8uYjRmJaeYnjYYomR5wugC7JnEtvJbgpNAHoMJu2GPNUfaZ22qLYxxo7twFw+Mt
w/nVToPTI2sXQEzMcTZ/tqQryWZgxEBxz3sdw8v8lBONR5fkshq1IRrbXOUt/o/H
mk/vkk7qmkEHwAMQUPyNsbcfGg798iKQwK1zSklE2eQ9Sz65WoZX5piZVOSAD1Gi
GsdzP7oI2wFwwGNGIpc64VR2BrHnT0BQOT8nvnM6bjzyBlmq/KgtsVFwnUWehnmY
wILuEK72dPcpKwaksPg8lj9qAY9sTdDhtdTj16wzU+YjnbPnVZfvBQ0D8qlr+56D
krnnk13/So+sfddgeykuMtveqssI4IBonyW7XEk05nb8j6PiyV7Bt5drbJj49X/8
wrXcjA9isnsiy80ga3vSjWMy+GXHqihe33p8tj2Sf/fFA3wa3Qf+OKyv10ZwZQn8
UqSXdGErv+rqrlIG7ZoJ0DFRTax898bRk7oYvwtq+1NRRNsAN29US5O6jogeXMWJ
EJWMYh1gPx56o55NnGrKOvCbSfx2NJ8a73h8Q7w27n6v0hYEF6Wdw7GX4V6PLbXN
kZsSjXo3y1XdUIMWPXw08iaY4vYM2spNypIisJYYYsgQEAJaP+UYnHRmZjQYG3US
MzwadQKdvCL9L1Y3QN8VrYolAp2Qdje5KGLMJ4PqeFuA1k+gJz57NaOq7pGKm0BS
Hikh5BofccXAz09FZeNJjkGPRlrqRQ8dy6PNh7iHQzXlLrJuV1IkA5OHWaoUW3s7
LGh1GangTdbK4Jt9ciBbO2IA//m4eRUlKE/FjDUzVp1RQu/JjNgL2TFMnORud4bv
6MwI1qS5+bvuREYbF0O61svgEOmO3IY98A2sLQYBW3/OXt892Mo6z3O8baX8lW2/
ER/OXMFKQJ+0J8RGCbaGGJ5TtSeTSUmrngZriH0ZG/TljD7kIOyPjeRsO5PxrhX6
RVieqPa+OR5KRqU8t/G7uNIl0I9m5QsXXZroH80RdgZeJOXauikngAKkIP3D9iOs
4iX/t5Onfj64elRNfAYhNjAcMzgUUtSJ2GQaPhYuFpQ4nCbQJCrCq87eLDQ8xYH/
+qi/00YEfHflpd2TlNqDWXOHqiqnFnSLfSs3Dkiv4IlPjpYTjcP1DbgT6jwsmBGb
SueW0REvJbNnnzDm+mFveUQdMdU1X4oWg93bcUyknoqDJ8fnV28qgxelh1Jkby+9
jRoUmlxMXORILemEUqgXW92eS7fIReUFzQ6x6h/jyHq4n+gMIAbjLF0+l4SSk/2z
DH37J8aNfLMIJVK7LUEJVJ759JiXFb4H5PEU7gkfdWzSJdd3SfpDycbu3KiSdFyO
6+AcYjv2obNNo/I4AnNaosqTJTqonYAwnodsOzbsLbSo8UjRV2osctW+NXdL73QD
WEsIKEchxiOEPPHvsEMXs5eo/qdeFZUpgl7vgSofOoqWJgtiFZaBTweWovlNwzNu
nrjE5PSVdJgxhrkCC2XnklbVNIb+CzViOuveWKrGGwsAsBaXpjjD0eMhqgyeE6Zr
B4oAEG25ms1yIp2mJ1sjMqyTIIYcvmuBG706rpltrrN7Z+JXDzAv6GhwDUyS3NSv
2SQTeEDJWFpQ8olsYYswLBrUxq+iEIIGuCeMqg47ZNWpIOfkmuaSs+md/zMempID
Sr0p4/pIEWU2sLyy56TXkiaOkbFTJ6X1aND+SwGwhFyOLB7ORLh+n4QwtfjijFim
c85iMjGPaAnMWu6lJZZhWpl/clwCRuPcj1fXLryEtOs8OhrZVs3ETS3DLUCAjNlc
dZUEBQXxOB1utxzfuxgHWX3hQyt/wsozSWqbm83h2DmenJHoyu57AqbnE7o2sT/w
SmASFwRSQ1AQUYPYEdCAt4jOoWNnnbc2sNfKhHzezu2tDo000W80aPd+9CXSiKRg
szYluUYVld+G96YkmgRSxPaY32Wc+7/5Gtu8eKA6ub4iJwOx2aqFuWbuQ7QxQOUY
gyLDbESUggHGAA6t1VMGSUn8sxkGSAEwAvwb9uumky24yUQZm5yctcv4nSQ0zyEg
PEYcA9YbqMhfEhVi109dBClgUSG/wEIPDlM/LYLzzxbdhcFQ7XWuTgt6+Ajpbd+4
hgiY7Z/ScooAD7STdmN3JlhB3csit8X+av/KBElXdBGTuEJpzlflxhLKveBCfDEk
4Sf/HB0bP0bJvwfNlU7/9CJjTAQDM3rn4iAFXhwX4iEaU8+cIHZC4T+zmemEVWwq
R1d/EqgG0JKA7LcFYlum4G9LvNC63CiA3AQw/LxU8F1Xr/v3qGBbrbCXkJRGhRKV
f94EVlhqyelJBknkCyrdWBWPr+QmiclQ8mOWVVqKT+G5P4atiCX/L0u9asZvP2oj
tQkvecWGFPIgHsYhJp8ksYQwa5mSmwt+mLfYHuatq1uy22dexGzxBw7pIwPFNT4N
0sPujrbUuLiRtayf3j8NdCN7okOVQ9OjlOhzdhsbDqLUnwblMGTm50A6muhHP6NL
BNqw3tCpxDTnKwLc/OESwMJv8Zc0JV87tcYL/gEG3bMACxBeUeCabo8lRVzSF4Y+
uJsTAmTZnHT1zLaKKC2uc4YhhTOQXo9xBTi+grQadr5DldJ0M3zbKfV7roYKCN0o
fe1cFG4UuS2/OCmWhX8ONCS1pX+Mq2SiiYUQIgs8Wamv4GinDlk5+TAP+Xmrf6P/
09PW2Cwj4Q/QJ5IZOmwZfuiMyHIWAY2ObfttgE8XW19I6EwB6sC5VvgldOAPWmYT
avXcVCb4gDfKgw+nEyxDLjgHvnrYT+aTSxTSsjj67f8Wj/wOInleOJ9EDSA+N4+A
KKU+wxDSt4eexlwflZeWdsivtfJh9m6jWvwGLA4D5RHEE36+3r2QqmXaX2etD/na
mxqTwnRzwRvvd5pgOenpupzpbH6xFc46II2dmlrjw9dUd4iS3ITwEGR9G2yCuIOb
jl+A7sWD6gC5zko0/T8U7TUqkUb8FW8c3vRGgK7F4/zXIXEAkyQ3IKo8+nEI2eTW
3hggMABC69vwhenaJV/fuQdlkPL69PNbfng5s2resAw4AAhXqx58LgiKg9avrKw1
4aPWoDWBTbg+f1KHb052vvSpdYq+CWP+8/MMggdMTcecjExolUXRg6zJtWfwWfPi
wy8JjJ3IFJ2wkJkAtd7iq0nrbhwyDUcvva34RXwYxie0LGdBzFlNM9gjZoWopkac
gVyARbJsI+uVPN1cYKTWs1MNaWK9QRnIBhYl049XPGG+iueHdofwguBXROgQbDH1
R2glB+aFj90zBYSrhxpG4oOs9ZHdktewqOXgJxFE/UxO4LIfnj5i2/SFyXz12lCO
nzA5tmXwXr2Bk9XXvmH0tkSNqfBssUfT4/iVQAu39QZKN6b0rc3UxttpnmDx8q9x
lX8f3JK9PuwWkkVav/X4gCy/sybDt/L+QBSDDOQdEh/1nXE5bDPSxJpwk03Ofpr1
pIAf/dH2l0gGxUlzE3lpFBBpDCMRkqSKswN4mLFilQdbV3vW1lc1MxJT/Nog3MO/
k5mHQabOdJwxQfcJTxhrtYGZmtY2tujww8LCcmrPIwiM49qlU/tWrJ9rk8mNY7ki
WLFYZF1sjx63p1tQJWnlCVUMiMe0AriZAeqioHKqcnJZ5DRyhJ5pEnaIar4M/36T
nkUzLc2osQAn/YD32sTZaBjE0DXqAiKrORoyy0f7M2BdFhZg0JdcTYh2kKq0Mm+F
dkCnyRsxgkdwiQfJGj66BPLjggwIHo8W3iYnw+Gb5NYlBjrhdSoC3LxBDVrkAIEy
2tWbogwMIwi92Pe0RAoU619mQtH8KhUibzU1KQxjZZaWv4E0Tnzsqv5UXvTUgJki
DZaoHpXBYAyCrqBRDeviVLLyLfWBDL1eowyRa4HipzYE9AiHA6hcaiuSc0lqg6lh
4dOuEqcI5+ESrN3GknjC1nYVdkls8O1d0FwhX2WItQvF79MysFlFjXSJUuabmPIh
P+/GVDjVST/u0EZO5RaRESXUFHVr3OL9J0pHzKthC3NdYWNGjp0Wsg/t7UK8ynv/
T2drzh4xcbGxkJr2Z388WfHjbbFZm0hO2XAkkzeWFnfhEGFCtT6e93XP6wNOM4C/
mng5w/9jyi7hbTb4vUPZ3N3L6+MaubOGh+14937KjBpyjuyYOfZfovN5rAx9fzdh
htvrcHmzCIn2NhuRQE+V2vLbvB8svsTc7xqGKdsffn6tRAoWv84PuYtOEljIt/a5
AxTokTtwxczW4S58bYdHrL+6uo2/WX7uW8P0S5Tlw16cqOIk7zPk0UZ+Dh161Y+/
7A2TMT12FRyoXdTXyY26E/01VtJls5oK9Br2c1EUIbQ/PptC+y6khLStni3Ex/Ye
aRqXLfO4KJ1Y2XWHHktCzD88jU+tQmE0z7hZHzk2O+07tHJ0GhhKO3k61z3x0zm0
lrhjjJF/MYJA5sO/+nYyCSrEosts+CcQNEzAFMT4pOSiz/Tsr5OCnF0TYn+0DsYv
8xltiYNze77Hu9osB3qF1DTlZb0ruQEqEHG0hjLVIxqH75GjstgcSsT8gYx7XtrF
P6JXfnsO4rcEOfrDOoGMjERxX0Ot2kOODfazAuCtqf37eiRAO/QH0ZtZrpVo1n1Y
Q8Jg9JADngqMW7deV0Y9PrHojXDzQAu5rBqTjC6KOfeieUOkTPvuezXXsrqI9rAY
g/WsPu/a34zAHNf2K5J0MMGUMn530PB2dEZCuxYsXCF6c0liMPVMfLh9GLr1Tx02
fD2ed7YdHnz2XA2z90jmg4ZqPAwNN+XO12dvHsG+VYwiC4pVHN17b+ZDSp7BOOwa
QHQKYrCe5IB6BlSsfyoAl7ZRIHDM5fTtllGU12UhAVQgrFVXjii05Kr1cGp+iDQb
90p2y3lYxOkiscthlp38KiORF98RDtVhziNBsjmk+IMQ+xrE13tAhVDSIy4jwmrm
zj0F7yYF28rnkR8/bRdDUhk4d372MmMKrE4afznD6Yc+Hp6qqfhU56CUjJt4g31H
Vgwu4uf3NLRwjt2GAWhex79scV2Nrv5WDeW7D5IVhKK5gEIz/Cub3akNc1eDCwvr
Jc6m3Gzr8UU9BdeFgfrzcgl28S6XDT6bDf/uPxyLA51j2/rwfuKaS25WeAQVJs1b
lhZPCMWA4lGFsCYci8m6Ywz53ifrSvFZ/i/rb7eU1YWjwNy+NTzrZ5TZ0U0qzR0O
DhCaybEmt//PpYlCRXruALYegjx/t6QL8WfUYE7Askivy0QvzQmdxDc+MSE5g2R4
TnaNB/TnZpj36UkiT2sp0AgW+CLuwiGwHTqUCDtApFbbBGGla10Opcpt7Yc+x4OX
dUBZd0uU8ODHJ3TgtrT9eSUHoj1Do29oxwvXOYIfmcLMQtDAmrFxDCvqGqOA0bhc
NFfeyIySVJ+jo1qdvz+IR2csAZeDeIJyzHRT9W1zyapnzKgx6xCE/wVcPUl2aHYx
gAtMPh8X4kKBOswVYldeNWI92MeI4Pb1KRxW5JO8SvqjQxOMQdPcnM++wNC5ILBO
Alx1Yi6Gky6dn1UFLs0xoxdLoRJZ6qaTtvUQkJ2bRTGnB206Y7qDeC7sXXe0AKX7
l/c4b6gtDCVATvJnujy93ne8a1kr1N5b/EoEdfJj7keFt+wgokGHWyQDp3MuP5Uc
IaR5FGc01WhrXf1e0TlzZLtomPwUEfCPPN4IeeZLdvkCx3rXbt3qbqyAlhYh7D0t
b+F0fvU4t3QmpscUkAaGXb6NvY55VZpfr0cA6//oxSGLsTBSntkpdJGDSJPPEODe
1dBWKBS4L6QKt1hUGmrcgX/EEd66T9X6dYOqdFyKyP7JTG3ls7Dp9G3DLaKt/15Q
d0vdOpJ+beeaFRwTiCZU+mB8hA/WlnIDYzCoc58VdjpfXo9/BmrHFrL1JvSs2FQr
pltwsUCc/7C8PaBj6ZiRbLs2j3F3W8wYfeylm1CWCYqt1S81J3JpSQ1/HkAT+xbo
kcUBcfZrimk1Ar9TS0aIsUv8ZE2/OmABpSZfxvsIdxX8emC8JvQegfOm+etAhaHX
fSttB7a+pNx5qSsdrER9r3HGJNu+DhGi41KZlKwInvi3dBRcQlw4vTGaSROAjBqI
pl5qzngXuGzeMwvGJntAq2QWOqmKbnaKqQdyvGmaQBui8SkncgVv4eCa8kYZc+E8
3uZULn0mHPTBDiokc35gITnNKCyAoRDU4iWgKM+tyy//V0RwlT6b52q+1tvRd0g2
gYvCYNHTZ7rHvuEQGa5QyRgiNcfSXP9wsWj/IiMTee+lUa0b9VmoSHu9QizM2dDl
SWJ/ipqR5isw8FGLZAcd6zRXGsgwUg9njRVPrZpcpr1IibJEK8ZO5Fy1k6kC042Y
2qCH+lfmY02kmUSr/KFVbmUAla/1fRKhL1kSJslTaRhnfpdz3nVfHpc7aS9zqjBe
F8UqVjgr4AIIXWGcT7WQS397JWKcTH9qnwTJ9V86ysPBiDtQ1t07pXDEFxNm0c8K
qFYXCRdWJZ3OMyfWEUiDNbDIH610S4rM8c5Rfw780AcjjPv6Q5JGt88FqtBQyZ7Y
5LPNlGH92NQV4M1uTxsJd2FN8RGpVlRzZWRQA+tDr4tap1CsQymSsN/90NaHmPIM
6vSBts6BtvJxYdglylyxBenqTHYl67Zu7vPYBZ36KR2I0/DGg6PwCRTYRPbAEnKy
HaDZfqJ1BwET8gkQACUAcSy+C6OJpliuL5CicxahbBCEBUxZxzz94DMSGAiuVBx6
hDQD6O4IbFgVIyxv+HuK50pOgGbLchs6RLKMY0c0BmWJ7FHlMLpmujrU1pchAItC
onGJvsuRdHfHdAkNOugle+yiYP6Dx7i6/KBWd0+vo6YfGUaMQRyIlp+1SPlOacfz
z8uSTmrcimxyDqmGmm8SFm/vfO/3xNKYdLsQF+/waKoTgiIGaVsO+XtGie8UZ+ke
qYhxRob36u0NZB9sjxAKId5e88yQMR71CTBu0ec9jCVmy0vy1TmGlK1wV1BiOac5
8Zzy/s0HxQHtXhyVJBgOlv7AES5Gj6oql4I88EsXeVB79FHW9cbUKh8XhAbJ8SyJ
SmCpxuuq7OoIIi1hB5S6O0/pAk4F/qy8PSRlwVYfvVP6wjlpowQwNfDBfK/YSk4B
2BFRBHXALxUVPWZlyaPSlehD25Xdi0Xx0qWmJcOGndu9/FB0NSd4sahLaIItUQhj
tb1n9AHYC4+cpUqNoJ/LCJcf1nlUQQYhve2ESrNw0q5Dpd6imGOQ65BLAx7RS+HG
7QQtBeHAzW07H1FoRalacpmFsWB1qEjNVjIcxql6ioum689oImpznuwNYYiL2oqq
+jGpHbwo0nx96bfCxw29Z/1hhOcINiCvvAEqJwkAryvHMmB1LRbzGa6IG70yBM2b
TKDcIKmb2j7BhxQclGG2kb1TpU6Dlj6Fg9ELOR0GgL1GsWi30YaT0AlunXxB5VyR
GZXSSYRjvoTj8L0UrYYBZHlnsKdiPUXa9rIh11Zqjw/ctnKJjIP1uhJZ29hlDfmX
vdl7uwASFHpyWkIqddN+Br1z2y8wIEDc1Xp6Ljkw+djCZ/GS2vt6LNN3LIoMbBch
frO3RWGwQtEMCcp2+IUPSzR2kA2HHULkf71q4RnYz0bGBrMuEaMf5Ql5UfFY4xFb
NocWLHhKXeGdJ1o8LpmKmA1KpcMkqkaZaZm8C9JzPkozeiTauGoYBucb64jjV9iH
r8x7phKC0mh6nw4lonbIU/tsoLBoZ66xlM10BcKVlV3UDzJW376xsSfbvc9F5pdk
BLqBlFH66HvNgGZa5i8LBmjNBhsaL1ogxeZ5/ewL+kSUvopt++iXEcRQmIvtsSLN
eK5feJgO4YYDIasImwvATM0zR/kyxcO5BgEx5MzFQv7zwDPSZCDcEu4t/Wo5fvGy
Nfv8l2uvP7vPOUcFh6WUmn/yDvgsEuTXS8hChLlIVTRf3lwgl6gPI7FdjvG3YRg9
MXQQLRVNd3lM+OMhfmlWk7o3J+emMSVip7XMJEsZ3S0jsPnDOUurfAMawLVWS2Ho
Qm9X3V6/INxPIDLENsPge9tX3ktHnZk8SUMYRe397isTatOquxY5lLie2uNBbD0y
V30/vs8mrfyJfH3EeBpgqyXjs7+zHNCevHrLvv5L3wzH4AB6gyvThSDOzn9Ah6kZ
YMkIIsMoSTO/kGlgfJ2ARom5T5meDrWuH6Dd5rxajsnSDUhHC+gRkBU7xrB9XbuF
LnmiYuzT+ZGN6cbldmdLmEH6UB/Nktlr5DmsZphwai16HcSawfjVy+D7d3wfqB68
ovBn7hp+GEw3c6kpVmDVViFrkqGB/zzMT/XstQIOtLHTeDuI0qfIMTTA1pSffveK
IExYZ3ZcKJ8PcKX8bLYm9xzGHR2d+1czLDGHATHahK+LBFwwpaHWupYJP51LkS+G
1RZjjx9AsUNN9yAgvf+X8WNHZZ1Ne1ZNBUP+sOVYD/RHtil+pzlFMDy0MHGkDxwW
VP9XOJo7taD3xxK7XSpB6girXb5mZY7M+tOX4RcrqRXizRS6om6gVz7EwXsQWzoq
5YsJ3D4EhLb7diYImQywCn+XrQU7Wd4mJLfv6QROBLjQ1RqYHjyMvHnBloSNfadY
3JYcpYUEAQZBpbEVNpurDKv1oy/09smCCeJm6ErRIp1N7N/PMxFwhy2lZMtOpJmq
wSCPPa6/QK1vLr4of6xNx59UsEV6sbKJYKopu9dFIUC0kP9lV70CrpniPrAhPADj
P95chrZMMsPhliz5O17LSLhCEGVy2NdWDascLNqkb8QBbN7p6yLR5fcXPY2StM/r
t0UHAw/OEFLk7V//n0tGbkdwB7hwH1sKIOz80dZnIfrbq+twiot8sQP5HM6sW1kE
DCa4Alz2FnEag/4aJo+RdGSetX7NCa92B7mi6Yxd/wpCr/Zc3etDBD4BJOGW90AY
cy/F/kV4NnIUSbzBg1pfYH8DU8FROE4AX0Ls7sUHDapYqIJ5zraQwfdSzleo6ZBA
Sg2VT0ZwtRL5EUp5OuRDD7w8vNbLPJx38X3gI7Q07/JUz5i1zFVHaU/g1w+WkChM
h6doGQ2fmrPsqS/N9qXKezboZ0VOH85yH5dQYBYg68nlu7PWiQMwoFaEtsp/wIz2
3hfKXe0Co11t9tIYpE3cdKnxK/omnypsZKp/2wMsHXLysPHWU2TvRlyGp+kgMwXk
k5YeZ+MWqewmEXvIxysx0eHkUKIXIEfeC6cjIQhynYQjCUtIZr+G07C/3UP7uZMn
ydTs+qJVlg7YIvvlAzrhPFiLb+GkfRFdGqBuOzMQoRikv8a4BTruYSJFWm8CM64B
NensXyK4/DN8bywk+wnB2LDDareZMnC0yo9IINklLbujgC9nTu738LWZyqASJQKg
AEZVobPcEcfTmMAm8hUZ519BzRn8hVue36QoYcmT7CwNvnoa20CLc8QiF18DB6Mv
rnYffPSWP6P8RsHQs5v7MfOR/tB4dhCegSelA5UGAW32kGrUQVE0oapFdqwS1Vbt
w9p3DzzbnodCOk1kMxyD963Nj0f9wlehAu0QpeNqiDM3h9qa39IRPsw0sESPPHNH
E0FLiGLL0Z6Bbnty+2hIOZmrQdMcvJJ74E+8BDwss9wJ3e8WvSkYCpZbYkx5mrZ3
JYW8BK4tjHdv+7a/Jw4meWWEfjIkk+yu1+lCj/LAOQGYflg1U3dHB6QfBy/0WHga
OSyTKPnk09GVW3ldTWyNEkNT/AEkmpzpkXCroecQKg+fNxEebXuEoPLmFDTXEdKv
f/PHh79YwMsOKRgFpGAeTjyrJ2RKVrwyt3UjYxUOFXlt1x/GRUw1YENuQOVSP8De
y/f3OfLNFRFxBzds9/jr1M28Eip9A0JfBnDXfUB5yMVtc2b66QX7viCACnoJZgvL
S0KqC6ZQGrz4P+JgoyDKRXwrS2QwdQnQLEvN5M/RX+fsmOM+yx1I1Fz1+0HmrHsn
vM9sZKnNz45h5DUAiu+P/xE7oiiiFT5ZDtGRPzah4YyYJg3MCdD9bR3krZ3o7EY5
y5vlW3ltV/qC5ux3Gatf59ZULe13h27tQdsCkbVefuOc22hZ7gwy4RGPdPGxJjyu
a7Ex5DwTlGsWTnIuvm1OFbSnlPlPrgrV8QknxXSR+S1qgmdVT9wKI6+xigBJAnZF
5riO1XD9ZAhosEG5EjIKvE0cixEeAoRAI6cDwVEDtsjb1eTB1dVl/BPMODCcxe2o
AQBua8V8rKHtR8ui9Rx08bzD7G6ltN+bBljoPjsCjJtRPdNb7K7xuEwvcPMof2Sa
WAqNN8dIRfoM2zY8D3QS69JGlvBEU+HDx8x4qn34WUbKknMRg7FXt1taJU798of/
PdaBNGPFtTUC1Usx8I/4GA5+ImlmK0/uu7D/m3wTKOGbKqDbV/Bt9qeiMvBQs6vZ
gag5Uy4Uch/B4g4Z5rq+0y/UNrtox6YwWwbbAoTj0Yy9qsvrQMpJXs35kZppet94
/o2JPzKao+bFaNHidRS/EWmRyCG7GH4Hjs7ImF2xdF7rXbjpjBdrOr9nEpAxhmN8
Z8svLKSPqKHgw0yqsPic9dH5SuhLycxapPWR/8qB4VoIvayOJwXlUNEKmeb3RQ80
d72vMqTyikk/2e1HI2lqKgHF/1TJLXNnYmgNm9a+x+Ou9YcT6+kiLoP6CZcfg15R
hTSeHt9ksjYVHuVnJVMtwPVBhHQyr8zK7IYzuHLIPVEXpp1aDjRwrhu2Dz/YiH5r
FcgOMceSEhXhqktAI4y99b60+Qb6G2l7v1xtV0lVXAmMVY0cjoI1qLPJduebsv14
l4iPCmwlz2vm2Kjj2QPRTmjfF1/tif5+GDjPYD95MEQDGmSr2idLB9vvY7L7Jh2H
IBJ+v7vk3/HEO0g4zNiwRKQaDuAGPVLiGUkpuDC/RMXQqOz/vG2bJLX4C9qwjz5Z
fr1SRdaNIRkZLghU8qO06MduRJijMqY19TR7A5wjosnaE55Wiry2mf+eXVnO2V0y
PK/92XNaViSvgDQd8gI9x96xMFAy7+ThHJba56o8NrcxeYfwuM3GNMchJ4EMKm64
jf3p7kse2zekxxR5ti4fMI1Os3lORwKnuiFtBRKKmja47vMvrzIR/IEeaqQ4TXkn
NPMUWY6hz1AAsDpJhmUtQ7uga77XYE0yggJkXrX0Esd9IdBZ6DQnl6/4rLfKmhdR
dI8pN+8AW23qBiJuLqZAC1rSe3z4YTPFWg+xrwacQpnec4DndkhFkt51d0UiZdZG
gmidHvZBLQ3L4gQUTno8LlgENx4glRS7JM0HISdJpPTl+kcfWjRh5RWEbl0MxlTP
kKyCF/p3dgfUwiDJ52cqzXGFiuupFpwhiEm2jyQtKuHZWy5NG4d2oLycMtQUGs23
ulWrVmsAaK5Fsf0q9mXq0vbZHyZa34FQAJVze690Sq0vK471sGYPuXN485Tiojwh
xzuwdbMsukegcQcvSQnTWmIomozKWpGFL8qJTU9JbBs5K0r2/ZOy/I2phjzg8E3s
XSvP6QXD7cACQ3ibcqW8HjK0hHEWVbYdqtjfIVZQxhXRVDAEGrn9U7sFVckeRToV
SW1uSHeVWzsWVIkKX+55u/8zvYcTKgsegjJ8Mu0yQoHeHZWy5qCRVS3I1HP2x/H4
WKxpZnHI9hiew4O0MaJESl7YsSNmmBytwL4YSmSUtFhW4Qe7r10bosET0zsj9Ad7
XOwgjlSLvSe0FJ4Nregbxe5YFx9Urc0uGoPYXqu4jzBoi6vUSG+QebfnpBzZAMRw
va81ZdyrSAyKLMx4cHPkCQPp0T16J0TbpHtxNa63XM1gzLepHUY1zIopBTnTbCb2
2jqTHQBWbvigr8Sa/zKgOxN+7IVXqNi2BLuYZCf0UYyG9Ji0s5MzCxZ7fAOuPJ7I
BAfVsmJTi5kFIVOGWB3rc291jhI0HrJylxpMEQ9XSZ7eYVCCZHIbMyX17sKd77eA
yArToxrwLJ+Y8hrsW2TwroWe4UpZvB1JVxSPh6hrgrvTfgrXCp1/I1fm3/ydSXJT
EG72yKgfPUQa+QAcVJcJqKLlacka3LaXhEPzbHKk0rizeJ4ALnYRR4zfd5PhmX4g
rFJOsPHktgh8MFcRywmQ4rkUTsD9AwRJtwiHs+NJt1Mu1s09XHiyBs3ICYnRKb/Y
9XqIGp9IRNOIIyU75B1x5WfPUka6sCE7k9pUwMqqLa02SKIUeS2PwJICkvDjXkWY
Ko+iFtM97beiEMbEpVZUa7U/NOAJC/8RHvh1vQ+l8jQXxuu6gLXmeHzwU8Pp6l11
RG8uRcyVytf/qW2ryMtGkedD+uXS+ohRS+PgMiLdq9kRqRWqgHD+JZhp9G97xZhw
322vG44tJZm+JrF2T5PwnGEsCoXoWY9eaff/KrTqJDxacwpcQYWMB9smuqyi4utD
0AdrIcnsbZfJFRjsyPUOtfep+ySIxRhr48Wq9DkomQGxsW0diSFJ5fr9xt6UZkRd
4qStjFCeOhGoWIn2dTRHaf/+bMfHPN92te6He7bjApcOWtjO0plxmYa2C+YHfRlW
I+2tcR8L047gIz5eS2ARCJ9k/dZXXu4bfax07HL7D4GMNcBsJkkdX3UHmPqmTPQY
PqvVYEnEzkzIMfQP8dCOfxFbr++g0D0mNrUPAbLlxrUrpEDsx+bC1fo8cvTxzxdr
hvDixhZlW7Kj6H5W6urU6KmFFeWG/q7UhFY3tn3kxvcYrnZe+FFFxsS+Y6nh7Re8
htnuwsDo/CRwV2XfWg/MeTIfoOhpA578LJk1EUkWE1XzcmQkNOybDhGVrN4TAzCP
Yu8XVRNMEY/9fw6142OJkEGzrgW+l1R4ON3p0CFLZSVFJRstF4yB08lbLSIBNS2d
FxXBT1W/P6W4F/KpsNbrYf7a1ve0JzWt0eb0DzVVkbWRpwGJh+J8AqxnBczo7nF4
C1nBaaUQ2rr1k83+uKACUpq6EcEqjhg1uVHgDpsS1VDwqLO+NpMDrlm7vyVWUbQn
pc6w2EfLM/B9UTTe+xNhVZaVEl7HaORuCKoVOEKt4XXLnHDvl+8Ale4OSEFVCvvn
s2+nc2WACPx83CufmenAF19akY7hONeU1r2YpNP14EiDfi+etIf52b5PQ/r0pK82
keqntmHokdKbU8IUoAnscwmeb5RD7wtMJvpX/q2KGl4V9A1srY5+zO059Zg6rWTw
fVLj33lmthcM7mLMuTfrk2vzRtG79htiBC9eyIkaX+tcNIitZSlzi6FeWe/1Og/z
yBck76+q0U3zKXTv61mJmMroZo7ogkwddKlC4BT95B2KPxc3uhxr4DViXyJPLOcE
HVHlLia0OIWtLqeaQcMcuH54TnJg72noYLsCDNA4VN6IG+uXa75z1AtOfINzAAiR
uA2SODkR9sONEyQl169mW4aUom5NLLKkGmYqRn42u+hF0JbCfWWTigoKhO/gDStA
Nn67QbyQaVje/PXUQ3qvT1ZbLigK6OfAibAMGP39gfL9TnbQ0a+nCTirMbx8vJpQ
c/BmN8G2y7DBLIzfK29k2JOU/PiaVC1FVwRZLkmIudJOf5S71XrvLilFzzQi9fjp
Ps8Dkc9fuwUtalY1k6NNonGHTWkTlP/2F8bqW4WyT6+2FPyaP/EYRs8ujm2EYz7e
uCdpxwKKIEGuRLGPcyNh/lpzFX/Kwjpl5yurw4XYrsBx/DLfSvQDvcre8WZToNI2
lAkQE107a8D3kCm9RFsrxqmQPe4mituV5TQ7DMqh94rX+SClT0mNiEAxruJqLgrz
5O5dm7iLfczZva5tpEgZ59imH3Gu8CxjsPdB6pblBU/Xi37uuVqy+8gkI03lW7j4
d7C21FwZCX1zbvw1QvMSTfuV62g88H/wvs1JAt8SoHOWHQO99GDxQuGKxhRsFu15
CJCMbU6hztA3Ci8nrJShA/cjpihzWPN0tv0Q54dz13NuYOK4kyU0ybZ6tTSmSrXV
nje+/DQtegvyJ12Z7zxq02WnAsMdTO0TKqrehhN5FlPUrhBI79lVMgvMWxNay/Ht
PxtFTXeTBlo08ppqDUM/F+Fe17NXnR8RYffVKyb7Xq8PfT/TKtf2/DR8GPp4ZOB8
znIdyhnVLHrmkXpcbb0w6/NIn3nIUQKtSenGg7Z8xmUJAnYSJT9IYy+tURZyp8U1
JSsUhXyi+cU9K8aBrsHj7kXftTkeQgNSbRsXboM/cib5GOd7q07zd158Us6kV9LF
9X654QrSQsrZ1TmoIFPmzkFHqaLwh2WF68z+AS9VEev0EUmJbpU83L33EDCVpKAQ
8veaZwB4vp2HUryGW8sfPjTXKnRBd/QSZebtnS8U9unCfGbLLThhL+dHQwySOi74
vlgcFOm63fEDHfJA6OwluJRFYzpGHCu5rIsLTOnE2w0gPFLEEqfibHYfcppoc29z
cYenvHfD6LRk0xG0x1JqlV7lvNea4tjmD7wj7FfSy8/PoItTWwrvnUqijS3Q4tYg
f+nbdpwx/PUjeOl/RxUI/AzMBbzIq3WTQ8Gcwo6G/1CDxbt2US0PWGrGnkrOPwq9
iy4zZ+iIw/o5H5bNlTfGQ/Axlczc0oOiA180GF0aA7C2quRbkCqxHNKNmiTA/8+d
QqPVU0TXFCt3VAXbgkT52rPNFeY+UDO6netSH8yiSSfQ/wmAGLKwi/VKzTYNKj3T
DRp8e15sqrBpEmauncSVCV3LNraMhxQqXMR9eawjrAHcapHLu428vINtkGCMvuC0
dyQdPAUXIcJtJWDUA3qrKg0KoTMafbXGzDtxyo3vWimKoOPKN20n8DtiKTpMhndM
HhvrgpMmhaMO5ejFa0Q1MU58DgOp61SV6Aji76oVY9xZMhRLKx5shJDCY/4t/Vdl
25vddINWw+Ae4XDMsctom2rEuDpKihk9alR59Nq5M6aQtmp2dg9Cov440I+l+jYc
bo+Sry8oGSx0CSY6BJxKFCt+Q+QbrrBeRGinwhHzEH1MA/8L9WSidG6+pCviUM4F
ODjtfGSWAyiSRxZ/RlNWKk5261MpVXYTBm1m1vWkWU5puVZRqdbpSUogubw5Pp3U
hJWoL5fhjM0LSjCASd+1d8O5tdyqyHpiUtWE15kLWOtL6PvrKDKLrLjgW24GZtWS
//0ZurIp3YEH0JFp1sZL3PTdS6tM3c5YK9AYFigIvyEsbK+V7uWZKdhjfD2fQPjP
udY2FNlk+k+LvT5wUPDoYT21rDItPlXCpwWcwirz5R8Bw+PzDWmVOXpvKZ/3zW5D
NG6bjDPdGeElHXTzn5DOZicYxWYPmVi3dSFz4bQuKbcO+bBqtF0iptX6kviP9z2t
4SvZVoq1HwdVuOMNQDil6uTptx+6wcmwqi5b6V7M7Rc2ihdBJN6z57kfbTdeOaJO
0UnauGXgGXZuQGxXkQj8X0M+litmTyoLgY2rX6s75K56HkcyAFTRsq5am+5R/RjV
ICmf6JSVo7lO6rcc3EShAmLNZW6djIWXaFNL8MGrG7RLb6myuiqbwQsqlsfu7KG1
F3qW+GZuuJ7KH3B0uUvIDiV9rkBWn7gdvTl8sxyvP6gmdwYY11sG4XKW29FpOfUr
OHPzN+XzdRX5lIrCmBs6u+X5BcoLpnHHzglZuAaeiTFMUYDYZScJTB4XmjSUNJGs
7xqcQhA8DZ0NoKDzre57sbXnXfpBputXUMI64g9NVLeNRdDo8RCu/wm5+hzJlHil
4S+taojluSeHOSmhvtCDsKw6XrzE/My8YVYutVvWizFNz8ILgopWzAa6SlF8B/YX
gOBveiztU6dRW2BpeRl375ExomyF+Ov98mtdiJ73rKb6OUZDeUFN60/iIfHEhhg+
OSjAVKqQF/hF6Kn3RKUdNUX9RwYYjKZWS82jTHAKuYLdKHDfYoSJwrhMuJ10tthy
Wp5zRsKTPBgU34K8Vy3vMy0m86ojqk4b8hYqDTvUV/PoosggS41Fy8xWYCRFmm+H
x3aWwaBW4bBrxouAev/ZOoKSOnend5w/TO20NnKgBz0tGD/Qx/vhzUO9Qlmla+xT
gF28QE+Y6Javzdhw1avSuXCXq8lnTVjTRfK7qUZyocOLWTjvaBHZUV7I48Uv7ed8
CmjoKn6W2uiBO7FRMGWu3KTjBq5XFgwrcXLZQEtaXi9stKnX6cRz4phJHNWQb5e8
R8pJN/FmPbrlEsdmNOQpk3yJfLC8A/R5zKs+kDYJPijQfEAsqQVqY5SKHfIvwJSR
qEcpHu9TYL09FvA25xtit8HHAk5NcQE3Kn3SituAth1EN+2WoTphwrLOYAE1nfQS
NraLOPaLxyJ9N1U+9FDU2ZjbaRQBpv/Ha5sKFIPrMgrKaOZYbL1cxLG/EYG42Wnu
CxPLiZ1ad2VJ3y7kP6Zfx/0fIGmeKhUxef8PqXokNwFBpH5bdyVpG8Pcxz2xNCo/
0PEAfP5xhxycXU2LkSf7vlBkq+1DkK4RinLT2GIYbu5xejJW8/594V9rn529W3pE
e1O5KpbHasXf9TDZXU8BOZqwtaRJlxD0AplxzPKEArp6YbDNVPn/b44v91kgDx4+
grRS59FgjCokNbRTErunLsZ8W47HhUKeEgintTk+RL35/Lb9laQ10RlrLqhIYroh
2o/bXGDpMaMvYKTanmc58YBvRiTTUdEEmsJywcnMf+l++ceU7hVdVG9Z7zWPyPt6
BBWB1mVESnrrRniCpUxWHE8krJv/RQA8ruTrhBuzGwwoBn442/oi5CVKQRqDu/3P
v2MCh81mN5/2bFULx4djOzjJC8Y6AO94qOE0StOgqmRsJv6dC6Y5XY1tiZ3/5RP6
yG0NvLeoyNzqUlcnZhB+bSPl7kMOggn+ZfIolC88jfKPQZjAoroz/f2yWug+Jmzs
LFCZZAylKiHqRyE5uYLnnCQD8hlDj4c17/OJeCs1jnKJ/VtyejPK5ELZoaxtmvhw
QvgQhqtqrOtRfrULoNShdo2WrKoxlqXOUCyy29HfGcsQFc2DHzD+05vBlyNKRyH7
9H/rSwGOYbpJUKngVZ+Le8znhT6UKGggdO012XCoaSM8l7nmUHe/u8I2iyoSoViN
L838usVPNhUqfg1KHMigI7ZcLlIDh9qVuQ5KI5xxgO4kKnXnknm/ktoioNC+L1bQ
epoDBb/3V39JKwcPJD1hHJU1BwPY59te+MmDrSQt76TR6fFELw051thcaW7gxFVG
X2dW/S/yjOA0SWFwtIH6OB3a8pU2+4gdqEq/vBkP/3xIH2QlYRE9XSQ++CiosmEb
PmVl05bz5ApA6h3LUDrabghnJFKEszaY9uH9BSL4OdR1XAsYtG0MgSN4JQXC8hnj
0fIN+9zos3n5JQ7avKznWoTPsY12evCmW9R/zJbeEZaSIF1kBske/gU+Yc0b8gvU
20VUK0YJ+0gKmyZ9nm9Zy2zOp3ORCh69hs/Q+N6lSxd9iqqzYlEmtqppsJM1W4hP
EPH4wUFKk1jCHhb9KO647R1TBKCOTSuZptM5aexmeFxBEEQL3elsPiAGJgn2rJ6M
nx0YGhlaxKx1SrUCfcAci/WYV7jSwHYRZBsDnOQErfx4R6mYeGmPlHRlgPITEXCB
CYnP7xUEx7l+v+uzX3okZfOq/i7wWiEXJc6o8Wx4f5VEtO+j7SY3clqIcC5Kwp2s
gNlw70yWrxocndNYajldZ2Jt0cRHTkRFY9HJvjRdy/sck/Pzw+8JWihMuPFo2wuN
3zjHzPo2ix9roiJhjo6f24VGac/jsg8DklxjkkaadH4CQbE7zNZlQj38w5HY0Uia
eZk6s/3XIWaovZVMCywWbd0sqQbgIi38SyfpBGR6EWEhBeuyMTzYx+w+UAkRHcdv
PRP3ZSWujtQK+Ww8jPi+qljzsoTyQaM14WGZdzGn3EpkxeRswoEP7li+zRdaHbvy
tz14Jmw4tz5dU7rQBE49lCu/JiPKP3RLSR5bYclnDoZvTOeFOw9alMQoVIhtX222
zE+8/j3n1kR9ZEonifiFsrJn2W9qXnhYh6nRJwmOhl2+syBj40EeOt5cUBkVPGHH
zX2eqc9kpwx9PaTWtF3NZaGoKIa3MNgJmh/IzOIYhscev2MRCuVUr1oi99rcPhsJ
7dMGCAo/osHe/N7awbO9dtKkL7rVd50neSRbXZEtMCgXpivCqB34EEBQRZYeTpdN
aMg8bAvKKFkl4X0mWg31q6PV2bV8TlNx5cnwM9QEKFaCt5nScgR0drSkF5zwubKs
+AsfxVM9B73nCUo7f48KdPiiVNfaQpssCtXvfbTEQNOuNXAas0Dj6XdUuVwbOwWw
y0J1MYkpNAf1ixj1cftIb6HWP2DBMvlq7eCjYO7tu7tWNQ6pGQE6QBoBr6o5GHvK
XDwzOXQG/72bY7D6d0sk6f3zNK8LOPtbXFEZMoJ/2+iLudS1wH3o+3e1smplxUwY
fwJL+mmz25NeqdZTonG7wmCW8Kth3rQUACGn7/3NALaT084PY83bHCi4AFsafFTm
EgMC4lrV8xevPRrligUmaAVzmLm7v5/zmJabsjaxTnPK11GqCcRRGse9Gu7cZhCF
zvQsO+ZmTQagxMSMC6ORVw7BU8xvx6/GZd0JqYhTiTwlK4WfyzssMEiV+jSOFI3W
uwdfVoYtHtUpWb0lWVXVwGU78nSJZJKb7T9sW2S0jJ0kUBQK9Xq+R6thJBVMRZ3P
/Bjyh54LHs32dzSvagBW3nTtrfaniMYqJzVnvRsrSTYeKbgwNte9QN7rHIPBxAgz
8sFcIqxLHhMzhqitNQNlfX8DdCSaZYUMH9d9eUPjrafBCL6Zga6myPkcqUW393dc
zBIW/mC6hsxa+ZIZwzyP0hh+OAntlv+ZW/K/UjOcl9xd48WbLLUSKPTaVMlIn9jb
n5UY2yDn3HkxTMDpdWcGwJQLz+7vv3/8Ozi3zYekuX0DFu4aerrwf+RrRZYqEVB2
I20nbdhZIJcPGkWWGAK1t1hmvyhpyDpaXbv2pifIoeUi+NaI0Wd5FIY614Y80rp7
AJ5j2WQ99WjEvGC8SZPMKNQERULO+3oYCO4uOA3pXUeLvOpAn5IwGlBkL3ZYSBg6
mpus0XIAbtFwO+K0ttSvPkDwq04t2rJb6w+7Hnsi/MvkR0/BqQ8up1qc2pJ7nPaC
/QDHNcRUQIlGoVjzbd5uo6kVbfCOELhlXWKs2ryvoyVJag+hl/zz3MMWL/nqQNGH
gBmiMNH8OoxoRYOV5QpTV5qkrZMODzw8HbMO7wE3wzbjc8hEpZGRL8CTkESdzy17
EKC9UyJ5PNYsfRbQKVk63FUMW3ecnz3RNgSayOdSu1YD8NGp8Gk9PKd0usbrJYVH
qMuNvE2ShZ/qAkV7H0QuIhA1ifjUj3u8eMu0FhI38emw9UwdN/4Ep53cz3EtsL5P
OzG0q+wNZVCTXWeZ21SlqnHxzhidIiKSSDiuwc+JqKXBw97xBy4I5qj4F96k5Nu0
8XL+/6r3dHEAVFrDnbjnBX2mjIGtFsTdbdxwZeIWBFTyUE21rRa4JPAtITPv+4tp
xEXOHaBqbxoA3AlilqxX3yrubGSJwKa9RLKs+N+HBPGfuQhzjXna1bNJMmVdMpoD
Bv4XpPhIoZ3adqWqW09Az+RUCEPx0Jm9oo37oSVjkos+eXS1oHyUprtj2fll8I5D
XOcwq2vQqxNX8a+NKDAJmuqQwgULXnNuE+lZ4s7LziywH4uiQ5RwBrqrf22A35GT
AcSON/Lm61xExtv1Dg2PuWYq443c3xMmyWhIcQ5WSWDfg1JehGC8dQ39th0hjesp
wKjby8Kt6117xznow2CJdT/qUoRzOvHyO0V4frFEdNBQW2nJ/ls7quPkS7WnZ63E
WzjRniHxmcX4V5q2tYkCGnvG8K4bLjwIX6WVP3PaRPohmzxEI+0TzJSY54cnC5Yu
3TiBOmGyVC6JLLnwvvMJ16THubTmQ1HVu9EibyO+vzNQ2kmhIHRhhkpCeFnSV9fE
aUWlsxU2QEKKbba5zfTFHTZh+HD0g712dfCiR0P9W2Z259JVwpHB+aaB9Ug0OCnK
XPAaPCDymZJL6c5aBYgAPGRSt9VYb7jPasJ/6tg8j9vNtFbCi1o+yWfXgaA1p+5y
adxvmAbxCq01Eew/5F7pLWfrtkwkPWrT1+Wg63ISmzt7O2feTL9M2S1da3pHkrDV
6d/uMGYBBBTRwyoath8s6TJhBjubTwrPUl6+nx1h3ouawTD373jdq+/Cn5hOz6Sb
u8Sdi0+M3rjHuWb79ClJM37OMKIBs8hBKjqF3cQs54ZDm2uWLBuylhBj6zwICd5u
cj3Msv31ARI6083fkig0PcNGIV1xgmtGf5Nton9m590N8ig8B7rOa2HwmJn/ssMS
RYUPkwmXtYHlzsw+RPeya+G4Cm1Vph1D3j9MjJPDcGoFwDVStC2CoUngWauQcLB2
mK7/Tu91aWX5EGNrfHwGVKXHxvycqoMp9F0FFDmRa+yEhj/Mrjyxo6/ERWGX7oSE
uNox093swFi2SVGXX5HXS7jdcKz+d/hO0n5q8oOjYMyRZw+V6xSGqK/3ohtTx1au
wA++vseNkcPV25HRoEQHDj2/3lE2Uqw/6q56nSukKSzk5Ev6AcFqanZ4lZS8S1bb
XyBkPHjuJGNLpdA0ZdaerydRXfKxfYO/hXiVETYKZt3FoasTCenB4hEv701hJKuf
5C0TH4cPc5aPt7jf9GpiKUvVbZDq8bM6kiHFW9DASFPPeikWG7+KER6B72skFnw5
EPrV23gwhv4FWAsXdGZLq73gwg7o10EJNlK/EtuHmeMmH8hApJUqa8arhdmdhjc9
0yCwNguVKryxCyzBsMgElnDdGLZzIZPBauhdZjvfzkYSKTVjpYqtBd17GrS+wVZi
iltvusm6iT1OxZwO8WjVRI8PIcRBRgWnQ03PqhYQqD4vHRN7wHKSzZw4mQOb0CdI
m+rC+ctUFNYudWpREwVu7bflzSma8dXB3dLr+VxSJmveex0/WircKIV96nnXMTiX
f6MfXSWIMXX088pTkEkcDTOwJyYOCzRPvo9EKWgKyYZgYj1o4Q3/VE7GbG1gDNrI
563zT0PFpUlA9tdLltyaVh38ZIEsSgQSrylvMCyUROmt3xx3Ie6xjznl68CQ8QMS
J5JHvEHOFcmlqq7g0w18MnRnuK9EUmM6G5BiP3l/dk+vdYscFldDA1U4IJrpNSKo
1Pm5U9uzZqQ/7T3yLcBr2JC7lfjB4psbWs2UVBW87Aoz/j/7FsobRsMZHVpzheB6
HCtB3pstLUCGasyb/awAq48BqyOIBmo/mLLRoYZJwyr9yxmE+OhZ+Z1+PWMS/QQz
JVC1fhbMBbo0wNZj0nb/xrjGNOGNI4E7q7JWU9/9b0SYoih88n6FBbCO1Q1VVcGK
PHDPQZjFINkWSCqVFwEHoSrBGiWHCttss8Uk4AiexdWgc3ztlv/L8uhva4T1jSR0
rIsvd/E8tvcMbJ/kNsbgkhOJ+JReRWK1hBAHjTo+2EWhBr8hRe6QrKHBp/vxQANv
dOrHeA02NOL/EVQAp03hBpQvd80DmNpcQlCgp0pJrFIOcQ6Ag8yugDS5e0Tb6jLj
oTTGEabudRNBFVHLCDJeCo2iiNx835Y4wjktIG/LNp3pK8pW7tws7otjG4J1cSgu
hqcNKzcyfj5VCGh8mFFeq/73rQbrSV/rFmuASNh/eBONo2krH+x+YsYAI5oxpAAf
lCOM87fi/X/08D9pHNwnHZ5og/Gj63y0ZKRbQp1cwcQ/ma4MpcvOyrB57/8wij8R
YwiIb7WHOhg88N6Dt9X9ymrmTj0eOB+r4vavN6DTjsLRfVpd1QvDle/6yBpiJ1PO
xi+R0k2MxU07dXKykg7WCiCqH8/0OIiXxJNJLicQySWy7DcJr6W/g1V2KXs8vA44
3JJVyCDna7p8DtUy7dFgIVBfKYxAgDatbthEbk83AspBQE2s8jvj4GtxXEfj0PGq
NyNWTaq8wtTHMwQs5+zhLo7r4JKfzaTTxJpmHi3+IhOyqSkJ5m2rJ2Uw2COB1rEQ
Kp6QAEv7ADjOwxpyeE4S7EPh5ZCVHVwmixBqDe5uaK/OUR2+cO+LU/zAbtFaBcrM
91UOdPU85s08uNfwKUIeVpckMVFnY8oqupAO+HstuRGPiBoO4S7HGqtxc28N/HNK
10glBJ9RTDYKoC7xp7cUaefvmLkiN3EePEh/+IgnKIeraMwWHQRNU+VGHu42QUWh
o25EyNcFVEe3C4RRCKIl8Z43tfY/3eTyBo/wKIqAbyksLMJ20QXe9XR2IYhLdp8L
A32HB/n3g7MytdtwyS5AMku42rh8wGRr+tBvWpra3XfnxagpA91fmBR9Here0GkH
we8MXwovclaXI9dD+8lT4hSiBkL21182CR+acdZgM+rC6Hzjr5PXswFzKiJ8v5uD
pci9iEsT82pE+hXzeYbxdxXWAGdZsO6YVAp3X5JOs9EPozlRi57FN5MOmSZTm2X+
JWxqHtF/lvoX2EB3E+t+mFAfNL1EOdcfquAduXEMAiucfLWFnu0JkIdIinu7/l4i
ZUNganpcGMesjfJkqF6/o9URZLCR2KroCMiOuCGgDj0uvU/IRWNACk4jMOttz7Bm
4Zl7C+rElSgAOKDdJevVbMcf3Is3bZPnmAa7PDtSWTXxdPePP3OzVZiUb1rtfnPt
YBtwgxZfr0vcBihAaIipUSAdRMi+I9WZtJWjWJNUTAtW3iVSnLf4wAMAsa1O2Ukd
o3DJbHJpxTVKdwogh1hmXcyqMiO3KhU/N7OjQLQ/bs5tu+GrJgwISAISvv8681Zc
0t6Rw/P0SiR1rnEUAftGTHeqowkbkHHTzwNLCc8E+lMk2trUHk2p+ZxcxNDc+NpK
Vhy2GlBVGr0XzeteVG5vCVmX/TEzZrTBJfPID55PpcIHl+rfONoo1voJaPWnz1pa
EoAblANBGsd/JTVDXJpPgg5j3wvY9EIj4Y/hcfJXwNfa+KokRsu6jwPuNyGUzWTY
vyqLB4NW9Cvv9Ce4kb5rDkC3u+QZFvsAEy0dbguYXOq17Tr69G29cAXfHD+kuJ1J
/ymYm7zpFbPuzGuJ+ETkpmLAxhhXVeXtDRqOhFOmFEA1RtX0O8EfxYH/FqOcPtTI
uyhZnMf0eeb71XH4oRafioYm3B7tFYOHOKzq9cBZ9O2dJTp6FXa/qCz4L65/+WVk
dyAkbCWUMdTXc7TsPGW4ANOGvEoXklS8vYkCxnFv82fj/AHCsE3IS9vKNRrAu7iZ
fZamRNRUwi5ULwrhbIMWpIc5zLrjXPHBVTS3PZ6V27o1/7XBWbhsGkotkRku2GWE
GM7cRYIf2ama/cVSWKQdwQtRdwiu9yJWk2lxl7JBtRmnUjJDkQCSErUDuA8nKMsn
JNuiBNmJie0Dwfy/FFPZhEvwgaqCQ6Au06EgKBn/EA1RnCG0V+tauA932JhNoHZW
J7+2dfjFhGekwzG3BOAEn1/F7zmr6zGNi4gi+26gcyH7JRoxvdljnEYa8n7lReKN
ZsTKR+/isJ3TxBCUtEBjAS8pqYlTH5pbKM28ktPNQ4XeJZVpAF1R4cpfP9Xa3Jva
jiEf87n+3dQpXXieFYiv8u/B0iAxqIbf54wckFNzfF9YTA8/QbdAhMbvAbMxlRmb
GYhcB7k4uNlAfdRAkiAjg7uS1zcT3zlAxtzTVbaFRRtd8aSW3GKO24WegoDcuPb8
FB5OUrM0RKcZBNLTCoRoRBLY0DOyb9SrZzk5ZxvMuZxO2CneWo6gfb19pg00J2tT
Q82k/kVVKR2iV+yFaKrovvnd29B2AqoEMtvppYl08gxohsCQmV0zIf+hmySUHxn7
Gl7mHUtcnRHrl16J82GysVeDthOyRSB9OW1Rdgvr91cFN6fuNv9aTN4YOLpHn3yW
KWuJEQHmzruHuyv5c7Flif+d9Hae7m8FFPp6Yh43iNlmQ321QSN9O+gkVIpHQ284
jsVj6qxzIMy2Bz419ht7ttGBbI2F4OheNv1KZ0tDE4UwIvEk0ES7fGfFK1P+5E0N
DT/hxq8nI2DUjnWx1r9Ygx6+rrgoSN1no7Ra4/1KOFYM8rLdT6tyd0QF1ZzGLNE3
PN+BaLZxbrquPnZICSn2ry4LOWX4fiNNvsbpnS3kqW+1DJK9DdcumaQa4PBhvjMx
a8aniPuQXMHa00b7rloM8RS/Nf/hzzJbSvU1UQ4YwjWnv/Hh7Q/dWLFcxVhE+E5R
EcjbZTBPt3TTTJDKmKIcvG985YmtWt/TvsRhhLrsQxcz1Wpcb8gvaxgQvHUzQoX6
5QjQcWtbtqyzT9e5EZWLrq3QrJXC7p4wLbYVw5lP+G9rtX9Jv81rMvEsta7noULD
30X5KefyX8cnXqHKXOTMz6SSk30UH9bdoMJjkNwhSeE33jaJCYHyudGWbdhxOmbI
LX1lUWb2bbYAg8gbcROudJRjd2DPWZF/xoN7+9ydtegOQNfUlo9Kn9oIu3mGf3fp
RrZh4a2G9gx5M2D5oKg855rpBUi/1CI3B/eO3CH1XJqlY87a4PsQyi4YSgH1Qc6S
XNhvQCsZxUjZy/GVfL65SvZLABXq0JBwpOIUSPbRsVt8lMmyyrfkZ1Nx26lgGZtI
7QdTCtlVMrYF9h8ivWNjcyAqFU3M/1KbWPWYo2HoOD1NF2L6uy9vFrhp0C9KLXZs
lPUk1R4+xdm1YJW3gy2aXDskP83MGv+3d0tChQrc6Xvy1r9H0qscIb3ItZzm2/YW
zcBrapqq0xv+GmaBYeage17VRJ5JFmyHO2Al2HbshPSZ/OYeMSDVS0fOFF5S+tEN
hNI0zvehq/05yxc18ek1FyCUgnBCv0QTC8Kuax6835HAkg2yywiDzZt/8jxmmz1D
/5PcpsFNDE/jhG9Np0aZzc0N4XruNGDY4yMKVWnMNQNiQCBGfecgNHbpg70rL8Ie
Hmfb/+sx0/vcSmTeTOLL16ntHIQZEZcRaTRn0av65qJjSf1cVfKvbSQQxrE6oDYB
z5iF9J9B/OVbliu0rChHa3cXu8UNku86SUYuMy3Np4+KbuUUAxpRnEvaiiVb/DI7
uOnzdNN/9uwSmaP4FdQK7+fcRWaMS/JBthcf4jRt1edo2rU5+NXixd8IaJWx+kLl
Y4vpLlvNPL2JXxos7nr/RC8qV5bTubawB+eVw3UGZFh+43gdM5Pcmqr1gSQlYamK
B6WN8mQFPcgJIlojCVcHHXdqpyPkKmITI/7ng3w2edkxj86VYgefJTI4PCUKM60X
a9HZK2IS6kL6P76hContBrfWSsa88GYrGgODW94ufaxsLQQYnu7+RNa9lTGyS0+F
TqmrmRVCo+hFrGzgj0tvKA6TNwjLuPzvTAfW8jzcpoiABzNThVsTDVbDJA31o6GK
fxDaGeCYVbedeBHYAw9fasy6YtG+VZOGA+8pL+eBB6McNAweVTESqolOvLFyM2km
5VlR41B/y95az2wFIYLFEH+P+FRfcH7DXo616ePazMmBvPQnsz1+ShKs81byHLfj
64ma5hlBgYiENphz/Aya8c+oSJ6dUjvWe0qowkmKWEW8fP/MLU5+ePxWCpXAXN+l
BsLlMtKIQroRQnMJppmJPgzBmkmTYVow3bmD9XCLemMrjAZ7ka4lyDxP8fgU2RVP
47+A6eyBKCZoBKrO74ab5GuqF25tIa7RP7z/gjn4iwkbyyi7+NC5/nmFBVF0DLX5
SPRba3NAGS6FXHcN2Vg8jTyPL2kAK+w+8ArjDyixhoBGY16U3Vhag6bPeAtLXusy
Tfc+8VkXSZZtt6Do65K85wCOkJiB38OxBs+mT1a07JJ2SVYNYeQ2FYoGY3Gtk163
6o9ltUW4g7fnYVbG9y/aV8XJmT1XP+S5nlbGSllEBolKI0tV2MvUFfFcQVySIDO3
X5OIlLPRKugEVYGlvIVJPgtuwYFEjbqi/GW/FT9n3oUn2s2kzR7HlSB5rdq7gj1Q
Uwi185zuf5aMCzNjVWkaD0bIlHLvGwiPn5P7XnERf0qchKulqNfU31Vp38ixI1GI
n6iS0F8lZNW1lbYkj9EBi4Z01X8bLrdR+ajQlan6pB5O+Eg8GghBAjz7W+SNTj++
I01aQQiFPbirtdMfux/xbJ8IjGQaACYLfRLV6dGQ7KzzODsKabRtrbI9L5dkmsE5
woZu+cqsaB1+IsxLqfQ2UBYxzcX4twnx4JuacDZZ767BlXcI9jnYX4dX/2rD289p
R9XGpwtKwqUVOtITt3yRD4V9D0Begkk8qRI4bUH+i0FFQPjOietO6r9QLBtT3HNB
jCXv6DPT2isI7tJZZaqNvuSlQpDQBIH78LhVkXXK/J+9AJlj1BZCSg99LtO9LPC8
DCC1//P806Cos8sLiNk8bb/aadOdkNhwRV41XRuys8qWybXJtw+Z4ra1OfnRTA50
cAHFWBnMzNc991xTpzaeDwCZxs22feeUpYRkCyy3+ALRUpTroMU7DEWK0qDF9NKq
2ZEcAQ1GkDwZFA01EBlvjcJB4gD9abLz+vzI5tjNkSyieoeEfU5vVmeBHuk1tKZA
LZuzfOB11c9h8yjitytOwC4rCfC36YBbJ9brMz6DZT9x9kEVFEiBBnT5UciG9wDH
yc2y7/mzvPfHoVLu4Ac6I7zzhjbrXAVHK0yTwfc97vCZ4d+98GNbT77Iw0apoR2g
XDrT4kaEgSYpsGHZbmRJL3C5qN28VKdkfipx7o6dhccAYPhdp07ZSVZK+T4/d4a2
xr/jDEhAaxupkimDyj1pgrd+JDLnn8yQLENEBeLcM8Fg1gH58XVMgHBvWynBoJ5J
ifhHiHolK7gNLXl3WkXM0ajz4L6qHx/hS/xIOW9mTZdbIu9fI+4WNj9VjH3UzW3N
+D7JtWd/Fyq1QTF2gbbfFsKUtsFJ+3lIfX62lngkzLKjVLXxI5HYi7TCHqe9yNQ8
PoL64QSKYEoK30WY+hGRM2MhIy1G0OyUEgJuoL8gX4diuGph+hY8jbGXGyoxuS7g
6WynR6xNoZ03KjgfSkFTViwLS5CbUx7wKGiSJDluyhD9CfgsnRtXaWPNhpyXSzGy
nJb0fk4C54t5Xl4xKUHKYNoi/HF/8/BDjgBkb+L/xtGQs6+wnZot+DtSk90M3RZf
nPP6lCGdnhHcci37iRA3Uydb7q+A8g6S/z+2C+WYdrbN83XEPe4fejhePT8OfX6Q
MCYOTjBuIETrm1zVn4foUnpIoYzv5qOF/JIiRanpddgOWT09B4SnK2GiF9r57Meh
ASZn5S7LimuInbEy6r50nf998JNNhDColQpbeH+aWGO+XU1zk1bTVivuEPva7jqm
xDwWZZyPVfdqaDkY/VOdHeV5XQ8q9PCsT7tgNzdtrFxSv2rbSFIX7CQoeiU1tD4W
B+To06fXlQ1OTbqWBa8P7VGEV2IZcViu2CaPY4pmAwMPhz8/0i72skk3hvou+HGW
uE/27DX+7EUwQcRKYvHuagI3NgejSkRc0zhN7W18pV7w0LvhcFKx6d9anyNNQpa/
/iRgXgxbD+8WTzJFmdFH6zqSUJv8eTH28aEP5dyMhu5jLdXSlWyLkJrI9pDwmrwC
kPWsVL6q4PwIwWzJL20GNGe7FAFvoddxdjkRi9GdcX6vjsCTimSN+uShmLn8V1fC
tWydXTBvCioaqntBXU5CXvYzh8pazE4VEQWcDJJ6eEBvmZ6GiLZT9WAoqRVfPdrh
2BCcWPTbtmVFiLHBIdPrCCutZo/Ad0IlEXJGrjwoxvFEL0l0Lf/XoPkzQg8uFEYE
lzWQrG7+ehix5TpFrhzcnpBYVjZ6EcbKifnMTJk5vk9Ydh02r58CQyfrpQ8BwJVG
5RRtGnh5/M7sobInvmt9oSYBCWxTkeeM1UVoVihF8CslDA+T7VgapbKEwsGPoiGs
xFu1pAW7+lo09oz5zY2Uj7febMI7n+IKsqa+w/JBha0aL6Wq+xeJn4laFxUaG6S2
PV45QLrtLNaECT5k2llsivxy3Q37X/nwLfrwcQSSsu/2VJZXtywkg5Ripqmd4Mqv
BMz6pH3o8PuwRcNMkz3xKIUtWAOjx98fMoGNgB1wH8WpCqLWyhtPnYK9U6BLFHCM
ZSTnncayRhTfziG1lI69wiihbOCt7hi49LKrSkDPUweOiJ4MIsjX/AZj3bF8Mgz9
XLkkdAbni/tIFPWIa5ffGO8SAIkrtJdWzSo093HtH22eRgM10LsCoAgr1OJlSzaT
D2mv5R0Ed/zmRutkr4y9SIhyNdLomNudzKG2qROQmH00QpGttz5bXo9yVJDuJuhH
zzQl0NlC51+w9803BvC75ZD1l82uk1SGJqezCpdOV5eWHqIsUrWv+H6TiUymHmsH
75+dGm2/GjcOMzCdtKL5GI7VkrnyeZEqM7D9yFFmmTeR4ajAMOP7yxCKuh/NVfaH
cfHPCneXPEuOm3td4AwUJsmQBAGrZs6UgSulQrEye10N3/CqUfVUUn9T65Lkr7xq
NK5+O+1ZtMlAu5nU2HZrkVSYju8pCf18ljR9leaHD4Uh5TTJLztD6azR1VhCHKfZ
JC9/I7W1GQK44i7uDoa4+dpUMp1pGDrlngCytq0LXn2wB/wQpm6Lj6L01U7urS42
nqIOWWbEcpAt7S+MHjt4m8dctzN1EALUD294PlS98S2wYmKNwc1hkyl85cCRiqdh
VMZkWD2mcC9cBTYYsR1biT/zj/ITA9nuc4jIsOZZPZ/bgMlZXVZrg5MOP6GlxGvS
iQH0Q/W2vOpNklnjvlIlA9iN7WPxiUqWbwAPfnQUOIdSaGUjiu9JhmdIz7kyzxh9
GFDgp9wpDXKW0xZJqvm6Y/SgCeltd8VlhGGPdMno+kPIzcCXJGvOD9zz8xaaxh/L
Y4ovAtbEDKB4W7KlLK/vzlDRUal908VVryGpdx1QrCPXDmjZ3czXceQbTUyYJyUB
R9dFy/jDv2Xakf5LVZcWWh7a+21BH9gMOcsM2uvalNaVdLRWgeHotKAFmApvMSey
JNZqUGJ6neMrBMkjnYBSluAaj7NKbggafptydkTzh5cn6ootSoxfSFNT3FMYkMtF
xWBQ89tSLPPkjXL2zFO80l+Xvu+KWdJq9MSk5Wn0wX7RhYBclotR+k3FAC7SWyot
eXbwjvwxBwuPYmySFeEkLLpF+EaVIrCwFb0U3c2CxuiAxbixdiLjYbhSn/49wpnj
ehFsxbD60xlZ2qEH/GhLd9PSjqG6EJZAnLmD2KXZRhVrZRpO/g8OQm/yOMrITcfL
eLbhoT68UmauzFdsqxszLVXid4wVgPBwe0UT3KkaGHm4uS8pHhCRIHmlNwMrrubj
sEyOSP62lCNKMNsFfdAPHJPAqb1gKxP8LCQ+k16gSPOhj0A1vtGMZ7T0CyYJL9mv
yVGYdpE4nyx57m4OZa3sTOotKeJnzOYUns19ONN8SjvXMydQ7Ki0cJ7BTwX82MDw
sdRuTWqqIEBNTgei7N7IhCKoZMeOn3EbA9xFs7em2YWD1DkjFwc7gObgbcgPStWn
FHMyVGZbxIOc11w6OCxncc6BE4lh7BHSwhwsm5I/05UN7BUONYwS5YOFDEBOE6gI
gCxeO4dN1U7MNIk9fRbeTO2J3JB4U2TmXg54Dihk41KULCRUkVGTJwjNRdAMnXhy
xZ3iMb5mSd72TGGFASW2Eg7Gs2DCt0nwUC2YMuCkpRjNLwm90SdPjffATVLaYu3S
CBxZOS7LO5JWAUqYleN2cHQPUimLwzZ42vD/FPuTXMnkN8XvNdn8LJtKDuuKyGm5
cPgBQHYKKDEiOAVj/zGd+cqsk9WxQs47gzFBVt+VTNjU33TwO5Ge81G251iXGv6c
LcfHEshi6VFZl1eRuu9lq5NJIbL3ze5bEnuqU/W/rnhCfCCeTpHediNmVfezkQSG
DKtYso/AUSjmmHNCuaWNz98J6jM2hh+Y4QCrP++9FYcNSZ768GXeIfxRdWysZvs8
fhSa9Vulk0No09PgXp5jWTyoMQ5gBlvtSeU1ET0HPXqYq0yJqeq2UDvMjvQlv/ab
nxbskWm1kXZIIWp6V2Nc/+C85EhWKV1QJoM0nqjSvGlwdzwxQ38uZ9n7F/o+roFr
B50NQiKbZJK9N4rZkMVSzV0uGu8LniJB7XoVRD1G/GKVBj/UuvtqoNzsQLG9hCzX
7EdyJ0FCzsgTjh/4AwqrSDBCYHG1QrVEYqmHLzh+CLL/j49gWZbjtz/d69bdPSLL
aVYPOoIOw85ztbkd935FQ4jPWOTP/OzaX1xppyG878dyLo/RfAIsRILpPNc0u+li
NA24oOePET3JLtDPRjeYus7Knn1GJLe8S7NNDEUAcm7W4Cs+wTsd332IywBXKzS9
R2aFgwQAPsw7X4d/SsBxxZctO4xfUuFCGEHTmo/IkHM6VQUrxVj9eqv1poysB5vR
5Upy8d0Dr1UpU3k06rSc4liIJduW+45tjJPLkAbq+uNTwlRJ0i03tT+MNETz63RF
tEYUUR5cLXwWACcz4NOKDRHpCa6ijX5r8kbiyzMJITJkpG5VXsNQ1SP3eYL6VJiZ
IDxRWyaZCkSeYt/ETbM1+t0Lrec1yYKT0//gK8NmSI3i77SBHY/CM4ujRDop13Lo
sD6WNLUHp87ot4N96opxlDyIzrIOFfCD/vXTjuUuwJtwrfcXPSqP/HAUjOaimoQK
qc53pRpUOoPWAdENqr9Sde97y4KLnnE5Bw5vBDYCHdUIyuFhQZyzETUNw9H23mTN
pTjQazkTLaxrkrHY5c2hsx8M//a1B/5hJSny45mCoQ9QesaytHLkFTmi8ivxeO6R
DsYjAFw2+VV+Wf70q+q3GCn7WsqHMKXwaJ6mD8R/ffqo5Qo+KaMSpBGJF888c5AX
cOtCPzDBibBc/KGY3gDDUPX/hs0SEqULEJnfBB3xYjR3/abMBCMQuYrBuIllWL7Y
fop34EAKZN4I01Rvc27BSCCh5nMSHWXFAcmQzVKlSfpIfO/83rs9jWt4k0UH7AIn
nH5HybKlpCpA4i5j+NXqqJYWhXa6cF8V/eTIbIeqgpVbZtcCyongDpH+lfyrfIh6
tw1S10azR9EZP4flWgzr0amxBuRmnGfZsJNB3yuyNuQ0K8CKyiLI+Dt9I7FkGFgc
ZBd4gAcvBRMNSdKYSzSG4AktQQI3NzVTIdAyQbZ0ly3qR8Ppy8ztfmSFzt7o1876
9f1LX4e3jrWZcyD95zofrE9Tj14JBJOKGQCZrx6eWUkWorjWbpZrFhuw9lkLnzEW
YWjvjTJ7mvBhLU5uR0ELyAnTF2z+Zd31/90uvxwcyWigCB1b0GR5plef1STUFEi4
wxFg/5FSoe6tx6GI+PexWckg2H/gOjDltuEBi5PuaB0qlJwmPKoyY8KLlU46qDra
CoawDyfnR9v/TW8mWNEtNcpwmbUywPqa1EpDIYfP/srooheCAOqOPsvEw75vWMvZ
vS3DqFnpLKMkMUpYAIht8dp+xZkCME4uamdYZUqX2RGtPa3ufyutnSfhim3OFCWw
w9vevFesduwFyEo4EViB0cOeZwAs7urhKgt6GHRZlvUGL8TYUpZq0c1arVJPDZ4+
ERfHU575cXzhDDXc87HrsY2R1AyAGmVWue6tRlcT5yikWu6J2bw9K6moPnLcoJIp
9pEf1WkTLm9xPiWaVNPCdcOJdlQVFXWcK50ZCzHsMN/N1QVKT6SW5zqCkSSI2FiN
QteoRdK7OVVUHV4qW2OYErU3whI6hxpTKvCawt2Y/c0bLyomI2F5aiKzVXl4OQ9E
8aNAETQ3Ls+6msdAQePy7CzpESFA4GEWNa/Mblp2RYW4iC3Oh/NeZJIhAhcx2MBI
kvdCRUBdkFEEjuhZo18kpQ22PMoUzY34COtoOPpUXprrac1pI0hvDzpi/w40sJlS
35Dg2Rbdh1kE4T6/5pj7dWrdQ3JtsedjetfRu+nT4zbNGypraE0kz6xcyBMTw9M+
Wbh0bw0q7HIeTIFy+92XlsxRo4jMo8DfYQ4qWKE87C3v1aa5SRL9vePUYhE9nEVW
WvzTrFvf4TdLq5EfBG3MOgwjOdUPPbSUTzt/natqXNuFtFiC2RkRKn6Dq+FvAav7
Q3DpC0Lq0/QeWJfPSBz9detVuajdVMJTASRPLXnLlZqpvO/vBVgJ5l4GCRltfywG
YEHc222W163+2p6Geree37wDd3DyYW44HzDuSVVj3Al0qSkCaYu9WZB1+bOfGfb/
yXzk2ljhwBSyJjBjsMF7ftt8zl3HJztwiKfgrwYqXblwZnO5nPAKmLh39qwu32xb
wcLxKfwwP9V7tdgSZ1h/r+jquFKMmYeI2BXML5tg0psksYCEJkpjJ9EE5NkQaFOc
ryyas4zBS8rlKwWJzkmxKTcGL3zjkewIzr626nOnAPVlZA1ARE1RW3uUznC3NAW6
D1B/JFz6YWgiOyUtc6S/f53LRrKSihHyJYkybvP/BRNENUFutwdLBpexn+n6MzHZ
vdtaO6FXlIIRpZf+IwDtFRY461uOj7ixI4v33pVAVGUMgKs/L4PtkHUnk8f115t0
TZPPVPKw7Lp2OfzHfCN984baDkJvPWjIB4xw4MsLwA75c2cYLtuTnOFUaqqJDFCp
U5Iu/JEq4SZJa2sPpOWPUiK1wZHdF9br/7aZCKIe7z1Z8JcE/mjLue8ky1hEAUvN
eMrFmG5t3Nq1Ni3etY+r7TPLi+7ZjGRtdv00iHo0qL38qR33QqT3RB55GmKz82Xz
8GYcII43sLY8B62v9Ty+HL2fXwi1AYNWJp1OdVe2J+RrpKFofrCgApw8Tg2+0Fyq
SeD5mPDZAPqeUxYyHN0dhs+oeUjWgygPqyTzNl0MnsrnNZUR3ad3AN+A9L16Lsgn
+9s0HqVto9Xw+b0+efv+pjx+o8FfPF5qLD8dcknvAU2PaLe3LpU9Jmwu2kqx0UbL
7UqoJV5oRn3OO8j23xYeE2AKa8k6iEBR0RHSz+dgNA6Nc2LfwEOX8UNcbrULfhmQ
R7/2YtF03jEjwN0HtkOQ1QtDVPrILUsFwYNdIWHM0VTbzrqoqeHFTQ0EdkJiBda7
lqRw64XSLXX9mNSUPKks4xk1YGRjs8vcOjicfAmWZVMGoiBdvQtetPqOCeEy220l
/DdL9Gq506h7+Er5KG3jwe8sUe/+Yvrdbbm9d+oSaqrRHyoKpLsNL0ME5FGEPvBW
NWihJVRB4v5BkH0CJ5g13129LUL4J5r1Tir6cUcZvqnO44rH7BTY1AfGSHufx+rj
2BRTIZ7IVDARADn+JpZn8lsL5xqwxGGL4+8XzfbUwC4W1wYIT/30cAPvQIA/W702
RCJzWzsrUwyPSaLcrsvesnx0wM+Zyvg7xY/WMMYwT1iqtfk+JaLpUNrCofp646K4
3eSpWPlHC247g1A/NllmVfBMjxVBeoilbJRL8j/b9Czb042rau2ehZQ1aZNU652o
h4KMtrMJ7Wj66YrdwimI20Hcs8EqWbGY4mv3O/AlTQZBdv95fYctBxmkiQ3iBTSl
GLpCdR4VX+dJ7NU9sSaul2HP4+gjipD1yeCFcVgTxG2vYwFSQOWhYIVp+APK7jLx
tuvwkgmKWW1JniX4EIU4p6vWED62zHKakl84w/a1DEgUbQzOEc0pNqrE2wGRZgOO
JoP3/Hjb/1vZbHhB6WFli1U3IYKqwOG4uB+eAOiCXrG8OR60MwNAZ3s0ObyuJGgT
ffcbzVNjRRrjFzSHxHqgMahKmAScXNeAI1hUhVl30C8RIOZKHMiXqoSpUp3ovRRC
p6gWQMq34BirSyjZZ6gf1xmKjtL8ebMJR1IfmMAw1uefMuuZce09LcGpxtAL1cyg
kT7q8HLkkxbjCmNqsDv4Gwg3Kw5D309CPzy9yDVik33fvc9MrR3n857wC1z1P/XC
pmBrHhnMPEw/qtdDAHRAt+ir0uKNDvHOX6kRpRMsLpfrSr5NPwXuuyX1uxcHk9Y9
9zXIzYgf6PJrs/T1WqkUGoSzZQQgKZHN/Z4dLgGhofKTwCaNqGXx001AzHTQj0kC
4avMlRaWtAbnKb6b8IQqsxNjEWsYnGWwDqI/QrrDY4JVx88Akc/1aESUY8ATh6OU
GWRteVYz7lS/l8aRw7nD8qFwI4UEMAt5Zsflr4w279sW6LJfuCgs/mqZaCnsoxhP
vkc9216tMohmpAjyNbEvDQ6mOVjm2u8whbca0aH1Dm18yl9lGKYXSsm5UpvO6KXx
ai5dEL0l0j6RWyRAp1BNFvkLEsMpnedfuh+gIrrgA4yCiUSWmteEX5w+7GHzSHY3
A604qPBh5nfX6CZ4ZqR8cKIgdljrf+Eci00C3q7X+s9+dLhseGRRYxu0ckebFCkg
0ge+32TCAHD38YlVgRe/GMd9Uaw2pH2DEcXiSU1AFpS9jAgQRwYJ7vkXVZdcp7ku
L76BY/MpER7mP+7eXTGq0EX3ngt684pYW2+8c1jwwWRveY9WAffuSaQ0rkRoHZyO
2oRy+JmgKG+Nut4t6kLMQT46Z67fIPbyMvu3pz4y4KxOmN1kofuQqeqK93B7Z168
sLl1VTjHJ2J9Dl7Ks8CyUN7xQ5MAe1IZ6pp7cxJZ3ElpOa7bIU1EJXwqsz5frmMS
XlQKapn5iOIdERpZqiB+VMS0YBUuArQwdvTAxpqafb/UEfIIVz40H8+e8FGO6U8n
pvH5a/XquLmNUpRgOu5h6lLij+UxkqGuG3R3yWk6BPxUGfTTvgYHfaGa6y5Q5/Tq
ijO0O//qLahkks9FQF0dcqPboO8XhJl2KgRx4Y4YNLyqyffHPodetPeUKp3kc3vj
qqN2dJnfusHCh7odJCAVVUZSA0zEm2Gv1MyNIfzKW2WgVubmCJa+buFf9aL2Pa4V
rTtCxewPtys8XQ38M2OXJpEQMm/pdqa0WvRfaRaZGuF/7ukQIfrFZJpdr29d8RfS
nIy1gmOP4NNaXME89ZswAnS++DzJ6BDdsG16pnIdc8gzKqo7nwvfIkAY4GDXM596
ez8qnAOSPg+bF1LEgdzeea1ADzUMQbDz6C4oPPxmQdM0i7aJ3ilV+iVjxbQ+sFL8
JkNbhZRYAUQMeOTBCrUHKzmOJA5AMNX9mu1MDFl82CvqOMP5QMJKjLHSCJQ5HPis
HJHOFY9Y6+4JFfWEdsqx4X3NqGH3TU5CEPyqL33/xaD4pBrmI4KATRwA8kkiaJ4/
4y28OFUDVZv3ynCVLTrv60XXL17dllIhEiaMjQZQ6TRTkyxm5qKkNsx6mOxyz8vE
bwOQW1sHK7r3EaUzv8J4sVvw78kxVRvOI+D4M68FN+EN8cgviZogiCpSU43BVWzJ
WSu0DKFM5xd1Z4hV0Uu9B4vt72NIZwaWFPrCRmPQOmdbLNjUX4+B5wib5wnNXw6p
7tAaDHG8X+ILDjkOSGlILP/5czz9PnlBPJJbxs1509GF4Hlf7CgfynoArvgWqyAf
vwHAmj+PbDxYDz2FOApDxtUr4ec2DREbqBCZ/DuyXhu/VxFgHxgOQk4HcgMf1oVf
vXQwOoXCJKURW/oACnYjdsPdtXMPBBBmJAXAQUGp812avcC0/8hU+xNAHhSEIMGs
WhyLXvrxZPkvtc4EaiYQ+roBUO/bHRAc9o5z+qetnxVLI2rPRzNcQyrMPIOGUJRn
qRSbI3BRG845CGRPDhmhgEypFMS0WW6DBK4SjP+cJVCY+8PLFMGMCMQ+5tlKoxAY
AOH0+W+ZslaNfW8A2TWMfWz8H3k34HKkysYa9XhbPLdfoLkxxsO61cUmFwoNdO4p
AkZiWQVVve4233a/xNKAUsm+fmpxHms4DZdnqpdZx3iD/smmCjZpSXlxtcaF1AVE
O/6DAYGPajdNhyOWigdw7bkktSafYBa+04UdxRHveHR3N3kDWcEVPRKrkEcnys/q
so7fF5+XiEOlfHTW+UAbNiKjJaP83HyakLUjVO/MiVaWepfJQkfjcWPLf6ZbGe1G
DRy1tXryqqAUJuep1RX7ewFBceFSmoGM8OU5EfoSPEAqq+HK4lvCnM6K4ohmumGc
FSr1hVCvxC8w0kB/VdfKXbzi5hmxRSQz9FqVAbSZ+PAm6+W+1aww6F8K0oC4jKFQ
cBepJ1TNApk9uAAdt/oGTWgsJWwmYYNAjQwrh49t+tZF7aeAnsFGmwtmQzP+fpFq
vXGl6r8sQqpnGoD6M+BNPA+qQUYKDGrf/akmm8DaqbMoXvyLlFHHUDjCq3JoQGmD
CetvqoJgzqxYtdfa8qAQHtw+oOz9aSGeoShTExL/iRTIXaImKz0/bSROQ7QeQCh1
VPcOI3N5cIBUDSfOwPx8rlERa8+Spt7zcpxEY0EDgWC4SkUf0h+89cPt5A8mX1lb
ZKLyI87avBRIMsxwa9EaIfBZNtBTrHXQMrNMWkHkvHcDGbU8ocAp94YBGYhVYJyY
M3mjkjdMcU8lQAXhumaozxbuBgMgWC9OWso9Nxn/mJCYz/So8UbvZIYt5oVchWaQ
5lIeTZo4pyMiNRZJEFiQsUp4+yvNhkIi6UfIrEAOhrlv4B+IKRC1rHDbnj7GNUpw
L4KfCbT25rA7eTXVCSk9X6s6lCZSDnEAPb/NoOX4mJ35LMVGtWxtCfmOvR/WgW45
Tv6CN2/NEnQ3oF8jEC1Dx1eE0UMfUBXOSC2ASUFBpPM62+NyOntlmNP7jRVO/+ql
/U9VKeuD4UfElZ/LODKjB9MKue8E7p6YRg2/m56/hOfZlq0mIrjLYWNax+IJhQkl
XvsZQLSu3T62j6AzOgh7TeAXtfA2z0dEONfVbjEy4AqvLoqt3in4JMsKvD+2Lu5Z
YbyvD/ZakCTrelKjyDumM0yoaRt8oqm0jPJ6xi07i/PHdQV1/pJq4YMYikEF8vEx
c4+AkX+Ei79oPyWj4F2PXY+jT90C+qcQVbRGuEHLIiMYn/pCfDXxntjgXzH4ysAN
ZMD3uYEzAoC+CGrrSLRqxmGSvYaJ3K00Mzza5frkv5p6LJohQBUXItyz9WqO9PDV
6ETKxv/mz8jBPCn46sX3vj1EIpi9MMTF47DetqWWvaQDUfnXa5uvQvzGxvbxeKbJ
yKK5ee2iFpbeVK2KoQoFGR2avvVx5O23pSgxB6Ztxay+lXNtTFu2IKRmu9ex/bS2
IYegeVjHz/FZy/QZzpAJ0A9W8lZvJf1KVmPMs4zzl3Axuea4+Avc07nrH1aIU1TB
PYLE+QgaKHxO/HpJJwhfo+IOW3wCra/MFt+shiBpXToa8b8hDJydbbZMOxitWexL
/wfyQu7x7d3IUavXporm38GLfkc4T89rjs/vD+KN4lE6mmOmkGZxRY0O1x1xDkPy
afMhQGGVRai+pErp++IgKOV1hsiMzquoHGV1f/VoExMW8D/HbV0NmR6te6tEBOlX
bP4wviyyQHihz+MNCDEnWyv+kEjrDLko7nz2j7eKC7h3zyFo2rDP7x+Hn9BQ1g7S
OdB2ijd2wZei/yhkIw24JkzQZEdOS0e+W0gL7+lg5t+f4sCt8TrCmDfyyKWu6jfS
7jMsnpKUwE24DLbRmwkv0/o/QCe6Ucqw0ayMrQ4dFdT/cLC0zb3jFQgj4wN7GWH6
yjz3bjNcTI2Oy16LqogImKuBBz9gFzB5YU53t3GVOLuC4/9Sl1g8uyvl2xQbCwYF
3cTUBI+NjG/kjLiZ4f8kjwvFKWZgADsxtn3cmWbRJLSf+lniMhrWqJFRXkJrH4ac
THIGiamV2h4LvcSO4ix5yTQG1mnBT2L+kHC42M/S7r5QCgkn3fjpPT6SGZP4PGYZ
1kHmmXuiHLKETW6iVNoOtYaaePNdDq2782OQl4zE4E/OWodSL9+0HTbUt8BDQkG4
q9X0nrBkbdREJLecQqv9QgaQK37D/kl4etA8RN2UsqkKQATzKFKhq4Rcvi1/p4kU
fasPHR2BvH3+zuATgmWmHh14G1MMwlPvSuZ9vr3/SXhIpo646oJznYQ6PdlvXQL4
RKlG/5dISosJPTeKzOwKupLijBsr9wRk72pF91Pj8KLlHeEM8OLEn1TTvPcb9q4s
iJhvvPATGGKEDL4f1B9NzpJtUaeimgvmIUep74yVW0wb+Lh0BvYz2wHKlwVO9Rh6
SCh/8c5fW0/badk3R4GIJKMLputjrVOLBBejf1GFVpYbyZdD2EwQ+woUZ4HQxZ6V
NK9Oc8Wy1+PsEb0tNZcfkCIB3L9mzpFC6DFZfuTldC5ziwnQGhD9z5COJ0C6mSN3
KYjh6WWEKy+ZXHDGMw6x80Uzf6fO9nUnnLlRkWx/jtXmeIVmHwPdrN3I0WpTnd9a
icqopyiBOhNXFXgWWAPdAFfoe539menPMUXN1NJAZ4Xgy8pvp/4nV4I6Jj5lG0Mi
oXE5rgOPhIB+4uOQOTQZxCUN+6hxm03NY7XhbXMxGECSjPY/H+ctb/SoQC/YHPfE
93LY6NMfn8TQHaM0bmSsaTGzhjRDTJClzQsuHNdiecs6BkAC9BqyQF3H1TiPo5JQ
v7Wnpaxl4r21bGKfbO0YI84V7k+StG1xZtaOM+SUzTBysxtBtGcztihg7OWw1ftK
Spim5iTZjxUrgwQ6LO387GOIC7AkIbkw1Fotm+YItXz+zEhfq02IxlTCEJwWxHfM
gwEeGpjBfo2J7V59Hy5m9EihDuVm3xj9dqYAjU1ZaGbkPhJF1tIgZZdIHKWn25Nz
EGmd2RcYz+A8tRKClinJQcphYeff9tNs+5g4Yh9bS9Jp3e22Y2Grna5yI0LBuOov
FhMc5E9+0Z+9LZBnJuznsUlHrBMo8cQNEHd+isL4eJaoT6aUTri1rL2J3d68v+a6
h9PpyjPqO3E+yhYL18acv6dYAsO4UI2QEzwn9mJX8EPBERI6kR5Py62R6qaOvX0p
AMvuI8Aa0YSnviNM/CXTZpl/Wleu07vjBkGcISeI7hu0Ofy8xyvzFEpfbk7PytqM
VT6gDfRyK8WCmVoeC9/b9LBTgfgcYl8sDUE6AtJbIEcxaqjZKuxwN717wf+EZdFG
pV9h30cA+0diXlZQ9tlc+x3Cn2TgmsVsRlFcKCbKOh3LtpwcF2RM7P0zj1Y1BhTM
/fVDNbHbelUD5W4g167zUF61XfoVkgK7NbAUPYfM9+qXs7/uMo2TRVP1YM7pI9uG
rh9BEpChwI7I98IQ/ZfzJwS8mLbUDgaYwCfjsAD8g4ASOlo2w1yuYy+px1TQMIiq
Er8QVn9sd//Pa5xUjfkeTm3TfaMABeahOJHCGZVqepxxgvj+RqqgK6AQ2svYUxnT
S1eENTynTSedPlA2196es6A/XqkHmTgQHxn4xTjw2oOVmBVZiHWlnOv2T331u9gd
MEj1/S7bfaoZ7xAqnDYVMGzsYHY5CoVkVdcukHo0EmxuWWSZjIApE8U7Xj930FAw
PYF1Zweh/PWGZuUKhe51S4hkCBQNy9PKCxy7NZ55WTFHhXM54xuNjUWgYzqzein6
ojSFnS/dZOP1ADlhJr2t4sjzI2byxER03CiYtATEAHadTpG9RNHuKIKGqnYHD+Cd
6fDUKIFOqofu0i6oTlQSrxTsuDgjeTcqNtU4wQ19qpOwGH8606flVdQgF1eGZubW
LQ1l4f7URJK5atu2hBdE283e0V0brtKIrNN2xLVUTnKXBOA6OqupE9dO65riNivy
Tw+053bww3XifADIjKECMJy39+BBzF3wl8cwC+2EfI+97yaPFJ014vdiRL5M5nil
+IwdgJy5KWg2ZrmwIh+NuzSHo2OXuo4khUd8iHT0jl5fLomkM/yFxo/gptdi9yP3
uPaKU4cfrJGHn5d+gio28rhy/fwrrmO7DK9UNfYl3BXTZP2zPeqjtd89xszs5L3h
4d+Pj5n6gdrru8SnJ7TsuPlCXAsVqHq9SuHpnllxS2Z72XsKxoZMPZGhWp/x4VaU
9NN5mptSwKc+b9+Vta5SSWUV7hIBSwDuWGKHHrouXGyvhOi3zaR32/Q8Bu3YpYkc
4Gzh+Yiyg4lidGkYesPRzszlzZ1J65XyQnn0VLL+Gs8Q0fyk7DnqR/BL/gvlMN9U
8JT34BzMemULTQ4KUBJYW1FTfW48oDF9LoMsB7fBplvqnZU0dR4m1GeDL9kawhZ3
heeyDCWWrB5mwxvSz/cWDq8mIST2nF4toE1bh82ML4iycIvcGjM1V6nBitLMxbjZ
CXpsvM9Z2r9cWUknN+vjVELihB6wo/HRmTjwxgbHM6A3ZLhC0xAtXcllrn3zmcC0
o/yO271qQK+dMGHqOH2YpejMdztqDyD8t2gLT/UHekCz7ZwU0H8UleST7lLi4Jx8
LVvWGtPTHiEmKAGUwZQK6ZrE1GIwqPytbLSy/tux8RQ38/H+2P/0nxFzC9Fjwlt+
FbnBYMe9xN7J4QYJ5HQIAd4pAye8YvWtBB0xxeOed/s8XjYotu9zv1+C6nDoyodI
oPkWE1KrBlTFSpCgC7ZWwNEEf7pWLYBjt5djVeNYgY+HidiNCYKWuEq/YL854Gim
7kBaMMNnW1IjJYrAdjjXyrhSBx2XLpQuZWoe9jWIuqdoSICXlToIMNSWcP9Jfu/5
NIbXcmqm2pxlR7YXPXcVUfrKqQqb62QhEkGiJlAbSfYSYqf9hBvesbHp782ZXOLT
/gg/EBi5XrlR2MUZzL0pyrH2wMbR9YpvH0hPTkv55m7EDjraMl/LPEF2AIgF2z/v
eep2/RpJPD6tMMdTKcyk9GDwiQhzlP8YVr9q1r6sv4eX8Q2nH71q5b2A/BYGb0AM
S8MWerrlqxqBML3DNzuDorudL3FV9nJbpagrNUHiMRYCec1M1Ltw7t9PipJJm7Wm
wcUyT1tjDvCep+UbkCbAf/OISSu5EPV+BuDjTIJsm63zNfS8J7Y/12KtAgm1H2VY
96GuD3I3Zaf9jy2yYgCvaoiMdrGE46ku6PlvN3LMmUEVEhtPoNeXcrpviHIXkbRd
56xYWC7Uw38+vufbTpo9OMdsc7yulhrKQJPdVs1XzI7YeEpt3FIjMP6Ji9qojdgT
PBBB03N0LQ7NClFeMkGdAHMucoQu0pTemsJQc7NK+upapE4bMDBj5b/aYGAJRiat
DXtJz1TMLZiDR7sFreGc/VICzTG9wChK6dPaNeC9xtRwLlySMhgUXLmOpbVtzkgz
8riOHLN1CQTePkHcEGwNnvOyANfOf2+rMr3HSsLqET14RqOjw7Xsr/AOjEyPTd9b
PQovPnxarJ3dT/uBwUksAhP7ES1fdWx6aKNqUxzhtSF7SyUUS+IF+ZBN3gv+S+hw
zsAm+0IYKLHOMiOHl2oS9lk5IFviCevAxdVSaH8Qgfk9o/sXZOkuiuXkkJuJVbqo
QDZpGWxxcbIbHNsdxhiNfrdCBdOs4L6CW6PgXc79KMgiHwraQx91tsOE4B6lUcLt
irPOXquIJnyF6m/6TD5Zisc+UdX4xMvdZ8S/bLGh1jd7sfqvZiutC8YHL5Hi8f+d
lWknYgmu2nbs6IsbolJyXM0NcTle6JbIlQMA3ROwFZJYVo9ai59dTWv6LpAa6LKh
qsoXZpK+2B/QENeA57rnNZQkOOz/Kg9CoHZhORnvX3JpEHyp8v31oleDiRX35kmN
kkOfQszltfW5k9MdMFg4xObo/05nAf8rtivw5XMteHG7/oqFwe01OPHwvuqVu2s1
DBGbQe6WmjpGQj0hhjyYPt1L+5nri9Db84xmPid7bEqAtGb5La0Rri6/jmLXCBgU
nFCgWbNe+UGvtzD0VYEejj7RSaXV14QH3d6MOHvgFxGDSU9n/M9Vq/7EirxE5hT5
GrDuVs+2ltAlOw0ysPgZ8p/BaWVvMOngpTUW1xQrP4OnM94YrtGiGRPUwy64wZuv
94dggeuGqba8jQmJmPVscA7c+0CUKplY7CbaRS8ZMAQVQ4uSTjFoxlYIkN3EPwm0
7koya+GgrXTyB4QX5nx5thD5Wy5287Fhc5YhyaBseZyiwGJWUQkqljASyXg3y0JS
a3X+v/h4QvGH5O8yVOqKpRXFnrjFFUqNtzZQHaB2ttjPp47NZEn20h0UevPhtKup
tAhNZkd+413y6SzgQDpCP2x1lWNg1YexY+ZNiA2MgIimRMrLH85PMO84vWCfEwpD
6both/eRkR0cavpU8/Zi1n13QVrdGsSjtPGAP12pORQ7nkwM9ew4lhyDbYwTo+a0
J2MSrJoMd4FJwZyznvKPZsVO+/V8R4AEEICQrSh+fH5NaYF/pQRvPyKezX1dn/PD
TEkNotlfEtgX7T7/y2W/REwakg/FuLeSM22k60DXnw4L6zCGNV+VVacWhyWq4Ubk
FAIsmHiTZwxhvd9SrWJQCKz1sKacTs6L95t/eTGyQV/f59ck7Cct6IiWOHIzH4ee
6UqA4XgyCzIIoOuuKRryMCSCchd407y4AYMRbriEV9j5La+S0yZaKT44DArvSheb
ySFND9HDhRy7DJpiLM2gLw7MJMvyWFAvVYdzTzCtW8y/JgNAcCYqAwRkcTLbhqVQ
yuHusa97rvhKxdO7AtenJpuroyF9Y1CWLGwUW5Yg5oLVzIczyf6mSs+6c90krC1f
6iMnFUYUSi4gGbSE+meMyG4ahZJTKTIw21AGHzRxkoAxB4oSo1OcOaV7a5gwxDmf
6KpurKOjD5NZcc+YUUTHyqMtWYEKtnxlFJNouQwNRipmnmetHfHmlJGlJyjBxGZA
pS1196VLOrGQm47iXa9nRehgs1uNenvIyON+YpJ1LqI549mM8MOscM3z8cDOizVM
jdSfeqpG+jHp43qseBrwSP4SHOxjS/Nikbhcbegwi8qi7bIrYfl0Mx9AvZ4Ve6TE
SlzoZxQjaSXNMS512qRZce97ZAc8eliXwfTrwMmh1H39erFRpMjN+riiRA3dAOEM
oCGELKsoaMbhvyUB3tAox+U0WXJIdJrsoDhHY8QhOmuxmvLfLfkiAeK0ptYDKf9C
i2kkwSGhRMZVkyOeLFCEMpmvjYgPVMPx6sQbphGe4WizPns2lp57ajXUx/xLDhZN
KvTWNCA4lcn03xiPJNsZvL+2jaklqn+J0HoY5YNzwYGSp3Ev0GjANkePfA/jNYbM
XKZLTb6RlkxvFb4yEG0Bzhws/Y7k2S0qzo8yx6+dd/s0ZVUrAhfYIKwKf++bzwJw
nzFt3//hkM5SjJqxj/eKAJZfEAqkUsqBd4x96wz5kNLxfsjYyCsKALlaxVSFrbWt
ByghlVEMr9Fzd1jny95MpHorImEcMw3ZbUBf/To7tpMTQGKle71yIa9paZFeqweO
ZMri/SpiF7yPQ6TaMtFai8DC8Mf7aH0fFi8owSOIFaXapOYKkSUmWqyvLQZuRAPH
8nKgJj7PBaPXGEVtBlBvRlce+IHfHiaDNnafuRXXPIvbC3hV0JJrZ7MLzI/Yn2Ja
YCMrQzgr64n+ypMSN116ihCM4LLe30BxL/mUSobPAHGpDXeiJQrD6ibK03j4E31h
yp8Q31lh3EbRISwMIevYYsE7DP8qgWOU6dD1RgolGAngASFCGbaalq0elF6uXQlJ
sgy2uit8fatB9PqoAGQXBRKZMqTnyhpWdSY4rc1SA0snJcnBYe741UZASn54yZ0L
+vVEgygnt2oeZPBbT9WLbcjwJnycDUcF3C7W1S+dVSHBb7XtQAYdzrd6ETQHH61p
CL/aG6FOVFtQfuxiX6TJaE3Twu8PwHVkDKMzb3FSPplFcVHcm21MoTy82BGbjjzn
cJjnym5gxSYdXbwe4Zw6esrhJrArT4kYp3VD9kHcfuaZyyjfzqFl2Kb8wPgIKnO+
3hj9g/aQ/cwtdyBMIcIXROpW+hb5wueSXNmH+pStVk1+lxgd/lE9HHT5X/JFomj6
lFJIyeJzI5gr63lDaTUEyPml+iinUEBTZUkX3OqKUvy0yfOF/J9FigTmAs24veIo
NFmtOfxrajWGoHjBxGFszg+EXoyHNUnH6jm+Jw6tuofIhpU3qBTgIe678hSqlSTR
fdYotkYoSQKiKNOtxuXQcj47grixJleXbO0MgEJZdjca3bfrC4Qn86nAa/DzdnYl
UVmTuqmgG/3EBmUbpr8g+3u2Ug4D0bBKD7RqiqvPVEh2y28sfq8KTellnwvm8T84
OL9XDbgxJ9rH5poobj99vEDzmOUq4fwmvIyRvIoL1m7tHTUcGxF9Hi84F8HpyEGj
LHrn7gLKKmwv8OehrhmTLLPXmkPurhBOFiHmyvSO9YXUYjn4RGcOsRt4+Oy211tT
qSqSnntzjsjsWiMTuL7xbv5aFLqg/lMQUxZ8m14tuvdiqPUxGBYb5JGaetSCUbXn
5M1EO/HJQrUhBp0ZmPz6E4w2fyHmNbeTXpN+D7iiPzkdumiIfg6KcSgpEiwHwvVg
snDYQfqkBRNB/yauyECbKzL+WoJG6ksvS8T+T5Vy3Qp4ez2dnPzi3IFtsazHryoB
R/Vsl84fv5v9sId7ZRXRxGMMME7o/4DmNhxDNnChfMgoSrDrc/hLDRnMKFJBHEhh
+cpfTdVGtoBX5pMM+u5bjldtkqO82mXfJOrRfCsV1tcCVL5NzQzgevvCy1rGBhsN
WXAnIsDxoL1q44o0nU/4CoeHCtPMg1Cxp4pi35fgfjMd6hMnfzq8G6KYOvocam4H
w2RQUp4HNomnTDyUi06nMC+vRBh9wXLHUdSKXjDxGJFrCYFsBgRaWyyIdtEDrbPx
DuEcBYxsmMHFkbdLiBAMQAgQh5ZRL6TsQD28k3ntDtdBPEiorhmT8cnlqctEABAI
3w3b9Z8RytXLJt4gYLowAQSkvpdf1pdJj92eNijrS/mjqeOpjqu4SVi/5HTfSqvX
h29qavtO+s2OdtM0EI3CduO2ACmG6UAnXXIuSCULd+OG9U0Uw0kwDPMzW+USUmt4
onsNX2kF5T1x3v0+D5C1BEoFEE6AMObmqtxdNQ4y/eu3OFy2k0ayk6xVQHwmlQya
7hrAcMqMUvHg9GBotwgnozKe/oFP+h54g/l32sZczImHw5TmjULvYSrucJE/iMJn
rkeVnj1jpUUTxh3DEb5EsyhvzNCeMfG81lF+aBRRDdrdlKPcmGt+l1+8a9gTDAB6
7mw1L62XD93igr53BDRG5HvZGhNXgH21/tDkixH6rkaTL8kTgoUD5tZMwgLWc89Z
luZjBqTEdeS7tw/Zt5wuUyOIP0BNR9ypD+tRUba7qlrsPwpozxdKRrQqkaZQ9gqF
NlrlHbuqaTT1I/Op1H86/1mjcH66RqQs68YRvWsps2bBeBRRF/jP0CBB+mzaeb8k
PndLxdJYI58qHlFcnfYzR20AXMmSChPzS36i8Xnhmay7SdF6yaw/IqMC5oS8VINq
ZEXLXbSk3crNt+tBIgEfUbfDwu6l3cxPaY0b28y9LhL/Z5GGGnZyxaOYnxtkVEnB
8VE/okttDfrY3fkdB0dldzxDQ91qs8Q29ilDSLrjpDJiYbaawoM7G6KUTK9lQRJp
WTFy8cQnadSgvJ/5MeLp51wtl6eiRjl4LXc7jpzOrnBlwc78Vra0fGDrAGXr+Pij
Pzm1gixiXrtuKiLQX8Je+sGeuXkqDuAaYRYAlzhgb8mEIVvP8DYknVY3l9QeQWq1
z2Ik2NLCV/+Ywn9YsKA4qlX34GD9Mpu2q95+Qr9oNiEHQakdvEG1geYS3sUVoQ1+
lhYVlV4JfyDNBg2ho5JIQIS9kYFED/C5XjqdHvwMqhuYNj6JYTCDMnXMkvxvkEO5
VgO9GjcKbJ21UuZOKQ4t/DkM7Eu0+ERXX7NlAVIoazsDMclmDaM5NbKI3hycaQO8
NSZVbBohZokchjpAE4UqpxUHIC1yGk94fLi5bDdHt8WVEgwD43GrZhimfWu7ldub
28TOpffrl8DhF+v/INMqHGbGI4Yvf5/mVSv2AtEVilBCq4RE3X3CPyEM2qjXwZNn
VuiUaZJzkOLZUssEWzKsBSu3lt/JRMEV3JdGNszGJJUFmWaq5lpENA532wjQWW2f
CNtXXAe26ao63wkUh11taN8MTUZcFjyJ0wVLx29rQyprOIrWNP/8joWTrHpSWmtg
1xMtJGRQfPmOa8IVmD1Wa8HOuuVFGEcDhGHLmAxtsTABUu6HoJnR+flfbritoHUZ
wuP9Bva29+IMF/xJOCLMqAAVaX8vgdA/l1HeNZufF+Xr0fGbYOmvnCQ7h7yDeo3I
GbJbgO+YHhnEJKqlpplnsnjPixPQMxf5jyuLs9XeQJciTxmg8b8f19Ii4YtZupoT
cavegzDqlBXoxHnRVY9VyNyy+tg9RzPlIu/xhwr5ZdP3B2UbevUu3UQ2wPtYKYmq
0K3/vDFByxiQl+u5vNsxs3QDTJCm8A4G3Hqet/KW/GdtNNAT0u8xdNR0w8h2A4tX
ToDh9vdUUljVkRCtgA2ovYCwonfztv0NpXYioWdA11PybIMw6MfAe4HirMloCoAp
/TtvsBjfiVniSHVuwhkA385Vb/8FuwglKeEaKya8YnG5Fi+0UGFOG4mZLFteDJ6v
FOxs1j9GQYuahGKcvF0InUecdz1FqxyX90QOYrE1n9qjqJs4TwXyNB+nqvOd+7S4
eGgQC7vtvsqX6YOgOu4kWm6eWvXa4ZY24ooFurWI80zExbNAUHw0pZ83uC49w7rz
iZyamOWsyErl1JtJoOTj9eNmljyzJUPxyydhBbRFawwjA0TsWgmuVpSsgXPF7D7R
M0qS8bqOlmngM3gIfSHIXbiYypvsPCej3QGmCf4gmA6N3qeycZCc0j51lhjiPlgg
biN6F6C5f1h9kSYRUM5S4Qp6VsbflFGNWNFzZ6XMXd2B38Qm+yUpS5DonO/mhck5
KLLvdQPfDEY+OZ0ayOefxDzNDJLQPVKEoxaYzYfupT11VhvNcoAf+U8f00oKu1Vz
05CIqH1F2UCz5EStBQXtOc7C8x4fAQk8fOoJV8JNE1YFrktfSN7uCSUuqydwuKvO
SJxOn6CLS1cQZIpzSIZHaitNrh6ukiMQEngzAYeByPZluE2q6Z3WgNIU1wy/diD9
dyPDbUCQJG5RUBPKqgKqIuYa648EyNysUQgy9kPXYg+9f0VRdXjAVwwXxLkyeQ6i
BipvL1A64+W+Pz7nEkdRqZvcxMzD3xbS3EipxkOgqv+Yd5oj/4KHuifPlg4+RMQx
ZMKWJzvjdDEOy2vNyqqgg6EKgtS3XyIJr/o3yy7m9MrqJ3TmrXS1IjtGi27zA4Xc
TgOTq5erhfKKSjRpqu/xk5pXxrwM24BXrK4shfDNPlj+gsP0yV7L3VzHBT3Sz+Fq
F7DLtSUQtQC6Mc/Q0J3SsgyWyRXhwtPhik5SvQp2y9Fr2OxE0MJ6Jkgd9/irGn9S
D/M6O7S2GZH2qLb+5bjoSdda65vPifwxwS4whZNuFzbKlMidaBydvIf2oWUdsza2
DRMYOH9rCTXqMnbITOgwBttae8OFfSTAhxc43Vrmai0pGylf/EjTZK6sR9julIt+
8dKocdsGAJ8zoS+bjz+/Nj2bkJ3Lbbkm3b1qp9E96qp94V8G3YvWSWsiEeS1MdSx
3f16AMGnk/9X0BeKU6A5sVIsygXH7sPWRGNP0EdGs0eW8nt2+x77FEcH0Qzd1q68
OTrGGfBXJFdXMW1Bn2IzurUroygFsR3fWHRqAnrbIkIOCPtcvt4C2r+77Jkc/Z5m
2A5gveOFVgBMVEI/ALBghes2/aoDSq6zmQ81RUwvgFPrSebkV1JLmR1aIX/BkiwI
Src2LdkYr9VYkor3z7x8U1n6qXkflSTAa7f3sbzp4/iAiW38QDAYzVqxO23UfLP3
IirLCJlSEGrhoJpUFgn6gmJ0jD6zIMCH6Nvzp9/d0PmCfa0Zk/zU2XB+M7KH05uD
p7Rcp8wKRfxXt6fbAiUlZNaF+XTTpPmjllOdPrM/IdYM4Btv7fqLyQvp0tfIh8SK
bl2jWgWvSe6HIRz3+ZBkdnztk9VKYy6MuOsAh0T6Kg+wP5QBsbNioNQACtKv4Rhe
SpXhNxVzXfkJFavLAjiBJEW5IiTN7hmEmrCrhuwdFNzZWtK4CNmljsGQSOJ0Zh1Q
0NhbXsrr3tpMsbvv8YzQ2NzI72vPe1AUhiFwdMy7UdHZzwzA6rsv8KvTD1fpBDUg
17V7+EFLSjY2T2ro8MAQbU1EgbNMrMm0Rs4pwklITJkvjvJEWHIUBp5ezDhnDMqm
qvzvzUap2c6wZoo3HFbivXny+ClErnYSv+D4Wf4CyZ5CDfWFwlt2KTFrlSCopTYF
Eb7Be2GtyyoOl9HRlcA49w4aQ9Yhzya6nUuHPaKep2icz9TxCHeXpg3I1ck0TfcC
4grU1DGlBmzaD5E3q232+Q1Nen6rvqM9EYjUP1u7h10ytH6F7+fkIlgt6Pu96Rfc
o3owHgJpFPua35AmIQ1hiWBRSCsARTwQ1hHp2lvjCIXVEQUVIcb+rXiVfrElrEXS
QfddAtgqO/WQW4T4qVasJnT7MD23VXUx1q/d5CtylXzOd1GDgbXN8+IwSvJo0RsO
WP31qc0kj7DvzNbRy1ArXgLOJFOLS2Q3yZFPKGW/rvD45nEhsoPTUGe3OUzFhSri
/LtYfGR1+NQJOqkKgs9+ozGm3l49oeRIypXzJuLUxRUW2fwfmxb6cQ99WZ3MXezS
piPi72dLLzuLPAwoCejf9SO/zTNIPo7HuqIyPryej2BPNLohfU0hxgm8fpZ3A6RQ
ivlI5rLIeABrlo3sX/CkUM58Iq7GADMXlyHwtOrwDR3lxvoUQpltVtUCPyTP0HZI
EKQf8Nw7WkJKCOUFoDtVoP4Qb/8b18opSYRrDmNevEINrCpU1cMF2xVIQfeaiwy3
DNRECPujg+5+jJufVjX+4ikWLKmpDnGIuou5aXNZAhmIFJmo98zSTyTXXZP3zpqa
fLXhKHjPzKpa6KCM6JTxJJJBem3Ko+2h6AZ1M6c4PXTWIJZi+e+J2F597NukuTBp
jj4uSylhnlxWkky0hoB2f1kD8Jdlv8SC4CjGaoWc8XodSwJ54Jdw10kOwNUzVMH1
uNMCdLUKkodnyU5K+1Wc38OP1GL0zKVpKarq5T+KWeYZKYV/sPFMeMJ8wS87yvgk
qKg10I+D9j6Prh3D8y3QnYz/4uNjCmWk3Lzq0R569dXOWZf2iH8C+ADESouJGZdU
Lt+ytN19Z3PU+LuvJDg7iBycGrO7y491vuhWovIGsAOIUAQLBKK2usLnQO3DDHuq
oG3K8RSyi/hVx5sngr4GFcf8ulL+ixAtFz5OogoGzOBnYuGNK1Mn5VMxgYw52ZEG
bS2JtM1xfadAZEg7xHkTO69rRvdrke4Lb+y7N6lbjq9HKfn9/515T36dfQb74QSE
CDfg20MXz0pkWDrma7UwIsolqAi26bzzukkGeFaOTVsRZbP7Gz0n5/mz+Cao0AtY
z9MD4ltP6LiNH12EE/W3riXRUVPJX9KOntsjQNhrLsAtObioObF62RRl4gaoC8za
wQgWreTieENryOAUU3UB4MNxQCnfqo3pVUwMCKTDqFWVTc6XJka5FiwYhh9nBUBp
zoFFA0y0AbrkwVQjwumgcgQrtUdg1POn8rzWmgZnJ2j3cIoq5VZdQw8i3SMhpTOY
fnj078k9Bsg5CBzpqqi8zpzsUNGf8r2xVALaHtER+NetWCqQcYYb8XxceGtJ1OrW
JjolHew1GfXPIdqBdIdNeQUB94ihwVDVbwn8r50IC/0zTh/5a1k+fbPmyVgBdAQY
z3GzuCDw9yMq14HLJVo13MJ13J+hz/uut5xmucIV+6p8q7ODMBFuS1vCwWmjdp7+
wEGgkrVHbMfWo2U8XivbruSoAYwYFf6xZghdtddJRfFdC7XKQ7gTjVcOciidSVUy
o8dOFUK51i0ppzvVcIoRNRSOc7le8CI/COiQPwMI1tzjUaE8HK/QZXtLwB0e1nC+
mMEB0vFkRRRsFyoYlcGrxW1mVBfRYijkfk1ziNpi0Dpw4R19Ryo4kiaPdE9KKZqO
9ezY3uTAeUw58ZQ/GeiK3In46mUrgw5I8Z0hV+gbvPb5xKbbSUEdyVdCsEzSBBpj
buq/z2AbcItq3rLEWxd5veyyGlvwmzjzoHF4sQZtz3cw+RIclLulAPlubimBWjWU
EiAp+xgUzuRoVcJe4LjAyCNv/+3xM+4aMh8NSWLTM+RKYFy5dowVpnQWP5Uc0f6s
HapHZ1swZLxvikyrDuBm8eRi1fyyU8vezB8FFxYIAA2vDGtpgYM+u2CVre0QAlTc
xV4qXFcFE7zlyNtoiYR2/0cDv740GXWKnMMZ6KCLAJLjBXrGmvcU9cgx1rOslrGl
769oN3dsYAT698gWwTrWS1G89/8hiHNtngY4iQ7Jlo1rCoVjWPpRrsmZu/4UgMsj
RhU2TKC1xVKMs8LoHFLI5Jyj5AILqScsNl0B3KI3mDVakV8hso4/er4JjQgO3Wjw
g029kYtztsM7ThtaUndeBzUR81UehDCr3S1i4TiZNu3maOyUOF7xwHQaVJ89ZK2p
CKLTXWh4wc97j1HhuLisToXPWZJIfYiN6xn5dmvxDtvdjA999VNT0HeNfPsviTW/
WqqkQv/ROllyleAVZ2sT5rIqPtv0htg2l5a6FAU46Y4JEbHsMBjNuktf8XQ9SZ4L
/a1Fv0EG8DkH7pNum5mdNZK6FptFDT70tKfsJT+YL+JEFH50eSSFDYKLmHe00+Iv
lMJk8DviJ/nTW+sY46CfGfIKlaU+CKiXWt7nHbx/VX0XwqFQFEgnRgU5XmUb1WB8
F6j3Y5DiE0hMA6Sx8JJM+4zsKi6drjhqGPJHMXa3/I+JUdXTfUFDJlBFP2+9Rhob
HyPpppcgeE2qdz/Q2qvs4LN8VJjFUGzJRGF4AyjYW6gD/CJ8hbbLMs0IobUcavUd
UbI1WQjNYfo5lkLVtb1sX/hKCW/2r6YigXrYCRpwLAGLyUHTlXT2WWooqFv5SkP3
JzRhOGRzUFNP4w6GP2tv1iIQHO19fRFNedRTCuwq09+TpLp/aICZ8NqPG2B+AAPw
iNuZ84Og4S9pE7Rq902djE9CjeEDpfUwQ/B5L4Xfy/51aiCKf6TaVi6aPWphpv0B
BwVKi1GooWc18VSC1Ke5pMnVCygENuia8Ss1i75qtFQGdKgWshTArkcAZBSd2vwm
a+Gft1kCaOPTOvf9qHLjXhOHV+PL065x/ZL7daN0+vRoA8rkWBqFraS/IasvJQSf
X5Zp9qWzFZTK/ol3Y+Xiw72KVI2Njey0Jct5YoAvDt3RmA58QeDZqa9ECnc178Dc
bexPzQf/tBNcx6Dk6xPMP6TLJMrY8mTJZwWRbWzc8Ap144ek+mUkyRRc/xoHqSpW
u1d8HAXOhSiAdC/uyJT1E5ea/+MpdUn0o+2vr+bYYVE/J04aTTLiF4K6S2t+2ayF
SLCpQVOjE5Qip2k1iyx9sW9kwshVd0Ae01ykCkBRSwarhszN0folxg5cSPVsBnOd
4FKK+DNqdkYNVn7gop3weeuUFu0kIi5GvulIhx4ObQ8NR5fCArMEqPsmWFsR6W4P
/WT3JRGSOfNDdwx6hKPYGCRu5KkYtsNwsJlPy/tAGDhaveSJopdvB5XOOawCuzJb
I6YChIgBVdXI9sNZrmX85Trt7PlgiZMlGezbKVqAt33xr3kaNMaolLQzeFgYlKKr
b2AjMiPUVELkf3i303dmNl9j/vs4QsYPWFjsa2fBCp8OzXKP0cr4ZCDXKedCq6HO
2gWxUpouAV55DzidbsSyBGbpJm1uUG1rGxYMoMzFrDaN8ROA73aV6oXyM02nKfhz
7rGIHqY8JFrSFER1flxtDOLIv64Sxflnvbs4nEAutCRWvDrJPm62WlTmOel5v+Bg
L2i0vIy/zaXcqlGVkNzWHvDqgtPVYO3sD0q6Map0YBQWnz169PUyRUMrXv8EVjqe
1+gK6vdqQLfp9c3tgYP0S+1KRThgrkBmc0AxDuoByhgsB9MDKSwqnNP3Rqu2qy7i
gT/gfOOBtaUDacqkO0FWB3OYYj01DEX9qzXdse95xSet5sUASdViomRMIpYhhPpa
du+1ZGSen6/4jiPu0MBG5unm+SKAD3JoKYWZpAj/LIMEr1/xOOlC3gMyQGtztokC
UPMmqDNGOnnZJspJzbwhoj9go8ZYesLBYsHcLXL3oI4FsoqMa5TGMgarCJl5IefP
ESyPyp9zQSpaUmyLY1atzvpVW9/6J6xil8AW8EANyN+9+iVRLp/Ty1gaobDMrPNW
kF0pLEdIXdcI/N0zOH1btbjQZbObEcu1WhtSeRlal0oLLrAQL3xpremokvu6JJk1
XBi64qIp44rOP1SNt4lcc3u+Rd28whly+pTewCwCW6fywQwoHvDtSFE2TXudTKkF
6d7se43oYSM33sNzIR44xdtuX1PxXDcnN79xkFK8uqbOfFYbTtfX/l/lJbWfk8DL
T6hgcbGMhGPdhtewYe+LQfVSCmn6bkG4VvxRZL+r71Dan6y6Hlt4YPnG/9Ts/Toe
BUPJoBAnij1LLs8U7xeGIIh+Ywy7RS6FaDVfgNiG/TzDwwEp8vMr98Hfy+2jMjeb
muHelK8K+pyKuba6n+RrcmbmZzF2bQZh2Aysoc6m33CEsXK1p/bkEVVdq2muT8Rd
BWrzurhFRL69I877DKzxYZCs/wxL89W2ji21GEf8ImZb23F00rn4TvgFI3dl0fM3
sItErb3RcNjIbTyLRQL3JoTb2S4mzIwwIrrRvJcYJDn4uj30xM/Nz9JDH/Z8LBrU
doH1gkwzVui/w1jlJ5NeSffPjaJ1jvNSRZUv6lw8byo7GI3c17CFhHBA/paXbaSW
bVcv+06gwMGX9SaiITyqyq53ECAMb7QYOgShXzbWoCfnZCaPeO1LpqAZLxWFDV+a
n7u18L5IUnEsQl3M/ktLi74QTcVnUm/S6rPT1Tvl+nX0DvYpFDc3929+tWeGeguq
gXkqW/d3h8zseKF8chqvv43QYUCEYOOL9Rn4NLEL8yathxJSCqMbk9WB4rit0K1w
0Wcjm0MbSLSo+OL8Dls5xqv/CbfVUkqaUomRWWGU0CC6YU2/uV2gMMtwsDoYySIu
TRDTCyQpAbz+0RUnAXzQv0+lsdPzmcpQaMt+pMVqnyEeFI9K4UjBUK75CVoWjvZj
t6qootfgBV5F/T5iwCtlX1haIlm/BQty1YyK5qgO+skpYaXnu6CfuCd0igaS2Y2w
D4ViWH4GWqoElyaI5EDmILtlJI2B69Jlw73v6V5vb9u0rrseju+doGx+/NTNS+Ip
6Fd417qE1n442NKr1fVmlHsu9pyi+VRoSrncrL8Jb/Mh8Nl2aC1uI46aSzIWuFXS
t0d2LxP92jxWnObkbT5+UbkaeC3sAkyUuNxmAkU1IoWEfFRrh3FeHwIbTuIv1IAE
jKYtyVD/vBx3lLyIDyBY5o2kIHnBEn5IdxaeFtlPjxefy5jy2DBgpFYnWH1LhS3D
qgaiNDx3/+eITT/y9NvfC+2gJL5FwnyqHjD/JGsgCcllFIA0xe0v7JNRzqOTkW++
rABDKug8LOIoXigCXp4o6hG6THxXJwQU+B11ytksaTzwzXs868okTLvqHlZ8FL6p
sgZEUbvDF6885+LS+ZbxhfYSzvkoUFsI/dzPEDHxULGSam2Jx4BE3T+ToADCbxVv
ulz1jUb+BlwxxLCT0f04h9QUsWdD4F9gG+z9z65m3g+tKPR3EnNHPjAtNtzov6pD
UFirGA+AK7L+b/2Jq0s2uc6sqSqOyNC3Q2uVBjITajeuRGaL0ZA/dbXz7MSE8BLh
cMeireeBQaSyZLNN7bZk56ED4YEm9HoFPqpORoi4D/tBzu62wAAFtTvMvVE5/CeA
5ITqkSGizcAAc3Se+f8JG2RCFX4SQTHEOPobh4MfyTbqanhtlEa3gkBKjo3I7ALs
+X1vsBHTXURGdTPc7WUUpakVuufWqvQfd+uXhIc+huDutXT6H9dIdBjdYbxcBt1E
O9nmK6F0BYAgufNXAcGsJkB6cJpAHAVI9JvIzMBYmJnkPqz47rnA+QCTM6+Wiy7t
NIDBMexJ6mle9/N0KqqGko47XAaxT406LNzQLjkmMleEK80Zhdb8Yb81cj3Ym44n
WtRmeDdhS11kQB2ixTS1NDZ8K8n5954OUM03HbVwI+1Fl2tjR9SbH2bMiXY0lpcY
yeq9uWVrDkj2yjD+mU8UPNXhV/r5BSSvz+gOW+7wOg9kUlJFbzSeka39zmQLGznS
qtZbKCpsu+7/w8f4TO/PhQ0aPIRpCtKlbs1Znwb+Ub3/S1E5eEEbMyyWUCUl9BAO
MfYMvYBn1GJeydm38yBwnVxYXIui0ac3bW4T1U/oDyt0lMAkE9h9IU4LjnuIiLP9
8NnQmAfDbQhHx6Vb5XOBDarIy+YQFiOVkmpJP3ArNgIUGtD+2ft8SyPfoy/Mddnk
ZHTFIdMpNsp+pIkxV4T/HJ7urjmPMEYZm3DB3MSuU8qWepK8BQ8Zmr/KaqiqeOTk
xbZyAaVSwBy9DRxDT6Ms/FrlqVYRems0CcJ7meLmDdMMNdvZNDF+eeoERjDGt/cb
XBKa2OwzhKdND1RkIPMjgSlzbQ9AQswU9iBYGkyjT/cPnGzrRyWBO4ftVQbXS5WY
fSSD9YzMcJOZKu64NOqU0ocYviI71PKhDDgS/alKa5FLGlpKPJ9hssfliFdAGoG3
Rcr2jiUw4tP6jqGBOT31I5IRKo2nU3UZEuE5ru5u/U3p5E5dfWE7BekXdhY03lSY
aVz9XTnYZqt2rnOtqoyqGO11g1wFqEJcnBoXsPZTzSq/gPnftuWAlte0mKpM079m
+a1/I49cR9Xfv12Tt5yFUOhn7FiMKBinWdUBgxLDkC3YPBE406rjpWUVGBKlStr3
Z2whjxTNSXco/0Ghk/xQwMi5HK7zeU13pT2WpZRuPS0aMER6GKOsAfu/t/oXcI0F
OqghY219QvuJsmbAQNGGI4q8Ee5QQ0RAWU1Myc3QMy5UcaDK3k2Rd8PqrPjY8Am6
TOoyNIo/GtrApFneEGrzB/lxh2evSjdndTIVh7hq4rplCDPGtY39zZO9CWqOq5mH
SdBeUzPyECeyJ61DG/rGswzx+2BV2o1MCRlA6XQfWHGQMERtXRFnG7hDAuEepcQI
tXWZX1UkGbYpTsJddwhTtmwpMQFruBpvhQFRSpp6B6//XEOM7F8jbfy8rE+GeXau
unGmHIhawnUExawAR5xeQiyfRe7HYFkq78GGXd8LkWZORiXGnFKBL2s2i/uvprLj
a5zYXDNMdu40UE/If9FCdSCMGkgPkfk+Okm13xTp3WXiMjn8myb2gwJVM4YUGh7P
zV431gkS5Lp2sfjxNgIfNVg5uk28B1uJ7Jc+ZKe4/+DHFKe3WSraV8TwN3aunJZI
UqEUJDzgQBgj3zDiDJHPxoswNfJ/dOx12v52pL9YeWMg88GFjM3ht6CvSe0jNREo
+d0dO05qEl2l92kpWmF0GP/r4xDUFdl+srHltTe7Ar1IYeopMRzqzv6rWkW2ivsw
CbrH+4cs8KuksSEwfUkzKmPDuwxS8Q8jy9G6VXTdNLCHeflU3XP4Iasp/k6Q/jUC
8rIepzDs3422tzKJfA1P949S17TCbs5pK3aUZLbjSAiGJExlb4QCO/CgVH6A3kPk
Piv7tOApHlak7qYvh0EdYc2rChCMgr0lFBXi0+JixV/Co0bcb2kCiYwnJPuuy/Az
kUxJasrPfwtsr4dyeJdgQ13exnS6PDSjsLfHC9692Yiyio9XssExRTGBB0WZ9bnR
ykHfuHXs1fA9n/OzjGXl27HSzYFhs8t0/+XyIwl+q7Xq/Jh7yZss98LIT2Rrxxsq
c4TdcTqKk3F9YtQdM1ONXt6IVSqMtQwHnyDWzarsS4mA+EH6PZOLHALANf7OlqwJ
IoPqlf/SZh9zJDkZDRkiNLtCUUEJ2F3gvB0xpeCMaUYpc5k+oU1vSxm9WVcp13hW
42kX96VpgkVfNysEmgFfPPK4wHL8ckh8FdaKpIieA8/cp14O1tfkqoxqkaUP+WeD
aiTdAcddXwgrf3dqzvfXQ2nvyuOJhutxS6+R9m+Vmvb8l9zAEXbuzZo+VuWp23/4
cY5uh4A5ScTmEaZozXvCOcbh9YO4cCTWLjc6vjsZLP0bMEau6SL00gZsurCeosQh
kEAkzz/EkBH9P8Z3844PFyTL7dfZ1sRFbpEvE+30VwQWZKR4lBCUDp9v+smSqIV+
yH8zp7ilLHzg0xdtriRjGaUW9gz0Tp3gx9RCPfqABfiwc7BXcKXSGSnYC4Ee0KWw
+iFBv7kAAcChu81Ww5HN1voWmyjJQZzOFwnS405WXv8uUDJWgvjDoZjaeEb3jWlQ
l37PHWsXvZXnzNS98hwPZBBASr97N9A0LT2FcBpunWcbhlz7VJuZP3y6Pxag70Qa
gqekxTIIHBLWF2sNHYehMnMJYeGexUwxpFJvOyPn+VqhEZx9SNotFwYh0zN5zuwk
UBoDcj19oiBreZxrxysXHQzG1/yzqL0+EoSA22zWhhb8ald5HwUsKFiX6weBqMds
YvcIg62Ja4ZmEznkHuoeHSQ4HXeH3XnCakhmgT2NXxGeKo0yeJInvaHgj3P9ywUI
VgKV7hco5kBWRBUnyTtbOSjJwGGWuDP1q4MGt89LwrjnlZ4yn00E9N7ErubL3mvZ
9fyA2RHyQB1NpYdJLWhemZQAwE7FItJ5TX0p6q19qIfgbdMXVedefwaAdBgtGwb5
NN+eqLId9kejsaVLR9oYlYQvfkk9IYrHnwOAvuulwA4Nda7hdX1FSmu2Z3J0zjzX
WNlbmab9TWbq70zsNcFuJ3AkEROltf/fPi6CjWAkSOQ5kUmEzEg5uabE16sUGkY7
n/uT0DsfuH7mIYDoGge3QtHzsK9W8uJsrlY4RS7nvCahBHnN5OpyJronKbzBo0K3
2MQrXiJA9buXEXmrlVoC5i4o7GS/FM3yWHRWTGavAoFPrgewNkMWN2DDroAarQLU
mL1rJ9y77B3yi2Ry5BYlsUNrYt8wDeGhUR0PKJ9oINadI5v49RrO2XVzaKte+ONs
rSto3GAvZM1bGFtDWDMNU8aIb9KF8Jr7t0V0AcDttajMGIMaCVQCbZDdGPZDk8Lt
8koN+CqEm6jzxrUq2Hq5f7adeR/DwiG5s6DvZ8rQzw6qttWAAgXM3fcQxUo3i6OC
64QoyT8XZgV5j4psMLsZQ+lAR+dvG+IzQJsgmMx/sBvUq4ksJhwWGVgk3a5WE8KS
bSHard26egKYdipzHHzdh36hquu8mVa/J3g/FGLROTgkJAz83E+rC8tliPXjeM3w
ne/TG8ksrIfakm/gdFrCc+tzOS1XUH09CuNbA8Vlt9uq2V9nPLBp1XU3FjtTmr/8
mBdTy1I2bggllCChSRsIaA3rzO19lBioK27IrSywK+IcQRrjSG7NR1SDBX4YX95A
AolO6qalmsbvjWHMo+APSLMmQTOrqQwI2nJMev6+E4baVZyCCVXpHTGeNOf3ZIkN
8w9aTq8Pwcr8NvntTEXg4F0P2wlPk5BWGukWuPz5Ai8MWgp0CZVEPrkJ8PjNQOey
WeSMJENRzcgXXqPBkNBQ/0AVAIrf2lHnnz88gGAKlmYpOwqY0RY6HPkWyu0DXCGL
J+hK0wIjzDB+OtOI1ifrJhccyLlB/4u8Qv7MwHN6LB9NQalbpshb4nFXgYW3jjP/
Xevw2BFOceBZAivfO5s2ACql0G8q1w54np9T3mVjiBZfkcJ+x5jQsmgwQnEf+MJu
A5mgbopsXjNqzJv9JA6yFt8szUvO82W/6bvhKmrpB6WnGhTpRyBcdsLTjf9d9ohF
CjBdCWuH/YTzJZQ0rbRN/jeY8qYsqXcRuiYN2pNyJXvFuQu6LPt7Mr3AzyGkmH3B
0jM8seLrwzzX9V3lDBAw15v2p076ICbZVbS6xbr902UoUK8zJ3hnsYok8JdsXYSX
6fkWG8qQjeyCq682z1BPl9LBkgnv+f5Ldi2KphHJh/99IZAVl0kBDgI72Tr0OOke
YeBp1hlqiUwo2WkZujI/ExEKCi2bUka9bHhb2vxnU+ly5rx84Wmsc2QAdr0GuPcJ
WE0lNTtUBeeM6guLIfQRgt9DAue3ipgLOk6wlB7qv8B3el1Fe5NnZRWKP4F/T317
whZ4h0kFxj8XremHMkS1+py2g94n8xfcaddcR7mCbpiug7VAPqzwnl/5DFjS+q5j
mbyMsDbidQgTQFKAN4LqonPBag4OmdJfXAHlUDBPCRFM2tIL4/CPyN3cVapdwjAH
v9gtOXqyzcq8iy1nMR70LF7EX5U67tvhrZBw053z4ItdseH2ZPGAMv2/3ku5D3e/
SpzYAHsOALdIPRah6VkLxCHwCcGblgVnrwCXS6ja4xaPxfprK8xaIYMXeCgk/w+O
FPcW9jgd57/Z+eLx8mTYvtDFzElBQk0vB05Mpc6EX3zgtZ8LqUh88lusO0j717+a
Kw5onSEZIsCdNi5Qctc046z+Q4g4E0sMAXnqpVaXr7VKoctzGv3fhZymrhLbj20Y
dwaanjCLRLFns3tdYMH2NSjwLkapQXKe6lzsZxvyAqKC99xABB+BXuamwind0qfo
NTFNlOF0n8Ce+h8NEhTZ7AalZcGY9U6C6AD2J3DVD/nTC+zYcgl7QL9djvEQ5lwC
TlHQtglKyI3MiwhxG4xDCfRvVeg1epJbFFnrtAt0WLGRY/LXbGImGL8vAX5RSWgk
qzCDXhNshBRv7bMy9Tmzl2yTPpmTnhZDRRoDbvgR1gwkvBaWmL7+nEJiteaf/eLd
BQHaGVGuZLWYrnkJQd9Qe72Alkrrcc/iVbER6ezmkTWLHx4YSQkpFCBABBtWxQBn
wSdGzD4NQiCnnD2gRMnJvW+AeRCCkmFh98I4AaSJ9eprlch2L9M3B3K8ONRF7NLo
N8XxDrZ58Fvik5Sa3RbMTrRYvBNMa5rvxr6tDO8Q/wB8IAG3Eq0IwOE+uFUKogBR
ESg8BEAtkJwjx3P0iGPivhXFYegYTpkl8uN2kmG5yvLfS2AHMWohcDkwN/UVo0sP
fvtBKB3zA/qtJq9i76ZEgkjR8jBnwCbDaxKc61HiQVYxqnaJRN2FTtjiCrceHkfn
1Ee0f/PQZ6cKq5nUteod+JQQs0LJ7YZlOaVo78MvWpEmTbM2Spw5E86CFL26i5hk
/icjimCjLBMTTGj7LT7fdG0wpgLIfmHTBnUV8zTcHvTDSiEjyZ07ZtvABMj6MkVR
apAAeTDyueUuMh9CsKGaaN2+rRF48F0j1YufxQVPNXR5f5R/lYVGoDOxcSq/+65I
kkKFUDtvXt0fNflWmaLYo/ywjJP4ss6mIqejKdgqC6LTxLLrzRqUSeUmcf9rq6ka
zjObF3u3XaH6k2x0sFlJk7x5mYAwjaChEGOwMEKs2TY7g/Q6lHUVkW8bmIhHcXp8
teDj/hwWRYCL7RG/9cgLVcp5P0S5doe/koxCHuqdoDn2cia8Zo8WXRAtw3ufkNYH
EoPpB6RwNvQpFBbKw/mpnBDjw/OyJyUVPcBizogA2nsJJpv2p2AoO8TjY1R/g/XW
Hje8UvGe23Spl4t3qmznxVrlLBPi7uoR5WIf1xDOkLWif8M72vt1oN/dl4fE7kVp
G9XfFRNaJ3BPqsOt0kbasReebG0bptbcPxgGr3vGP4m8MKEaLrQHO43qeHhXMdmH
PmVf/omxEOYaQx8p4scq2VUkMXsfHTRCtsSksjeEd2yyZGGSgyqWXh1AIzcXfkgY
iZWGiCzSK495N7DiEltSM0Wy5/2g/5ZnEsDGY04mU1S478rtEoW/TIGlus1kbwSX
l0B7vdVEk+OkF8h7IdbKYd0vMr0EuoO4mXzuUPUFCbTI2TYZkrau3sUqs6odms2Q
5DQ4mFwc2YWvQ5dCsnXM8B/Z7Xla2o4xoSS3DoRTqkJfjVpFuV75dJUG2MZW28Xj
jyh0j9xy7YJ7tGSm+H8BJzfkVdOUniVA3i+WKk/lK56Zwe6MKURM7RG/dp82WibR
6qrgocSRSFyEBD+YLdMzrQs5KaPvIzU5ol4BHbnJWdP7K+tCN548JPrTdjetUdgA
DTJVpS49+nZkyskwJUBEi5xz6gN2WqDRUmZv5oFhL3lkcokLo9QLEijMR9yBzK3l
8TjrRXK7D7+QNplWkeIzmdIV8uhrQC/DYD5eqCItNtGlqyFVLFv9nhMDVqZ8oWxF
IcVlgeUhr7TLpy8P+vAPHPpd2xz/5xTSNKXo6CpBd3Gfvysc2AogyLkFY+mLPq7W
XN3R0aIUykCyyXfeqd4QA+N2JR/quzPbSQlqF3m+OTRoUFrnTrumuUOkNA5gET6y
/Z89FELr6q/EehPlr88A7FAkR3k3IXhl3HyaF8fO73ZyYSoY7SQAZY0PcDnD6uQc
Hz4QATZF3ioKIY5DfWk/aG6n2eqzX3S8DA+yGtAESYKqNRjQg192ONQ/2g4xAJmM
OGavvZjAW4aZsiy2+6EGqSKzwpk4WVnRxNldXBdEpWKMitLWnedI+9B44J/aTuFr
lVjiIhefh2tpPVKilZdXtKILoJjRrs2IcIyyanHHVeAigRpFJ+Hy+h5UL7/A3ySt
d/craKp98mMp+tQX7V/pFEq3lsL2NylxuAd7n/3Ut9J5a6e27uCenBMmubT2RUoO
7/NKQB3S2gNkpLRnoVT/9DMrnZdIY0ffiUgmu4UM9MIIlCgAuzZXfU7BVcMS8KLI
dgnsx8vWbT8cSTLC7KkwduCeJ7GIADdQNumC+QVSwyCE6zFA4XyxX06ZEqCsDdMZ
TniAap9w7NU3N0SnF/vFcqiMjAwA7EMIP6n6QH7BpAGlV8aXanQfYjc4cEF/sBMu
yLtJ4atNIR+NWQj7tXw6QXKbztA9ETVKs2/mMK6W7Uerr2INhNZVXZRicp+6x579
xyxnbIesFmrnOEgmvH2p5OqrxvimOLItw7JQdZl3AD3AKulb7Hy5CZx7wOaWDpdt
RdK/quCR5+ZFDgNpT9UWY72KLBXu5pnfxuVGzEJYpTBSGv9Nry2cttFYIRVbDL8l
ptF9EPh/OzDP6aiC+GBKClCnOeOjz8aOlukTDsoHjjxRAlrN0h7IbQcRdOYNctPK
jwkE2Fn+W/kQ8f0qBeS4V1ixLPSLw56b5W2Qke9MXWc47nY1ev9GgLtjFPZQH8JF
4SJ0JuSvvqI4LrrfmoPU6jUmaRUDIPh+Kol7gxale2GHlpARGJpj/XOaqWB/8L6z
9HNEx2ni1dQssZWQmRFyIY57nbATfXZ7sngYjLs70hQ0KhDdFkiwcB/Ta8wPXxuz
d/3aCRQEMZ7bZg3rv/W92he2r2RCMkVBtZlrzHkZTpUmrruxpWW4pzuzyKsYyJhL
uGy2Rz3M6Dpti7l2PY3q8rmYyXBihklDH5QZs3GB0if5mltqx5PvOqnS2EjxiDe4
duUqjsoNzdThJNWZd5CiJP1etNDtH3oHwQ9mVI+2KtzWGPuoPu+D+PWQOExuaVUe
FWmUF1c7fk9U2bCiN36hgRkyhEgYoegjwXVbc7cPC/Ti+HGNUMyYTNX35d1wjs92
9Zk+kJ6jxGKbJR0vrDzQvtEQSxhlXgo6o3/O8FufaNiWn5OVS3IV6U8BFxp2uFTd
v/fTSps/C1ErYwPOAjsgYHsWXbItPmBUHPT4WPSkP2zxUSHGjWbhTXvWtSWsvFNd
Wxsyj7sr2m0MzFnGVWqe6Zwt5Vi/F7dR2rrvfuKUVzkILY7P1pWwES4dC3zh3U+o
x0EYNeDCczHiVLXO+aZFKu3oRaOg/NbY4jUWEH3OFPwCf7H+76T9wTVLLtI4ID92
31U6XmjNw2TULiCRK9wTe4DbXTgnm1zjf8X1gTBtEhsK6Cg46zyEOUUpqr30cjoj
8xaa9vqjE5wyRV3x39HBK/pbOJHvojkmzR7mLqhBgqRADwwz8MWubUVqZeLznF9t
7G0Y40MN9RlMurd4lzb/ngpXea7oV5nTl02oA84D0rnbBHfMpPYVexgekYiKi0UF
M/PmOUNKhidANG67a5mIcbzA70Ia0stUUFQN884Aq+Zpvfi84AWdy3mK0H/IaQm2
NAMJrcTuhB9LAtkuNBaU4iAUtjM7X6MnxZZS5ajd5RFA00hFJXpOQlvPVJGmWbZ6
xljAYFSGdBlF0UyU0rHGSPFrztrFziAlWZYIDk5PyzMg9y1Ro+ZuCi6mYX5igTLn
ZOEgYJQWcVIfkZyCxouI6U/U5J4oG0+Zs+T3j/t7HV3NGBjVf9kK1Pz79p9BWM+D
Qu1freo7wxpluh1foNNWmxRnHGrs1H8fPr4yp/YUA9wYSkVEq7a3RQB01v8eTTln
TkBOhIqabfhp95J6qYxeQbkd0e9b+lKKC0aoLQPVKo03aa9jk1vYkVzEOhz5cPbb
QPeElL0kuuUs8OCoLeh336HtWmHmg1n4N0vILjxz6NUeTv3EbcMd1APD96m8CjkT
baeYhcLHeNyvoZNFdBiyKux9ZKB0119zY+4xsI6FlcEEpAKMEcw4a0CAzCbrroON
8IepCnSzsozyfczhk6o5WRo7RjMSZHNvnFSpiqeNlDxB9WpyE2ao58ctVtLs/+5o
OsORiialLA8edfcAcmWA8COxcdkRq1FdlZoik7EbAu3939ePpD2aXu8zTKU+PIrd
OugMzQzMTQfJFCmKKINSQBMl6iszeHeA77d/gdIGDFyniY6mfuhxURGIdEWX96Ph
BEnU16orG3FKqu3Fg9ucj8F60ql1AKGENvQR3qRtRhCxS75hjsiAM+L+N9SBY7Xd
gMzSr2a7nJQoBq98SkSQjSjFuxX068l/D3uG+9RzZ5Ou4TU2GTAHw7jUw1NtYSLo
cmeekRWsoC/t7B4bkYpQNkJn8E9YEMV6Q+VI2O70MpTvYz3daeRObMXbJ/4v+qRm
lHZI8/WySZgh4CRrMpggj/JIOPReTDR7Bzno5YxpVIXhOIN0Qpxvh/xCx6qD0phF
AbeyYhqtFrJ6e0iPjNwHriGD+axeEY8arD0d8m+xl+YvIjMzSq0VSrufHvHasrXZ
j3M/fvw8xlFcPrmaKUnQBhxPEE55HdYvK62oNFx9L0BL1pnhoYEM6CwU1aODqjPt
mzFUoPZqQ5RuFU6wQ4WK0N5wLWJDDqUnjqeyv9nC+cTNgBadXrKAo2zLQYhUYyVD
qOTayCjMGiu9uHdtRiCmb5jWE792ih2rGaC7WdgaYJcjNBzVT/Uors8YPMH35FWW
lfComisC/0L1uPFLjcWFhmFQOLIf8CauyItgllVEtOI7NA0OhXMtwDaUnfuhemh6
BI63FNXWSZb2xX1EAtXwNP/qXN6fOZVpMsm4+xBCvtenTkY5s2EBdurjAd3N5ZfV
+5o7JdTcKyszZZ4vtKQimtUuw/UG5S8r7vVxZP88WW6FsnyRFqz/wG+wMv2tDsfg
h1ue87iZANzlexzC8AvRAJxvz4paEdzCo8qTONSbkyXVzvXorlQuriIWsTyt2Bdp
LJoTXvcnnSH/0Fwru3Km1qaIS+rnEEAfNOvE/ZUwyviBwEv8NEqyN236O5ielWSX
z2gS1U0TbF3+Qd5znJatdQvC4H6YKCkW3kt0iyQhRYsubACmNTE5um44HmSTILzT
8dVU0mvqZaHyv7XlgeNfodh6esyfdeSujA7Ozc3jhwn8MlA4JAJgAyMSx2RUBhu9
irqUafjq0gZe+FPaUgyejzVKOv1tvxIEpJWK84hzWXERvUu53cV+qdDxTXYFjlVF
3F8m8hCBa5lbrc7TLLzkQ10BMcChtEe8Vi65xZS0wCISMaY5HWHhqvvDb1o9/WTM
L4emQK2WqBPHwwN4XLMMLRfYL3X93w9FIWp7z8pTeYZCNiwxuyDj2RlLQQ+f2N/A
7FwaX2MGoeYg7e7dk1JoCby2PC8FZryAXdMx+stOU5sm9e7pjv+CPAUoY11/tJO8
yQIkLoOnkAbyoYj76oWgcpVYBLXFQanN1z8BBm8yAEIrPqv8KBBUiNn02hP+9Rjd
QSpaTS/h+qdHr7FiGj2HuibbUUHbky63YJqRuPEnQFqIe0JmBnQR9bIqAEzz/jDL
uj2lp1XhSibYigvhBkWEUbTYxt6of8LsG/yGB3PCcYap8F6TBDj691MtG0o7rtIN
wuBo2M7D0tcRcW/cXNQx3hDNyMeBtA/639QGU5QNWNABTmViTW1ZaEupyAai2Zs7
P0kZd+p4/4D2hR4v+fH1DZpnZ8mg1yvhHgwJ2ZmxZLflT29PBYMk/8u+BNtlvZ7r
6qBtByyZTo+tCGSkexZcAGIQQBn2YRf68ohlsT8MD3MIN7eWeL9fh1gwFXSnwmLf
exAy2SMUUlbjtiySx3aRRrNvGMub1Y8kITrL/9yBnl8oNQH2c0CO/X3Ot9QgpI0a
s/MGc/ACFJJU/HsUudpdxDGx+WHDGGPeujKEt4nkYsfhe8PPlKI0bAaFwXSaoXjz
I935XemtSEOOhqZiZmrNXqYPZNNfqyrUb253w4X5Birs+adSQN40hkQoTo/g5Gh5
nNs7eS2ZfS6CwZDtq5fIpDUVXgKRpP78rgc+9Kz0zsRbviYAjDXvhOhCbL5q2/T1
GXduUwcRMJcyCUvKTIazYMHEglhpE4pFbRmiFuVltLYSzaowu274BIv1r3WfGlbH
vq7IrwDtqRW8tObI122J2bpS+89H2wCsTIgAfDIr+EXapfdYKNgVIuzyNGcUYhMn
LlnzGUOaPYUqDCbobqfPA2YiUrVUpMa3kF4wzLXokNWL6ntUXSbWtNAPrQ+9o0p0
I7MV0P/2LjjoPNC5BwVXlbBFUBLydq/I7VGShw6GGYfsROk3U7qfJ2z2rzKRQJuG
MncFG6BDR7bYs6mkbsqRdNOPPEybbm/We8DUTaZ4CaZC7UcQuYHv/GHylsGpcHSQ
yc+EkjOXIT5usm96Ywuoh6rU+oBsrp7paZbsrgIycd8waY59mI/aO4MRTqg1FHLq
ByZDLv3Ng7DvQ1T5dnaO4L2NsPWpt2LUq8p7ZPKy8rt6S3YnuTQveCXQptQPQTny
qnETdlkR15t6iWgrZBPYS8l2cqMD5teehKqwuShJ9/PWapJI2sKFPi0EU4GdLQXw
INwHyQpdPtbGnuMoEnYTsamswF2mhIWxdOSzkqnLLsm838QD/Zh4KL1Ix5zx3gwv
Y6tMHPOnu5BqhrUhMi6YUfVAGr12z2IVtcVx67xfzziU7c1OL1ocojwP0QGlSISR
CUeuVSrc6g+sbMC5obHP9W7yrUlRfnJeN96JFNhaCPJZ5KGomYgrTlhYPRJLm6Rt
7VxZnu8nZ+8iQYJ7LVmKERQfusgPtsVOX2GBQWAt9GKTCKFHjK2SS1P/Ub+ihDMy
MobKkb1w1KGnFwKQSMxIZ+edkFe4vUcOAX/gfuWi/fu/yHj5V/4IZCUZr46Y7KdS
w51NniD3f2C4rK29UueJSDOJ5LqifhjJlnkWhTZh/uvABDj6Z7ewSNFvGOdoR0Bg
OJiHMh3W2weuZ+GCT3mwb8rT2kG3tXMY2h1KE7KLK9xE9IjB9/5JbrvlyJsEjiay
eTYYPRnqAqVUDyp8qEln5BJMLNZWWE3JC1y1q+4j5x3i5d3KmKDMYPEWeJJks5sF
ZYINS6c4+EgXU+8BO6emeD8J8w471tgcCgvCsiKweEPICVi4rZZGcUI45IISXLZp
Ev6ecFf33NPdvUVqR+50v+cmgi0Cefh6iXYJV+pB7F1syQBCg3XFdhbevAZz34Dc
XO9rZLVlCedxR4nIQVpsik9QXE2oMFuO/TTFgB9CrzSZ2IdL5rK7gMWUCq2N3dA2
mJJ4QVfRkVCLziqQaE+c5yu7cBzpvlhlwGSv7RKhR2hVIGNxROy6VpVVfu6ku7xu
D6L2nqCzJxeAEiebUEql811DzaGQRgYKpI98gU3QKW17iyyFqU9yW0mejiVW4QLJ
rKTF1O6tYz560vkC13jUnYhAAYADzEsJYbyC9oF4TVXbyarozZ+a/0bycuWjRQ+/
lMsCtEDqWWkScLhkS5y3FtQjJZ0ln8aIVRH/3M9wP8up69xV83Zh+OtmLB+fn0C+
JaUv57+FoEHVCy7Ru4Ux4XmYkZqdbVC12Ud5xDJO88K+uobvEo7aHjE4PCZCmcPV
S5PnB+FfbKNltVCXKg2M7gilVnKma7o/iKCf+UWnEHDVmoTOPwzIrgRR4e7/QmGN
E/WjDtdf3Yx+v94C53+5eAItqbF3S6LK6r0JTPmFFYGcKEvj9FJ93i7wLBW5PPw4
nWv+cHUxssf/1VtfP6NJCTdEz/WVO3/Z8Q3Nd1BdkZzU4fmRhl79ACWktvkLQYh3
HPMCgkE2/8mqboIKXAfqZQGWtM9tuESwr4wt/7IRI2fEw/qkGf89CeUyOjZIGoeE
NjcvaoMXoHkWfyFQvB3vQKfitklB5fiGTLnVM5DCf0qdfhgOnnRZam+SfY/oKkc1
dJXBZkNpG3KtZYj3nDSAqEMJLWPno/lUoD70o+tFF6tXhOFI7tomtM3cD4Vt1rms
Q+ahVd6U0XNpksLcYqPDE6hI+mL4TI6zlRNUejaAJL3XsUSziNZJ25EEQo8pptL0
CEtuMdgCVOvb0wWio0HD5pFmsiVO7mnwNI/wtE0k2wpOOLh0eHCzNdm7w7aENt4w
yuXBvvdokZ5H3Cu8tLJiPmL8VeCHwJW/kJFKoYZzM1MLO1SNt0Q8XdfcWdGK4iqO
9lgGt7UDvuMGKDGhTFFabdPyX6utlisl9XlangGZBXD7QonY7fdQpwQiPr3GzW9a
kHRGvHKAdM5JQcj5lda/KNv0i0+RlNsQC9Sg0OJ2Y9Wa0B/4lMtoNzd7Ozs1Cd7l
obvL0fDoyEjLJUbbADQa+P486lzqZgJMyhOStfMMUNisnOuBhbpa4qRHQGVsdW77
6qmFtYEUWHSl9ZLBOvuGbkudl52BXlKVpT8VW3jL2fUHNLrkkoX+PafABw0uXiVS
CrgFv9Vo/do0qVcJVPXGUW9kwzEF/nsynEMT7cT5F4Wscf4YUY8IrHeqaTLDLhcL
IZOnzPcnv2Y2MQoqV1YZ7eZrdecgCVEbK7whmkEhhOeF4yH2WBF4SXl/eP9QgzuM
tIxzfmTbuC4ovePGE3ZBnJgQQwD1v+p9zdZMnkFqHqFnhHxfj5tMKMeT1UFdxjYc
xwDqPKtdJyldZCiCDLqIw/KuNK3opw/TFT0j4gbcGYZiOtaAz9Oa9XJTsEsIEiBr
cX/Wc8O/LGIU9pQiZzfKhobULV1RUuxw5MI7KGV4YLi1gXJeOzRDFj+ol/WzlDwC
h+EUo1JlWzDMNDx/DM6JUqdEJv3711zrOBk2VlhyFWGIjesMECeTp/sUGS+SxA1E
ZBoj5z9ZBGpwxKuMp1m5MaIInllj/pj18amGS4exkLJpp1ACSyfoAMDhqSs79anq
LxBE7CAMkcjka5XRGTQiijYQLqWtIN6+bilubs4OLhUJq0WbNNMK7fiAX/7r2F3k
Lh+l47nfjl2vsn4cvQwWKr/DKGsNtdgjkHiVr6G1yRATQtpUG2KkeaWEzuXNK4Cy
rjlUVL9RVGIzWiaAldscsg6vuW71rk5FaOVluwkp/Hzokae7/oEQcqY2gxsVKxaZ
Oqairpclu75j9ZZe0PKjohIP1UatAywJbQrBwwWwA9cW+OdwPPTgKhSTKsem17Ns
Vtn+4wKZ/qXeBRZfv1F/3T9wlXsZKzCQ+S6K2l+NAzJF3cUcwoEY8sHnFeml7DGw
/4RSjZy/EmDcvL3g3KWhdzSC45ooh4iqdwoeqGJe6ZJY8tHKLmZMa0u1FjWp9Xqi
llw7Xj1aacSRJHgKCkugRMfTIAwllGfug6NPpybXOkWfaOm5fCDRIvBdw9xDk32d
j8n+eDbwVsGTL0NKdUI6TXKd8TyuVSwMoLxrBWnQs7y3Jg3e70gGRxPJRV1bWJPq
mJXb0Id1Yqn+ZBaUaKqlP5pNHdgFgqV9uCFpZNGkP0LuYb2yyK/SBAm/o14N5xNR
tB5HmE51PlocEHXwRZNqnF9ZqoZRTSLf3rOLlBTqGGBQZlOK94o5693dp2/lTTy4
6S8PtWDFj85MVDKIhZaxyd2OU/PPVkZm8ac1BhgmxF139G8F08dO9GiO0EZSWvpd
MYD+YOaYbHmCKKxi+XFVrs7UYbbCbgyJOexvXr7VxL6BF4xtjw5qjwOwKTOQ0CPb
Ylwi65L7Nz7iGYrWeJFp7Th8Etj6fEhdmShWUkPXujnf+MBGmTfB0ShYsXNqVtoP
Lfvk3BcHp+gPTqfh77lalHKxzI5EMMwRT4vKKUaSvggwjNtz4extT82PSPTi4s6+
INF74tuLkuqFMzq+xoBm7iOuA9mD7BKEEWPl9blik/N2vwSbPk/DuF21kJ/G582Z
Tls6lltwJVJogMT7ig0Y6gw+DtkaTLZeUJxku3QisFfA0WWUAjk/0W4kw51JLtj1
ZAT7Jhh5KKHsSpzv0Kt59l7IgRe9iCukwXYUumP6gzdFjayJGkUMBixuESMZxQHN
ua0NZ3bmQ+dA+rpNwnqt5wo9rwqw/D8/4xzscudeYjEpI81Kn3W+umwUSPNNsMYD
NRp5rhbGT51vWAVB4gm13mk7t8LF42LVbMwtEP8ATzxZ7xhMstsgdTdSHqO6IWEJ
nvoFa1/3WDOgDIYHwHOniRwb8tHROXLTl1DgEbWChDy89MeXv7ecje2DRIqEkxlf
0W+H6atRFPx0TPlUOGt4Ke/riTHTIUomEZYHpEU+G3TyHrZoPRehStS9UFujgkAH
aC5KJVfjRuaT7U49STdc1tnUBrcBqj79JA5LFLZbKsFKhQVISdeP7yJGxmMXEeBB
UWvinK+miWJTwnE/vOx5KKiIwxeSXnn2YzfrBkcHCdIRa+C2MB78eF96qS/zZsDF
nm4L7TyhzJIogsnfcEWqj3Kss//OT80HIYVEtoyImr9e7oZOAAW26I0fohc5eiR2
rNn2NABrotF68cxSwkqJEOmaGVmoqc67X0ocEej6dmJjafNSmRd11LMeTu8QOZnG
yQuM7+7pGvOO4prZP7VUdaCPy+Drz4/XbKYtekqNhmnX4gRkUX3sLtpC0JSO5tCs
WJP42jGxWJpYQ8DpT5S6tgJcHcqy+ng+8a3+JRBBgqFd/P9zC7j7BClLze7h+VEn
IWweN/LBzxh/Cl6nmVUT8NDU9bkOosN4igLwbdryCwcflMgtnCv0hvkuvfWzVdO1
af+dVMRqhHnBcGMAj49SG8vHlxd6luDoNSgURj44wfyW3fU7sMtPiw33NKeCHzyt
8qt4o6ynN/VFZvk9/3BaAPgZaBBbXn8wdUiEGaX1nrSG9Te0EaE+Bo3l0WpRLD2M
3D5UT6+5vS8ufgHLgrTnnsrmSv1gS8KE2ONj+H/FhO3ty3QazGbo6zBcoFlmypR+
s6zjvtP+kyto1EXuR0z/a7TbJTFSdF8RhhSGw84M5NCCGG/yPP8+jWGHXG4B/69U
FzBapQFUi9HkUcRkuTPF/TN+PcHrTs1rsDN6o6EZjX/lCbVRx9Si2YqNWEJo/yE/
hshVz/zpF1cH0jFhhhHL8ByTk01YsjajkSP8C3o6xElNimTI5YNpZPuQ74F5qe1j
bjGUzdpKaL0KbIMw5BT2lZT9WzW546jTgvwHgnua3qsA7eHmGhXmhbdmznoyNZH6
Qc7lkRPBsjDQFK9Dba1Yo6EUsKezk5/8VRy87MyBs4XvGZJ04eaToUG5CLdcJk5E
Ay+rLsfWJ98U4TrA3+uO3sf3ebcuSaJJjy5WnS9oOHHyPm69wmFPItqJJ0ygHPfz
LDHeVYGJ4x5mftclljCPYKfdsGOnsnOfQtbSUPqxiN0Od9vfC7K01b4yQ9uL0i7m
4wM43Yn5bMGahPKxcjDtYBQmHmPdC+iPBhkP+KaDaTW4z3Lh5IqAXJ8ulF/xIBE+
zGy5yCSIS741Pm9v1mA6v8Ws/FgcNvgW9PGTNn66M4qxRhE1V4BJK4av3RR4lQ/H
n4FRUdZQ0xeTP+7C5+j3dyvH7HBkd+No94wNmQn5WoRTm5kK+q/ABIgD8a5YkDOb
NM0Jm6HKO+hC5dvRAhZ3KdZZL+ww/u3Kq2pixA3WPec6kuII6jq2nmGNhIKpogY/
JcirLgCmKo4B9G46wsFjhMRf62XXlwfFwonAfBtsMAlFE04UlPeqXZmaUHGQdNUT
vTb7Q/jwR+bJUdpTkylPACdPug/PeV21mjYRiRnUUo6NdzTFON7y6YURR4VNxW+c
CgPphdrtQ/L98HEU9iYKxD8BfS0gnSNGEEVoMhNBiaBEw0NhMGFrtu9RnmXS9nq4
00k63aO1+RFitPKYfxtrhBDvQ0l8YE65pyzU0N4gITxdQMf339dV2d4wbNpBoc9p
vrVsZSOSgut8rdRcqjZiVn/b1ZYhGKs29WfIzRSv9cS+z6mSWJB16bwO1hTnBUsF
snCM5ZHz8lJSVn6+oAUquua0R88OlXeb9inc5NfahtuJU6V+Cd9vnfnv8OUKaBbe
cM5tNoD0/Eq2KPrFd0CgquXLRG5um7jNHyj2ZfhVtzQBCfBU0vhjeIzumH5bCnfq
5P7I13eiBcGPISpCjN+nlEtVawsOY10EHBn5V2hnt5zKSIPwDZLAc2D1JHN5+gQT
iAUeqA/k9QKnJAjADU8e64BmhRWRdPd8bxJHyf1gdONvcoc4My7XkmqhtRDPUqem
0LQ65wMv7r2xKWwQHEa7e2uP8apBvPxK/C8z0k/5gdHfLe5wUOkPNZOCa3K2Md8W
H0nK1fcqC+l4F7NqlBw7AI8XlR+ZayAJ883PoyQtCYytD2I3qoAnfg4wNRZLZt8O
pH8G/KyHPF6RB1GlohJ6aQGoNDSl4J8dFiQJuz5kAEQXpRmEZtnmlHD53Aw8yb9d
c2Nqu08dROR3jO32qvp+EH4MEWgcMgahAC0SgJ1DOwIzaalBpZtGi5WQaErcTEzL
tWU7SRdl846OMBJ932CE5VVYha+fjR2Vo+N2AsCSpItQKlvNlTZ1OrKIDJPjkuW+
Sjuo5ChkF6ZKoe6DFm3BnmgmCKrOIMWU17vmATqJ0RnR8xeHfsYbFQuL+tL6hepz
QKRiXOdGHzJA+0SxT3NcZHN6P7jmL4njnwHjt1j8O7j9vyU2vXluFD2ThHLrFuse
NNz7AhJjRivTOaJCPirOC8pM41fNNted60Bl4CD0wFWBR4tceOIyMlO4l+gzx5cS
Wap9hCVTndYie2NsgmG2m4qx8EGLiCLKuGtiO23KD7tcU/q8LGlc0pDikQWhiv8w
YlzeZYanBDz8zfJIZDSJyJ++nm8v7H/UUku4MrpJVhDF5UWoJmH4evXHXRBIDGxx
rX5oqBglBro7XCXH7Vgvvcg6c0hOb9APS0fMivodIm2sGbQFqAZ81BM7zlrPZ5rN
+Li/L5LMvlaPlq2fAWGpOuRxGqc4TVIBtzTgi+Z6WPcoBmEYO0yBU8BjQmNHrwtS
uqmW9shGlr+MBtYPT034suM2UHXzuCDHCfCcNL1LEtZLrMc5h9zu6TO5RLguj2gc
HaDz4Qp4PHdxCHzruWUlqetwage8pOSx9U7OJbUQWlqydlh6+zYUPDjZrFOWJzxy
l5z/NWNxPqTPA2d3I+1PgoQHvaOgz+TJ3CH/XihYahMelja50UVOwh2LarNq0wvR
NUIz5xv4LOPqi2fhkduhUeMPCBYfaFy6dKvVwsS47GZo4KhI0wprsTfXYEN6LflK
qJtQJTI2Xqt1F0uLHoq+Dy9GBtV2/WcrPpJmCo23/yFDilvaY1LMWdn8DSJCIHDZ
Rzs8SgEC24NKXOL8f4phMp6IMw9hL4Cs3EtqhdEUWd1u/9VpBttpVQcI9YTrtB+o
cdQQtwYT64LSjrY15bCg8U9T/ivfgkVfhWZnNuRthrsLbNFsqVk994lKI+JiJ5Qe
Aq0/C9sb2+58q9JlvLPeVhz16hXNhLVi8JSI/EFqGcM8T82W6T0TxTp11kkQl3iI
IYb48zOCSDTZW+Ux1AK99US8o0Jf+entrysyfN/yKn1HHUVK6acG1fY4J7gJJxbv
Oh+bwv+F8lMc2XHsl6LWVh8hPrW0AnH8hs/R9cytC5WIPcDCT8hZwWXr8AWPozVU
mXyD986NWRYeIbnQdq8GGxIXrjzgLzHGXGdpULITJHBUCJAG88KgbmfyJDpGDe5Z
5FiyrHjIAiFj7wxAr71UHJ/7Ib3tv+fPXmwcLYk4/PYx34P3PMXgPvej3oaaX8Xt
sGqJaMrqf7jrOWCAw+NPvnuHhy8S1j0ujF6udSk+BTB9IEBbAtJuW26f58RvuOcg
+9w3bJ57GKQKqS0J0gpJ2VkakWPPui1073RNk+krv6s3xXCTdijEKEPgEIkEX7pN
IJHHYv1AqfylS186DXVIBBYo8UvKOCAFwmLSwQ8LHE703chmPfTB9P5Sz7u/BEz6
lhFN5zw4KbJR39K/WB02R/8rxjmTXYQYGOnDabC5prWZKJbDIBDwittYG7HUudtJ
2DfZh3B7bB54jXMj0mEL7gnp5HWJ1CoFCQCeNhIiTqOwLmetnLj7GNzWvaYzZF/m
IC6CNA1fUBX3gYLxruNbMIDobF3Bzt5IITPTD8PiMdeRQX94/mqn8pq6/kLn3Uw5
g3X/mAmAvcD9ZBpOBYyTNgUWq1jUvYWmlvM3GSNjGXN2safVv2zPXMD9JBpFl2X4
uNWhjf/2GuhtlQUNSneki/l13Mru4p9bkujOBKhMzxJIDh220TjHZ4BnGS072hF9
rFJ78rYaadvPCJVIHUAOOGxyCvH1rQDI8xiAEBLy3j3ILdiAJ8wQAbu31DmOmZu3
PKLR/DBL7WSzLVfppjBAT/20dPDRhDcBf8Te1jhowZPTlFq5yUQfdHUzl9o59wxb
2bSqgqmtJPk2ipoch8t4zATiWDxY+hbj9l5FhdMS3XgcM9BVna2WMgjKMzdjVku/
6azXV6IFxX6eUeyS0Ofl0QFiNPI6F4LWtzMM2Qto1GyYEkUSNC//wIDet0v+96u6
weco3hpi5Ln93sZ4tfbZofMij9xALqlWpsTr4mQ0h+6ga66Q0CC2YS9jsqK1mJ5p
jHn7yS3hzCwhzkqLu7p6L1CPOw7VMAJzpBTTn0yswp0AKOIHOAMJXYnjmFc9krmX
OdeRW/HnAQt5eJla5epFBbAvIe0mhA//p06oKHwZehXi6A7bvqjuphlYeORcvLGL
51X75gXAC8nCsenjXPb4IRfT7TNDiQ9AsY7AVeP2oVHudIDWJiTWDDAjGC/c+Y4D
97weQXXl8NJ5VHg0xhDjgTc/ZcReE9hmvfpAC1siedEj5JnxCsWTIQAiOOPi2CAk
mdF5OSpjqFcEckCPXdSPJC6TqD4j/KwX+R88+UB03ii5DfKHio4yWTi2a9Fbma26
DETwDfO5SyDAc/wsJJ3Yqr/kDQB3VtTfM4lgWTLc49fLXtbMUY0t9q+s7fB3CiYp
mg61eKLH/4X7yFPIMUWawRW2cRFr4ZcwG4xbf2S1oXKjhzs2vvpW1MijpMLuh7N+
oECe/FmYQthHKGzzuWaCL1qjA3TDgBVk0tlaXFScJRcL8pcIDX7oEMoDLDLfMfqc
ukE9wo2aJVkTvZrxrEZ8cg7HRf9pj8XH9TcxkqWrw3WeZo4xuF0JWMVZLi0p0SEz
JCMYrQ7IaPWTvptPH+4iuyCmoeozFsYxeltDVI+1pNvQx3lbSJGIhBTm/5WNfule
wuDMpgPp3C1KCFaiMBFOXLO4l+SH5ejzp27HzSZQ/T2MCr4c0in37dNaPy6rL1jb
7E5s1oJyidcakgZcRIEAnMsN3k6rzkDvVcbGL048wT6+oMD7duxW0PiCDfO9qfjT
9pb9NGjbcFdicISXZMCG6WiQrtS/b6jBh2WMqV8r1cK/jamrnYZYXlXPeBZ8vu58
LfDFulre+ltHkkROzxrC9njakLH6h5+frSnFHzRteg+z6n5fJoQzd0nOsMRaQU2F
zRGCiZv0U+xorVBHGgZPBLIQCUt3kX13fHdxVNMAeihLNLcGsCAUxcvDX4tSMrcL
wqCyoKPfT7nY6+IUQ65nzDL9SA82fKDeOOW6RRMAEIUUuaij91RwiAOb47Z/CbmB
acvJO2JhVZsn5SSJL9lw3dWnFrTLo1cmKBKRXcdZVFtE7P80c7E9pmKwWzmPyA5n
zqrlzMfSPK+9Poawpq1kC1D2SB95I8iLSzG94zsCPhG0Vnd4uqcKFi959ZAWOv+y
2Be2LGomTw9Ynz4ssENa8+uBBWNnIQamwwIX3bBtKgjAHE+qocVJvhMFvDHPTn/0
5Mn/X5Yo8HYm7uWeAJ6vjKtNhLUSTouD/TkK8WG00mCEhdP6BOqKx/vsETpaKce7
osG70amAOqDZ1od37kGXSoJVE5Sl4kz1siKU7SP27OF4g5eINmWj9yZsNiusjioB
qaxwe5VnCw8nb8ORfo3aTADFOzMxys4bgOhDzPS/VNtWfmCknefq/MwKQK46XlUc
/30vM7UprwXIKO/OdREnB3Dqn193ICFXGSZy3FojhFUxlUVhBuUXkMQJkXpKlZ8P
0e5XBr252P7+FkYyo8vlwtBeXqfZCQCmhRDAmt3qxx5jVEvWybIzRCmyzPWpMiQy
ARYTdhNk6U/6JUQaki+x1L5qrJbcWZETlwn2+oSwecsEpzifagRASYNIVuPzXPIb
Q2+mlVCC2aEhbHzKVag5yfafh3Hl4erNdLh60GVKw4j0xvFs3E9BWZEWelCmZZqe
wY2t9bWxvVm0t1EF85gDSce+yqNk5wh+QhXZQ+LNAohD9fOUYz1nYbrWAVLgf1Fo
jEvSNM0Ialp5GJ5CAtgPfZZ9S9WFtYW3iQf/AIS8dDXefGRY7Yv1vFKDskGg+3TT
yg+A4LNhXkOg7+EEEmczy1xrsZPQTHVxE5+H/PSV6BPU835iC9e3KQMCC6rGzEss
9H4trlsZj2tS8UB0n9rXZ/DufNE3fEFRWtkRyZzsTLPijj2/hZjQbPePAto1olzD
wrW0CGRc40u8LKfDrkd6R2BTfXrTWejkAaBWFAKb0NR1ruVb/5vxHbzbmyrVYg/C
xIy2MAFKAe2QVvMnT8iv9DgcuTifaiSE6y0hl8Aaavl4UBQjznmKLAO5EIL9KjLg
mNg7Wja02hTgBzM66hoM9Wl18LiJmsJjgdZFs5kHKCY1UcmufxYhJQucfKhFDRsE
TISj2NsG4qNWJw7IHKWyhgur/I36sMCsH4JOl/QPBDEGxrMgFk19ijIst3GRKbuP
aCB8C6zA1iVcab8U6+qgFbHXG/z72gf3NSc3b4WcD15t2gw2a89KXbRTqFv9gYGj
ZZlIEpdUGxMPxooSnp3AvQYeB0CLMmHVro9wnzJEQRt1Xoe/FXoylW0nue1MbHRg
czupTkG7oeGt8TiB19X1xNXPworMtc6GMshO/3NyLzYNbi7KlefCn3ZmdZW8+JDe
E8af/q2UHG86gIOj28kliGcbjRgKV3O47CoqTmeZ0m7iqiSLiUNd/ZummrNvwAE8
U2xa4uFiMeQfRXUPOHMe4RNnFvNr4S3aTo72wV27AMNrcJO6ed4kDpil/Y3ifvcI
0U2h3njyt3WQv/TGK0S5D+vpQqKXQIa4ATaHtCa38Wr3Qvmlpygp4hv3BCIia28Y
UN6DExMIIDHp58DH8ll+qkSBhVxsiAPMJaDVPsDh6QeM2Id7gqtryFRmJI4wSgCF
Q+VtqFJM+vwwvdE9psNqfTfD5cUA+HrT0EZQltL33nJUWecw+n3ONzJxDnDIOQ07
lTGaRc9yWso3aoqeF8R2E+U2keBnxS1M8ciiFf8VVzGlriiA8R1+8ma5B3X+wJ0+
/m5itFKQfwlphffRBGKmGx//Gg1jW2EdN2wVMb0YCOWDnaFnkclQQ2D0q0VGsyyB
1R+dfRwtE9bljAx1YLN1+CfUD7t10VzW/g0gf+vIpCw1//YT5jFPRRJ79zm6cLCh
WOreoqEnP6NFXJai2lY2+Otoj1yCTsGhtKRQcSoy+FUGLz/SyDFCEgkzwyuYcNol
NCufYhUQuX/llchQ3CPZWemVKhzx9Zzr+6kaoCB9qMq3vgiMn2DVlOqoth1/xfTX
HvmTKoyDv7lmQlJRP9coKyTgfUPhWfLUS0YSN6AK72HlEZHag1F+AKWHKX9Hcpbc
jvIU/yN+EV0Otp5Vy6V8m7hPSy0euEi3eRGP9UfbH0q5H1o2KWgOTfGON22yBWQL
e0XM8rPR6eBgTPyZ/g+Jy5bfjrivgxOEtgOQQWQkvZ+vOrqdBCQhpFzCdHrR/t14
++YkUAuBS403HDgTqANw5vJFcsQretPxiHzWmWhxXz9NjqiTUYCeWQA4KKeg4mso
1ww2Kwq0tiPd7bKEm0M1C6vQMYHSS7wjN0EXIhbtLDp95Hc/jB/CvRqhAPw70m7f
7DjHH4/2dMarH7/OEr6avv7kU+xdKRhKlHOBTLp8gf2EdZZPd3QjP+Ka+ZcoETgu
Ug66aQ7ImS8XwkaqSuw8ydybZjmk8ISqffb+12CzZlqnXhoC7IsbSApl2eTd8Ax6
YhcEUIqwtH12mUkg9rVHRhZqMR+G++E60Wyb9t1V358isnYLwVLHBOHs/RQmWyVO
2+2t4NalvOXxTa40W8EtzjTUNsPNObpPhAhDSGjX5Q/6wCrZaHMwP780+m0aUqez
IfssJvWp9zqCg17IuP6NioaraMMbGePLRrOU8ej0+x7RBpjlspGQz0UiIBIn8SAt
x7HLyWhkgAbYnWnhS1RuSykL4yWOdD22ucCwRAxNSK7ldRrp0/ihVvIwzZMaHYWQ
YJbauiZPN0LXdGiiuioxiYsC27XLvHr7mk38B+1gjTH4f+cXjz++vZN9yihNH5h3
JKOEgBkKyEgxew+lgm7434zbGG2nvGjioudWLDsKy1cew8YKjqp6bdW1DYGQYkme
bOi5QTnNRwfCvG4cT3fw2W2wQT/PCEhhG+AobSP9eONCbwG8ABkmBFKGsyrsLy+I
VKeHWbGmU7Opg7Ms4WYf5SCjB+Qqy7a1IQfY22b8bTHmeuDWhniW09zW6EhC27cs
VF5YLgHoGrEssIVrNVPMXOo1xzdqyqzrFlD6np/J0EP0eFGtB4uo8l/2cydUJEOK
IECRFyC+zUxhNdWpKAuuEloFydLaHgCLQ1PDcH3eZ+f5pwLX2UlXaZHq3kXd+WVS
OX+JBTBV9ADLwqnC6RrMckcgV79jCjApgqRZx3FHMPQRqFOShPsmMBQatYXK+8YX
zfVAhzhEFHCTXb8byUHfP1lClgD6ERY0LndwBmjefX9xmBO/JJUNtoZv8/Cizk7+
1gSL+S/2MgaFBRWLky2Z4PopwTkRKv9uWQIAHDtRdoj7QI9tRZiybhYYYlnFIEVI
fZQ7hb73CRWEJ0sSQT/yuvt5ITR2EqZFRV+FLze4MLi5yI1WxeRNi+K9uI6KSxhY
emJgGSobdmE476xAtBLomNTsEmvH0RAcp7NJ5kQadRLWY7ObQz/1u35PsFq7sz87
pGh2UE3HqPMRZoX9qasfGLx1YGasVdXTx6WHywpb8YKPGttVAH7jZ4YFaEDjHLgV
FJ2SxLuOk55wG0Pvbq2P9/9HssksS9vmFhtdzQiyxEi/dPrfWP1EdB8wQ4ub3Zen
2FG5nLfts9bZXdmWwkQOZTojoc30x0cpO4QVFOBjzdsUNQRo1Z4G1YoPZuJzOcd+
GjRqtgNdW+UM5UD6wnqlv0eGi2lm+L9DUCfvyQvrC+iPnPWz1dhhiDDeKvjSe1P1
me5+Jz6XRYfCARG6KrwmFwNvJIlE9hVoiRMh4gBKdopQQ4PDGdXJCn4voSlRDwL2
BJPCbG+XBd3etLzrJmZzs9BKkciCqV7IkWOv47dXTsHFzSPniO2d01MejLG3GqmF
AdFr+ipKHIVOgfYbNCKWTGfJltu0r2Zri0eAN70lzzwICnfMy/yZVjEaeaDjVvI1
tiybkIJbuLeamFbWvjBsu5tnCwUzyjDk4EbpHnVQQxDUFCg0fMw0dL/VQPO30h+U
CjMkL4ahLNZVywqe31RB7wOSKkSx4kbIe54sfDRsPL0TxMFWEpJ3L8t7JJ6bERrW
9Q4bFu8eB8l3tYJSkeTVyqF9AcojURdO0zqGhIMS8TBO67Tp8h8egggo3HOuhl3c
p98JhdrbR/vEAL4Ya8M8ydnrnhSesrVuFQt022Rxu8VO4HNCRZx1iocHxcEeB5sy
CXRtGJN/+H5/8wp25mpzysud6YKD3J/KESQa7mzgvarYXRc7UDE8gtoJRPT+89Vz
KsbU1piskiaFgVTDp05vxS+YvpGKRP/wLDBwa1T7Aeoa5BL+TOE7JglML3BPxNfT
hLSePOkPjZClJoWhkXhvGXCCaQSFB4gPcPNVqt/nP7tFc4gL2p4KGU2gjXAOxnlo
Ttd6k/Z7Gc0KFuhjRodZFj03lkkLv0DzGTekckgqpu4UlfJTQXH+HFqJXCoAGsMo
CKI7NvoVkfpUmtBS756+SSniXoxAzL7ewD/x290iJjJaU+YwaGROp6ovRUTa/4zD
GX88zNYB8kX6TbGPv8bCK2cvSMIhVjE3oMTJtXczg9Qj+CbBs0ulsH0xtuDADff/
12tZvwq8eB9CVG4yBfr+7kDEPGUFIb1eNoUJCgFXz69vfsQPUm7RrYoy1runpW3u
B7eKULCd6WA48YtXr51w5nMO7j5zYEr7LSJs5q+k2f33jJ2zNSmCedu0CbpRdPus
AVsorkWHeT40/iHTpNwELJN3YA8rWa4JvGzG7m602I/Que3BY2P1iRCgD1i7g/0U
14AnGQtd76deW79U28HV7g9agiF3T7kRjb2FAG0P47K/ihyJrMiJUFkhXwvfphSQ
vQws6KGAfOzVPrvM7NePEBuWBCLgAd2u9GUiSY59pZq8npnufm+QfLQxujn7BU9o
1omxZyRXCTsilM47JSIokT7Mah1BPEX89UHqrN1KXCVy/b/sI1hOoMLOpvsPhw4D
sEO1P/2Eg907pAaqRrThJKx6CVdIpYD+P9vxgcO/ZCAfd4wQZlDTaq6D8oHOCeJi
FqPvWLYuD8YsVtbJZrYEoOgYW8USayK8nMWKkgB8U97/rYdeiYwRkoconOqnrPQl
vuqhPMg993aREqXGZRtE4Eh3qERg5OCxKeUBWszjYvelHRxvMctwNnosZmJpVZHz
GkpEbm9+h4bBQsrgjnDDwreXg9gMX0k+pi9itECzeoboRg5J69WeultUZGfOv09l
QGhB9nw8uylW01ja7zlAu4rYeOTcYaNNQxbhus44186hjtrlNHnQSFdjBcKG53vm
xLRoU5RczcJ7sSfb5IJ08zj06JAV8sd1s/7T+k7TpNOYs5W7AdMrWowJyERpv47n
rDIFQTZPQ0nEMro6yNbzv0FFD/mclvrB6sEn1kRp+/7Fd/n1KVRlhYCd9IVNsOmf
cr+rYSMKIO1/piasohD+8uXxckmseGEazA3nVEzg5wLvfD/tAm+IAR8+pTHZIjhY
7Gfn+Z1ORjeqxmy8V5rkv5c/+AkkDUJD7ejMM1u8Z7mVMhgE1+ToZoITWBgXbrNm
zBPEjL3z05/7v9326tKVURqD6gydzi2amfKbhYytXxe8AqOZupWI3AhAFVUbXYK+
pG0q+4bQ3zriSVJSksmBBZA94vs7jGp1vBQkbpN4cGS93n5Qot1C9ewfL9AsUWvp
ay5drRP+qdM7X7y4xX0dKzhTU2xa0jGZAps+THAaHWi0C/XS2q88kh6XRg7FYxis
u65NtP7zbJukVdwcI/CCvjVWuLd0KU4YyTHpKqhXC6eiiDpLth+53no79tKMo6Qq
/gmauzviRrt1/UOrT8fB6hqvmp+Ick15+AupZoGUmMJFmIIBKm3uD9dunR0QJcDU
8NeIyzHBYJjg9rQM5vWktFO5V3zs/pgPxXHHmBPXAiKibUMpyCKGaQ3spiq3JDMn
qrjAqYC+Gtp8oDowBVI69dVKPBAgtuQMtBKGu5RMW6xZpKcB0Nh9LZj2aznwp9gP
fWnWt+9HNTPw9YmE3FjN1qYdgdMnvC26yYBOr0abITTs3lIzqboyOikAl8bU8+vu
1soq09oa3ae8adCjTrzkm36AFEmD6lm/d/vr1aj89H5dzO8fqKds545G3aCpkGy7
QyDA2xbsmdiHfiaiggQ1i9KGayFsldsPMjS1mZxbG0UqQXKgO0ZCFsuDvqRFHlB9
A0yOiPH330tD53uQRCDnW9TNNOEAt197LAwgtDqXsfeNdwQvBqArWjEcpM2D+RO6
S/Jkg//Hqf5rBccHBdDa+F39rzkENDMILNI5x0Tx8R0VJsJ8ouAY3UEVxpCDUulb
6PD0viX/4AynHdoh09FyI4SZQ7Ig+UJZIV3sn9nc5K2IpcdrGPlWJuOBM8XGq/th
+uQPVuVtRHoFOEF4pZs8a6SNqq6ffs+ZIIEYHu/gejlg63kgDASWVRylggDaJY0b
gqsHnHw5HqVC8NDcH45GXfSL/pHEqAFDytVPHcGRVjn2POw1uE0k/KjGgH5eUByW
7gKVJ6+HDFkP2+Stb4pBjnhUcODh8p8FbKr3SpYck+ylehdI2c6r9wnTVIm6sHzQ
gp1YoRFMK8KJ7iFUlAPZRAARys9WRQs49SOTsfUurzqtwViqknlpFulTjZxK+/eF
JxcwzHeSlLixSn/pPC3Dfev/DxFIDPDEVhWhoDcmMVJ4e5vE6XKmHmDp/vwTv0Ou
dnENKPm5WnF0E2SlD8/qbWG050iKvVJERPv8ZjVatYsWR6JjMtmSvRagDpsK6IxV
6BTCdZAABocDO+Zqt0T7bDwR4UBvg0pJvJHhdCoiMMVU7fzJXxqgGeBDtjaexbuY
big94l/rqrUteticQUKR5bssekVVaWFmsan5aiR1kA92cshzE9R9vVCBWkBsUUuc
aLxtWltDmjoeq/I40p0CLrk0uKWYlZWTN4X5YuYcEY1y2Xn8DSjXbzEEjaVV0w2G
h2DMmNCt4yGNE2LIfrzih2OWkDnZlbvKfgO35ohEj+hamUoo/+KoUv4sDT1BKW0J
yHeIsmPcSr62SNT/jGpKzHTyg/5u/r1jUv/ulZ+fgaJXCvvjJob5xV/Exmp5shaq
byeU4RsPh7oXm8pH1Cji9nfiKWVb45l4zh2FYvreONZLjsVKQ2wiw7S363T/Co2E
asalYcul3hyX7M+dhwymfIR1pROqpZJCaHJc3spCDT3UuASYTA2WfWSnn/IucrZA
wQclwVBQxHUdv9ONobIPPvSf/LKSUeOO6L+WAQJHvxNTSDS5+1O3dmBBxBH0gC9D
d3ZLJgIoRn2qIg6iij+/MjOy3iE3ZUtU61pjuXS+4RSQqbKdg91OvyyiiO61j8vh
gum/X/YpnpPu3BHHlrv/OEQ27EicjJ+vMzNEzgMb5epKfux3oACZiyMG2bPlubH7
UGA6AKLRUSQFh4Op5P+GBdEzsZbuXCpSxa65jEvRXSJBIDBiemUm2c5Ctpcl8mMA
LOCYfQjCzb4nIFI2HRm5AuPznEvEChxvi76Dez6oWpDPcTiNPNkl7+4FfOmJ32Ba
Auz5meICWimWQ20/IYT+R3EANbUx+aU3HF5PSy4FFJSwwfLgi1uTWSvdezjAmY9t
FmIuTjAVMHYB77SSHBOoABgfAPr/h5fBGv1pDOlRJVJ/IEZBBkPi4R4LQiSffyKF
8k2gYJckZ/Lbs25zAHnJt26v0zopkSxV/l0eEJ5Qn11nd1n1s6uMJjo468r8NHO4
jDOkoC2FVgWcIBV9kdTQC18N7ryR8yS9QeCzY9kW+tdl+oiwxvf8yPikqMzkvFmV
mv5xJEVneS8KLBs1WxVXyw7/oQ1w4YognoovzRLzUfKodnJJ6nojsuuaMpz3BRIS
k6iznVVfzDDYaHUALKeicgYdoZFfHPh89ZNu9JacUn3flN3kxq7sZlWYVhaerN2v
KspLEBgOWD79JiWJR5jrHXcL7kmaRJxu2Ln5gbmiAp7SV1oVVWEqNQeCz7CYqtyO
MRMm6HMaY2jS8kFESTGgevjQUtQB7PIk1f23A42aDwxD1jvPLgk4C8mPx/mdDMo+
fVcoPgaoH90nKMvbeIDOebX++LfPisXBv5tlx9qK4oAIgUscj2vMo7UHreD6xz6I
iuFC8HbN9pHhgJ4pO+K+jW65DrwnhI7iebNVQYim05TD6xk5fbA9HMEg71b7I3xq
9irEEWNWRpFTVnEKeHSqpWQQSTuCjPlW2yl2h6m3axaTwj8jzis8h+mjm7UATtGb
xNmvK9Eg0p78plmsS2GO+sVEn06/Y5idlLuh+6phdsHZ5t70BlbWLX0VrA+8dokx
RoosIONCvO67VJh2tIAPu9O99JPqf5zL/x94AbXeK4aM2MLq0GJsBD1SJl9Kb7zY
98jsIVzWN8RfUkmhPblk9KcP4FgCXxZKaAhCLFkueZgWHCRZ8MJa7zdBbIWL8Zne
R8NYoWuzSW3RwRWs5Sft5r9QHqIPp7gV8Ks5jlrnNVvqypcYUQDOjl0oie0YlGLx
zAzR+l3Ulc0zW/5u1A8imycFEX3r+B1GMXBIl/c3DMUnRVOo2jeCi5MivigwVRhK
LOnVQiEnSVLQ+khQ9IOa4lK2vfGsEq6sZkeMI1qF9RRjYCch5mLeFzouOCvkBqg6
IZecLkaW1lhBt0cpZkEYLja10rDPQywpsMAZtaxtVTC19fUL3Y7wlWgd1OOXJQgu
hfWYqn1xyM+rlCGJdSTgKRgOI/CZOzq3FJgXC0xQ0dAeDnkIjNrFoXiKk22OXP+M
fTkVOBeCJYhYStpGvb50xjpa5bgvf65lao8qF+9HclYCVuukXbRGtJEORqKCSE2f
AupSi+BDxHezrffuEGz7SN3HP/XUp/jZs4EGrdHIue7m4VQaeW3M8bCgnBx8tNjL
pvYCgoNLSDavFuiQzC1wcHpW2YS2ukrjJMpAKeXrFPx/S9IWmF/ojCNvYJd7XyqE
LqlmaVE0oC7/EpZLVcjbWRryWMCDqQ3gXuIt/Xzovoik7lwByDeufNKk2obDyE/N
bL0fPWvKuIzgbNp+LP2WVcM/SGrQlULByCbN9UWA9Gj332y3E2ZjH2uRJCPvItWz
Uxa3nMQCpdxF0WyazPxNkEi6OlUvtmxJ6HnUMNSfNIUfZdpW1T7LMoufPYDkGlcp
YWEd18brcSMTYAZJlkfN+tPbTHI3Eq5TQppA3Z8AGVwL93/1m2TX/obFo3Fuso9p
E9rxpL5O62Zf1/BWwz0+++kkqCUYbDzek+MKg+gi6JVOQUY7+4tj4qMNPOUGGGfb
xNg3XgV+ZlFQSvmoYt/aeUEmHAN7pcycVwWma4l+8/pPYVogdcjSO2tF5/HFpPyH
6iAI5K5MgMDbDeEOU/ivgYL0ap0vV2ouALUliDY8S8CCc7S0n1nNMkW1ILaXW+TJ
0q6UGkwZ67n6XlU3n1xRPr6kLsgyGw49JoSAtsfffSn/hsQ0NkNv5hRn9OzPizNu
cSN9vobOb2PdBOy4ZnTcY+JeC5+M8nf8moeb9n+yORv0PyOzTgPK3vc0nn73pqjV
2o80vU1mx7IY/Ksz/9Dda+mZcY+U+owFtdr87cZAGqDg0jaooDewZnrr05yzbXDL
Aj+Jn6d8H9bzoNvICcn1PN8SMmftpUXElaPawBP124/wscGK5qC76Ur6jQtGbf9D
GIosE/9e97Y0NQwf0f9Qq5/ky9dqut+Iwlfpor216QPO9oKdS5YPlcor9dRK681X
Vcdj3tFFYIhF9YXStKp4E+Lr2Z3bJ6ngriKRN5z0GgLt3ISxztdfuveoWRG/LtRt
KZHa+6t7wzuFl4wBccrRhGG+5chYqN2QU7KjPWEajr9hjKCvPCkdqIcmAoqbSdEx
IldUW1CHuaN98kKBon+/tTaE3SXmBJpFvp5MWue7Pb+Lp9C6DRaQx0C+8pDy9pYx
5g4V15y6Pk+siuuom4fY5hkHIjRjHfh4NtxquYfD62jmF7rA/m0Bp77Uxhk8lK4/
K+xFFo4jsI2CxHmP0KhlEefF0tbW5iEK8Os0NHXcNjuDD+u3aK2lbTR2t1wRN9sA
Oeuw6uS+eyJO8vSDcGpxT3Y/kcfgcew+STGxaIZmiwkheqhf/78cOsGatsviaUqY
uPP2oO1nOncXQSIfBcQqaPYR7AmGt64Pbsu33dGcS8+e3YmVVsKI310L0CrbgXY8
YF1gPakCU8lALWgKGlFZ0cNvT1MZp+jHh+GMUJcGIPeYzbMJMLleoh4Y6vKNiG1m
v8TbtMCt1eTMj9TNfszZoujrEtEkpLdGj50g7oiRfzgEWOJhU359k6oOYWVIBXhu
F8qKgYUOqRxj07wBblRrf4lvSdMwWZVyY+1I6udVOu7+xicxS3JrQkN45wsYsu8S
i1NKRu4EmhCpTF9V1FDeXDJi1R+lZ0LQMTMuPxwdLMt/n86m6Tdu908X0MSNntHg
8HHgDaMk4MmiZ2F6pPNNtqHErXuk/JvQ4TiH92e5OzHCMvmHrl5/3biXH/a+bOHx
q3Kf7XF4Uy0k3icdjfcEKqs99qiDfjR+N+0lB+S0tgEjdKJKvp8jOUt+9mik5cr2
6BJEwIBLD221QSET0Bsw5S7Rz6JAlESj+KfIfUj/vjz1x/NWtt9faL/FCIN9xnyp
qhHI1OyaTn428D4KuXZXNzRaIV+tBsOHk0yHmozcFcGFkLWwoMPhf+1eOqdgIN1Q
sJ1M0zzpg/wif5t/VqyiD/DbHsfJ0n//48BlEj0/E4I891xKt+xavxHWUqj9Wm41
aET56zsoSdA9cwcLn+OsWwHGMg4HxQvtP54/EIUyOA/u1hf0qe1HU5yNz+Vvh+eu
wRokI6k3cNUdjb7r7aVqalz3mF9I2oqdChKUyvOWGLWocReMsJmlWmVEhavMgtMF
rQ/ecgOhjAcWiD7PRRQB063zv28HCFshUAwI2n4EgYOAi15xZ+YfQwNKQ3QChSWn
/MYHrPO+KLmtuJteJyu765iF0dYpO0TavGypPp89AabgfGgKaZrDKHFURHLhlWVJ
0kGR0hzKjm99VPz+YjhOoAoyPaRvGmod6zPkKq3oMxKAdhE8gFweAkkXlcnzhcnS
hPJvsFAS2/lG83HSAiZQtgzIdFoYOgZwnVx8B35yUVQcwb0frJbURQVi9prGHF+a
w7Eoa6aq4mlijr8SLsnt+s/5wMIpl1Vxu3q7I2tE5BgXWLBWcOt+KgVBgamBECw6
6kBlWv3OJz+meW/lJsUpJy4sj1VYZFur+cn5m9vBANwtefJ3BCRLYJlylKeRsTVo
CzfZEOXATrAEiptdeDLxxPS9Id+eloldtL6bSCrXCbUbI8Dr3DqtMs6XKxPux4pu
PMeSvw2kppPyq50qOVIyvUOEC9oBtgsRXBmDX10wHEfliEp67J5te0eWrZ/hdWUz
JlA7lz0L+lFOxSGeW57Xo/ySqqy3PX66oxxSL1pzWnUr0Ppgwkmou/BDKxKey2oc
n6vR7tVKMj3k9hSs59l8GHbl6zpYXmFIvn+arvJou0bvb2v+sUaJQjbGzVa+hz4x
y/4R5L7J3uMYYyQ9unuO8EzbXT7nK1JbBEQkUIrtRsh8O3w1IwM1ed7TvsnmOJX1
5Inp1vgw92h+PC1IepmYRJhT+x+7fDeVzWRdugFEUD4UHLVso1XI12+ClvpONILA
ZP9NMEI6g0LqGmiwV1MC5q64BL82ujJwvbnMw/edoCzIwcnqj48vAwg1Agke0DmD
Af/dV06mEREJtooHWFWL0Wb5su4vCrdsXcdz9cU/jdV7uWEQwnAzCN4uFu6XIgJG
GSFlOj9DkXMPkCFPZev6kRXwJ8/d+4k+RKyJ7Z50aX/JiPDhXJOfyytBhnqPrmWC
TaziQpFU6l3BxCeSDuRkhMEvT1AdS2SLiqEyqAQWjkX5j/jYROgXkPA7O20Yg/yK
tQDPHSp16zivmamR/I69T3EaxM4O+FnsTcVwp+agkpo8ab50U+rjNJiVFps+kBO5
ouXqbNYKQHVoCWrbLiS1h0EOXybFI2zYduKqXqjoJt+6ughcbpkhgWIbfTvGQmzR
DlyeUecpVh5gkUjBIWixWpk3SKxHhvaB9pymT+7MgvaM4s6zdSd/46ddD4h2l1yU
y2g5yS1DW/YeTj9MIIMWdeinUr6MwGn1asSyrL8N6Sb3OAUo1+4MgfkKVUlUiTOq
WBBE6IL+r28wjgwQrgIIB/wxQGoCPOHYzc3sZYP/R+7GoXRgoOAYBvFbtclq4H2c
4Srz4f/sVQdpzBxHUsXt0C8bYDSGvBy+xqsfCHpJfzjaZt37CYTzZgoRIenSmMA+
eG9BBrNoA4HhgBYEZkGhJXHx0pLArNXKBGASwRPZ+DBA0G+6v+HwIXppBEhxtmR8
T812uoO8v8qCXfJ+KZSNjED53iLAFrSjXGyqnworhRsy+hAjbI+79QuFEhLGX+Bg
zfBbYCSJ5zLOS/t7yDn61d5GV8bIanTQQC2u5pQrf45NVqPloyg5gA5FDNwBlqeQ
fk/mVymOKu/TuBfEk5efMmwzxxwoxABf35K7A4pZYQ1Xs1sEG4hAYKNBtVjqDLNj
UfUuMUoQCTY3ZxDs9TruMtlNMwVHvY30832bdtShxGa25o5O35p/E2UeyMwxt69l
vHIl0U8V/m7+A+ToZe6bcxqRO8SxG2dN4Szfuc7L6x1/OZTdTd6zqjCOUR4dDbCC
99albKRGcl3ddFHxrVS6jbjKtL66JOaFARZhwYxcKoZAloz1OwhYGSWGAGj93Ad9
brmu0YGyiC3Q7zqnLGx0pnkCgS2zmqlmXaJEuTEPU5vHAoKSEDolj3+oxReb26Ru
4kmML/PePilFwxI2NTHEyYFpNovtr3JOu1BrSNzoeomDhu4XKBgAqEbtBJgL/bpy
gHeqpfWWi2LdMINssOpTKB5TUPDRTU/ASbtcafdomLB5tp8JLA4IJHAUJOke0K5D
wnaA1Hv7sZ+VF1M62+f0SOGPwHSr5bhMBuweLQFOgvM1+e9F+sCHiNluhtxG3aX1
QidTSXZXdXidIJ0IQUYXkA+mzHSZoscya+289v3MlrQTdIQVUJGu34LK+2Ol02PQ
WPqy76eyS/m50V0j8F8JGCtk3kpcsPkRf1ccaMzRyVDUWOJ7B65G8sar+gRP1W19
X7uLoepFa8afECacrrFXUyOwpj3AUpdC91bwoecR4/HN8O39E3UnAhf4BJSvs7Wy
olCQhTqrhVYTqM8D2sHkINHMAQCxltR1NDpJILEPY10BPjJ9zXh+4MV89eumK2IJ
xGrbaopZtH641F0epo+UXQLi1nm3NifEWJXhMrPIi0h8oAdF/nNStl9XBBrSuzM1
nmvmslFqvmryuqAVvsdWSstL3EVrWBSJLyCl922yEFALVDzPAr14isX1yzNI0GNX
FceYwX2Ca9iHfvpqOiirzSW9kEKT/rdkD0KhxPJxXZQwNTjRjLjC3Y3UXV1gH3jR
RSbBSzVy2ymbh8rY4RVHQaVqqGtGJYlp6zbpYDgfe4L1WLyn3nWK1Po6jwquO3Jl
TnbUglLpUR80ngsqxiC6EMvdzaZeW8Mvk0n3mM/qZmFEHQaA0oh0ptXjHQ5U1+Mc
5NQxSgsdsqLDYGuWXiwswC7FpTYO3aw9N18oFS8d9ykfnOKb80zfCuLb8eyaV4hb
46TkCIsOm2XBc7sCvaCs1dbXVS8s0zyfHXxopGDP9LoXBNwTjMd678w96amUvvug
mcABjxR9eAmYfJz7cE4j4LvOeVKAVLs0XBLLqyEFGiHsjC+2INthgBSs7LUOu/mb
k4Ao/BwERhmQUxbZJ9L4ZyLDNnlNQAPahg+mL+B8Is3+dpzawz8DBzMxS7RG+d5g
bxMbxfUSXquDgKmIt2YM6ahGEseUphhRwYPvL90xU+5HtjL3wZeY4W1LHsOC+Qo2
Y4gyb4GLodAvlFFGWjI52A1h7GjPY3z+vQ3HsjoyaCoJvTt97I2Pl5FUgp1Ak+78
m04RJ4ZAanrt2iHz5+NunJ8fKkuVtXgwBNkxVoX/8ZqWdejgDVtBEfBx5Wy2+PSL
a3x4Fi7lO8SlPdU8ajiEIR6J1r1k1lWTHcb2/XI71D70P9ifKk4EpQxP1kOLXn9h
KlZPEtu+olFx/p9XCDq2rvUFYfYfhwdtqrY+ZfE7rh4P3lDVq1TEWpgD8aTyY/pg
TkGRakhtfw2V7jIA0QRo16ZbWjcW5xzmVrr+T/SjxPoUFLibKKvqCTRuiaDzBeYX
tCaBY2ikp0Ei4roNHOwv7loQ6sIIOuz2EGjCUqeFyhy1sxA6SjJeezbaypoqPSB3
M3meDcucOXqsK6qhXLilLo9PfnKcG8S/Po4WY2KbvFQqrZf2BrZn8ND2rGgKeKRI
2AT+gh7Qq4iMXKz2uuEiSq/gpRLwPvslm/vYEE3phtwP7HrKEfy8oJgQA/HMsldF
YfIPyRnGTBAYrvgdYRIDHCvaqa+HDaD4WYPCUTkUh0ACxtw6K9zjfqWPpwTToK6/
I0knQVab1m5rsyJwa1kJntsOQ+ZD6kvPOhj3wf+rVbI90yV3mFiY616SkKsN6jLV
jl/fKWTeJ/B8NNL2JSWKhbP6z3pi6bI5Z3tdjcyt6V3SIRyo5sYtB1UWMYZWh+T8
cz6WWWwNgWZsMOk0B8oRAao+NWBNwBcv2XdGo70QbgzoAmpn0PiHemr5ik69JZWw
JA+lRBoBGxL5J+niiDY+Une/ANiPm0WjQWwF8PTT4CyUqmZyLiouerUti2W28bCp
hU0wTWdBPFqe2fkFBjPswpzxR+PAiuNUU2EEGyhSgIWpL+YZUJmjLFcUykP/WTKu
DO8GD1GRQA8w7HkeXgUt4IteY6QsDD/5TndewPkh6KaorU2iNx5+L/LNPMo2sqh1
vUEL8kLqqhSf838LHkRSphXLreclyFHr6BseQbj7vjvOp5T9XDyu+gT+fWD2jpoA
xcjbQpoN/9oga5iTcquPfIgf3ae6n9HtJ0wgrP7X1bAkPDY6KP+2ZTEJqyIxW1qF
ouL38X4AFCpfcTcu9kye75TvFK9MdHPSKRf0jhQHUAab7C1D/sMokaTFABXnZBe6
xDu5+s8FPzb9MR29thZ+LK4zSmR9aAyzWgf8Ezac67psiWfqlU4iZZArSGIsWAEB
fGYxKOLPLYMfaQklaNTGugQZwayW9yrVcGqAOn7JnxoaKgVFh9egpznt8HdTIb94
kd1+uVX6+ix6xQjK/DxOjeeRcOn1xKdo+59CFCGeDAlAJ58EIsBsxmafH4oQzSDu
Yfs8ef+0p6no+HnJbnBU9tY49HUVb7W9LM0MdjXSZViNK6dN/hcl/mXCdG+0AS8y
gfCt+CFzhEW1YIwfq/psoN2WrpCGBj1I9nM+ANakUBCqLrR64+JosPZ2BviUmk4M
szXPZKtjFiODpQ25VzvFV6XL0CQlQR7rjTE07XTxQMPz6pZ4na9MGsF0b2afduGq
Mb/F8Agj5nbqTITPUOTew9T8KHiMLxnPaH9yTjOTtj9W/1UrVFw59l/Zo8wToOQh
dPsF2vjXatCPxivgMCOLPm23p/chdXLBiWBICA2dnEgvcJ1x4QqRg7OoqWWhyrq+
aULE5gUtjnVvv+OqJhmPLnkINMnruIZ8ALFsVBX5hNWPjYnIgAAwoYtJ7Bu1rAG3
CCq8os54WLF1du+PLY5Crg7nTcm+gaEPlBGAmDOMKOP9ESvhudTg+6qNQbNXSu6+
V85QdNzN+rYGOrukAidGxBxDdGSQl/mMD+RJe1QO4BXoiH84l/5dTIZydPrrBs5C
nF1Ajza9OOIf9K3VAZMtjNVp/bDqiVXlwIJSm4eg0foqAjK0h0amjNRWRCtNCISf
q5PpQeagIPCgI1pd7I3wvKlIAge6tJtVI79rnZg6zNVQAZS3Mjfx25GWQ8Y7bFsB
oLL+BQw9mQ66MtKqV3avnb8W2dvTn0kRUrbDlfqqYhnsmr99SuLbMk6K1mu+qX/a
QYAaVDlF9K7YnWusBmiWC80oqKoadA6EXgCljmqlFyHJlHHSTOEpyicrLBdS7jiC
hxE5Gouwmlrzq7R4nTLRYEf7tardFO7oU2iO8KJ0yLzczOsp3u1olHnRsBpKbG7X
0XLCL/P56L48S0AH1gdPkt/YqwyokmfOqS8zDJ+p8bzwogFKGgeqtWaQynTP1ftj
LtqkN3D18QqfeWF2DcZGr2WVHiBGUEi5wq9FpujQDw9CdvLSZchV0b7Xmq2bwlcA
Sb5ame/gY1+tK93sCcZrjDOUnW+PTP9X5nuPRL2dfTI3z9zcYWkYvmwOiReJ8+95
qoYB9dVhATFuN3/rGwbHHt7w+ZWZPnD9vYEngld7NULGKCLe3XJFJwFczpic/Vhk
lOT4WrgSOkljoqDD3rdq/1skDWe3UNPU4tnUlGEuqZrF6c1Z4lv5tYdk/QEaDvnp
axHokgixHuH9FHFyLAgd+QABmqbXDJWgRekXqHNJ3G+PjesIXvIBASpQ3nSXKDIA
NeiUUt3u+lPJJ8hkAR8Bg5mYgonPX2daPiEQLXGiyS6nNoS/IJlG076AcQFDqnwv
LveFNWnS0MNi3UAgQje2NHIsIN9ZpL5CzJlGD2FThlpnMNcgMBA3orU0CLmpzMXc
Dc0xsjFZX0kcQKYuwt6yOb+2sshtw8rdq7iF0NFb5PIbz8s4/gnEQ8mUpO9WvGZ7
+vUJrqGeuegk+FWQ9K1o+F0DM0ryTJppOV1ANdY1v/4QrlUidgxUnEBlPOZ+eWQP
4RPaz2+IE9KGs6aOaTjLOKCd63aAdmbG8GxlvIc89mEkgxCgK8+vSi64VWhLrKsg
r5A4xKFXBXb1JPzfKL6YwMNh8oQqcXR04adRr0+zFuY4K4qDG0CS6wxUKBkq0vSo
WwuLT9AImGM34ltsO4/vkZrGJInV3U5cOxj6ZYdxy3BOE75+QvSOvPCF61fjntOm
smZZQYqrxVuLrBwt9tYtSymB6QKxmtsG5QbmcEILOl4s4ygsiHFgwA+QImoxpE6Y
4Mxo/as9NKJ1xSwUH2oglHqGLimzA7OdChVr6UqQss67zMP/RZdyqKj8OjQIhc9E
xUfGuAl27vQi8nakppMQJqEFNuys+NKbP9Cy4YrwuImothFeuAKTnXjZ2FZ3VD0c
Rc0D4zI2BNPMGIO46zRpuOBqhQ7uW2Ku4QBsHY7EXQHIrRrzl2B3e6gSTuMDDx5D
Ukxl+NuYYbsQN3hRVeqjX2M+Zivvq1qfHwzYdJqnLm45uJ6duH5zebV/mtubh1ED
Ov1p/dP5ZXP1Nr4gc6j0Jzj8KjSeUASrN3onX1qih3NjBY2LFD49ee9G+LwhGZwM
W4Dyg/zVJowiL/pEz3zDL18qcWNh0vyk+hZqqPhd49vl1PWmW2eIbwD7aEESURI1
1esjcBAvBcbperuhASJYSowhbfEcjWkQD836QSgpaZEw0tWuMqmPRCuZs13P+YJz
XekS+Q7f/KhNwg7qbpriwHZxLnoDS/By9MXjBo5GFemc/cuz6OgEMgTXaNwWHTzl
BLI50DXEVoyFExkLnuCjaOsO0b9QoHjZeHwcFHrqzOi2RfSjv1YdIWSXeujsp/Sb
4SY7iITZKfKRe+kINZIzOkA97pNjoqyqEqfHZWRTT9BcDQ68QBzyhLo5B+3TZrci
xwxzOcBhonZJxnBsRpRgbA624JfLvXVPq5D86bwdrD8iOdUQwK+nBagCnKovrzyG
kuRRYnPgAbk1BVvlXKvTUNyj2L6UYCcHB1cVgmVj10IRx5Dk96wgE523SgONzGTT
a7COiBiH3A2WBkt3vmMigBvfAE8+YqnHaSEqRTQjQmPz/q6ScKX3/RKofR0EN9ss
Pz5tArOfdF5+dXIFm3jIEyST+FWa+PnJUuPbM6qCbuvnAteTf83OrPsYRtTbHh+F
ZXf/cMt+zoAGi1QZNTp7G3CJDR8n+CoikiljEDlkJa1vBhxlh11eI+HvH+/t0Bl+
+4LQgGgeDiMgGjibABzrX8AxqWtXuQkd94TCbXIeamDJIhKDkC4t8zPz1a1O2TZd
M1Ykg4ALLsuoGVlMm2dwCTCXV0pBTkxuQdNBgMyctekwmgqs5/UUpFhyYjlMOUvI
OHYExTNi+E2r2gVU8RTn7PYmW3NJgmuAKgeuHNBG3M1kRTo3cpeo0taBLDC+7oPi
xa7NNHrenlEi5mZlTGgJs12HvpBmIxLqxh42RqTpDBZXk4Ay9BkXEbs1kaWf5kjW
dzNCGPcl4ARIB20rerODTGpGdd+ttHrFDBFRaS1/z7j5bZKpSzbNUSJJ5TIhfGTF
vQsYrvb8z/wQw7UL0NdnC1wy3j6t5MsY6HXGrkrHz7I/Gma/ourvLXpfTMdinvnv
YanISnyXltNjQ0+gImCL1GEpCXk5BAx3iFisWwY6730QiKK5MOWDRom9suMSUM5l
mpi6jTb4H7J3SoxgdmOt9ETRnH5aCuafDoCSL3rtBN9TwPvTAYB23jsjeWc8B0mI
NRAcSkDFQ4jhbw/jexwgwmeJIVdiy2vZlzZb3fg5VRPjDJr/kONidgacPGYdgb4W
BLXkJqxVO4Cuc9IM1XibfhkKZNYG6C1YW92F4Zz2hB1+CNbBAgdW1RaKVPmXpBds
pJGYl5pjKr3nXNVPpbFPHdpVrGIa9pPMPbnObVmlxcbUpgGV862F3aMwqtjO/Yhg
5jk/YxLyHSV3fVlka8JFNGGqfJ8aUztMTrbf8/0F9bgEOUYuuQ23bn2Dkx5x1u2+
yfcmWNYSZTKSRcWrlm9VRA5DLO48bZzQaGjiBFLqQVHYDoSJFKFtYvzFarH1USHe
FgcgElfB7lHkZEVc6OQhjKiWaJSce7JMdEVTxkyDWjVAd3dLpI56OT45RnSlAKr8
PaOnx7Rve8fFPY1LLLV6zlFQlsaJWCTPQtuI+8WeI7FQ6D5YLeOr8UeR9H7HyN9t
ebaJsKvKNdfbNzaZ59B9BnjwdQWePsioTrOqwMGR8Z3H+iPMj5RVpIje7f8VJArz
Z1Qp/Yu3AXLzcFB1wgRQNczE0jC+8jbLh5S2Wm5XrR9q4mQjJPmtu48n/0DZFwJx
iJ+tUfUn1SLy99zdezo6hPS5g4VcjWz9c/GSvEpHCMeKLWUXsDmqqgDYT5LsGVw+
Kb0+M8IOHGxfVfYPXUjM9Fo6jxieFcyKB1rs7D2XU6sk//+jQNKM8wLh037StdSt
zojfmR/3D9HTEUe2Ri6cTo0BdN5zjSVq1C6RMKBkRwnoWn4s88st3IRtQKoA2C3E
fHl7WgY27dIrDE1p7fSRI/fkm2IQCzZmVj28T5rZXKB5A10UNgISOjB6xtmCqE1V
qRVOmBJtgHb91MLuWpCTML2LqJq+LFW7u0C+mGld5jiMjarmSnOQJVWz4Ni8fkXJ
n6dE//dCOJvVqf9N1jVoUn7BDOVrvox48gJ7Vr2uaa3Eg7PZyVGbMSp33pxahPNK
bxKKtkY5DNAf3RCp3y9SqdfZv9zdPZ3hRx+YFskPZmjt2ndZ5+hkBJZAAxO/kn/I
YmFS+GvJ0l6kSSD2Gw9AhghH2EAoOtXL+wiKhM1wIb97P65877OMmrffyPz3h2WT
Ym6EzIxIZPc2aJDQsnZ2ciOYrdrQeMaTXDbH0Sctu28uIOuw0F/g/rK2Q34PnXD8
4pDG/i2CwL6MaSLLxYMLEjvZmIRvzP0cboa11x2LqyyFIWVeulDEubL8ReMxPtFf
2MHeDxvXgwAZQs9htH/MiKm0hh4W6mLglpkz/HZr73m1sXxvxqZ0Hbz960iZuDfG
AmojIgsrf7yFmRU9CdcXfpcdZQ4vBhC6sWt/ARaXdC3xnMiNE2z/kEMqHi8vW8CG
y2bfNKno2U3B24xXj5ZpG7ThFFWLJN8oC+4rPc44RwB1jktCey0RyWE99axyrAQL
vWSVoO8O/AenfnHKlwE22K1lkfud+OA618bwuZEa7QtYNPgCiU/57MajJ8fy60F8
57zZPMg5aMB4txm1wcNm6fYPivFDBnaS6thH9dmsOmkeJjQ28nmeXLlG66yCNqe9
sfcAk38IzYkEN9NmJ2uy55W+jq7AjhbiPIyLMSgHgc28zxsn4n3ZJ2ObaU0uUdrz
ytSLrPQnzMR6Ap3XfX8Ik621IGezkk+B+82dDLq5WhvcKE0dzarHq8is9OtefCyb
6KB5gOkU90tUipZk43dzamd08RV1/nVJAHUEXUm543qQVReyppKpnjmY2B/7D9NE
PsSmiX1oKedDhLLJpgq0sWF56qrqYrDRvTX9vP0+hCvG3mlaVsb5cKhu4JI57gJA
y8rYbAwMvINjyWV33P7Za8SMaOLxu/D2YGqdJuvkoBF85OVuuEKUi9qO5ai6MB0T
e2c7Cmz0lupQJjjANkDFR+ujoFKT+ARmi/OLbqAAmDbBnvAA0eLRz73cZx3anoKO
PfAsSYYQPSUN7fHOdipnBTgmLLNdVMGgyvLdSKWKKsqE3UIQqxKlamcM+WzDjohA
1lVH0BvDp6GkVA9Z51qdn4iDc2oN/jumDFM5RCP3vOE073jZhMiaHiKE5fb2Endy
dSOZkPr67K4MW6/uK+hUb6wR4CRxsp+2BkuBGaNUkL8zLSzpNXp4r7GM36AsAIvO
wN0gLOLV2ZKBCr0zFSsj76hzUZ2KYv85i/opn743NbcfRZ8EOZFCcKiVgYsZUQPu
yttX1dO+imQS0i7Z7YK7O4ch0IIpsiflDJsPW+eACjObb9/rU+dcCpDCNJixZqno
gsZ3PhhxJa8U7D2/eArlEXPhhkAZ1olPiYFqlTohOnXZUwwH+Ai9i91uLRMofur8
z6OkmTcAU379jvEE87rCYD1MmP69nVGZannlZnhg8svGF5HByQREX3jNXYg808SV
Ejl6P0UAPy4PbctPERpnbzDrsaskPRRVAfGA2WMa69m3FFh/G/WMWzQOZaJqQzyE
06HII4wU7vIhhlSbEZgcu+QgBtiIu4LRpa5ey5Jh03wVz9Z3BEUxxG4hpaAusBhx
uOwyFC6JVlcp1mBjiEQVJWF8D08Ztjh7zfAC/af3eqlSxkSI0j35O65ccJfQacdH
fZ5NJXuA0KGhAcPdd+WjjI3RVcuJuGZcu7HwVvcwJsYaQjA5A/mEo1X7OES5it0i
2zFeZOIq2gzzsLVqdsPOkcgdTU902UXO09/jXvyfkBTjAG2z50JlNbdEXtp3jN4g
AiFL8Uxrst3yxhyofHVvoaAXPDeHrr2m8km8NhthrewVxYjZGVy95tpaThQ7J9s5
749JT1jjwqichmepCOP6fTJleqzbOwwfOx3dmIegCTEPl8KiiUxa7N+0kGXE1Lj3
TP7AXTAzyPehldjDigldEADcNDyUpw1aqbxoEl2hKkdgnoLpxAPI9IiWfb4i11Hq
h8d4WrOS+unIOtc9rjrBPfWGX1yesX1YLLPZMpAyY3pFxVqUmsbY58bqdcdWqRYe
NJd2i+qd4CzPKSyHoQW/Icu5iJ4VVJAR+IyLYyXT/fXZDyOLtA4EEdQDkcgSG4tE
LfozVcvDcpVxwbeOBgDXY4F1pbJisB9J+VpBHT0advBROymBT9pDvyWAnxNje9Um
DHJ2ArQB7E9uCxmH3BKAeobk+jcmiyQieQQA1MPvsdJykfDtnx0NNnNowQzjMa4B
sJ9B7bwnHhUZM9i7M4JaHvplnNcLAIZBuOVCyt8wODUS6KZnyTzc6RDr5c6J9Dgm
LqM46RlvBnILUkK0rKRcT/GqzhppfYpFOBekAXpoym1NrkSP8eKWa8eeKPtpPF+m
hh/U63hlHf553JXF6w/kt9/L8Vx4jwkp7dNWmER2oDK7Ata1rEeBgS8Zk6si8gf1
3RBRRTLt079IKpVtAlUgld/DlpKKkoZ+kgjjp6uXqIgJWdghFQJuW5eupVAXpnzA
/5hOfjbyrIRf6JFLN6bugSetrHDt6MDzg9jJ9vXr81VD/DHgpnu6Z997uiL8VTBj
FFC79I4lERl4KKfXuhktDnebrjsL2E9siEPjMsCnc6/EogcslmtTbJ9uNMBSfDqZ
RajfICilS79CyIbSzdZVXuGu491bYb3lG0ebp4SHnoFG8ivk/EGzSWT4m5M6J3FN
eJ9AJwqyHWNZ0wyIncQfsXfGRjnqKVGrCYLDdwbSAFE2wJj9KpknNVbqkWYCAlOP
17X/Mo/xEKm1aVtJ0klugM3PkuPzjJ3yW2hujgHzhUSeXIUPzmReOIHH16wmUwmZ
lnJVSm3TCgr7e9Zec1N5WR7LJL+ZQKsSTsVui2aHx6NhBr6/5TT2f74pNWSs7OtX
2goqMndM3d0m2O+Y98KS77eKTJ4A+BLxVoGUvmVWK/Nu3YJ35M8+aeTkIPZpfIWI
v/xEzS2cYlYNR7JXdQ3NoHGhKi0RoU3ONPLTeoUI6im2vf0S0lynxc/CYyqsSgdZ
FG1zG0K/G+0RyqJyQGmdpfOj02XO6NefR4p2cU6FkLWE3pf2XQ7RGd6yfoFjBr5X
FyvxFeY44p2Wha7sCfbJ3gt4FI/V3yeF8d8Bs3w9r7eSOVgpZjsTcdiKFckwIa34
0UnoM0vAJqiEAeOemXms3MGar7GZiAXmMCgk3ZKILRCq4L5+iE2pB58XWt3JjHcv
fecAG30HlVmh1LJEtDHUonSsqDlS9l/4kNabdtGtaB5KZpjdofzql0hzE8rhyHrr
NwPWzFBJbb4PC+vnU73WKQ4wC0JHotmIka5o9V1qMEzGHf26bdp57Im6QOUUW2LV
pkBym67nEdMpE/1Y+4gP6Dd97rMc+NWIgFqPkEFCxIJgoV360fOvR6w03Rn5FthQ
ZDbtjQ2uAeoP3POCG8NTTZbHFD+LKoIz0C2dgICp2nIjeSX/FDe2j57HvRja5yRw
MhdkZvmbi6JPYqjubo/7DdgCBSUzDAz0iaP3aA1rZcMRi2epjPIBNBo15f9bhIK0
EYGXMFSnR6pjsCf6Fq9KWae7tbZlyu5iOwtJvpdvZPTMK4oDel5la6Ix4lAHhZw+
gFmEPZHU7eBZ3DCjaCpgho8T9fF3m0YzMARTTKMpCgmYP1fKe22Na0Df0rTIQ+Yb
vgEeDjfisx1NJXMb/1TTRuAJbH8B+ovpNSNyifCq4vkSQblnbvClsbvbY3GHKVkQ
qoiHuBql4LebkDiWknJdvLb5ZN5VHFLR+eq2DiJ0eDS/bPov+/bzvAoJq4PZnSO2
ngnOCSuFqXQAxrF6VB87MQh/shiiKDIW0eQu8fEckFGlPrsMTrHuuqIMCSyElk98
HqTv0J5v4+ZNiy7kAH2jkJLyiOnW6PZ38YEtRk+qg3bXKq5P8srjV+BYxD/lLGJC
/nBIyzZ06Xpd4k9TPQByMjbFQ8llEtMmunMpkYIkWCaNrLJc9SaHqWCQqHykGOSJ
XYyNN3Un5DWNksVU8R4CklCvP2A0XH+tHDC96psk7CKHgi3srpQc30RXptedvwPF
0uTVRomCRlNJ9bct1J+d7h0pvwKWN1vbUvUfdg+97+3D2blxP9gD8onhVVtwYRb2
sV+aqrETT/hg7f/vFYk2mJXaBvcqGTqUlyFEypqlRmwcC9WoRsGsSwtWe8zS1rFa
F4YtIL9d1BKOWND+dQb6jRR+y6Fw/NgFgbQD+fW8YTmS1TXB3+i/d3dSQ8CR34+s
/QPKZ0YXLBvz6L7v144F2B21EIht0ZwUNBkXfWvruNRaA7DsGnGMriw5w04DYmNS
embUXDePtgfO0cyg9ANqF4ZIHPHAXcu+jmp/ATn4qdWS5De9XUHir0l8eG2IOvCH
wLUAgvnNMx1MeqWFhHtGeyJQMD9fAbcgswLnyjaWPcND12cqejRuO3MqhEbOWtqu
n+yL1gjd9HrbIw/wphLLB4Ym1eVz7SUEq/TO/WgF7W49/CkRqhyWxkYRctgRivIC
18Ri269GDKTI41CJDrR6v+JV5g1vJ5wBaK3VBCX9yB1f6PxR/ejoIPQoQ6FkUpbJ
lY2/bLMWGYs9WiMzQBxDX0AjTixlst0kz+Jkq+AYMlqIFvyQf1bx19ZW0YMbYqFq
TREj7NlcPBt1s2WmLQmdpEKiAD0R1+22zWg8y98A3nIr6KRX3zSi4cUadR+lAt+M
5dncdxzISX+pkeaEBRBYL+y/T7ccA4ibmnVFk32FflBhPBfqZ/RvTcqTIVpeN1RT
dHBQ8+WgBHYb9OC8Ogy2LycdC8tCDXk2XY4Hf5W2fuIOQTu8AgGHs6oCOkOeMruA
G5GcsNkkiO1a6kN+jUK5/Fe9GrzBm5UAmAqZnE7JZP1AI2H9jTfZXeqo+1inP8nV
LDRorNWDbzFdWvPeRBrWnrHoInBl7Mq1qGdaUfRIU08w7or+pAYlSJi2Xp69ehvg
J8KCGw8xtiydrbg+ysle7hjvkrkQcKHlQB6fosWtejzo2gxjKsnWukM5eUvfWhUf
Wr62+wJ9/kmWjzUedQDV2b1iPqX0oa+mTH4dNgWQpqIfokkOz93hDwSNrSa1GGuS
YVCF9UgpD5PSwK+aCpLOMSYUMBb1/+IfMdmUjEVtWSZVuSjHTmaE+EdlurgVu98X
jJ1gWW2aN9BV9DjdcMzlcAK0mcTqkmOKMqYv4uY5pYgSDZh/vxw9ZxDmgyOgyh5G
kIQfQXcA2ExncTNnsaXaxydFJQdT+Gt/+l4rfxpl2jUuTgvyDZ0aOc++SBjDqKKp
qVtdMDSCbeeX7nzhXIUNRyNZpuFenJDRkqJyK/FSBdheqX+Dci7nCOqXQah+JCsn
vJRbFnOIFRU7F1lT3Lr49bAaDkmjW0BemECb/7C9XCJKJLKZGo/UKxjC5o/3lBLE
NYxlXur2RtFXLY8B2O7ZJisKCBP46VO7o6wn/IhqXTDQzJDCh4qvzXFYGXItGiMo
UAbVO1LoQnlZP78d6I27lhQRPCAgPMwKc6AII1Qdw7ShA1I1fjAGObJDzcEunYjB
WgAVVl77f7+S52gANxT6TF/+4brnFVqNmwCG6rLuxp47GaswOfLpU6kXvNtMgIIq
5Oz3M5MEGZkOl/cb8r1fwL4W3dWLa2kr3vJNNKIEhp4z8bNCSWvw8YaQ4uqWI7Ws
vYNNKM3FOFNrWfFwk6txBS5mEdb1PmeHCJJXw36JvqUUzkUbtxWo4RGRAqrWZo+U
/FHFbZHI8HpnOh9tnLYpP0DhknC+UwNd2xSr/175wg/O9VtSZj7tm6giw8ykSXTd
4MQ6HJpHy8/KIvvq3dDauA1g2EasdFFNWJnzc5SqTm3Jk6LWBIJR+TSsHF7jVyOs
lcbMAADLn9Svoy0rq6dawel+WSuJK5ek213ABG54FU3NsLuMiVezLO/8YVk2M9/c
Mg8C6/WqelJ0NBmMGyjeBGnLinLzXAbHEc+GIdPB2NAogakvAW3BNT4fx9KjgJhM
2OtkzopeUo0ZgN2ONSZonIhWwnVejBIKEtzdUbgBHQ6HwqzODwY6l40EEpOb68UI
jvxH8rY81Apv6QB5axsAdJscy0ZSD3A4TBETU2AOT4dFk1PCvljgesxYYmvmwsUt
Py4Wn8+mcHHLcwtR+kD+r4h3VOvpwDp8ytzunXOwkjqi4MJVathJna3C28ZlOOBj
57NVbxfLdel27PLxIqtLQa/dNGsvpkW+1xeLEwkeJiI1OFUXw81vk4fheXxv1oFH
bbFKcXfSnGDOvN8WTskN1/gSLgGL1rc5YszFcULOLSys1fVhb/7tYXGHGfFYVibi
cTIflrbtg0nH5iQzxH3Gt+OZlzSwPKD56kTyu2uTNJGAttdwwVtgMeB5XAtmMe5d
rhh7PPGlK9yco04vV+VqdqNkIVBLfOYzkFyWgT8VDt6feJV3jUFSqGdVmMpAuWxl
N+tnqWB6CMh1JvHaecE5xzmx6FpGEm5pCeDtYPtYRm5MQQ3983sHfi8RIAXTNea2
kKuBJuv7Kfy6wShSbB6F4pZSs1pZwaypSBLFI7HI8wVGaHXofk0TbuvTBIHERb8N
ZqhnnTjj8R8QHNU3J2+EIRTJvbNnusfRTRz5a8FEOsFn0OARRHOndfWC7QJZRuWJ
xnOKe/pALz1uLqYqYChIUi3/Xnhb/yIrEoHUvg9H07eEB+jdR1OQ2IMPR+9kpAQY
9cltl414AedeWfYzQLlKUsVk8OJBadoiBpuZ0KmNFW8aJagDijCQzC0y9Mvn/IO2
4UB+a7fZAMu5yGpUWJaFj8V2sjbA6Ud5L9/TILKhvNI7vQvCubOnNi4d/JCd+TeX
wSfEIwYADCod/jd2UCT35kOsJjLCBW1w4GXo1rxXYuH9gijB8O3RumcYkpizbNlW
Y3DbzuIJc4YZJUrKJbXaJA4uA8rDYbd537LFTxJhCKY34bGPD5x+J7qSWf/CgDex
gueRxI4AaETe2bVzpNCsJm8f49CilKzGSxk8cXqZJvR5ZfiQDcrSBPTm3VDVUU9f
Cz9pFNzAIcLUq7YSuKHRR+RUJFejljrJGi1cFNKa57y6tsjf6EpkARl/K4Mt7pu7
cvLdN1L6kS6z0X5xabJxVQMtTpR+6XHXv2qkZ1zPctr5wMOuZfSry91XFviVpufE
7uuneaLXORIhWmyVQ7ufOJlnhK1wIGnpFoyAY1Lzmy5JCmx4wuoUjtjmym/gV6NR
+zHjZMKnQkfYKWxzlFfB6cKqnuW6i7vRASO1QDTwxxcOfHDwvXlrO9KhAGUdo4L7
BM5gnW8lg0zzTkZCWB0TWlcoEd3jRY+m1W8+Ov6w6ynFpp2Rn85kVrC4kn0uBJ+k
FUg5UbFyt3/Z04/o8G35shilSlZHta40MT7zrv+MjIS0jrM3u+ZZpWDyGUMsnHDq
+cohhv1qaH8Fcy1xRg0XmhSxMLck67mpyJSRiPHgRQyQt3FFXJNc2UTSGRa4hFzn
Jy+dvNMCY7gLcRpD9Ruts2l7mp1S1Fta3qdF9eGvGU2VDBheMQIwGBaizfUsUNui
L3+Hxdo0X1OknixbpwZzLG4ZFrpI9wjOlFNITiIUiC5smy1JfdwjaZ4/9CKW48uJ
DNRFrsY2nhguM0hLMUPlZNc8FMApHOFGc+4eucBB2pigjAUikJc+bih3g243ZpUs
mC83PDpTBIjITOBVOXHaIFFrlB48xNwLlR+NyDI+dMbD3q1adiohUosQ5QHkD/1A
Ub3Ku5i3vAxYLU+kuonR88XmimhXAGQBxaH/G3ywSs8SCOaBNFTafhQ1//VBvVli
wWa1JSalLk8KANNzJg2AlBp0UMO/C8h3UYIMdYfwLvTzkz2Gux4nHLcxckiqXjBZ
iTgULZnOllXE/2Dxpxsn6nixYGW9H7QQJgZ8mUD4lO930wWNZa20/2YjrxMx1rBs
Ye3gtpFMNpCJyVGrndL85dvHYkueFwrdj9tlp3effH6fnFJ8mqSfwR1HOQrcrrqU
WMv/LFUmLRRnfn1s/77XeHcc7J9ZjBWSOAPLM6v+dXqN4dcpEoUQ1BSbCkYKz36R
GwumPHMxJIj4f7dxnx5h4Zup12l3Nv06Pu6tkKdg9N3gLA7EdmiqIDyZM4lMu3f8
eHplrXb7q58FA9cL+7s+VEAxNYXmkxWrLpLvUusgNDWWNOT+AGpUlXI37vf8CCK9
KDdyuEJB2fGo2SmJWOn1hJZ7EiREqeakRaqP5Ddjiwxp3klu9/WBRfSZayiOs+JE
9vpKchVWnbNO/5jGxxN7l0gG1O2wRouIPXUipWMY30jJ+A5tPjy6ZMiDxt2btTGl
cZdWdF0DFBqAe6GQW0HnOtHN6GYuJlLDzK843DqpmEOo1wrVIdk0pFw11B3VpBm4
OUwiGgTzIVLCSTJMrdOGl0DzjNHZrEUOijEidinYQkdKpuNJx6aiASEWroyZRDs5
upjJhLcuvAk2KVQJyga5yYE6dbrtHmmN3sanupOF0RZkrGWO5e6N31aHUwfkKHu2
yWi3Z10GroTzG1VElDQLZOfdot18fqZS3vgCjf+UIEB8aLbjQgSfj+e+UfU75MhU
6C0xtrK/wGAZQ8PZgU20GpN1ygr6WRE6OXQ6fOAkgaH/Toc8LSNiwq6836PzRExp
ZTL5KD3mOyLBv0muTM65aiczc50rGBAEj58ixVaWeHxSwkMnIbhUoKUQfP15AGac
7+37Ckvq6uqFePZCH9FLGnqKupPpP2DI60BNsGNDEFnwR/CPi+WRuut8RFEDKgxz
pE7bGIdahXogS5aFnOI0qVxzqvMU0XDPhnQOhBNbgG/S1V+Rc122T0IwfDcAKJmU
9DKKOXd2lHPbcwYbGgWldSSHU1wHD1mtl+BBJQA6AZzQu3p7p15sR4CtCXU/CBur
F6cFMz9u+S6lDJevrId4UyM4i0f5aS0dkwC+Leujx1WPHK3Zk89UfOoT+XmYYgQM
ZsFhiB8/+0m0NOPXwEhLDL0D2+WSQ8wF0RH1zLXqu8jCyfISu5TxkZfIsGGXvSAc
B7vnP3aqBFXzQ65dQ/XGFetQARXojeoWiItBJq1WNE1gIilMtCf0xsxdwScuvOXG
lWc4D5RdVGvqFCB4W2Yj3TfgCC9yWVtdILsalA3udkNshTeEhRLCNAS+e2p0CqiJ
GUtTctY1L8e6W58Yl3m14Gzn67UqFLw0R27vz9OIvK0nHg7AahOkV3pZ3cClUpbO
5ut+W63SyYoY2SaUw8iLiPJCpkOIhS9vnWA9FvxZIhNX+4jWQVBCebmyES1d5mR2
cDsqHFGGC2x6j97ul8HIrNaTH2+hzxyIW1y3FztIl8MWOenMB+3WG/JeZ12DCjKW
+xaim0/2EK3VHLhnCyYuA9pK/xIPtks9wAARqein8wxzVP8hJ/KxUymZRTf09lZT
u83R0L7M41fk+jhYOCMWPV0fwYVbMFGyR1AQj50CXWnQpfu5zn688peqGNMwLFLg
HYtq2FEIvJF+1uRBvwq9lqKWc4Poznu9eEuJqRfsG9qeTNljQTSYIiJJZV87H1ZY
xtaIO/brQ3xaU0lCr37dWlc4QEXmhrJIupTCI5NwaJ05+Mjr6Thn05sGygytrWVO
FAvjAFkp+Tt0GPiFHyBcOsu7ZJLjXgr/oKurmvhpgDWh2KGYpQVaOy9++tnHiPNM
BtKFS6WG6iAoUbw9db+JqleQcb7WQlzG/AOHxOW08m/CPSlUvmCSEH+6nT9s42eV
PwAmyuMKtmx6PlfQiVdmf8jSeruMz3oO9XLFubye6eQdbltHnWg65zoXGBT9PWSN
Z+Kdd5IpunCzcDvB9jpHYvOXwtKzBq6TTsUHZNgZ9IGD6Wsoi9LDe10La+raaGgq
FHQvh4+/xInYqt6vl1W3fnlLVfmZuQ6z3ZKqfgw59cglnwVSqZSJuD1CwRJoSBW7
z6/cNaLNQgrfCbJLzsU3U3IilKdAhFsJI0+JPkgy0TZyfuzrVO4I5f+M+pdkPAfD
IhH5fY8uteKjYYrZ60emybvmx43xiqzSK2Wp6zDO+jYToAaVw3NzikRIXM8490De
+g36wRPfnOQbgwqK5Ns2pH51BE7fKgtHXCTnAzMmKeZwh/h/Z4vLnHJB01j12kI9
Lqd61GhJBwBpcZLAP4BUU2oh8nfkxcTmEbDXz61JUj7NOoicPLILFLh2gMxB6WCr
uvAEJ5T/zJO+oRP5QDgMgMb1KBanJFZX1mPFOyVFEeQA9S74tDXKu4/HPgBTa/vn
SSZINXvRmE3CXuU5icIKcvFEoHKsQMAYDcPVk1OHyPc4ZKYBLERvXGaWuVC7j+qX
gv4DeF7hLnPfZJoP3pVVO2PYqqEL3E4wXxllAw5zmq1p4S3y9DIy3sqE1VtRBp//
h4/CwvUAVOWbZ0eaeXYnqTCwHjQfmTUreXXTbp/XAl6Fp6+JSeoXWIatnjosLc6i
KY8SQeYgLJWaNDcYG6abnu4bJFTKTtduK3d7bnFKvweJM4jd9mDysK6TWJXu8hFK
AUShYZoqleVG/reoGeKt8KSv9HFyJ+xmogSr13Qx0mE4ydd38+S6Wg/hovQ+XWHg
jnbEN9HuFJO29393Gc4tsKGJRD4eym0pu4PytDB16ToTU1AIXqUUZ9y5b8gdeOd6
hIjCM0JM7FRLYGRDUnZSGbKWGYTD+7oKn0lipkJgSGrnJgxVI0VZpiXI2L7ZrezO
uKeYYmhkfTaIGOeBs6r5M4GHlKhuf8Zfw4vYYFIA5CXRX01VlwPIGPqXEPGmlP/W
60FFgyj99rgq0aTdCJcH8BdqLgzlTkUrbokbe3eP/3Ekspf0hKeksnr0P7ijB7QV
7rR+BQMxWkxNDTOpkoJ8tyroAAEKP2WmQ+IhZTRJZmg3c4cDIJbmFOJgAF2lJZMO
nMQF6jP+5KiYY+J0QLx/29NxSrfM41strGnXsvJeKYamCy+oqkO+RQ1yNLN6O2km
b3CTh68lAU0Lile/wO2/IHzj7jytPKSgOPzQcoQhQhBMQSfNVmQBTVii7XdzfDKu
TTnMwyn6Y2tPQY1I6Ljh5NIfC5X/egb79/ccejVJAwqhvpAGcDhAlym2PZBJZnE2
Pm3/47ARMmZl+dmOZ0rFX3L9Y/PP10iqZjnzbRtapFZ0iYoPGycAHmNsVaylTmtI
BDpQTMNcDGveX9EWpvvtbPt4UokYlHkjMGran3Mm76cVO0GbhPDv0mQmf2/G4Tra
GpZueAny9HjrXCQeXDh96Yx1zr9BBHnCplykJBSqc3Soyvxu1YjZo425jx4pjtLk
APT+sJgSXm1RhfDr1JdWQTbJ+FzCmlwkItRMlY/DFObI+ZPVqRXU3STNKZqxTpFP
v3KLob4EoccAeiQYOnDqp5Sj4GXoiKH2T4dQDmAZ3dlCRkgPg9e8Fcsm0LEQhaVR
LDholHxjklmh43eq/4u1fytGWlJ3OUJQ5NQFA458EfwVSEFvXy9p5ran/aKbtScP
PyMfY0Cr/AEpKSK8tg0k/myn5Pdg8hOq98hy3tCFBXFqgf4tHbVyojpe3Ixtm/3W
Mgvz/bRmiIW0LUgy0pwwTLuy+3gFemHVO/7fR9jC3ahdUp53hDnw1Jrcx4esHLch
ARRJvu0/Apry5VA9hC3CIctlKLltctGNUcWzwVNmlmfHEqKCcQX21rKDerTMzfJy
DdwLGzhoeTwrZ6SCW0EXlr5+OYObJDe9FZUVL7QgasjPLlHrjLwpE7TWuuVkGDvY
uaII9dEvUP3ZIWZcpYgfW29qVKNycBZwnnb59Go6LoEjB8nUd7XUhwGowlxNsThW
pA8pUUPTktvFiE61J/Zttssnuix2KTeEuEYBEUR++wtyzdZQ+G7A+csmz6w0RdFK
veK5ekNO+l7qiNPljUBgcLNdvHvGVfsc3w/IFvvIHB4EqWjryCjMcHjM9hSemLya
VFawYlp7oesvvJajCrrSxgfSVB7olyrzZKlwWvbXAXylWdxLGlLsu6O3Kz7FAFG4
Pa/vBmZKBLu7OQeTxwR6SG7sFM5LcIcipaqOeIuu4PPxHB5036Of/dhlQtPKRpdR
8FG/XxNOlt1YmjLc3etu/h5a3LdVyf9sdkvk+sOqq+M4WhAfwwcfeNYUHz1TuGNY
pu/U8crmmGG5RhpF8j3qhUevJxnRxLpa7gEWRGve4xAWPO+Szk4x7HXtn1Q0bpka
2unkElJicyTqXf6RI05G9e9JtYfUKXgH8g8tcokvnp2xGcGZmkmXgYz+h7SrUOXd
ThJI9CW8gx83ZacZr6x2T9AzRNzHtzn7kKoxx2bTuWSHjB5paPTe+3bqbsaoAbic
c5sb2WyQv4CbEjaivwBSYPZWtnT5X0HsLpg1nZNaAZBOSsQAqIQpl5lkkJBzN2I3
IIyqjmqkSVGoWJ4dLwLhmqs++b/gurslIoEOE0NKrU5Hmxk87ixDRuqeHSWSiTyc
REeaHoCPNh2iYvd0gc8fPI9NBSV90Lz5n1Tye40shjKpfCB/06ZcsYzhSWRAi2j9
y2TlxoTLThrtnQVnhWokK0SxLPV8k6LwhgIrJtmMh1e2akI/1r/o386FjFgwQDhZ
NMie5Zd7yrDLBYkRFX7r7c1mv9kflxEuvst4kUirEkypIwChpZJtGiqzHEdOgCLa
92j4RCrYpWEoAowr02cY979HYOlalxbO/bAWOrBJLzonp98SXX17tov7Rlx6U0Z3
aSzCxLfLHpubJ15QF7wBNUrdp/6WrrqBpp+RLLwk61GSu8aDLwhDKc7B32tzqKVY
lA/lGIIFheSKGP8DXOIxDqYTNyP8zGJ+3ABWJcKzp3sncWyujwbm3MJ9+E8FSaX0
92SkRgdPuOczUC1A9RvymscoU7LTq2A+JSxIDgDBXdpqSMY4jS8Jt2iNa9K4/0Lk
dT7muvOohcGuOxFXHaR8NzYoAxq6Ytp2nVS87padz1GIcMk56f9FfuGlXCgLrHMg
gnkMkzF24qe2XsJ9xIG/9NXD9+TIaLxJAlIadLBI6mUD2AgHMbjJHX1rozNK8I6r
Ytu5qQEHPnBGmV+MfNDdJhINbl2TKkLo0p9vJ+jDyNk55rd7iHiNKi46kTFhdy3O
vo6MdNzmH101M8+/Gm+l8w2I6tA9mSHJjnKoln0OgDZerwCpNq95dIyPRjv3E1cV
Fapb39ayA/ksVaTCzrv/yk32awt6NKCAd5suPx/OLpdTfeiYjO1ILdAaykAvityd
s9un3gesVX3CsVPqt4Q4UzVwHhJGHh0oOvDQfzYWqWQE17R7DUHXezMyL2uyRm+R
sHQUcyoPx5nYmCxTiyThCuLj1SoCeq7Rm56CoEcIrSQSFf6EpO/Kd9qFBNVPMrBK
oJBHq4K152Oac+vi2BFolbMp06gQS/VJ5iGEEGepKt9vzNKx2HvtonJOyvf5NXFD
dHUcojpaILXq2dIRIJhgq1cJzkusmlJWdF/mt/Safnb9wSNWxQawwLzL4BzVasfi
BY8619Z8Hq8XnaCLXzQYtu7WESFUR922boubD7WMPbvNSxNxAtM/KU4gIbNvSl/C
lNnyJggG/ykL3fHMjJUK9rcQv5Da9uwifFu4mWOBwSbnJBZjyuB1bwRy6MxDkona
3M+YPE3zxipqN7kQ2vQeK2FqQ1kn+zTdm/VkrqViZBJIwWAu/vVt9ZS0CDVgM4IK
L+aGHA6F4yLKa7cIdGMMUOlf17dAz/qB8tvv1uhwh6no8SzW9Z2SaP+zkYMGZ+ER
eMkWkOoqu2tNxytmSsPulj3btwDyeKMWwhrnx8X9chRpPbncbEJsPnhBc6bGph0D
7AA4SlKXtNjbBvSaWqHNj12GwOBEAy6YUHRF/TJbl//dl61SFjnNQxZkt9XDVG4A
untszzW9nr7WgMxL3bk/LBB0Sn+RdA5cDHchly7b044FiPj0e47DBFZMbAnotMCn
Tm25V2quo8nSCi0YL8WpguEx3V2pGH36fJTwS0xuZKdlxJUO8d1TQxF1cPkuTxBo
hk5xgQd1RKnsrB7hM4WTXbCYTqQyyrTwWpRHno7U8x1RZT70XgrLdAJmg+hfSH94
uVqfIBCB1Q8YpJF0EPPxfwsQnMV54x0F45keq5UXTBRtcq4hHWkaGZTHUXMTu4lY
i2dDdyX0nV7JfTMfiGeuYxPhq/qtHkRdvqTY5Rk1Os8IEFjkA8UzwQk/nhCEBqTe
QJpcU6fYXzqDOVQDjbRptdGOFZt5BDDAiFtKzDBPauNUNYYzFNwe1sP1lLRGV7RD
1Ng1RBWINsBPO9G0h2uYNJIQRtaxJV/kXUf5pzrpjb4Bu6EoKVfDi2zoDka51BIi
wx5hO4gLJTNCN/S/d80ZyvdzPA1O++FBQzLo0wUFqo29FuQ62scYs7ZYtb/d2Be7
yBcHNVleNNt0Y+xUbeBcTF24YX6yJ/IPNcBqKmyILFjHIEhV2L/zMCcKvfBG+aUq
YW08R9joxLKlPeVdh/bqxYdeKwtbUMVeDMbCPGxhRaIbhUb70yQk7HYlGUluKopn
OUnC0f9H+E336mkzOH50LnbiTgHU6ekTXdZotd05iygSrnv/r4vUhMNQ9W9SwxWF
+dFTFtm3YhHpBEPdovuc2WOBsd/tkT/bdC1xhFb1srA26T5Evsuo2ZDyj4laQf5p
CRRpGBq3dHc/7YCdCr6BImdw4tFwVQIHWtefxgvElG2j7ZPdou9Y9jUE7WNNZCSs
QNRUxu+zbA/CKiYluiVx9tWR08vBDkvMBoyizKaDGo2VhgLJZI3zqu+Hgj2kK1S3
odWNAWpOP7X34fCB1Z8GOYYAVqTO+9ME7mxkbNInHhpnJ/+glsksQsxL230SSoqV
sJiNPbTMWoNq0eOEA7bIPOy9/ObKloaQDpmqGvb5WwYUHy5EdcHKeA4G+m50xzYC
86QgWI6z5mfm8lbjr2ZSWHK8AX7zbREbrW0ROwIFtuxXtQleYdFmwvvWQdNILZLt
TpgKqxFguRPI+D9GO0B30CTv3cXZYf6nT0Njoj+WzJ3yYBMhWGl8uBBP0geamNFl
eGJ6FRKQ5Ra3Ag0K+T7Ca2wostqbxW7GdiFTXU8bUDx9Key9KP8BsCTn7dguVa5O
ONlFlSiH/CXl6q+MG6+zMMpGTON8q2zXNmUR45UnG+fO4heFRhwyXj+Cs2cxa+t7
yn5j+KkBjJGMsG0KCz7NdrKs8jCKUu1jXgx/pyWYRLhs0zGJyC2y2PZFlcDEoaNa
7FnF36XAQqyHZ59mipb5RxS0qYX2bbOd/hs4nmZsmtzpJtD2RXQYj78Im5hNeog6
ytIRiqOMUtpdXa08BKElUKwjz82i+WQ4PjFNcH8alr5qinHwN3pOWqZmBAx8awkc
nxdNbmELAcLfGYyQX6tTbKd6GaQK8yxCkkhLTkMqsoopAtPZdS7O9oU60Ctpr3vM
44P+u9edIVy3Tgkr3rMWTXU5BtLNLjxZ0E43Ppkz1md9veduJlIzuFWObX28pT6S
vHSgg8hMviip38UvpPDNpPgUSab1APQ/6LM601rC0/L6dyvzmyBmWHAt+tFAKNQ9
usJru5cVROQuMbgnX72bvRQPCEyrKf1XKerO2QUnO3NsgG653kZL/FFXHj23b+uf
28DvlBs98ckZfWFTmWGBdsIxfT6JCa8ONhCpssgME83HsTXjw3dIom6tMsSp+k3Z
2mFe6yoY4Gg7x5ii5kefojpvv4bsp3IJlw6xnAtNiqbasTwcjoyRQObCNfpHjs7l
Coctr546lo9BYmad8Aq3rNufI7KpL+9cCFCOoWKMgLnenLOWWeHF0iIhtHLNIJf9
nGNRx5SktqGwFLU5qsH9XekXhE0WpE4W41gYdaEyAzeOHvMM/Jbc543rvhM2aYtV
1hmLhiW98i0YRRrRj7O8ieJGNUda3CaUQX3/UmRDHJoEuCr0+z+jbUsP6ySFsPHl
wbsCWWVA1U4/w6qOh5TVqn/xpR7DxQdTtNYOamiXUPPBTIPotkNXrmTAmri2uouh
HJMIzlKwHMs8bxdB4uYGiKJqD0HH2zPv0KMiGlf2FGIriTIHe2Yx6bRqJK3lMpFv
cEjGM5S2azauMKP8H38c2AsUytTgprUJKdTw9Q4jgWXYXTzD6qUuMQQ5WhQioNFX
SXcDnjmcn2D3unXxB0gJ87G+9OjlhHiWdNs9cwu7IM8M4LQnwu82TsjtlZTeVMyb
FUVBkfK5zCalaJrcPSksdrN9YnJFCKtKlD5oXfUrvlMsnLAk4HLCrO649/QKlCDF
ZJ3daVO/8YdOSU2p0SQ/HkM9RYshhQqTm2FTq9zQ6XFStmnKKbdjAhL6+ny35gTf
+Pd2FQR4yrOU7n4kZoBCB4dI3xvkxncga8kpCIKJ7QyaArrJJujFvis5PvhVlWyX
SyQbJrntBPpK3Rc7aj8rbGQ2Chpj0A37NFeX8NpVtgDYM/UDNrZeRsznzo365VoF
y6r2F1Z5sqhtm/LChyWfd7ugxST6PEp6Tuw+2Hdn2R4bDCS+hYdnZz2amZpKSWov
23A3wkzVr7e11YDe8839t5ICLjSMY/7v/uuM5ZkbwAMcikXY0Y5KPixC7/JYm1BL
9Z6uaBYMFrRWt94a9gtErMNgNB8QViSgfJ3v179cA+7ASSYpL/9Fy3DKSB93Ff7u
Q16xRz0XnGu3bIj/bRkjC2E8gkd/4ReyI7Hz+RxBUN+Hq+CumOI6Y1Oy/EDznmpD
nrXTCvBGNCMeO3QkPK3u6AMzx2+ZEKJBx0j7kwTRitUJr/NhleViMNtx13HbeuVk
EuJMtJYQQ0yhslqXOzBsEHtlhH8LGH4F2xY1LOwF3Aa9Y4za6q0GYV9uhSmdc9r3
wwqBT3M+8yiy/y/uQyoRhUPQwA9Yclcm0hBmC71kDWZHv1Q+a17zjY7/AkCxzcgj
65zskhckDjYM3QHdGTklmiJT4GRRt5ocahj123VaKggN5GjPCbKRHy3oy17awK1a
33NgJY+4El8dmFbxDCYQo+JgMmP7ypy9VNbBe/DF5wMIOBwf7eMziumard0RDK6K
mUDg8iicAt9VRjJyHSh4cu/0CdarF2pQXrwlgNFAeQRlgoNy/JhRVozzc/etmnVW
XEcnNRjaaLnX0ZQmoUn+WVwiQ9KFJrePPaxzyagD2ze2eFt0BuLBMgpNPnyc7epS
y1X8IS89LM9KP8IefDJKfU9Na22WDPh1zaqj1cH2D31kwRX2ltEIByKLqqINqshc
zfQyEL7I4shtOjz43TcqLY97x1p/6KLjV6GUqcFHucEu7qIOB98KnzOE/lqX1KgK
nAD+cxDaktAaw0yu2K5lR5mLfDjaMZxljzmMZbbgIYchiEa71clI8OiEhZHRMXpx
Ejgy5buvSJQ4LJcroPudZUw+3oMuknIWZK/aZSgisVQNBp3/vbp20ametndrU45n
T/5jMUiAuAqR0imgDtlvAI2th8VbTs+iCnydOsLmRtRAx2oTq3Cdk6i8tVdVpZe4
YxKntLReSR6wUMiDNAIZ2ZrTKkQ/VHG1H/Aoj6nrOdTtefj7tWRtDi8IbrQz2q+O
JJxY4WmU0jpUV9PBtX83KQmhiK0lNhXvSLZet1DUBT8bESEcw5Tl8EmejlBmGu8W
K/vScTQbxJIYhCiAa8l2HBN5yJffx0pM4tYQYnDntWLQNzjMwz8JAv6CIG3UKwph
h3JnXkDD89EEgCJRkaS4CKCPSua3oGLHfM8cZmPc7e4kQnr8tWZ4YS2su4ittmI+
DMST3v6Vajay2HAXN8Nj5cgTlgGx/SMtcuZI1y7LUQU0ybfwwXTj+jlwRYIwijJO
n7+k+HQuOBn2YXpGG6IYOEdvaaEtz7Ybkvg6KYRkBGC/6VIKZp/Be+aBsi9h4VQO
+odHp8L9MxRG43lHcSDcvDZBW7Zstok+cHz5aF/uNoEq9vIGrkAZ0avw7+oWCwcw
/oDNOJCjJ/NhiyVF5rBs7gelTFY/j0jh8jsPgUInSygnsG6vdnvKxvRWUyaPRdjJ
UBOoczyg/bG2Tco9DK7xHi5m5CaOhHMiEKTkktgn9o5Z8I9816vz1z+D1yUzn7Gh
oG3LUK47xOC29EUNJcpUY6gxbAPJVjr2E5l8SsartRPjcCUCWy6IwOv7zV2y2LT8
5SHM3e3wSr87VLAmON9+5T6ncbssPfK5tBuvO0erTXYRbvhW3OtImDx8ka6HFT0+
rDoZciiDNPxafFFHnw79wRH13GC24kd64ok9dVV/oM5MBdtrarOdqC96iNp6k2HM
4k7LJw24TiSg9MnFtm1AFoxCOyN8+KOu72IIPkpf3y5D95ut0MVVGIy0keVBR5Gh
/eCdHY8s1sKdcGkUbF0pUqHALdFFCQB8fhinPFnF5b29e2kESPiiwdQqx5QWMpaS
4cPmTL+Tr+JnBik32wEOCTFm+1oD69wUA67RPcXmZVfntzM8XtO9PjEyoe7zkfaC
3PUPUleRnT/ZTfD3E9Y/O2i1SZ28ff7YPQ2GR69xORYSj2vjwgfh8bejCMoZFLgz
ofTYpQ5mZqcA3GCGx+fn5tt8rPxbNBwtnsu7t15FEAuMW2gNTpf4h4KE2o/ioi2q
PUL4efFDhE975SVaytZ/j1lMOnZKMsXpk5DT1o2RD7z4OWoRnu5zrrMQwqLHhz2P
8zejkPqJajxOgltoCLMac8UrWEopXDHUBC2MU0GY4nsRFSTmNQK/4KmjaQHOAeMD
/LQuqcDBVvy/vUP7Nz3HxXtndueiCuGvSRLZwOGqM2uIlr+xWDveb2uijxAd1AE3
GoIQ2jZd9kc1l1W2u4iABKenLKHQm8KxMHS/JEEhSEhVJOb+hvQhQ6X9dzqQ2FYz
XTGsEgz6imJDBpgySsTHEyIpWWP2M9ACXsMbACWVrDVsM0lo6IAREWhGWdhnL1cv
nPGDtDEoBKJkp1W4+hbMuqbUBBe4FT6POCmFhUPByOmRKPni2euB4RVLlh+aWP2P
vXtEcF7iy6u9n1Vx7JuqOyzN/yjn56PAHUzsODc7slkbQJbZsc4HSOYKx+tCnsSe
FASChBayxJTop1TIl14V3vRq24m7cLF8QYAWOACmTi3dlQGRt1rGeUAJfUYalTGU
ooTAtievwdpKuVGrMNUQTGkTAos9TNR6Wmviqj3NJxMU0MtiC8ovUS4hrQ1XRYEw
N2MjANwNpQ1tozXkIbo2upqpd3aAuKdXppmrzUoPBK3e49RZoWT2Du/aH6CyJoaI
sz2ZLUNFPUlLkHGixOT2iMx9faSLeMkUP5a+mEWBht4gfjXRZBlV44mbryFaVhMu
bxpVvJ4ZgLhrDvNoDb/BqCadtWohCBn3den84qStD3q4wxA2SQn2GhhQIj6X1Mm4
TDHFTQsX5/1/nZBvZMrc4mSOET2v3DmWHMVkTrapX2PBXWzLonAPvXzakzHR0ysp
Cmdmr4e5DtcWHQZ7snV9cm6jRVpAzuf5rTbH4t6cal1OOiDh4u0Ntn009xPcUbZg
xXZYwScqGgvwseSVx5rv4dKeML3js/g+bRLk3Q/4Kg4YVr+R5w34JBALGXbfCNRR
SrIDdQFk5gJ/W2JzXp2nNZqSTGVJvmaBYZ0tGVG7ApVyj3UW0e4N4t0jSAHPb0u7
h5FEqdl12YPwi4MKGSrqJuqKzRVn/ffD7Iqfhun/u2bIZSH1yc1lcKVdeOQdwf5y
UjZdMU5Uu90X3K+uLzmjzDa640DgPGwcQkqvTkvFLtqEfIK8OGb6kCr1++ESxWRk
mSmOzXz39RllQRDS12dUnXpyXF8GKRDtzkYZ/Iqbb77rwMrAQy/4WGLLluk+62+9
uJmqEmH3ysoAW6MR9A0YE5jvqEkrWryDBZpPSotDZc9QQsIINnNlQLPh85WjBPyL
9XbSsYCsXw11TJxXVPfKdmLAX/+XleNqCw0ymuZviM2y0exKEbDVU8VrLnBFmlGP
uuYzO7b42bDJT/WZprBzGIW8aaLfO/tsVqGvXi6Mgy7Oo2iNoQDimjrSq8eK/937
eKJfByIuzr/+I6Jlzu/XS63vMGk9CjJ0Bxhh29OOd6CJaB3skT+NpKeizbosxrC/
XygqyG7Ij3SN5ylbfZ+uzATi9z+37UETo4GHNf6xzp+nPpWonRowGvCid33GuPvl
QVAElV5n9Y+NMpCfpPoTveTQuX7ZkMAwBoByTOVA32dVBhGTcTYNEUrkuOAoPaD0
xrABdycsMnmHWygtC8dlamN8COmSA9+z2vBUkUVpjrRLeJTy8nZ6D/qsGA4U5POc
wRYhI7oiSXeKBkv7qaUrnu2PUiAm3S7jA3VirIDPD74YX+1iH0KHNo+jK0R0NY4a
B/dUnL0ZO/40oTl66WzByRz58+M1ZutNHIy7nUlUVFk2ho5nZFOLgn30fdC1vslE
paOEBt4MpHsB4IU/jOVZ1fohIDqBRXjPOujJIg28WOTSOhDqLLVAyo9G99IFqtvX
+Y5eXy3Hhauek0/PJYGRJ005g3iaqYL+ynqkB52YBwombsFNtrBMPFrcxG7RgCl+
CFCZ7gJE+purgGn2Th44R6NU8RNaacb8LQPVVYQ8eYHN+k5zwleT426W9G4Woniv
LUHmwSambDFz5DA+/+eyFjmWWUJ8O1uNHTxcROMgfVSqnrQEY2zp6lgMG9TYbUDj
G7veJvq92NFECWiE25MADuw7H2sDbV4A4yHNKGtetoSIADUt4f70naoDFs5Cpjj7
VdUMcQcP3qzuHYBOvnZHWq8hUkoj1qZnNiXdeUFYVhH940bSObw9j+ieFXqMuXvG
mRo20AWZLoteTUvnGRUWcCQg9hpAzdReXdwjJdTCf/iRFCduHDC9ySDwRp9jN+ab
MsnmF+cuiQSPpQiKRKFdZP3OV0CJ8WOKXaTywah3r9wLkxtIz1yPeV+cjq5gA/0s
f9ma7Ij51eNRwNxi9HXWSU5y2/rE3tKefGACxJ+k3KHh3pRe1FN7P6MsKZ8nwlOb
TtHTkZM5PRk6Y0dCe2rtuYnptsorJUqSDzX3oMUjnB3BACISd+tTvhCcvY3pCGk3
nsZ76gEkbZkQYUXM2XNizdjAu8QakH9TGKQ8nBYschc4f57Af0HvmnlMVVTEgr4T
wQnqJ5oYdHE2vazA8WLn6JeW3vEdQ/BZa9FNmhU+tZ4F+fS6WGXZK5FYdp1k1tzH
DnOmpuQ3QMctUrFXOCTqQHZpAMDaMbSrTl4vLB6qFAqXbXRLEzbCnRjJpgMxY87E
Ctxnszt+i6YocP3su1j9iWrE7KXHxoOgo8zOTRe2T4POCKtYGUj3i1ZOKcIN30u/
FE9pAYFEWBFvAdWhskX9wtbSwxXObHN5uL7m2hKtccsy36GG0sUp63F8YyxiUYYM
YoLKdn4cgPvAIXy62qBX+B/Em6fhEA/OEnmcxuSp2hMDotouWhKb9pWUCWrGXEFB
RCYDqhUs66EMx7kKKa90n5/bSQulLIgsyDR3QEYfFV3srZHMQDSh6F8x+Y9BKXQw
Mrj2D7h6kRLz0uA9ord2LfH4aCpY63V8TGYicSZdzKzXNbESy/yeCOf+PVTMFtN8
i1SetX2TVLT+/L/kF5aTY7rW6LMcDqqVY5dw+wZXIR7p/I3atk/KYw3Kq0qgBZuG
YP3MLhE781W50MshlYSmYNn4qBw/013dSs12zbZlytXZeJNSTw6tMn+JfFRL0REA
6tukcBvyM5r/dVqH8BTXZYB4S1kTaQS7XGED1B+TuimBXaJz6jmXgB9CWTTTgS75
v3yUr3cP3abZaZgffaBwq72R6ygGTtx4Jy2udsu2sDPCSvl9lOwdlcYTAHpp6UFq
eMjeHVUHkYSyurwtZMFyHPLSyrkkNDCGgRMt0I+dtoe6Tex1OJ7RywnZ+ZyneHrr
kna2v6kkSeNyKe4TJECxJBk7tg2ROaed/e5MwqKxOym6k5tO/hlUtnrEY9fryk0k
xLKF2LEh63Ymp18Xr8wK5zmyV9XwA1ywLTlswaqJ4fj+YgNOUuLx7hoRlxyg+GWR
mtF03mQNat5ucRx3RDC8t/m4q+lOkxv1hCD0BXZtdzhS7mMDRdhoa/19S50eD2YP
raa2gRgSAgAw//iYk2JBcav6rHvnGkux5/i1RjFf4VpOpZSj6oP1a4kut25YIKA6
LJd5W/m2ZU9Q5dk+toQEVAL8kcIzqNPWo0Dg4715yPWfbWD6KBMjGF3NZ9SSJhSO
8G6f5LG0U60x2taJnSTdJjakb/BH2bGDU5XqR+ErxYuJrAjoYD1rqE4HFg7R2PHe
B3NUvYy/JChX1bE9pX1N5+vv6vJlPPCWGxKSGUnMNe9gp9K0I5rcRxV7PfV3hEak
mhNWxeSvXzhb9B9A5jjwc/BwjuKQhepoGWrsvbHh6dmduqKsYuef0B8PIGFDGpQc
4r00EfuAE65pVDYqBaaQ4EM4os5ocDUaWaIZKRyJ86oXCPimkcGNtBL8z1xJhYaM
Z7PLxZslrmSXWuzkhP3SFcC7vdlb9CoRM3k1JwiGDgnHvIySOyZYCxXp2KQS8Y4A
azcQrbXrJk+SUoCmEUvPhwCYPi06HGG7r03h/xY3KSrZqdJ7v3Vmatf7EN/gbN+b
C87CXL98f9+a21Jnsz3ipBePtqkWS5RRrMcfhZwPXbofoONncsT8r/nANMbI5tKJ
5PSpDumKc5MKjjK9XKrEUo2cPgDYoBwgScBa5TAwiSt0fZh+abQpTbT3hveXq6Sc
z1X9S74pq9FTUrvb6l7izoSEwiEiL372ZkfNrftVlY1cQ9RsOhSEw3v9xqyZwHFU
dADujcAGp8ExBMLND9z0Vd0hAvZ8f+MFeCO3a9UQ7Hh8WkQjFcLZYOZ+T2cxs69O
H3DvCfGGzCpL2BHciOgOR6ugXVjQotFx36HUt7Y0EQ3d/YErfyOWwrMSj5ZVSLBR
XJErXay3Vk8aIRMsgpvHRLL2P8f5pixB649098ZEe7Dnx5yoyAW1P6FKgTJA6NRL
FuiHmwmjrqK8YkjUahrDUnHh8XaUPN7/WmquLuyWUpxukAJsKBwonDbdn19yWWnc
+LyxAflQBm3En3YX+FrqrIMWIgzZKqZ3CPTj9/kc9lPWBfwXSr2InTyRgkiMB47D
ARaujYOYmcHYrRwtxOOFYgdTSJvpQ3IUJm6gdiGb4YujPSFVR+l8eCtc6UeYsW5o
s6b0vIDTFaVJUAoT+keSBup/YBD/2RY7QRRRWYI/NKjBSaVPWXzQNZgH+6ijsjCs
Wdt3I1JkB2dwvUd2nYsKPfS8j40r1veBlV9v6/oX/OJaORt1wTpvb3UXxJnUj37g
QLHiBw2TkCkZLiyUm6jhm7Vf/h76SvB45HR4qM8LsfCqLxziQ6FaGAy6/hnCONik
P5T1bYnVibjPt+rPF3XhayF8DeCBtQ1zGpvRCc+nmuO82VKqxfzgn6u5XUv89Kr+
H0ZPfzy5EiP2E6w0aXBpP8IUUHM2Dr8l/N/rqaOWyDYLAxCS2Nhhio6JTB0PbyOa
MsIsfd9g4xPRdADELVlz2Ncdu1UCbBht42sIXfpmAygRqoAke7VbdvEFJbF/u2HQ
v4fu3ZMEU3NVEgs9pIag5BapLzIhzB/iAwBaqYJuDoGpZTr8F80hoSR+OOvQEWhm
Znb1nU4v+gLMJy3Wbqm3NkPtVULexX+h25YhU3GdS3WdanBlcSFoEWqI8IB7NM9L
0nVmhx92Lo0ksHKYsRIVAYbXxvSD/NpbCpGa5pOce7u/bxbaHVQsLGDwLqg1pt3K
oBeVtq3uvgyvTNOALWT/7G7G6SCdwtfuOAd9pIX06xnb3vxUsgtyyVnCOQo/IfeA
dav1kIv2CWBFFe1sPh0XO/Ob2JMJEELdmXS2wPjbM2ioPqN5G1XldbZcCRKuD0hI
SI/C3EEORIjObwngS9gk4n8DvdI0Jx1hsG/wrbvNVk+u/pqDz1p/+1yZQsukLnhJ
+pZ/+Kfq6UXnRectHGvc8jTtOMkLv8dYB5tAQSwja5QgnmtTft8g5YFUsZEIMfZD
c+iw7gUAiFFGHRSOBXbsZB6zJw1v4qSbay42/qVtWPAf4YApPnRKZTLqmqcfT+0S
MAexsZ848JSOB/DGtUhlxARgjCIZnmsLlMPxDpdte4vrTAqf0+KD70NzYVAsJ37S
TicjLUPnQAqnAqiAN+t1w8guDp3kHYGnyWwsvEZjTiZMRBorLPvZxW0lVor1VINw
ykuPEbXh+dp+wcXEjeYcSu9g175Om8t68S/WOJ9MfruhxS0pgFn7LvgdQr0QxJpX
jQkromogbpuy+/iKHmqmIYvp47O5/Qrqhq1E172uNFl5mLfNVtI5bEu07nOP/3qW
zRye/uDAC9d1LZK99b6wEg7nnXsy3yC/ZLc9MxXBVTHEk1n+e9DzP7d8i06BlS3S
1dpPx/pjxc5WMaZIrZMOw5xWBwesA11NpEd3hKRh6VGRSpHukoUuijKXgeWLRyxE
fso5vJYn4t9qm+iBx0dlMLxx/df8MJIGbNesu3YK3bvb0lsAb0OBUIoNp6WI28K6
8PDYC08QyIcYfQdeh35T9QGKlswhW1bDJqwCjdqLJQ3W80spSo443kmsV+F9aCmd
f0rcqa4S2d8vbV9peLUjsh8KQjw4X11/D0BQdiJgiYQ0Ez7puC0L4EW94igdmam4
X0/xNkv396qFq3NyB4HLnky9bXSXHBmhHYCsBz8mYMAsGVrYKMpGxGtr6gDD+bRQ
TxKN0bqrLEJL1Tp23iesQB5b70FKNUR4Sm85RPEf58Q0z0WUlMMc2qwqh4XUcX0M
kPviJMWLp0pd3reNCJkvIfGOqiE6j7T2ieGxdmxv/P0KW67Z9tidMGkpjq0jmr34
nNLV1NPB/47omUZrm9CGh5Xq9LiAMHJJETHi7qx9GQIwW2D83I443ZjQshvlwsYb
tgnEz+sc3/cvHUHH1fCOsAhgeJwF8b18Rugm3DDCbe9PMqM6mksFXPDkXxY5x1dK
rz2+GNrHeLPMaF66Tu/TuQ92znmzsveu1ElRUxh9jkx9sKMzYfTwrLhD6FHlIwo1
BxZ6hjRQ6yVTA+zUOnG8JVrhElAUXc36hWhlYfDSNGXvksN+kq5xHxl4Hjf3RTLi
2gjLZUOKYmMcbdNG1TGaIyOH5d6lpJ/brMNvYlOXfd4xbnC1mOuLmhLOQnMvNtOk
Ma/dru/Q+6lRsqPge4d7EBYi/6yfaNNrJq6FnMiKk5mR9NYBrEuUd/1P8SgYtYxo
EDYMDTGmTNCT8smOU1aMXzZt0n0DrP9oxNsdKs/JRpRI/lEIrRuYdhZBp5yckEq6
ETtrO3Cnp/n4gRTx0pUeR0ZFfZPOgoa3gXlZdj2a4P8Y8E1BECa2ty5wzbkMs8gi
SMOkCJCio4oRxRc7tpqCniVAygC0drJWXbse/Gby9pPP9MpYn0peC+aIZvaMTLFX
KsfpB4oZhOsW5geUh8saeqJ/RFXLeTfwkHce3ROaB4HZNFrSW7kg8d8qs0kPG+kP
yRQEPILnx9SbZ2Fmi2b+tg4sCBU8/fuitFXzG+5ryVK/L6sPVpAedoM4t78YTVJP
B9xkGXO6OJ3A7l33X44dAhhkDdAsaqgg3qasxkvcTfQmcJ7Fxm009PT5H2SJkk21
BAQWplxJitUIDypSjr9Dhe7KrCjZGZseAY/c1U4swPBByUo6c30ulYQICuCVs6tv
6QlViN7x02K5qVZek/NguTMWms9dckQs9iePTrVF3s47JcGgui075ETX0IG5Jz+Q
fNXBQvfhG3GQ9UmZNw65hXggsRCR3I5QT85SWIzzNVh5DOavgNqXEC9qApXSaIZF
20bDD4gkw7oz3fNB19pHM1Qc1vmnsNcMS/wbIlA6+bfu0LE2gQZ1cjIVzFXyPPaR
tpRY09y8dj2baZFN8z+Wzd44/l/9TW7L5LP6fN3r5QwhMT4VJ2U0i86YG89lgtaQ
rQ8oDITNyBofqcCo/yzIt10G7uElMMqeG4LYJNQvcO3zdu5a4g8DEwbGJL4PZrbG
iH3m56gQFUfJoazCGTeRDBD6Si3UnHWnEAn9v8d5uYBWu5BwrXQfWqsfj5jQpVSg
4dxqD8sYpoSaq3dEvjagXoKwsNdkSYXjROwGIZQJSlcmt2MCoY8gQxwF39eCvaeL
rP90m5wuXwcCNxD7UwN6wbnQS1S/+TujEQW4Jg2QWgbB6mUxtXNp57Lmw9txVH0Z
Qw4Nib1uoX9e4K0mkNC1koIFkS56SIiSIMi6j5QLK1mQyTUoeHdmD3jtwsfzMcVK
8RPJqZoos6pQvQB4QQBdgKQ2XYUaox3lS7j6lf8bdFCFU5qHfi1zQ2fkNnDi1phr
lg89fSY8VWB1T2+/5mQWYIh6cCzsWVYu42hXRDHGrE0wipwhHHEsAR4QTlWwjW9H
vjUa/FdvK9XOt7duv0+f69vv70If4rNwp/JTUrxgaYE3AaS2bHsRSiAF2iO3U4og
2HoANqjLivDZwi7AsH2HAlFfAyqV/ZIY7ioNVFzfgjmnc2prYbOfSwqSD5iiqGpB
uqKoEMJLrsu7WWCffrTsNEcZHZ/o/n534gcRdrrlQo6wOOZ6TTijKiXj1wbnqk7D
TQf6FkBaPVh1IVIkoyp9eAf9LOxmzOrPHDEriI4EnDJTAc1hFVB/0SjqptzGGkXh
5Oik4Lsb98hPINuHzHhLuL4jO32NJAmq550fqdrrTBzJ1TfH12/GRmTdQ0ihbFIP
pdrRXiVGm91SXJvwc/9fLOJGKs4mvU0ssTh4vlBVZeWIL5rn7e1crQEEGlBl/tDQ
AFjj3iTHzMSqHHZ4uqRUMTrASUpnWy+TKJU0SjeOpK3JSjz3PYbuBPGHSXiKxiAQ
LGBpg6chrNpR4OH/aU0xs7mBvlq/JXZFehzX8JbqszTWxYe3ELgVTFudRKizfzxP
UbGk80YWrilrIHk9KGWFL9MsDdifmr0HQu4+UiE3oIgbj5Rhla/Li2dco+SmfMh+
VEh59fRNJX8j7q42TK1Zcw9H6p9I9x+cVSrEXDR87BPfNQG6iFMx3dTMdzBDI9Ai
p0ojkboeQ/5K9Ki7YGtHi56uztUHvE+si6WiF0wN/ePAvHXDfp2XFH0uV27exfPz
TtjH4MnwlC/i1fxN0KiBUt3Tjr741tLX7rELjIG5St+i2xd91QolWw9qxKYB8itH
EvSN7wcXUfnFK31NClmDncFdKLJ8WAc2DDeuU/omsu7TlGDdJxH15vTZGEvk8RmU
FAkK93wE+ZOvKGjGrwrvqu2RfMOynhadlfDbU+LlJV3JyJSbpHwegQc3bkq9QK7P
bGfb58J2SQT6wFLgejh3E1ofokxTD7A9k21A/zY+s7Ioz8o+CUOk2Hfg09klIkG9
hUq9Rd28xU8iEs+8ZvDCEDMnhyyvzjmnRfLbrn3Uzls3WdTN26smJM07u/3QyxEk
XmLN+jpZ5/kY6G/8Dw6RHmnVeTP9IjZdHyO1aILzHw6vg3MA5FOt4ioyTh672vo4
LH9dA/jQaijpLmF2oKeb6gVjFDyPlY4qRt4SWGUTw0RihMAT1IMyPg5gCYHnnApw
K6m6ck4C2SgrSPJmtf8i1kXbnjj4PmBK1EbSLZgrB7HIxtHdiDHT5j0bHASqUzeT
JsHpTOzEufvU2v/WP2YwISjtV5mVwp13h4w0k0O0hsuTk/0FvtRzufZOAF2Mgt9w
HY7/lcFYR6yGq1oadpA5k33Y0oxhS5XfssE3h21/DfqeZOn+V/3MH8sGv8/61Xxc
7UklYC5vWf1yHaKAGHj0rY2636FjClYQ/5x9uOpKSM3wiDdQAmRlQNkP0/NeUUXF
hhZzu78b+Xw0FV5qcYeSou1yL9L67QjZnapHHHywWM96JAvC7l1DMHLd0y6RhX38
DAcBqn6Dkr8z4tRLQUwTN5dmj/dnnaIXW5s4rXiEHTZ0hgiAdjm52F63J+nkV/jb
QDuMPl3XNvlEZ+vJfE7fi+M7h1NWv5QsVvIBXORrSE/rYesa5V5YXubfI5Z6iEep
/Vel6P0QbC6Udc+2HzDXd8rtKahMDjhdiEBu1KTUUPRf8ZBszIfJWYKQsJq8filB
+y3sS/MiZ7QuteDUw9WLPCCLbXPw+Y4m/8IN8HstkL8UCjBzXEzTBsJT+IDXM6XD
6H4Zw2WBMgFkKSF9ta4N1+Wn4aqxSwyKOWE2HbmOKaolzeTwXPja5q3S+tEG4aWX
BQ9r42uqnVqgBwbilh/a0zPBdGwnPTWxbQn8gNIegX9sQNzrDHqFauP2LV1Tlxuh
VQ3UrhNll75gdqdbdwcsLm/NoOlDaJSHsx4Ulo3Wwb5EbRf9gNX9Odp9kqU2wHCj
oEskyH5VxFc/w7jG1SXDyILwEf9EoJ9UbCM0oCVBsMTRDZ5FuUJXITB5pvrecOPw
S/3ZDY87xH26Ii1dLDWiqIEh88iYZI70l/JhrNVKI/aUcARaBei+8h9AIWv+kRtJ
N3Za+5RnW6W+ujB2hdZAjDVn4LYhnD9UrCU45eFdis9KrRANf8e09+Tzz59SDZs1
ZMI/hIe2sKX14OyGupAzCAcP2ZM8ZCTu7q3Q19GO6TvZwhFX3ryN+XMtU3apSgrT
NbiQ0sRT9aQQ5LNznknrZMtl/HOPSU0W321fm0NMJlX8guZXiSRUuz/JgCHL9xNH
OLjI+Cg7SmEg00RFBBhpLGbvI4Q8VXeiBLEA7oPGHKW8lhSRO4qAFlDb/+PG5OeE
r9GJh6qDL1ykPVa/og2pNWzQm2FcADzj2xxoX9pwd6UY+Axk0f/FS8ld/qRiuIuE
zDV43JwVd6EAqVo5MqbpNWzBoT5YIo/71fdzm8B49931/O4CZykWvxryMx7ezV2q
GBLyQVKLjVVTkTy089MVsa6R/rfcBRKGkQ2L1ApR8S2vBJNj/RSS1s9HcuQenbII
aKPvlX6zdN77LYtGOi1hVyUWtcX6KedyPat6srVzSdTHjsqRoKGDesaTwMkFFAKp
4i/epnkkARYO3772/jW2VdEWAuKBxaCodTL9of17TNSQnbdu0yiIPkjxb23ohiVb
ZmK5LWHM70dnSrcaVMScOTqQO+ulpdvdGQqhKFUwg/8eOoC9llL9UehcILNOtFZ7
iXzYn2OrWQEv+u+LI6bP1XXOCzlgnAu9sMv+WLjPiAeB8YNWa1ZWsNllwrmCfnlj
VpQauPWL7yGsyvN/5EdBkCHt587uMjHTZzbS0hDYqbzB4xPnn3s/UBB6OkItPn6/
h8ibBQgBdhMPfgE/ZznZwauvFOtev1K+7yvzNFDigMf04zBg0TGASwCBaRFhX7zs
SYKBlW9m6FVmGogj0YBKmFFSCTSiXzNOTuD0FU40CicG95X7L5vRyGph3VJJnFzl
qsAOoEWBqUYaSPwCXPtEBQxq4nrWFI9LtySaQauSzQAQDPF8gzd47KNhWQ9EAQ5y
hUB3OpnJIE8WCdPpKWBhO0zebehUEEvgCuwaqy/y5hJ16u+2NqHsWLfFFqDKto2F
W833ZlWGqFsa/fbIvfjgZPLqswLtqk5c501kjjbK4uE67qlC0FkBZvVkWRjwnjoN
XCKGNGE51hxQo18QKXlTOQgSqrqHsvA6h56tVni6tR8tFbDJAwkrgEugOPSkvt5E
kBA2RVqb7ce/lDRnCLzi5yz0UAt/X/ACzjNQVIItJ10UefgyCri4F8ltMbEIMkS4
GFGgzt+WwCmtEeM452FQgUJfoxwAjd4KTGoWUmR0/xdMp9wqaD696s3nu4btQcaM
u9bn3vWVsYIV+gtHjzwZXPEDOhWeqRI871SmKaJRcDqw9Xm0krk8JNEs5OhZaAX9
yKGrcuxx3qtVa7JD27ePpdYek7U/WLhvP9ZdHZACQ8Ln+Jloau2koJDlkgGGXdDq
LUEg6EJ4kTyk+xkySElDOYjOvQLHpeNjYSO4j8bAewByoQ+BZX4VFZUWUSDTrOsn
K40QBjfjIndgK6ZPD9bRGn559yXHgaXws6cVEkzoIKtwPeX7hlTsntb8zKyAlmEc
R1lQ4opjipRyZWD5iXbz+DKgdeZB2TAJX/oyh/oGV/LM+Eo/+AvTHjU0H1Ai9Jfy
USVXjQy211jjA3P0k6Par6P5C3ygZakap7vSHfEORaF3CUTZaoAt08CkThg76rJz
s8QrYdDMz3bT/9vJ5b4mmFXifGz+XRvYBCl5r/Q2bGsZpsilrhxf78h6a7Lh9wg9
LAn1l9+sOCv1oEorQiEiYTt6TC4kSZ/baBtdguJvJjo56HnUgxj0rbzsagRpxh5M
77ljtgVjfxpBrSaQZFxu+NASclxfA3WBrYyij/Z7m/XKJH8XLRCjHJK2z//yNng+
QuBO3WWqmyMYZKmRwZKVeZJTwBQJlJmRMbfzdyHkmCeBlJRQXvDbEuKmZaTyg/uV
O5XYIgGNc1lx33Ke825o1rmFFSJiW16Vq5QESPIBv6nZ6VINlqTAV6ekVE5pQaXb
nBKpdvXxm8QOnwvXbc8YN+0toLNJsYDkSwNacT8LV6xkvdasj159ns4rhWQu5Vp3
LlQqMmovPRPrUrLVHfndgFRh1b42niMXO2/rx0m8F891Q2gZXisMKWsoBiA5KxXw
Dp8hkVybMTfjx7QaxTM4dOnjurteQyxFsOSEQ3/iBfCPLPMPzre6MnLaRUViQ4AH
oSN5VpZJSMaEUN8ZEzBlWrK06GAIzlDNXkuDrxJbz859ZGEUumSkOX9/P7Do/h1E
IOiPNuvRYTIyCn6e2nGsYT0rW37xTWFOk7vFEt4VRyhGKq1YvvcJkU5//0y6RURT
dT5YPKxH9Wy6Gl5mHTxscbuW5vshI9VW14SceE9p8IhoQs96YwZqH4mTJaItHHWi
PVxtYx2nqTwspSwvArPOIiuxfEgm5eXMNGh798rFHSI6p5Lua3WUfU7tBj+GVfPp
jHWTvzAvdKk1rMIb5ctfqL85X8boRDRwAfGqojBQ7/2JhGenLqS8EkLNKT5BsWYQ
lhsyAqSKwk2EHHw9vT7eDdyp4PFK21HOcFdQmDI/xQpgjQqYjVucZ73Kwv/V/l8/
8FtEe4qfUTf+S2t1y3c+gAJSv0GYmbPZNwJE34kmCoWr62ScybxtsxHJwCGEs7+D
yNpjY19AKooCtriBGnrMzeSWJZXcGjB4PukNPZX013azYeKtq8S1nxObkfBK3E6C
qVkecqP89f6Mz0Am3A9f1hTQhebX1eq70b59sj9HhYe2ZUjBIspTCTNiARO7ZvCo
uafegbsYnS0affaudpGZkd2qfDTrIzBpI3Ja5F2gErJNVBHRXLsN+l8DUsrFP99i
5e5jO4UkbaP9pPT5y0As1RUBlORp6OCbgwAOzVjRyZ67pEAeNgK/jDGHkF3VSw2j
MJG7xFlzATO5SK4TgNKJfsYH4fk/KFyqHvpt0yRkd+WO/en1kxH0cEXPzRpRi+Ey
ZgnVDz1mHLEP+t72stpaj296+tfESnxi29Z2MZ2KU+Xfkh3/ljKk8lDFYzk2WfTB
2CKd8PRbIvoeg7CYYKbX/RlpB9vYj1tKRkVgn04OGheBmbDNBOkRYPTaAuNxC7PR
lN0+UQ1JARWUfLh76hXnxfcOALzAds5zJBwYKrlCTgr2WedRtM8YjmDoKCDcwoBF
rNgCln7XYB16CS62fqK3SNMla5kr09unQDBguVC+fqbUdGzGOUZY/4/J7YZFwC83
3AG88wAvkRmnbrZV3bFZynI5GuKIB24Za70eU6qyLTvWMhJIlJvq2HggEgTqjJbV
EHAsuTQMjyd00C5Pv8mi9incJaPeCyha3le6t3L5I5PYpOoolCmWsyJqREd9WpMK
qNnAS9qVJmxrNuiEurAsYnR4NtjoehGXt8DrdJXOzlnjTmO+VgByD7sB+8tbt19B
LoYUTxJa9LtFJm6L27snSOPfNr1mbFhK5Yt5pgPUuDjZKicmwuB/9dvdvZDa792k
pL3lCb/EDETejQ56eTJ15T6P0m2jeXLZsNiiC4hEBARJfHz3aWgx1x3LWJwqAg9i
OYGN+kNj8DypJAYls5LbTakwIgirYq0XXlXOFO37S2v6dmCkn0uQjD0GPZ/LGj92
cN1XmU/m8aFTjBuF5S3IzAWyFoE5KrAeJ78dEo8RE5kGM4xH+C4r6TwS9gumt7pm
WkH67CYl1AGlu74QHjDTpBCflKUnCXOLTfXt342+PMs/D4L4TecJdcL25WqFkbp0
SwMVkAM0inmP7Ep09d4riNtF+xa1DkwPHwaOs31fXF8rCGxjHxT/eFaNpnUoaiL5
vtFxSDNQqQOwiT3eH1yMyZ/1o2aX3Iu7rQGD81m2qXoFN0MCdvOnaoa/xaKqbc7F
lz4Qsxy9fX8/vnwG7EQi1wNItOwEO8zH4afxa5FQTc1q+azF3BCDftVhXFmRelWo
YFzA0iwTgbLrPViuEkp630Tzvl7ZkDwsmsChdTt0t3XGAjp8inexfql01rhz39Kb
m3Az62a//DSKBouBxREsNOO3rDwlC3c+3dO54O2/8ph4E/FTHFRgGfn/2tQYD2t/
qjRv/xBCe4fY06HDAWU56i/roi0CwydpAE6FjcmCv+IcfyKfH7/eWwYf1PEeQFGw
0K3Bwv4PrCmEE9I8W7yHetqLfBsku8nJZXW71A8+HmNLn1BftZ+mYbeX4XD32aO/
DnWQp8zf7YqlTJ6iRhLve37JbCGjl6gKlOfzbkvZ/qSVMt0JNHRheuSaJc4XE9Fy
/F+G3WzcI3xIa5nv+TEm+INTQgBHcu7TbpqqXQ7dLJ7zgvjxtdjNkS9LN0q0Vie1
54+vwL8KmBNwXFUgtsiGsthDYTmcdavsScRTGcZL8ePfUq4V4MvF0SXTnoKRPCgb
mxs1baeS2WPJ8Q+u2lD3WDPKH7P4wULMNfn9rUfBq7+qzqCRO0FWmESvrUnz637y
mfTquK7fVIIuxw9IH6mm0pQXJFpo8QPqDkmJiHPx3Cn/h+iU915qi7M4IJid2SGu
+oDLq0psAfhG5+SjhhVy653LeoM9TicE2jWZ/xJKr98CbKaB7bcEGLYktKKEWB7Y
WHRtN3g7ZFBswwEKU2sjdz93eqyTaEf9saKNhpS65tUOEBZVqNArO3YI5GVwYBMZ
q+N7Cuosj1VrbVagYzsvJymfb3CwMfFwUlTUYVjdMDIaIEqhI6xoIjscA7b7QrfH
stsMiLdxvpE+pCLQz8xYu+T4QITcdlcg9dySn3DjMS7u2Dk87Ih5mCssydAd8Gnt
0/ADAtaJPGEepEe2O8gD43qQRRinVWSSqwsjRA2XBoxBaPMNwuKl9NP68GWpWrxP
2+O7dNEqCKu56lu3VG8ujkpc+oFYdI/WpDRRQpKo8JDBbfsUZ3WQuhYX8DVsE8gt
+hNd0DLQAxngFb1LER0IJYhlDgTDilPBaQo2ZkZFCUDkGXoDYjlH2t7dVLvhvXKi
3vm1oUjBg0zU4PGZRfyAdlIZ4nqdvITZ13UOW6PUFLZVmUhfn1zjKE6joLXWEwkL
3urY+o+/EkVlvdM9DIpFLGfWjNlPNCTRjzd9UT4r/ivYNZ6GHowANaFe6LUWYBhO
avPlJ1A1QfOfSkV5d6ZOTPdh1oYhRoEl5C0P7aQwXAwfpVsEwHEmQAAzC2dUZS3Z
Co1gcrHxNJP4/HyZEBfb4o8ibJh75GV3fbDywqnsP9kDXQW0A4Xi4mCQzintGc+c
oepAqmYzGrn6Q7GH3chMqjj/6WWBSKAjunqRe+kdawnDVGT/glmUkRDTW8DJF6DG
qujWQmhYMoP2+FYlxhDTnALtAZeMSeSdhfR8n2L7dAP6Jp294Np86GCKE8Z/js3K
JPpadxWSk+pkjOHs1czizJsESDq2i7esRkVNFd5vesxLzGj+0G0BoGKa3kXyBkY9
qDXHCdjHmohnpMG7Wmpq0i3ugoXhb/2XX9BbYGJCLkNzJZA/bf1Ex6lO0sltxUXV
KEec3fpz9R/6xGtn4pCLTspFl8SmujRZaEZ4XFs5hiKlip5gyVksuhpGLaeAKk6A
rBnVw19QdsPw5f0TQsUmrZhSuMiCzY3oT/rF66ioqxWklUSFl5BZJtumNyuOlZQe
M5ME3Cmj2g077YsliRrz0Mr75UL9vsjM4SNzv6JJqJmPOps270qqWnVUbt2QHrUG
RA+IGibmAUyEIbAnXCI112A02y8AJlYSifKli26E8Xmllh4pxmBrAyiGnpE+iVG4
/2IwYaKRCHAEb6aHeC0TZNlWmCDEgim0l6HsG7eThNcyqrI9+PuPrc5nyaSPtX5j
FAm8K/hWj2n4+xvGx3L/YQzE6z6i44Fqa3XQnRmyZbqkXCM1vIFAWJ8sunRpqEPL
19p9NVF+HWsVNO5AFbaLa+TMc/LPb6ZoCoYUs1qiV0fITJTEqnE31e5esMoA5Avj
gl7mMvrT2a8ZBgyzdZ3+mlKGOYpHBqp+v8OR/fvMAp5iR/xu5g+ZCTInWD8Ah6xW
1100/N75EiezBTqKaxyMyH4lta3Mwd6bd6cvka+D+lGCcco+olIubGWA8mGoVtbE
HXIQnHlox2ur7YAZg/98BA2AIzpYfzoOzw3fMGQAQFxAufU93s5kQmfMeODcTDpc
T1G6zIG9c8Gy0M9VZ4xG79kZojFmKNG4XPjJcEAhdKYG4O4f7BtK5EjijbR6+JE4
UmXkxY1pU2lYuSGHbcucc3ARdEpzTV36KVewV5UI0rfpaSKHmcQac3LTsUYrEf9c
pfumja06T3FnK9IgHJtY6TEvmr65fei7mtt74U/8tmeZvYBeqqbcamMw7UC/Yivc
p194Bou/AeySWx6Qgzffarhx/WvuOspG+4+zL5VcDTW0ENxDIZUe/wqCifL5bE5q
SYeMdlFmLRbfd/IZXOG0LVQvonftq6WyMDwbO6lakf+JpHlfI9n6w0NtDIxNgj6F
KawbvA4wHwfNOaARh5L//SUONKUJGDGTfDhTh4gIiQliQwINARHhOebwBY8WQQ9T
kLuCfLwZYIEfgO0KLmKWdvLQbGU4mgx7A3GcAkKULYJteg0lnAIejGN56gXYaUEh
EalwFluFcr3tP2V9tyq3zwpt+fSnNa2beNhX+pX2btOV/xa+WEMLMcXjPPGrHXRM
J+qcfcYSHfvQwMkB2rI1XfwVm11RVkI01GIyb+fjKELab/8s0amPX1zNdBFdElja
i5itxsG3FjPa2DQRhrPbkJtXXfFN2dbf0mxeOr5LljHiGVNiQlx8zuJV7eV0WtkN
yFH5Tu9f2OrITgzhmPtcTXDfnAfOYyoGxs1Gj0/AKw/iTxyis8MmRVMUY9xhv1El
7gacbse2D6HqpbzPXTuZzyr/k9jEHcO+0noWfyAQAVN/p2lB+fqeICf4+sM18Va5
p8KYgPxE3aLKm/UoFwy8OjaxoQqw1SdXZ16TP+XJOBcOBRWyt4YVnzXEAnv8+KEC
90VcgBXFiBV0y6B5IKSk1T9WDiRL79JGZD6he0ET8f5HANWkOYU+08qj4vnMJVwA
51vaW0OkBmNmET+JrS1hplVZcAx66w5A0G/rVXKT6FJNEG9NxfAymzjnD/o1nTvm
muC7rajvBTOG4xcbZncHYNIMJi3n6VTD6dJ9oL0Gt13YYJZuZQrJeJ/RAzXKxow0
lEuoKc1+bqrpvb7r7BKv5wjL2VugCHTi54yZthR3TUjppzmaFYGLfLmrBSzivpdQ
waWfaS9pbqT1e+spGvv3JneEJP17UbktDjBFaE01Lquk58SNGUFdmGT3SiuH0r9d
wQTd3Vu4MPMFacspigICoH3BDixo/OKhnDylQMeoeTWXDfuDEIV5+JO9rEq2PNEt
q21EslUvgAD82yL41KPlTzgRjK8G1IgwHF4GgR23T7nTV6Cj8mCv5SaLfPjGFpi4
HhBEIZfdPjAY5D9vfbwlUO742pnCeLHUJ/e/vYw9Vx14EHcxzugwggn2mXRjpMF0
8Dm4wQdPh3HJsatt37azXxMka0OwCpbTcBzsn86lzyyo4qAJh+/KAhRYk2SNvsGM
EaClxNtjEnbE+RB6lkPWys1L4EW8wX7MCW2Z/GEIzumA0g6qEUXFMunzc7NquuAV
3dqzhpnmFxBLCf6REL/2vT68c4kD/ECUuyGTNWFCPbRP5fUIMKO0sZ8SPQnvLJvr
IcF/dXfAC+wd5YXc2hjrl5QKmwpDcfME/TfbA8OUAQzPJSjELVhFE+JUe3IjZB9X
YGXha6/aLGVaEOTRnWBBPIKcWZj3LOc2Dp7p5To4J1YpO9E2SMnhu44sDAQ2esHF
iFNxvpcs+KaPN+7f3r92aWfvv0kxy45P73votUq8dJ0o65yp6jgmcb1FoS8+oj+7
nxxxZxpb1w3fPmUEs4VsxjpbAiBnW17gmH4gbRs8vRzXpCliyLfx346AZ5sMv9Im
OOA6tUz2/8Mn7FeA/wCQnhKAjQcWWPdzyPzJdm57/IiXD+K6Lm3Xc/I0XMhhGetD
WRCo2Pv4cy8bmjmlq7VLfGE4iC+S3M5F/mgKJ4ETYAqV7a+KR3/ita+GeuO0+VY1
H9uhtQdFEdlnes59WrpARIpECX4Q5HgjSsVljdkFfL7uJMW6EfQW8gaoeERlXaBy
pUG2h7kRmqDynZays2PbTj2fwK88d6qLVGb5Z+8r22HtYuFNaJ7ftV+MY1EXj2fv
6knJCHDb2J7KFB5bTq3nZx7jM6CEdKduju7Lt+pHxkpZHJ3CBkcYeVAlfFYCFTdw
ai8TMZ9O9N47K8SSTkFJI102/sOKCGAvqDGhguCj1ll7VDoojo+V4KGL+gbq6mWK
XTu7yHbBzYAR83j6KKZTfHfHsdM4HiAThz7GN3yP1hT8O1oJrMDM8vJfn77Rxcxx
a3oGsHShEwYJkXhNW1RE3531TkZTrVvqlOuZuhXQUP9Vx3nWdlhVUKHW/ffIXtld
y3R88cvB0AHm5AVMR3N8qe9UgSx8rDvkeIm/lcP5ZoQ0ko3IMjvFQQ8xtSDakprV
Kdut4eK337DFF1FmxcEzro+cfOdAJ7PeM2cBwjeRFNBF+GDKgDBN0+wQ+9wDuMzv
GLh2qI8i1Dw6IpuyCri+3sM5oZghHGYLejWhwMsAajEtTkF5iGROHIqo6gA9nbEa
fRsiFZX4onAtjqL0Rr2Zj00WO5j1HKNqxfHnQ3EpJm5s64VHx3hJqwCNXrE2YBUE
jXzrXhqmHJuhOKWz+3uSGVzJqrhzpDSwXaVvB+dx/TYK0bXzMYXjdTN3UnamwD2I
57GMVj64gocT4yteZd3tUHeNp5XmgmD4bj4Tdf2FpQula98ymX3jyVcDILvEfYyB
bTP8IX1TeiMWeayY1fbx/P3ZZW7WHmpBJYdguZpT5Vk+vOtcK9No42RlwmJfW/yr
c8OtjC57IyCIcSHvg6cBCdO3Zcv8jeT1JoJJLzxhJNDlXkpXnshnodS9lcqR8G63
fXzrOKs8tb2jUVBDWjTfdvjlDeo8j8bjTIcbUW0aX+zLodsMBhMmipLPwmoCzMQ+
NgqnqCzJu5HHCNpCLml3EBb//e3S0z8phsh8XqjpHxTKdCBIQGNf5ryziMjdMEow
Kx4PupO3M2q2um/3qRSPAasiVBiYzXFQWpbQ01t2l7QHIiqzDbJukBeOAMWOrDO0
sDjdBP6kJ/jU4ucRT9lACXoYTri4fcub4IS0rbU0a8gMXQ0OsftiPR+20QCXIuro
XRog/tJhqlQKR3QTFrGPc9941Bc7j3D/c44Ua453UK/ka43inpKzksgdILbZrbXE
grm8TP5Oo42KxetytBmuj7OCCVj3+tStkmCYS/7yDC4hZ0GJl8B1kc81MSaZaKWz
CThvTuLDwfQ0Y4OFUmw/7IJn2Ak6b4oUORNunVPNTE1bBWbOpLCZJ1u1U7sqMU1s
Z6+1h9Zk6FQRijB/avRTzEsH7EIYMA4LXcs0icIIUOxzC9LPGGoluOYg7pHWSrvQ
HjaCETWothjnfPqsUOcyDbrzYSxuM3fGuqakdfdAoaPLFEW3aWbgmeE5dar4+TLp
RmTlMKo9NTK0Lz4ZVpm64ioxs9gMR3wsYRwHMDb/vzKkPZg6DBPCMBXxQ0NUNcLo
1pCP9vqndmF+N9pilbAAVFc2nnTT21BfAC5j7JAzd5dIzB2qz8zvkbJ+Kid9l7TV
EVWblHcrfY+q+eVc8bQ6Gg7jXvkPHHRWxK2PxHxxl6bLw55D/+ZIX0f9+hN197ga
UoEyoZN9RyRfV0+Xl3b3g1jy5Lj8AUFkugHjrvPenRvTqPDuPu3AMLEiYSbBhLQv
t+XkmipQnXS4a4s2Vm/b8fUKWmW+Lz3nmUceoKKDkE7E4A5vltIck9rHesDcU80a
ibInKL+BwD/tGPzRLI3rSDYcPOE9mr3NHevXEmId/Z10Qf8fFM2Gh6bjwu1+MUxQ
G49AEi1qLBF1EB9kaQj6uiIgopNG8OHhribMDF8Q+osirLom6AhgZSUh203/Lppp
/fmbiAJlF6IdLLwvj3YzTDRAChaRgcQOifoTVH0CGRvXz4xEroppUp6CehpNMJtK
5AwgehAet2lyPkkE+0Sn9BkBsUIxou4VHtGsGBtF6XN+umIQE6oOeNNQjpmy3tid
oR94VAIA1aOueZ5fvchWIxHVz2Jhkbxzu+57DPqYcKd2VTsDUY4JorSEgbOcGOme
ROh67n4HKIKyOjuIcK2QxFbla0nKEPeC2d3jXlF6Xot4DJC6QF2j+esX3j5zafmW
GG3x53J9Rrwo/MFByfcC6sAWskkXwAFyQqmOLcUhiQmGNEeM9ndyzNnpRYa32TKR
/5Z4iLeD3dkK6HdRHPxbJfHC1dwTuuyMrYZVjXBc6fIFhrT92V+dCDg2tSjFXjWj
B2HCME95OlPG2pKNVM4UV2RrD2wZWg4y329HDVw5mkna7bMvXVUlLHxejBTHcP4B
Idd9C458GhJV+Ud/2XDiWjfCXdcwIYemAlWY8JCcrGEawWxvy/M4mkzYFlVL2cGZ
/j4VOatXS0yZNU7G55SVBpVdNXynRIEI6qgtkXURrGZ1dTAxX4GFUNxAxEeN87Rl
2ISb3T73hv6w+PVVkHo77zrAnDfHHgFN9FDr3s08lt4PoKM9m+wk0y/eCG9VuG9b
QtWSVHXOKuN1gyZ45XlqqoS8aDR6ZIzdI+Hb/eH9fvfH0oaDSCmPpzrBe4PYfQXS
SnreuMJsqROzh5bl7QRgCx3kkR00pmDkcC5n1S47yKlhzmxEKQjUnxBXTGUqSNDV
HKRgHuXHiQB07JlBlwiX4lL6tc2K1WLWJfiK/HM4guHiFAp688HoV9mRJuufhaaZ
RFjvD3HRNzjEuZtAwk0pB1NwasHububkX/h+RAD6W8RHDfTKD4K3+mbR8aQEM7MO
p210uhRAf6tF5sOavP0RvZVOfFLiVtJBdfrJObu+LuKRduoa8fdJvlnrQEUr5irH
a7CypVHNSaS23HcriN3XoPBTq0k+Mz0JCyZA+pi4q2RN3m77j1kJDTysB8+iv9Qw
H0mXfctlrBtxY6l7VgYwXTJ/uh6uBKMeKOATJImZ45eKO5ClhsBFp7SFOpwh131X
g+TI5I+a7uPgwId5p6fz/CPCLz6m5qzrqPl/Ak/i5hQlU5YIOIBtTfrrbW6yHa19
3xxKf+c5vVr/9Q+E3XjZ0UrM0++HRHIYKn5J5UoKZ7GZtoXrR22fysvpN+t5gY+C
AlAL7K979Eb3ETzr9VrsuRF8Hauh/W2lB9xUTFsW4ayjy/oGwh6mz16GuL8+RXV+
IqtCcymZVcqEW5F1r8ER+3/7rhhb8Mj39dglMzMZFbImMAXWgrHOKYoaD3ZnMKtW
xiBpUOKPkUaTTTQ5+5d8GUTb9MX/uUAkVpATvWgvkFUxNuDKvNyOzG7OesP0ucHO
zdaTKm6EpqDHG5rB9pfrhrsdnEodXKG60WSufe8Y708NJaReLC5fPVF09TszQUKc
smc0FARqFDCX8EkbsFq/BQ2DtZOxwuHs4szzY77otDqQWNghWmLn1H5RB/j28Gzj
yUyRwnF9Rfjd3HwJIMCGjDK90XZXWcS5Lrdn3/Tg984OyoJ1KHLuwDMCVfAA0Rmm
xxcqsn7LA44ea1mJrLClsvaFq6ceVAM7FiZjFUdPwmqlfx4aFiXs7qy0Foo9MY3S
dx+3CCtdBSQHtoTjvLZJHyuu21Rn128Zw1znLaZn1vOOF0By51BfS8Uik8EU3Wm+
wbByAPvfqrJab1I7q0d6C4niJqj7UuCVkwZCUzaQrvJ0vquVmgjcEjFltM30Rfzk
gBVSjWSyvLZYl6SZJhhQOIvbSWzogE/qwyFmGxqiCEAaxPInqzXHALJIYrLTy6Sy
o3KsVCaxUZFMVSLdyj7E/TfsEgQ0kn73EjraHZhpGjwVi4dBciFKI+RcnXyfzReN
MUGWVtFCjjWumN18Saxe1wsawjqxitHPAKSLLp27y4ckJyGrC0/EQkJndIav9+VB
C7TD+Revv4MApRVhP6rFB2WIxg10beasBaqANwNITEBtrqX+rNajLYr5F1M3nj62
0h92D/RnYhh9w0drH5072c64FIuL1y/K8eNek30hVDTirGK4kwIiEPeaTr5JqTHo
Drs2x2V/zikaBImUgonLTWq+dGWqIiBjnX2/EBhxqtmfGAcF0D61uAAjEbTKfQkn
DE4JLQlsklkxyhvHr+ZwesAdISuWMQ2WoRhYoBt5Pf/b8wL8Pq5EsErC0pdIxS+x
06NznT4Fjgt/05L4HHvu3640w9ukxZbdpmWxsuPYXJPNmx7GK5yL/+lJJ8HNvqvQ
pxy0SbHkQhW+kNNur5BAq0S6GcZosop+CgKXmGqmQfeZgO2d/a3096k0mc4JiTZI
MhyNV21a88Ed60KlPDZ6BlxA4Q8zjaDF0ghBCm6YNN+iNohc6eGYBLBdc1H1ozkW
Q+T4AeRdHqAwnw/1mOeuOcCyeuloWcbcW3siOVhmngcg0dIOkvtLodoEuiUkjSLg
U895ZCvPC4SkD+kLqZrNcaUkyD7Y87FzaLANsTG+925xSQzL1aKT8o8nH7LENrvI
BfqJjSVZ+f/pX0LD5rmjJfoctMNd9YpyAiVBhGb6pyVY+AnLWMeQdGjJ5rvomvf6
ExzCcYMaMsX+ZW2F7+okLvUz9WjlqLVK7jsqKfN4dbinQq+T1f/5Xv2NtPZ6+NDd
BlHvo2e0b1jHroj4j4sIxa0TwcYJi79hqu3v6MMKcCAN4wwtFMbj819RFpw0WBT1
RuYBBTQVbbaUMSa9s/bztyBJDwk72mV2MsKgkhFgG+RNDBS4Bwa9zroSis8aK0Jn
8SMA5eOUhimSPed4FM8a095+OcTXKMtnteq5LT1yay18ba4ZqGLD92kP1AOClUkU
1z7yMd+Yi336xfB8tvou++GbOly5ciQolf1o8LX56f6DpHolkWndTO4xbIUrzEhp
kB/xkLBk9DHeLpxmu7MWZloWZioWXq1vVXKlfg6I6fV5EBzDikruqzc5oALmnxlA
+oWUQvyFsuChAnPEgqj6t6LDt2xJpD74DSe8X2IjsF6MqpMqWrto/C5dCj7nIiBp
BS7woOiR2b7RG4o7zLAuDqCz+w2NGRdaB0zn8zmPd0A+GGc9Xho/eGHMV9QsLqCF
vCO/A0gkuBk04PiEAhmj72XryOyk9oOvTGah9E/ZQMlWy+sRBfwc4LHJUVWsABtI
UwQRa5E8ed4fmMaDtu40yM73ArO1s2Qxlk5WW+65Fi/yORvszjjGvAXJbxscjOo3
6Fhdli7aRzO/CwQBv0ZoA0zfkw/qmvqH05mWoOg2p+V2vHK7+KZBfAe98fPDC91X
U1mizETsBFBvyuVN5f55CwSLDLYvq8HvA11WHUqsacQK823dgLWx670ru2GH9Mc5
QtHmD27IeFKiiMqs05zXOs6ck4NRH9NCDTUdlu52s/jjHNM+3LRZx7ldN0Nqrvw9
xGuQ0Gku3re/x7sXgzMOuWKK88y/wAZDtWGn6fbFZa6KkUxxTkpsKty/R2047KDa
1teW79sURU+/BClp/TOELlT9SQttQbpfeLwxV0MhquT4XhhsYSpReONAf1GIwOoC
S/Gs2lbywAWA/yf57jtyetUo9naz03q5lwJPdAbr+wFOcDTzCtgCVqhzDfOgREan
+vXDRxb6fron/H3N0pYUkvoOVNXWYaXxj9eXPjfhzqxej/dlmElt4i9NRLGeNARw
n5d8PvDKbT+oU5xNjj53B9WHVt1Rvwn9SBxnsIcU+e1HI1nkEmH4Sm3l/U0hQ1ZM
1fD5YkT9C/vVvVtUBrvc/FNFwkbQ/Ub4GbKxOHaD82Xthlml7d5bBRaICnH3AXLI
WH2siIMcXYZ6k8sY1vn1NADIkrgVSYa95zBIQmc3FRG1fiPceiAyqUZRETRc1tSF
WmytaPe23atzTrkFa9HJy0SyhqqhjbYeXh3JLPnVYMECVDFehpmGFnp3LIO/E0L6
3l2jDo4tl8fbFIM10+shbrndWFthvo+pxS0BeDpa0qdMfuk2Ve5eh/eMTJRrPJJx
lmKEaoZ5i43Fh9DbiHRbx77gOzAdzY83570nFHQVjSs5rPSnQHufpmjM/+jW/imE
dz3sZMupoQqVSwLmJmAIoBjPjKssKT7Lq93dc/BwK+VUeZ1u7dhPF575mnrWY+07
CcFcIAz9W4ZZiOtINv2U9dfH0qv6ENu/mHyMsRsHvJIz5s4/xfyyK8RSnJUF3/WE
zlzIxX5zl57Tb5qYoed2FjSDQTY+sXsBTq4+aWJq94/p/hM/4cpdeHM2jX2IHJKB
j1d4JA+zW/ObH6lbMpGMHd25abTD3KsFU918VfqbpQIpSMT9ks6NNIrlj5indirA
sW0wvkDooorTjKieNWy4RaDHELSbve105x/z0a1jDI4Pc0RohyXbfzFsGbkHNqBn
kbIEziZcIbp8CHjXp5hcnI4qhy98XED/PAWgaTZY1L5j34FnAHMWxqAR8W/kapD5
o4PHUzc8OwBXhRLT+V7e9S5cih/1Nl3SkcNHU1nlVueM9IqLRLfKD26nqhW8CN5Q
SfI2ul/tbPP6q9TZcx90IlCA9hBqciqqo5sRxNYJuywNvtbqB0tZhQ1hXJOOuWxo
iWpUjOyD19grfup62CqphQBJxvvWhEjhH3nRYhDp7fY0apiCmoi3i8Srorjo3MK9
nm4FO4HrlcoRzsXtS4D3uR2/8CIczCrosOGYVamMv9DbFSQSsLw0yjJWn8Rvd2vE
mNTO5NFG3z5G7P8pv2JNvfqG2NNvFUpXLp6SVMDgvk27h2UZJG5CXRiCrXY6HroA
Uypp6G8pgjLCAKc2gc0a78x4IjlrGqnQ0P/WWruMhcf5ZWLkggZ8T9t7pk/BwQMB
Ak9fTCCbah65CB6FuT7HSM3TLjBj0EOct3Db1Ak/nxjUikR4ySBrb9AAUdeXAIYE
aDfbj7zBm3K1qUopVi+GOreBb+B2jdevDT6eO6BKrUTDx9R4RBO3N3aZ68gs4u7x
rygbq1lNNDd36/eZAtTi85VRmITA5fOFAVr+r8P1jh7BeHfyI9Q2XgDwYE856fmb
FaFvyIkFpLpDCpdZUVtizNVphmS8kjjkk63g/A25kq4RvR9oKVcVuM0N6hCLe5Wc
mPlcQW0a1iTnXlVpk83Jas7WPcdji79fmen78KKkgOyz7xxdsvsqFfySBVxbFRHZ
ft/TqT1RkMFUWbrnSopNjRMKthQZIjAQ7ihuBPX8Y+b6wwwn/Ac0N4tGr5AQEGMA
M0fXxXHfejyII3aZJQcko/jelQZrsJFVRXLRHeumSLpnI3eoskDqqo+Wro1JyBfn
w5+jEK6IBff0iH3OWBeuIEt7JLby5cA8en1u2bGSeZ2gFDvqIJu4/cQ35arWw048
SGXPkLj6wcSbt+xgu+fzPtCLhtLsQacJZ/kPRtdNDtPdKbdC6+wplH2OGin8zGxJ
2OI/CwjSNFudaF6H04TDQ0C5gxgeXU1J0EdRZIFnzks2T0eszz17Vky4k4PS5zAA
rz2fllAm525N03GReTyduguyZdROIUAibIsNbX45JEFbksAyoMJ3+nQq4pS2g9/Q
q9Erzfnyz43ULTUZRaoRjxev2fbXADrPFziOuklSUE+V8EFnwGOqh4hbQ2TC+GnA
2Iysqut1yckOYamowSuN0Txo4UQPzccwuqHtUAak38HXh9Wtrtpel0Wv8EKF/yz8
YPd/6wDY66+MJUOg+pmTuxP7pyoox6bU+nP+11Tu9HpvuNhDrU1r4GVTA2CZwWOT
U549QpcLB3WV8layece7gyVXBRswuFTkd32NB3Xyud7MW3N/5FCNw6lLejkfzxDh
PDOTf1paYIPdq5BbZIRHSgMggAdGwdjfWNUOD0OxIGNGnBAiGewo1icZ8SEhrnXF
oH+8Q7OUKrEf1JniaxJOVu2j6G6kbj3Z9FtlpoPzYeWV9m9JwY2V12eg6eEqlrtD
ZW/66A4cTatZMa/BVs803T4vxvY6i2fZclM16FW07rUfVvW9qFRJeYdq9ainkzKf
pegeRX4iEluY+OjpxHE/xs5zZKn2/sVf0BzxuQojYkL0HtniJVnFunTxpPk5jeEq
sVk2jt+QHxf5YNUgblrEOd8VKw0iVnp899ByD9+t+dMWhAmgOvBQqsWFrWIlQbsp
P6Stw/4P7x1mJP80X/aPnS336XShT7AdoCzirVCbTMAfbW0vqjsZ5GkxXUOQi394
olOQZua4SHeVcjVU+dSajo7ARuC+j2uFDF+YB/vobzQHRHN+YWzyKw8ofr354pdb
+eUos/tLU8QihJ1P16st292PO2EXa6XLmwmSzJqeFUYXzy8r6iHy2fYZ9OOa9oaW
+cPLGoKVueG/V5mmtiaBUDnJwnfdqc/AiluosmNdAg/kGa6VyvFtfN/wE7HzCY4U
H/6dbb6gW7tzFAJzjOJo7CLuv/oEXRuyzCVsP5V+9hb/UVTjazRdRA4Lo+f5Sh1j
TZCpeBX3mF24W3C3cm8hEbMVXQys4jAWZ/JZFIfTQ0H3N3cz2l+QwBvWOuFlgSej
KoQ43bkujAyeXtcQ9ggJantOgxgbCG4UoGDiHg3cG2fvxXd7SU7qBvV3Jq4Z1VM2
/wHK2o8UWqHjr1dzhJgEjCFv9PnokI2GqehvN2Kxo7WKG0lwYBuKOHtt9kf6yYrR
KnolI2POeROdEf8jsqUsocC/4ImwFYaSDNYbnLlgoZ6+bvhVpFNwDvo2HVn8/vHU
1VJajmsHOIV3ZLNqs0rp8Z8XM7ZwehfbzkMXgIUFByCKejlNC1aw5fUW6VoV4YAH
ifzDJEgU8M8fNTjjGsfh6XDLRPOGT4qo2wRm/Bkay1kSW435ozLzbUSYDII8USSs
ETLH2RELybuhaZKWxtY8G2teeMA4h2ctIIvN+l/YlfYXBe+p2uHzKM50ex3nF9SI
osHHQjmtDvoxjvQzvjFdgFR9Me/4LcpwIuKuD3zeTRw6xUvjD4mOsGakuXRbDg8L
DLtiaTjpXUrC7JF9HSRWW3rHkSA41/QVBSGgzcB12ugzm5nWOjCOY/CShQlZkLM3
KsMsgszdUgyWFajDz/zhvtjdi/6woHRr7vV97cIt0sZexm9hleB5/lr6g2fhw5Er
awrL4/Wcpc65ulaTZjt82KVmo6w+XYBFZq6Oox8r4mrVYV4umO6XWsYngu8Xwp3D
H+1A+bmgJ4jNRgeyhb95XvIxNRobDwdtzAVag8JR7cJZESTMs+YkOW4/D2xS/cyO
fx8EDZOUvptbEzTySBe15gGv8vpUIxVblaVc9xmO4PK9UjafJiA6AgyneE7GxKuP
rIUm3iqWDLTt6r3cs3FQ+iOEn+kl66O7BCqcTPVkLXftYNvKVIfzAJD4+6cz18UP
HzkSG2mqqye4QCMuHgvjNl1IdGvmW3svwV2As4oCWLbh8AylSDkUXbCM4sJyOW8/
AkO/TC85Z7/rlHu/rc8EvZK/WAl5G2GatAE6hOryUk4cj1zPEhJxFBItHBZaSHjS
hGSt877f8dZwIUVQWjIC7Zqn+/f8jb1WMkUr/+v0ExJnOOQglckZf1l9kWtXzI65
HIYEO6PCVsXzYbPxHUe+3h6BMLeUU8MHoLjHDmnseN3qe2Fp1Lhge5t3CRukTxT1
QAK9WH2fqTpOgwL747jPgUnDamDszDngVD9CNj1X2m2FNzSuHylwdJ7k0Vfzj8nN
3xiFVHy/sKN+vdFyzzRz1xuQffcOKmHR8xy2yyF4zKVujKVDzr9My4a4DFgWGrnz
j5rOoLPgcH3FzYej4ypHKKiKEVvf+NcETA+90eF4V8w/xXGwC+I9K/G/dfr5FJoO
rcVHUWgxIeQKmW7QFpkIZgr53A/zP9R24oC1WnyqrrNjF7PM0DBtYTxadgfEAytY
j3vE7IZ9Q9PwUx/3/DejB35OlhwElhIBuASfKB0RWWsWEh3+ObLhSc5rXdJBTue8
Yl9w+d5m07wEvoHEpv4k7bR+YFcefr6I0YH90QhUY3nWr9ZGfN12dM484tqHQD/W
sp30hpbTBfmnxyPZBT0CvEQX4yrN4Fpp3e9wxGaNb6UqIr1dJ9PMPm/HfbDRynNe
/0yaDdOm8JUklFn3KzNYQ1Pzgt5hbZnZucZBTKPlH7W1EqCDYn5UfSpgLYOwsVyR
51BZSQHi+YbDMAFE2sRLxaCsmLBvfWxWDG6ySVxbQ0Z1w+78RrVP2vojn82ZaAV1
JYM8ceJXcwEUSaCBoi3b0hUyn8vW6BHqFbevZFkNvZjFQLvlvI/i3J/BcZkhcSAA
RAW1rM4tNzYC9Kb1sEZzWjqEjHCIUbqU/zqV5oJJQYMl5T2kiuBQLiQxq7k2zdAe
BBh+SkYYoBkR04BMU82KGBtdNuCcjZAyytYb3HzBCeZePVxQrqE9CDLG9L3/P9io
umWpAJD6yciAVlaRLlx3IJ796phxZl8qS1n09ZeEQsa9JJgjRXzoCos6W7l3/cqx
w/oYlQ0X4ixBMI1re/8adRzzyefdmQBuPH4hpLheX6Bk7zWWMdR/4vYpmX1pojYz
DfeTydrbkWIUURYLYt3A6D+heYqPC548ZGgxMRtdRlO2QxMRcN6fiZwADb9r7haj
yOe0Lm7I2o9iACJei/5PP2jy/U7Dn/2u4XlFJch8KlHBrCVWZaWBLhn2KtbLJOVH
5T1dr8FJrBw4gfAskrKzNWHuwF5+EVRGL76yR3yXNmlBg9+4kza+aEhoL7ZsGX8o
woMS1sP0+aur825Lut2dxJz4NwBcwqhIsVYXe5LaXsYMceof5IZJZokjtaEfxFtW
XriSD13fyIy0TKY+iBbCk6rDdTB1u4a04asfU75sdqr38a8ZWVuErPjIAtd+UE55
mrKJrssCDgGg8kJKrjCWGtvWB9xNFVIOaG1uyQgG3EBVexd3HPDM1Wj9sHbZPXjo
qNmAsF/dKe0NlNAlDMW4uJE+1uJLe5YOAbJeTT0vNZ4PJVZEe/Z2k1T92WEYrfjg
Jkut2BuITGBbDOuWFQ0CnN6u21TX7JR44G7aXbIArRZThL6/TXmaAX27B+ErOGGk
CVHRlI66YqA+s6nzqK9UN42W7weBXiZOEjpESysSKF5kY5zCKXr0vfjH5EZxjZ+g
2ElfvqObCOwqfZw/1lVETBshDecgPN/wZJ67vHVjM0T9Krv++vAUYSyun7wzoBwp
8xb6Gu+jW3WJ1yZIE6m23nXn92cTUxgdaNZNkKKc5O9tKSik7KRhMA9BgaklynTa
Lsh5cA+MHKFgsOXlNyb2XR1x7LdkHslhlNA9hyVMHYNcagZ5Lu6eXnkgZ3gLF1p9
YO6tVMgUl+Gzby7qZBwMywIJ1gUIB14TiG6m2CKO9OCh77HnFyY1YzkkuqAIz/mf
xEG4L50PIdmURm5RtJ7m87YuGsKS5QVQTYO2DPrTuQPxzNrKZsX7NY579XLvKCUu
aftM2yJ7h+tXzV5LEQZvZTHLvXqbcvvnO6KPtcgvhjtNyAJz/ahAW/6FNkvkDxfs
zH1vd0fJb2IPSZsjW0HgYZJx0AyPu9+4M1B/kQsJ3DZvrSIs8Vy1cAD9Bpy9uaw7
QIdGzmmPxvJ9Dq09tny2ycDFeQK1yCuRL03hFGFYYnL12FfupHIfEWAcXI+23DME
EKvMKFoIj+VtxauVTTzllLU35NOl/sh9vXtqVqqBXg3JwvBMfZEpQ00fBBfH5+no
mxjxuqiHm9LlUtvO7tXSZlPf1K4mRdLC0spX/vmZefn/2vBsmFQ5GlKu5359u5P4
CrqFMde2iAeW11s4V9ARqfi8esLwncEnMmhTKH6sW4q8Ps835Zw9l+XQvxIZdK02
RXjjNxphFw6AkhLOyRPVyKbRW4/3FA1iNsYrFVkH3J+KhcVu7OxAbiIw+9/E4sl5
XpnzjTSnnJkDuvyRGmtDsqEBNsxJDaYVQH3z/IVkn7rs8Bh5kuwdy7J0N18wlGjQ
p+QgYxsjboI7ecU6dZ+/Zoz47rNYS+LUsgRnxffaOkvbayfheh4vqhccQdSYeuma
yZj7BSjcXbpMjvJbL0NUZBVlcmwR7S7GLu1VOs7Jae9BMaPUl88TcsyugSgRkhbV
Q1r0uOLcfdZWZNUoybNO1eI8lmdL0fkbRyxl/dqM00Jbn644v30HF/lfAxvjpyP5
ykktdKr7nWDjShhbK1qMCXp2T4BCJOZfykm5NcBVoIiZn+WkNp6UVXarWyaax38N
uxh79jptL/8RmhTfr2euRnL/l5BxEKABU4U+oNiX3CGba4w44YSkqYrwWUMY7gpn
NhQPv0PvqjtNvS3KgVxCyGXlDmmm8nN5Rhitif+Hn3F/2HJpnt8xLKDy1G+PzKm+
p5gvUsFvTBeTfQ3J0hd8WX+MFK4EtFtOBAlJ060FRt0ZXcsb+ncnAgNuwg0eryv+
Q9CSB46gSM0UyTm8abcWbQTWNNejsYO7iTZiuwGNWojHodf/yELVr847us9kfkR+
WJj/r+NunEP/OeyfGwt9KRBaXhYXSVBGVAAjXpyIi9S9iwhru1E3o+h/uMdU/Kcz
FjLZ/JAfuReLj/noztv3WEsu57luZPrFip7S1pMdy+cMSkiiO13f4uGA0UKArErj
XfM8zaxJD7TU1dPGCmpJXTzjeAJ7ejtbW+ODheQ04/1e+zs6vFyPFUdqqNv6jGle
gDQ7cjchq3cP+CSAx6PhoXJcWbmC/AYBtpATusxYgVvdxZeN523GCt4n2KDMUwPD
eWMs8jg1d5XmmlnJzX/V8x0IFexRmKgv/6kYWD/qZJHTyWG3dK9P3ChepgfhPcNx
C6x7ntpoQiGSSB4hvhNUmddKh6U6nkE67vc0DVX1mdFICv8Z10oR0pM2FTtkR9Ao
7K/0qitTTpAHa5vOOpRUa2de4k70CSnvEjeCqLjfxHDLxyauvqj6XWq3uLnDXZ9/
Q1fBSkjMuCCv6iPqRrcIFNkx/ymAXjzPpQG6U6t8fAWi9ljinuLMSnDKiPivm6xA
EJyMVliXPmXYEFP9zkrVLea7bX+gSPipMr40L9nmt0eCzni0zvy7FGCjQ7sGv7Kw
XCN/5p7dATD4BFluATYI7796SKlMq+R8zGAv0ORfYttNG+lgqi31LnA5AiDFpxkm
krJJ59zn/Iag9JRLiY4Qo4+1N2S5GKbnT3firB+tlFBQsiekWuAozxMm6tmKtHRg
T827DUdE/rE7UqLjYPG2sWb8rJ8rGmR5KyXju+w5KFQ4UwW6QQTgglDy1Xlpx+Og
qoo43KdcnKRuY081FDW/lVN1GWRVG4oZF7zVYP/tJelIxLOf0BO9cbhUQsVeIRj4
CaSZsstN8P2zxxSpHmMPsYfzcRkTxLWx98qsTWzZpWFbRxgABfYrcyB2a6pOh1in
8RF34ZDEAHRReEV/4BlFM3FtWCAXi7M7s7eDdxNvBDhcAhMWGN36foK4PQiio0xh
iUl9m23qPrYiE1O971pQc7FJtnV1UjF56oLAJmYDMIS0ZaFXgBpeDU9Lh24sKvD9
xMn25M61BPBFW3pkJnBIYZ2nfMNwoNH7fhXI+ho01EZEJpFU4lt+y85qd1x2kP92
wqUgfh2qWSyHEru+x9rSV/WRd1hKw6ARH6kptFpwwdKfKI28MZDOukptcg/k6jjk
81GJ8Lg4YUVTdItw0U65T46TVWFae6A2RbFO8wRXXxZB7W4vN3pQy//rID9WGVDg
Tv65xXLfj8xSugSY3GvzMtWN2MqFNFqGC8Vc8MCKB/D5CS85zOwjtGti0FP7QXz6
96+PzYwpRMHTbQUV+mPrCxsTHtYfG+vxmTgHGTlTbO22QqkBOkx/rvf+tw6rMGL1
9zphyRIeuhKykJOkSY43I5S7L04yaFLyBq7w8IINaYXJZRKP3h+XJdDNpWNDs0o6
/hu6w37yVlEPcSAc0bGnrDYmrQeAF4iJoep/btWyTXOSsOPOzHlMs8uaf6IydHDx
3sBpoA5LbkFEuwFJ2Vdfj4rxzPWeUymVrQUEjtruWz7fhGUFnI7tyJ1713TzIWmm
DYbkJT+6xyPI2cFS6rIByNQufxUKWHB/4ZkY9+DaOr/y4vPYT3wjuvrQ4FRxZSYV
pqttlNZCgNhj+ZblQjKvi130LKOW0nRp6RK4gMdNlZStpB73iHZEFt5EwFhJNxRR
SNHM1+Fnt9ZJz1BFZJSZv4NzMTQU5jHWzcRgXXtdfaYnPGjhAPgLNZSmk+qHk5k9
kEJHda+8YSG4QNXIgiCuJp40FJZhQYLrsJ7/+Je7++2ZnpFoEwR7XfJo26dhEoj6
vqHKw0JEMx/WNHsaq/yF1Xx/J10jcH6uC7jaVxx8tKbMht8b1jqJmHh1wgBSDMCP
eKz52zxkc9GVhzuS/tgYthgZ1QcLpi32tPSAJBGM+atSFd+8tebnj1WIaudrLmLm
f+sOrbDwb4TXhieS8MURHysBvRORfJUVI3QxGa4ry+TqMYJx+HWH9OIS+tOASsu3
AkeuGglcwDkenEv+6HPXEPbOjgeMJ1iz+L+OzMHFwxMZyVY2fsagnkpSma6IH41j
usH3C2K6On049yrlXRj2fnhrCsc2Ns2qGWasQJTiXm0n1BsMkppLnWRvBkCoE6CW
7MLaD2yjQTV7ZVjqjVCQ8yIw3K7Xj5LeN1zNtrYRuf+hWNTjQwCRNG4jmSOwVGSk
6i5H3hirFA0ZITUI9uwnHyU4VirHmhLCFGcvDDsQkWOare+op1JldpkpfPC+cVIh
p6SncD26nc1MctOLC73Eczp3zWocL0cubEHOfbNX3PVLiPSZCtWTVVCVya3Ia/C4
kF/jU0AkT9TByyRh0hP7ItS4A7Ite32Ch1uW7tt2b/z9we5ziOqkezD42iiZmOzM
K5AxlTTR2Tou3Vkxy49HqEtySiNtlhY69ML3rvCiOpn8HOuPQkhFVyCpPel4JA15
9yavl7A7Ls7STMIhVqVN6b5RsaZIeb04mRXpBdvwvR8dWBONAZUvYMGat+q9ZTKN
9aoqUnUr8JZ6R6W67avNSLTA5S2ZsHmA23cyaXXdLGbtVgKmdFw7opjxCK5nEmb/
rQ8VlNY+Ddpf0wn/UUrL1oTyH/KL5j66ZawdEfVmK2d9LxxIi94pIzrY4RxNAZ0Z
fOST9uiaZdEyxzieHY3daY05hMwj+aYJiFJ2Zotq5lTidGS1zjJ8hpuyxGDNjJtU
snCOooXy7mgVz1uc0PAFlGRf2NL7QHCsTKUn9VQF6NlU1dSIeoZ5oKlzXoTZgvSl
1po/ZL7MqGfGC4zGpLhvzGp82QGrGZC6Xuo8AKDfbmzOhocTJCiE+KOPWYqxZECj
asUKQMAesghycnXzLkMumw3t03pVyd05mex07OsxQLFyNyY7aaWyg8Kc/kmhcBFF
A3imRxRLZLXKCTpieq2SFOgRN7sQ7LiuIUbhBggnfvVhH0wFIV6oHb7S4LIsTq3Y
suOCyGG8AhhY4Fy0250mDv5JSd4di25F81vyoV98e8+3+/huSD1UtkxZS7kRTkvq
hPta4ekr4dCTBglrY3MhFnwS1lh4tyZSPFg6ovL/2DjE9PV2959fYhsxD0duBwpO
C6ADus7HCaTQSIjdIQ79i4GjIA+uxgxLDpZSNTJH13UaQqmRF3ElXh5bGH2i+OhB
CFAjSZAA6ycbgrgBaO5ZU93wPkAZQ/JsE5kZ7b+CoHrhXeo4mKTUdvUnBELiYL0H
bwCAxB82JRMvcRYFTq3tT+Ox3GgxdpSvZq7fP239XDf4DMwKm/IR+L59i5Q1hHSs
AhOU7c/uCO6rm/u26zNqekbKVkFHtcckoptJUfyEkiDpHUm/SdKfrojX8mvHP/Xq
CJyssF5owNlJ3XqNOyp5VvyuC1MWT5AW4CzHz4ZLyn80Pgae5PTMWD7EeYAe1MCT
6Ts1WugPQYvJFj2DsGv2VNPSsofQWZsMFpMmxPdWZm/xq1OwyS9/nI3Jqp9rnquA
pZqSWhBm4KOkTcTtLr7jGNeIGmOPDNNEkEjwvNoJ0ZztzfEGpUhrV3tj/8ZM23aV
kFlSS28rLORKv6Y1/0Fgj064bu5Is3Q0kUsKGPMzLl8+Zh+AJ/0Z1iljnnoxnoxW
+eu6cxGZlwTU/y/hZHmoYpiC/ozwjC8tg7fghCsNZ2jwfD5I0K0Iwa5qs7w2aoSg
nJCQYhMaIwygCISPRDwFoZHNFxV9OTIj46bnyuUcypjKw4QEii1zVRiLFoqZU4PG
Lu33cPoCJ8zTi0/FDhlS1YKky/couMeWDezXbMW1NVInhZ7FqnSqECmUFWvzeNqt
wvWTqGSAr8wnEUdmueGr9if5PVnwg9zUsQbxGVzfkD9O5XAVL943+3pC7xEJTe+c
S/Ipp8J/Hg7Kc2rE0NcbO9RExE5nH1IK8auTsJeF1Dzap9+iuNx1cvuOYA2/kTvf
byWcWyK9v2PIigXrpPeDSmKEF8epM2PkovfVPSrXPYqD9YtvWjBuWNQfumpjanmg
oQVywaOcki61W8h/BJRmmSe3ookFR4MKPejxrT6M2F+FpsqHKpMTITHf9vClcU0l
j8iH6dVbe+ZmBqMMpG2wsYrmHrkdzDg8rTnfMTN42TPyRihQm28ehuseZLLXsK5y
uNdjRD0i7qVXv34/rXAnB//Es3Z0gsfEDL3c0J3GKQeywboVniZtA6xIR24tFEco
P2Z3/P0cirssPvFHi2VN4a2OuEWcibEPUCt2HfMCvdvt5+xPq7+OLdqMr00z01KL
eLRsmPdhsry4xbn2ER8aKuoVgiBA4oK0eiQ9x2ltd9mYmbL1RUtsUGqUhpcVICAO
TB1H+hYGE5H2brutCN63C4ENTJAdtaK4YbbvrHOOV7/4oOQ7tigrALJIZqjOcwZg
BYob3kCk4P5KtNjMeJ/Et8zQSS7tTkcPoFVwG6zk/o49itWY1zQtOzp318oRFnGK
xwVjmSJmKS3sr8tvuDQm27cNeSQH0Ca9Yb/RjXcDhxUonTCir/9SY48iS0Ky9mzm
z2lUxzOrDJLA28L+vK0c14BfytT9CKVIPTxGVrhIb7OEOe4/e6pMqc3LFnucm3rq
nGL0SjU38ZmKfiiQTvudvCLrr5XVaZlGY2s3YCa9DJWaQbejZKc8IGjpETE0nJPk
8cVj6X8I8RImCp/D6eezWVysml20Rh3DeZ209WkNM37j2uNmbSKiedT4C+yJu2eH
u0jm+jNA3+scCti52G5PdqRDZuTgtz4z8aGKFbipbaPVk15L3+TFGveHOsBEVuOf
ZMoqxshMFlKGY013ZlfYFu5jfW4d+heepGH2wFR0kRRJuWYoIZ+BFZwKJip4mpB5
+1QNkCL38kpcgmipRXpDHKS7dtQVYQYyoUGzdYRU0G5vNuyZjqaJe1Eo9AnbI/9G
YpQEiIrgAFqNxY0phcnlBJBES80fHBxL+3kovBMLDYRX5+RuI8IjCMlBuu6D2Yej
u2+yTeR8b1Ei5loAICui8/C1DwnZXYJFmKFh5Zfzkphcbhn0SxJS9sK8lhsob1OF
tJ/xF0kIr56nbd0mLLXhc5GTZqDtqvq0eSx0+cYQWeXAZj29lJppBwMwUIGmUaE3
ytc0P37hkHhfCEBYOM5Qv5iX9aqbGC9Oans4/aNK0h4ILCgeNBCeGIPSsvqL5W9K
nzWSw5bnt6zi1R7LFBOT7m1NyXPYeKe3Rb/VO7O8dOIfwcoU1AQ0yZ9/q7e88QTT
efkkQBD//t/qRYfS4VpqIiXMmHIZL5OP1rnFoNfqBOeSIP6mpuuI5Cpw7UP9TD5k
B6tsRJjur0sHJMZQfUld8zX/0+MGlP7vx+7Rg10753EnYvFMbo7vXta6mZZ+WWQ8
1LSRN48leQuYeohMP0XQbZ/s7GjAHsbXQJWS1oTMSP3tF7Q8w2YtnE2nU0t/d7Lt
la1ryDhKLxznRusY/Cz8KP4p/bc4JOyxjuVc4UrJ8uNVotuPeQOEtYub24HhSLAa
cqilQnwEDID/8PeQr6fzB9i2Pved1Pdw/lMxeg/VFPTy8KakxBxdDr3zu0tRwsw5
f53Y9s+L/N3wR7cXKODEPUHaEtTm0tjOHJ6RftX+0MG/Lm/DYtqlE/EWd+scDRD6
hsKpE34Od3AD1XsFV1NPEibdHEjVK8woeVadbEIoSX6VEnvN2sxhr385z1K2jI6m
zyqJm2GV3rQI20Q/OB2s5C/t1mZ2ZI6u/BYs56Yp8lxCAtjJf2h5CrJX8ehJ/bs4
tDq1Em4GqbUfG6qkCrhetSrQal2pUjwNetG6sRrZNAybcW0Yuo/PJnEX8ZNSriIM
pZu05TMNgzRJSuneIAAJajOHNxI0tPYgaDJrpWCMdhQu/U9OM9mONutVIPLVuDuC
XwaX/K+bDbbIiozMlMKr28yEz4mD11sqV/vpSCwfd6gzCiV2ZzuAsAzcy3EfNHzk
U8hLGC9nD3r0Cdk5h0VV0gwIzOqYqY7aI3QtpPc53IZqtfAPm1WE/994BYdP7qYv
e+Q7RcEgNrboH/5S41BaSib50HaOgQjxLT92NVNh2g4jpwp8VaQKzJhQYxL+qrl6
2uG7VPDYmN0mA8FiyDgZxURH4ExmY1oa3YOdnp/jBRkXmF541l2PkOKILsh4TGsE
XZDh/us+/2IQC3Gw+KZsgsZiTBja0PuGxRzkWxbu0cM3uF/JWgvQBeLEm1hSpC6m
RTUUNrIliWLGj8LMhriU+S6s3QACTtKcgZEfp4l8gxjQcb2IdgyUZTY/8d/xZUA/
ztGwJOAjDkIjgGsSaR5I6KOZz63U6CRRMAJV/AnLUqiqKwmclrcipwfOihT+wisC
NvHEv186yVnvx0MPHLYJ5PNiRV8n60EB+mJgaljECCBptMF8Y8eeh9J7K04UTRWM
kZBYVCKynUhiRpmVl4k+t2znRtuF4dQJZ9Q6bZM+FSjtbVhBBWIHFktpuNjRCcyB
He00x2uK7+XqFF2vh5MBjF9ndH3Gm+aVYZqf44WyLDWVbDIYpqLYRSu4qXXvSo3V
Vk5pNgqT/ox8r5WXlLI1nEdUzfZnFJcE/ItmAbqkp6fRl2B/6og3UFwYWgxh+Co9
KMQTrhTixSh12JLFKgni8W2dU380eUS2CxInFa8ygIwHziWwSoWBtcU01F7ooqNV
fGriwc/HcGTEv4HFm+pjQ5fL1niPNl0HM4NAapHu+PPsHh2f1sh3SI210XqpKJOp
XIq6Yo0MNKmfaJmxjR5ffoa/pgtxXsQERkFzHfqrtMyvHZJL9Q2c1Wsyxtcx2qk2
9at1IGYq6kmk8IJF/YYJmh+9Vp4OZ9FDCM/BZlM8Zi8BebijOmx8yxna+BwexKAp
SSt68p7xNYnD1KLdd2V7NF6Fwi6TJYPbbBgiGMcH5nfErLWeheq1gEx1HlIVIA1D
DQJ37GyImAd6qmmuyz+jzcPLT8qT/LYQLrNq+KFBw6ZKo5QhA3rPUBa+AICQq0tx
PO7SeIpI+ZBdBRTgkFmli99WCAu2dJaaKlnAkyUXLEnSGWg5e/TMftKjRFy0H4SP
DeFb1jHwB0yjmG7If/LX7dv3rkMxMLljroNW51JzO9PSGnELLTruS+TyY+pG1Hx7
nC4PE3RTyvjBDbuZK1hl+AU/rbTjcTZPMHdmisbbFRWFlGpYDa+MClB28J8g+dwg
lqvLqMtFe/JyXPB2h1bcQo5T6a0qbmuqUYgFM+Dc8h+QnZs13bHdUW/sqV/84Ee7
nzcvlX5Mz6TUC5zMyVtpzMlSeUHHj3tTOt7hQscIhJlLlm6LMQWUKD3pyCnTpe80
0Le0uSLcjBCVHvpu4z18e5wPk9m+96wrMxC87bdcDyN2TvCITqEZTsN2XaS7e60h
LDga0zqqdzuVYpAwVI6NGF63wcwiniaXMSQnrvVLcaEONLA3AFwxL6rKQjvdjprJ
KdiiXAVBSJI1EZ04To3IyTcfn2H1CmXEN+cXHOZzNkqe1hFMPeuxQjhRIfYSgrOe
q70oGW89MKTLArKs5uh1tO0rW5JvXlySKYLrUMTY56bLT726Bx5tj9q/gwtr6Q9m
QZovg1POwFMa9B6h0BxW2CafkJGRHUamCRmgODeM0o8Q1FeBWjgoZdEU2LP0L8Nu
CzH8p28+XfKEuVmIKywtQio6d0KK2p7kq7hso16r6u9wGzYiBW97UQPgpVZLafWX
NyzKTnG5jdLkHXELK7g9tJuEayhxbR8d6aYwExP0xa/VO4+YAp4Lj63GuXFfC4g0
zQgTQza6znt4HoC6vbje9osZYDJfMdOquBNyHLJ3gUI+KZpufUeo40z8zGnbBALx
Lz4i0y/yL6O5Dv/i/tX94tkjN0QCjzAnDjydPoJzgG6AUh0aw1jzLma97EHCGqhL
Tl7VWCvalukbsj/EVdGXqzZK1qdu40yzTYNsdAKS9jY8p/t6nk+ioaRNtl+RW+m2
58AgQREUAFmLa+76d11zNtTE8jK7S1w/wle+AKkvR6S/DcXCFDFfJ1C9bGK63E/Z
/qR5cBxTU3Rd4qIJA6YWyBr9dXhZDJo5o4kuoniDbHO8gWQqqp82AOsj1wou/EL5
uH/s0Ms3SmCwFlMM6T577FAyPzIzbF+GDEEt8YX4QX1wR7zOBXmE7I79pAf+a8ha
+9ADhHBhWVNiv4Ejsi5Ws0pqYcXIe4VEqQRYS2s3IQARnM21qWOyxNwXltWiggFj
e7cYg7tNGFh1yglAcT2NNfs9qEIWD6swqEMggBgJ5CutYRyBgIi3VY39QvZp5Gf9
uPZ/IsNS24zYjxaID94j0S00GTMVt+4Q3hZEQaUser9OpUuTJSEQbImPTC+5/wRe
RwYXlcVjbl3y3PrUaBmbt/dTpI/YhTKYiKfb0dFX9VsSGQSHPS6nJRY5nwkR90bC
93bjFWE3QaDlq22hyttVrBxMDzv7eqoAjGPKJpUXdgwS09djqPqyA9RjY33n3Q8U
Xw1bNZvUbFRy6oKiWtpb9sqdSfD/JHK8ngunJiaLZ9TWwLnh1Cs3W56t78r1bjlE
M40Dqb/XFk1bW3hufhc+mKy+FFVgD+at8FOO+Hk/G8TMPPlpFa9VM8gkddMlfVjg
uv1DiIuXbG8ya9pYOSkYGv+CZdLozmi13v1fX372BDtCd9P1WbVzV7V0HB8oHp6i
l0Pn08y3Ge3lx/4I5XU+E+0KNHrD3gfrPiP+KJIDHqO4lTL3tkOJ0ZeU6+dfG3wE
+Hj+Ho3yTOiwW0mtMzZ0A/u9JwiRWiWs+f4FE3MyVJqyr/8qi0XwgpOVyMXmbFs4
EFiJPbVSFJd8/SQhy2/QbYLtzTy4RPmSZ8QwKldE0Oo0eOV5KnWvW4zAlThX9DsZ
RpHGjkVlYVEQSyZiBaP2uOxcSGWmzl0cWvocmiFxZU1YSiLqfIxeCONM9pwgka/v
cKPzqfk5aRIY+OQ7FzsR9I1P1ymnqvArbdHcuE5inaa9G4N622lDBdHTlwOS5mqH
oDH9k/JNqg7kPGHMZ+h4Gxd7ss11xbp2nHV5n1frTN0EVYBJw14pu7cXM6IQS1Aj
uCGvqeHbTq7VjB8DqfWF8tNSC/ghe9eqz9l7hbr5e8h1UFQ6n7/Z27kknlU/693m
FghX7IqsF73iaMduThCLQhJVbeVjW+5nGbxboMqONOLWumKxKDlcaqHY7jFjfTSQ
V+8PyIRN2a92SJ74oxFCfYJ+mQsIze4Pg8bvd2VnH4JXFv9dHmPkCqmmxmVotyUk
Fh0sFfX6/H3c2NVK57C8a0WTiSn/JvGSLYkC+ZWrQQL275FgwVrES/Zd6Xqn5ltA
fipV3iYW4niwlkA8gPupu1OhNgPKaBFGQdUqQeFVwplI8hg6jIBqx1RKrrLuGnd3
T3P2ipUvPNXeFUyq/62JGivE8AWuv+LbehipdQ45rtlNwCVYxz0+ry2Zv2E07QmL
kt3h4pe6Fur3MjXvTli2Ch7tU/BgTTcTEV7YuYCD94sDJ3Ibui45db9nJVYkCxDd
9cevr/sy/QvBXGASE/cJvehVqKL0F/ybzqsJKfjQ010tI9bJ8I6sWNusaPKrCpCp
ww6pcMBRhDG1ix1TbNL+NwAgr/+uF6sk3qQ6A4l4bLOYfihePVOzQ+adfh959YKa
O+t/DhI3uS3NrgzcMhQmg8ZbbXFodXSx2xO2V6cwFWB9J35wwfCYn8aBXGy3A87k
jFw2KZNYFJzXbbRIXInkJ+Uc9cE0YuB0TaSXCaQ6Yd4mXSMnc8T8+S9TXfwLCWaF
yV8o0fXucZ87p1xbNxhYaPYLRcnpfwVnb0akbggWM3giDCJbjHUErv57hb/qQJeB
YhSI1n1SC3vLWDXzmzzjqTiInQiV7Z0WpE+erQzwNTgCEsKbgoDNfguoN8mbBxnp
LpuoEnWgOxwGWRzGdUFVXDaGU5SkSEzi7U63nxWY6hLQWBfd9GZRnGLsmdPb2Xal
sakopA84WFrn/MFHH6vDGvYpjGxFujCQm2QcyEdekFenqkf2HDvBiGHwPMmjBDyu
LFeUVmhWyRWhKzCGGlYODSdRo9WEBafO+JsAkoHNo0zVnX6ohWzaGWeF8sRxDymK
eP7fW8ZW4kzXZFHphWXgBPtbWSSsF1am+ErBkNzOm2m1nq9HZYly+iY3u5+9VSo1
qo2esrMqoXon5zCrsNqm0vUioR9Fex2hHL4F9zBExvQ2lmqucRQWpHkEZNmSe5hv
g3Tqncu/TGUmAjpDu+vgsGcAx2TFNFiuB/BAa4TCEP6oNCGCJQT4DYosTUlNpYXH
Et21zxnXIVknRk87urBeTdbYKaky9W7lAoQKiHRcxcngGmtF0gu/ZE4xDzruT4Dq
MNB6tdgV6n/H3Z74OFt6rTXGhXMbZNJNFLFfWpf/omgETtKf/uMruRDMpEL7zxne
3SxMdDNanh35O/uDc1SFu0HrhraVtIOvrjMGAiAOMrEUvFR2/qCFp/tb+RwC+e/g
OO8K4Rd9gaupM85PdfVkNy6L0Z2sNNfCKxjnkXm34r22cga0/LJ6m14ttQilqD0Q
qv0UvuBA90kjetmwA0gC06tAQBPL29kPn0UyyNwl0+PMAJvxh4XqbaX+dUjUSCIL
tq55SyxZ+Jy/LQeyccYP3MlHyOwLq6l6Kp/Vvrgbdt8jE3k4YgKjR0uVduav7dWR
7ucqUPb09uwgY1FoW7iErQNPscdpf6+IybfkAz8iUY9FWBfnSEaHZESCrVAQscHR
znhtidKwHWzPP9T0HJQDlIIIpWpYZCybZ9mUiZf71cdW7H7UmZ3QfdVKYxpmlCna
sLpYGD+pMoQOKGxHsUvJf9CrXf9slarKOHBsaL4kok8er8kit4E+dwcarPUBOv1s
LhIymXgrHRy8fcpHi+3zP8tv93y6Hpp2MsneIu50kkidC1Icw3eLEgo0jUykzhv3
IfV65+HrxRRHzYMTTWRKXX10kjeX9kGVq3VZ13Qw6QatBVmzLuxsuHZNdU6y1T9F
ip0QzHfIH0Yspn/MXLg4T+dMyvAZ+OGaPuvRC2y39uzxTMV39BDnMOPZNaE0qVDN
UIXVa8iLo55kjYY15//zHnjPXFUwJ2QiPx3FSoRcXBv4z8GVeX09hqi7B66tWzLV
/A32DpOl8GnSmgHFiCbPDpvOx09EQTn+8Jtvv+GcgD4vsOhsJAxlsuux+r0E9ydV
FMm/S5LfaJ0pw0Yv1pLLwsuTJyhN0bnYQ5dB+wh2ZXoSHjTylJqWQwIzQBq+hSrV
duGD+Z8yITSo6HSWgUWPmckNuDuFHaf4y5zKfMORWu8oimP5Vvni23Lug7gzU6Yx
uuViTW4rHJpd7NDdyAPYN4thlx4xb58WSVLSsyG7fST2V59ID4O2B8sRwN055vdf
OgFlhrCvkUO9hUlmGF6XT6opa4EAvIc4Mo8ITy7a29YKn/NTXIr7p8oa7madzLL+
6oDfYO7Jp7qPUR+fUbmInIqb3fYKW2GzDlgL3ncLjJh40AH8SGEQeRMdZPHGn8N1
evWf2eHRcqFx1dRr7OAwsb3m47RxhWlwnAJdlHCmNvWcSMyL8MpSJ6kXGt3rTdfq
4PmzVALL/zcch3lkOlnK4HK6gJdZio73ywHHcKKBfgovEEDicC7bMP2EsCRfT7s1
2o1bxORNAs3lpYLivQIlsC2+pIprPQhOANX5/VxXyobJeL2ufxMWpnw8MKop1tX6
wyvjNSBTQULQY3CH5HfNL1uwE9H7ifpq2BI8zuiRbAqwOPw8COEJKIncWkUE7AWG
dvkGBl9wmhUAMrLVD5UE/2fXpz0/Yy0GX+40SLAA/xE6uzaeGLQz39tDS2sNaV+a
x0hWzj+dsQBRl+qKdqopbbMWNVrihxbiQ6qqpRF84e9pgHIQfuhT5Zbq+VBsXKAp
4f7KShpBNE8fYsMsWoN0DZ1ObT3ZH7PXCAbGxmrNXXK6ezq0j9Zj1Uq3nKx9pljH
2KsAZQ+iyJiXXqQlpVdN4d0pLTTRQ7YJUybJYU1sm27Vq7OXKPFI7Bl3aZCh2ixt
b9y6t+aHz8LW7qglTdjyXRTUfaTnah6wvfXlQRGto1H47Gowcu45p8uoCcNBtQA/
SEemdMGicE5Zot3rDlExPRN3SU2fR/QBxZ1446tZAPbQHrpNCUrOaf2l0Xdc7h4+
3BakkLh0iI6YBxs94rMBUO7vQ5QnQh6acjyJ7mchftisDL9dTE+rEXw3qs/+XSkh
/oZltcHrWPt6iTO3mA4M+aaglFEOouWJeP3M2olGa+vx9oC8S4OXAqzd+j2wDHiE
Gie/OTGu+nSRTrevhaUNWrkD8a5ATvNBMPONzcUzTvwMgyVSunA6ZdqywT2jC2/I
q+ZSZ8EY1N5b0DlrOxc7nMC+aamEbU/mB453sultEowFYekz8LREJNY6QSpVhf63
q41XEhyQAORXegTB+b5wGoDhrLXzjornArqTHsxDfWkgP1zDBJ0lkLIXQzZ7d1S1
FCIAyVYpVxQ14jRm6/6yMNWMMaxYp/kQLmsbZrAeEijW4TTBjXO8lX6QfsjUjAuT
oXKjxTR4Q/y/iRMTmAtH3/BHhqQb5uJ1EimbCmdsr/x/Q7whdtz8zBg4LDOsl95G
wJtMY6r4QG9nQGB3y2EtTRB1QTq5cMmk2WgDmjjV2d+BqZnpyeEWhtHuQAM8hYRt
peSy/mnvAs/7iI92/oUsRRD27BVyGV4r3Ec3j8myeOnQ59tDNv66UqrFkxBx3Ie3
Z28DaVF8LZ5Khvi4xEvbtbCEAZ3EpIhux4Zx2NdSFXm6otWDH36XQz9ISUP04QAa
VrNmifT2cvmTAwJGCwJ3ysq4fCyCAB6KsN1JgK0jrC7R6a9YQxss/RrXvrdNA2zf
OXl47DgcAO+b1v7VmHwCHUncBPoBxvH469gvTGOgNk2VWDtLtF0BpyvJ9CVD+I/4
qaplePGVT2S/t21iy+GcCyZ+ft0iYr1wKQi92uTqGukpEqvEf4F9RKdE7JeYaHJZ
MO58eLVXoMbxNGl3zzxnGsjCjFrLxpU8UU2CSRWHhgWmKKDq9NYZypV8hFmGw+Uz
x9VUai1JSvLXmT7ketQlXIdYM+eBOqCoJYQZV64C85THhwwG8uzLEdbrkfzZ8rrg
dPRd6NbLbOgVTCXvps3Cb5zi4EsV5edSGigxyntTgMAwFQarR4qK+Qq58N3kZkQL
A/TP+Avf9UjVeM1RdDmbKCUdMAVCLSPhLF00gQgmy1nhDFbqXH7/9BFW5ALHvUZ3
441DlaSe/9p2xM4wzQEWhcl286wOeCaUEVhwrwqskRohunDTNS/19KdKKsLVk6/I
sys9oK05EfLOk1LGYIKmP0NKLiNFLtAxLNeoeW1Op7NCKZLabWKb04lVAwEVcm4w
lIWRgJRiYW996QMbrEay41wgW42NZvCqwvU+p7hy5C/7FXgBvyoxxrk8dBHgQuj2
9VIs/97EKGctUrRqkgg8KZA6f+UQdFZenbFcfh6VgdoILplv/xDSjnzktZadY4Zn
l/GtzPTrrzmU8XxwNxdHNMuLQiUdFmxGjy4rBUoU7A7W0zWrwtgCb9IgxGiw/b48
zka3gkU4bTe/5+LZSiPN/2/v7JnSgGLXg38xLs3Y+zgCgeQSmg0EFRATZb/Wrfa6
ajy2LiSBbNdtnfFrXlOwCJbqln+LUtMLr/+vbCjIlNXJNCHNcfGdiM2Gu4/otGF2
AwOfkeQtr3hkuyrwTOvQj18umCuuDgyyQNJ+9LD8ASlCLrE+Jc4pQdk793l5q6Qy
586q0GEIlTRVSVbCgygI4zT7BdgxAHWqQk1yHyScP/XXtJSQZlRTpm2IZVuAGEh6
fSW8mshBEZmznJL9zZOSGXGFYeEbpbwBbWSvugAyf/NRGHnHpP6yRcgSY09HzXJj
ZpMgQREO4o3oeigDbGnuBTBiW4zA6DkhDBOKM43h2dhIJqALCgfKhULxQK3j33yM
/pBk4rp6UvW2KaaUNq6b8u7uczgKY7iK8Pc6v2HEUopx5hfmPqboenrEbi74EH4h
aQpYliptCoRgGPeZln7LGDO2BUz0T3bv8B9X6Vqk2BVJaGxtSwRYAIssvd3CJpwR
DEOM5yaWCQo2LHCGObNF0Xs4CckGhdnLembjyeMnmHdz5ZRjHDhQJ1NHFYTGjNTE
XUqe/kbxRutuSgCqPXVHwYCl8C/O5g7jsMz0e9t4UZhVUjP6Veh+eX5WxbmDHHK4
iAiUEWYF6kea1/z/SWsXkctsNUw3qYrIQGMlTSdXdU8qxlo/TE69gnhb0qzAWJpG
5qzTKObBtOltpvLcu7DBaq4aXi4fAlcbv+IHFvrygyL/35104ZolwLZ5iDeXwSz+
3hoUv657MVYlHKJRcmr/JhJKIZb4rKrIkbuuUb6RaApE819pbAWDPV1wW2AiZMR2
aYIQxqBzEk+L+N6P61ZZnsfNThk6BL8/h6TVk0y72rh060tMf/He+WhxzXtR3FE/
q1VyJwNU2JtBnrDIvI0iQbE00EVi3vGMTjWnJPagT3t6mBkjpTfmHEF2/vB2HK8Q
WLEzvllwJDgQPDBCWQq1G3dQh+Xbe9Nw17blulbPwYwKizlP/K2HFlsn/eX3MbiQ
XpjsVJF+vUUKh/Wjqbg/aqLIHqkWPGqT2B8zqqrGXpY2P8mral5duNPPAxYd1Dxk
pn/AxchEXHmr0btzsWNmJQQ3X2FYP0Gr1xXDih81k2zshMJfZvdxwXwmGIZcLlM0
ZHE7RSAOa00NuusTBT+eJxNPb+E6cBKpgFUOOIox/zZNjdHclASNCzOms+OqwNO1
rZYEuaDUFeezav08nvtDqM2hvJGEE6SV1pzBvO/2MxFzNykLaWr2uk2Zgjl38hl2
xzlbhha/INyVbf3KOk+kewJKXmO9FsIW+o/o+FH//qwe4mJan0L8Fm6zuAa92n5k
5o5TSK+Jr1LwpIe3zcK28whNen2Fa0wANGl06U+9T7irQFT12oP1kOdjgSRm+x+p
9m01yBg9axOA+loA6Py8aNwJ1Vt50dgWpFdYQ+xQWzJSNIkBdRb/IDI40U5U431d
hkXwDPQa8SjV+HHVurESA/3vrhm3j/eKrbZ20CB0wl3mtPzMrBzfsP1a7zej5M6L
hECpWrHPkzHpkIEl5rfWLIjNFC4ZckOPMoOex9sc78fbTCjSwlvLcw4/BVbpTL7S
XGJigRlZPF8ASqEjN3r5Wk8R/4JyZxtMIxoemM/iNQRVCvvOi0EpX9eRvQWCBALo
I9mv9m+Vrf4CHJLhTovCw2YcobAp7ZtzhAa/AXmHOJnMyz3/BYFvZn0RkojJ54Ak
mnOok68TvJTJc5pJULK1GnCxHZ1mmfmAShQnx4QiU27Bjzs/9uaJJInQZb3Ulqlh
m5Bvh7erCFe+LtBjmrzYw1SKXA74MxjMz2SdSFEmAd34NaGNh8FEFhLpN7dbcZDg
1CMU85M8/VyPsp4xSnXmvcb4ck0EqbXwBkeuYhyjEvJBrC7KBThuhcHdKdImBADI
jYuwb2FOy0oHqXwVmjeKvsWUn4vfNteD3pcM3+hpYwgI1fITw8jtUYzWg2L7BGcG
9wkaK/7az4h03846nEc9d9Jtihx92aJ//dauOHDBDFVYso9ApDBk4RfLSt3a9Fwi
ufup8v4eJ5tMJeCrFlPVBihAo+VK2IJ9yeFgN0Zb0R3HPAAM2R5/seFBA1OpBYuh
z4xO/XlQj56P8qrS73IM6dXcSqrid28fuG4d0RjiqaDww1QgnlSsVkpJc6KwYbrd
fnNOxpbxp6udPeyuqMBxXyggKa7TFQp9yDLwzkbpgX9/VMdkoi98dKDrmrW6CTxs
XCeUfmogYsmc2RkYlwb6Dp46YXMXDRAJxm9Wsric18oEKWAtkFV4l9bH4at/wGXT
UmmM6KMeFmTIi93S/7wP2noSpjlc3Xep6XbXtmd5fwJDQpBi4rmrxibgqufD05Jm
/mGdq+yXfbZe2idfKL+4Dr8fo8e9W/nSsfqbbesb8vv7a3RXk8FRfR8do0YIaqMx
76IEi59a4VDY3txFTWooA61RJ/MKo2OHkhS5zBF6z7eeQg3H6PKneKe7ODHcUdDJ
uy0F/gYIT/oR//ZruXigy9oDn+m2aFyDO7spdS3wIByszuKBlTEMu+BaJKPmC20h
OIHZ76XUFbs0kE8tg6WToOdxNXHJvyd3Vmu46E64Ci35gSZaR4PB8BjwTRYkdrBL
Dlm0zDWRRtaxcwbY0nmJB0B+YdMPz+e1nj7o5oUN2uvAbYzVdeFWxDF8rjsosIqz
U1yQZgeA/R1DAadv0qrWprUrRS1JM4/u80GRV3R0tn+s53j0DMZunoAwdouXHEZs
dnbYiPL9cVOdmvPV8NKxCkRo7kYjreh85u6weLpaR1vEqHTUuwcUTR63LnFP9HD4
BmFodwTypYAF4uVuDDH8BwVqVt8hOb1fUzuPvve0YYcoMfg5FalPaAUU0W98/Oyb
z4JO84+HSU/8OrBoOI8P3MWtV7anjisD1qWwQhYrlT2O6hFICiQXGB7LR5ZNT6ic
GvqVG2+7P9Cnd/sx0uBqzTfur34Nm6R91Rldw76DJRjBDOHm2XFUInWRMhdOrTMt
FB7/gZGapYDxj19xbwi2gCThGkApEItBmnfYOb+9uqTjqqWuGb4eliKcCsqT2aLj
QXWCx3RtdsJ6jCr3VVhnfrppG3jqNtLCFQFIiC9mo7EkCJ5uCbmzjX4FsPGfl2jw
t1DonEXZ76oBu/vl9vB9kXWsRm10xtYIhk5Z7ZLNucRlWE99igIFMlGdVy3Vdc52
yHTbWtjJWK5VhdMcwFNI2SPBVJ7ANwzAurKddb8jP6pCjhlDVkdU9zKk5U7iQYRn
pLkLoPfcEI01HBJRk4z+PNQcDZ36DexhlkCcFVQ+lkWW0f4aB/RAp6qfNddZ3RjL
5u/QN3sgi7IBcn14rwe6xnxGsF5kcOywA1PobaMNqzBUa+8zKL8j+6poEc/Kuv4y
xNXPk2DpXPDYJ2/t896duUkpG4nGW7QXI/IN29keud8Od0thLth6Mx3oSzNyVhVb
J7Mxlu8yPIzemg2ySqcsSXISbBiElDOm6xo+FWFGg9XjqNFJyijmTvkooNOVD4pO
Acpo6UrvGEl4jFydZQfKdPsFbEAQOg0r06PSU6cuuUN3LCwFk5oRnTlOi36k0vem
qI3W5GCCVhP6XUE4gWLAwuNGLhfuE6sxfjnJ7tVV3i82gBUZiRRkQ2GvpoUzXFoE
fpVLKmzwN9AjryeHNLR+vSvgVcKrlnsd3ZhrZEkRY2myndk60gIk3p8j0Ag5eo7v
zGg5dquN5eclthIfJwg3gbp5KswlV2W4RzcCm2C123+SM31whyi1CT+R4XMdL9q+
TkWUVx+ougJ0wGDptxpcUWG1FgQTOiBhNWK9mbAYgzgxjaICQePFJkmDYXo2aZ9E
iRMjAKw2zA0XWHCYPpQgLHaX+V3XGQVDLb7ZT4ukO1IL+Oqe0omMEwiHlXC0LbQY
dPCCUhFhEeGIXyQZgpmoXiVdA8g1il1N6EivFjgIXk/zcYRZJezjUBU7gFmW8vbI
tphTkBUc8CNN5GiGOgImyMIk3fbGseWsJNjctUk5kktnUM7R8t22b12Qzzz+sRy6
BXZeUuSnW6asey5zGSgt6B8QJH1pOElua2OAuqA+klaE5LvMKiwVC6MdujpfBKEq
eNb+0oyVWVNr+GeMoO1TdzUK+i35WdlNFEH5SiTMnNGCQdw7cpGExjLokWoLpcqf
lz66EyRAF6sxohohm5WwFfjjcm0+L0Hb1S9SYFmK1vxfuCcRrZ34eE2jZtqMk4bg
ju09n93WAsXgNEOusIuGvml7ZOFcUK5csIr6o9NAxVIHMKfCzgygC9OpwYs+/W4Q
W+radqYW4jSzuDxXG2Z22o3rhJiNXsxF8dd5gOKZ4E2HfCeHHrp/9MpIxMymo/Y7
WvLSit3vM9QwytumjVSZRNSeucorlFVOILSeXTsfG2IkA/qiTBtDg3z0XNDjjHD9
uX1sU22G1NI3RpOycb0T0p3s0+lXu/tO8Er49dYZlzgQlcGRwFW8ZtI2gB61eUDq
hkiMUBcPQ6H3vJzt2u2bXrusaepDLHToIy4NzH8UZlC3cHXt43fN/ANP/Nd1D7ba
LZ3bF6DPLACYvsrioK0qEyuqPGNJ/nXxMCSBdrq3XZTesBHALM/50nfKPo10RAEK
/Ct+db1hei6p2nwouc6XqXJUlNOZ+eifC8NmyfD+1gyj0nlUCgr1QlrfxnrzXvNI
+7WV6ene0OV5F43bWiEna4tam8rsWsbApFVLljISfKzOIC/Qw6wS+YGbHxn9FbjL
+QE7GGeA1odc+b84Vz0m9Z3uXyfmpSEq8XowbWguQq5Z3HtCMTQj4HlV/sgaqGV8
prczCDevHrJw2RgnW5t5VY4Y4sliCwwo5CL+1YkdQTRbb6FxOzCRlCsMsYordfL1
NWm0Esfzws8x4wuKkIJaHpsdmDbk+9XMP6CPII6nc2RTXwU/SFA18VmVBl3gODhU
uWHe3wtX0ryWnCmcynZpuvl1UlVvLEvbOCq/YcsheJm+wYR3qiamuMOh2UJ3yPms
EgVNZDzDVQDmR9X3BKyhZt7/uYFqvbnLDXDqpDjp+/2YJENxnUjYtDO86tBaPx78
Fc96Q5qxHSvZKmD8rudQtRsqnRTdvvd1E3HxvXV3f/b19lXnyeWeAKznn8+5FSbb
+kMb6HiGAme0uGnUBoSMsQ09Yl4AbuWNh7V18olRLX0c2anOz8RhDt+LIdW1UCUL
rd32eA74BjvLluGzjxz0vNjbWlb+lEucLNKrNLBTRHp59McW7etkyvTfZYl3QVa7
yg7D/VfBoLPHczb4sYouRG7yKDzG9z5nWCHr1X6RXF3jydSLj9mv8uQsGvz1qa4p
qAmTxDaXOpLOUKt29ND1NUmgaf1HVUmmcMw/dIoy0coXbUmJeR/GTFje5wNOW2Ia
Lwvg1KifSZvdKPRdOMpDHGTQnfibGsBoise2W07Sjgl5wt9uZyPCJBNJufarokoj
0XigQC/K49G79JchS/R3B6H+YmwoRNrSzRVWTZMyWAbd1I94kAICYZFnRhDHL2uJ
VKFP4wl0W1UyitecZ79K8vejuBkh46a5Wv/MFG0vZDcqqksOLLm2UTeUt03GbVpU
9pKc3K1EwIzFCkj2t6DXbvDrokEz/fPAK/I+0QkOU8WOD7aRhR0c9u5fr6g2oQQz
qtiWg+CsCwQC6MFCGX04UGkSFzgBewzpJ8KQFnEeRBHqNky6yqZJj3oNMKwXCNJa
MWJVNU426V0XY4v1/do1rZh8I8EmKK2WlJR+y8SXl8eWWHicH3y27THEFgnxFTLj
75WrOmKeHGyD4HDa95idFdZrbgcz3r8iiO243Hc1TYeHqLMXNy4vh1UBHup0EYr1
0cN52aiTfS9ib6f1jGCh6MJa2iZmpMULssdk+chGsL43azt3PLqTLswQDV4fmgdZ
nu38F0HlsLmF1dcER9v/2QTvWkP05oUpGtJTmEpyUXElmLgka5Xphu33vrn3E/kK
d5EkaZ5/4Uo5+2ESWruuA4mZjEvxfhB33X0EJEYctYFjkLVwhxbk03Upm8hICUtI
aFYzeRw872yaYIpGBafHqrZzT8z/ml0IzobCjkTnUNiuCn6iZtWVTis8n5l0MLSV
0qcLCq9Bqt6o6E1PaFnPrFzHt2CVpha9dMeD2b7RxFrXG/Wb8GY0BqifWa3004k/
APiVkzdWVNBUXalLtSGooWc5M/JfJ58+K24qWwnWA/6p7XXT76TUEzkoYTgFFYrz
0ZR0pynUbnlwA7W0Okukgopr+Qsqj3myZ4SF8OFnXFhB+1xSxqHcD3n7qWsoYRnn
LkxeXS/oeC/CKWroAycU6M2VS927NbOd3akVlVCIHKBjb23C9iEgggG7fB8adEI4
aysENNtckKAWmz3Bhkjjn9OzM46UsGJOoSFZeDcqkMeinbsrAB2XBM2QLcVbjvKA
EIYApDZZuRRN30SYWnftWjGluf4Of3GcXckurzU6mvc2XlUR7hay09msONeP/abG
9YyNp7I8eKJGXkQHc3Kzn5EUypc02TbPgKV3HK0a2i4XGWd8G2v9Lgwdzwo12x95
O4R+u1hCTorZnZXw/wXsla7ePKgVp8iYPW14UUIjp2CRa2Emdx7+IXoY9aWuTr9P
OvaL2yjlCKr9jolTy571t4Ao4HE+G6hj7jnth+vD53I7BD8N7nhCdMZgKtvldaZD
ONLwLTIfZyBdx2xQaxTioUmman2hgVAo5nRXxcukDIFa6dNmnlaLmGannut1aJbw
Xr8E6Hz+W6ARjKvMHIrNcE6aiTDQMPu/+ObkJ3beqjVn7gxLqZC7HuxQKp5PaO8O
8In0it+srdQkVZezWAisuRlHvzj+AaoM8/hx7egbOEeVL0NTGXONI6/nAVpYhliO
tVEpy3MU+FM5tSH1R5ndOOdfMhxNp4F3Sfj1i6VVxPN3OPolEfPMDhN9fwu8aCmZ
8DeviKz2iilL2IznouhFzrsPMS/jMZwwMvFFcmgp+DWkSsjZ6y8aOWfVRvIoIcoQ
jQU13CCe9Hx4pHKXecfMrPcu2Eq2RTO58KDPe5IodQdz3qMmytW6WSC+FwpgeeNT
ORE+OVXMxdGxVP2g3fO+9CDPGh7SyMOKjjUArJKnW6uVMUlPMT75ZOlqcGy+MK3A
34/nQFgLKkr/wqv7y7g+i5RFyL+m93ACUmw4tnJFtavdJxHPiDBYJM9bFJjpzI3I
uPSQrfzO48AQ7/pziQvCfPlsE/CmZ0TT7l+A9ZyaRxroefcz57GpX3bI3SYhQBGo
XCuyNTKcMQpQevk/8BPm4AxXDIb2vZtwAPwbLv8kdwOOQTyj+PBcG4U5Qrszqqul
kP5EFc59BWwiZeDW55RWNQxTs8HWAlaXpP8vWUy8Vz25DNL1Sosju3rCaI/iKvyO
V62HrnHZExVzwIB0nuDnVI+L28lMhQqqVuBuj9Y/DuKnyVm0ABY4kRGgryXUWnk+
aiTeyz8N4nUOVvDHjcxhT/vpID38QPkr66zm1r4OCNymn4IUp8fcirySN6bNs9YF
52a+WabD7K+niSWs0LxOgXvvQEHBxNgTFqk5P+FSxuul6hu5qAJPEvNNEOoh/56e
FNl6aJcW9DygRH3GyhV4mJZofE83WBFjlga9jHPDINV+Zth/Ea6GjLI3XrhFS/TX
WimeVsQ1kcIEn/mYOh18PMDGz4nTfRKPEHDyYk8g9CMJ1TqU7J9aCn1lQ4oTFBxi
s2ldtjigkJEeRxigQcjFgPx8Bn08aVM63LGHe+/N313D3rncgaUPkcDD3SEQbqlN
yBGFy3/8YOJ45M+6grLr9C6R4SOdvR+czS9jRczItEjnHBp5MMnApRQcAqYICSbR
yvzfRyMlo/S0gAuT8SxKxqtTxB+3DOELkfZ3gdiR9TlIrkNlujMXpkizmUTm8sw8
YOsYJSyTg0blIu32/7rNxmCsWteN2bbvEWTDLFQz/vO4jSPAByg4OMuZSRqW9gkE
Va5uHMIVEj0cS6f7HnywVpkOPLv2lKSZsXfA8eAs/n/N8CLZhLByoWTsaR4C2/WJ
bbLIDsdh6FuzKA7fUeg98IT4InabCo9uu0wQnOhcN0VUy60qMWxWIKdPtYkItRiO
hCT/t1jF6GWr8NO0v1Nyzmj+sbtaYdeROuymjd2LvyfnHsEYYYmAWKQzCtB0rMyH
Pj4NkTsnRu4IRuXK9HoFfnA7/pxe9leaX1ApV++d1kjvPkf9RdB+15J11PTdngeW
Tb8aC/+x3SAFFB4egVxZCHq7LhnYiP73ZOYxQVC/5Jd31vTofymPzSYkFF+B0mGG
7Vgju7gogV8y3F3MiLDVuoCFPYbtA3D55Ajaf3Hp0cr3PXbJMAvI/vqs+ZykmMKv
wmTtzUOgCADFp0LEu/mofJ796ETevMa8KBNYKl9PKBtlOmiQW6t7iswN6do6Jwtc
QspXa9OxgC3MnWfIOSBLO0ukKO3rqbUOkqkMsWK46gNggvrNRX/nTvI5oxzsAu6d
JUNDLT2xPb4SUxw/bs4zsBzD4aiHBffS1we8Lc0Wj5afxZ/z51aO8ubcPaVDiBCm
k885+arNMw/tCYVzOaoNZqUiI21xg+4m1UZPwQfanlDFj6wRzcPgDd8i4DScEHYj
dV75IwDBnrv6sPPMQttNg0M9bi4sW+JCJqMoZE0akIKIR/Llb10jN5rIjK9ymRBo
+4D4Al4N2rGmPftUm16srKqJ880aeK9HMfMx47OM/LIK4Ao4if9TCG0RkZEhv8KW
/vQFXuQg4JFHN4V49rhNRSvsnWgc+7gQbAljtzzY1ugFHD8AkB2bdf0P59ZEiwq5
ezHj5cvfpNX6Ix580+Xt7f8c2tBULWloc8L7NahyvUazNQiJkxLlhYyMAzUDjVgB
N+9PSf8lUpuZk12FE7u5KyEmhlJGYeWJQ7NKtaYxv+5F1p4UjfHrURyhMFkcOELI
9vTV4uzu8W4rWNzYxRNo/hmSESQ0IVuM+AdDgyHo3Ncld/9hzk5Gzmqox1mMd7H2
Kjzq7/afspTPLpxsYdhdp/4c5INdJ3+vxC1iK5WjzIwDqFm2cqFh79ZXyrhUXaKg
HaCe2btqdWQFiWNgT5MUB5zriIr3GOwsrMAhVTrnP8WzMKKun5eYUrD4FQsXFkFd
dRNqTZDAOKJzXqwEHcNNfbMURzKk5qQ+hE/qtVGfbqcqW0ARbfLHBqn7ALs3bXVy
a9xn5AQ/NAix0CfC02QLoWFND9ciFSplWZGN4Xt1RXZv4azVYH/7ZrohbN+0Rm5F
OpKY3LUDqgV/bpR5/RgfnNJuR0D0nAHb8PJ8YYnU/CIyl++2Kx/+7UYxkHpSmi6H
rM6XkeXfZ5K9fm09GHJ3x/LGLU53ih9k/A3ir+uoBTsU0BZcYp5g0bsdHdwYNttl
KySFY9DB6JCAJ4KQbROwrmacDxYXV/ZAKu0bE5A8XY4oAePa5E/0TTUtGuTsSd10
U3tgSdUY6HL9scqEj4G+dGe5WzvNyzzH+9MYd8pQEc7Yf7IwPBa4s3NGhe7+sz5Q
/vFyonPTmd9ympgd7PbeCtpabW7qsCwDRw8fPVBv70yd0clVq/zR3uylh9n4ZylF
HzrC9zcXNfk9z5rrkp6H0BGgQ6bToSpvEN7m0WaJaWlYq6vSVEZQ+tGqlXTRSQOv
lp4K6eRh5+IvAfsxeCixojNWSG7tZh77jBmo7CNeh9dNEAIrpj0VR6RVZP4t4dbD
vRRTRLRa+2xFHzvmay8S4RntYOB1OaOt9bDtZMiBnM8C7ECyRPZjFLuhkeYBSz/t
Tpv05N8sOwpZGq8fxCFVNNp6kI5KQg601pZdRONpyHd+L1kykx1BJcJ20DY8xBHN
TPxY9V9rg5EanHmn4bE8ZbIiMYBBM4WNU3RJGjiH2Nb7B63H9+szyVrAvlblJjf3
o5XNpQYmOJ1hIZ/o2DE9B6PkC4nZMxcWAK8oy5PGEJJdGQH7/aakmJbqclSNMiQ2
Z6jVNPB2ONlMVBilLnix4jVh8WknHgT1H8pJrGOI3VnhSdf1thh9e4S2xYyOlCM6
sexm5Jyyet+wjC4RI/wCaAK4k3dWApXuK3znbcN1+1YP3kg9vV+lOV/K+PPAV+m3
dYCg8TdIbPGt+ek0jMS1e2XKpP+h84E/hFgGJ9C6BWsSl8MqIMHbpupz7WvnAiAR
q64scmjwMVnIoTc6Lv4nfjlF+m4QdKg/QOaoQZC6F7R40SZUkB272BxYCy2p9XPA
uzN/TlvEsGqDhYWBprLWiZ8uxrv7WSGy1lyEt7eP3Q5pTHGF41Zy69Ehubpisa5u
Fqz/CosH+Qtymfa1+niGYaTxI73jmxdfAfinS6WQYHHYwtWd5JDzQdVkzUZ2wu5R
C9EadO9sS9cLd0/BEr/j8fXhndGZK/2Vf5QS8ew8B9khFHGBtUZ90/pVg5nExqvN
8AbtMykFNIbcnpFkZrVlgmP7s8Y8xEQBrPrTEMsjUnwz/0R1B//uFX1mnR2+h1Wm
TaBzF8JFJTLHAbP6DYlyiA+DwTJPp5sCyz5QUzSv0vCtG9cgxuSUhiBRr5gh7e8x
PSUVBJpvbZIkcVYJHbx69T4x9lyawdkLorFEImGW1U/K0nsVXMo8ubow+6lCxq2M
1XAmHz3Gr8yKVpqiSkrPkSWezAc8U5tc2FfvR3ZY4hwhF2/kxx1r52dv79XRdmA4
RztvrE6S0AYPI52aQ5rTRnX9k0gXNHe9qFGewg+Qd3/oSn5CqzFbWQYJQQpXH1fj
E4X4czPOuu3FSCzrhYQ1eWF3JAkkZfs3tgdNCffKkNZhMxQjLOZr/n/4tAj0zrts
JCsYB0emz8JaMjns4tfbvyyWfGJpV12mXEfSzDJr1WeraAn4Xwr9L2UqhP/lppMj
bFmOngmll95cz/ypxcaET/gFXG/0NZmvgs2qx2m7Nb8SxZyoEjlPs3ieJlitW2fF
vyuE2d1nVsPK6L+/jle++cResd7tVDgwuHa0vMY3UaZHd1ovqvKgU0c5/mdUNgTx
o0g+nkmxVWynvzTt/QISB1ZIGww6Ly+3SBxxpYXTLi2XM9zl8OGmu5m2lyxMX3R2
cyt02aX1u+0fRGZ+Vkb8XgRRhimN85x6LIsJ5grTuRBmAWOaobBDJFsI32fDFk5C
9giNhs+POolY2tWdUUVJILG+U+g3sGN38n7gmFxdxa87WWRItV76eU3QGS7su3J5
jYvDgoXYUhyCv24vlex+/UycyB0n4Omd+7Dime8fOY3sWoGyUDE1Xfy8x3ITG0/K
+pVY+GIivzU5jZDJsZ4HlgaPYWajFFh2UkyRYUqi3vu5ZEgeG7969HZHjwnlnHBV
3X4XQpDJA1+0lUcCcKLvthaVIk+1XmhqivHKT7jqueTycNHpObPtUBVcXFHAqjov
PVz0MGzX1uh1KrrXLJ5Yq8F/nO9dRweNugw9F9TXwRfs5avDPtd0Ooj5LEl0CVyc
3HtLiKtvhyXRNmm9+F0UT/c3Vm0UTwGK2EJrQKooydgAFFnzp/YTBWHZNrH0CASy
/BLfeldEkoLT+UA2wZI0Pb+osJL/wQwsEVZePLdy23g1+Fd/heV9IH1kpG040qwG
H+yauqN/6OFcooYT7t+vR+UeTV2VCT3Qy5LRONBiTGM1bDD7pviaSwpGD5C3i+cE
lcxfnqLIRm3/n4oXz+O1jqP+s4f+whMLKIPpYWPa6pLVrh3s4/5B5r9Texk2eYV9
broc+ZFz6D1r/oKJlsM0VoSjoD64nLiAAhCA4Kf7WK6O3UuU6aARtamU77Go74ef
MkpL8dxY0fX9QBVxVKcsyJR87jWKnxpuKp95kx5XXqCAkQ8F5DrovdVVYaIlE6YV
ZRBOS90jA9VH39wsS8SNfq4C6xoxjIx1xVXz1B8/Bgh6R1Jrc02GK/gyBHkEXwxE
SBRkCgl6ikIhiyIYWwF+1dQ1OyjJDtBnPvS/UycOze3xUwLKnkoS6q+RqbsR4dkA
OsW4eDV0nUBxBLrc6qTZI3vAjRcLiHl67jAHqnwSi4EhwQkC0UmWYgcmoHjRV9iV
xPwY96E6Ydh/CjpEM1bic1nfAvZvMJItqoSy2VvEuq79UPxZH2FmyTcl2jq77w7o
4VgcD+i1vhozJ9DBfBlnH1TLWur9tKgnwJJu47rhxzrBGOYrjeVJhptB6WdwGLXy
q3gyO0XdsTqLjCD9IH1c7fajB2x2nfeo7s5Ocs9WU4POYF6zBR+rLNq3h+WgvQL9
Vk2qEUKnDAQqHSmoLdLFnbugSwfYjeGUlIAacIKelP4JGjWINM9QZ+JjdWSUwp30
qdblXCxtbTRXrwPQ/NlS+KfweO/aVx7hdg8f7Onlgcwm+jSlVl+ZVSI7/QNBpXqh
8RNMYCBOLjr/dcqPxujJHVkJv00+XLoC3dgsXyWYQpXnlfZuDGDDyn9ndb4Zc0F3
vbm0u62GuD6Xy9g7X8EBn8dccpDbHkuk6AIPOg205eX/sX56mQQhJzSNBFd/yT20
ZXQ6OJBiaYOdp0YDHKC9ofiP0vfF3APzlP+NPwT6dmdQKkXiOOwboYrcOGoXVDyH
gTYBu00PVREH9U6GddeHOO4Rdh6TRsJjx3n9p2OO4iQiuRXYuPA+suVg2f+mjMfU
YCEljj3ptOv3NX7nIVYoxM5EP9jBVH/MIURWeMZYxUgJunE5eQOvxyjnm0ZbFn5h
B8s2lHib8BfQEBEy+Ui5Oh7zTvAViPyBzxR5VEOPt/ZzsklXaNphludLK+Ysh5kF
JYKsQPHopCX2l27zNP4QSzLR0J3Tn/F8nuBq9tqh3btizDNqadyIldbekAP42qUw
fZkkdiQkFnw9PjQVvxbGWf/NPFKEhwJ/ei+5gElQ6iQ6NIt/2G5dfBDPnWSY6XxK
CxgqtAPla315xOe1GQ2Oxc//CROlpFffPDA1hR9xvRD69wHqOqz9K294D2+LCaw6
4hYhbeR1IFb/7qGz+fuUgpJqxrea/gOtjrH6n0Bws91ooP8/vCwiQMe1zdhXYGXo
Bjg3h+j0QguehKy1Nytsw8iTmlBNxUcIhe43P0aSbKt3UhIeGdUjt0fBU8zgoyZb
6f8FUlF+opXUPKsvmgCAiS3JYgOxsgjfHXkV0+rxHwcR4PKS6pfQTuO3Vc+wt6RF
dCvxJREQ16nflx9be8rm96EsIHcXA0BBa4xSWsqeziaeKVL7p/6LuK9v/Ljb6tn0
pJgRQvbOxQHSOJmq3PKifvi0489kf6sCmKIsN8B6DidLkrpp1B/DhQ3fzv050vtQ
v9FKGGA6E8jxT1iOAzEnmS64yQAAtKpJvjeXaOB7HXQjuUZHNI1lNoOEplAgPgEf
sGsmXAQKAqizDClP+pzxqJqYqXQpyioLZQItIaVElcvzBw2E/9vx3APScGQ5rIGF
QG+AlSyJ+2F1nTHtJTu2Nu+eAbsyC2AMY61SYMa7eevgzW/OETYTKMCh8lcAjrRx
HlpEIQZaF7BfuSukt2eHJtF81O/e5MyVDrmR+DMHY36+AxW1HeU5YZgGCpEOCEVV
WlZf4N2l/p5gP+lLxX2exSF77Pmc0xjZKQU3ciMNVR5GYZzgccqV8VV7TGc72FYc
EDrTCLxREThz7XGNRJKmnJTBXR4mbmxcqLI+OaQInxy8uUn09776YfnJsBFxbKhI
Ov6Ms0cmikBFK3whojxklkpslMoJmjmV17rHSG8l7OogXifDkZoG2TrjU3Ah6Gc8
6cc3W8dqNIMsW92VoRv16NSDGTAhcdbFvK4Q01UpmuRNZtJDxnxYo+GnaoSt5v6H
Z+O9jaea77wCS4ZiMSIj79Ru1+gbeHwONI7GGf1gHt3WUeDu+8WZWPbuVN1cUwCZ
uhFQlILz82FPTRiD4pZQpTKfNMsMEKAftEY4TvfDA89Cc5Re0i+JF4GXYFVYNy+2
DTu9JbZgNB+USDbZx5pt7oHCf0cc1HP8nfbcHy+qqRI0aaxXESVDfA84jhQLYFJU
i4OVH4udKgHDm1+tetoJVeIv1noyYnGhGYSUxF4xj6ezKlVm4ZUg6VeI1yMiiEWW
tsWgCuarIH5ESkHyZgAhT/sT79ezqYjF+kWGiH+D7pEF4c9hH7TG++qA4HzJEBNv
JWBcXCcMWpZxdmQmN18etRSBOrS/QsRKUo2iVgpC+rtxgXIdVVXlEZ3crtQqjO5V
qBHGAor/daFbDD2JRkqvnQa+WgIkMbyk2Z6nYBAXGKYqr50V5M0j4Gi0ND44R2HK
4o0B8xgUPBlC9uv8BFxGQ0oJ320ob2KdH6CVOOghuVUyJwXDahD9mrWvkCKj+wZM
cjl6irEULnfroq4AjzkqJSfBdQpjG1E8X2RQCfEP+OnV/ATVbtNbBYonQjKUN71z
EJ/01EMHZhdaIdtu88hDNLs3ZLDG18yFX4PjdpatTUUhAdtijYyR67i+GO0o/VRg
WX3a4EaNZb7tbLcr2AHaopQ1N+j2cJxfYlEm8EULRhp6PR+oi5429m2isIrRqxx7
m2SAMpdW1ByPRMMSp6azSqxRlXI1M0Sd5N26VZnqdZsM08/Ot7RaOnoGGzPxeav0
A5SwpJFPYc2T993+yklFbcz0kzXDLbFTuD6616evaNCXXMaNj68qeOUmH6gDzvZV
p87ZCysWMoupSMczNx28vDC4Q69fEFISvKF+kOPkPthvruSKMBxhsJ8vR3VS5bSZ
suZzczSVVxk2VvMrxx63hBqguQIXKSge43UDFwP5nYiJ8gMPsLle7HyYDFxE0Ptb
AOrTP+OU7r+58TaJCiRPfcWGTIrfiEFz5bE43/TUTzYsQqM9l6opk1XyrKJHWYCU
wknD2FUWIJtcJNtb6cuDR04RGhigoeTo/Y72Vt5cZm06deM7cud/1sIx5tEP6qle
yEJbqeqjioKbmWXvLsf5SAvmbaldGLsUbtTd7qo3Jmv3HxjKLC7a+LmVWZDdyZuz
0IhI00oy6vW6GBJb1ofg295DRne0rs4LHr+bnSZyMbUnQRKyUlBGvplIUcEafR+f
4FFUNPJ3lVRZJtBvYJA1yViJZ2l/FKLLidfdGz61YSEvp4rITnJk8gjM/x9z/4od
XQWCSIHjdbZs3BVMVsV2+1h3rey1K5Pkwg8ehPGWtGbl3r3ZTgpb5LN4jRyUnmlW
S11UVl9fPA5iU5B9g2J1sb39YCC3B5osn38NENJgoyS5Otvu+xIGoqlQ2DQSKQWc
2ZoHoEgELHjGDE6TeM38QjycOvXjuUkilda5q3ALZttWywwpDvmUhWy1jKToMJUT
CiYwZdjwwOWKDoXL2Ly0p65y52T/6r0LL3RNPAvMFR37bKcLMVwqYv8wnyopWjeE
aUFaXVp1D6JyrCuPxbodgRBfl26pBbnBUQ8h/WmjrTA2X2tngnqdbS0pbKuiAyYv
TampQYIjVmk1Ou5YqfD88AQLvCeoqemUCkDj9Denf5EjBngzpVx9WCPOLhvH8O8V
N7VrpIYHZF44pqrOs062HtLfamDZeaIUPHl/o1ucgozIAUBda5TRhQI3qCq+KMfR
7Cx7MdG0L5Zoi6C1FlawrY31Jh9NKz+pNDsmKNkYnu46/umwIvgN/HwYCoYtE88w
Tl3n7vjOmsGLNaMvtwpmpzcWo08EdhsmGABYywoz3Wen4tZW4noRMOFfsIpZxRN3
tHDdaTVa+MfTauasS07oID4qI0MI5HcOCWf+MBhewfYlY7iOOl9DkMILu9HyRQIx
xKfkKLawuCGK72gKGGsx1mkqrE/YJcsPYl14k82TuAmnesSjsZvcDjYD1I5WDC1B
ZK43QRtDUK1y6/VhAwDECAUd3KbZFj6FWSOKuNqNIFQ6pYFmfunEq1ty0IascZbq
7KgyR7K8IKb/mtgsX9rMHqHtV4RfyavnR5StZNptJUXRlw4ww9MrZIEiUnN88lET
d/PJF2xOrdMruV5pQT73AksZhq0bHJyHUtKqeSDDLIF/ekgETqqTQhcdw0WAtzkK
c2yQe9XGy4p66Kq0HOXZc5uyXvJY5OQ1xVkz0QfRRpX3ktExTXeNAoT5HVL6hrmR
4MPF42oNcSr9zo1tZ/ZY14rMFjOGj95LRhFPr17MXIMwNNwQ9OLPx1FxzjDfQu8A
qcbsd9BIwdRQVxY4ypI+HHN9N7ETDzhlogGLmTPUK47vl9fwlL7NWiiawleOQ39G
ZyksY/JVW0HHcaT458z4+uIp+Sxw+9fY8tdpnY3TLf+cv8fm0aKdvxfNhvnnXtvm
Sku83tMelRJwUaNT9xgS9wpZZkSafmLi4VikabTorGSzOt4n8HwXcjameZBh6pBv
OVreyiWjoYKJn++f+TZ0i6cm/bBLZq+/z4u/LmBwLFZGTV48cUgBG1uYSAuqATzA
n6QB54LF48ZUxaYgXiRl7tiaiUWU5xuVPfLeiMMEJ3SYtUvLFBRVaEqjgs6fTpxy
XFzSaP6icsP418RRzaeO1+b+rQotSzsEdIZ0IQLVJVoap5ccWVp2Lpfp6Ji6njEP
Y2a8fdwxlWmB6uTpIhex5E96cqW06bYYiDikyltWF7KU66KkGfSaTb5lpofb6b5x
a2veKxwPoWUzqvDMC7UnC1MFwb1anKWB345JrLvqS75w4BhnoAw+HSBykjLUAug3
P40/GgY0A/STArTrn2e5OwzMScACR1YfVi768cgjsbE05ZDK3d25epXEPded0iEf
ASSJSSUDmNaZBZ6hruZTkVr6NaVg6UBWwY9hLmGNhvZHt7HGVFLTfqgPSG4U1RzP
jKsJx45M5Oez2ay3fpafbzmPdNRouDwmToaQPWt0WJHbQzmIgQVm91PYDotO3MzB
T/aThiPspBKvKLTXd1QcfwtMmZHm/42ZgOdDlgHysOxsFC6L8MvjoJn0sai8H5sL
Pk2rPHUkUaqF86clQ25EUfKfPoWuuB1eoWQD/UkAbxSsa9YhNTV1BDnXLP4WYYsK
OFh10MPgLVuYl/9cY7BVQ+OGpAuILP+i+JCc/5C+5ls0OuQxdFCHzqm95yb9KOPx
8g8kwiqUdENt9V5RWrxPuavmHBEwdjtYsG4jeFFRgZMXj/tw2e/KtL/SsqS0X1xi
cW7nnNmTQrrUSPkWIr2HgFfhhdvCf9Ev2/6+VNkH2Q3RZAX0uAIRqhWKlXprCHG7
/pxOeV1sAFddEEIBp20vd5gdbsNLruOxq2srRjfUY1Ru4CsqhrDRdRpwnS7BMyRX
Qs/klPUWdgdvSMqkEbiOw8lis7rXunOJ3JO5BGSIYSmZij0LWAxfXE/l1A6fc2Zk
MV58WskSa+TUnYlA8ev3Dmmi79NkfoQlGvYH3L/bkv9FsE6mPoeRlw6dV5iNuoPC
4p8HBlaLk5il2RhGV3rDPqM2HMNyW60uPbMenA6vBiPf3YpTdAsP5/G6+f+CA/BS
S5O43nghXgoe9F0c8cB1UAkP6HwzMawX/VJJwQq+slw1D4YYqC/Jmq8efSZy0HzS
y8J/ZA9FD+YxiFqcpf+QMmXrG9GF6O32GEsuZauId0mFBZK1bO8UhjCx3IrHHKth
wn/kR6sJBXsI9gGjLMn/JL9uGb6Ms4KFMRkKcZg7KVa6ESdqvYRoWrPzLnGgpkjj
qg2vMgqqxG1mq6QGL9aq+q3t8ck9Phy4EVDatE/C5CJ4CglXFXHRmroRCvqTSHSK
JEmyD73WMaT9nPt3lsc7OSBvn6LqnpvHvSNL2/cNuyT38KffFfAYFMbXjD4lBEuH
AlzGPu+mTEgZJAAWo4LRGtGvgX3l60kixZMXwDJGZuOC3bk20/uP+WJckBEol4JB
u7S4fU7mJPmgOPDd2M1Pyx4tVmntu8mWXYA8Fs7itSZza/rXsIkOLkUQ5mMaFv2M
sj40nvWChQt8InGI/cym9RhvQt9UDk4i2jgxPj2pLSRodQHyl5M/s417LTGWzwDf
87SKGOv2p3msWi/4uNUu2TiAgYGe4AafbV93yaYjq8UhkD/Hpf23v8ddJRKfXn1i
OtamGBahlP7B+qozRoNPPtQxJx0hkFyryVVhbMIH8APz6jWnwjQ04gDVUySdLPy/
1T5d9v6ToggU9cmyG/YijZ45JAamyrt2q1qCId6Ls9yVlRCxMOD8CbDmdesJoVVY
u7OYQCijtzwfaLzSnQC3w4c3PQG6on5buvSHjEUWLHpGFqYAazw9rvS9czi4/toS
tZWF7Cee4PBJ+LLhpasuANc1Xu9pMskrxbrrYhyr48S5B6q25ogzUncTSyio5E6X
GEvJ9AUBgswiQrcz6q6UVh5TPugl/+ldP3CZ18zJX4ZmzJRdZBQ1dDw+WS6H6QNY
GYL+ZtnTRlGlP5rUplj9A86HKdN0v4zyzYgjb+wXshKbPD1AlqcDuRC4S8Cs0/7K
JNPyzmvI2hlFKfQsD2rHmCd10KaMioO1WLzxxIXBKeKdI725aFIXpjP2Qi8h9TDf
UEOdIK7pcB5nwAKwIpvq0bIcIMMLgEDhO0s6PQYR1oEGGhs7kK6jdDAnpc98UHvg
LwS6HJgvZ7oOdOIHqHD9+7NXoq1BwVkHJaMOCrbOpwegltwnzCRqyiRi3UoihpKu
A+nvgVavZuwCS0UKaxpncebbXM+tTzLh/MN/WSZwHnGHDgZbreQpXpwCljftvxpX
LYTMySmYgZN+pbAUXWMyzi/nAEk9SpeCq/2TJQhKEhziav+3PBjm44ifP1GmxQbt
ceDK5TkN9rckcwqHeqNa04eTO8goGiwSufCiP1VcDVx4a0osf2VtYd+jr9m4hsDc
p1M6wAp9SfqK8cIpkOWJLota5RIRik9iD8L7kt0VCTzA8LjpL0RJLmHCkHmQxPsI
OwGKZ+qiTVYhAjnze8Xiw/p2IzZCjKZnfZDNbLRURbzXo8qLP9CTcHw+01DyMZ4N
Qj1vkd/Ch8YWsEQTTHsbcyCkzCAdEcVVJ4/F/WZrESrGS2XsFTTWjp14uTe8uvlO
/g78bzczuhKXn45lqMGDITqKnffeyUrTI7dy60akTU9CHVOCc38wfT4L5YwFyXcJ
mU7QBDTjk6Oz7xlwFaaFGNpwPEb8Nk+V6SAsGeVMjnfjkCOxj5k4ZqK3L9WBhUAo
f/YYAFx1Oaj2kSj5P8QBmXKoo1UbQLU0JO8g1bGXgkdTyFao29PN6BZnUPBWMM5X
wF9ovVPcHuNbZIBMQ2K7CqLLC7KxQ4QxKuewKwo3yvoCFhNLIrpfyif5SdWtSsH5
HDOj8ntJRBUG1sjUafQATzvT05uVGIN2IF6cGmTACH3eizCTfRIGBk3UnDwDa/ZO
Q1Ui8bZ7fnKR5NsdAS+AQ6TMV7jTWWzGwCLMtoTOFBrtvCYO77SipdUrsklmr7q9
T2m75Hf4k3xVZUIXkjT+dQSMcmnsPpiWKDMQahXfV6ZMLpTIUksvlPrtu5R+Yamu
T/JRz6vOECohBn9XR68Cp1H5s1kJvGPvixyqP4i9G07Zc0mt4sDW1POWhpPk2Je8
WhuL5AH+D4uBWnpotLbGbzWWA9Iga/pnymUbc4kY+0EEj+P1EIBogqzOXwqVDexz
WYboCvDnFUVISPc5H6lg+HSjkiw3wofp9ymVeHBJa05pJiq61Slp9lPb8YaqU9fd
2mr41KGC33cfFxpiyRO5GShihW311VICmG78G06rdmZoDQWUEQ581kOqFsDxHBn3
JgiJYAQbcvYpct3jmoWwXNfIJW/4OUwcdVoYDPnEA2ohmVtFbMpYKjQnmWmMvI+N
U8h01q9yRIINDIv3bW2eHsyCvW8i0dvqTwwVQTc42zIG3lB6s6UsFzZuod5YB3eP
z8f8tnduPyV56Zvd0IbDHrz39H/HfryPyLmGQaZDglE/dZ5EJ7lnmJaQRMvsItW1
stRP7eiAdW/haK9WC0XKT95hUtypKUOY16dwXgCYJ5Nrt1e4TrQJUwiW7jZ043OY
WM8+zuLV02+RUk7/bvlGMI0DeBgfeONGwfQ9FNrpXWVFMazOvgKtL56rgWsDrAoV
/3pMLzoW5v2ppPnzlTZc8Fii14U4CYKiVQLJw1KcTWdqYtq2RrLykHT52LTXuqBa
ofE3x7errLvm0+nnNJ8HN/VYAGaIvxtevT3PzkcC+PFyCndwLpLtuYHhikG44JkW
DXfZVGoWNTPZkJrwltySpnZIDmMRoA6PXFoGtXcwvluQi+XzNDq34hMpaQziqmM2
eSxo74H6/Cz64b39HFf5yBsdLJR3VZyuFCd/aRDmAmJrvCTGZPc/XXhAe6pqK2bL
CRyT9OKLhusFUEs9nGFUsL5bWlsAb05YBnzBRW9an7IM4W68WnTIoadHxwC0+Tc/
vJuQzxaB848kau0cqL/401cMGKyRqKH39kS0nG0RT0Nyli2D07PMBLDqb8NVLXvP
w6glwnWb7KeBz8XAXdDwS9R5OQgHsVtP0G/jfBcO1WHxiUY6lWM6zzDYTPiznimJ
ZXU8LhsT48sqYOVsHxjz/cVfaICYsmHaGH55etWUGNjsggNu1ugNqCPRAUqvREt0
+aZ9hMr8Cinci6aaXXh5KYEIomfmZLSOdKN1k20HrM8s19wHc9A3qHJ5RwlgOFpO
DTxqP3oKiXP8j0CUWI+fdfzAP5RsuYXWi4+XH4sqZNTAQd204nU23il0df0WHzKr
+z7puOjwv3XNCnZhu/XC3vMVjfnOHNSbgQ+/dQihlJY7rcGTMc1gPEHWn4NFkqOx
wD1aMM2ADyNEQmjhSU3UsQzPyMSL0Xp0wSBgVLbd8CXuFwACVo1B5NEEcCVftN3g
mmiOz6T8Ia1ZnX5iA3Iq7ISHWs/ZoQai2T1cjYwOR+dTlmPJ4Bw0eqOjjcw0GlZM
+ielHXXB4N/PW6F0uc13/pwwuLvBFiLS+ilUgVGkWH7otY5rPRDe7SOLkMaefvRc
HW6xoTzo51uKFqnXJNAz0JqxXXmbXH5rFBQnysS8MFWT8cl25H7uSF92G8XshoIj
fpFfFTuIs48G8amUZwIxHxzAi15Xzl+nLGc/7uIpe/5yo9OGUGs5e23tRXsxgYhC
VJbYZJP8sT7Qmjni0Sybh0gZMevA8uyaqD/6vsSpD1+iM+TcPt2lyAy0HPECiSbf
cOHrgotS0onN2jO+QkpBhVtAYxGl/hzGzPgbz39ovyGTKq+E+YOSiNvOKD3UTvEN
RHXl4v9a89EMbL0A1Wnl9qr6MbIvpQW91oPpkjfJM4TCRXe94oDi01T6Ig7qRWDs
PrlkKbXMKWSwaIO0cZE6nbaBDh3xsF/QGD7WKsyi4/YY3SJFbspjENelpSwP31ly
LbwrhKQo5qOQs3md3vFWHsoxDEPOEc4mNk8iffA+QLN/xRZZt1gN2zpfgycbpGR3
vB8UxwiAKeWdwsWhaeqRH7VtHVPDTwU4FiMOAD85B4/RZC/gVQcnDJK4ek3ec3nU
jz3Ss0rgkenl8bqPLwLRVuA6PaVRoQ+qzQyIXR+vKAXpZMJzyK4ObPUudXhkvO4v
8I0XYdnPMz0SECVWmAmCzURbRzJL4B6NNs3+ToHjg5/J8wuAlZjMBHpt9aJu3vaU
oi7w7x4V3UxScCvMfaH0+TRucCJgzRubF2QnEDEUIM1HTu3osnoWwj6ZrjQAgsYL
5U+HgefhDRiiP0PNeME6ys7QHvF+Z23BYbSB0Yd8t9I8scUH6hQgWNemdvKl//k/
vPhR0TmXIymjeArSKN9qn3/gJbkQUWHq0/v/PwdFKdQm5oZqBK4QDnrThYoXhikQ
fbmskXzk1l26KDAq2slFZiwsL/Xt4uqaf4z3pA9mBZslZ+E6/37rgBHBVW5m8uf0
VtLwfvvEHnMxHkLj4PJagXhmi6TaEv/3+Vd1EpCr/pJC8mRsIAmYBdL9+xG1Gr/k
8uCjchjc+zlhyTSGRrcnnC8iecDYXnjIUk8niZ2dRX8fjpaXfeT/azQK0glldvzF
LP4xdPaka1fBOpnxXKcGUVCbstNlBdQ4xesCYL/QOuU1IwTn6BmSfSspT3l81kQ3
r0d1InkGvacXLSz5OxY4NKHLPjmVBRUURcAdY5ZZ5NzJKwKyIrNq+4Gpjwgb8ugo
QN6YQM3W4LuH/MoNffKFTB3fnN9nHM0up2AZuZ6AxH/NaSFqYTj2+mDT023iACzt
DpFwEYcjcWU77sQc1wOy/ylwOVG1y/rrfBGCnq9PjokPXAkMksGh8VffoDakCP/I
nTkzhyN0pGiW+HIPU4/K8PcwbZwqUIcBna4A6mqQzYPemewsQ1opTu+LqZ35zqB0
h+0PpFpJrNVZvktZJtx1oiNi1mD7AHpVnbgehCoKeBQpN7JkIqzogrBJdhMhVcDg
NU4+5fLez/eaFF22B0D7drRy5XC9GD5i8P5QeWBhRs2qhgKciFMSTyrXutgLwQk5
BdPFmw61Ib2QvB/BcktRnlZdR2o5lQPe4rmBUZ6vU/eafUvXdqczGFQEecMaIaGY
QI7yNBBwn5KEi2IyUEp5L3IxtcIC02GZNh8Alc16qbGOvaqSWE+A4YdAdNe/Aex4
SKHiQ5FvDxTFPZJHroWBLo+Ms+MaSgIxgfoyQ1cqfv5ip0dUnNpnxB+rSL3M5zeL
cRbheGXfljR4gNjowNlHPL7FvZU0w7yVl1l97kam1MEXnsvbonp1wUa7NhjAoWbv
F6LegasFBNAya/7lWnsrCeItFsYGMn9iaMmgI4cIIil/ZqJMeDzfuhKEdAYxYD4G
YBSOgc77JU3avXOL4TrQLO6IO/yrqZxmIvqyGoQ55R5oPrEGNiiPSQWY5T6MCGes
GyG6+nvtHolPyu4lLxLuBDcBXuJmB0Q+Na9b97EFXX9DQMijCpRCO+YhBywJ296P
zBp/LyW6IjN3dKADSTtqugzJTkw5BO58DUybuQJdwuMOLoZbG8Uyv9M4uVRQ/vil
B763nrMYVj1fkeLCezcJbuVOXX1XL1xFrgALujaKf9L8s5U0kPb8WN0OPw1HPzSt
XALIYdNLF9/Ut52qmMpVHbUAuaBbavXpaqB47v62MdD0GiOkMJ7O24ubKQdpjWrZ
YsGTeRlmSRNwFvbDsdZmPSNTjCSFl+DHjutyd8FsoMd3J6RRDVqeBk+nNQZ7DDAD
qtNWEgYmjec7tCPJwbb12SYb53/e/fXs7Q6skqRVFNV2zI5llI5zkIUxZ/Z9IY0X
zS5+xOfzdjC0K0uApiC+o6gd+CK9uPn2rt4I1WS2AgBuXrhXIhQ3O4R61sYO3pQB
aV/X639zudkndvkZ0uCMSbnBxFkX3fhjL/AlDnQgUtvqOmDJHWPyFqIeq4zjFg0h
1Ra0xkg7VO/3eNoEMl+kVsYsBSLuwsTaWPmKDgqI6TT1cpJtJHcaispv2zNfQ5NQ
opfrEM6WQjisuwB0DKDsioRjvXfYfYPYcTqSvfGGa1PlbdFoXCGonHkvpkcA+smc
ZUduaVqEVaiAhMgEY5SL4MkVtWoHMEyDCxCvZVarGVh+LwWTNyCRS/0YPTinUzkc
KBgex95Cgr+B5JjuIHojP2RPd/nws+FGmMr/dIOXwv/jrKloixKdto5phsCuyfEa
KhlhD24sht3JQkzZB+n/JS75hj2OJTv8aCvcCt2zDpwY3zGcob7BxhPu0UO2k+wF
YftG1jdQrTDYQihP580aeOs+dIZejzVD7fK26wu5F0EXgilHGDTImiWjEhK+16kD
XmwsHMl8JAokETxhvqvWt6JUITfoh6xV/j+JV7JAq87Jo/9HQi7U26pI2qMl8gE7
dzuoda0u8bu2oeczkoY4rpdUrzdPUmcDlk8mc+P7XVzLneseSX/fs8bDokBOePs3
cnWLts+pXvE87Kh/2v4WhzDYXY58zlphakbREiLvwf2fZMAdjIBtNPoPAATOdv2O
yjm4xd7MBnNYQzgDxYZczZ4VquLemQ8uHs3gdKw9CJzRzCe45I9EUCDZZ85l/4Oi
aJRzJYqGrDdUbU0m5PodDR9RoCPV61PUcB3M1U0ZuEDHaH0+G2R9EbVsAu4arJ1n
VEaLTAEZt9yt2lSWJo07NdvmPjk16Dt1BeOpeJXF6I+v4Q0zll0O8oZj38a8SXwn
fkHQpp79+utMTZevrQgSyAUH9A0OqJUGajTsNh233J4scQb2k4RSgFxGZhp0JN0b
hzRtnZnyY/HmS/Qt3faRDxbyyhnD++RqmwTg8DRNCwGdIOrKo57BqCxYUzJC+5PZ
QCK2CtmwDeFAazSB7wokBpVxrdpGmMLgM2HL8SZwuoqTZ0cwn0vBEF6eine/Cvs9
9xt7FemL/xX1thoOodLdm4LR2piR5UPVLqkEBoWs1lABoPqfRzgZ04bP6NIx1+cb
SJJzkHUf1zOONR5jkr+t3hp67jOrCUQJ3Eu9AahSB3K+JXtW+9CFtgXS4/UQ4qk6
QQuLn1Hy/T28oq56fecjsfnLYCF0mSYo/oHFZpBbLLQAtI4BgmDSytlEtCMOY/R5
t1CoT9DNbdgfEBnOTYKRyh/STCUHIbyGzXSnAPixWTj4oF3lA0m1eKQokN0cWYl9
DXVypqsQpEWqF5CFnWJnUgMYyCVk7XMAFtu/jy+tlU7Laq47VYd2xU1jOw7IapVF
HlcQnGDFV4ybHl2yOFPZoz06/oU8rdDsXsWdNBmJXRp+LWXo0IMj75x3noxFTqDG
vYiGcxdCsgMbtWRtTSCqktI7rU+aBitL2rVo+t7lqMVfo8GZjWLv3BOYsTSlgjDv
JbhHSLojw0sFNaWuzd2kRSaScyU5s+dB2YqpOLmbvk7nXvoOmINrZ7i7aYkzBpDi
hGO2lNI2X3WG0/aJLhv17TEYK0WJ0V0GBoAqRNOtifD82AEyanQ7iWQTyj/TeL0/
OnWLyWTJeccKy6F2IpO5iQ5VUhQRQToqnWk2oF2Rljz9LHggM4ZGSnLyaBEXg8xg
1dQTIRq0oeNcjgkLcRodRrPEOfDWZew3Wy5SyqiblWXplLXE3fuN1tBEgirQIGg8
pAQ/uCewQWAeYiVxeGMJqIeD1jklsM2fclEsgZi/+M4UdmopzXwUz4LDUuIlg/qs
lUaIMB5+I/8kt9/kLSl25hfRZkEvTyfymMy9zGukl/DtfbAww0IjWce66JgKH2zO
BeFmzzLjSdVpbqazjFqilVX18VELFHhb3oe3ifALXIrjswQzCq7FzZi827duZyoH
EbeywbrZ6pwzMFWzuul7O9ESj3dY35xie7gTEDxtC9qC/7jty2WDFbNJ8O+Z+OdX
L7Hv+tecgPPrhYhDO6u4uIcKsboEhU3C/LKgnoRqsdk8h3dja5xpFIQsonaNcf8L
pKb8Si93HiEOc3nsYOABqYWGWRb7BSaaktEIyC6pQ2qKUKhUFJSJ5E9UYHPU+E78
LaCQqZNxPt+FHGQNQ1kXTesPR54LXltSMoWn7NMyKVKLEhI9XrXtzFkg9jtEHDej
3ZQxq/BJiL2cs27ppm3KyK6yVsHptixsvpuHtNRSNRhsGLRy8yl1zJHIAXzPabFL
uQDWZPU5Oj6lVZaiOYQvvKbm723iTQcXq5yzN8IqDZ2P6QmA85y1avY2nk/x0T2z
R2l4Z1SZ9PSuRX+0p2T6zp9Jn2GBxWiGpimh/h2LdlDsHtS3tT8n4m6AVSK1PFtM
gPX3avQDKHL2W2jrVAo9ZlzwI7ro12vToEXX8XU7x495ACA+WILAsQA1VqCG7cEV
IAhmbwwMlhUUr7QZ8SkQ5/zeUwbnc8Blo5NUbfBb6AUwCxhhEvIU3Y6hLAj1UeDZ
mxebzuQMc2mWG9Y/5fwr09Qs7sQhutgiMGyBLXOftb+v4VFcMSb9IWWTbu6BHuK1
/oQtHZ/a2yCIk+ZNSVpS/43o5IjNLLEVd5InlejVw5w6ai73BSny3tbAE6l8lkiX
GfJCEf3tprxvD+mrV0O2Ve6WyVQqCxcikvaJ+BNUh4aNB0dwS8GZAEJLcvsZmgJ+
BKqnpTmov7xCMtjMAVhKH2kBOfDXqJp1H4pEhoRECgX3yWBi7TeQnTmLXoXwH8C/
ppOmpI4tSe0J6HNFfyGO5C34wz3lIhieKW958A4RXXEcR0ecxYDezdZ/u9eURdrO
p9CiaZB2IekNwJhoP8Q9yoEMXXngYDl2LYr8YN9F9nuLnTtS0EL+d4bbUPAjPjxr
jiDbLcnrWRyICaMo9n6sx754zAEwH4S00lAggEcG1jUbkVjKpumO9u48FEB+oICM
waEpxJpFjfO4VZ/oT+bSYOJnk2kr9ciw2VkfycJYarqOIfkAkfDL1WGdQihlKgq8
sih4qj2EFuDadNxkoMzss6HvpNfxIp6E3xb/3dWSzhsFU4/J4VxVd2ikSp4XDeCq
wnCOfu8ZtX0R7EvN7vHw4XCm6AaK7Dz7+vKMnKoltE19t+FvABc+/+tgfyzlaaY+
fULjYBN1co7d75mOT5dGNqRAuQNyFd4roVIFF3pj09wz7mG4btx0Ai+aTUIGfDMF
Ol9lKN53qKVtWU8J1EZdu6b43v+w8BoT670uwUYgimmNNuJWWnNvzdUZvw6jefoF
TwySV5z+Sy9qFq8t1D9PZsR8udN9ULR2yc3d5PtqVEsKq6mlSoVfSFZRaW+gnMvd
NmPe/5pzQPrF5CbXvLoyMIoY5HfPGwU4Klj/rDHpHOAXBsfu12yUAtPMJlF6KuvS
/T1vLPOdxzZvUtco5ke1I5UysCyHSgqwR1uSGKXj6OWgQt/Y9y8x8vsgYXH1BBbQ
2IUtpOAYIq3BuV8xfC/s5vBfrABpac0T1Md4hdp7/PLUNZbO+NCc+SBojFacEJSC
FDXIhDvgQdsyhnvMNG0x3wjw0YMMSg36xmwmOI+HQmsA8nGFy9Hf2X3zuSVawzja
6PyyOpHYYRPIWm37emhH6jSyfrqkTmFUfRSfzZtIWT0c6oPp2UI00LWCGfE1Sw/z
GQi4AfID2pyv96uo7rt0psr4NAjWUyq1ci2a6/t+J2/D78IvtrtXyKal4fhPpII6
eDvjcI/ab70E+h5xlFwleSS3CwHBj7Lt1P5BfJATmHMP1u9Fr/wWvMjgjsdNwhlx
GY+oq4Hygf0Ey82380QpBaOJglGm1hu5tfXiFxj6Iwbgn3ItEPKTOoEzZrzZ5DbP
D9T52vMQ+wWp3ID3SmJ0JsKcdajWtwBT4/oQrw9XFzhv/aCzgixUHIV1x92tsBds
lU3gcJBINDnSrZUOnt+Qqc+ovgEx8Ex6bnMERVThPq4IuHvJ8L/0wV7PuR8bCCNm
umcJLDMV1TVxr2O6OLIW4Dy+5vtMu4KyQc9m4DUXEVePqDMEfwE4cjEJD1EOFZwQ
u3c3iZ+pFNeLz8rMMvti1iJWh4kTmZXARJYHERQ/US2NL8JjOo9S+4D9QCDcepo1
BYwuUNLRRj6zIAfxu/LbPYRoMavIoICZhEZkTyXDloWV/83YhYvbPir3D0ppd6tc
Lt+qoE3lUaReBfSFMvINaGjbRHUTUnaDaqOtSSSLlxSnymct3CnHStcVnhmtTRDl
tHO92faOSls7Ut+JhiWSDZ8FYzDh9SJAnij5RtssJJCtTW6w80ohro3aS06OdTo1
IWiF/XEyVZ0imZq0q/sKEM4rrDI/khVElRtyaxym6IORJ8oNp9gmecjVe8CA7u06
PhJWTuslbeYMyHWgBFIGU0blH4lC8V+QM8vQ0ev+dXUDcQTe/u3JvOCdkkDESgxV
GHQY3JuZlnrAzr2tmjm49Kwlj+KagxN0wiSBhn7HvlAL/WhbL3pnzJpx6J8K6gL4
Bo9Nrw/at2Tuy09GGmIJoKZwa+qnkPPO+bnM7DZlACiOiXGvX28cC5+Nj8tnGXJe
Fr5wP7DZUhXtYt/zCa5BrG65V8+X3Y68BaLn3E4/AhwV1GmhpMMIdo3s6cmDZ/dX
qbnPuGVl0rsRIJWWeR9lAYKUUagA1awG6mtSUd1BetCMa+1Q1LhII6cNKUJtq8fv
SH9731I7kgAlaC+zSe71eJxWvMOgo8QSMVcoN8bbmRUbG+gH8vCxGHTU24N0lIK6
GNh3w6pajmw7E55pySqfig8l5Oc1ZNsbgRQlXnawF1qAr2OFculm2SUMqikldT+8
Y6p+f+cm0PTA/76NDDBD/dXve5SUGCJtedK9erg8TsWnVmvYJCb9ccK75BDvm/E3
2V2VtBkcHeWvebXuzxKE8CARBPcglqJDBCDb2xkZGfCU/8JSZHSLHQLzMFOChsNb
HZVBaepy/RzVmDhHNBXF56c2vzme3KuxL9TtlpbKAO0P02AsfcMGxwlohaXkHvxP
JpV4Xl//F8hIHLLxjqJ/tR7lrtZZdjR1uCMaszf9XyuTWazy72WJ3zA4roZY2ZE7
Pj0vt5LvtbZRsUjH16lM7960mGtFiSYirmKSvKcySHDufY3PcLvmdf+Uc/sGDK3/
uTaMpw/lnmPypvkTmVA2IlEdMoIvRuY/eZY6FjFZInySCt1SKpzUabS9yT2sybyy
XO6k6Ma0gm5I4E0xkcYcYYrlcT0aDxIhuQ8d2hcoKufD/YPrmv+ed/QxMOoVZUED
yqFVCGqivzrXjAqep7jmJ+nPL/Lu/2XHrJMnhOANWEpFasmD1JvVbau5MqC68XpP
WO/03SgDa0fG5k+FIS00xC/g0QTVDko06cWp906Ch8/qkdTLzlSpXOxC1RUaa1AR
Jj9dRovRdnhUE5NZxCSCXgbVOpuFRCKORDm9TlNS0500nqMdHcCphBYsu6FKrzdr
HmPbIfPylTfKyULgpmgslCQFDXdLZ5yZzAGv5tsmuxbFVBdWT6f/+bPmBOLSJBZp
mNz4NxwxKugADGb6DFqD/Ao5tXT4l6pK5inlCTd6NA6uDvGLHzhAUMmf+sOhIQnM
qhUSqwXmljVY4W3bGT+jnGOpJleuXlIySxVnFdruAU+AkVf6Kk2/L6GPMexxfxmM
PkLG8ecCxMzppKllyrq4YREmUMKsskQsGX2+02HUPutbLlqi3Z9KSdHAzAfwDzO+
RHRvVMkmf3wuETNimcdVtBzKy673uNWxtz+n5gnXm+zmog8o4DnYYpCQ7fFMooVz
Z0/KVIgrnqMyxM8AmR4pmxvb65evVSpniTi/KwZ03ttUKuafsMVhE8sjbhOCGsjb
cs68MwqfvxITDX3WO6YmUa951L6HCfo7lzZtdHLxmhGcDA0AvN0apOfghPGVH/MT
e1McriRSZqrhDT3fLq5i/YPu26a6xY1r5DUEL6h9AtXbJtVeG+jeufqSTSi0SHCQ
yc/mxNYGrjcSHiwH7MxiAtYTKWbYFQAfeVp+RcLSR89hxGuS6o9K2eQNB1vmohEe
7n165pEAYRd52IQ5FPz/9u9CeB4kRfqeuAtVOq8HAfVqIfhbna9EVWZ7nhIctlP5
qIIMd+sMHFeHiRn84sbaJFsbQNl0TlmjVuaBAhUKPRzylT3Kog0mWyWAayF5WQli
2PTm8d3orVRoEiIPWZw/WDjXIAvHReJLN+0cTvOKHDrW+2qzVoLjBBUvtZuHwwX6
H+T+T7hgPw29kFaWRW/xbxpp2JIZHJ+iMPbFp3NI5+mb5mgjwdxY9oZclilzkj8l
X+zGUl5I0V3rTDsGaunSDqV/KvaPV6qCE/kywyxRTHlFPVxhVSsV0c5BLnJg+X4t
dFFUHxwC0QCrNy2rlxFWuUwexpxUvq81fOlRIdD/Uomj+RxWdq/aPeeyi7WZ5Spx
3hPSeEYJOT848b9WQHGK9bFTl7S7tqofwvbxdtKpncn9DeLnFb42JXc2E0HWH/f5
uPoy6ZXVrqRv2jTZeeE5PkTlzLBJzJFUMSP20Q0Vtxbb5z72WP64DMFOVkfXZwVZ
50E2oErc3fYNY4wxx9XGoLqyFdcspBRwDCwtJgHD9tBsG1IKEqkDpsZ27T40935H
ytIrDlfWTNmWPCzWNM0EHRtJU0XKD3MfH8nfmWYXFuMcXsc0PjY5/MoD07BKKrKJ
SlwNpqRRezCB/DzTsdCiXc8A1cJeUHHSIF3wowEdJOrva/hLczJiyb4yLXUJejbX
Ews2Uz4V/Qx+H4Eo2b59ESm5p3HDQrRYGVazNqzNpklDsWSf8s8BSOVmqF2JJEZ7
dYp1BHGw1nFDJ+BgVNMCM+G7hHvZmx10hDANfcU/RtdUwUy9nmxp0KNlKM9LKJb+
vbIf74sT4kRho3kcWJxtbrDG8ULfNKX24lKyvn4m44Errx92NqzsmTB2qFrc7L7Y
E2E70Hxjk2BOa28m/66rmLf0YRy5bAYCMSBBZDsKmZLdYFnFSF8d3lVBwJC6Wbr9
sknP9kjW0MNK75o9OZypnWDrj6or7MJxrWEYZMGJv92+7A3Ra/5wAc55p48IiqCz
9S11zHZi0nI1rAjiHh0TnRtqGLanIFjE/wwELWFtYjypxCOi48A/uZcpG3ggRGgU
DlZusUvlR7YQGiMpYcjPKdJldt509UVGEWuQM9hn3HO/0jkjw97RLkbt7v8I69HA
sicprfE/CLk/ZDDvdndCT8sM5G6R63+di0f3AanLL87ZdY9bX6rFCYjQjYwMIW38
lxYK8gRSGYs5riyemNAj7eyMoNxJsW5DMJIh00a/e6D8Ajh/8ys/cGEF7ZKinWZ6
x8t9at1O3tz1BJnWjvk+sDV/oC7zgUqVBjsoMIYRXJShzkW1CE9+VuT+GOnavzeE
Vm2/tk9GkAHjKOMGXgxeUOSVaiBMnmni8QrUvJN0WS0y3IKkOHDkPpy56QC8R0CC
Ev2LPSWzwIjs6vctRUfW0IuSB7/8s3jkfcv7auRaTr+ET8E8qUoUYWPZ0pxqOjD/
uRo90OVl/os1KQ4YJeN1cLdIDYGeX3GtcH9Xpwebq2baJvWHJESDk8XO++eOlnQi
vgcjI6vsLKEbeb6A9SR2qlQfn8MkBs7rmeJlecap8Ln2h9dNfpRRQ/aCv9y1ZkX2
OTS++hpGmnSVrSKRZeb9dL73AI6o15xc3YMK8uOARHw5gOFw3G6hBEDG3A+3hvgt
46BC6he6BZ+s8x4WzBMXYZInyRs1n2YhJ1ty9lFgLMqTs3sCN4IW04EyHCNv4kwT
DmRmyV0oUYw+QRDnrV0fNiYSdd9NRAXirfekajtSo46wtnN1EqBv3Uafj7udF/3O
qiDX7pw1wc5rDPscEhbilWQBzdcBP3BGO5d6cUVPkOr+U8r6MKchZ0Gp5VSTO+mu
mdpDGthW3Zt1j1Rz5LdCLyaKwUDOMRv+fcH73XKe4Ld4l3GRbP3OjJCoFtG19R+X
SdrmYqbTp3mY1XryZvRFNrrsxJyr3CLZmTrbSPZAFAARNG88eHws+EdKRAu42l4D
n1Oxchx7bKx7UNJQyArf+JL+Uxd/xdYHGMYtCdxg6vNU7UF8ZSRzViwdujd2goFc
LLm1Tip026+tyKwHB/CDZha5XXrw9JH4g6QyMzJL1nIraXBxmuGfvrSG6occ+5b8
dL1eHtAytQnalS1GMB/xaMMufpgYQAH7SZYiCZQ8A+rPzXBwOiLYeugF2axIcJA4
oa+mwlbRX1syh0XvuvtNVyePI2diasSPo7XuNh3UuYAQGKb8pkS++I4MI1Kgv8XP
/CzFAXsrDNowddolJEuIZVICmahdMz8sM0UW+TWnUIjmlpCikojHMUwJ7zy1m1rC
WLmHW/XKAMwqLfFNtxygoSjWPzTUhl9PQ3otPPzIT1rf3C5n3YpAl7wBlST2Jf+G
Rha71wzmEe1ATzko9BrHaV1/Mx2gsMs1oJZiEoSnT6mPUxHKIP0HDx2psnzIaL3w
7NhFSoWRfHbqvC2mSy2w1lTh8zZeWE+QX6sDZuVXnwkZuwm+yKvP2485UqlAG/VH
pb5TlmofATMsSjHdUAbtIAH4TutBXQcIQntk96iDTtPidufoNiPI4hOKCaJW3/o0
DSkfb8IrTYlVbs2shjO8olSKJqy+uuDRgO8ElzQVNdlNpNNmd5iIsGhiYPOYSgzu
/HWXW7oE4InzJ/4s6YJAZd25t6d8BzmFTJFZZnHalYkveCdfnM0ZtE3IlhXfuNlL
pNOH2PFzhqt1iLF0J6ogo9G0pQgEUe4etfXwtwXfqIYY3z7PXABmnl1vqb7+9jYA
EjpGMVphdZvyeKloHfIPutrfqCC4Wsyg8MpuQb1DasXoeGnPxtymqZiEjDaornCY
OV06vesOr8rnP9C8V/7hgj/0PM0B5CVnl3VYMe4iNRM0ZhUmtCPmh5lZBLrZWsYW
P7lfXfv82BjHnNcPI6Vsv9kRxxlLdflXaoGbZSXwsPZzFSyMWnafft6BjSRRDVby
zOEVDG0mVuRbLxHXxw/ltCzO2Eg4T5V2ldCPa6WzKOSsJ88qXSaUaHEBnFJOijIj
MpPHf/ksJqKmI+T4I7p04eZTOWPDbQwVc9Nd7Qy4zUHqFU6pbiu/Mh3elG2MLxwG
Jq8p2jSYRXoUnT89HI+3dIYeVqMVJDAw8Sfd72jB/kbxgUXpFlEl9NOnfWT+1RTT
3hBB1upobEHfzQDl3mD4Zf7h53ybu2z6qBHpAZtM6WEmI6kEa+n0F12Bs+50SvMT
HzoIMsAZQsop/9pRDmvnpxB9s3dsyNxKgLWJDOFPiUGPxrIMkse6+UpecBazHMmc
oLh16TP740VRglS4Wuwu/PI8iH+wFIBkEj7YGIP0kqZO05yfahTprMuLF4S30VL8
jRErIXWB0KW/vbEGFC2C0u+v9gUEg7K0BjjErrJlmMUmC7Q3Qsa04HWJ9iVNcqFH
ZPmrz687BQZE17ub0Z00Bc/fbnSBJIbNalJfir5wW6fjABpbceZCrM/D1BGWJbmE
l5+354NpwZqT+IBF0kuhFlNSYsHAilbakKvgR/jnUDoQ4pl9Bt24kCkg0QGn2kCe
B2XT7/ydfNMxhxnwOz5rFF+E7MZGmpEPp2IIToSq5+qFAyEElos49GqRSBIW/iP7
TVrXE4tRJVzrVxJrqhz1DOlJibOhKMMnMdMpAXG1GvhTaHIzJHXVzHpUIf4zeapN
Twd4L17ad+eB9WXh1uyL8eWkc/+6HETJkDNJNr19jICWadcJkJf1j8QADixF/yZ8
p3ohmgRTMWRd5Rxp80kqnjQOCFz1vU5rZROdaLCj0KAvOymssPDU2g8pyaS+YQu0
80dgpQDYhsMw9Sj/3VbilQQ5YjDq7whkPhJtkTm5qo0+kY5U7PO7q0exTdp7Twhx
YQgdLEiVLjyPhSeWcYDxbi82Y5SG2lQLxda64Sd9pKZ2XzXyx5K4tGFx9wsj8A5S
gBJbpsqdQiRdvLa2qMJ+/tEwLAiE/+RQetzgxqUQ0rTk3v0IykdO0Kj/6OhrU6NQ
K4kWiskM3QW9OmMx2VUtulkqU4tQ95huEwiadsDXF16/IZQguXo4BIBJ+f+Aog0V
CCMZjxwLCQMllhfLjX78G1mcpbMAPleEsxObQQCgaov9sZlftOpZK9seEYrA77Kg
nkGdifdUp79xcLl6PAZFaT1dvwl1v36h+3VsrGYwRmcugt6xtyIKJvfrcuT9s230
UNo9cCBSFbFcMMBMpfyEM/Vzhre+ptReGkjthKTflIkGBmvg2ObGrhd9LV2tTa28
4/FIPvFzpDnEaeNcZhDSdnNgDK7p78Rc+tPcYN4UI0eyrNk4ZQeJoauZ7i5RVLJw
hx0yBmKC1eQM3EvIVs3ECQztH/OPM56oNkblgYysCksDUwfrgrzw3RmgkBI31yOz
LTRCpdKiiL8DNnEI2RIiKI/J4Dv+AGSgyNj3Exoy/GQYKWMlH2aRaI+XsWu6yDLQ
aT8fceOMOmLgPPuIzzFXQ4SYBTL/kI22WB1WeJoI+m6NZ9V58vDF/YawPh9bKhYz
mYebQFurtr8j09NVTrJM0sTOD/0/qvYxROw9+oWCNgiELOrdXzEvQ2/xxDd7a62G
XEwUw1I9QUD/pZMVnWjiK56zQ1JvgsBF2xxQZCA9af5/5ohznj6xeKkEJfxYkAkL
FEzze8nx/r+zL9Se1FQAYs0yXArXeT01Wf5/2ZTAUJcLS8RTXzr5nm/xsgRNTsCq
sobMIzdGXrZ3ATVHlqy1gJif7lNrTMPHh9ymzv0UU7oVfJBlwKMtxkcjH6adWN0Z
wNpApwcTM4UD/QAqENfgZb9lN9SA/cLy5gkasfN9uQX1bzD9slpfX65ntX6t+976
IasogyXa/WCZ35bxreez3l6GWNlkDo53xL1rG8Uy0+3BZ/P+CmWqBUDMffXbJT7v
tHlAD3iMlF/45y+tZvE5IhshuPYEp+18c9XL9QsaDdvROjXHXG8czzO6XhzjzlFW
CtuOpd1fhLiVgzW22BwDLDjwKrZ8K0AeHCoam9Y8EobV6JCQqG8e3W8vYhVGUjL4
kIf7rxPo0sKFQxDGW52etP3YJhMwAjm34/JKAMtOGTAlAYKAMPe92/UNO6e0kNEQ
xCLmKxTk0IK/+UtaFJUSebda4iIGUm4UZtM7Vy4zDRvgilwx8yOOER2+yEl6JxgK
WP27Pi8RLLqiagy4QcKHFXZ9Esf7qzkOyKiBOubASKc2es53Y9sq2X3j4vZDpMGR
cpclSyl/Qt6JNlrwSU7HjkZv44CA6xfGkn5BELv0B+wj5Ik03JGuy4GMUbf+ULuk
jJ8DeRjef7E3AMn6ajPp1C3OkE5g0JiRsK4v0r7kzR2x5whR07p7Iav8+rHvgu1t
9x/8b+oAm3I0AQJpagpc6CB9+Z9jDl0E/8UbGCLpX8/jGmmLhUwXfNqsHEZ1Xih3
L+5i64LHhnHa8uvRlFHF95lYPpWk80vK0cRAfFTy4GY5MWqbhNScMIV4L3EWPoQk
cA69bCDXs22x3pO63NsvaQiaWSaLF/1Req8UyDpBQHfUT/NPnGevy3dBBO5Q0xXu
36lNe1oprf8/Dhm5aZUKpGqFqakw9AU+D19irgTdJNQqSEyDfV5OEHsCwD1lq6OK
O/6ZJm6SlblfdPJR/ZYrh0Znij5X8vLAPFA3S9ArSjPd8ap0VBq4yQBstFuucJsc
2KwhYPtctB7OYjGceQKBCYLIP4D3ouEAwK7voor9eMZwa7GMl6qBsnG+UyQQ4qbi
Wl+zQDtxUHz9/S7keEmVoD6N1WhGLlHUw5GogyNmMQU7B7NRKS6hHjm6AL4waR4R
rVhoHUm7uEJBCDTlVKef3aGCxJznvO7mUd8tgNMAbXcu4+7NzyibZjICEQ26KRfB
uzP0zM0PKb+hU176AVIL6zjNVTSzK0wmNF3pFPNDHH9hyawIJe8Li/UbBrxAIRLk
T23x1mC3sns2v2fSRNvr9Us6FlTJ+S7x8xs3CE386DZ8tcZ5vYHqJi6kq5u4/g85
RT7rRDkvGf9EfWOEZdcZ4QBpi00cW5glgaXpmyPjh2apPrPCQEMtBW2sK8pYA9ZD
e4JZ8BZxI83lunBdYTgOSuBGFAJU4E+9K8tevp+buHBTIgK3VRBmVxRj3rW7RWHA
e91zKtjM6ZnmqpDJ3FVy2LIHfmc23NsrcluI/CQpQvWQOnT8+CixVQTZS6ch7Pw2
XDnklP6o5CXdH2jxcw79Kqm/CPD7GblQqAYxnPazcraSFE5pXohWvzkydAK7xmq3
ByytlQpTaJbOyLSAGmH05/d6ZelyHp/hbGmYpPfN4GaGKnbJ79Zk2SFNaVW8+JJ1
twKYsF8ZCwdiO/e3VNVDeaq3pIzFzFjOS25Wqg11Ezw0n+RHdO9z22N11d4U9H+Z
FpCdSZD8c6C4v7YGMtOBX2ib7ZLaCXvD6S6lqShnXlK9CSVMv39JOtJdHRhj79Jy
F3E1G/8XErjXcOPsLoVJe3/kaMvTWMyFmlBw4YlVRwkNtnpUoWnv2dloQm72x9n5
txt56YqUn5WwuZcShOIByrnmAfYaWPaa06OS1hNG7CxvgUe18/wuWLgjUf2T3QY2
v5JuE+qXUBOfQkb3Qfy9Eqmstr9i+6VnZoLwjil7EAUw0ulJPuBK8mw2isATnEN5
WnT0mxzN/vf4CVGjWB5Gz/JtgnmZ2tDMOJkyj4sc3XqIs9aho4VYTqB6T61I3VWu
49AO5i7nSOtL6ezxgHVwuPEs1scsfV+PQgwuObBZFKqjUrMe2i8DfAT35FToqZLm
8YA7OmahK2tD9+ZhXAPfzySnGwzBa7cwvF0fvT4Tje/rq9fNiTBMIb4/ETmO0gPS
DnfpnMd+A7iuTHFpdInoG/DCx/X+VS2Z59dhaXiHTME22cQWo0PFmZjtT0iZ6sjM
/GKCR4H6MX0SoVW6G0uXivCVJEm977cOHqlx6YOvC2QZ9WjnqHp/DqR7nryLj2mH
PZ1SwRWBeXoL72dZhMWtKxH4Wi3mhg9fBATN5LIE6vDm99UprN5KYXE6i9md0oKp
IqpkCi9fyvMOUhuQWb3MCcDhRerp5aV82f5E1BV5+HboZIP+a0Kd/+BSbq89loxe
whuJGurVQGpUo431BodyCKfD/I07oTwZLsx5bzhQyDck+Ar0wQQndtl654indi5D
0HzJe98xyyugDD6P8aa1lB13tQDmN4QPePptPKSQns9IxUC8SkfXg/wRD90/ScPK
/fY9RXP17Zw4jW4YMG/FFQ/CLHPtRGlwUSPcbwm5FYB8XQ+BQqO0JnvoFkVRH1+1
d1xfL1pOQJ10qmxePiL0hW1cPb1vziEi0qQ+S5D2q2+zBfnISais8Wq7uzKCnrdL
cu1AB0pxDn3kVs+z2HhhzuWY8ZIkJCgxzfiCbnA9/mzx92GPgnLiftGj8n5ix9vw
lYTkJv8hFxIhY0JDX0dgGCRM3HMTa2YwhdPpqKTiDkSRf0R2pPxvpkd37E538HeB
gsaHZ1gcksSQdrBRzjp9166HJTm9QPvTLbyaaDXNDe3LbsOuiXZ0a2+K+owXhKEA
OCEBeXv2oV/8v/0DwVrFelBok1lIUywndk5iB+yaLRdayItS8KERRK2RKI7sjlbJ
fzaQ3QYMzp/Xd8nkrwyoehBxESlYQv5tSOu0JnxAlOfYXEqWq0/olHRopalo76WE
+IUU+xZDuoKjMFebEhiM1IkwhV1aeBgBF1guZwGnFnrEtjICX32zKtrZwuRe0COX
NDxMBprMl164tPGPO5qngODksuX+ZmMnqdBL6uVfTRYBq8BPm237zhcElaH7UL2Y
O5ffEO/9Q/dbW+J0y0G6sP/ml3ELNK1lumT26V0gzQ2v2I88xf1vc95n/ZaqClss
4X1gBivYsdeSg7Sai5fF7rGayY4rqtSk83W8z3IK9TWG8m+A4vzNXZNSN2dhYohm
SpH24g4l+HMF5TQ2gZwvupPgzGape8FP82huRnm2WMCFj8wQfyYaFzc+k7rtenGd
Wyq8YdBO/PCdsxYxa3TxsySbKYK59kR8NVVdTsCB15QBX1O0tk2NeeH/ddk2YpGt
WGx994LKSSnUbFS+ZtX8KDaxoFavMMSk2KNwrvS/yAHpHwzU3i43k78Hm8t3kTQb
i/5UtfX/Fj3dRLEBCjeg+7lizRQWgezr8Yj/trPbniBoxFCln0h46MIJOLrI2Y4m
hOJkLznPsfyB6VqK9UC51AOgWHX+6L79eSo5KBs2SDaq/0mqVTUA6e1rA+vPCuxF
dBvA6e4NXaNPAChugI+ahYe3x1LcZVjC5v/w9pWY1qBv5EGQz/gp8z6m/dMgzJBI
M56chz/I6Ti1gqhqOw4QB64824hNPX/fSRYB/Vc+ksan2SsFNK37GZi9ZMAx+9q+
sN7lakRor6Lri3stdrQ36KCKa3uEeLKNqsFCgQKqPY0qHB/G7ZfoZ6hD59yac5uo
CmDhso+qep4PDr96W86Sz38M65PdlUPiDDFSI1NVznMqtqwj5RBTHXvkI2U3N138
Lb5rqon8ADOtOnzz9u9hv5Iu1uvEMwC50CZrp4do4RMB30mXt5BvHPw7KuT4IWNx
I5yi4YSN8ar1sl6+WnjTmaD0TZx+lMcsXiQleHKkP3eJwFxQ4+BBsWqC6Sdg412B
d68OOr692OH2Wn1WITP3XZaHayVXqVbS6VPB9flyJBj/Sp3M0AJv4GIcwXVDenRW
Lx74GokZHyr9GgJFy3t/ABGgtqArbGdBBwQq77Fd161jb4cxKdqVlZl7g6kWcBrI
KaQWUehImmDEdIde4+3lpRhQYUUJklRzVKoX9vnr3hzxx42mrGrLizo14ujPHlcG
7kuY2YW77oYZ0FnFc77SrNEZOIGMhtfr5Ez/mPveTqaCiHkRDJr+cogiDAeXjcTI
ul/5GWc5dY3405jd95bmo2cEyfaZK4BqCz0U2Iekoa7fgYdsvZ7rtFjgERMFbp6s
4MiSLucfXBJxJJH0q7Ct3cJW3p48j2FOfJOJHsyWm43o9dHdj7izqrG58uBromMO
/aTWi6vrG9EacM5g3gwKSnqGddY6n0+gU70rhyC/3leU1/8SLSDVk+uJAr1iGxOe
Y+DCOcWqQBFzPpScZDxH2EWQraItPQwUd4qPW3ncE7pzp6a2K5Ls71XlxOrsLcGJ
7HWxiMcttivU/V5EE9UUK3v0i7KOTNITWY/T4NPE3HmpOfUh1ga2FGMx5vBNvahM
EO94JuFuYujbrRLTu3iUzYCgO8Wo1dZ5vuDqV00PsXvdMjQ6aCcX2rpqW/hAlY/C
u3brUEhxb2hYi0X35geNIE+DiuSFx5ocHBAJgXF8kEUkWbFvZBeTyyGAfWNt0M1M
k85HpuO8n57Ns7uuJ3PcmoDXIRPYdNnY9nh/PLCa/1c9WnDXZk48qK+1djGnBCNh
4DV2+nrgETFfIF/DgqRCS/EqCzukgMwa8ulzqBvH2LQslOCxS3fdnYnMT5fUwFIc
Eyq94Dsc5gLpemYfoDkBf7vCbVuysGmiIcPXJkY0UGuXPP00VVphkmWd0oGH3xOW
mVQsGimbLLpPnZMoSWPulPBCpSIOKv3IoubiikZi7GZqyS1nzjZc1JW5ToR7fX8U
Xk/Bu8mc0zDXZPOzksppV6W3z1J703qBUapu6Pw24q9IljAATXm78njNeaYfTGwi
nkVhl3zkJHtpX+aAhcAbD8hbWkEYX6Gzy2I/tjBDnzlCvVemMJSEtQP83Xo+t2+G
La5c/CbGt7mdh1oNfrfG9DMQxaVJyGB5ESDxia049Lc9+cmO+6zS9lbL2/cv/R+m
v8b8TiFUgVl71ag5p+iffkbOyWRMkCxHv1L6E/r4lfuVya3KyjFy4wRk6PLod+mR
L6OjOWVPPnJpG6ymvRaW3yoqKoVUwrTiLHLjn1OGfDhT6rZ5THQgRWIaWdW+Jzt9
Qn+RAfXgSKMbdRg4yZbaEOLwbD65SWcGGMyYdfaHRqvvvhi++suIJO0sBeOyWr2b
T5nQRIvKOGpZvC/z245Q5yYTG9IM7xV48eL+rf4s+DlLATtln2q6zRAFbrhq2J22
ZAJ7T6cvMuMXdkhdm6qSAU66Do+ak5OMwD/HKNib7OerRT+jdmaUVPLPBqyjLBfY
m0piaqRAfMoPi8K4FWvSBJjWogUYtoC62Bqbb0lHQJvBuJJMCVQNYzdGdufkLea5
qLaq7mf6cKe2a2dSjgdaD3lKLs17tXn9Xc2KsZBFNtzkY85Iqs7PmOqJbAqAxWXU
dPuTICirZZAoX87e1nQVuVPALRLLa0Xetu0xyHMtoXXU7VEr/duJ7l61MwFrWcTx
daUXp+0kF/zYt2+QQ1fTo9Swy2GrTKP4+IjNOCaLPhCBSGw0f06LrxVjwfJjYpLb
UN7QwM898Tow44X/EoqrBARRX1jSmmrFMkkbWGvjaG5IKk0aOoRd9JvCz1/o1P0G
djwuGJphqRUz0wgtxSQEHrV452CeRqhIamJ7aGdw+xGpQGixhkt4Uioa2oHNzZZg
Tk1ziP9Cxum1JqT08vzumYUg3Pe1R2T/PrZksfC0jp2/H5l4WgAQsGthZ/jQzCj1
43z3jZnYuEF0z3HKweeJIPifepeI6WLa4pwM6xTq7r4HM8O/LUh2tybYPOic+94c
ktBlSMAYBtpzEP43dTLdaEGGWQnsBBw5lVKTFVJUJSyrdTaqB0LAPDqo2fhv7IbQ
KRDdurSVBG4WCtgPePXzYvgKA21xeMRel2NqoP0ygY3TcV+ZTxgPm4hvOpsF5ypQ
CGGTMDUxUZ0dZOEDG3LVZOc3LMpYU28UWifuOTOW71oJiBhPbjXlTqte/knqjQWD
1jh8z3GqUs9CbBPqlNwIFM1SIMGbNP/zsNhXQPkGJNyXFFxIjBZiDU4PqMWpAI2W
af5iEMEDgp2zhakcCX520TRaNc6u1WKiZdaWjQDI24Ef7I/src5FrrRSBbNps9hv
pI12VSjkZNSEtdw6GJjc86pKBvILAAic0YUM3r4YoLNA2deYUIkrrJ1T+7GBTMv1
GHfMOptlCXPentESVJpXdFdlL2mgeEad23HWyWhGlMQyi0CO7oAJQTCBI/Flph5A
FsPv/vOCXJTCskI3yxR7En05x8XHArVKmsZK1LohVBM9G+AmA4BJxgVtaF+mpgaj
ef5Vca5QBi6xX/2SJqEkpBU3qFLL2VfIwa4JYc0N6PKITx2YzSNmwJYNZhF/FHO5
iknhkWcY0rs7ncXJveguxZi6lbnE8Z5ViOEmF1oq4+5GW/bsag6vIeDDozbNVL8C
8izq7mWwHBDPFVCWn5wV8DSdOcTuNtHIZYC05KsSwhScjPW8Uo4OdPZNkqT23nYH
IJVjbaEZlRhszSNSIQOR+v9/dWtqRCsyPa6ZnBJYqvnDS/l1Mhk+l0CEwh7CzAdg
rbm/K2EgkI2PCKNAAOF/gI/Yyumo0YIbSlJ3aHnqau+zHQAOIcFEZAaRaQWLi7q4
oQ/YoUZZf5tpz/e1ULPp8a6E7aY8Fk4ujb8C2rr/RfBwP7vjxsyLTHym/S50+hVx
BdOta3CfDzThLWIXjZbh8oLvljCRHWoVA5WUWvZDtww57YptVC5NzV87/vnc1qsS
ZIeaUrgiD96JFUuZlojVHYsNpOMG7rsRiLOuSL7bqjHvnkea3Xk0zw2RNJ+xGFjW
1Q9Qx2H83ePj6l01x1IF83om1V/jwTQY3EWpU6pO6xwV6FiWIta5hPsh5SS6teYZ
zAq1b0a/Ql00hGIUBVNasDQ1EJFOyIs7n+3GERVV86tL8aw65VRZQ42DpJB2c2Wg
SCBL/MjFnIcsXilkLQE/Cw2L31WmG1+nAI+uWItrT3jOwcuH2meaSM/bisX31NeR
QAvDu+zYZP05jOV28HsXxhPKV4ZOT8Qz6CQ83m10lYyZqIc9YWQ5yVqWBH9Q9Ljh
BRS7LG1H/19xyrz8JmQYhClqSIOjbvv4IainfZo1XR4THnBoz2hahy1U1uuna0//
XfEtNevsZoeVoSJuqedax26rXN9sCB+ygn432s0s6UoFy/s4JuSsilsnZ7iethM1
LeHebvGP+wP8Hx61qkTi3eKM27LV4eyppGsz+GT8c1CS8NMZqrmLk3Yx7LhTN8Cv
15O0Is9v3gUUecTdUSo+qDSVnfk4xbNDiyD+KwsMV4ge6ELm7ZYPu+oeDhqdEZ7W
30TTPcNyc23fDAxUb87EcqJwOWTumjAJ+SpjsFkOIcCrIv7r0c50yahzIhrfnGdr
TnGN7UljEn/SpTBt7WtAVde8lqHugUnYCiOVOTDSWl8Kb8uKGMC+BUSNXZm1KdBw
JDGg6BP4Uovth0YtDX1Rui+BI8FhYp6o+4Bp9K1/iBaDzFLMxxlXLgxV2jTa2fts
Ty1AYUDmVxVRsALMc/4kJE/u1wzd/t/B54w2EtMWtlBqhzncFXzCtIZoYqHn3NaB
vvQLkGqtZ8OjMbUjYo85+poaILXpX3Zn1bW3f4jAfdHHjlSkBKB+jGJW8XSkZ6uF
/5ESGAufbkOHsf07PmUlZ2UDlt6Vep2lHHssYroWCMJ47+FGSAx2tk3lg0GDfaWB
wZP5BFbnchYqtTXBeYAg0gEXaeqVq3QoSz3xI79TEdzTTe2fi0lZA/Wh8eu/Py3w
SFQvb3hBzyOW9vrtVYACk4xZBgO0VpO27Ge0e2fXqVRWHoZuO4w34DFE1A3bpxA/
upokXSPgv8AABUrwijrpMnBR0JFYmiEA4KNwuG+L8JwPmKPBBUgNQhPadOfpMr37
tX6ff467u7CSNcAuBww4cleYT0f0g8EG5cekcCgMW0MRAIwkWyCkfa72RrXFdwte
6uuvEplD9F2jHmMVP84PrJLL6DfH2pmzfScMo3WwPtvTSC+RfGiFbb4fk0uxM/rC
fLEsZEfvmOSxtXpyTB/7tWW23/8S+jSTlR5F3Kj5a7y9hVeOH/YuAOP+7KtpZ+6q
dfERbC9CWQ8+3lDw5XaNzFe5n1HtrPXDgc2ormN8wqcAPzEF79RFp1dLGr0Ks2B/
UzkFiOQ/rcTeg3XIV47hPXfv53qQxw6TuUcvXmA5ydFDC4+D9AOfVTCyW3l/vFES
0FG7hYbPJpc+dfJGi/2KemOj1Q0I/EsJz2yH64uKsD5deRsVgx2731ZuBAC+PK/q
mxr0oO9pIPN+frKe6mBmrXi60N93Kyp6I0ZRUWEtPcMPTbhRorU6njsGlEGL5gQH
2xlFJ+7J/YBtYfJQcoP9k5E9fr3iOBnWvGr8fuqpkPh3cXDfm29ogHJMCiBklXJo
9bWfaiTRZBAGYvuxuXEIYLOCNQoexh6P6VxdkIYKKbhUQzWT+l8jXAiw2XQEXOC6
2ej1PNqB4nK27buxD72Tn8JmOepNpehqJVIoR1iwRHF5OcmxoBZdvlE/NX/QACEl
Bp6phzyQAqlP8cnn5VhDjkryUTJv7FqCUKilcagh+SkPwAA7tyE/f4XtcDVW0xxb
gzCbGjY1WCKYrPX8vjf0Wpgb8OsZQuf3HDIZyPv92LKFHyfsPgzVaWXE4MgcIyuq
p8HIt3cE3JfxLFCj13DxwVwFM14cHz1lK04OSrpc/opjMp9BeRqMgMoRyHSa6Ln7
+qHW7PfIbvf0VWXE8KE3INQEYJDjC2TBBMNV84eWIbR6fBknDAsJGOreyr5SyfBw
k66J18nsFxPE5JC7HMqvCAmWl9GHCiMtREGX1wY5GJUf/xj4YyqkOZ9oB/lelu6z
ceYbySHzCUFvr0SDLA0K5NNT/extxJxvUFge/WWckI76+grFi0Bc6r/ok4xCHpk+
hnAgOZe+0CY3kXU9tt4IqvLjz3igf1wPdjBb+O8yb35+4lM0VdQ5DZb1zjkWKG+M
7myzFqtsbWLPM/q00ZuR9/Tv0gY6wHdka3Dz/LJT9CDeoIMwnDw027B2quNj459f
gGwKfZYqs4GdaodJYrLtIyG5vREKEkH74rRvH119LMKBIchH8p3CP9bl/Qp3Na8B
FocW0u99JfeOhU9rbjl+lCcExCpWslWcdDPjVXglhE+1ExfO/O0G3AdrRrXB4Qhl
tC52vcZ4rgBmXKHTO6yl6xCsR4jdb3MBuXL9oOJ7vD15OpJZKX+IrvZY5C/uQV8w
pq1cpgdcIcFHKXit460jQJ5bzJrSf4IBZTTvTeSoSIxiiTFGaz1CRec/TtfnArRe
8Bt+ZfA7ehToq4ajY72x9YN1bDfWnDBru80aVAhm4RTfBm/kFWJLS6OG+U9vuZdR
zMOGutxdZ/1hOtmOrNHaQrSM1wLB/a2o4WRGg+UZejTrnYQq2mKMaEEc41f3nsAd
kPTZOPLqycfkufQDwR0GcNMXwrwRxIBVAUFFzc5vfmz6YDXyP47KBUzy3b57t+FA
mB/SM1x511YNGdgUKngXAwRIFb2iKBhrhzEZy7bhohpg+vAuYAN90AwLxnASX1T4
FqMkjOPy0tdLnmHGlKR4cY7d4hn7XZsBZbz2UZckozbxpRBy4GvVF8SupVDDUj+v
jpJrE3YEMbuYJenzVHRXf+T4y4wjdirVucdkxTLSKA3i6VE7iKSkBRndTkcst2DG
qDhCpMhGVTWw1TlBAgaZqGgRmnlJI/WKZpHCnQliLberCr2zFYjEx4mPZyGy+Axz
3QHdTCuurubegL4eH6OaLvxIzLG/pdsOYNuRixKXcgmnqis3kp3P2v4K3DlVNeIs
g6Pntmi+BwcN0Ion5PGn7WwU9mTd7W3zvQxB54HH3V9e8IBEQOCUkUXjKkvVBrZj
wEVvO5vqStM1UE0YiTHylZyIwEHuvYjGfWdw3MPtlFz9RJqVpDyf/91fOJLjt9FS
LeQEMfEmD2I6quMWHy3JFMN/t+ABFHz9A81+ldYgPXn2ccth15cQVsMoshpsIfzS
GFuxOSN8WaxEWiNls+OKM9/4AO1t8f8PGOffNu5anh0AZi/NtmFJBFT1GbtQVG4E
wxXiJItGrQshDLJquDhA3w7JAoeJfBsyiHpiRuR8HMaAx2ztYq3+AQP/mK9tZyt4
HYE6m/jetgtQrpsdRBH1n/nkfkAvh909NidZYE7QzeM1ZQErOg0W9AhtnycjxFoC
NH9e2EfLnZ9trOYhSs8D7R5ibpH/VV9NINFRxIOx9Gt+JA3aJdABB1sBLTP6qrVV
5Zp2gbX6JjaASMiLDnmULemp5X5pj2qWKRXB3gHFyvMOzAkJbzmG5aLC78shUpMa
qEZsoBUuQDzbvaIGLmfLIsBjnzizechSbxhWztUy9MNo7dmuVX5uquqsWg/9Xs4I
tmcSr0SUPHUEIupINfh9l3ORWwQE1QWSTISdB2nGWZi1VUvIM2P8Tw5+6TzH4gSV
hf3qUQtLAHhV7MHqRANGsOJ6jwetrx3dshBDcwXjPYCvXlc92A0UKqPXJbMQ6WPg
hbCmVZ6NU/mxWJDs1pufsvE8reyM2VpE+6bFw7Ljbffc6vA1HYO8hG7+NmTiliUw
hNFPSqWCFKX8cy2fXTPpLrwA1PWG1OJdooljzx+uNzoPKwSC2sMhRQbJjB94985m
+JHEo80f/qFdiwscc+Y3kldJDB1QPx9V/BU9S653X5ROBQJjbZcjul0r4zQwC4Wa
KBBq8MP1e2vZPOGUsXXjeWku0Puu0FMAM5ltqj5VjbjkBC8onfj+LqLFUUOjGNNt
FjfJKauQVtd1TPnyxkRcTbgkZPRRcHj08Dcisb9jNFatspP7QONHRWrsN+quDRsb
t7lRdhFEtTOyZMWRx0xeIyieYiWUj879xCl/CQ0owIwxtiXitok01PYb6kgcancY
AseObm24UV+fYFdc5sY6VR1NAcxCHSeWdNEM/R7lRyNuWxMguEy+2trRXfgy0Ekk
ovJ+SLU5fQ7f56J0m/Vbu9iO0t8BBI+NHItGElN1okleyNPpzvuNWfAY8ITL+UcZ
TjWesB5fiCPm6xuw1of+PaQwrHT0JIDcZxu4FrYRaeXStbxe/SXq2Oy4z/ypdr0x
puob56VuYu8dkzjAjh3svWLiSozGwIWRAiOmv2qn6zOLewJOUxmcUyKXcoHYaiyr
6p6ZHkMtsraWzjFt0QAS4397iyFXGQuF23H1aWzOAyesUhyBVYw/zTT1eUNBCMoD
PMLylIPREl9FFTMLX0c/xTihsX2Nb+8qyUhWLF9YKocgzfWgBSj/bj4ixHXjq6Bw
Y66HgUg+pWJYtGFDAxE+9ims+4MiwG+dOZUnonrNFN1kch54MUW4XOtakzXPiAx3
61YUHh86olc/B09AXaJe4QkSikJTRZMvvaumjXyAOdX8OoU+8/s/qTbZhFxhKhbE
ktRdHwTJDz70Ihg2QsbBXilwQxUUAkX6IIkMgersittQMsrb/SRlCfXg99u7fVp5
5G5hCxKZnEmqVRUsyYwL7PsQiC69I1/gZLjTT0LKDl1hFeZ3AkQr8eo8LQmEP3R7
7Dbf28skRtJLsIfHOfT77Ze5vv1m9jwEyLT3HKN7cgO3ch4JAbL8HNHKCXlfMInF
tvz9rpPkXr2xGgsUJmqSgeG7QMAQrDbrON59V45ZMMUFFo4mQU6bYnqRDQYQ3Xsy
Oa1TDZLb5CzOXBWrXKFQsFUFKsHvmjw87gX4UBus4IPzcCEBjjzaBZngQAZNQU02
rWAew8e3WHuJJo3Vl8aV0f08h3+Uy7m+XBlfMG9Xy1KXHs//iOPRCta369hKuKNR
lWD4+d1iyGcwDYUOS9Cfi4GAkkrT/JcHx0ckDtee+yM8CIeuJMrXwYuxW2QT5i10
qfjUBSBnyTKw7Li8eC2ESSfbH1dme/p8kFX88ZUqVO803ejbnU9dCaEISDqY7yg3
t2yt8JFBva72voVgbDlE6QZqSSkmj5sBsqLz+MlS6Lqx0ZXaHPCSIWYWOIztnTyj
w6/5CWGYW+Ow4+YcZNwxCQc2xazduCGHKNBcakitol/2sbF99x3QGRrtqGZZnoth
coH0zoye2uS3idUQkDp8SYVyA06CAZv6S3a0wp1fsvrJiE3sRDgS8pnWQXFySKQM
HTdxbR9RZFHpk/7K22I5JxLfLoG/QPEtpOkjxb5nWp9KD3AD8sWXGuPR9uuFkJTJ
WFzWU+YWPTD8D+9vRT2LKmTdDh5T3pK8cM0AIE2hFOs3qSLPqSZz2SgGudY61YGu
4H6W3XLLZRq4NZyZqd3bp1t5ISlIUmB1lv/9ELH6h0SH+2KYvoXHsGBG+GTJi4oi
fmkkjRjKOxmheZcM7+HoQoC/H4TY4pmBTfgrExDUxz8d8PmBc0EX2HOAJmVqEX1y
VDF6jBwADQbRx7zpxi7p2qp/mCXSlMddmdtc9h/5AFjkGkbtPuRgBNN8oSTzxoN9
NfvDhksbhn8FjxQn+PeFVNqjQqvn/VgrruJdVXGL1UNJ57rQIX06P0jgUTIJQWIX
NKhuSAn46aZpmOajCgnHrsO5bAUHvz1WHCSp1uuStSFMA4BorVIfHwp/obwtvyEQ
L17iwEVPwC2WWuM7jkw0T9LLriELtOzT0zpRcqx9NN9ycwBorGfY3Y0O6+Wt2hcf
VA4CoI+LQk85B2HrNv5wjLc/UUzaaQLgkNcaSdeJX15bO3mGgjQUmsxN12VXmMOX
gpdfpfS47FKuA7Sg4Aac23YyZhamvQzyoEQvC3OQ2MeRG+c41Pb3clYDIaxGEd5E
wdJsWq6D/Gdj9e2dLeGeofR1AeJdpXJYf8JZJkjAoy+mifHXKNagCb15HppusOfD
Mp7e8hj4sG8KdpxDF0QPoBArnCVhQrCVxnIUseef4hMQY6HVu6MqKko9QemPOIEe
H5DXypNNJsAoU8dBx3nmy7z6k6B+RysVBGNcINpgjkjXRRs/bkkf6/Qtiniq5ira
6CxqLV9XJSmWThwEUQeFNAbfp9DAiY0CdLW+AFxqQhSpN+KLTdRPN+naKHwlOcf5
VTTcnCHFUyPNiFOqwdUB5u4tENWZwCcBbKe7A3i25ZIdEnhP0diHLfr9mxb5Krg2
A4oCWzLtk8TTIjIrviKW26NgGePWe/GvmsTCLa1ceyagrqSFuq3xznY8VehDYgJS
6lLj4S9LmmeFBZGJkPSfFQYVnAVQpqRYRT4wXRl6TMZ4YPaXnkOFdIU8UvoQr6Cc
PNbty+0kEk7DkGXlYL7CfXLUOWjEn1i3Dk8HZAYauU4ulzLPSE5ZBzKrgg3rWJTj
AbiqjOHe/WC9s36ws8xXwUg5yRPcxV8dcr8EGJgPV9acVr0z5bA36Qt/isCvh56c
9gn3QJcKkpy+dpj++f6TEfGJJMOJWDyshX+3wPW8jqu4swnJKmrFtBmy8OBRLnLC
YE2wdmJbxKmW49BXl5gs7hCZiQcA4vb7zQyHVKtCUgdb+PUSfMFgpY3YVXl1wYSr
ESH7K4dwW9Ircior3YDovvvEuxLbHFqhyL398oO/QH1lI8gMKqzjWv5NAW5RZr+W
MHUflty93F+YmoX5bfpCXon7ZImD6zmJbDkIYS969j7SHT7unb3YiaXGPcO3Ssc8
zDIl/EADhHIepMXa/dHbUj+txw7pi37HiwjsGpABPxin2jlonswv5FKY+uS7r/Ax
/1HVLZHw9w5vqVSP8fA02mTP3loRjrBZVJ0gP6NJYgg9ofBAW7dJM23u4fHIml15
m1F3tJlWB7iOfnVjG7CNlTXg7nVBmnODr4YXoCgMgDgXrBcjKWF7R6yq5ZhPVzjS
uSl8zfnKp61PvkJ2tgaZHY4xHVKrRj5UXsbxpRjCJcPDzBTMxmGTrYQxqofW92nd
MaYTnsyZXkSb/9VsWuAgiGtmvtvEQrLjfZdZJvmjMCRvZ1hAGS/2xFw0X4XWVor/
MOoqVVfVk4F7HB8CzIUtKZGDYm6LToFpvOK6bDn8ZeoQAYIrbn1jhvhezGpym2xh
ce/FYiAQiE9Orag17IjlnPqJLdyUrn0786R3zJ4fkcKcN5tX2ZZbozhSCIYpBKo0
zNmKPXtsyr1AZrJA30eQlCk/c4YY1BrUiVv2PcDr7PQQThnpELiMYfQNM/LiXqyo
bE9IMVAIhZpeqnSjMXcyBbDAbPKr3vuNzTropKVil2akluakdI5pvvRlH+QIFSa3
u38OicaewiWm0PY7FudeW7bDrhAvjBGTZAYPtScxh+56khyZlfAtoP1ZtJ8ZT5wW
UXEkktBcaCJ8RCQz4qcs2kdrj39kBE8obiE+jZA7XYmyYKbZodpdJN8O+dPOoMVx
pE98b+LKvNguBTXFqNaMNbWZXsfkxpZjIq1S2A8Ugmtz2SFbPQbOtwKV7ZlvKJ5/
Q2enmi2+Cjq7Jx5cEHy0fRorIur4VSiQO5yj6Otm76KmkaNQHxRLHAWFIPpAWLf2
EszEjcIC9UImPdMhF3xFGdMzP1gJe2ce8eXwb96HPfjFfT6g5Pe6OIlPkwg3Hx1v
weKEjZmuxQapH1Yf1dhKq4A115gRWg1t3KrI+CJ+SxGRbeXsEnqFYTl8D/8r7tr7
IYBKd6ddaby/snjF8EHlMd+WC/GE/cLcwmZKwU2gL9ZkMTVeprDqhphYEj3KJ1fv
CXQsHw3QbTTV0aPdXzJXnTe5hFsWi+T3xd//OnaLykSDSwhzQ6YRa5g6gCKRHbZW
5n9fycFxsRylCpdYhxTAHH/y9p4tHKN4U8Tzd52/rnxGGKSMrYRxRN9gBFkK+dU1
ov2YbTZbAXBw/oX+Pq7t8UfRgcWK8Yrx9C2cXeXbcn7JUpvEhccTRxWxqBV8ta5G
rpRLQ4cxA4VIxPYXDQTdVucKrAmLcolIFQeprfVKP/mLmUdB3rrMSXt7DRJcbr9w
/L53boLKeyBo0G3TnnOhgPz+fFCeYpO12gh8R1V31rcBN4A7f2O2uxZYnIqtcqqa
UitSk7TEccNa5Ih70kBk0aVk5SNwB2y9F4H6UuApzNUZLOTZtI5QUungoXcF++hT
r137l1P0+RHCFx590ZbqLVYgwGzzpCpkh5YkyWIRqAUen4R7E7/oSOmS11guHjc3
UK1W5Ai+Okvh7E6+aFt10GUR7D4dfe+K3Lh4zm7R99uLP606mGbOgppIbjlx1yUW
bedyTdd89gCkNZ6l5Fdo3WskfDAZAHlnx69NCYDV+Iw12XDTFkTlGijr4Gru8bHd
3pORgXnFmWKwQTrwV6tUxcSjgt3Suqh18aq6dzk/znsAvvGH5qTQaNZ/3mhyMQdA
i9jeqLx5H2rg6Y64d4eqh4gsxBF/CVVYdlnS6g0pDsT6q4rV2Pf9/QL0MY86dmwB
ubDdsUyPhluEnN659zmJfucYTlQxX869Arp6yJCUmdaQCD+Nw+lZEitHdta/H7HQ
TgJnHrBnAbMdrNGa2+CtKvNIG5unGxkoWteVRZ4wJfoxm3gBa5sZ75WvO7LkUF10
V9DGRK3bW8fIdB+aBw0I3Qo/KU/52JqqRNFvaCFmBrYgvnn81M/zy7vXoZY906RT
IrEpTBGCJ7hdgIkUnlZVMima2CzoQqFF/RfA9CVBfjVoQvD16y43NZC+eFsiyvxG
/3cjcwaHz5OrHJq46r1lFzohzgfLrQkVj1u2XmbgBqGJ4t+2Zicqp6jfo9Nltill
bjISxqjmI3sw/HyRPCgXRAVO+xFjobNCnLaGktkhqv8lK68G/6tw8uCL3m98Tixz
qCdOzDOOkp91HovsBH5dclsL2G3vLkonsE7LWxpSpN0K54x/o+fkZOpf/GxdjFnK
q8td7808TEAwlb+sji4JVskDYgpsYAAjwd5CjRkpR0gtiDOvQjAYQawB0aJ95BqO
hfVXLirt83b3ikVcn50Mvi1EVItmqF6k5vodcw9S1jSAAvxkTarEYg/xE3LGTvC9
niLXsRzXX9N3GHbMDpisN+e9AyBRrT0IpgYDAgJuus4GPZD1FyBhryWe51DMeCC0
k5iFFlgFaZpCCBbaaO9q8BIWnkdyHbe7o+D8nxJrhEBtchTfBll2eOHa84eMLTmB
qUw0HQK+tHPxHT4ZtprdlQdu2dhyq8TRt0HEs+7Q/tAjByoMX4u6LoAs8yizlcLV
KkAVoe6vTxcBsNKqG+O1hJLT4qBMKaGfpTdDXjIz6kQxivv0p/ipkjcj4Utq6HM5
ayJaRKfTQxt5a5i3rwYQydrw8G6VoFew4Jog2lmDhTb9xFiaF4XkJsl8Zc4So/b2
E5/xqlBrJ0NMD4/PYhlPx6VzfP8Xt4O4W9Q/PaY/w9RhxBjBpBeKzdqlIGmQVHyJ
ZoBW2e8jNCKEFGlv+vYOZSw2IdUeVD2dhP5o7f6ckcRF9SRxlQ69BP0CNRTja9eZ
6Q8U6DCCWPQeqjwkPrHSjcuUgHBwAOeO9Ee+8OTiTyoJmOWzq5dMUZEjG/kyPgZI
yEK84M62xgc8NhsYQIe8v99oV7n3PfDxG5SITzX/6BIn9DOrC7FX0CilOpQQnfP7
lKQd6r3QfbsjK0r3oOhJ7R/GsnWSfO8aTPQLVRLIw1JK5xBRAk8UDBMZvH5lXij3
IPEE2QQH0NAnUF1f9wKP7Tg7VmURuYfKT4a76TOjbOYtmzrgj9MrJXbbIWRdV6kg
jQL5VZ7OCSIYVyXqULIXEiAoVXql/VPozp4GjzoUOcLrp0FYfgkaJVo7vTLCaFyb
JxhQSP4jHPeOTwa8f2JNu4kIHfGtzehN0F+s2bNdYI4+sCU7jmBHFgQPsSuy2igK
61MOphLr+tHibFP9qFcaNksH3QIjQJRdNktd2F+7p8ZIZ50FErMPpjGT04ioZ+iU
2RhLAtckonpPAETBFywo6jYFQtbMx6F8cO4hVBTVmVZ8ogOF1yUn2JHshNqoz4KG
TOp+qCcrJZKU5+IEMwt/hHQ6ta3xqQlBUbWHUBE/xHptHP1yX4XrB8zeczpYNsou
y10q0joM6pmfDnIZlElrtFAAt1PuHId1fQz+XTY+XBZ9H2qcFn7FlrN9ybb9LSpL
hdig0++YcU62Y7SLM6ab34RTOkD9kAR8PmgDlQVV/9P1F39iYlsRwtTwamIm0aMO
BSjzYfz116gjoIvUPlDmVHsldvsj/Lis2iCzIImIL5Raqdg27QiWKtE4kQ/x2F62
hpkuURPFc1zu4KXpxG6JPFZexRw+FyxT61KElyjbv0my6UimUw3OH0nw3gDFZ5GH
o5vqgzEfomf9IGKCW/sCfHuTvIGiKBSomGCqw3cMBvN1UFQCvCO7m1vkAUzlzvWS
PabiM+/l+cNRZoV5WrDtEH3MKQW6wDwAApDQKH5vNfm8hSa8dWHhiNMlHIFyxhkD
d2dthJlCN78d3LeG+zJFZ5+uxgsOvI8nQx3VV+BslBeu9cd56W5NOmD0rLehucuS
vGsMImTJ5efrbLlj5d63m7sEOy4L4iPW6qpipDRGYV8/6xej8WdycyDOz5ZvciVg
A7K8Aruq52B0RFauhNZmmDCusKcasl2P5OyFsX8n0AKUqhAIC90iFeFHc6CO02jc
WjWoZj7Gd9RryZNylMIiLyD/OihCPAU9veHSXLGmL3Dvrip/VcXVducn0Ac/0s/f
FHfentA7B8UkXahkb6OHkDdv92uaX/Rx/QT+NGRYiPVwjtDZMHucQnzp9AXHRQ9n
81Dl+YzKsVWyY6hFaUaGR6oEpyy8OLh6WQKoy30WIyIMuUBOgwZu+erZJT7+EJEA
MCoSyVUEHqQ6YR/azo6pXGVvhKyOeHJoWNuLBPZk3wgCfnTG5mC6OFsz8IupKyAn
ahXSPXy9i1M1eg3QZeZcwPh8exasLFP84rXuegiRYYQbHA8oPxQzedDD33muuihJ
ocYwSigbOGXlq34cfVfDyXLw+3YsodHIyDgvxPiSPk37IrdKl3HxfVy3CkfZzdNe
ci1+CFyS6WTzhtvExZM1lDnphmNpUfObM/QM4mexKKksnzNkUJ66cBxfWDB4q1EH
bswA0dWHlLvTnx3aNUrincKrOVO/CKPOLpMOySaPvt45ky3CQw/q+b57oo7nPzM4
09NlHYzwNys97ILodxb44JhURjUVP31GcYWmMH7zcwfrpWBRX+xA6Gr+SUQ1K3OE
kSpZ8oS1v1BWqSrwl2IXWO/uOF5dUy2nQYlt1r2GxkZ6SKoQtixc3soNRWtTIUJT
MvZaqN13YM3N8GLu7NajisHgGg7T+G1IF8y//iwpJ2LcSvFtoRl7ygHpw/+ywLYx
iy2m+ebeKqmPtCQ5Z9aecl7vjwa2RRiPDeFt9c89iSMUhb0OnpqaNIcC+28pue5t
DIBEPw4bMFAEGzd0B665J88fcWpe7zqWvFvog900GMmreD5jKaQ5CRfgPZDv+/8D
P8aHRdTMd266ypEshdjt5i0/srrI+VPhSxWH8ckgSvYY3hR6d/vGy+qCr2pZ7Td7
CAQk/m+XFwMXuwAMYZuZX/fo1Ks68p74wN16UR+8REs2A/heVJDXC8cJUQk5/uhw
gr5QiWsmihVKdlUt7a3pnLGzh87mG1w14sfqNM4f86atYagUaAFTqbYQzS8G42sI
HXFjjScWAndc8DEj7hah1NzzS4yLPBD4Ij8y7aRzIdvugWNF+Zi+yOI5n93uuzeY
sP9Q0jw/32gxiKpjEndmu15nxjIqcBD1comHf0hJBbuc2yW/obE1UK2dF4FKgVAm
FaEu4K0o1RnBHe1WhoEUFU3mqFKgDnQze5axc6F1fAenQOImOBIp4atnGffYDsI3
4+Hkb0HNRLgjCWStKyOIl0TzNc9alZ0pv10209Rmpt4yWEubqvv9XJFoeRlH4KMU
vJW1x2lBlLe3ofOKYoJSFyZe+dQkdLFcd9je8sEJsnifxu1gKECesF7K4GDy3v62
NE/GSwXe1mvC0D+pBsXlkGY+GaLlYrVJ06OuA97dUKmyvqiHK9zAqxckn0MteNqY
Sxs0J6pMQUYamotLkhfgf0B6bnRi8YbTMAT1PeD6GTdaRsp7zUQ+KKhhGbXktTuR
ZXV50KnVQU0nh9MYOZruHP8JWkwbFLkfbsRjpMAC9QnGUyOiTGZPHipludskHPET
FOUawTSnsIjhnRuAIBoF6L2Y2cbfepuJ5bmRpvTAezneS3hTEyUhHoGatu2VNNe+
2i8vE3ma76QnOFP3e1ZiLSjDTMgLG22f5Gq7D1JpdW4tPNmwkApYLFW37PYm8Bem
tlGMwNf/oCY+Na3yPvP7/4WVGf4c/+o8ptUJCfyI84PZWr0+pNIyk5Qh3CppEvD3
IqtSBBPYJpCD9LJIJQoboR77Z+rrVy7scpyVECg9nuBnhAj3NfaVh1Q0SviMZ8WT
OU7Ab9q0fnp8pKFj5Ip7nivaPIpqMQJMHQMYrz2eRmsKfedZ1/3eMGq3xPitDk+L
0hY10hDs1s21fUgR6tJmC0Oym+5vksR/uLp2mYXSfHJtlIJPgeob7S/FYsVuW1lI
jLpIIb6KPWCkeATnChgaCzke+ZC1iqD9nvBuogTWw6x41ybbbusOro3JtNjnbMye
I2lVPHcrggdCuByaI1jXZjkY6Teiz0Vrj9psA93eL13twKayhniMV+d8S6unB60E
zwu2mOQiW+hH6FuWSfS5HWShqbEKN6ZuSTOB/rPRbA7QHDoIAJx/9CN6q7+xt0uo
YuTZO1qxGP1QF9CxCYz7cCr5Mwyk1hbH9P5e70mqv0ewxTQ/GZzJwnOrrGQZgTn1
NKGoXhJE3QzdNHkBHRBnd/0XEikJI4JKYlNxcUrGqqGAgdOx8e6Jqrl7sndFb2k4
7ZxYgqYgY8jLQcuHdikkegaeahK+raJEww16w7WekUQQUatdAwf/2xAKeKxUQN9f
i3lSw+G5Vf7S0WcU5zH5zSIOnC6iMAJzgtSn4h1UfQ1wqaC0FUykSF90yppB5ShK
0Kqu7xj6JdbILWrwx+EuN2nUNadiou7LUCLXQkswxSCuhBuf+or7f196uFIYyZho
x9Y/jRsTvr0/kKrZaJuE3iOYW7pUANsjK5wkGJ1k1DSBBhZ4FuqzJCZ1ikXPYP4j
yK0rocYLR2TMS3wEd+eLB3ivEhFSIPnYEtf4bohd/Gf7aWoIE+Yi7GXuG6Wo7OsT
mHYAGQEgRJ75l2t/kuULtr7OV/+RIcw08Z1jxUBDbqbB/3Eat/fGeak1cgf4+Qnv
WAs3U8uY07QPz36/0gDwKfDozSITinQPpG9t+eUClJZ5gJWUIZ6NIrTfhGyZAfbN
VtB4mA5ZT45DSI5FjL/ylhehKtrgHJPtxF0GJRGgVfu56KcqqSV+Prme2PG3GBlG
SC+Hk3fs09eRCRkNYOO1JuKLwH2rLIHDJHpM5XIe8JfDYR90H9TyIBS/X0RDs4+X
w0rVM4lBwBNox2zj9L5+0yCzW2O60ETQt7HL1XejKJRSw7crV6qdSzhuUz6aWhmW
GlU4IQTbwS4mJNtIq+JjnAW9alXXcl2YxhXqCnKPn0XPLcH3w2FTgoT6xO62S37X
6Ihy0ocJ+yaY7HK5kz1UMhUTMCtLIxp/kZq20kfESN0q6xIZprN+4cgP9FL+SnJ5
jZEBpd8wViGBByM7sYbWQSkTC8XwINMZVtc2zcwPf8FLubyn0/npdkQc8M2RgjsA
VjtgbgjPOI0TcAhno7U1BGepYDgMsbRYf1oqPGIfIePHLZPsZ+ce6c4NOFc7WDlw
aD4IQ/wCcCQKJMARAu09m7hJ4dXcyiR8l6npbLVkbgrWJIUayWDbTJALviUhRRvp
63bYfDr+mHp5+dK6UDkiDN9HA+nC/QFkCjnREgw8SDH/ZffUas4fY3wkJYw2hOxY
TmgkXwXbv1WpJDI3Fj4smj5j6y+YrSQwLWLgN6tMw0bQx8ztexhWOtrHk5B+O6aO
PmZAbZikTKoT54RD/R9tKdT7cIbbUjrxlFKoJHgaiQhaUzBownFpRRtQuRAF2phZ
NOHYAKRlrr26Xrg5qSc19XzZv9y+gtXg65T+AM8JJxaPFWEB30TOxFkGbMup+CL1
Sllv9UKx0gk5arjFN6v16vOD+0CsYqfo5UARzFdBdEmMY74Uhwbn/EEmmP4DB56m
AjACD85b0GykOixiu1UQS3d0g37HvB+/MjCrkOnBV0scx3V4HAztFxQkH0IcyCQH
dpjll8leEeKEn3/QYkSZty91rnyoYMrjkUGnmpw4xEpZ3wnQjyHDm33FKQQzaq6a
GsZ4UjlXTrmBQdqZhTMRMZ+C0epn45xm9St1k1wF4ROCgV4bXxgTki4it7OnttsG
qwbpB+M2exhEoWjWoA+dSN3s5P3YP5DgjaerWtIEBZlafT+G5vxeA6Bx9DMU8ESX
yfk8HiYkxJd4u246TFFAGvTo+pQ0Z8IdU1S9Tt3O+s7ly6kaXyoKICSMxZR2AB0X
U8CSdJ9RmLF9QRz67E35g9G8HJZM3jvRU8RjSHqxcaNGPL+qZ7Gh5WKfjUOmPlH9
MYXKWwAABDCq2Gbgw0R/mgYpb7E6DTLg08hCs39Yziyvdo/mVh9YyAUD6Fogu9ZP
7ey2cTTBZc6tjWGWGNPTgwZYXX0dR2pBaJ8s7xRitqEnckvcP/YraVLjMkEcrZao
cr1qx3wymBnKP0J6jl0Aaag0dMPs8Lvhg3g3iz03V9+Xu6Y2d5B0jJ/uXJhEZLTh
3XL9g56dpqerX3zTq3oSoYcL5n1miQLEFpb/UcbaXsSK84FOoX0nJ92TghqGWSvV
Z+KItxHFcKAxGON6jGQRVq77fR7/GlcBRIQfMURrkQWZejPPq/tRvYYju2SWBn0m
JDBgpyLi4dxKdj6o6A9+7cGIcppI3i7qgKcKcE8I122M7SLwKjy08CGCqZbkPNZd
h33iWbZZazRT1QaPDRc4ZcFBgFYCKfFou0vPzCSKw59mwODl/Bh5SZ052I8s5zmx
vFzKS92RM3xzGL84XVf8GyvTfelvSEuEBqI/7j0ljvKy3M9D1N4BfEht8hphTIRi
NtWAI0im/pTVUT7u7kQAruCkjqYgZQ8pE+ZiyB29lYCv/aL/QXMQWDGY9fQQg1XA
qIhy/8YsA548ihABeorJiL9TY8z4MbFEUu18AH+uwwGGw+JT0jFDFNWotGTH85Qf
1/03kS7rmaIuel7vL5IldSReOsa3QXj5yZQs67so3anCYe8MMAtx+9Qlskyck7Ei
LQooJ2aPnx7W959BHDUBF/jkNDQV3rLTuoS/UO34zko7ZVlPmy5PEjbxPNnsNSie
9FWa/jP18HD+TdMFF2sfJyTdry9O/oEfhiN1kNNn9YKkUj8ZndwIeeZ24eyJbTGQ
8CjlSKQsx9JdZ7cHo8bBiIFCIItEqxB+ozxdx1zfZGxj+vIz3bjUp+ZrV8WoS4vt
y02MeSsD822y8pGsQKAeiwoytFyELZGTycN1UuXO1mFl3gfvovqjXeUqy7hMvUbV
+d0YNTb5aMAlhIo2pbITc0GqvYhWnEMNEKq+5T10O2D8mJxlAMHweTE7Av8ViQE0
M+jpn9vLAA4vqmyQc8doW3bhgYS9e8RdNL5Nq01p2QXufd8EQfjbEhbHEeHV2p2Y
s02peebCLH2bvOwse0iquY8kVgOo8wwTu9im3ptawkw/snObHzjTDDx+QrwPV+6g
CfYNJyTsmq/riJinSbPAs6z/neUkCtAoxtku4bYzXJKpRAedbzkSd19onst2IsKr
tulJyEdGWAJaQ+fEO+//Owmy/kVJD/qUr76n+t2J7fMXkf3UovA+DVWtiDhMInNE
lOeNnNBxMcbzucFQYovw9XlvzhhWoyLP1k8I6IFIJ5g0iXaMVaf7cDf1gP13+nxV
tizlM6tu7b4UbjoX3naiowBbk3JfxxtnEVnuyLoOqH3DNH89JoQSORvuFJrHwBW4
ydKQ136Mivyn4kkwRpHB7dOxlQV8XqTB7+a3DBHr94mozcC5JU4LfALVPumqnwea
y+NjUaa7gAestabXLCjt2aJ15pQLfKSmNvaql0c/jwzwT51FulcndoUHXL7916yA
BhaWVFzRfHyaysW8f22V+Vfi0EVqwEQCOLVt3xelCAq78qEQFa1ZFsdAgTLw1vfg
8ol7wG3FZ3i3v8XKqZAy8pdutAz/nLWPHRnn64FgcAQdMNQVFcgfqoUTi+0oV7AL
J3rAO9qAKt35yQE1cDUrjq2fupM6WmDR3PCgrUOoedGI7b984Y2VA7pcevdzbok0
BMLUfXDv+u4y1pgs/F6At/VtR+zr2qEv1KKc9Bm/FcTkwQySkILTuO7jWuQsGye6
885ZLue97ocmVKUUtb9DkkU3MHW5OIXv1Zx9z4fCzgN7hGkKeKMPowUYPdQU+VDM
cWdOa9xWPRzn52hfAejv3xpEdY6xfZ61U/Fp4TNrjxFGHsmOxnGeQT8OpaNE7X9Z
x2ZOOzDeUbE9LVXK4VyjEKjn2HR//IzFYp5pvpLtQDbyOOC5/Zbcj19n1AXpMKmd
7GCe8GcYuYayLZvzpVX/tpu2feNsIRob0aVFpqP0xiqpRqpAbCs7SH+On12HSohk
xZHTxHKqM0sN7GdfeZAqvv0Wb7+K5TBtBjT+tssEnxCB8qv/iHo+6COF/56QxcWH
WrWDh1pDIGyNY8pgDnflZK3MoNOXjLqrUEjqk0loexLGVugBmyEK60iZMAQXToLp
b/T3RHKXfWjqPvgP/WiIyGwyYpms/66uQqKBQ9P2r2tYElyfhJbjyldx/ad4AhoT
ZZXiotdjM0OBRo5BVUeHEFQ6TTFW1N6aWPRNhRdBnUTdFas6+in8VMYjP51wsUkn
mijEnA8chW8C/cAuNNRu/cJ7Ym5H5meyOXFZwmuB2Nd5+lv6WnMIVbgpqHMH0Ynm
JxdCNN+n5azuZXdL55lDBL8ncrGTn+kWdRpaxdmYRBg0hvhgKzTvyY2pLY6Z3Ksg
R3/Qxq08X//AsGJaIw364V2PmSaZsfhOiN1lqlE+kXcol7hJTIN8B1Xok7RqA7IB
dzrviALKeyNQstqCdkrSaoqBlSPnsGcyWjApF6wjoj4p6c3KViJjSE01PkHLogJu
2Cgwn/+U0/dSUY+rewzfSddFMuFtHcD5BBAsIP8G5YvvXYjR0vU4V0I0bFKSN1KT
t1vwtQchvT2sPZ+t2+xhevbsytPliB/86k4xQdWxen1y7gaWc02LGHXHmUxVuNa9
oeTyi18n4bfn/4cKuLnUwAe0oI1pBLsgEiRrW+tNxpXy6Zq3LOZfYhQKM3XmC/BB
QxURZ/7FpSnhz8KIXo/AXTppWQO1is2MD0zYJ+MDsmnx/814+fJgFu9Yv9hTrl6n
x89Al/G717faayLNhCa1wUS2NBSNPNQPPKuxcLYDEISE/yVk64UgnR9NPOwkbtSu
BgkQpvE36x4W25m5HSezxfJF89TsNDj6p0WZ3atrLu3Qzyf3tw9cz+n5Xw6TISi+
VmKJdLhrwVnSNFNnlsZUfPi1DFAUyma48s9q1i1XJZQzhGVe59hXFz5VimT0pmJ+
2vhMN67Cx90g6gF7dIQ+bXi9eSb7dnN22D26WCaxBeNiNYSiV2DMrV1l15F0me5c
C9cJME1VXzNagftsIrpfcn0Rc5DhxgYJxVUIP+yC0h9loH143XiN3hGj+q9Hauyt
NpHcEn1NUHkA1CEITvRHMgsx/XsUuQyAuniuoAwyWG4XMNP4YJhUUtjaDDx5f1l7
QD0vi4hdAnOZ1Jp/f3dkvx8b2QgXxtIjlpxJEHdqmMNOewUI3U5EiDjLMxR6jBSR
9OW6lKLlNnUiOWCi1vJU/OVOHTKOiKHVbp026tRNPzm/GeWfBZaNuHJkcvanH+A0
MLbX8st7qFTeGSstUnFsZ43lWRsCFunY3ZW735IbnqtufDopAUHqmjBMSGyb/mHP
/y7SS80w8zF0+VF4vGd9bP28qSeA3SDJgLaNxpOCbdKrhXzpJQZdIvhHsXJpQ9nE
KsdfJIjw58AA+FX3ty50rG+85a30tKCEOiwzeRx4LlFT2kBdO6t2hPXqjuJqaqYo
/9CgEsg6q6aAZkURfqgIJMxzGfi9PQx87ZRH+EqH7G2ruzBBQivQOPu4KJ6eewUU
2wTN4qzxChUtnsDeJxu8jMaVgJafgdudx92Hn2n+r0C+1BqASk863Czz/jOn46b0
Fd7cBs5JS+fRpzxmKYlMZrekAa9qLnkhGbj24h1EmnGBkGMvxD/DRauIvRqFKiyV
vvJKyt0ME8RkM9HtRNmSEL8uKCgiudw60YhI5jqZkeRYQeOg7GC7HGgy0CXrup18
Y+iMbHLCMifqsH5Elj4OnmUlx1Oxlk2lcuUxIVOuqPlyj43KYfujYH+NPhJDoQbe
gY7/1DeGgatbgmQmASqyIV7OIQXjkmaJRPLzeGjsHFNVQOkIdpVWpqvIPzCA1Sep
UwuJbQQM3Z4ERQcg8WCI0DiJMxIPJA1tK7TaM6US/gAjTWYdcnneNiGef8v2qWtV
MIckVpBOCl/xilzgT9/52QtCw7MS/TTGNnbi8sFOHmM6obaeEwNhBOYr6yVBtrUA
XEPm85B8Zs3Uf06tvXD0LKwUGM7w/f2dvr7eZLgfedsedY2zAqX3JQKdlNOblgf8
OynAiIv0M7Evgr9yxj8uLH3eQqTdW9CgYJcE9j0BM1dvbt1E4n+bWqQY5XvB7vxI
Cu8P5bgfikDH5+5aoZuCkt4sU5qLmJkd3AXZRY2gmyaxwCO5WTwPjBoVrMtc08XI
E1P4h1VrHmz3CLxfyGio7tGU7MNVMKdS64JWguVcwuXkNSfofNZYEKuD+J67/jLO
IU6GeDSmKCDCysgtskJNfHL84JAV5gkcxPd/y8hA2UasNeES+ihw/ZXCs9pMghw8
eTZxeXlA3wXUPnn4l885yaBK9pytORAsAyOE3+bMCGRckluAcgfrIEvoAMWT6/iq
4yQugT1FCDClRFB7WtMDFy1GQPrL6xai8hJHdRIdACmZhj0WI//LRDj0yThV+bs4
PyYXp6qz+7V/+eEj4aEPru85xzNo5AtuoRvIbtKBfTY73KJgaOxEVhqYO7fimXw1
lSuiLooIpz1wa66E0W6mjgKj7OUbddMpk8H/BK3RlfTy66AyPl02CGnAxRK6V2Ix
Wy2/m0r3IiYBRSIcZ2Cib6pv+1xaldeoC32GNFriet6qXABPVk0S9d+haxszNx2h
ZXNAozwklqbllPuK52ziLN+Oy8BeXM4aD8yGy4nkwEA9n/FAvxPJ6/139Sbir/Wu
GiYiDkxl/cNjIOtGZ7Qc0Oy5L2Qozt3z+OZNhGw1pWwkfHQv3O9ykd2KzBL1+NFi
l5rr2/0bI9I0W8Wu9q0dXEmMUfwk6fw9PHozVnGW2uOF6n4PZaHG8oijbnybF+qi
hiu2k1dppXcxmdS7VSyYL4Zj4XGBGfJ/rp77AzugsHm38y8RCrYwdKXtdkxah+Lw
GIbuCM49frSQu8x2BxdT+3OBt9R5o/NAgaWe/YvYDhGUoz3atlBvBAPxCjYvJJQS
5FXz6chOMWfV8XboElAj8ww+m79RBEkloYTW+hgPL0H5E0VY+EFJzKen5iFO33gY
d3blqAv7UUJGGQe3kwTdA9o2QhJAXoF1eF13fVvHs0vm3vhG1wGiEhf8SWqTXtUu
lPYV+XgnqImbLhk9tjItn26yBl0IdSkn8b2vTWojACBS8RDMxJaW7g2qwM1MfDtC
8jDral+RGyiMYvhL/t5zuH8TcsV4KA/98kW8EpEL+yoX8J6vl9434NQQcAF3liLw
Ug7X/sYcmF1VraEaJ2GgF2tM+tqSDmVW25hdiBcDdJ4WaEriKwwU/6vc00iKzyRt
u13nT2i2qT7l2qh/GuXslQ0/r61SB1t06JCiRaH1SNcubdSYZnesTfCTvLWLVBW2
INg/6Gg64+Ll8Y8wddIUik88OUnXuBLvFe/cfXUAxPcuAXREBH3F0v2fg+Km+9UU
+uqnw8UJrwLzrs+ERnZLCh09LeNmHrmesV4+fguwIbz5eW8biJORbEXl5mwb/z1S
pPIKhljVwiVn17muVd6OTxqvjM1VavQ3bkXd3C3g8kilwfRBy4ARKLdnUfkm1Kf3
Q0njcqpYuC66PWyhcBZExXMBedgtzHCpvt3KzDduAFkXmVphe2SO+K63eAk1JhAu
ESLJpFvuJu0pJhM2vZiluNY1RCtv/R8ctqjxHdSp6iGrXNXl2pM8zS/M9l4GJT0+
by995U7+OkoVS0rvFbjSq8dWZOzOoiQQZ5/dul9iiBDvgAeRbjcyuqT2BC8L0z8O
TkyrRwmMxfbfF76uLMO847c1ucrdD3HAPjvdyTIiyq+jB3C//y7d9RLE3fl7ebNq
8TlsxFZwoZyGIJuYCKEs4xvoiwTkRon04+6rJbo6jX/8eNJkGkUiaFDmHQq8tTwd
EnH6tn6O5vuP7sgPUv/qhKbk5tWNlhqFNyik+xOeS6F7vy34nfZsYzSnyLy6mZxB
AaLBrmjU9z4/7A/zYzypTcurz1mw1M77Y3g9+MqTn6lGmf+UyY5EjMVkCLSku9ri
r7wPpcq4cbYiEN9yD4HRaei5/fmVKlUW7Cr0sWIaoeMsE7Wx0PR+0RkPOF0iSWEi
T2kyj45AN56n0VCN5L+T1UeTOEvctp1COyYEP7rzHAxlLjZf0Gfnal/94lpBHSHp
wYBMN/6S/tZbSOoSS0cIBvQ7/ppDNj6YlVl7jZT41sxjvmua/D3R06eGmHrm/MlC
8Ouwy8UMPpuRjDjjNEJvzU55uIjcp9SMn5qY1meEI3dGodbnjKxNxoErptdOrv49
5zxSirnaFIjZqsimg3x5k36rtjOtc0hl0OgXcoNr1HtFZUEG5gIcVUplPyqBzWfX
nwX04PWyz6SkP7HfRIgrKVCaddvWa+at/mTeW1EUlouLh4kWrxrvTzDwDKVC6xFM
cMExX2/NqLZsJopjpSTfDo8ALioe3/SbBf+H/PQcjMXkjX76Zq2HmRt3aFbYvJi8
P6avwRm+g011kxb1SqmNgNew2eXiJMej6HW+3m9GIV/rsMdONeViSdrY7fhDIw2m
yRZIZYJU6jPabRnqitXf/410Nvyy3g2pCZaTLIr0juALbHHbkhc6bSzlIxe5tS2D
Y/nMLqFkhklg5YhIXtlr9sKYJrqgtR0YMwajVhsswKCyFIoDbsIlAbqpx6u3EcJ8
hBEein9f/3NH2OhoeS5+PPai4cGD6lu5A46kAYvqkzPR/R/TIzrMNjoUZkPlhN/0
zPwuWh1CIyHSuy1a8Wtsgmtp/iZ/QrS9hVaNu5QPFKoTTWPSKG5iqkQvcFnsVE9y
YiSs2t9Ek3aBsCGKP62zlmVRPcrvoFK6e/l8gxP8SyHL40K+EBAzSmyd0xg79FK5
CUYAZI6aGO3RGReXgHknQ/au9d4Dew9ZXLpTKaVf5fF0cocnGw6aiVs9C+MxlLDB
rSailn7zw288uXh1aYHYySsylNXVs7m0N/EO85sicbRyKvcUWvZ/4uh4EA/kcl6z
27A2B+1T+Fj4p6zTUM6zOV2/O2dJ0V8qtfwCFdcKouezO7QM9xJE3eDuF+xQsLiR
hcb3ETE8UHXCiXmxu+hs/iwwi26JfabtfsvF7gsWvwQa6vTo/C/EmcWByKYs4UlN
BYBXZZ3aQVFW8w2cP4jhAh+APvz42vPO18p7/sfgq5/m/iRjC62yr22MZ8BWHFk4
8duFphwna69vm3KA4xhkvYfOCBpDf8zrCHXsKjY+pVDi1+R3TG+0rOeto3r7SVJa
IS972zPKEI/CW6nHodTZDp8S1M1nxA6RvZNCBqXPL1p/k5V3uklYmciaI6q2obmB
cpw0hPLUzo8ZkZhEXnZo4IepWP3/U8+nKcUNHiyQLPeUk2D/+oKsBvJgfdLbhovi
6EAI/Nz1ga+1btzPfzOxEP7lkhcSbhhBDQXlLhMZLJMIltNYMjoWVMh70N7rCdR0
WAhsNa0VOiLC/QZJ2AOWuazDAvgRMhK80Q2xgXwh1zzx/58hgLgMhppc5nFHfvr6
7i4sCtdc5FpjpaH97icudQSITF6gjUTULKvOKzjcnCZHOuxFP3hpZbTvYCXonoXZ
VXJwoxDudS4aZQvTjfrs7EtkgNtpsOUuyvhEzaaP3oAsPsd1tq09RofFmhsEw+IU
ywrrjPKD7UvkMnCRyBJowkwtQdnuX7SRyYgijbziqnA2cvlo2TYwBtWksibIVTiG
b13n37YqYwAOHoablecnlWLC2NZ1pdP24YDz6hW6sht41VG/kb0xW9qTmSs1eJBN
oEUOvpfiZdDBjZErnIz0Dq06AEOk+/JZ+6py3Lq2dnetwlVmQVu7IN7edHfGmGxD
7tj3UwGJZHSdGl0gZchV/nrfXeFYZ+k8JjMUG5Fz5XjbaG1prQ5H3uR4HGPeGQw/
cRDDqErof9ZsL4BNI78yIj+y4Y4/7bUxcpI9Ilo17GN6Y973uQaGCFf/Qg6YVHz4
yODG3kDZBP8qqnaSsbBLQBaqYNQVXcLM9ajMqtgumJ0htozCU+5MlHD4g3guWjmF
77+KNTTX9+CAjIQk5XAm4ZdXG5Zmn38lXBg+D98o87o0IupC4h1A4w1TMrCGlOzw
6QOmhNaC9mDAhKiXAXsgmJ6f9NmNPWJ0DDkfYO5l+rM07m+QDKU990r9GGR/wbOo
N6zD8YrIlj1ZNcyQ9JdvgE4+kpbQ7IcpgVQBJmHmY4i2TVRCxuuMrnHiyfR4kZuN
k3eHLUbvaGtSq3lb978BHbAm0fkKUJ9Abb/J1RZ+hzaNB+Dum/Ry8QgJrdWOgiaL
Djl4JInMIkKjpQEy5XR6LCEgkJCi+X/4oVEZRkvRr7EyIbKCPGJmyNppbhF2LDPf
xXgvVcqGv2DB8iUO3cDbXOO3QSbBNcTwvzMPAD/LcyyipBkhnAOADM/O9Kgxtp0z
2anSf4fZ3Fujha0BkEIK+/4rD6bnWDK3KbKiwC7ydtC8prOJXZht/7JEl+3DOtS0
c+niHlvTbkHiQnEEYA4doHgS3m1YSi4jM4TUyS9jCaZMvovvg+kfANbGYPGfOY5T
5YcfCUpZC3wD7h88SXSIWyi0q7UBvNSgOmsx7AfihH4QPO3+scWkw+UgDbJLj6vd
3N/huY7/AOFQ7MMuwT3P1doDLFt1RExdLeTqkjvLtdsqNZOFAbPgWvm1acIRu98k
Cuo6HKphIRCHwo58xwNlFT2uoAaYeTP+AVrE46dsaZ9aj+of3hd5myvtYefXSXqL
sCZ/NvLvJut7EScRNqFi7O16N9lUVaoFpk+LY+G1H8+/PhscMdQMoAP2HnfNhssX
LzPy22li2fda2hCvKvH+NyYnzNnFGgGnF4eanjWeZ8/Lg9SChgLh5kbtwEhqy5QB
aPDE/wCWCEOX4CcdzkImFPk7ARtJxfBsdiRmOWd4W+vGMqJOvZf9W3E+LHeh9Dpz
hNg6u45Bs8lfciy5CYNaPsZp0iBVXJ+c4DGgYjW/aRe9zdKMd3Y839lIgp4lg8dR
xPV4u/Pwm6k675VUMYYdpeUxCKvBYnDp0pi86uNiIxM2rATVwXp+bG9mNgQrvcc0
mHUnnIYGksLvJbcbDPLmYI6Z5ZfVD8aKDEFU/lCnvNCAEC6BGsVw+VYyZwyDXEkS
0rI2tbUrxSK8GuBaFbXYT1mHrPrKRmdFKEiVBqRf9R6zZLVgk5dmrLbTNh5OA1B+
MdYOe4IDY+/V+4gQt8KU02+67BjDPlnVPRcKREOUyk1OoCKlFAsQ6U4FfkeMoqKk
XA5yuenQe0DD8eQy646NEQFGOT9JTb1XyQK1o331ZxD+z6uYvtcJFiKza57b6dUf
oYBZ37NpQCXfzTSjOXKamqBWbsd5Y0Ti8cBSocMBishs+QHp/XzOQBVfi1UKLjOG
g27eeRLH4qTdqpt+outEjF/X6+E02jYykkxn1YoTuhZ1GIA2DeaCVttaTFnuBs4y
mbVz1th04Wg9qC266x+sTjwc2TtOuJLFphmzqECp8SV4m+l69xtRi7avFV4+H9OI
N4wy0EuIOGPOUTz6oVFbmEpsVfiNuIOYsZ8OOqroV4Adt25IOVlSySmSE0+hxvmI
unNU6RjFFp9tZMkOGv0vgVdsAnrWGqtYJlgGeLEcIyy0qBpdCb43OaulVZzbsfmp
aYh+CHVjWRh/t6ZLj946SkZYx5shRkV3ME6zNwHgqyC5LaZIK5WmrJlccWByZ/7K
NUDJTpHgwL7s7huseQsdcMMYawQn3EPWBZ6fzyDOMs1YBguPFuBsZe6Zu9JLIbxV
MjAVqETUwpxAd3QBoglSCyklNxOpjh3atxUxZ3vQJLlDroMuTbAsgfvk0n6bL8LQ
SymhU43sXnQ6ydR9m56GpapfigxDfNxx6+09CakDCXbh440enJZnM5VQTX1sZSYF
/hGeP+tRBf0dv83egP1kmEek++VDsRJNyQvwdkQK9hrIkSb2NMvIMriJ196JAi/l
7O+eoKK0hfUhK66Ry83wvvQ+6JAYsLn2hANlXp+IsOR3frSIbX2qhzL8hu/g1O6M
2Qf5VW0i7wcdsKV410XN13qC/QPk2qWgafK13NzsBBF4RxEeuG47ICPMK8sji3eS
+Kutt9b/fwjMzVROarzQKfQQbBtgiukS8/KG3a1+ypMi+kn2x1nY7lorhJcUqec4
/x7Dx697KGmX5c79NlP6UHYd4yXj2arqEAv6oXGtj8w3FFIFJYPWaValCQ1ZdxWs
XFPezNSNS8nnVWK//CZJsJi00bSlsXxoGUHdkJXbnxjrbeXc4RpMMTdXIdy4drS0
+nzLIwHuH2/pdpgO/DRf/nUe+etYVGuDsVyBsNvzfQf3r+D+RRYf4RmHCZt5YABy
FXtSgv1k0CsRTBnkJw30Q5rY9R5nODVCr2SKRA5IG5Ymh9CWWIGdmF6Am4BUCjAC
wkgggk/LtuJ0q9qfBM90qm0oRHRe2kkVUQ35TGjRTJvPc/huKYv3xD+Fb9DvULlC
/JWPlm3CsXrYNBeRl5PxJE+nLegRyLOXY8wYhmJES1fYMV6iYgg/fxa+xoHTKIfy
bcKPLjAlc/G5/OXvqzZRBdjeyljl2pMLI928Nw06IDz6atyUZiB9NZM65RcKziJp
v0EO9Ua0OcSIKa4UsH26mGUU6MtuaRU5L8+K1wrF9dm0LnXDzA77sIIW4GpWq8ey
5zFADyDL6rPJpoZfyZ3DkMcBmXu06eheUG+FPTE62zxcvN8fMmycBtKt7hAOcP1M
/D4HMnz2Y1ph/AgObrt+hIOOhvdPrqIGVfwmXOOEPld6MpO1Q+hXDHpsmGhgvtI3
T2hSFpH7pQss2IQ6qKtGLuRlMIa5stFHd0UFLnbAp6KwBOeD7TlaeAgRWr4y231y
KGc+JGQOS0qdS6yANBUfIO6Zibgs3Ebw2340u5U8bwdP2JDKlXJSYxNyHf4DmBK2
p3zTT6tSS7ioPljj/9uke53u+WeqktpM+jEep2mUzFGkFZyCswpKle2SADReyyL7
5UHRykAy02MatUFk9rwtGzc1pnyk1suWNVB4g4V2U7OSB8/2UEWdEGTMoXIwmEqP
KeKqxcFX6sIH/zcgtaILm8IMi7MXCV46+ecJYNKUkCIUjlLV9nn59lq8zGQVVros
KxM1Jy8qp3EewmwM8gPiwDYb9zYhJqvmhnzIW5HjVTKE59kFsNM6NwVjXHhDEuOw
8z7fCp+vQr6RtikDpJEEN7qe6v4WB8+Gk9b/bgqvElwvcszEIzxebMER9AwN25ro
P31WyMOhCcMgTndV0R48Lmzeb1ATECcKMQEtbPt9cb37GS49nn+r2cdWU6W+z2rD
x+mHs/p90xCDbNRfPmRmDGo99ziyzoCD+bT4iVkhBSrPymhJW1aSMHAO42v11OyS
9qcoG6miDyEOMhqkUpa3++hoxKzYr4W+wV+c98HDLRg/qPLUqBl7MoZry4Yl3RQa
UFlHFvhf8Vaf+vksZphBLr+JXa6h5sdkDhrUvtwJ+NgY40NJe8jKJQQ7zFIU+1Fh
bVr+yq9NM0Ht+AB7i47G74T0vhq/KaOXzqi3FGkUvWQJ9HmSxwkMmOWmD92AFT2e
0qOhUUHhhGon/b696WV/IwrmNWHcSUy0/BinYEnURfTlaewdqYoXa03mkvIr/QTd
ww2b2sDVz6ue5BCYycvUVvdcMOeX3gW6gqBG4aT/QGaC5n/hZoYb4GmtxGGiiGgE
xnmJVi57cq86PLuBsqs3KP/U8RZnpRpyeFcqQmMs3ZwDq+M6wvZTK3BmdNXB6htL
vMD+xtfWYK5CnPV6BFy7F/JLif4EhEXMzQDdX5Y8SV0dpBAyhvfWHqqg4IKMpKgW
YyK9f9sG+q0hgqyw6q9ukQ+mPTI6wWlNUDcYHk7FA+LF9BaWaSZoZIsO2SxrGu/G
1I3a+za+1kxiObal4EYeWxIgGQOI/SuBITz2xqaZRRwhTep5OdlRbF6pqf3hWqy9
N+15Z8WA29nEcVyLnIuNSMea0/F3rGoIxtXRBbUDg75dedcau3oKlU5AlXHO5B+a
/oCqWu/BFXgHg+feNfBdufRn6SlVhr3T1oElC71ys7il7taAaNbt4/v/ATUM85Rq
H/m/X/sczzsf4TisAYEm60C5OUX7jk5XAX0aAvqqeMpGBX+grkOQIj0MvHreICsF
LLhOdahpNaYFWX+aSvp9D6V6cI4C3E0oJVNOl/jKL0gyaXZrRzGggguKkxhz1ohr
GiWgL9uNLreLworgPdIO2KN5ojTDGqn9YDBHpC1IDXD3KzhO73Q9mGZbAyQzVXBl
jWqS53ODNkJ2XT/6TubhbcCQh8q1KJjl4iLRpW3C68s/0zFUKPVVmLS8jUjDhCIa
cXg7gOw7YFUFLLBmUhdw6n8o1R1hlCowKyvYOd+KvBMhhepSairmik7sTl5gBclV
8As2/HV8aa5N0S34isTGCS0zJzIP4j7Zp2uSC4vjNi32CyQqaSGrk43ce4Jjxj9M
etSgMjzwn4rmscXDMswKgzndCZu5l8nno7qlVzT4hgGVZYREGk4H9pCQnE8oaA6S
6wlED5RV7rK6SjD7BaKrW8Y1iZ0cld+4DwK3S7aP24JSMpW9F7EgxJ0tGve3TMtG
NRT6zZ9yq5ttbsDb8P+aY2XSN0hZ6nRMkQ6zhegjO4zy2DDIR/l486Dvi6MDHURI
trZLoEjp31aFEX2FgVzmV8TnfrW4LvzJ6JeMJaQvPCx89KIXJkgL+asvE9Xb4Msj
KEDAFz1AYgP31cWJC2n86PH1cjixU8HVI9dfrU/nGKp26CAHe1bY8AyRD9FvYj93
RCijYlr2s5c5Jc/Qen9F1Y3Jv3wJjZ9oMfw4e6WxkCsTM0fO76jI/VmcDSW7y2nC
OGOSCLIfyJl2T3+zHtIn2KpYR1Er8Rb5AWYLuVdyA0g1FwerqxVkwo+NhA0syx1j
1UjEKUe4k5F+xh+EX4g1zKJ6DcG/r5BCgqrsw5NqsWZTKTkwm6WEjNE3YZ3zh/uV
YwXJcI0A+c/3KGKPiTZY3Kwyh3IbdVGvytK3A5RuILxnHR3YROwVHMTbfcbALmZS
kJ6PIlRDncBEtuD7Ws3A6oiUOuIUqX412sMEufYzhDi/RpBxzpvPPxbnO59/rXx8
TUKjFi27qSi8BIX86PdSIHe+h0E5/w9yQUk+91TinyTlo+D66SAjN2th/NjO0Hdk
cs87sOT7TSTaOxyiL2D2cEegm3tLc8S6MAFPNp8WO0+GA96mlBb8waDcX95A65TI
e3HfTXnDTZGh1l7N5FVruWhrwLI8IoIDhYjzZeADhL+tjItaAvMl3inb+SuDmiC7
lm9siqfP7kaNaD5+qgNLug9K37MU+QPpWUnDbM6usd9aqqxsHBgMBiCbSOg0dPHl
OfvxHgAq1nb2+6NkzCiuimeB0oxpBYB57rW6Z6rnbKjtQ026rZpN8bAZZ/+pWode
MvRDm1wH+ymsoB5DqFXnrVAEgSUHP8RrZ/rzeerxV+giEooAGBdVENd03aktQ6lL
wd82Vj7Owfcnvh/48/gCk9qT4rQYfYortqVLL1fMJbaLkOwK9TkNVrbWWWdUI4tz
mi01/2/j/Nv+k8GMSXDu5rluD/5cWNMqOqUYHMEx1WiqCgVtlqrKHV3aMjYiNsGG
VzCLxEkP5zNk9YWeUucH3ysUNgq30cLs2mZoKD5SygeaCUbWFy1aGPFzNHYcOvfq
F6lLWYUZ51Jb+4RiTrpboIHteXOHsGzY/A8LvbSdOP0KdhlKLz9GOTFBa/Ot0GAw
8AByFcZ7tJjiBlAIU+CZtlPWw03veqsOXEzIZQCxY57cX35rlz7rDDK6mu9EEDKb
1zOCvcJqnJxkDGRiiOpstTCL++XnXXwWk4DrtQrDpKHrEjC2dxhgf18z1F8+g4f2
tH/pWLM3aHyO1y7uECHlFk38ndFy1Db0d66dUrWADMMGnRGHMSXrO51hv4Of7eMV
m/WjZNM+UV8fLTX8myUtLqwJ40Ne4tnAd1m41bcs78vFpwn+1KSa7oHnCG59vzEH
DM5CmLJI8+oRJFIpjQ7CZC3XefR11vZMqeBAIXgMOGmQwIp42fJcQflLABKZfRcY
R9mnujKkvBPRT/yOZUc0H+LJVPK5GpYnzlph5/BS8SBhDqeHeXsDmZKoJlVDbA15
sQ8T4500M7iEnuO4a/0idjhUx+8XqrClVdO0/5ZeMMddoGD73GTKSgz+uhcViSnn
5qbQOu1HV5P0nshNTJqfhgXZ38ekV0XnV8gWoPmMMVvIanVK3Ta+QZcp0ZcA5q0w
gZgEeDs51GKfLA8uEemu4G4X/DtN9GfuDk2XhTrE2PBiF9nc0gooC3S5xo0AeSDb
jkEbfG80TppViXWmWjrwCjjzLQ2z2dzHpe6dMsUeXQTaxY6t4Y5a71HzZxVbLVg2
BCf6z6Ng/gejWoBq3XLt/9tnv7UbuX+ZRDM4cE+mNQlFtr/B0hDfLXsLB8bXhKvJ
9pCRpXApqzXG7hxKzvM6faMTXYRgltDS9azfci8htPAsXrp1DoV3Z1Htk1g8SYq3
RXBSGy4k2bhRWnkW62mDgZooNrzPYCWEMJImCplInQT6ExsnuIwcc25DiAPbl24O
mKJyINPG/Nj2EUIKhZrxlJjI8myMXDVULJn8qCERWT+WqnLFx/KqbLbyJGdme9q5
gCIJH7UwF4GIRiWuSLNr109bo9BKj7zUal967mz8iLNwPBhRu/6f+oss43q4h4sd
4t+BVFn+g5kyxIGLoIbZ9QVZgGdFeU4J6hMYBSxklhzd6Dpaiz4FBgg6E7NMqcDP
JEIqd3VkMl+CH/XuNOz2vPEbdzrPWmZa3yXdMFdV86MtVi7DD/eZeQ0+lORIsUbb
HBKjw5AKVSvZJft7R+4jvgNEIHcrAJ+sN99uBiRb0dVL0h5TfQAdliqm+of7txKQ
5KpqhVJANlDp8P0uDIysA8YcD0B+2Rt4KrB9jC0RZvlBsK0tmmtOVJyopbs1Lsj+
bC8tBgakzGO7unZq6GshKiwrIJki5Uu/L2Mf+hDYfeGov9xbl3DctqkbTo7ES0k1
MA6gUz/YsD35lDg3b1TtAWLVyN/td4dU1lUMiVQULuJn7focthdC02eon5eU06yT
cCuZPWsE16i98UfBkvDVryztrkVQQoHs92jqx61kL/JUSH2DtdZCBPp2Z5Qpn+bn
Mmt5IDEnjoctH46oBznZAscAZY670Y3GD74ml6Ajcc0pSoQwstBiPTRz3OOZqCV1
SmT1UE7jniNe4Ogrp+aDXH6Ap2aPfQYU12pjRMaWWYiZR0f901d2zlgomhN5U5pt
XZEuinMU/V4VxEvj/JG2+6H0xqN7m4XiSpECeAvhgHdd0kSoV45a+lU+ypMNH3Gv
kgunAM61hxeDEjFbcPbOy94cL/isd1jJr1xx6D/TxS2AzaionUkWXfEtr6iF/VDw
8dXQ3uwD7y6lQXsjqF55r8daF7jSvsJz95YKeTQAsb/EB47dHy2OGinT52VFdt/V
DhVHqZuGK5CmGrIUqpR8gjWZXwN4xalz5k7bGHaIUtwcKb8QWVefW9skQ/QR6nw9
qOFFeF2XAYj2rFkSJLR6klXU5yuSevmKfaNAHF+uFDPKFc/iho/eZFLZyDYLdx6a
R2atXzZ/KU32u4Rdg7uS+0eMubcRF3K8WqM5hB4IVS3nPOHHX25CPELE12rcPqZY
m+lgpW04puWz0ZIfYNq1fOou0mZKtLM0mzcv+IrBwrBSL7/7lZKEBei2hSXgNxRw
TxLgEwOfI7O8Mc3wQV6vNdckx8Iuz669hTovSj2CartVMBmhqRTMEhVdKKoIX8Zu
NYSbpCv6nyEgT1mn7pDgYgOGEQ62t6edFv5lhXaL5OzPVPMe1YZu4o5DrR/wvk3G
q6DmRQOhuNzciv08ryrwbGdPu0wvRYdJIq+aNVUnTehqgEe7aiNwHQaa9bMwZeji
+AlfV5LTddQPRWEqMcjRA3iXHAG/fcrvNz6sL4V2ay4FuRNGZRh+hji17Sd2I56f
7Y5nZ0FF3B4lQFrM9UL1IQcMNxYHqaKzDEpyZXcOZZydilXYvSn7LTBsHl+REOaz
6Vf7QmxmehBeLoAW9iYDJ21li4DceLISi1p2B5ximQ7IQTd02++s9Wr+H9G2qHE8
6AoD/KCIpOnadGyF7YRr+fBCw9+4rUca6H38jq6QEDvgOi2y9f8c6ArOsib9e+fp
BPrJh3mvcB6VGB7oI+aHBRiij/JwNyr4NWur2KSJf+qvfflHII+Wf+SyYeOWLXjt
6bHatHwXAmjt2xebge81+PD43OI5ZUZsqqwTtA1w1oYjUIKPEpSOi39KvqJSExSM
+6F3FtnAb+jvjBN2xqvqKgEmpGrCS2ifRYON+YbJB1zlUneYOfREbz66LpPb+0dM
cadsRLoASqgkN8MJmAht8+f+yMXBPAHRGnW4GlgvRaWhvc9UNUmozUcpoCc4gOMV
WvlIZdNfpG3jywNQg0c5W4kTI1GUZK4gd1QQYSsYlwqMhCKIEqRKVN5+W9tQ2WsT
D/imhfndPCImNZt2/96PhwY4/dxHZo6yV4JK1HOREfXZpvYVzUXbRjajjmuJjjgs
jJNGbi/AdR1OWd840Pgcn0DyUL0z2sYp4OIkEyqEH7gczp+E1Lw3FwtxbD8RshmI
aBw9l6TTPDB1HY3sssja0ZKPq4zca3KMFIH95XeRvPdzIgfa7OiLSTGOmPnxqf+1
Kt9d/B6hLYoyy/M8/bnkAmeNH91Ftd0OgTnFloDG+Ht/eVxp5NlWfIXybAwDKRNQ
g8O0v2J3XPvsNxE95/NhCGqXDMleFcykV+1ASgy3LK5quJuq2FK/23avUyM3ca6a
z8X3+knK+fvzuU1ulyVrK2ss6Cc3Qv5mXYGEV0kdZn3YZ/pVVi9xcG+N/hDp5Xr6
6KT/pmGVjLizIRfhmXDFs3pxEggTTkCJ/Bp6Mq/VlqaCdX2mqUvIQDUkzaxX4xaU
Ktsp3sb+Z1ALpl/SuBeaSyeJsOhvt+3/kyUtB4ht/Mlr0Y23fnDCbTPO7zwe1+Cc
moeDpgt4nJJcPiC2TpfR00u0YhAV8clBwJ7FgoLquB4nnE01UwOaoUPpenpzE+n4
upQqjA7V1o+/I/ttschLIjqTpfvz91W7ZlaTUxMKIcgyOI9YA9N0HVa78aJJTbv6
UAVm3PCCkfyapEDmDujYbfdB2OSg9LnSfq1FqwfxCKU8qPAwPBs5dpqjAVicULp+
qVN7BmjPSY60MwsbomRLwI9ijSqRiO09AJtm4GCBnyVnr/j3RNXO8tDCKHJyqJR+
iVYRz1H6QSJt7I/xtXHDyE3gNZlpLV/nqpQhPD8BVJBGvZuCqYoy23exOxanss5C
eaJcWl8abxF113r1KouzD4JmQqPOSz6VM3LxHHHfB+FhMUF48vsrHhH7EX2XXM/A
CooLJvJqQgMCzYqZ+KoB7Hvrk8PuSfZvZfpBFKtfV9E/hj2aEyTe7LqHKDsU3Kn+
CgHTC2AvLwwA5f5HxkmIE5UGoph4XAk5CtTrSvig7Epi1oflSz/OrfQQKhR6esac
sTzxqqG4cntcoX5aGoDgWr8jUDRL3zGPGdylrq/0TpGv33WNJC7qeZ7y99Ps+gg2
A5lPAAyvWFjQI/jgLd0rnfMS8xDHmuk+ggsn5+ccN1QSOcrGnvQjIW0pctQC+eYu
tW7FkyekuEXBCSUDdV85jcwOlq4nlQCXqUrEnrIW5Ptg4WrsBftK9vJBAfhbjXWq
cheChLYhUS/27m+hjHbtRV4xmNagG8jyxVGzZYUlusmFCLz6V07JUktQFQhk4kUS
LL+07m3owOAD3wO8x7UELO/Tq4GuK/fc8XzBrGpSHLeTJRTzxo1Mv48qmS7gDJIq
GFROC0Kobbzo9Alh5KfNHZi/8WCN2zKmt3ZKmLXdhwxRuNS+a2u/MnUwyB9hQmWJ
dHr/hnNn2TypjTw0N6aJ+DWpAB7aPyHvmDRe3DZfWocMtB8M5KFBr1zYSkDsGNuP
/NLqh36OmfsXO6BrB+fF1Kz1onFqCAccwlK4bnSbYSwqg2K6MhuXvd5D7B58+e1X
QU8wHmcLRJzTG+gtqFl2c9bP30EABSqdoq4oOD4IyO5GmEdkMvAjZqN6mOVY8Sdt
U/AP4Pe9zzFVY7aUNriw3idTCEfjTqubgV1xaKkhUlLTN9aDABzq9Qla42Ddk/UJ
QxbiTMk7owTn5JUVOrBgcOUcNjb37tmGITxnu6ZjMacb0jR7mEVYjhnvulFwYB+o
KeKGGegUxVhdd8ca7Tdze4B9ZFcFOPqkbc8+KPKs6TBZsMbyrhy9+Q4tzq5TLkzx
oigJofhF01H9z74kkXh1cVvLqSu8H2Q/6na+zqAa3CJ1PlEg7GEjwijgdIl8JNWS
xADHVkr6JFRM26BYNzjh39LY2foanMnmWB8h2YwIAXWdhv7jAVSneWy+5Iw8WAxJ
ZtY7BcUH62p/X22A4eOUigtjaCXE7LOY3NRwH5QQll7YQeM+QUSmV9TMsViMtHDZ
LoHUXLc4Fd3BQEzDcmLfO8FGZYUhuBB9ZVWTkm9WhJsvsB+tcdS5mE66GZ04wSoG
GD1JV8mDp7AfVfCg24YMnjnlw1C236FuP4Xu78zef6GZJjSgs2on6AE23r+tXb1F
+1a8XkF6iOLlm3j+YhkEZBd6LZudTI/QJTkknl0lOIFJTF3wikG22FVLeiFp4kZE
ZFKQb+RXS6+8UXVC+kIrDw13kjtCn5Z4Dorbd56QNRm6gt4AoXRAycxgC+zpds+x
KOzU1e3cdWX7HUdI/f82F2KMrWjurpOMudkLe3hkVRIhsHJJOPPAVDVDzOoJXHGX
fC4H5xoh1KPRsx6MBkNQ2iE42GdNhldOJxLgTpn51XiEkDSQuqWdIs87LieZLyF7
fAZvmvLk+jJlGgK1+9NnzbD/4Qeclvhuokz1BlfsW96qdVZxDkpQ3P0+VgoW3Y+Y
N5Ku5gvkETUA7Mf2KFomOj7RC4adlytS0q9TfvvPyZm0yKIdtn8cohAk1GHiMmOE
cuvPqu9mJV/BxoouaRgiJc60WBdSfvcO17H7v2rncEv5Z2405JJBFaZq91w6peKu
l3WFOcW7Omvc90mnaDxq7dA7l3yTfFpi+sZeyuZrLMtOYNGb2R/BPoxldNejcnJr
1NapFRnDY9AQdD9ud7ThJ1ROEgQdCQUh6ac6YeDGn+PRKgFv/Ja/WG5NZ4YAewef
xBQ6FsZwmmO/GH5H/UCxijlh6ubHBcHe7rekjx2ScPqrAkGZXUE1Z3XVLaQoMVH0
6mcjQjjzarofBinRGGb/RcQv5fc2NZOrJAXEIMquz/6Mtl/NV9YgscDj2ag7pIKv
xl5fRYSCtP8K/h13jwCzRQqb+dHkMlkzHgnum0tmeHTWKh/VKFbhhO8H5pyIWKGe
PURQYSlm/+D225fClFIfZUVxl6zehLUH7COLzzDK3ZyWId+0gTwMUrGOTgsSrCdV
X5NcojDo/pIRI3DxY7cySugWazGeD+z5N+PriJzGzUHno50hjMgRHQIglzI7YEub
z9tMFoRtxxnmrDZGEWDvkSrr/tkvhg9DjCKK2Zk6Ab2aLUT/Oh9DxGXg6vmHKvn2
IwtmXGWzupTg+HSnPWMM0Omi8zwKCDrh6T3BYmL1UsDMsSbMDYej0UBeR6Dh0o2M
glwXAiY7zCbJjF83zJPNL2RBNo++EW1nc8b2FJVzh0e48blCSrP0syYJsRJ7dtEu
3ejJpJMoVAXx8njG3P0DBZBaRAgFN13qYKW4MIjAeglPEDutBS3v88X1Gi/zzlkc
Zhw6ivOZA4Y3kVhl92zPCSpN0d32i6W3kLu3hXNe6u/rpPiFHdO/mWLSFzVPPfYe
03Alma44NG1ppMvZryJ7NXDvxWLbcXT5vOQVGso1KBXR3BHQOng9iw3A6C5x6nAh
xSl+RciWk2GvJg0FQLEsJdYHeVfS+hZCYvIdszKEf74lCJEvVF4gqaVS4SfV/6rb
xSZyOJCdeNPRV59TOx39v6j8aTLKUlFN16FqiQh1nYdMcATe7zFDM+yb+QydyiuQ
j8jWWi0qhA2yW6Ilgbzfl8Cb11QAHDznjDFTm35aOibQ4W09BvamyRdBOPXPI7/2
M/l8LDLvn8xm6SeQja7DtIeQ3Hxd0o54iIUopgLcIiSJQtWLNZE/nLzBwfwizEcn
c3rxEEML6jhw882/tkFqu/cfNaXSJbTGbpAfNFEUZY6dSw8D9bupVeFZJgbuSRxf
9FQRkHtd+4iZi+cc+27wD+itvcjxUHitwDeD4zhgwFeCd3asC7TdcV2uAnfCCJuG
xwGAsVfhtK3y82vb/+A3mgt9sBYJraf4xOqTC3f5aVfFz4F6cuBVRGlN8LH1U6uY
OksBmFMdfA/4IMOucxHeAY/D7vl2gpzO1NZSfKL6RRb1UVLoiUpY/LrzH1lKj4Yt
9Of9IST/aRQEKJmEzqDnDZp3qmJh5bwZr+2R9Eq8AC2y0SqgUBPdDARWWRP87fWS
1+iFxym/tCxoKQPgZrzEev1TBAi/X3qNuv/mYVyA5by18UKsFfxnFWS0KtElxCMP
YZRBha9/+1SNW7vZEOkDrOpbze2hF+j+sd/Q6UXcY1gbmRBgV/Zz4aXyIRGAWdIy
18Z0S4JnY1EHFytzAXgmeHkD20PgCl+sLUVuDHOipLpoyzznY2FPKkli2OzMWCGz
LFhY8BhZFBpqboXPa8ByUyHIsCeWwxTap8RDoN2LiVvTEbwvw9dhqj0+a3VzH34Q
mj6+kqD4Iw6Ecuvbf3CQE998XoTQP2U0y+PcIghHVxHGpN11GAEC1Fg6/LdQcgHA
3zyHBDdObeLraxor+/o5y9omGPDHwjoERl7i1mXBirXGUKQrZ40cBZvJBfNEFbFa
m7PsbvYA2hCweMiCoxkF2Cf0yDbErcad15eFRunFDvrjq/LKCL6yRP79LRU/nJeN
AMMRrrTPPFUuS4rFkYcOrKZojMfaxr5fme7rp9LFmJEq0Nqpu0Zp3WAC7/DhrJ5L
h4ppoZBIXynyOEylMD5QOoleg8bCENGl8nSL5TuSRiMxEfCJTwHY816ylfAU2fPb
UR9NNQ8+XnOFbogrH6a+LjTSdwOYm2qnmQC87yEY00eBshRzgDdSb+Htat2YQFoo
DQwUG2Tablk//nAszue7kPnu8ocLa47wtLAPaGEIKSoawDiWBLBgT1XRtVAt5JXr
FNTfpXKfdTg9cDHhuAWLqyCN+6dFZUN8SlWABEk5muzjY57tQxWiup7BfCygkw5Z
ZmM3xIDotWOUW7/77M85gKuH30cEDBzzBqEhbB9Sw0Ctq7XP3NVCEjrqq3DWTa2c
PWTWGR0+8B5QqLl1aDQqQLgEj4soFs70R2pOpFQOFNfTY+GkuwaccZdIR4mq8cdh
WOZzHMbwH7ItT/ztOF5BAJEzE/pNHh6n+oi55iDTCMr1lm8t1A3HlAj7mu/uDMak
+dUhR/0lt9XYgJeIzHIqfGPE1i+1J3xupzCncSQ0MRZvE6RolBnHlK2jgK80wRjL
8clH85AMgsBiAxgB157DD7+a3Pri1xIlgCtBuIqkmpdH5btBFrPdT4faG8snrNf3
GlLGRc4xdnSYKBytSnPA6g6Rf00n5R/XYgA69gx4DZZ7U+CtZeiuAgUPM98bVCux
uJcDEGP7E4jjRVusZUFWIozaA8xXwFZrJ/mX85SNChP5t0nL8kvrU8ASStmxhBR2
5nm/h6faLdFN2XgNFxaWMjviWHhlaxHFgpMjsby5dIWcLkLnTqvBWA5g3tt7Nnis
b7b4MQNO66dV8DxkPzSG/2c9WJKm1Z0c3P+PXI97Xf39zfWyjjdq61PD0wV3LlxJ
wlYwlM8VaqiEjf1y6PYRTz/SSrC59Ov2bSxKNwxFWC0eESyX9ExP4Q83qI6zhRS6
/s2NriuH+e7C0Hc3Qm1wtCgXTiymre5RiWtPkQks3r6sha5etBRMDyCLTKP0aCnU
YEg1HlriI1eFQlP8/ls/zvFTh5Q+Ynba0GUjAavs30NM0S86paKvcwli9YqGZjeo
DBEQ8dhG2AOqQOQy/I4u88wY4tV8Jw77EXjLwyF6cZkoIzsmS2fffI8nxZa/3rdh
Ml+XDRJ7viE8AE6HrdplblQc2ZeGk3VbuMFutl8DIGzSttG1CFIOV3PehaSbtwxI
Hwsy5OKEnBZvHbFQshcPEPnMxhcTADKjv4vBWgRAFY50/cU8PnS9zQoGW6zyPEa/
vD5V/9XxM0Qp0j5mLhccN9rQCUIhllP8G5HH/Ud9Ph4ZdS+mnm2S3Qbk5yIGURs3
uQ2g3PedxjExkTv4OxVOzytA/Tz9mAwL/duMDyVhRNOTO5ktqQ+HZeF2unYNZaBd
rA9qoIg2xfW0EPT56gxXdgxLEJrcWl3mdFM0JzqWcA6oY37moVf54o5f3QpNUU47
a+imGtwtadubBcplslktDfkUOM7slWh1dbK2fn8NpHa+prhF8W0CKYwwN3IbfZ13
ECZe40MR8Q3Nlfs6+Y0tTK8ZLsCELtJ/fgv5BTt6OpRV7MJSRV+XXuOUr/gQ5Snp
gkMTn1Q8VadCenM1rjLWPKqLvu0kKaixzS6lHGmQL/NUL1zy0/mZiDqklPgOFtPe
jFj2wslSGm/OopghKzH9YFe+yyvNZN4M3re3Hg9F6A/Blw04hVXsORaIKD4sxF58
XcGODY9iXUJZLCnvZzQBdq7BAF4n1PEUYcgfsGgKmoo7QcpdT40ePUBdfETLWIUd
NUDcunvygyEFVibS0YtopQLxruJPl6FYxMidCrZUxaIh0wm883VhoLBEB5DeaeJP
SfA1ZgAnDVhffBNT8zlpigpDNUiHX0avVNTX4P3Y+9ddPdRHCE2DiGpXlJPHYbNz
0RRIQuUi1Qci2pcc2ukG9+4UE90gkh0N+YsHHG24PSrpc2fU9jdWVRlMQGFJsw79
iYS9yBqzSNmX7KHK7sepHOKvQEIgPlOwp/8sVx/P+GK5vyGtsM/K4AsjYgB+yP4t
gHXduI8r+gxqnTNkGQm72qkWi9X5ODCbBK0ByVI0FVS3DbmdOeGrkD3xrVQlLBPl
aOPC7+9NR7xN2hUeOGw7ayRU1OQPo5vsnJydi85NtbXO/NcABmV1mkcVp0u7k6s3
XDDVpdjMBX8352pyf92KqAnfeCNzSk35FtOhrRoUKzvnbdeJII9QmgB4EbO2N20h
Jt7UitP4dffPaBmwLZ70Rhbg1GcOnOtXNhYZ5nvAisxLe9ByQr8Clo0f/n4aptny
RYa49bGs+dlKXxeBnhmlMODzsZziLyX4wEn+zQJyonLkb56gLXV9hojFEatDmXbO
WpOwXMSuI6Ex2dmQA3E/Z74piuT53QCthF1PNJnwrqoavxDLqgQ5WslahGRpDGnW
78TFer860llV0i30qX1nTwkc2NHPlFM6vNfKtThyqdvD/jglRndrfdvTY3fkUG/O
FvXIAUMocRnxjRGYXO6MqsOzGdCAIa357wlutuWFsDCU3IV8sOGMYRQQKjaji/WV
fanT+5UpFIi84l5DRSs4V0qVvoy/MLM3RlucIoJ+qdT5a6tBXVTuvjkLZRn3csIn
j/Bg5aTANu2rwR2zjjWxboAMlXsD7CaPXi/1/K4XT/IW9vQWPK5J2eNWZdfJsQp1
ySp/m5vDnNKHRNtt7hxCLri2UakgzpvtNwBS5AJr9ROqZYjvN4lzyoZSGoFsE+pi
SUtYJRSXFJm9TRvncj4cg8jTCDjFOKfUFvAdSCI6MMjzsBFgdK75lHd7mCh3mrzX
VG7aVFvfCPZiGqPXsDEysxLfTAN4qYz4wXMehKhB8IeWH5Z6ztN2hnofyfHaYVS9
soojLCYjT3kxVux3b0yonI5bEGPj9EDJkTSK3+saD+HCqVOTUzxGIgOEBQwOQwtT
YahyfdyVFRj+AuSOozmIUrD08fCF6QV8TVy9rvt5QZHcd4XSk+TksbhsWSc6zhzN
I2VMfKViYK9zzrCIfblZEC8Z3VCKcK1Y3hx4zE/7EufPdLr09t4/i1Szcd1kpdyd
IPLgLPtEDQA/qUmTM4pwSgt6vMPsu2ZgC3m0FzBqtNiSY+3076Yw4mtgSi8PaRDB
k3dZ7lyNFmh0JGwQNwEkynVhzz4dzVHI5FgDwIC4R0lhhRl0CVuJWvVhqU/HXO6Z
9iRGnRZYec0uM4IQS6Nsc9/58Az/EGR/4VBxitiyPvhzhBA4S0LaKql6LmKMXMEF
LtU05cGmae3nfuRaVTYPetYcnNrKmOROa8DUsFtms6XzAosMJ/Q8WrkkhhpjN2lh
C84UJBjdrDh3jYkINhm+RNnswbwVHrdFeUNx9+0zvhXAp0B/ydvrYpe482DnQXhq
iGwAPrbkpUv29EquSSj2IKCAfxgP7a6yL0XABO2Ct6pXRXD73MfEPVFyEbd2feje
5tShxhG+W0/xSxH2sn4EDWdG8Kj/XYvn6VS2vu72iS518ActuwV9huaZRs2UhsDh
OSZIgEuXBMRaNB4rj3Gqgx7qMJDFI3Rpidc+Fvg4Ol4zLnSoB7LJ+8I7be1hQzIC
uE2RM1PyV8JzyB5mWj4G3nHI9yGpkYd5M/SvpYozKx8ZhGp8gdBxNZc8drKBxssu
HDi8J4rr5GG72ON1VS/tPEODEiQXTq/otyTGRivCBynzERZ+q3QtOqJ+YloteBAD
cAekOrq+FVI9x6C//2Lb+EeOWH7ovi2HdGF1IstC2rJ+L6g9UKKi3AOuDVR+rIlq
KsWDVfdLc2N/9KemwB3JvJckFdi0h5RFGS0kfYeXUTQ9ZvMYhJB7Ibyb50qSj0rp
jogzrrxdm/7wP+HPP75cDTpZvF/0y7XZ3Z19gWddlArgJjWXDE6yWfDGbUTBoA5Z
1CPQLLMTRV7Wf9KEuqurU4WT9kAeficjhK61+sum4kxr5zklrHT/hBhif3GEMDgp
jx3Pau7gBdu3VW4yYcd2jfiGJ+8pdY1FIewlZ6ZmTCHLOIi7zXs2yuKSFeAgtI9l
2UIo8v/AxspWSrVCilVh4giYkLQ39cVnhIGoKulE/N8ffkglxkzqjjkZML3VlUJG
fmkk6gWrYKsVMn6D5xCYVcNepjm9HVX8Kpi28PzPqM45rR1e7hTY7FTO5C6bX44i
Nim5lG67Uy9jgGalDkNJRc/3nYOepV0nF/NzB8RHDvKitX99dVyykq3akmIyCl1Y
PXZNLB6by7d8xDVtIMNRNzSyO7LoeX4QwH/I+DoegHiBRL4x2XSiHaEiVIK7rQh3
NN//oVt/Dgd1xrap8tGhse185LboIjEMKGm00a8VoFRmBzczy+4jMYVChxFu8Hfo
V29NpmphDnNxq9nJ2tTg+7ROinXmkTQTINv6euxUSnrZMxDXNa9LqJKD39fP/2wK
jGMd0hzY586QpazkHSZ8W4tYVAnN0Dm43tdGDQM3p1P1+wzE16OLaZCuVvEhnb8j
r7Tojfgw2mTnNqKvftlqriukfIhetx5ki3lvrsED2y5Zdvm68YTH7jZrzK2fi9vE
tAQa0qID8gMTAJstvmNvRpYztxYbBRdCaI5SCP8x8/lH0xwM+tDErU4QM/+szaDo
XFYMPjWeUAjV3xKlkF2GpRq3SUeOURpF+ekv9Akavut+vOuKtqjnba+hEyuPPF4z
Pzp48s4Pm1kWyB5wCVjmbBDWyZCoV/MdVWXxlpfT7/dJc74iIxm6PaxeSgFxvptd
I5Gq5uyvTKGaVPTZjs4FHp+hRX/7O+cA21ltcuarqHVa5o8U2JnIco5gK5J+wgf2
s22YMXlyYiiAQrQMIRMSq52uZv0nQe8T2Mk+zoYlcKFGW1Y2Ik79ZqxHJZI/ZXg6
kGxicWN6ZSu0Vr8vLOK1K3hO1mxzFMvIrf9wQvrMLpwFQwhCVU7998b08zj7Doro
nFJ2XJqYJ+7XEYL5GohlvmHmAiGYzByyN0yFIS6kukNzZrpepAeKbIlgFWhgktKp
Jw0xy5o7be7aXG4zIsaicDHbPoS2pP9WuuT8CFFvlmvp/yA1KZ+tnCcDucaGX8s/
elQu5TFbjbydzHpnzq8huCg4kEnVkAcWFAgEv1uZFn1jzAttoTQ/HZ7XQQOgdVja
BkIamloxPRziPhfIC+iqzvG63od/fbQGvxzS5DCk6k3GCnk30oaVsEGzT92h5/oA
7yOlpTrYKe/EqhxWmEK5rgXOMWdsABI5URqYZKnOMG+DYj31B+zURsHSymIUG72z
dwJ1iJbI7Lhpq7Cjh53WQROxp2466bGdCukNByXyyK55nt7XlV2ISpP4wC7fCUFF
l5XS8wM+VvXq5dePbccovNPnJJqO/8USlSdLel08L9s9CRiweR79pHHqS0Wsz0hm
yCFxh10T6pMeSXe6uSaiSNHBq3jMmftGfI3hQQN8lxNPAj6Rjs0bH4B+MrjMZvn1
UTFpQj1Igup2npjaIlM9Zy6QP07td2/R0jP0qXYjPjgTilTSDJiCJcFzFWVPIXvv
Kqb9WLcAnQlVgrNv6fRC1nHa2chDIVPabfNi1o+bVdn7Iet4igzXVtw4b0/it3QB
n1p4LhVxIDenTjRp8mmpBXkw5gFh+dOKK+8KkcOhdmo7/Z8CXqIlAH/l/oqsKV9Y
eFNPGqGRneMQRgrYIaIOnnVbA433ue8N+lNJDd8HDzB2kI8hPgFThGWe1Y/EZxvv
/C8DdsATCyW7Z51RFkvXvO3iTdyODN7xCWkWs06ZrsFrGD3jl5EYDV4i85HZ4CS5
YSguBgQYPoTYBti8ziXobOl5R87aFlnv4oOfT4AO/+ifKu9603/Swnq9KWz5xhrs
IHevlo1sZ0YyEWs7D4XjJdTi+mUXYk5Zxlk67pK6FOgJ3QqZoYtKpolpWkP4obmn
ObsTLytl85KkT7a6/18WRcCvWlXWCPTz2SgbtCqZQfWeq5bf/A+ayGNobNACa4xK
WVdUTtNOaF7NLhl9/F+XN4aQnU12UMPHXFa+YG7Fl6zukn7D1NBklIx2jqtVqKIK
F1v0nbSAr1F+vyRH6+Y8XWbvw7D0PhNdVwHOcnNk9eI32Z4DIEVGQQCiGT9f0mXc
NVWho4iAbEXZk/wXkufkDSWwCJgnnqPrbORnf3oHtxX8C0JhT1UWU7QjEw7qL1wN
+JzSwPjnSeYX/QlW0zqA2XZGM3au+2cZU4rUXKvCIuJZqim9QYmHEpoozuvTHXYZ
TO/jUSNcqDaZA9gHRC8133Tc0ML8nYECG0JOA/Ih1o5b+38vLI4RA4SQiolvhh0M
qD1gtKyLtqac1lT3p9TDME5eSRQ5Cv0Ie/HuKlc3Abf1KqhuPwr35n14Kli1OJjl
FX3K0y9TGLwvdvdYUabH4JrA6gxsPr7N/bbG/JKDKWxePuhTq8nIPlnSALLTDVRf
PF35SVOHDUBe+hOIUd5IYQDVUIztTfoSpFQyRjV/lGTREJ6e5AAKFiIgkOtVr5BS
0FbxZjGiqXIp5amotJye2W3bO90B5RUP1lXIs2Y8QFONIecoN8r5Ghyr/0mRwytV
YO14xhjtpTQ5lSNDIAHpcZhsOuR/dZqqL6aGQFUcFmYJvag/Il9kQ0/WxZ1ZngpN
fxnyKBkmoysAyvNXV3DTaRd1lN2+F3MVxstaTLKB5Ux/O4DiZNcdOgwAjoEXU+DZ
vQv2xIcceD7b/loJHbGovELSy/f2F3cxwVGh/f8iZxAcx/z+8cC2uHejIaeXLxZ7
e1pBNsmp/P7z5TP0qi1Xsiy6h35ZPemXvfgKsOi8bhL8DIGZBsd7uGuXXIRKhTu8
bjdfSkMZMdxBj4LYToUuHFWrsCotqaiQfCZiUWdeYS3Ruqu4N+dB6NLKRcsgiaJ1
KJ5DX9NqQz1IQORfDHOfIJxHG/7MgqvAOo1z8bXdRL1EfW1pOKiHaaR/CIsuGgfj
37UYVIi+2wspo0DQJkYmxftfQuy+4Bk7bazYKJ/MZ+7qZW2QNMm3jwKq5JKseryj
ODffslj3XsA+mPCVWPJ+0McIFlU6sBwif435FEP5WPnRl0ag1JFxrZQNUMCLiyFP
OJjC5F7rnrdvgJbWK7v/t3G/feaa0E9LZYBOu55UtSoWZI0rRi+D/dt3H06mjp38
rzu/S8DQ5S4Yiitw0VUWeQj5qQ0HapnMbfgNOm9yR2BWdy8CUWNBGdHCBhf5hW3I
Ohp05lTZmRcAmv75++hBSjs4ctCi0QUy1Lm/TnblR97uIU1iFsUMrTXTVwzOZbPd
8YaqzOTTRRP/eAbemOA3sUwuSS5FMh7JrqCs3qQcqSm/Il6oXS5MgPWMA/s6JghZ
pcr1vYDpG/tt6Ce+akwpkTCUnP0MAE5eEca/tdLBWsA72s0CIdUSSzebbpmiGRlh
YyT+wvFDElY1e+gFR+cvzoujEM/0PnLuQZ0esI/aa0q2nnH4CYqPwgbdTpTXET5N
1CAeeNq7qpxwZTm+H7oddbq9ooqpkVP9wTd4iGTyEL/yddUBgwSZYYV8eP//KPkA
UirG31r4o7wgAiQmZSgjJSm2EjWaS4TQ4s6sNQvUHbjjlYmSfaskjEchaJxAkmSD
q0rEvr77XjrSBpMGqaDySvTdIgOo9Vof+J1QQZERhHOwByZ+DX3RDRozfNuLiWGZ
D1BrZrSAcqp0FVf89WMbNrJduAlqrlFZAp5X3Y/TbGkvh6AI4DKWlITOnLGRI30S
3tWslA4bNmD07vu6Z86YEpuVEC1W7ODtoqE9tdNP+LAwOCNAXj5uNi90CAMFfCos
nq8FjAx3p5Gwq7vbmhC2+dLBll0kH5c3BoD2U5azzEMc8z7cE9lp44Ou+Hcnn7H1
2wQiypvrZWeWQdb2aN6gWlIewj7xrB4ScRFtEdHaG/FQhqbnpbLOlEPYuXWdmy83
xBOv5jU18fzPAOlccSF/GZ3zR9kesyRSDDn5MEOiF9T9hzaALJ2kYmALt7120Txg
yvzMikcbX7jflg8jfMpox5Uro94EGO9Gv6D//XhRPBbFZxaGIBjB4xqFC0Zb840B
TlCieSyxScTk7TbGJqDaNYkO3CKlyKQggH0KIuYI6x/icenG4xgZrnnyUooQL2KG
97REoj0HF5CtSZRyXxm1bKZjrzrSxpWuCjsJmM87RLydKC5HksOKGWYolvD1DiRs
yO8wu2YC0cNFJ2LWKbVtTsF5Vv1GTokfK2vssE8+6PZ7dSLf1hBuURbClriKZQAF
0gxxxTFAGiK8CKoBTArC3brflABWKM0rVXPMcTC8LOcHrxtSY+BKW+WmKr/FTIGX
TsGZ4lIMsVVvB3aRZk2/ymEUMz3zmOxxLidOg7ueSHdhiPJ/LiwHLaT2Qkp4Y4az
CWlI43x78J+DsMTSOoHItyT1a9GV57vVYm42hLUSqeuzYsxDPlonRKBtLhxROVUz
8kNu3EcS6ab0qGX7UfcVMbXELCxpGf7MMcef7qkSsVFICtD+MW8p3QZyWm4yGdFV
MvDTyRzdxukEzXhAMfsr44LHwbASMHZEUSi3U83r2mA8c6ChQX5q57yLylwZOZII
dTsyjNX+0eALg0Q08epUgRryXWz4fJ8qOScGzHDImBtMFI4BFTt2LAaZKmQqf+mV
csx65CydHnp00zSmEwTCy0DGApN4+TSpHjzUbmMfz60HLHvenEJvPl/kG2HAmGSJ
L4o8NOfJN9EKav1op99l49kP0dREyth42YYSDyCLmmDnuJ56F76Nzrf+n4Cg1TjV
F+dkRt+lLoKGNjcjzTlt7bRegI008qCrnaGW4u5alvClop5fU349T+gjb6Ex4YJ/
udi6A+A04kxNhH7O6SbOIyRreDzf1/Me3GP5XqFchzfd3RAGfFvQhurmRdvKJafp
Qez10lguxafpBnzDlKXwNwYiYaKaTzSPh1wLxuYE3sR2/fu1TQL9peZ6NHJVjMZf
JwB1ttIwyLSROZyPV5Y0vY87nFoKWjt7Y+7Li9Qb/122NolQrEUeNWXLeP68s7b7
gYWbo6zKECmyPsAFnFawcapn4q8LdX3rrMyTQ+e41/9Mi7GL9tVB/MshDqP+0ZRB
FHo8LyQdwpHk31NPZDgxrszu/jdYKnPtMVA97RwU2SpScMZJJGroK6w1NZi3Iw+d
jQoMTruwzzeeX+e78fifP/Y/qbyn5NUtLVAPPSA6Qn4rdFC4FS/o2sA0xnWNlMuJ
B9DibHhf6UE8hfUUTzEigFAP9Jyfb8L1TIZxgcKQMavftYeMgaoFDhtRZ5AqkTNX
Tc0S/FE87eyWUMT49Ydi5erlUR/kYg64B9d+gyMt83YvK80S7G86tEwb2L8giRAN
oWQlv9GBQhHbJvf+ugNz5F/0tY1fcz6xVnhuJakifwFHPemXEAvd/JTYK1ryD6UQ
Qhe+ZpFI3BlNARUBHhBBbI9oM5caczWOeGTmqtdFnvpfWPuqX+sda1WJZO0tqiuL
Q2Ed/5OJwemJ2bhbX/JyDmXtH0NB/lTCkfbBsiMhxO2G2NNiFU9zc6DPBuharF7P
GY33bVPHtC0prO8G17blG+IMx3xhURRqmAQ8aw5JbGlAKLPTnJlUkBQVM4XPHcL4
u7W8tW2EFi691awMa6knAFG9+I0kmoE7oQd7L8kG8kuOS0wwuTsxSoQV1hVdMtp7
M1nZuJ1ZoH7FC79Izn1KGNQ7abX/cdq/8SXZPkb0om3hjLdqVS/59ZxCLTYN+Nqy
0CXVtu9pt7+PhSAbgZa/B+2T5jZldsD1ZHgKH0sTyc4Fd2RPxOAVXVp8K9kejPjj
suQ0zt4JLxfwhpbkHLxjNLkT0aeMAkP5+gN/bznfP18Zf8GtiGvG6wctHkX7aO8y
/9FXQ5d4HOciJJSgQf2Bdh0UrDuOzWrhm0RpsjT1kMaJWjxa+mYudKm9CIEnVnXY
k6N/qeeswPy2b0S9je5jkPxlI/1X8Jjo/x4wUqo3ExRVGufxQxS+zR01v0PB9u6J
1oWReTEVpfm+/P5KOOAMbHLOsZBcCjE2cq4jtL2vdTXZj1AAsTz1ElWsoz2RECuR
3wp7gQKeRS2t89tdWhhAhXxk7GnQvmemx+xBYuq7tXow48PocRPJiVK1lSF0IWN9
A2M48GmVHavSpjIkSxwyYFx4ExYTRHIDpfaLt7WUFoik8gHyoBZwVwjBrFwyUNga
0in8PmBB1H83/YD1UQM29N9TLo+i7IF8f1EFnxVwWSpd101/YAPxvjzHg4ZXWUyo
FgYnf/g9RxccwB3c0zqaQywn/w1Qtz6OhdR5vCjTFFtit+zoLD+iq4NYP7A3N/bY
XgTWw3aQ01eiRPhElFosV9Ml0Bs+6BGrvSCUr5nKlQ7QKwLelyrHO0YGLN7BkA+v
hSOnfmLa2KSSuikkQxwPtbV69/yuyomRCpKcL8MbBGk1YenceD/aV+0SP+ho6tj3
Pjzcy3faoY8w67j/Mwkg+5SvlTnXTlghNHMApGK5bmyRGg7qEqVs4oYk72Vfp+DB
LW0D4+QiVu5q4gpCN5yfWvieV0lBijA+g5wm3dSw9tlxFdOLkPctES5Tt0tGh+l/
nWMRwRKXUufibuT26zis9SVsQ9/pTviKDJwBF2j3e4dgM8p3N1CFc1pKFkfidptt
vW1EDFsEh89owAJWCfPpi6dYymnFeXHsjJ4V686anIh0VLAP28LxFNf6gn2F4PB/
gKwwVg+Etg73n6xO/LG6rHSBSD576YawLc8sRa0Lor/nDjoCXcQNJPeXQ3y0fx8t
hR9D8Hb2bKQi76DqENU5+RxBy8I63y8dXgR/sFv2OrmtXC+Skvcfqfs+aSM8Hlcn
XnZeKz1/dpdE6GtKm3KIs3OvCsaqj9FX94rndK1kYkSB70nr9VUD9vZ2pTsJoZCq
cLQFSWV05pywWENebwe73xJ45Tz1IiwhHpxfOJzamBsPUhnxaOWMuzJcqJXCElVK
AZtmrGHxs7BmBDdY9aeJAhphcDBeanliCxmCFvCki1SirxpZjDkaCux+3a7qzhbh
Qu2V6QiiO9l/Ag+jnwQjM8Z1awH2eFQ7cKEdsqjZ/P6SO+SBSnE4xjpeEOKMHJT9
IWo2kCy6Z5SPCqqPoETe6u1R0Fo5G0xvvVA049XtLBt1tdoIHxagYej5wbzE82sm
h1DzgvmILCt50tGkdLTlQka1NX+9OhvLMy9s6wPC3UPqtjSfso6aXhtxgLMzR9RX
Cgie/EXggOa36xmmtVT5PqvBRrKPRX0sMpiBMFQthlQRo/g0h7YGYNLs83lMzmdT
SnadySjLehKCcWaDSuNyhVQlrQHW2B1IwFPoTgM0655G112okrlnv4G1HpKeikNr
mAp+lW+xFbLbF50ph+yGZs1JCfdSRuQJdapUfGmsz4W1OSVk8pTGt4F3STXDpIAU
OUvx8IGE47NraGSOVir96jB17yd4XZ78cjrnKzCm/AcseRXKbTpVFgihYMR56JiV
a6cfQBUBN0qIfe8gAFpj5s5bEyl3X88H5ldxb33gYsbBKSiXW6UbD1/TxIE2HEbZ
zXsbuaRAr8qA4YeLEHaeFxXp1RA9ebNSD1T22K0kkeShs4LgRw22/i8UGOn8t7jt
+sD81PXhVz68dR57QXHjo9jEOID3cEFNRirS3fO+O2SzULavMXAISTSflervaBDI
jrnrHhQH6e1AJy3lE51Wb2/0gO2aurBnGbvoFGlwzH4jT5EfVKL5AQ6a0/pPcDZF
DdO0sT91Obk6ge+kj3E9jSoZzBv9gPJjezTulNzXK1OjORySABskhbrEt6ATaFAq
b3exFAT45KnPi85TMegVGizWmLGn6Je3vIOL1UZIBj0aEqibs0rMcrz2rcUOsfLj
H3nnYtrYCkffe90nCCtNZlfCCvH04mW4B6XGDuQHaUvktWyaF54RvEKbMyF9OfHZ
s/e9HkRr7iTria3CzjqsIGBTLAY0Kxkzci9MFF9SGF6r54R/WdahmZYEuCnQZI0H
8Q84OxI7b9UjbwKtP2AaKBnnDst+7teejcXZTXUul6tR2sZtQJDgoAgkZXaUHwSv
SzbhxW/iRN+A/f2NDNOiWeRqTEX9NwHzQtju6BmaoXUVISCPJKzGISA2p6g1cdUA
XPaRo9FuaiG3tJJdMQm4Tah95PianPh2ouOrfikVcpkGbEj9d/msOAGIjpXfG+ci
6FflSA8kzjUlI7YJrgc/kR5Aoeue0O2lpaKY2G7ONRpvoHTuVe/VsA4GVNmxzZsx
f2VIpXFOgeSiYHvpIE/Jp6gUPUFL5PfDhwpb31QAQlrpB8cEJfy8cJcqxExgmjSc
rOMILnvl/X5WHL3E291/QID1/umzYJOkFSguSmnuwAibFhiT9Y2yeA0oMwo0FX0x
+6TSB8rww05OKsDHHmk8o7O9K1vHzUzrQPKhTpdJdUE6wNtBi6pNuI6c7g9evXiC
Up8nx4nnosIcTdfycuQaVxE2GBgFCzUW4CWlcXxkQt9dwDOFqK0KWYrZ8rLuQu9m
sgm7GJCt/faGHWpWpSO2QwjT83pchctq4NmDAATCr7Z0Q4jDvyzInXhMoDSC7mdJ
uTvfL4K2aaX+S2GozCg3f6f7bRl/u3Xgi2Sak5MB3i5dtim8r9AVPPF5Z+zqLzOT
dzWB/XwOG8PoaT4khY7g0GQdXVCyx0lBrUxV7iUXwAKxCl/PbDxQEnUtg4kBnyMn
0NDGkTLIVlzaOjlEojbRjQHisVhgR57FO9+j57DTUdSw5NuVo++fqxl+tP4eOcKg
uZnWZWHZ4aSjg8BvH1IwB1PdGu5TJEOqtrmLs/2S/qZNRHPMGe26Olx8fikk3jwY
ccWekDF/PQ/ox8slD5ZkbjvsnDntwR99u9nYlpq4Fgr394JtVYbPwT2NCObgtvZ5
lWQ08dFsn30SLXcVuNQU+eb0dsmlNnLTqfomE6ISwxeuHmT7hDKb/0wNB5j24f9Y
bqDHQAJvtZb9FUmAPOJ8PZYY/TRMIk+m2Wcr/O7O39+vISmdXgpEa91yQHQeyqOd
AEfCUZONNd3WfcjguR1I9X+Yxaq9Vim/gtrP9DaXAOTwcM/QGPw976f1675JPngg
Z56YngfnOquQDAMaZt13vGqwTMff/MDnN+lwIRbwCTiMvwO09zXUpzHQYEPlW/Ls
rgqNmiBe0MvamfvNRAlL/J0qz0QwcEC10hi7kbMGBmGI0dvj40J9o0kKe7LTodRW
yVOBl3ez43Uz8GAkdW+IM9cFow5weuLpl9V8wmAxikZbQMP60J23AdiQCALlR5AI
Xp7ZIexfSfe1YpfuC3tU7FfUY28cnHvL8dOv3o8jvo7VVU0sskw8APE/Ddz5wIuz
P5olThVjIBkJYQMf2L1D0BhmbxoR4tko1KaUz5pNhwoj/mSj1qJ9qAoQ7crI/ffW
xn93lOtb8HRvO7n29GQygvawfH2GXg4JQhJLF9gbVr+U4IDQ4eCwMFojA5b12V2x
eD603OA4ZUnpYrAJukj0nQLotqjVASvVwe0aXFP5htMjS2uKMKRDFPgpxCiiNQLm
GbB7dsaCjUIOPj3HeCJHac7r1awrIazXzAbZNcARm+tIbWAo5khfZYA6BPLeUi78
4FNzsfprY+yb2y20vBSJb0Kk+4MqZhUt8cxS5updwh9A2wFf21ZMvvwe1sequ9BJ
lAt/i0/XHm+YxvQhmbBobkGIvyzghFmqCx0FE1+L6EqlMLNOOvz9O0uZoRYErLvP
TsXLCrL08CFAdaK26t0nx2C4INITE9zPWoWucF9jRIOuenYc/Z+5Mndq6Yu1h/sm
vbhSr8qxo6Lb6hbwVvHbiwJv+G9dsS86FLU2vC9zpp31rfzjpzFA0OOKfN8u4QdH
0M59s1Di3L0UvyX1FtgcnXnMEGFEpynjUOms/LHI12xGzpqihzqnQTY6JvAHOEHf
LZyfojIlyThmMr65FsYjUzbK21330N7lE1iXc3vmujXwMTZ629Ez8t1NaizxnHB4
oxifK6ZiHwBrb5zyywqMqDLXfZ4I5Jo86Hx8Tb9awnd8dJ2ISzp7acmRmBnLVy+p
2Ec9X/uNvs1iaCS0Rim5f0ZD+buWdUy9XqytBfVoa/vF38ybhzGlpVYqtkS+/j6E
uy6ZsIdSfQibYI64MGkY/DsGBNwTiiYgNclu03H37q8um5tjUJJBgpxFuxoGgNTt
/0dp6hbnMppqY1kVzqUvauGOcU7mRAp530ls8BOZz0YRzxrOyTmbrHvPEEild7kW
jeLm5km553efXVT2UyL6abYDfTa6IhnX4iEvl29kl2hmac/gqxRcGXZUF+9x6A4/
ZYePpORrBHLj2+0s4XDafGNe6SubsMio6MHg8lP0/MZlqM1RldLYt32nzaeAXm/H
kH+6Cf29AvK7qbJ057giceu52Wv5/Dkb9gNbB5rgGhsT+NI0GEvfCms1yAXmsdwc
5qo+wOuouxHdjN06H1LE+ksLYjlEHbNZOPxGcXfRBVJzYBqoPul5ig6Xptx+MHsZ
5TJZXflkg9RIBLpQsrcaamwKh+hTq31v6vI9djOo+qEN3CS+yLLM7svK7Avi7LfG
sAQLesEA1um7s5/nE4SZxxwLV9XY+ugPAz+N0raX79R3dzxz9IZsymX5awFT9+Xs
1wwKVQwAC44c6PvSRpDywNA96Y8ijbNSzyiFq5XwkriNdsGD0EWa1AUsWGaC4QOr
cLiyvPlKdqLr7FqXOGGDZ18d8DIFlq4coOLWmXgUlwP9uCd1WQq9xnbc4fqFL7Tq
bye8k9XJl5Nd1tvipikZ6y8m9j58j9BWDG6JLdkL99MTVE5IVEdUZYySd27CtNev
9UtrEDlCeLRc6uHP/XyKAY3humC3UCYdJoGptN6GWi1Qj8OtMsASTnUzolvy6Hla
q3/OMOICfFxTsv2qSQv7am5wjZmYJeFcBxzvWTgceXnPEjfalFF8JrCt+2Dm5bGp
pnKilyd8RCn0sOzC4Lhoth2GNpuPSozg1oqAX7O3et1coUz0pNO5HXuKISMZ8YTd
MkBHyAxy1plKNk0V4tXvFLg9z+LyzK8qwomqKhVdFdm4TYsJr1PQGM4rLchimLZT
A67VJFA5qsf+TP/PEzU9XelrQoykWayxBN2w1bhnBBkByIczYoSazA9px2GM8ld2
NL4CffDf24Z4AS3T+y15usmNIPJyTwjE5Xt6mhit+D2N1pwxflRMGzpg7uvqHu2C
kw2sH29QNl1P77IYmcvs3JNG4s5mznEn1kUYsknICRiY10q2WccphigeAgsA1xma
2NRcxM3OMYRvdpjwmackT3J1kMOmqoLEXoEpDDIH8i4KXiILN5W5Zo0rzbu+vV+u
UNc3WXEr9v5FDdEZH417P0y8TBjY5WuPLm2AvSPgCjnJFYOkNKGGz2K33mbzytIs
vDTvqIOUyfipmNqtKZHHmX7cHVw51myMXGf8BS0cJ6baB37cn8OfQifu0QAx4EB4
wfxKwMwBlGukPkLAmPntp/NcyUrMLfow8/h9Zeyw6dml+G085CgIQ5DuJ+KYarl+
Ij2rLWld2uZl2n6p7qXZA+4NQxkPctq5x0IfwAjIV6uHAiXlzrMuPkxmWyAVmqBu
4lnBU60YxPWdZxpW4SqkUtUAhuT01eZ76lK+KtIlegLP7bhrTY49dHaUgSGzgSEk
ttXsd/EoKB5VdXrSjNE7mBeKtEKhM5mQRZjt33u5Cu0cFfbDSyzUUYwRpUPEddis
h2t1utjY52SzeA6I85wbeR2NFoO7w6KAkFrzORJPsJL/7QrRRSMiZoQCLwOM5jHR
ae9gryp4Qk5bfwaN8mfrYj/y7/5erjZHL9uPGTrYNuNPVwgqunYkTxSxvP/fvXCd
e2UshGSa6zshgcOAB7m1jUl4dGMbo2W4ZsAhM90+lrnBrhwGK3BCM8AeRwgNlrGe
6M7ANUbJp6us62Is+FAnuVpRA/GgfJ/HTNvSigTtIhw4aNhEMVUki+SRNVmDrnfS
koIg3mwIruD0ExNfsBoe23WvhC0SIg9fc7MtD21GnbDiid7DdCF4VE4BXlABTSm+
klTpd8GJlmwAFLAYMctcJoVqyhJcnwLoqFEKulpG2DIMK134066k2KGsu5zwoS73
/PIDjptEhGVRk1IyMiR4j8jFrnuFGdY4qkJ6r2ku8oyOvhvoLV2mIBZBjWoYbpP4
ArH/MVSA88HoSM6tI3yksKoiczai0wfXioxdFnDXKa5Jj98PeWlg7aQwt5p186nd
41YdpT9YlvXCnMPA4LTV6fd8sN6g6y0E4QKkhTdb8chbh9VOtlpRAOtltb7VMaWQ
gXHajiU7lmTsTzaZcP7kjXIJGzmf7feGynzQ+xbh1fvxzy+UYaBM4i+aNcCpQ4l0
mIBXKq+bpxQSoK8WYCoVEfgs91UKqPl71GF9j8Q4+3fUqMCujy5JDLZcKskiEw6p
YA/PsCKXKk3Io7ZTqN1MJjTXo9Vr5uGgHZeUPUtb4nT+IzGe5Brxbg8fjw9W5od8
lij76DyiQAxhbpeWeW4z3hISLi9evCBrkwDZF2yNDapd1dT31vc7bCIZY5ck2Vzn
6bsrwfg4QxQeAUhj2spTnEwiziiG6lPCSSJ8mwiMPLFKqO3yXvQ/zwisQaydtMT4
ul/haeow+o9mcwpvl5KpcGLSaQuhMyZUK3ITEV/q78TVcEX51v1a/vttXxs+T6rD
dTzBAHgBGiCm/Ui6xN4hR4xP7vmJzpDdtHob16tNLs6rMFlRD+dQ5WqxcPTKJMBH
gWXSqahFLeJ5pjcgkyRx2mRx8R76PEtIIFULx52KwMMlFI+OrnKnVqkD3AYfD6ZO
Wx12hmlLoOppREIyiso6jQoiJ8ox+gb4BKQyHzZF2+NuefvaiMUimSGJ2W12Wpy0
En7v1OM/gJJjizkMc+Fm2uwE/fdjHu+JGFo3CMDhDnBwp1TfwpZr6wrXrO2bUGsR
RkvJKcyjh8kJXSu3IqHzn/+7pbOXPpgChILUV26KsuW6gBDbpl89SSlfbJbtFden
c8ou7tN7jdwiqzCIwm3hlr5Hsac8GunHPunQqJXycNKrES4EEJ4KCMWpe+0/zIp5
oNCbwPuhOP53fUhnobBgZkgbHrmrzwTSmFbwlMJ4YxK7cZ9WJwEmFDj8+pqAeFZK
njHxTouDKfaZFKorKtOjsH/Fx1PWifW9sMXebXYI15f6sOZMYNrybfbIeNM7uR6+
lttgWfopxaueXyAwRleBFWbEcbdp/+U7mVkJe5bhQZ4oBflIE71fquviJhQPFcqN
tNxxLj5gUTHvq3ioWS8XM/5Iel0F/jL+My82INjh00kJVXeLZ9TlvCeODmnqRHCc
ULpqU+HimRElvgarzm1+j3cyr4x+3QkCB8fzyaBapK43sdWxFamUPc11V5XVURrD
JMrkSzb+Fe5AEnovzDjJZzHE5gZrcZ77hVA47f92+S+Ju584x/7lFVqcwv1wWOc8
j4K6g61TWWSjsVdMYDjT1O3ga+R2G4Ro7lr56o/b1dmQ9yBImG+Swhxt0x7l3/J3
dUc20+Cu91YrShMBGE0shDKeWkJldbudepjpFxQA40FCJAwOh+nkz3gvUyKwpKJu
zNm0VoMOHNl2XdmQGn8auovvwZDO4UxEX5dLX/KJDN44bOO5atE0CYSM+ylRZoWz
S3uVBNNmh9pAngW5vtFWhMtyveSeuXKYQo1485jjG5HroNhCHAPl8dr558XGDlOu
1xJBSEdONDFcNomfnsOK6q0lC/nnp8FFkDM3PkWPfWSOnPkAWqwkpBM/IBEBo4lY
uBvVHgfxMqJdnJxDSFZ/kI+Jw/SubJBRIuaihEW6BEUKcwSGn9ZCURZoQNmyoosc
OfS6LT0wWEW9wZQohDJ/7sUTXC6OI7eoAwQ50QqvKa29s8wLBM1x+r6f60ZpaNKZ
+2ME1FoN48zuR8uKz8eBaNnEtzgVlikw1pZjZGeFQO+2+1juRGx39BdW5ZvgnMdX
Ptzz0xqz0h9jP/4SBOndqEmcg+EDqeVRq6xtFgfRNaWKj/hexGpnemOHGyXkTlDy
qC4iyHzHIh4eeVo13XBp4TpjSOomoqldPdTE7MavRdj6+bLREiCE8A5rWPBi2MXH
3UlWR0364bsTCLl9Eb23BQupzK3Ykb0f4RBKHmunrq3ziNALA/MdBUKSrIDTwmc4
UDRhsv0wf2SEDExg+nq+KdpUSFsAQF3+Lna5j1+DC4iOzEvwi0ThjqXjzOAKIdgW
QtA6+ZdLA0C4KJ9nQuQrZO94SF+K0lcEoXPqx54VVgybpMfdacDbi+kVe/ZrSZtV
wpCEBc35CEhKw2w7oPaxCYd4YrNkB76TFnaHvzA9w+mTFbZoc+HBLsXUFHM1UTYd
NVQ9qA6RlP6Li3t8jfSNKqqK34YdkccMS3iRPBRqxrEgW1Jd5PilcyiNDvIglRDG
5DrlWRgEnmAcRvyYxLTaNUvZtWa2XaM6Am2qyg99ghd4kAyH4wJa3eqrgKhkz5Zj
IXUL06L2s+mR1ZgwFjx1L0zajU3CQ+HnUfqAMIsAUYkg7m98QoWK5lsF0bscnxwE
e9/GkmVykga3Lfa0qLjSJUxlx7fzSoylzn6G1WGDMxlzkhqSXQZVMCTqUVkb/0OB
c1RKTVvFjSd982GjTS6Be+0iME1KpXGfWb8IKPU/jNnzNcym5ovhjPs2y76ODXZo
HSYeAplt8nn4thG3/IMPLH+T+MiO/WVzDg2BMdflsgXPPmlS4eIQVa/j0+LV10Xa
eblmDm/cmlUPpgFF/EreS+qSGi6RaOMX8PcJthTVFzE1PoD9aiG/0YB+s241SkFT
x9LpTXqeAGGMVNfVR4dFkWLxpxYr82I7lgACHJcsHsV+NrliXgOTlmcMynGfbXyF
714d2Qz8celGo24LmvRt++jldv/x82soyRQK1rDGlO+JYHaCV4OBqLj+tk19PcQD
EpOrZTWTC1mTcDs9J1CbkSoBwXrY9fFPG0xlFe67CI2aMa4xHHobOoRMPsMHJNGq
lBacbEnE+QYvZAu1Zbuu2j+uul5nVBo54RCmvOyYwdnzeOaVVVqUqbl78cW5V8sd
L5GpdMOqqNtynu1bX6ayTXAiehMBNN4MzEbxY67vnNCUamDt42AkP48a3vQN83Jv
+XuT08Ey4F+UHYBvgcdxwAzXkJp6QFbdtf3wZPxh2xPhLNjMDlmJDkZffhwI37y6
1oX/EEbc9LKAQH1x+yAQbe8/Pfir3f/p2IVFYECdtIQu8jdCd/lBCz37l2Yewj+S
fv8YDSsJexj32i++t6yaSvW9BfjfDCYe81S5SpR3nBG7+VgBa07DSjegKZU8vTZw
Amahm4EBhV3sKTikmRVInfWZcpqugPwsCubeYxU8QkKRtxQsebLdTjilb/eg6SId
/eJlyXCNFI/rg/ll02OQB0y56dEcAbjNUPeySn8HXNZvhdoATTcIORz7OmXASy2N
fAdbt6GH9EKqblhnDakiS7XmLIMviB5/EeQ38MgYwmVHJz5xVK47CqoN3Sag2XxU
b1QLmOB2iqJz00cQhmST23w4sPYD91xzYswmf514pp/RzIrGdDW4MBzq9G5kngTF
GnB0n2B4HQfqoIu8cmzoLjG+DlU87XmDnQMF1wWmRsBL7SpaJO+5Ikfd5vKvA0qJ
ObiJWAauquoYnu2VQIWQ0mDwfPXtM7Rexxg2Osn95lAWqaofVLXgOEuRNjMfGV9J
XU3OOVna2c0z3r3eOrO08bm18T9dyFjhsoDXPdDnonitOFLV7T/lY40W77KmAyWK
KSGJwWSLLVG/kXiUDAQaU2eUxwPvBtjXk6nc6TN14sKuiCjnZZliluBH6KXn1a/p
evtMX0IsYKt7Uw6YK/5jxr4Vf75ACC23akC3h6flR7az7L4/hkOe3L3W9CalJUYx
RsTAuJ6tbVy/SMVb2A+ntQv4IxPor9twZvEbDwzf+/Zn9nCpe0mjj7e/eol2R6MG
OLZLNRR09S91Jx8SPYjPedQHOLPjTqMo5U+FB5dBzMoAS3mA3L3DYEAjzfqAn2Kh
H2hyqHcy5zcoz/bq97gDMJFUX5GNfo+UgDmBzaoo5Z76sNkYNgA/HfchXRT9L34D
TN3CjnjilWEz2/FZ0lMXA4WQd6XMwoG8n7zva4675WEKp1qPop7P5JbyrBB+VJxF
kZg30aOdLoqFNavew5wWMCyTfdQJEeLFhc+gAYx1f7UMxj/KWwxfIil9+MKASfDD
YD3V+7uqaB0Kpt6z+pdC8nUVSImQpIBjdHEcd50HV3gxqPFCotoRcTIwLLhjZQHO
/EXFZ1Lqmh1TtNcHuL2LKk1xXjrpFC7EvglhUNhXrkBoL7RabsSNo4vNI8WKV1Fw
tleqv+yy66RnYsZcDrfFPal/ikaWUc0TXhXm1j6bawbb//sb1IjF2BMGI9j4CVkI
ylGXGEpCDKJKbFDv7mWOknmCjIgW/JPXMZpR7A7beqx6fMrTfAkSh4EKah02RfxZ
HvqRxV+U+74A9P40GR3kFubhOE6Sr6+f2p14KnPwvbtoFr0AQ7qWjhvVNV8fm1Zt
A068gwFvAcKJovQWsNwwUmFks0wrYlMxKBUlpRt//hfS4asxnU0dAmTPVaHoZmC5
WzKB46CacR4wXiBlbxc0K6t0AzapXNJEwYMnoQBB9zkPY/+mAc8Pkaw34yhdhD+U
5Klrdc0H55wlfy5I4sUwooYVfb2gxlBVQRFsGIcO+na/HgiliPmodxtUonKr6o1n
dQekbvNJdRdVwxn7sxB6zgS+wqULiv1AVCSMD5MBTBZcZZIfFPn1edoO08RSFUOU
0FiUKgpRBW3nPxRZsMtCwHa0wrGuJut6EOKCDimhSQh8sKIewlvJAwUSoCj15QmZ
qRdBMWyqD8KdaH6+14irFxpAGN5BaKWa27oNiRs4oPpo0tvJHpOv/zgnKu1fpWbe
zz/rXW8qmF8bCrHRSwFkTDtH+rdhzyIHl9wg5p2VM0Pk1/2tdSKgl/1mqYAjAF9p
aqOq7TzdOgsF4diaymiLt8kYWT3zodmoD77minC1x81SYj5fZmGCmjhyDs5oy5vW
okvY3N44I4a0cQmCpn3s6ij+Oub8XsS8R5AvJGMwAM6hruNuGlCWvRZGxxJOk5cv
mFCcRiTSDvfNUxVEL/RUzvUP25qfC1kCt6/YVL2oobt9GFtqSRYXqsP9T8BzOEyG
UGVioq9pEQ/OaUFgApWmKYCuDPrNJw90NZW6t24d1uPRTVqxXvue1Uvk49Zu8KrN
lSKa6uJwMy+oLSzh6kYnbxfvhc3fgWh2oAgTx8NtsgIx0ZTC5ZGcwPXiMfZUxgdU
XCFPcicPtB1w8JPm/1APXsptf3Y8URBGKTZrfyLjTUAuJxi6C476qo3DA65uMHqJ
Ou+xtKBN/bphtRZp89iZBksm3tfcqf6XzcHmq2kYmtThLhXPC4y/V90hnvocdn4K
u4+2esHJVmyTbhUT1C2uMiw7rXWzu/cPBjZvuCxrcPBrTg1bRm5GiLoM+TCp3xzF
uCPslf8WD3Dp44KwiV5T8cWHXFIN1D91d7CgcLi4d+DIgFbPyWyn3cmZn999fn0E
KWLa/2mniKouVt2jlQlPRBu+FnG/QOZ8ujwaz2vnOfPl1Ws+rYRMaA6yaWfCxgSf
WMX6/K3E6ldCKyBhdvPIq8hJcOxj/xYoq1tvJLlnm0/U7vfaG1T1P/r/M3ZciaWd
a/Bx/672x4eTB9sm44dLe1m8Su9UWPHZ67I54UHQ/i0X7fP/IIV5FqZhMNej0faL
Ef5du7h2sKn9eUg2LDzl+w7//ZzKovhTkR/GDpBGD3i9bHai/TirVyv/nirh8TDW
YIAVkxtvJhAgvts6qW/Ut3duDmeL21IA4DPPmYteC0bVvZ6enn7hwjFUcJdantBI
e8JOtjdbS0EC4pB3Et6K/coEO/uYvk3G6oGGypju5TCZoUAbfK4wfosKDAQuj4ev
ivYuotpNEv6Uzspe9LysvI6sIQud/dU3TtbeECmMtHr+miMLu5otTPu+ClWx/zdl
b5qwdAuVHfOoGlNdT8AP1a9xmZSw6+QaIJSPPQdvXQtBpGZeMrPGoxsbPwljvji2
ghzImf6F7Y4x+C0C1ZDWqZTPoXZAmSocfoOGY71J+puVR+T7MXhXXiLv7h2trAhq
cJL3XHTXH9YgViMGMLqPjqEbt6rfGGYgBUQIRs9kzuCAouinBZ72bAEieHIAo006
MUSBvDu2m5y8ntR+qYECuinL/5aPuY8TacVI5OGcsbQMyF7wZvgvcqT3s0KKLTzQ
CqtGMtoTjK+E3fW/a8kFOjSpdN4Ejvo2OtmutKH2Tl6VTR8MgMVQZwxntducniS+
ADDFfJ9ZZ2BUz+s9EWbilzgP+OpwyFsk2+Hk1lbLfx3AsCN3ybx0hgyjyVeoAV3I
wQDiS1f7WYZmjMKSn1W2zXXuw1zcO60nvCM3u+VENZLj1Ies8bXClfV2vAKfGauQ
JNnqu0wEfii5gd9lcYdGpjKmeMHzAB/J8LHPQGWqtjqp9krXMYLBU/9+P4QJxbBV
XQsQl4iYLyNPbniFnI6fcaUe1d2jmafE03qkxjU/BS9szokViMe4yesSl+BP0kr/
XZImiJVwMQMHiu3oZW/tVsDaQryGHdREFffxk2mAHHw/e2aIL5ycwLjfjMunW975
KZBCClj+qzvUbo8+ux/FWK9VCcFzAZ/llc2AxobI+4L+Fh154ntZNyaO4R8t5hr+
QOkYT3CfKEVQYozJM/TqC46kXB6D8Ok0NXKBEPxAEvSWuFudRBxbcNWmGlDEyVtX
qP5ZEp/ddIauDzQo4cyz+C86/fUf5t+Y/pryc4VBvs0ujaax6lxDYWiq8lu4xD1a
t7DGc6sQZNHlMg4R7Zt0dfpn8XK/SfLcBzX7/KcjyhRPrmqCzJ27iGs/VEegKsxR
FJh8x3A+pj12vo25RcAukWlOBVO0BfU07wMruJm3WKtZYDl4yvj7FTzfNZTuC73C
wXkLN/Yw21hniTZK0sc1ez+WjvyUz+YuVjyQbOCdKQpJbVpOtQLF96Zkasbm/MTR
3sVnMkitCvcCmrpsELvOW1eaI9OY2//XHL+3dZGxWy9DllI39ul0qycA8YcblMhr
qnJXTggTQaGSe8FYAZZN9P3064XfSMJsYtPhJc9vegDHiHJs8FXPFpgTDK5XKofz
G2Qy5l2v0e9lRwGOvsLvvAbVQZ2PiQ9DBSQ5MsS3G6+VhEUAa5jqiLbAJYKABTEu
28bbFwG5q0h9t1ilSiH2dlNllN4WdaCk+/DgJXxmsmVYH+BlvwY49RFTQjp8TQP9
ZMP2Wd1qf6HE64ivJDe2kIK4frfjcQlwIbbVBc2vkSFzSHMGo/twLRQhb7A0sAqk
wcwWY5waBQh3M16zd0DTWjMALbIyVgNEA2Zc7WqAyhVcrTieeDYdixRn3enFulbV
ju7wuX7MxDWqGSeAFfZ4aR4VLCXlKcaVCjqRis/FhzlcXJnYwbIo6ZCMX/5XL8wB
kurmM3XZIY0NT/P7kBZ/RbdPG/RYoqzls7EgXXKplhenTdSBxUldPhWwlukY0ezU
fxcvkciAj94AQK09QGtIMDxJ+5wCpNguJtiT2NJcqYlSaTvamefnGYWX8HBgBQJe
IoX3GFAVx4lJngOUwnHPaxHVfISQpC8gndf9PTgSaz0ZEUWMQlMLpo7g/NwuR+81
q1h9FB4xgBPOMRq5tNc+c1Wxcrep9jdaJg9DD9UMNIXyoEVeIX4n0yxipbiaIaEn
sngmE26AKiPhA5TwKL42JcR7YduTekRw7XbjlFCxFgxKja09ra6+/UsaBmToSU5Y
7CJpe7MXnZDfwH5200Q205rj68vZt53X92Aw1N7cIBI13nfhXxb5J+An04DTHXH0
fjHDKJmWp1tNLznoKFrdf6I0qUVA7olu0o2GXuq+slCclOM3NSBgzlAZ4wlZEKln
auw+Ofli5jGK8CN5ipxbJ9tJAVdQ44xnYUiS8s5BxhJDdjEhG1omF/Ju5zoUrduQ
M9dQ9D5XJvZdRUvLMfkLAqSzPMRjo4TJe9xNisANXXxzZDc0589wCVmaAMcgatKV
qxr8F706DA5D47RppLIn9F9EtbnWO2EwArq7Ih++VL6uyDhvaQI8MbncawVOhyVj
kyqDXrD2jvQW8tpvlCoHpoLKSKUUDliSzGl08htzGO+o/AaITG0vfuq0NkCtyxCI
HukhMBicsSq78JwDmqq/wkP46XyDJyUkcq06SbCOAwkNzbkB2vN6Evo2xGwaz/om
7Oh0Mq/T3f5HHygJhrjstSkT7eIE5rfidzt4us62//3uu0kFICdi/quaVJtg/LKm
bbXMDxhdtPeI4EoG6JhlOYatvPSRdRZAGKXU3IVuue2iDtbUgsL9QaVpMB5gpdSe
4jU4CGIK/hTBOFcXRw8AWxb6oDzOY87I3GrF0Uzvfe8ieF+Xn0PNUifYsu7fxoqO
p1r0bmbjQbVl3VA04dBbiNP/bu+/3seqDVN2fUDf/q4QJiascRdRVYsH86BpJyHR
RJ8IO3QJzQFOejBiWHso+klRwBKcO5nkF4TOFcrc42eLmFk1U1MZI2MSVaYLA8uL
UL4z8WO32AlqoRAkBfJlWAIBdFerfu8dBsd0Sk0vYIg3JCfAKnfcc5nQEjfC1YUs
XiMBQ3Ef2ilJD5xeHWIpR9sJaYWDTvAPnAtbg9GrQcjxIZsWWQBJmqrcxMrJKacf
8mphPvpjDLbbyocENahXDVTSYbQ3Q+C4bSp3p1w1ocGKA95pIO+zP9A3LaeTrtcA
yGEda4SwaSvipS1zqSfP27RKlEgfg0SBWK2Y082K1GtnE8oyyGBXdm7kZqZgVDQE
kLubzkvDgHZ0x9C6V3BYCHoW+L2RLt8aaiy42TqLJAD/ESrOEMYSalO8HOIuSUyV
+i4HNeY8NMk0e4x4bXk60j3RWMJHNVcfRcy5UBihNB3uBUDhL26rkeiGOZS3gX45
rlP9QwMW63orKKl3UKvXtCPr8RxUMUa4l7d5dlpKzlk217Q2z8YhOX4vr4dlX1HK
ToyQHrauMgOoICJQeSTubewM8yTFoEfx1cdYsmvAwwN61ZfEDh4XJcwT2mxCgLa+
GjWQzJy+rylbuYLDffnNmThyMHcAaiXn0Am6Ip0TSwQvtuuOmOk88+kTkJfQMnYg
OzWFMVZ4pPSsPt37hzt0VC0vVwDxuGcCo8ZfSWWfgB4bww/85rfKBTuQYtFJ/bR7
GZWMdnLzosieKAW0rEwjfEJplYkSrpweEePx/CnI/sOqJ+Jw0ACkYuT5AO+39W+r
CU7jjHkxXti5lWFipl0omdts1bTENCYlGgRx/yiyo1VdCChIMobKOvNDzc3yhBFR
3SotfNl7H7QGJd/vjwfkqsZ2tvfxUApAWYEvHgbOSNs5XOSeRz1aRBSTAWtKQBoV
kTMF+lJ2C0/XMuBbl/NFGtuBMI8ocTB5OplLOBnMQe5fLNm+O/+c16o3jNR3gMR8
eOxykNWtQEHuOQToEk22MXsF8mtB4MEhvmWdUTM2x2qHggOLNDaWgwuDQ+9/FZh+
LMQgawguJ8vghqR4Fn7cGH9udIjueoOUTL6t0ZtQO8k0jfWeJ6inNU8fYKfdoOHw
cWB41lhQEa/o9/fauUBN5LMMR+QVRnBC5/6yx/sPQedpbC56dwnzo3ji9qil/kcK
tbypecDvk0t6eWQsSGHoxMiWmGEbpPnDtGBiDoslmsGKZZchN0eKM52xiruItxib
ynYCaDNM3fjnj9+mmz4Gz+pzw2ZUt1agLI28rxJ/v8tewRDHk6XT9JBG27DBJ5kN
WlLLAIkf1ldMTrTiJvlu9wZe5SYmXSs6MI36i+QaQTGe9TZ4OdjOdfMiKe2o+nPL
hRsabkkr5ZuFGa/Y94GylleJP0leIslHyMlmWYi6/n1c2ii1chcjlgFTyp9kFks+
zyFFxYNGpirEtOXuwWrYQc7hCfxlsDpqiNRWNwqjkXs4AGTopgMkw4o0iQYaka2Z
9VN9ENWPvDUVKgsiWpNrou36ashEaisxukymjePILUN9CJcDgIyIwBUl07O5USA7
MbCjR5AJcODO7+dRYD9BBCrKuFE7oQsNdaOoBTebYaek0CLRu3DHOEG233C/CaKF
rCCeBzW0gtkbP10cQylPvsZattayqw9BpDUz/HMUXJLDeeClm7/T71VPZ4zoDpvu
Y1u1uYp1uZtywrLM0o+CscJNRgRe8SrwlkF7DiUSY1Dwaoa5qAxxYsu204o4kDUr
3M3ZM1CpMkoZv4BzDuezuBCy0o7D5aOrdT74yjQp9998Ytvt/wmTXRpjEKMOloqP
gwvGcTGij0fm/ELni3Oxzu+LWmRgTjvBFH6iMmt0T3wzzAPbTmOUOPLjGYwNWLWV
koNr/FG/w1zjtFWPjaY5yk6JBi6opwt69g4HwmCqknGJLDARrTrgfJmRL9MvmZLW
HF7Exk7CRFP8W3UY/cVoAfmwQ8wDu4LcPY1b+MelAswkfEJOQQzYnXkseVdUMopH
URjd4cNTGH1jbD6m0B9XNF7I3r8B26O4wQre0w6DIyyvAcPyXD7U3iwaZUjrX3CW
D8cO7Qa9fUsD1vMR7SuW++pcUsTJ+4tvsqJcvMuYp2d/zsTq3uwz66ajqHvIIyf3
1ujCeO1nh9x4Cch7XH9tRoMBbfkKNyP0akwfFuDFEyDKZ9H/veeXNvCvp5VD2xAM
lLnN8iWl6FQCcubXTljBgXQk7lkaYgGiXzdtT0k+xw51MN+sXEXj9e36Lws8TKoP
uIUXiNJnwuoSKD/+lm/I3Rd0U2Sh+c4I4XuSj5DsHrGGF4ajine+jhyMgqLI+bZk
HgcBJqKfZ1Ws/s4RQIZmzUjAwWiIJiYc9VcTuQua0Lc1cPqAtP2/pvwNnut+k0tV
pBhpVqKp3taU+zxpo8YqLf6hGJXhL1G323Gj2y7hTDtsXMND+k/apEQqUK8mdmZ2
/oXqmgRlVaELUDjrES1OhIRrlq9gW7AgroV0HfUPwkQKFFJEPaM0K2exiSfFocFs
ghl0QEZcNV98xlfMdLu8A1USreiM7XemkV6EKKCYiw17PJ4IyfjEQibTqhIkcUZ3
9+MBCkSPwSqk1ChBUbaiJV3bpK+2VuGedKC3zi/qZBPjEPS8X185EXdZ1IoPC3T/
Edz9kSXXcI3GBZvU14VqkXJH8FELPrOxinaiLPFvOXKXWQ1BwxEieGwUT3r0VZaP
1HpTcs6AzzsuXjIU+G+BQJJ1r5qc3SZlSFazwlhlrp9qItNeAARbP8f6VljTw6xc
HRpQ27blVA0AHfIu1Ab77JOWxzS4E/N/nRhXMTRjctlOJ/ZOq7TiAa6kvSww6Vcw
LbRj30ji9KjcrAsGLHy2OQoAR2FTBUtoopOYS8It8NA/PA6E3/rH7gQ6EXt0XEON
guc7yeu6BwXuwcsQQKpDU4kAAU9RHcte9xf0W2/JopydmjRhfebwCVm4u0lFPrR2
SXHSJJkIM+CB85aGRjapCie5M+7WpAJQvewPNJQwxPihHjUck8ey2XDQQC5aEPdd
WqvJfPV9ARUiAH/XZOKjOhH2mBNF9Oo4Pp86+mCN4z9K+/JLttB6j++0R9yojxMF
8z42br0xqUgC6mwlvQxD8VBzFjBzYCNiGtx0C07KZXnYrE+pIB60BeEia2MawfzW
W2IK09DawgO/xbsa65NSgBPabcJ999imJQ07sKLi4jGx7In7XDtmgx3PJx39fq0k
wQ+xiMLBCXz6eeFM1VcKUGD78x/83aE2E8TDE4i4cEPM2127Gvn2AQ85r1jr20iq
+uEXkeCLBHjts6eI1wrvh6lpJkFcNTNvqrFlN/a/2+oo/MCai3fIZweuDoY8/1aL
rJltHn5SBrHriZ1eDmtZrGjq6ONkPkE3xX5EvSEuYnbi2dlsZhr0dcEVmus5OyoL
3HaMKPtZ3sgEDOKCkiPpMzbmTViplXXZvC6p59FjoGpUP2d8LA6kEpxbpzHraoiV
ueci+I0CjBWCSzb9f11wG7s+ELSZbyg4aQcatDBQMsVuxGsjXMFMu4ACV+ofUQR5
EYaYdQw6I+EnKGr4yGqSRp1FMFHF6JEbvZd3id+IjvN4vpfADZIfJRzouR1fvwud
lOrIJASmmlavl6Qlu1VAktT/C/Cl0vkzu+CtB99UOClig+9OhHJvznwKvtdLTgGI
bxmxrzUJiwK4DWKLpU86dC/60xc63EGt7kBIHMr+Cj0kinpw/bNZWcBqGNN+qGfJ
Aun8BJL9oqpZUNpz4znuf9Mz0Rm5cSg4by9XYc3maryi+dvv6xUivUtycvwuHCBp
4f1+DaVSLv4ir8T2uY7QLjL+D5PtKOMNz84KI1q9bRqg0HpXqwEufPU3fBLzsrO7
QB0AkYFKLMbGzW4LQ+bSjBlIkahLAkmfeyD+baICuSNUtHy2Gr2ptGJhWWt3jqMt
x5CyZ6BT8odSuKkYk0rKMx9ON6f/KjaCjYhvOxLyVNk8SI+Jzcti8Y9zsY8uc9Vm
D+k2AAXFxfGZ2MHVkpOlypDFxr49p89ysnWPBNN4jIbsD3/IqmeCmZR+RN0Ym3Du
QEsaHjHu/Cj/BM9/POiMm6IPfcN87FDpGuYl7cVDB+d7SQjxghBjxnYAjz2ZjpnP
4+wDFAt0Pth5NRNuaGx2gAjTISPmDnI1qIhSsvh8zC1eEWWyEmM11yoOTzCX/RT2
kdq62kho6cA+O+5lrtJ4QYP5Ap99HNSeV8iieZBlABxtB9zN95uGL3NDqoUzAiP5
MKyre2t9QT/f62qDnNGyS+4l0AazBpvCcYwvIDLVNkX6o+byk6aDJQ5j5Hc7Bs9O
CMyQDZN1Px7xhUqIeTMSJWplBxlyK1jsHxCzQGG8BYSM+KIM8zqwdADCUkVnXPC9
T1Vv2FWebg/808Z78nxXikzoRmJ3Kqpag6yIAXHatIVzrpBdXr4uHJwBXTQTRH0D
zESPTUAZqv7KJzGNYhF1obdY0uEL5qp1jFqFOovg1lcNc1+aee9GwDtWHziG72KA
zeLmp+xni7cja4YkvhxC1+kBerQNbQ1pvAzYhJbDum4MWb/lWk+dXLW3fdip9xts
ebQ5kEwDcP8KIpd9aqZcMEXEweO9Tnwhp2mJzpnRpCFAZlvCQopanfvuknXKAe9F
0rWVupQxnzUnsaLaZdU6D/2l1IAvGgheRzHfqU4K04y4B4WdfWnPQeixpAXbTfsw
CibX8F/feACNdMWzJAAwQtFmhzh+A62UdUFvyJiJktHVYzZAkiftJAcKtTGq0Hl6
VlD5OY9GvN3rfwOZWFAP24DXHYEP/AVKpcM7DN3UJWzrZqIhMqcKzd/tzywrAupV
OUy8zrTxlCF1nV8yw5UaiSX9/5UjzRiKz5R1wcCUgYGWzi24+foQGdpQH9F7gUi2
Vvd6bXy/IvxemR6DqA1W+fxmTia3ttxZ+Hh1nlvW/XOn289Ybeiu1mYgvDeAVUZS
DqvP2MRmoguVpt93vLaNuUUkk9LB4mcHalqwJfJ+toAiTKyRQIZeNouZGjBLedr3
+6jTOUKLs/OQ7eN/xkFILJfHJ87jUlBsQvJ1u3958NWQOXflohvi2yiVg7BXaJ03
dKYTte+SC6KcPQ76vMn/rQOKHL4xZPsW5txzitro6f1qn1AD0J5U2JINCoPQyPW/
eQAalXhN3g8J30UvoXAik9Ap0IV/pZuOyS+fZ7kciaqVxOrRLk4o46mab18oH/PN
DvLnr/vhyXAENOnBfDRZgRzp9097oHVecMpRqvd7bkysLfddjcnSwzg+mwO20/9a
OS8GgRDnTWjgXVh7lhcSrktWE2EyIijuCLcs8lRF0MDSgbFL/9Yto2cutnubGuiE
ySqnGT92AvrXdL87wI/37ca6xEmoqBGThoK2Fskt7NNwdJrj5SEcRxFmAMcQFwzI
/SQmJDUyslakttWy0MjceZJq/E0wyU/SF2bgc1+mMyJvCoEfRPBYN1SGWw2qVo9E
6iws1UoJ4OuvL7bUZDfL6qtUWYnEW+kUwoaln//TKHNLNojjqgzoN5N1y8YvJK7e
Rnz5xwka6x5mjiqvl8XSbfnupKiCfbLmGe7t4kp5DUjK+Jh1BpqZO3DPDervz2a2
8ftICAnIPH1vzG/XQpIfMRpRuZrD4OVvC85JBjmEOzH7rWpjR88Gn2ZAGxgS2J2/
uHkuWmjTm9QKl9JduUrt8ZC4qH7vvuDqoR+gGx3HfcN+D7mtGN5RtEHZWrDR1Z8Z
8Wop2n04//8E9HDMz0sXsQbDdATmcQAPN3YbnkpbCvv4gkCKVry9QF06iZC+qAoy
UDcRQY746HXT/GQbxlyCFPrlxuiLIPmafiLdYsGTkIq+0IkTwtlowbGdOh8F29lc
2uWJEfXFRoJl8duPPy00U/6divMXeUM9aOshe0PcCEuGR8IKKfu2nDpXFXcezm88
KFLwhoQhHLhl8Ki8yN4WPB3ZkwESSYIMgYYYZqjSwnyKq6KOMQ86v7KEEJUL6iPQ
R8gFWjM8HyyzTCjNybRkvlag+Tw05mkReGP6cFWm4J7TLZYO0WWu0lZXtkBbn1DV
KehI/2yYRxGqSvmBg60RGGDU/cki3bPZiexY8d09agY253ZND46/XJWR7ZdVuNf7
kyHplEwyS6ZvOWqAkO21Ysx/oIGb6iwI16uiPBZ9ODPcsoPTCFrv4OfIKjgV9fI1
wPVqtuQaTjc5kN5rtVCsS6YixfBYMH6bBAuzH7j8tAyo0QZqEodWDLmIyGZO48hg
Or2lihzivbh7zh27eGxPnUrjN0MJ6/nBcjBE7CrCma9peugPQMmuWLHlYgH4cQ5b
E7DxxF1mKWuGI8c1PzEL9d7PD/kfMpHdYkad9j6WlvRwyQaDR51B5r3dQUmZGZAI
xaiZ7Q5ncj52QJkX2X3Z8Ml0XNK7j9YA1RrzPAs0UkJD7mRf47UVQ1OsmdbrAexI
doZQcKGx7NlyjaIaoCZUnkUI9ceLewdGIrBMto4FKbzuo4hTZeHttE5YEA8v+hOG
xn+IKRtPgXRD/sf3HwkdeAiBUbr4Eh2QdlCOJxihgsnlst6WJv2wy4hQ19stPtTo
fo/R/sEY5QnizFYjFFonuc4HzlZUJGaSnTiJHNgPXJpmsBLwskfUO7y133BIERyU
2488MvxA3PztDGSfdO3alFEp0Snx2AL7H/OGI1iQcdvskauFpj3gc+glotjvlKUc
G2+cltuEsh1CjW+/u13Dqd1+rSdXOGn5EVgpdRlQ1XVLp8JGHvPj+trscmpCgQG7
efm5wt6m+sUN+j1uP645UkaKKwNUtRsSsGk4IjfRgkzs5k4QSuGC37xi2NDeaVnd
r3MJ2zcF8qD6RApPmfRwZiDwm7Nqj/5nb/VIoO9qH7++CeB00f0Refs2DuYAUcnK
jIhAl47qXOKKADG8xhTTsQjNShrHP4AMKE/v7ItEtsY+NgUZvKDhiv8KZFfOAeHp
SQcHZwQ5End5QS1ksSdiNksKpKJHtqocJRZPyKH+Mr0BcueAD61EkDzYQUm0MRAb
YnF6jtD+bg8WHQJzXP2P+RY+nJxRiNPGtWxkyfftFsmaVoLwmcqgWj5SUOzmE4MG
sUwU3lIbjEJjJ8WlVVm3z95Bha9rCLL2mqlDQLUY6+we64/FXwfADI3GnMtixcHp
icueeAJNnABw2o4pFxmORQSTMGgXFCC6I5KYgPnm1q1Y7cwdCXLRhC6472Krd1iF
Zn4mn6cfqcyUfAX28YNS78qyQywAkIiqATbcCkjQVi0+2IjcaJmlt3k0kutg4BL+
O2rI8ad1Vrd07n2sACrDr843PsL4SkhCJI2Nz+n1k6+220Cdeh0fOfYzwCmWz/6E
KbekJWEg++Rul8Ty7nXqMDOqnP2+UGWEfwgHwp9ZcLeUohMp1WMCOdk52AN+2SsY
0ybmwgavdPt4phP0rAFcDbyuCD1DdP8rX/98Aa3Ciu0gGq64PQqKKrK58BHMCKE7
s7wHglYvhk2jVIpa8EVP2HhXAqLm51DsGvfhmnfX/xHfGt+3PJhUdr17vGhZChgI
ZbdfSSSPiAaTNPG6gm2U5fi0sdb6KGr7jNDrGy4D19HvalaCzK8mHSlCAI1EwYYr
3nvO2s9LiDG1BdEyahnCrko5Ox5j7zpr4dibZo9bz+aTxCgoJ88xFDaBg631SwJ+
5JG396fsUG9ZM52N7gt4nBdyJFzAxd0C1uG7r13ndHGvcfwTQpMuRC/W4itQfKa4
mToZgwBKHC5BZXVY+tvK43HxrcAme1dTQ3xPBALQYUDP6bthsiFebSTzX/EKZqYf
a9oZoAVBQ86Q2S2sRlSTqg363DHptsJgBraHeo/n2gwoVca4Y49SGpJs1RSy6Yvx
T8CcrAU/GlQl6XloUPIROzEPWPrvBOFuzBvPl0zA3YUK7+7HKg5W6SiAHnI/j+cP
LcIEvQfAFKIjhJuqEajCluDN3EaVK5XJKgvP9YTSgFVxrgjIglkV3sfKoLsVu3q9
KPESiW4wm6vuZPGO58q08PwLdqtFUPjd0xdn8XrJY9NTzTA1k9x4g1Ytbd1wJWrQ
y/mIqsp5IGfn13M+S7f7TNpqda6euHsJv6bGG1yDqSX1rjiT4RALKMpmikqvtBh8
9mEGfUQ6grTV9OSh6ztsAtwqxM+TfA9MDYsGn6zhukNAaXyDhPaDIXko53bYq5hg
ysPjVhr13hy79r+HqMtyAsq4036BBXt51xT3MYO0jf9w0dyJ/zk6uYXzWe4cvGa/
LJbi53eYZU8+rPiaw7P9uE62//9Vj9cGDmgaLOewHSiyEWUOnunIn38WZs6mefTV
l2/tKaeeV9ZffZy6KsRFTA0jfE5RCJpIW2SXQsw7wQLj78+13zzRM1o3Y6PffrZB
j2+EWGh8/1glf+wbyCLSqeIQhbKPovg8yqS9/PIsefMSZuE/LbIjbOJMj0JitZ0Q
tUv13cye5sFos63sk8cUVFgHyUPvXugh2N6w72aJgCmvV8KpQOfCgF7Wgz9CNZQU
1IFNo3gXY/+VNqnXeTC6Z1thVp+t51o6v3hEVYphDwyVSXCKx8S3+emLiUEXhjsu
PnBN6VXkiIijGWmbCDIJamrY7yMbnHZ6ASChebkHu71qEYC9um3w/9WA5fgKFDfC
XtTctE052GHAc0BrMbuQIw7GcGjAvhBzF47Ff5uKsqlxLKzglvh+NtJKeA2Erm+T
/knmboxHcHZcRrwr4VTr8uZGuKkkSeuXEUuNq4S7opRqUJSjFNSwtvM03ldITAln
+JzdkkiUK11ala3hmGSqtkQ0YNv3Dt1URpJ0Xb4xjGoHB+B5/oZkm7Bgf+wXmxCM
+Q4cFDeL78CL2CtdjGEYi7fPs+hOSRyCKpseCb6YuXZQGGp2DNzOcrsILypLEPPa
DwAUi3fVgdDCmbSuWcdchDES5XOGuhstIIMbEA1BxJ2hw9OTowCqJ/crVhwzqosf
ZsMKhAv4taS/F2pW7dI3VCN+S7ePVXxUEcJ50nQLbUZu+VTWRmovOUQ7niuj9WCR
XrW2LsPMg6+pblWvgfkWCVSZklF7z91nrVRnM2B5jQ+p2uvfDTVPx07C4jIiP8kV
njwUcUTo8NRKVDC9r3upvZEKPo1I6rhAwWMbv+TR5zDs7T1GveOG99a1Qz7aCowG
yf/focDXkFxD3GuUxxAtf+f1TkGg5IkUBpEfqMSipmbDcPSrHJHltJ8HK+wFn5Ki
bWRs4LRRDs89XwWGMuevNUXLa6e2r2lPeOxRmqvOJSJOTICTbF4Io/ZWFFLrmf5X
gptd82pRt6yUPtpCZ4ms2NKMv/svwTCBYY7lJHBpv+FJRucu7QMqI03mwev68Shn
nmNhTpz2bQVeF75iBgiO7vLquu71TN8VdRzo3xKqbu0PMdNpJHlVJx586an14Qcc
F1cYUS9ayxdM04djWOZ20Co3HC5elmrgiIMDb3IccK1kpkNkBNOPdsEWEF9HB83c
MXD6KP0O9sQWeWZyWIVEEZWRvlqxLsKhcqtOHQAVdN21Gh2Kpc/mPs6YSkfqzVrd
cvyTFLVmwajYAqiQW8mqLaNlvdRzZ8lwXwExVCJBoeClogx/sIHcWgcv12p9Mqm3
n/4v+1QfUFDhVTTsHtNhg7DNbJeuqv5z1fDJAnKxaUTMqQ+M6O/I/wSr2wqGR9if
DrZDP6l/2JiyUAZeyglUYz+k2rKTAC6n8QMJdHPUn5Y1l9ZiEuaWdH2zpK64m7cJ
hwy1kDrytM0xVnD3GXKXmiYz6qnNHnlautriXLa7K9JF/tj7MG4VNfT0JPUVx/vH
Eyg9mBjysTFCh9qIeZ3nwJwbVOZiggzOLGX9WXB6dyMnwC4IRcrg5BqlAHrhYzt6
ABWZTmQFNHUOBGLyeH2YpmRcDgCltDF5BaQ9iK2GsyxqLIG7bi7VEypjxHykU05U
I7A8dgV2lzLL3URVeozOi8drJr2tdBF6IF1ml0Fqw44KXFBnxTfbWJRP/VMIgTv+
xR+gs4VxDMWG9kyPS/PlpIiyqhK4/6xzWKOTD8CLT6oXBGDyO4mf9htG1lOeaY7Q
rz5aMZ43zNvu1tOqNixrabb/jr8PzJcD5jFJXMuQEZtQ57oSHCyMvfqAI+v3R2Ty
8S4JwlL36lhwl9W0+Whr+N8sSl1dXaA7RQ3Doyr0dVqG6s6UC9AUStsa+uhl6HMh
qqDS1YDV45/QM2PkDL9qd0edsO6wpLkRL6hb6eBXHRiiatnhZbJ93xd+IKLViuM4
C85fcJgsJhJEM1ngeUcGkxAfqM7JxcZCGIS7VzWbspH2R7mgqIXUslcMjkIjOPh7
fuoAjuvcFM21V7WfCBK9RVMjsU338Efo1NGuOfYq2R+OSjj3eaNsEoNd8q09CMWZ
NPfWmXO7Ci8b8S0W4bVVpztXJ6t77BvxJe1ijGGtDnsdFnBqXKj156NOKPkWonfe
kc+LlJhazkVsct7drttjOqxuhXmTa/W4dD1Sw0fKK8d2lFwuHYkNFksAEBNKHkPD
57nulDQdsL0z8nkw1rgd96zGdQq0IsEJ/sjZReNSQ6J/XzcIYXh1H6PKF5HAc7BT
Ub7s1uZ9ZRN4xhJiiRA+RgD7/bdRcoxIr6SCT4TRHJAFca9YgYB8LppU43kngboI
+bqhjk599T8skezkcITbxqG2FWF1o8ncXyx3/w9i8b2BbbUyf9UDihILna2LD5Hk
87L/7e5knPMQx4QyYutFuV1PfQYdwwgJAgYOWOyxKKrLTVd8NTkIBjgQNE5iC7VU
Xdwomx/UKzmS1SrylMfZtZm2V4RD3o1A+hfzpfHsDlL8ojvAMc9ksb83wA0ff+Bo
ujTn/q8VrvCTXNnCFlDq6K8CWe//KkK/DkYPBgOFB2nfqcoYKncMCmmKkJHqbGHr
dnbOxzjXkZ4k0E8ZEPg+Al1ROScsYXmCkKSh+GZqmhvVK6fsRbFpUksMjce7AjfP
to/xaYc+z8FtzGmKqvt+1MRGqtCc+VqvDtsKXOkk7luzcDc2QJ6rHfbR9otJtkf/
cIME/JLRvo/QEbeupdf7w/nfHWkBxX5DJe7holyRrw9l3/JM8buB0hO2oiv99b7I
xwl6dESnYiZlqpbsaIz/5Dte0kNHtfTSQDKJ3YSpLl6nV2Uynd6nfnMVh+PIADx0
LWRn1lpymcWNPPHW/ZV8+q1Rr8lsXuE/hjhcg5D/ElDplUo/J1plxFKqUgQsw2uo
dk5HZAkT2FXPTzUvGGYodqcKGA2FZPYTWMfolk2IWY53pl7ObqvreRYojvfHo8s5
Q4sl94FeZuqpOiKs2eGquoKMxNPGMISxBaJdJvD3ZXTjsNdE/QPxnjx5Qdk0fnXv
LwSYSCXJjIhWm4s1+EifU4qNIx6pbTzss1YBTlceXSo52W1FVwvoM0hZ8+xuOKkN
XFj9JRaBIaO2bAxXDQIWHZH43TLqM28ba4iqqmQH3NrsRI7NywLukke5jEoXElzS
+EksWTJu/NTSyl0Uy3gMxIzTKvuVucsoGRLcg57IsZOKKU7M7kgujQ1m/QCEiHFU
OTbIYQOcSA4sPgzU4I/z8JoosHZS1qhlXW7Qcw41kR2REyhbaJIsflqWEiiGBU8B
RwyiRwvPTKmop932XHoWnEOH1Wxcyg0NEFRgY4ryOdjTiF32XMONvBZS4/ZS0nps
Ab0xliwgw3419gLPsMKc/WzyM1n5OGpehTLkqy65jBtxcZnTIgt4PgMgryIBJzHn
WnQJE4GS6stCv5G1J5kK3s8GRKlXaKpp65AXL3ie4mM+3VJVXHTEuD+l3AVBZUER
kEsbV+9/UOIsa/YNLqI+UaV1RnqRnHSTuGr+06RwkeLpSTDs/D+/wzrjcplmMgwK
1V4hZRTy74Go5cDNcXY1r9znEvHAgXOzK4vG74JGP8LxnRc+LBsbByIgQ3TaF/pX
L77HmjHU9vkeBJDIJ3QmKF6NdtRPLo/TEEGj5IV8qp359qchU4fSU7A/irBg5dW/
SzsZENJ6hBMBYxUPnTgyiNmXKQ6S/VLRBGvFtytzOgf+m9k4sL2/lH/7PSGX7w0X
2ZYt9DD1vGQuuqCBc3jZFmiyXMqwIXkqahhUx1CAnv+5UQj3Wnw+N56vcC1QqY91
US5xRq9hlgieEY7fnvW1nx7gsk9NclFT1A7bPwN/y/X+xtO1Osi62ibJSkgRVu2L
EwOYrndS9DZr7ROmE1mGLo7rXIcdhY03MIx1j7SjsM6iSwFMgTWDH8evNl1UIFyo
Z8ieMzK2jVYFAibce+CbF/VNYsKs8dMgtqV29i0BLUsG1/pcNhSKDqz0kEi5mLzK
MjQllbNFpSLfLpHwOQobNUMa5YxvFY6SkA3viHzUAC3hF9eXGcRjkTGZf30ujIHx
yE8EtQ62X+mndzm83TtetWtIEod9LJPCZrGimrV186ab2DtnnS61SUr7O0dezI1/
+YFowOyyQFVxQ2DYA/XQruA8Sv0lJtV2uF6bhmJ8GmSYQrs+dwlpBrQ0XcHbrLmH
wQC/ZUaHA6XIrPhoXWHhMXmU4DzGcyU+iKuWW5Q9vW+5isbu3bNhY53OeUJ9q/Dq
j0YuVpJfnUJDRO2peo+u2Fp97UGQ3AArt5eg6l1KF9Bs16vU4naNAQSM0ZwOpSv2
t2x8kNjeBZlL2NS450k51ivEEC6i6IDKMoVd50lyKTfCuCNOoeAJIfR5tNcA1+gS
rnrsG4D5Bcft1O8lFT5hASYX7G3091tkwpEtVMCM4Xb7tdJx3Wb5tKZQvwEoakNv
uWNjqAjZLOvqwZtYvfKSmaAlphtA9qCV7e5dfe95LvRL3ITCCISsixNzZEbpTU2l
vzBh4khQh1qGC4WRjnO4cjkdJSQoJZOK4e1x5bWAPUCG+YrQwMHuQuIBXga59Trt
u3b+ZnfbSV9PxSRZ6zDhpaAoK65HZqECAYBqqvLm9WSSNHhQ360xLfx6PxVbxOGC
bQRI/N4JDvi1InwokjfWQoyqnijSAtFAmB0ISNaSQvfvMMj+y5WM/Pc5VWGqs+P5
GzcKrw4oWCdca3KFGqzatwqfrDTyAWW5p9qnG8pSu7MS0e9YXLq1HUawuEEzZJiC
S9AITwMBKgbVY3679+uJgtXoDF9JV6JrTtUSfps9VlgKheX1fuI0PMuco9VtmF+X
l9Mgni/hAT4YNidwMCLvxXqXNx9916MAv8YcgnXebf1FBlLtB0HahbJisiux+1CW
9sDnP++UiAfiZ4bvosSW67ugRUZAtHmOft99PNh+Y2XBy7uX8aftT1imTYhRFkHS
wxsX+Dm845dNK7x7/vPDMQem4/KE5flSPjKQ/Iy1RfwYWR7HI2zxmwPbrBidhyiA
kxkELhXH7CUJq1coJT/nzKdIuxaOR8Eq4poK9QxZT3SGvZfRXIr78LbvhTPQvIML
jlbAlq0GIKkAfYxwtdZd2e/NomX84a8RoCj0VCNPjNSeh7AOLeIx835nC4SvDgSU
ripkSsr5P8Kuik61d9y5aYDLQBdUJaCY56VJCkXGQXQG5KjSSD8rqG7DJd4jodl5
l9BRG+emla98VKBSCGsgNaC4fTax747wfojCP8ihVEEEQ5aCGH00YL6n41dh5QJo
wdJoTKZ/y/YItOv6S40YJ3GRVXwbmykUZaFV8EAy0ltF1mPl3RGhsG2Z0YaIJqMU
nQCkCcb+NGjbYtLZrJbng17rVLhgsNFojTJQBXniAVy8kb1iyzSz0aKJmdRkT2NX
q+dnw+X6Wt0YIRPGp5EJ+8PaSgBav3ifM7eebKTKcvTLrKqv3zi+iFg/cDZDlsrj
yAPhkvpAPDQLCPNJLy+DmnpqUbeCNeAEWBRKP+AveWx/Q5jS7MlGJz0QxNm7mq3n
mohmeZauIOu2MMrLVxdhaYD1ED4f8/D8hc2rc3yxX8BWRvfTefuNxHy4v4wNhlIB
xARuT5O8PtIFKG9J61fder3XoI+4bTpiSWu3yVeZsKl4K/FEV2SJoTJUR81F8uYe
Lt+gDSCRW8Lrjg/1OAoe3NVJATSawoAZa6dbexeYwxc+MH51c2NcKeppKvnal0YO
Sbd/LPstJgT28AMd+VxXcVdpcVcCHGNGPIlHMBrSNifNWUxE9UXT/bcQ1LPuta9B
NOGwCDSxazC2nESR1tCZe0bVy07azaG7tuKlCKaTyQtn8A6HFvgvWNq0Ozm6XsTY
rfMmpZhQ1hGEZSd/Z1FfxjFCjJgd7Da8Id8tknwzi7HaDAuBn6wLfDKo7md1te2j
7Zkwl7b9hzUj1e0BSf9Ep+nz0507MbRQQDBQbQ0sPPTQ9lYhfkRW4B/T4jMpdnm3
yzlVJVQVlMnISj95yG3EotdSIClYdv84szST7GfgqjNy6iyiL7Pf6O0kyATkeLmw
pCDRYRoDrHuUywsCSGwB0P7bwNlp98RHyDCRJLZGU8+Iei4SFasdRtoKMqbwtXGT
paCB+NbLzHdBZ1MUMbHCfT2lpP3ko0tb2QbK4dvghJBCFXGJIvdmIt1/m4iG1sye
5HMP5LqhmztI2lBr3rkztq+Hx9xvWKyAuevYprWN8x84dUfr8nXNv8C2bXml+q5r
chntPMLDPz5lok4ca5yyeqelY2h9IdLji5tPNu1XxtUMWKP8xbeAk6K1sms/gTdO
56j4sDbKmQbVUCF2zitM/IxhE5EMHOnmDTQb6dLAJAr8ApJnu5qF2m00/zqwH7R5
uLlSthB9fCokEYxkyPRex+UqMbszuhoObH3eLVehQFNv5cw6vRDd8QDelesMY+2P
uQsMfvRQIA2uU3fBeLHizjPvBPO5hqjZCpH11Y3dIDpUrCDMyuuWiedOj78BQRJX
Wn+8iNmi7vD8TExyiu3gqVveamd5+YCMWtAjqWNZP/VCaBdoUvC1ANquKjMUPuOt
EKKcvBzzMSyMR9ABmGe7rJIMBlzArrHh4NFYf5z78OC8eCXaLKjzkBjFj4FSCG4z
GNymyLHfZ1avaLQlJ4IFHWJl0v1il2foWipoHDfTsex/G7n6t+98ce/tnufXEMcu
p3UGIE/lcDW+i9znArbzxLOLUQJzwOKdwL6OK927pdzaWjZQbX0rLihfwqosBtDl
jl5nMtNMlih5270u05w6PSiDSfBoEMuko2kdJs0izf2BBOgoNfnSELqJbk2ghZ+Z
fUTAzL62rG/ShGBXjxUXeiLnKAup5asZ5IA8lpA9USJzS7ixycAF3B1iT/4ysOyP
Prr+RTfOTSZs3XLabVe+zWoo0mtZLnGFRmCO697fHJArtDHuMVctPJAOSwsusCfV
cAr/N0nFIw1okFgWXNPlYDVyzreta7ij7WA/AuTgJFxmIcieG+YUVXpfdEqa1S2t
k+fPafCRzill3yUL1rl97z4G3A3r+djRbg5fiOczr1wu22bw5vjkS80ri8YicJLJ
Mf+kyyo5OXhBXgS4tFDnNNvAV66+Xwte6YBPAo8nxvJ4GpE4yceCZeGo+0ern1Tr
87L740LR9L3irX+LjfEI5iBtu59ld/1Z4THtWupp1fQQp2EkWT2jOWy5GTrvakAH
rk2WgBxL4AdyTioGkQ3+WyraZrjRmKPJQ5aqJ8HCSX+AwM1DRXm/9j9RfifzmYrd
u245Dv5cL6LvOaAeFDyqwPljsyx0WtOGYqEB68tqs7uPKriuLjE9TqlVS7yuJn9E
v0AQuNNYir+xU6Oz+x+A58B491XZ+Y7lAh9Pi/LuAdir3/M15RNN0eJsriQRvhpX
jLtqSt82sN1VoCz8zRlPk9SAoSMxET1Hh95X4Mx1NMGs4anaky9E/NvPMzK+ZjIF
0lKCg/AJ/RyFvWoeQ9t0AUWWKG0CIFckisFnbIhEAGj+xI2g91drX/u6YtrUNCms
c3PhQH95dJbeCr4mFA/Zxg1A9dJDQJdEPLimEDOiBC+LZm8k+1o3F+sDWU5FABl+
9JWa0jiUWn42xV5eh8+U64HGlHVSTXM5idNF0kdevtmbDfjDxOZMiuVt5k4qscYD
abc1pF0tXhKdB0RvFtFmdOjUjV7+fkwGMTOEfkDUkoMgI27CUYXk8DcLQPxVrIbC
5nTQNgcynzNozmZlW1zPhdb8NTOXjuy0bbV7Y34nU4b3mrXUupzEkX5blf18u9CX
p4UM35I9N/MpvFbCqBsUF6RaEp+kmoZ0PshV1QNdyZrd7t0nExpnND6X8OkAS55o
nEnpcU1/VFKgMFZkmTMwo1JsC5dTPoh8j0RKYJRdkETAq7cJLS5R7HIWyzQeFbUl
eh/kzIlsH/5WdFMUdTle9ueaxDXqOke2i31cpbq8IkuUgXFlCGoEKER4f59mot+6
vS8Sz0pxOK3Ivo7leXV+hmy/wDJY2B8Da7fBoBwXyDmQeVBB/7lAPr7TS8jT9/pB
2naAG2cuE002kvV4WgbMGEDp9N+IBI31k1CE0mr+Yjko++73aICDu5fdzs1IJvtG
UcoGTfEqwVUuOmhZ0H7ZDkOJSI2/2pt6C7XhaGcE0zNAOjOFgTq0SkawLIr40w2u
Dd+X/ZuAmeMqyQ4sw55pvRLTbQ3Q72Y2z3OHa/kEEoY1OjqCSdQ+WyZGt44sflVb
SYXOlWoCjZGbaes9O/KGy+IfN08aHwl/AXUAZ5arBExJj93ZkjvOQDvVcNO88AJl
O11bTnwP92T9YD15QMZbaFY2zJJHZlsD4Ua7lu5ndbzQLKL73ZnWReSPAEdo8607
F3QceOiKkCgjL2EQ57+EMczk7Lo2f0e+0RYi1pNDv6yZHBZgeGFJSbgd1sX4ymuA
BRmod8euNxoSvzKfUVdLHxMB8I5h14TA8GCRDMkPYmEU+6smKkHVw5DjzqUxGkdl
KnwIRaohlDM+TChyYvUg9/D44hFHiZBXk8TDMzBdA4FNOOdsGxUPHrLBGL5YkFkL
PmvV5iR15JJEQ/xpeRkcaw32HFoQemKHmX/V3vgFUaKX18EJpYi9EAFOfyE6sfZM
qCT18p1GrtpF+4UF5Do/yLGlLc8W8jh8S5qhmC1RzJDVnh+rvTCfZq3gT9cg3diX
Wpn8vci2dZq5SwseC1m+BiyMIbTTtx3YixJkRhpWzVGkLzxKiPE7p1P1OJcAPJzN
VcTbz/7OngdzRpUhip++1RXgvNDpx2HdyseeIOgKCsNeuknvLQAoFcME/Of+hHGG
g+oZBjDgEfZjoui16oWszeik89wTPOSqssIUd5uunpuPoDAEUU/KmszQdGqr5kVx
OhyajS/Jsp54Z0Z2eKjUSxG2t/8tGUaC/1XOkbbf6PYHJLWCwTa+PJHYxqSxgpSc
XiRpgT/3y4ElgGO5+irtC7O6t45k/pwBPMH6hfriZagMK7UXQtVVdSY4kBEtn3Fu
aXUOVE7stZQMlmpEn3oaNXS+rRnPcT/nZtKctru6tGdr9jjsboCVO8ZuQar7XpSH
U4I5n/bp0rck4Rdef7hAJx7aW5SZV1Jb3wQzt4FL0c116QW9NFEdyEBpQasjgdiN
Wv9EFBPMM6yZo4xp+kaoDcbN4jVdNuTBJ2JV2aJkvr0TCn4Z70TbCl6oaIUf8k1Q
nDpQHSBZsyueN/zppGE6U4LykO/B34r6K/QwwCtj8rNoTvBLcfk+zaLMg7WrXQIB
dhqgzdmlqcxDI0P2wSrfoCCXYueOT0w9NL9qlMG6znqt1La3QDr/5+ulGPNHBVkU
RjYFIi2vWAOWLuui18kI4GwBeVX4oegcy3qgYRk+QJVPtdiAVlUhfo8EeZkLIk2c
0qtrg+Npr/CZkhSRVfh+YZot31zuWJ5Os/0GLfOOadC/qGKgPo5to8IlRl5V+APK
rE5Jq8T8v0wdZ3gac2Q4A9cWry604rcMmFW+Xk60+A/FOMuJZubs6HMjiP1l/chL
qihiXS06i1/6BVqvk/lbuFkm76bCymNy1qtSHpUg+wXej7u0ZhBwYn8+Pc19Mxfd
GyjboVUvXKo0iODxEzzpOPURfNbemOp31t5L2TxrjWz9y1qufHtZTCC9K4B7Pk9d
siXaf6JpXTuMJVPZcUTeQZTYwweQdX2JVtKtHyRIClgXMxovAI2+2TR9zMa75ufo
Avj+JysSfL/h1VxFLv+OHO71ZBbAT/89+sDWnhxw86P2wIocUFuR9Xc26QiE/kn9
rEBdm5/l+mx7KZnsqYAxM99mYP6tkXwWdnpoJcLwHNh4w0VeyjgjzIPzV+RQMk8f
7AXtZnDMmjcpKSj2msEbXvquZqZ3vJqfcp+x9G6Mfh9/Zha8gOB1PzHgqDfbKcs8
XHjjdCryG6ZEBjnpGQvf46qmOVHi5lm4cqItVMTtNILsO+XI8TO8d3Q8WjLF3UR2
E3/gHp06NCIfOzpQjl17YejplTL0m7T2sSlTRVK+X5ZizmwOUemi4UeW/el1iOMX
sb210t4WnLEd71zCp43d/NtqKYTMod4l3+u+vUake7FDfbZ4J0c8tEMFJ3CKBtuA
XbYQw+m09JKVAqSc+aT7wA++urun9cQvW0WCAGYN576+ImL90xFas7apXvrp3JoE
TWFDTXsguULozOJXHqWVPw5OkYoWbPz7UXUil82DwlPPzDR3pe/rAUZVeXi/C6CE
aB7w1Q2/FXR/5Rj9RsJInkXLE/ijL3IC21fsGjl135dY14mZW4wWzqUfxsFHzuGF
pr9LW3jBJB3MmPxXBXbCEo3S4+ZLiRf1cEwwBWZjs7xuTzQZAYjsh7ILM/DhZ3AQ
qBC/7dMj44nQbxVUqqOiykIYPXtnNIJ0iZz5+GO4f+fabDsMUSyB0Jq36UUApLDm
IFDjmZ6lZMH/ZmMtXlWheKq4qyWKps6QE3g0OKqvFWMXSSj7YWqh9aLE5CABdhXV
pqRvOkNRbbD+tl6UlJjse9IlUznPBp2BGrUIAFwjto1DAcY+G+/V8SZxoQl12VV+
uT4+mCQio2ycT7n7gIL7L8ZE+JlAFn2LxcYh7IvWFw0+KksOxKqatt/9DrPtIEZJ
wZOXVSVMtKs9ihKn+EF2uvHYKF1b2Zlanztc0H+dJ1kqv+uoswtqLpXctZ7y4rum
sp4bQPH+c7glGURKhHZOEo0UkfN89fUmRM8nhRFruyDg8f07NGNNbIPv0bO0AZMZ
HvWYmWXflkwn2pPhEzUy32TRrjtyQ/K61CAUWlrLrYMc8tTSCL3Eac8Gib2UCroq
FyZMpR+IIhHSCdPZ7UOK7LNez1N8He66/rHI8shqIH+5PIt8ZArULkoUGvLBpNjQ
YDqkLx4HAw/IV+uFgrVMTdd6LaP2rOVvtxgO2Wnza23KtLLUkfXJuOl9gzK6Ehhy
lch5i3Lq62rtF6oVTOlPe6hCZ3b0FzhNCFRO2BinZL5vqg+J7JRjqkdFhuZMeueW
eAdqO6iT9Lz8axWkFfAcYHQxUYdTT4ywwnklkE6IUyEcwqNjGpRBvhBwHBzoUpPh
kE4J6T41FA6nyYvfiJfZDEZu31Ctd/qOoXYkKmzJUgh6wKMZ0NEPpCeR6lh412W0
7ZDfYMKVHUhTtG+Nk0iykTo75oevl8yEVUqag3Dt2G8Yz1wokAl+EhtHRrvygWcw
Ch55q7LeisD1Gq7U0NH9TSKOOOK5U7/6poO9rUHU0K1p0+8ujLP98F+hfcH9K/nw
7SA47JTQPz3BMDk7R0RRSW1Is6+vP8hF79zzrvxnZgzcavyMDBy0SsQB9Zl/sQHv
z2XCly35qhsgkfkVPvAJZaCnw3OinY8EynDGDVMdTfKG3IocPvVNKf1uI3O+xgdQ
oNZpH2I53r9HL/Tgv2NbEnRYYSsHO/fG0YcRAzTC0v3AOL431eP7EHB6RLKz10iX
hFrrKuxgT1MtgGOi10fKQ5mFjAbEya2YdbvRgy2Q1NFua+4gV0JI6VAYKOCUDoK6
QXGVMuU+CRG/eWL0scfOE0O2/m27FYRpOQQK5JmHUc9RufsnMyXMWO1XmSP7AhZh
o3853rsm+yi1GQojWxajRh5nTupdaK57U/bwcmkfgLUOxzsupwg7fb5f42/b2Cxc
uUr6yUp5/6bp9R1eG+8ie6LtyRojuN/87OqT5w1F3i5HzMG43PGb88cDayh7oOdl
mV66fgyN0dIzm7MZkD5LGcii8EqXPoa8XjtKg9ErJQnFCBjdo5/MLSCKM0bw1693
1LtfNDuMSK0YKmPihe3MRvIVwarHuc2qWZIVTdTZis1MOpLLX1M3gFWjZJlQTc+U
RAvSON4h1Mi6GbzXEA87oRl7bSCHqjlpj2UqAhGrDn88imha3D3SvSAo5MxtDvc3
nfXuaqXJ4qyIH6xL+aZD2U6FPFTfKbLr6/AXzxl6Fqu8CCAA1VTAptyCBLgX0WAP
MT164E1eR9VaAFH1lInArxVK2Fo2X/Ld5zyhGyItaHcXZifXszGBgjwn3RuBcP+0
QGWHgqwKGJzkSdJ+UphN4HYPS1QKeMN8d6fqjJsi9SdkEtMA7vUa/QAikGBugweB
AG21MMmglzHo0qKNtF3TpEbKpBL0RlnvFV0RcsEGPSgQb/dH7EPV8zXTR4r7G2by
fKZ/lMY0z5TGTJ+M7jjDDTBjm77kten06ZJ0sTpFniMmD/RiR4IUTa6BaXTYmtfM
854cW8191UxWBKSVppjJDpLEpttHP0lJ+ZH4yo9LCNMtuz9y9bqL4n1vISakhvUb
FxlHwp6qnTqS/Jf2vzULWVyITpNSQXySqD87MWRFlXa9GvJMTFFsE+cAR2jAho4P
W7Gwvj3Ufu5DMNVKIfKVNBPq5WV6pimWpN+yLiWMOj5N9b21T/6VYAL9++ISayHt
0X8yJ4D34RuuiWlPKAbdw9gWDGkz7+Q1ISZqmTvsy4+j4xGQTvAFieoziLrvSE7E
XxaL/f+GUU+96fpsLSSV5lntWwIdO0WDKyZTkwfooavxGUOt/H4lNqqODMb6iDM3
izNtgiH/k/qrivOT84O2TEG70zA9SO2So+N2aWeFHp5InRGhYCMSsY3ddRzJWjlE
OnFej8duCM1cjB2mh4kdYDTNgA4pzwnGFHMEZmEN6G0r0lGOhBI2nU5K8aSHpn6C
4uBDIvOXlGrz6M14kGA89e4l0ey4lTkvWE1pf5jiEwJ4zssL+rQpDUtnFGiW39NA
5mSOYKrDhFgLOrXLO4zTqJ1RC1krdaE5/D/PGaTlxAUo3BCn/kTsS37gEQlMwpHC
AMPfBOV+0twi2FuKtdvMMiNAft5TGWMz833ZSVlveifywCrGNkHLnDVPOPnl2GXy
g983nKcOf4T2+BMURaJ4XAjPyYoajwyTUznrkANNeya51PQyAcQx8UR6Xkir5gsB
ZnHH8+j7o1PELMtPXzjtJGFhy6Ciw0KG6pseQOc2geE4TBqwO1P5MR9BCEpU4kYu
JqRq3mnOPG4t+hnipYNrKgb4N0tbTLDZ6OFCDso3R6GkuB6lok9VZiMaPYnwiHfE
zP5Uu+DzazDo3g6p+wmuhBDJI0YJnfb4ErdqXOsu0xlH7BD2hYmda//cRDaE2s47
3VgZy5r3UWpzjih+gD5DP10QYeVs8NhdVi+abYvkmwpExL7TlWzliyGYLsatOxKy
G0VC0WHnXDw/NbHYtfwpkmQwY9Cnd55p4/imvX2iKjfHSBu/tlYdP+rz6KmtUxgc
6bNRJvAxywGLCFfSw5+EsUS21tdRENXmF8nYMqFbuEl/Em1Vwc/acSFFEFlV3Mrq
pAd7TSKUH2XTVIaNC7ZpM3Ab4NzGf0fmltggF2VYGIpuiDKOE3u5k6RSjeg6s7RL
X2a3pKhY+Vd5EqBsZUdqZ9HAkA4qgQtpVrTKEsS9yrr+NrOxmPbuH9JerJhW/cLt
aJIjO5108tMl4IJvRkYPO08Yuvksd1wlzTcVCKT5Twiiy+Kk9JxstUu6+rlIS68c
UJun3bH2PwKxaJ3jX23vSG9+4rZkBBmXUUcPj/32nUtW6PH65WEQhHlKxbm5rVRm
epzIlaOcwwJBmWkePLkn59XpBG6zHpuU7UzYBVyi79OrMo8Vc9Sf1B+AM27Mqffh
68/37vKQtQvk5dwjwVbzP+5Iw11NxLHTeR8qU7KxSQP5N2xAScjhTJj0ovtp2fen
NvpRT6vVs2x0Hzq4zsUuKKY45IQJ9Osl2HCw+Z178N5dJCQYQWWk7nUd/8ESln0Z
i3Jj8gR40UCyQ4VjXp2SUlUKL26m/nfy+2WEAU7EhwrC/yKZIWARc871gKAw2T52
Mg12vk/9sK7fqiudBz0qkSHaC1IuarFfOOrqRo5ASZnDr1F6ZMU21AxuKZamolxm
L+Db7PBO/kzD/zyi0Qx5DZbufsp8pO8l9T8PcIjaulgA11XAd1scdJ42+1PUANyn
2ZXldwwlnCGqE4AsvCiQdyl/daLj8UZyDHvmeCbER/1YRwinMmsGZkTL6fbWTwvH
z8GzXDhXS5e+EsyWIoAPYju23eUcw1z4pPmlQZ1Iz1lkI2MkJkEIXjUvLaS10R90
ByJHeWy318fb5O+jglM7K7hGhOL7OQRFcofBE3SmJYia/1oti3QQZcZpPN/iihqK
pFvn+zmDCYNFOpZaX6U+8w4qF74qkxBL/PbdxcArXKJMl3LsUyssYzCU5+yJvipg
BZUlLidk8cS0zJbS9VCgdjPUvV9n6/p10w/oVvdjIPWCmA98gGcbjP9p9ll/m1Bl
h4moVCYUdhRqecFqKS0VjlZ/3S6QwZ1fgEiUvGICVp1y9ItieZf2x4upZXakeBJD
mMgfEISMVys/OJt6KadZC31UMIDgYklfXK7MbOWIH+RyNZ16MNTHzDiHgg6f45Le
zca3wV94IliFj2IhW40gHVm/TxKk/ZRWbqYy/3rVslV+u/HdryFZkQkbA3crX/si
RKr2O2vGXcxW67efRT2OIHfvGvn5PKNNqJEGKW0BlY75VXJ216flRZrUqN0OfpcB
M6TjE2qGdP3kywuLvtjYdw32BNIwTim7tifCxhf9O321tHZtTGtGAxTWGhMEn0jW
eOZUymSPUXGjWkIcAsD9AJVG/FBZ8649Nq0yW97CDC2eG7DQSSZY/bp8NE5lBKJE
ltjm5pJUolk6lVEGBeRBNalMfdIsgOFRIz0laL1uUFoVxprHHawqywN9WsQex7Qd
1p60XO5RjTTUhMGIUKyM1LBC6BtxBhGrk1Q9xEFz5HBty3wBJu5LLPgHvw6+BNJ7
kdkSqhhNXDl16Z2kW+pWVrjlye3NYSmgWmuy6ZySRgkeXQUx4ftHmhps8KWZ9Ci4
eoVThLKWbaLmyVdbfpkNvD7e9onUfIZVc8RrpLIyPopjAaRUTVoJ8p1mMF3rt15H
B0W/ZkF+1Xu1EwO3EHEeVW1VxMxu66IyN9zLnC7O629QUv7ohu4L0nQNOKnXy9IO
gMvCeNvsjHaWbdPQpdGp7tXJ5BRAvSop8haJTNdn8CbEARtoIW0ZjoqySyQqlyir
FQJT2nNeMVMbDu6Vyjj4IaudtLNbPo+ifYJXjzd+CwrlyvBiFwiWIon6awsnc8aV
tmpYHoCOspnks1GVYRwqK8gLVLUTzWvGeFcgxZTZtxA1EbhHAf6OBSRbyb/g1a0V
k2YQJSGR8hHyr+S+fPyPZ+IsCVBrxZ+t2hOB+sjvaP8OeB40mshgsDs9ZERa4o+3
pphSzh0gSbp7sBbrmWOsTaOw+9tf9PpKT9jxu5VgMJ4ck5dof6NbcS/6tV58pUNd
sITlZfOEVNToivd5jsfEyuwD5mxJKe110myx0lFgoZVJO3cOwUiSuhnS4g4ZkzFL
oqu40+ezkkNIbPPBFf4GUpmZRGdgBjqdjF4df4bNFOEqVwZosyTwLOk6rXTCo/47
2OCroIkJA2AAfUgSjqiQf+SqZrXP7MSAoyhIA6sx94ZLayKd0pHYzCKU64J/ABB4
ytxYeqZm8lzfteRu3TlcqivQH+FEj7b+PGvMKAW9M9Qy8RXqBBOSNluyDTbGJobw
vclLeV46jgLe01rotEOx5oUcvvmHQManXNkuftbkM7eMDscRbeLZUaVR2RdVb96X
cN9p7fx16ogwM0EfZKeceT1MqMtjIbaeSw8rJJp8tZNv/y/X6nUzKmx5Ciwg6nw6
4DDF64lXMscaf3DhzvhpsC8IpqES8h7AF/VYvHiyAiVAS7P+V8mtFlP97mnCz+bD
pxTxsjRK+AtUjm0PJwX4SlgL/6UcMbVnHhDN1yIauXC13rFGZuSJuR9rapaCJ7ew
OxSrXQU7yek7durhvorFlSFny7eRSNAQsjC6G2bJwFMpxVVWOR4ut+AMSl3jiLq6
xyyirLVY0STvYV0cGbcePqoxpSc96ehA+xW0zilgwH1kuHKaTAH0S+lidwjuTpGK
O8JFhmYnsOHoLMRrGi0Cq8BCuRs0YqjPAMantBVSHfxw2uO1aRY4iAYmyX6LPbDi
qZKMq61r3FCdiMXhjJC+6aUmotNKm4zXO7r/lf0XLEgZ3Zop8rFTtZSBxqmIw0wP
BCdKzaJlvhvE1g1XPAoVG15B5uKndiJbE6xfAkaVCyhC17i3XWq6wsSJhEl38aVN
ZGSiH+U00IeRvBApkhvnozkCW56H5Sus6SWJla5EamdcOaTEVDnzP8GiU86wsNvY
4vBWganRXEyX7KDslhVgMLzhlcpk/teIiyXbuNV1QTqLmBBhx4ux81tsQlYsuGc1
sOSEU7TFrcLXRVZmMV/edDRPoMij8UQlodZYz6A977ZvzkZkWZMlmnhBooDFzBPP
CenPhG7dPCA2BaXUA3DypTC4jS+GXMOW34ipq5P6sIoylyQO/WJN7sY6vGytKpsr
8A9XyPNqP++HzMopoS8P/zhDJu/p9S7xhvNIkXliQQS4+PCDB0g6hpb6BtEyWBLP
FutOks0ixUOYSQNQpPTrvx4eOjLbFzXzhHigNb7cGrW9Yd1s4uup4C/Zs0JRZeis
sYvt+uclojXHigrgCb5q2d7Q3qubEWLlTlsHyGdiYvdUvzK/6Ee64O1y7s3ZyNQl
tkk5YoY/pk46YLKmjQD4U55L2j3XRTsJBEbmUDEjZ4et7P1xrZVnfUxeMIQH2SAO
Qj8/4WBo1Sd4ADgvKv/Q9jGoab2X27c2QnOEPmtuHrsjuQS6ReB8YMHg1C+Ut2Ct
5TPCs4IgrIXvidP08tD+hZlTJcrHPh0TY9OK8aGFAGhjqbRdvaQxQjdmVcJeTWnP
RbqztCYPuF+znjxOZpb4BVIG2UwIHhRnvaIDImJEjcTPkcf0jaX8cm4OLQm76CjY
00RkLrEbZO3DU0llOBJznP+teVih8SBpJy0ix1MISvPoqx9voYHlYvhd70Khv4c4
j8bOQl3jzX+25JX/ccLqJArsxgqmv1r+KNpn+D1G82EXVdANypoCdLz4VvuYYwEL
hEie7lQeBNC/NcS1B7Smwa1ImZOd1Du1bulsPzfTew2ZNE6wx5yJ5ssWL7cMU3UQ
ZJDIr5pC88AE5ClFhOKKUJPVgu5F4fKat2vyQRcKYuZK0RdGgjbuJmxt2vumjVM2
4IzmOq2jV1ztdVRRJhU17Ygr3ve8FfUP0MYGGC33f799KqAngkzppvCXENrDOT9c
uYri1xm3kqqeXv5tbqU/KlEt3tPYi3HJVybm32QiiHoEGNKgJ/fiDmHpAht43flf
7NhTFGH9s7yVoNkpiCalYATUVBAKRlxuj79eXij08VN1MCsEmYkYaYM4BmOKL3SC
ECa8i9G0rVTSwvu1VVfFbet8od93mUm5K5y6TTITBSOrdRs4DwmFhNggOLFzIpcm
gV3bB9i22BsSEWdWb4rzWzFyuH5LsV9dI4DzHWGNL3Qs1Q/yxplzByvknFIzvQh4
2KIK7/3/b4+pXtBJRes+fvwRnzd4Nd2yJ7PnsJFFV7h47/+MD2G7IJZZ9DJY2Jt6
Ujtg/DMHIv4ZYCgpGlrIcmZQczQZsmUSXstIDkUut6ivVqmA4dtjFDPKFPpQJlI+
XIYqY05/TtIL9vA+0ECmoQJqTDBdDwj9SKCnyP6U7HTCsjsl/dBDA6OugOsolhm2
xFW0RTvd2lhGrShSTng/0ENnI7Ldya8kFG6GKyXYDTfHsAP7hNwXp4PjXnElQ0VM
rOrQVBOVNQxqxyJ+3132cRH+JhLkNR0T4+s3OembL4FhJxsYxUopBhpC2S0kOqke
sWVBc4r4p7y/mFl4KwRO23MTKLV4aVzz8G307qQd873Y6lmcdLlfACX/isgXT3f6
U3xli5d2is3DdKZJpHOGE0YcfXPg8snXZSQ/fzXlwK3vddC0sM8NMW6mx2aHQ3QG
CcY1iFGUzGdDTh6bpUX7KxeCqy/S/+5rvZ3CqBm8hloDbjDzz9+m/gPmOt163W/L
CHxQsjoOXmbC9WRpx9b3sZEgMB8/tO3GCJc5TQmJmuwIlsp4x59EKX9SyEtP1+Gx
whDHYZ++x38ZoYhJW8SL0xv9a43PqIJWYnoaO25inBDhSGzeiLUBhUDsi8CABimg
xlG8ar4dqgd9BZnqeKLucgUF5806PXHuiDHzblqpPX7JvYvsGj9m6NGEzU5Gd/GS
AIYqU4w5TrmxcQOXBn1HrsjRNBMg2Qh+Mv6OqIub9GTGRXdcYqM+/Rj/dfy9JvEy
7HUAgGeKUTp9so03sRzNbtpygaORew1wdgPVja7EIC+6HiTqC6NFA2+hH+vngXfy
Add5nmKpE7JiPEVGCKpmNZNHhtTdp6017qXaCeA9LzexU+lEAVRyT1sGTwR9XV0z
rw5kv4cTl61/Vjza7ghHCLqdLvZsUUYOLes25S6VN581XQ8mtX2z2taI0nhHkJDP
vkZLx4OT7Ef+LxeiMk/pTWpm9fQu8EmtyR8V7+ZpHVknDMslH4rArDIswJAVuve1
t1FCnuWPOkElI0sGcSXRJHO6MzdvRkkZFO8QIuJFAc3rlihg/OBSwhIemgegGeAO
/d9Lw2zcaFBFvcvKMiVUelSz5m3fmLlXxscZMeJukX+qq+r5LFLRwGCtj3PNcHiK
AR/cJQ+nTZplPyBg5zixpnVK01J49DqE8IhlBOV9KD+2q24iBJSJAwMjK9Lex2wl
hnoGhmPVulcvPdem5mE31mP/atjJVNl/qkvXEh8NWZY4F9yf7OHZ7R+5XYVzp++2
9+KgoueJZmTNsmVI4ppSfQkevo7dkDOnw/Eud37yh2BxLodo5DsoVGLEutQaqnki
KKzEXwJ46+EesVUbNUVi1O967n/jqQKos8Ckda4PdAaXnPfY7F9NI5gKa+LZTEvB
hZ5R7Z5/XIMLcThZZz/6pbpqwfs/BXmHvYxjN4eGufq2JvjK0vm5VeITrP8eQ/ni
0psYURDtkZ5br9ZN7jOc2DSHUI7gsMnpFYNs7wCAQRwlGfbAgzUtjuMWvj+RVh/1
Y+G8ZwOWYosbpmWpEwY90xrfTZPtYZDBNuwfvnncN63bLHqxrXx9hOUOcwMV4vw9
BuNHY4PwH4YYFqXKzHvSR9Uy8U/7cjzi9TPNbfHWLGqO79lUmvmLjJk4LMR0QGYd
LKqtQaGaHAwzajWOsS8tQelvB4Fhq6T66sJNI/JIq2PTSGAHnkMby4VqwczoDdHS
ioWXdsGvooCkf59I2vZTB4daf+VRFISuPDpT3ckyVlwF4OU+u8CtQYhB9kV2VjjU
EQI/7tc4eISY8YTUkaQFaFmdPEwgqzPBtgQmc3Fk52euYz2xBUzx9pYzwcAqn4Oc
Zf3ubHbomm7jmj4ECMgf9/WEEVRIbCyMGkeiMOskwpxb3Lbf61iLmiXmQdl11uJP
oc8u11iG3dTFgDbzIGX+biJJ2mxiV1CjKjgWhu8nBkWVAfn0bUMflbcA76W4bIhZ
NM6DN9QnjZTemdB4FiZNc8thxvnFwdH1ji4eoIV7sY/mHK0ZU7ci+Y8Bf9ybC97C
zhqcBmscL79BOYOYFfenbaft3Iwd94bQQeDXVzsn4tt1ZxzoylT7h7ri8cXIvNr3
88aZh0/q6EDhHF9Uuea80rSMaWmfCllJplt/Sc0/lRxxmcPiKLgmueBjSaZu/7V5
T5NPfAg2uNGdozAYdolcWEZOMkL5bqB1z1ht6PENl4IFRpQCdYXacpURgR54jzFY
B+ES6UKiZpIlkxGuxZxfQqaS3YQk8J0OZ9PLLz91dYmQvI06GHjQjS4Q1QMnDg8R
Uggk20KJ4RkG9LTHCKvfE3JxlkcAeGsurkMotZyGoAYE/VOJXFUm4N/hAIZ92W95
jhUVv8jXK4XCsur+JuJIrMrQfDLjjMmkdbN5ZX1PtAMuutpzUhCQyGv7tj5cvxlt
qAuUpeaQr+Ig/qCINWfgmtnbr6fSWO9xW+NYGuq4sHa+lZIIIZNSFHvBgaIduLzM
9gUbflsmZkP4hgNu9T2aY92+ifU9/jna/r51upxJ/J8QhSQ2XNu8fDC3NVu+gt/A
0Zu3AtkF9cOgo6heDRSU4NwXLrNQnW6lOZ17lEMKv+vep+eubJ4RdL70Q1O1V+V4
vgZh9UaGVOzCdbZBdoFe6NEC4c87A1BKlAvmNsRg9wBeTqysdds1btkXADHOTRFD
A2MUjXo0PmQymqh9SgqgORYZ1Zv5g5TYsZj9JS+fVE/Vs0oP5iRUGC6/UOjs83rE
YIh3dZn9K44fEez4uV6HsqaoXJOdmBhXDzkPS2TH09YZIW+vD66QsJz7H65ynqjE
80+pR0lFGdpJWJU0msX0ott+uYazKFpbcw6FPPB+P7iLcP1zTnjtnwrcZag4itXZ
T04vDQx9LeFZ/lbPLk0DfRrnWrvM1HTLC67HNlhBhGydWjL1+1O83oEEyRQeVgKa
KtauSwdkKOFOMjpYb+FxiJIq1UeY3cfLo02FOGm4cxDatuaDcb6mrVJIBYkVxamu
0806rauiStV+jZeMwGdlvLG3Py///zTtwTisBSk1rzdFN5qzhay3Qi1/E/sQCMKx
Yl5KC9HGz///jmoIMRf2xfutYcuUC+qERO0bbSfg/zfIqAbuG8VdqnpaOenLvfkZ
OTSXrSdeh0IfpOh59fl2PjlUDnubl9zJDaWurFmElE/7etHKNKPuLN8Wj5mfuTHy
x6ISjsdaSItWAyxNxxlQda2kD63DsqRoQdU5TZbAE/vfu4nqgVWrf/cX2tAqaKBb
mSZfzwGC5LWwz3wkdbzoRSOwEEa3vkbFmpks9Nl+KWgq0SuFFd4s5V6fqMH3eD7d
bxx1I3I8mDxnNIh1Ov5BZ889s5Rj+xXrylrvgmCrsZo/K7neN5vAaWNr1fWy5exJ
ZSXuHI/+owLaPW01+jLpeVuJG+gwpVYDRcJ+A/26Mi0ALVZhWMnk6hO+zP43z8kg
CYGs9pnHuhq7nu7ktJzAieyKICAmwIlKeNkJ/VE0nZHmG0wmRTnGxy4dZfYCXpky
JYbZl0yf96JPcnSGmPL6IkTaxnb0NZt7qmyUXSNZcRjentYLxzhp07W3HRJJsVJv
wIn62sofupV+l89vpzvkM7o386iX65R/lDXSXyUMvYIPWmrGcrrbPqk3RgzqnCYg
EO5pkE6Gh2Y6zs9qg+jRgfqGvANha2sCGqjsv2L7XA5CzoAM6NilwUTAJVKXzE32
thWuL9fSCesxFBoFIdU9eTBofEG/F1Irwb8PxNSeqALv0GBTS9hNj3huBOilHKP4
BnCHThJge4SFjaq+vPVKkXFWlZw8dwhc5494lYPkB32/8X5QsGCTBamhjRwHs3Mn
YIHQzySyNQNmYrb/SUAMZuPbPToeT5DhPD0CDV20ZfGHedcEx2T7yVsd3L5CilgO
mYI5/6xnd/6vSoMgxee2nLdPyUwt0cPmwxw5y4RZAxwHvbqgubvQFmQCRSovrVSi
MZkW1gmjxs0TcBpTbVr6skGBIKnnYZ98cAEwGDvaPPftTXB6x43tVaSBtsFcctK5
5bwlTxhgS1VTzu8YcCyWo9jx757SVu/IUrBzdxnFJREfdqEd3FvkGPNtUfx+siB/
Nw0XBp316PsWmLb/N3VQZHPiqiFf5nwL6hpvCHAxX0G+habo0ZhiKivdeQtlbtLM
HDbg0yAagtj2WlnORxH/+RiQD6g2UdkblNJS+wu3QLqtX5LCaowSJKoFqBGFHKOo
HPSVKYVtBQoywg5nvPMYSDH5OuvGNu4C7PCCNxE9IKEAgm1p58anaXzozHOka7NY
wrbPbBHsmo7G+s4Pcck2kMk8Q28OV2y/h5n1waxtzRvhF+MnmHZxVnXJqX4T0j4x
H1xTESTN8qV4JdWTtwYo18Vd6rJ4/q+VXjVdAFPUbu3EgSdlwGIkHR5fko9LIwXt
Dfc5pQJyscP1SETEeBBSIOVnHSGOUn9PPUHB8Nz7lnwXP2xAAGRPC0r/i8budfha
cfL7onXwC/+HdaGEOL1V3K5F5DJB1XlJjo0S+rQ4ti+ru66AyoWY+ooEFcNM9IOP
UjnVuxbFCiKdSMvsGwa9RlYH5vZspb/ahF7SW68UC8gcSXCfZqoeNj0q5ykCszeN
LQwDd4H256D+Aqu3KbQ/ioSzAcpmLU8VfxRmLkXLaBnca7uEroRUctTiatf2YpCV
GMcnT26Gx5bAIt+ZyHfiOxiKp2QTZvbrF7KW86+A4qtgfQvVJXGuFqDV7TvO8Nwc
YzqN6OGn70SfynjFMeoZmDOf/HuuBy1fD8TX85lsv7SghKK19QlmMI81EjJVZHh3
9D6le3DlxTw8q7SV+url98goIhrk0CRK2K9oWGijIox5LCJiY/T2SyXXawIRsUqa
yweSN4iUC4I8nU9Z5K3In1N0kjGz5K/7VAYUynw2agQhKq4IewTd6oK72Vil86hT
9maK4Zauoc37Vzh/NaXSKqf4ZnNW+MTeRb3EPpo1j5xkdLdBFOqExGVQsh6i4LSk
mTBdjBVXNHnVf5pzUil90J1WRAegWy2weK29PAeyZKi1dQc+GiZiK3BamYzrTIn7
U7SVBWYcLIeMFE8heJOhzbUnWp4fpeYzOzpbRZVAmkaNfMGAlOY0jiyoLFoTnT4I
RmLa063xV1LBTv++2AdyL8ThU4pL+j28nK24nwtftCToOu42cj+cKltNETY68F2W
lMwltV586LHnI33RJ9URTj9q0ZQaOfD1VNlOIu52YPy8MSH/UFMgwN4PHsIa3PDV
Tn3kULTbkqqOnVO6/BOqSJslO2T2nOMFn3TCW+3o7mymT3aXSaVYjEfn6U0PNjEd
fnwm3Y6aDoMcziPJwWMFqrwXR7Dyo86/E18Qgp13WV42KiHQLBYj5NMVWHwyWST6
q6Z+2Kdlo0KvsSnxNTbsqlqiH0EvKk0hbvsX+N09T9XRzS/Yc21xrP68ZjonEJEM
L2kV4rHbow6z9y8omwdp5GuUX6IlcihqeDF63ep+FAzf+ZdkLD38QkPQfFtJFWbE
6sCcCMdIpO20u2/LUrBKDTpia8jWKxn5gDvNjxJLsu3Y16OnPspr2N901YCFjQGQ
v+5Kq9BuX5yH2jjeT21umgBcaUzIRU6GGS2WeeXrDlVJie/DjER8J1lQkPemtvdz
h5VieoKkulCuVPuZSc/23bmyPAN/fpzmm2UGiUbciIlxU6y6SCOiEHtCRtvO9t8h
RvgyqaAD2UPOb2PjswAL+xMgo6ZoXJqtM2YkDzYgUB0Kl2UKOeabXuYcIoZSzBwq
+dzGySn6mOgN+BaauJiTLHESMlYDCd1cPhK5PF9pa78KqmHUpo+8pBRzcRsbsIMY
ZA4Bf/9HeLWNzFlqJNjpc04Fm/fS3fBtx3EQ857AzxViv1gSKnIWyXnqxw0Ib4Ho
TTrE5xXSRI2UKOnTRNlWD2BBmO/HSFoq7jOl8m/zIcFBkoVJ8e0sm9mmxpvMa0D6
QhQ9tBS0QN2BjGzWJtuRtuAY4ztMJ2G6ndYYzvvui36R+lobadGZPiyWsvPWMPMN
Jo7YZxhiW1j/Cl1vlmZ6DPVHx+PqsEFY7Tja1oio3EKVCoKXbdshbcVqCNsH2ZFO
19VdFkTZGL04cL6ABUz60nmMl3GPIKZQ2Il1+TbLtwUA76fb7Y/BOXHYzjQm0hnz
TOJyN4Na3xA2uZMVleGbQ19tpuETlzsgeA+14/ECJFGnZi2MiW/s+ujat9YPY5/H
hIcfnmEfLQchhTxQne34B9S1dGdh2ysH9jzdfPY5GYYxIFJ4eRArsphjtg/lAVNl
vfyq3URLUsJxMXcuV5FHf9D31OmkJkH9V383RMPJhi2y+2Hrkx3weRqIqCZskiPj
R/m+HYsGSnRqP0IYqMsYIMgF2p8pXjt9HXJpeZa9WE/wo6LVvelZD/86Lp5ljD3A
J3R9pfCnNRaadkblef1yaorlZEZNcMhVkgVWxCSa1ccbzaUBkdzTXCm/RWptc/ub
Pa0r29gDcSflrdXOntaMe0UCx1pcOA9BDv1NTV9KTry4DpTZHy28a94jnGO7AKQ+
JiLOJNrZXQnjdGDdV+j4/C3xazEQX1edQoK0mh6+RX28kSZvzBOi4H4fYCOgeKLN
+CB5t0SfTwsL/tL49a/mUvYC1+tyHg/LCCiRnlqYmZmL2ryoGzu+VEu1htWIbXe/
Is2KLSl9NfC9TamUZ+4l0kcJcisE/ixLXEElAwErbPWyywP0uoR6UWp/sKVv/jwu
OparcgJqKtbnXZZ4s9IJJ6fc+kcBSOF/sONMjqgzPCf/6SN1QeZwGI0Fxjdfr7Sj
RsGrU3F+Ixz6DtBQu9UQgSQH+h2u4Sli0UJ9Fxfpi9Xz7dIRmXSBBsiDNJpmcvh6
3toUAgLPtrgF5zdlXbSOrdrnn/5wiM36TUd7cfp0BZiJNsXSv3COiVBbTwDyv6C8
fkW/wkbyhVKJrJtB2a6ngNxUTUAkh6vkabI5wl2a4W8JURd0XfOWNIpVMgyC4tVx
RKcRYpLyUgqY2c/N6y3LvermedBpMhJZR8RKC8dCCubU2XgjBdYAYQvcpciq2M3l
Zc9dDL1P2+uj+SXyv8s+/DEuTQ+QdD6qhn4j4jTjulHwCuvkKJbYu8gELYCXtGE8
XaQNG539zaTmKws0uUBTlp6J5vE7VC4l2uaZSSDGe6NQ4ZwE5pYXGDVf3jfU0XLq
YJurTuSePmPo5GMtEc/XMAX3kHWh967tEmyB2EdwirSoq/I2eTg/VMyErkwVRm3x
1ZPoat7LxC4Q8kKsOMcCuulLey4Mzh03LhGPX+Mtx1Ti1nOfYg6E/y9FZfST6Gmj
4z6RJ2b68ijoMyrHtnNkVKGibXkWfLxhSVqOaMO4dOcbIiqHieqZ4MTOuMYd9R5u
byEs7CrCVtyOphVj4YYfgW2YKsrfWABmK5+y67q+fsPWplQuI1OU1JITxaf9Ho1p
Stmjh42SUwFMH94EQv1d9PYZi+zX4/6+m46ll8RNm9TKQhMv2ydymtR3VA/Cofo5
Z1lPD1M9k3/QFHluuiVEOzsZ4JUryw8Ensg+JcIXyyLbrhwj8zQI1nCKVMuJEDxN
0T0vIOzMrtJBosgDR04YukyfBXZhqogjPjL/K8vUzhVeDQzbQlh/qz6JNgh0ubVS
hqsbeOHQpNYqGe4L2nMmqkupq6V0WukyT1BLAfBZljWc25FNc/Tp7kleYcmhB7NJ
b7pXuZYpOTzN4hxDX2hnZ419beGts5oiKx/ttZYYv20KPQ38vC8ZgMLoS9cxK7w0
rLEvw+vGM7NIaO+R4f5Jfq9EP7Dpk8vS0/1F6LHDvtfk+i8aA5OMza/gu0q3Z4W7
vQCRQ0dt9v+f7WFKEVFsJdvuCQ27dfckcq7euyIpqi8hATFfhQFUugwBi0M+5/+S
gYESG1BY4r+eboQIARPVyS+XvH9O2SwYrV4L6cdDp2Yq0DN3GlmZ5D9KLo7+KUi6
UbCZWvCiMJIiEF1Uy8ylfdZTJ+GcHoOB+btiy9P0G2FORZOfNyO8S0wNsAFkqLLz
+0M6OSY6r5AwOZC5IhWBwDudzuFnXImyIqKnQTbYlcbdG4A3qPfNs+12IhNcPGe1
q4EjzN1fDrtW1yCZMnACA0yyRQE1MdqJWXISK7Sua0O4xzIhilPpttH1cqI8/g5i
sViZ40reIICDlAe8w9WE7Thfzvo5E+Ee/VMOiYr0ghk4LH+WPgf0FWzM2pWfo1Um
lG9FP8OoOYM3KdJ++ojguLmXaMk2T9qt3c342/pomTaAJnl/o0SMOqXlwXrOCZ11
WlIA9fvrcVnhf0KpmKz53gC7w/hwh85GkK3g1XMXZ2YcFjrVzGAudgdGNnHFVkVK
AJYaFbR2Ak3Eb6FTccbR9s2+R+W7u8avu/hpmCbPzo1TJRiwVxDoqEx0ggFzky9O
mAxOJtA+wWXdfApJk0I8Sg+XaxDvOfj03Hrpbuv5XQ4GjJzUzwgO7ulsD8Urdl23
Vmdg+8d5EjeE8fflhNDjQdfk/lUPGlEqqJyJlfQBK9taHBtn8cIr6ThT9LVClmpi
PtpWEoiEhnQVEXEAHLCKwUxqgyoOuvA1bQAMNxfw3OcTYNnw5uQf8x0VBTqYff1z
AaglYsteeua0OpdxMfV8szZJ/iQNIgoKXSKT8/XVgAdoSU1g1gBQpguAnrJSXaO8
7cbvm2OXmD/+uV6xPTRQVR2cr/PPcBRp2JIEO1llNMzPca/CnD5yIdDygQGPeu6V
hsa3O2dyNgGsb1l7snz3CWIOOC4pgsBXmGil5Togbbls+vvJASln3rXXeMWwR0nr
FWAUjIbEEuo1YifqwoemhK4zQfQpCf5tw1EcdAcrD335ff8KJ5ZKc39blzdNJbBj
67gvneKQDC1FDFOb91usB2A0JNikED7Iip7AfqhoNCQjWrTLhfSXzTTLTZ5O77yf
vStGPJXRSTfJacfL33ZYxaIYw3okH58jgeiUcF8vMfKzKIuYQLYFV5AIWhtVIZ+y
FxBe+0KulezwhvuJAk1InCcep6kRuyjfDpm+TMiL/qAmq84AOeYVxGDcckU4/RjD
jCJFHvjaCvQmjveGqjMk+eGs6uTS0XM8IRY9MsrXUId/7qlTxzdQPqHAmORCslax
W7Do/YLkXOew85/pk5oVMNQAmiiM9ats308WQUJdlogTQF7QsN56P/5DkTpbiHi7
SO862oet4lfYtpTqz0DoOQ2veWpRDNkCe4I1F59wruzyW1P0dW7iq/16YM6lzRka
RrEp3g/0Azu1hYMwR8VTbu0ZSR1TwK/R9O60NMzXInhdbYcRBvDreTJYk6xfpRb4
QlNisRMkFV2f5IE+sbP5zYYMZiAt0UI9RJr2WCBcSG0rICZ4q4pBIia5KeAH0+gy
lFFvyHGxBpfL+HG3d0B2X/YzBBuVZtd5SoZXFT10N/Hdk2oZ+RU0hYc5jPPwARKN
e5WtkvyBdEnbYl1d9QjYlkO5z4u7UKMd34mbtj454l3hrS6+uGdNHRwZe9oB5eIJ
rd6wWjHrsboweWunvHg2Mwm7Ngvf8UJaK08GG2AQ3ALwltPYMCdfhntaXhESAmaL
FgqP2e2HLrYNcEfql2yd/A4L8bETtkfGb0JghrwJX+KeVHooUzGqcui5xW8XF0HR
95xgth8xzqhKvzwbbNOz+QtP5m2aOkNzBEEE5K1+uBFYBWFaphrMtg9s+sGrXyet
tIHdFmIV2s3CsVQDZxydEcdCal5y6wxcVNDL7me2Jvy2m2Yuzi0OEddFEzMpCz4Z
66taBXs/gx8+WSADqkMRzwNMtzNAjWRBTZH6sEztDT89l527tGYdhOHfwDbrBNfg
4nMt/QJtmgFt9rPlNxg7luQk69jdTvRtAi8szU95mRHZOxmhV/+KiAoCWsmntzV8
maRg+1vlAjJypUPqIW5hpxyLYFC/1hQ1hdApqxDFymtRkD0mPL8VxC58UUHkx7TH
bSDhDXNGNw2ddaPrMtcBdGeiQaUPKtfabIOK4v4vLdsYNDaUa+YZ4HHkNRvre/57
vp19bodwxBXxsPm4d1BOLQlVIc3Tqek3ae4hHJnNBIg6tAs6FFJE7DRMK3ciy86D
J7IslyMfv3Fx6czNv8ULoZgJVMIq1QggM2eKVD11Ut7RxAghmiDMuvddjsHvUGt4
ujTZzByYHp0WMD/u+WfNnAZHg7Ufd3shhqEsQm2Mq3wnVJASIwOVlAFpIXQsbhHx
vclcmCevdqdkEYU0A7h4TDPaFyltxrK7KUvc8A9Xrm70IG4/TlvtXSW6Bt3wfa8X
hf4jW8r6f3vpf0PMdIkJrBvXP06tPWA1QOT84kaZI3CJ8jiCTXXjq7j7CdlPzT1r
OKSPGdhmqYMPJnWnizGW0nsTq28eXL1eqzcJYRghXskjEaGbktVCVRUs+ROH4eMv
zqqWgYlaac6DhkrNasYgeiY47NLH1U95wPUOtBmEq2dLlvi0zc+7EluPDTERtIt4
w0fO7m/1Tq36+RJgmBvqNFaW1Rfdy09XXqEJbWSHBWJj8AOYMYKEzYd1o/R9r/LL
u6dGA8oFpyvpndJU2Bp+KvSo4Va80LjDkKNMBBL5SSefUkNSeXPeOj2SWrfH+w5x
3oNTg7kt1O7LRpLelwWygiJ3UDFKOZlPStXacGFUZzXDNCy2gEO5nVSUM/s69rS2
18k1q9ZQpCqvpuyK9Ka4SrKc9ZJJRu7rkVMsxTYY5H8L87kaDJ2QgSN8SVNH5Nou
8IzRMIhL2ub8xhmWiYI5N+D1iuIaZCvsY8sx9/STUsr7K6WBl0TD2BSpFMkhKpK2
3ajIU3ammtye4/YlJ4OURaNonJjnfwwxtLbVzKZDkGHU7yHIT7qiFhocTX0FT6NX
MptfdixUk9lCzZlSNFUlLMHPDsxCaZWtQZGEGFxHV7ur8Y8nhtcAFp33Bukx2SxJ
oG7uIY+aWbZLrI+8JHc7H48XVq3ne1RcGKTEne3fOmZNxCZeVwfJOsFj4A+oqCzv
zKBFfmVz+JKYtqYOUJHoK/HlaDlcoIqgSq9DRvNbNuS7xFu1JhMkU1tMrcMYFqmP
/wXkQyr09E81B4X+K9sDah9bkxyrL9C1ZIJag9Oomb+4vIrk6TWxmmVGRcYECwkG
DGYOan9Xlscko5V6mF9w/hogtf5sW6nA16YgpV+Y+j7fWoL7yPi+l0TjeGkhz2ak
LAWO/OiRuhuMRBJ5UoFqsBWbk30MlBZRDuun0kX4FWpYraRwgNvB9mxjl5Qsy5yR
SYNT3M7OB3W8qi4DojXR55kqV1Hj+LHT9C78cTYLfdMzSP5tbPILFvXdlTT1CDKX
Y3iwRHn1+7kJc02lDE1hgI5MwRp6MdQzG7S5NMVf4D1p4pJyFquPTeuGF5NSu9JW
Tr2BGvLodYoZLEIUbi9sd4n9IKzNNE9AagGlTncgf67CQDWuqh4kL/bFBctb7e9d
R9OH9QnEnfgNgEdLpxJh+XtZ/11+fFdFve9eWnF1LMMmNCnm/rYxaievKV/3bbCq
jNmgy8bjyTtiiVls0CAt9piuvbeq/yf//hNgoSR5z3Smz3L5HVvfrcCI0pZAnMrI
L7iKpp+jw0BrR/j7BffuF/FCLj+AEJxBnKojYoTaRkLIuL2qMDgkEspgXVUnZrHd
UFkA1ULIHZ3i4HGGuQIdtM3mZVu/rKtm0XolT+pMIQZV6C5duyMfLBAWLcop7fEE
LB8dwvQM6NhUKLh5erOM6UK3gdFeaK0sFoRtCNjaov1k5o0gFJ30jtOq/+Kq4m2j
emzSruoHyyNkpMPhaxgQriumNroxO3mRA3SRrfAnhUucPfNFayzUmwg2uRVuLbsu
+tcuyNNcAQ+XpFjHp5mZYDKLl0p4Lo8BKr9XSi1n/hBzBpOGUY7+pvcReLuEgUO5
XnpBoG7OaUaQFfx30PVVAK48ElqCH7nAlvNCvAG/P0aJjA1TOCaFXTRB4EeJAC3j
Gmq1h0FY4pJ7BuF3q1ooAb0yBLI7m1MWaXtc1BzVFTG09RRQ443okxVHiN7UaUmh
zui/uxkD5pu5mIZkHnD7L5pnEoOmof1MazLOSN5cpk1rG+o+Ac2pP1cWDNqNbYQS
I1F+2J86C45e7iPZnYlK9qS/43LMR/pA694v27HVqCkwuEnB6dYqJRksEuh91r6U
42bO4gFPVWNjUojsDmJx4BC5qXpu39H18njDNF/w8453Pg6w9oHlcdc7Oi1Dd38i
aOX7afMic2xODDvussibYubMOXOY+ygU2f/dea8qGU73PJEAopnzFl7r4ala13zt
w7UTTb1NyZyPAdKEFa50irMatOe4MJptYyluVzKjW8dGDgtc5kKumPWKoGWbzBF4
T1eoF/6Bl3iqGpd8Jzj/KYE41nxzO7NVGSs2+2SiUCQIywKPI34ykLH7zZSLODyN
fDmbj/750/udt640Sxh28+cVkMCtd5KFj5OxFSgeN0zd332KpUcgJPwkt9C/6K2O
zcMS8c3bY4VpPATaTqP1/tZ5cLaPFqfuLgJjJr8XAXsUrMBX076GZjHl0BsLxGfD
6eae8jtPLsmcqHCk0pigttlH+9CSyJm+cQolqcNt2DdGwckxJ9Kc7CVt7WX5ZvLY
fk0cWMsuFebMS9i0N0dlyGw2E2ckvVKTllyY4aal9as1VKKz4Pri/UcjrJagbEbL
doy2mG8jPvsJDo9XR7vE/qESGjj1X7BjpB4CGGrNE5/Ct26359TSLo+5c4zEzuLE
Aul826sdb7MkRayRPKfilJhDCYFdD0Uo16WhN9QLJOidQbq+kFqaF1Cu1WcyAO+j
kZLdzkbNOHAhgwXk8r+qrf612Z4s/5RTt31nyZADyMbVbV0OfwAhfv9DfNna3k0A
iZwkNl/TIpnyRJUQEMVIslIXEzoR0VGiciua2KUDBP4SAqnQSA+Ks9gVIurwhvgC
mtO9w416pNfFp06fMuUObNxwE4aO0tvaNqi7LapQLv5MwzY9l0WBC0kpH7zy69fu
DKbEvJ/qsV2evPcF2Zqo3RcRa2Aeg35F88ppvfsnyC0Gca4NxNf5wtStncAQMgC6
XK2Qtp/tloGaMhGnVy0MWAT8VB5+sau5y3X3mvSHif+rnjSiI26wnQOti/4xNB5n
q7TC4PrGg++HEFzmfmG81/Vgl9EE4NALUuxA/XfR+bew14O0FIPmo3lihTkxWJp2
XdZmFsYbZ66Oyj+JWUqlE8KPCHE7/fy7+YJHPHtMb/u++10tBruvaWJWGttXxMJI
aFmGkmMUTDo3bMeYetdlOevwGv+3hHHYqyD4k7IydO4cVLWEAk2gVAF761pHmIHJ
ewJ/L/3m1OLiro/gJdUh5CnSLLc6tay5d6tRzNQZ1QysSoQJMd7vGlwAioOWTkCE
iFZOE3yJ6FMUSv9QWhAyLATLxAELZKeByePXdyrluV/HAdt7vXN+AksvdUZxPtA4
zCWlRvvtM4YkKYuTOCYEPUcMEEUyPdgTbbqrW+ARyHWKvzcui0hSsmekBKi+a2l4
+MuopEnA91ypVyzLSkmymuSPsYC6CUqxDz8swFryRz+wWPiH482N8w2TR9AipMVA
xFwHFesPwrzeXTxV1a0IMG3nv2IlBMI3K5JNloi8B54x7cHMm3c13KvmMHX/zqbt
kNOsWqkfhKqoKg0IQhRRZEiatFl/cduoWbVVydedRf41qPIeA6DJapQ8hG0X0hOe
ullFZcKPRiDqQHFmWSiv9XgxfyVA0aH8x4tbB41WXNPEiAc7dicmeGIc1sqORAY5
BnJpzYHgEbxeluG3PtqVM09FbMximyefmSIsnHsNTL/YLiyMQ7B8ScCpNJyjczBr
MmvjZCA/qjRObKJaeWicDdyl++zrocSTY+8U8U5i4xvmweJ10CGeMTlmzcSCopTo
jw47vKpT/ttvLRGSo98log6KWSqLbJ1tmtHDiXOpOrjI0urelT2KCW1eyQgMKu/L
5LQphVGnDTa9eC+n9Uklq8sAiKnvDAI49VQHJppbGBulFdSbwCfg7xnq8rPRlddt
0cfOmFfs91+r6U92jrnkiDHHln0sZ5DVEu3+gc4rw4skGiCkAE0bnbEeH1KjEsY0
M/26Re43oPW152LlT2ClyDQNboi5QIODrgN6/twFgWoZc4UM8fELPattZvTt0xza
FA2jZVI0LKSHvu8Nwzeuqx4V9Gg+fgwPxd9RmHfFWyx/jxDT5SDmdtvt4vQEw/YF
+FzNBUMiGfQURRIgHThE74jqCvEZoEQDC0qolNx17gyVTVnxQ69Ab3z5PMiXjmf3
SbnaBQagstx7dBVhsBk2XNqjQSYR3HDE3Wdac+wl3PayU/WLufCpptgYpQ5EW5b9
U4WuOEkqEM3VIru499fcoYRPdrJf8JyJ2LeGicdU3j/TNOgN35tO6D7yIZgjZIcJ
se8j5+pMMvtKS9oI8/Zu+KCV4EfuVkctIdcV+yYxDlR18EjizdPtQ3pWIq9i/y6X
COQYpAaefzlODjHNuITMBKWV6r2HvWtmisxvBb4erVNf2XqvkFpaoYUN3bnG1Be5
bXF7/mrZDYmrRp08u8aP667W2J3Fv160yoHq0Ag5arJ62aD6K0Bu5BUnTOESdpi+
1nqBM+QyW2O3gAFKnG6B/EzFoA+LkSVjozTN/o7g8baFaez0yMMEh8p8bjyE3I/K
LFmde/8PeIT2w/li/Ezjl89yEuknKbEjiE36UuxPYEdFAvQBQ9/wL1kV9I1ciOpg
+Mhx9CwWtXK17M4Yr8UGUPCNJdMsy1CasYUEWIxC906NkkRxW8suEPqqNRv5ozuO
No92REFND4hEGmIPp3IWM+a5wO8FvhAjtkOA7KBqvJU9qfRzmxDsJ/up64CEgyAp
JP1dI++8C3Vod+2vB04qig2yLVxY00f5PCDnwi3PQP4Aq/WQHxY3YRnu5GFC3tgG
3+/17XZv1RvEZVF+WTOk9T2f9CQl9Vvnni66uGvGe4sAHe2PO99aIzlcxMOX4lRd
QLj6zm2npppNa7/65wb4OYPci2IDNwr/DXeTH8rnMpgXdSjNqfduRceEd9yYOtyb
1Ez6aXD21tClGcqcIc9QdVfN3RzGVoR0b4A35HX1MxLxhdR2hMoZVEDk3mL4ONhH
NFvgf0fW/uM3oyO65AxsUMcxPeXFa/lu+dfP5HCYb9s5rHvLPQ4RUg3MPc7WYpRW
er7nnx0OtyvQFhS7pSut1GGc2aX3mLryKkl7JOiV3BEd4rnem1AYz0oJfJEpH7EM
hcVqSmmlhJEodX4K0Jm4NTVw4Tep8OkKErJRwRXjl5Lsg1BMGjXsbyQLCSWG6ot3
th7t0RikEyB3l6axy6dmjcE8WZDSA7KMDCu5x13MVCbzBWbLCobq+mRNMKmMrYC0
BcfpGE59gupaGgrPnADs4+T+tDhCVGo5uvZuWlcn7Oz8XEUx35YN8ghs5jwRFJih
PgsaZu6pPjh+jDAJum6xN1+cLjDuSEnqSQP0kvapR4uGDi9McS8jlX33BluahfU8
CsgX2FWtRPY2k+a4V7Ugc5mWHR6Kx7NpVXynNH4OOnH56vmclx5/FwsgK/w58YzT
24F0QM8AMZq6vZjhJG4oDaXkluCuGYxrqMwhp0cYFQo5jSakrP4IP40nebS5ZlYa
nTWK6kXNZrwdiaXj+DKyqT04LvpgSdYaVBDlkIGTshmXWiMdMvB8vqaoFltYQInC
jq4r1Q+4vkR2bczFOCg7YvN87ijVE1Cput/vt6tuYxRTKX0JFq2p9cAKplP5O6HS
4+wlp8Yfr+Dg8BqhdNMLoznH3nDhOjseWEjlUjoHO4rUOJluGb78qy8WcY62yMPl
N3flnw93FUSljtzCK6z2kDx5jR9PDMl18chSzl68kX1gFTJxJJzKWUE8sbK3aOqc
1/213fj+3VqqEMbXk0m92nFTa44ReQN/rpSn20WBL9rXefuOYKGWrng4tzniSwSs
3GuDdeI8FemgxvskdY6hPGNC8BUFZRjN+PT0JwLrt6qv/MvWeMRPvW8dru7/+qES
0NJmRmhumfpf5RHll6Vj6U6yO/Q0PrKgJmF/UY3MVxSEOdjIQRLwWfurXaBU2l1p
gDUXTlLkqsF3O1afqpQpCZbeuzFcDLtZEx+GDTSyQJAG0dMfhtP+q0cVzcd9X8fN
oYxZ8t4B4Ltd4O4+QLGlqdFMcYzJYvA0ebn6xIveRsLUyFUhlGE4+G0sUh1ntYKF
liWKBwhCJ3bidPwAqWrwhhBrOe8AZW9Xisbl+jhxo5ZsahDe7GJ7ucSPtc429eSa
H0zhIQwCoqCjCyhMrppPR1kvU7q83PTrRWp/UCiFUbnPuH61mPjICnvY6MhvaY8A
IWe2vQrycy7M0qmvdK2Wj1Lkzsw3UJgo1YTeVr0+vviGMx1qgLudiRSpyf8+FOab
Ur9JyEPo9RRKprvoKGPvqKolsJYMjxLg6f7VVizNkL6nLXuzVzJx6Aublf1sCPHB
D1OvHuDfhqaUbcKbgwY95NyMcx9m4ThwQ+kd6kx34RLt+FWYh3+DC1Q+fI4iVmoM
cezuFObGlJmvJ6ZKuPIQB4FO1hP3TlTy3SNn/kRLoGS3xczxvz2khATu1apru03W
MJUGsAbQ0psPLgdhID2syNt1NqPIiOdtfax3oRXPp7TxXtwWwziCAVFN/MZn9C14
jGHGSQgIb+fgHzIiOZH0Yq/u0jiheyy1ubfRH9Tl10WLbx04ru2wOT/HNF9nCpZp
OtIwy9fwiE+N0ekeE9TOlJg5lXCXYIm1ibAQ56haBuA+Fst1mcJik7ceIf4ul3+U
qqsbAeQtH9/VeU0bPFS5SUD0j4AWv0DmE8WK1bsRx68vliUrC2bQD96yA/vg1o4y
TR31KZzWVWmZUFDVMKzeZTluGjxlxwJgtFR+AZC3Y6mfc1dX/s6I5oWCrt1ImdQK
dX9EEkNAWz9GrewHia+vgInGeelSh6d31JUPVAWspxFOcn2dVI9oVffIeKQsn2Mz
TrpGJ+l6rSad7RsZ6ucTnaSFN0pCaYmie2kyeFcHYJsUD4nA20tslLThNMvA/Y1C
OTY9kl2xZ8QXMvnzh5EHgEopjavyPENcrU+lfqSWXdOJyKwlwgls21NpvMZblRrN
fPjyWw+2/0V/LsKC63PPPpD01IkEy1KASxDxzmdSmdhw34re1ODJQpvmBMGhbm/R
DV7t12Xbhdd56MyFyG2GXZwRy1iBFZ5MPhPx2KWfBNpeB4f4z//d5z/yYtcBN+3V
tN5tfKdbnOY121dqGoVqG9LXNA64TCTNQ7J8xg6ZPxsqFgow2iBQFKxVsiuAvIqV
1hewUykGNDEAQX39avu6HhgzJOYi5XitsKNQcnbmFBsjVXrMLUBgrgSOu2UYKtYR
oCaJmWf319/3I7yoppZ7gX0meIgV/2CZV8Yvzb2TGtX+JG3umt21H305mnKJVbLs
fCmnXwNE8LdfV8tC/Rry/rcW/6vBswm6Fj1L6g9jh2KXwLEyLRYxSs7Ptr6IYSFE
ajMFS+16lQ7m87GMOv3/aCdBGx00cOsOFneJCXvP8f+tQmBNlHUKdTVIDPrmLKQ9
Ylzy83WIEmdfzPXF/dd9T+b5P6xVsW6L4Ul7xLKRtPgToSA2j+i4v+41n4X+3lYE
g2tXb7sCZjSUXsRLpIUgDr2b6VUhoUalw3jz2qVB5lBERdNSsidUn01wl+M6e8Hz
k0jzR1Z/7lz1KIHAg49MUbCVZ5bkHJduzRrZ55EISM+YBDV7KvfP/THmYrtNaWwG
KfdzHxFJ0S9mcM7M/E2neLsrNyR5nQRm4GvyKozqbEfg1is9YF8eo+TQ4p0ffvzh
Gr8T+4DfZ0auuiHgpPH1OVQOdCk57rzsCcxkVs4/syeV7a1p/3aKUBJoTWAnq+vl
ETRHm3vvxAIFO0oeTwnbvvemeVTf2fxZWDLHbrslQmdSBH+6qgID1iNdHkDGs6GM
oH9UW7Kw+1d/KubRNOPmtEGrHdtHdBXc5UC7ZYbRlxNqPl3afi6SGa+SdNsI37s1
v/O+UJ0b91TS50OgnTh0ZPMfoDvN5LawaUGKC2hEVeAvMGmcWp1OhuIwm5n0/r2Q
f2/JCq9mFJ1nQTDMMe81K6KqZtYqaaLA5OsWsvZqCLHTNvekmcTVMU0FSZa3zSxE
GA1nqsD1Mtps6AhSpdKLQNQBf8UaN4mZrOxSTlqM4L8wjBkcxqmpPjXSgXHJgd06
4b61ny4NzDoVbBw/MaCiPzGMgF3ZJcvtNgogfGAZGfLuxVBipJ/5xIdhfQXxVIQB
RGPSpbIfPkmslYW/Y2QHUnQEU2LzNvOxuC+nViM5QKMi7mD2ePRsIU7GC1lY+m5l
jBT68KLdxKAmzVJzcCUQZAnVovSPWMQ5zTXPRLgasoe8Reu4Y3K9LY+GVUt4DFXo
fFd+D0B4vQgGKYgeAXWn065PxJQv6k20KnjF6yhPAqvCXd+FGgvQY0Wc7slqXiyI
SAAYVdCRcwoTWAw5jOPX+kMjKyJJlfozewEfRQG0WjyoHpXkuTS4zCyuZWZ5Zxxy
zV5geNisrQVUUAVXBd0eC2Lei2VU+T05VQZ4UUNJcBPrniDIBwBsvMtG+jMMrgSa
y/37M+2lT8GkBVK8WKCioWgY8rtV9D4CTwZCGlgJnMULy8hzt1IhftJrkR/ec7SK
QBQJszS6jMqDO+xVzjkvGSZppk/6fMsyrpivqAN25gP0I/Tz3quYQ93aDoyEtrVP
3KDnmuN454XXwU2/zzgAAPPN9Csv9mX1LBnY18w/SMyrdLrDA/t+3OFmSzIiE2hS
O2yWTRUXffJyvJfM7H4C8v0BX5jzkZyGLZHd5gnKvPi7YugeVAOWgkSUdQMLYcX2
8ajpiR85vaXJJiHdXc9DHv0XmYXbuB7LDJ4WtVeRr85ibMwg0np/BLgkXadYXq+q
4w1o7wCHD+/hyR6qnrBYK5053dGHc4mq0sI3+h6tIQPZvJIYjusjkHJnU84pLaTN
km08uKfPBEU/6F1ZKuDy3OOnzFGDYVGv1sMQy7dMwV9RE8rZZHbMaWlGSkeZttzM
xgDaqYpMIXdoBzNLGmScLFXbIs5qixKgZp9fkRyvt2n2l52OmSDBu9JgAF4UiELv
/T21218VlYzlTNXwHoyzc090m2KpWK58SaS8o+zmiNFL2RBXUI5qnDlvE/jPjuGy
aBijrf2hXASgRR3cwPJioJ3WZD1XUTW7CyjL97AdUGvArpzC4w7XqRHsXmREkNmh
zOnDBR0JWcSDbIsM5AZKVhdJw+/F0evuIHV/25Lsoe8UmHay9cMBczPQYfwAgAoE
O/I0t1l4xgv8MOcbCj/vovOn3k4Y6+byickk8lcJQlfFi8MevWvRWmp81IgK2HCB
BN5CAf0u+L2kwgGrQxF/ajhr3oGlAJkzSU02RcMVBWzWHhaG7n+jBtxTjySKhmNI
f9TN1HVU/A1nAo09d+RbkKN8c75qzt5y0ekl6kWUFde7UV/yegUGhe0Q3ZI8dhxB
QMk6MEdrbcQnnyeypK9D5L/49Nn0+Jn+r7Ra7qcluN+hZu3APqbhPAFSfRft2/ZK
3upW7BAFIgM937tJXL+FNhxe/1zoQsMIytifePphMJj2sjEiUi958pulykxhUsnP
5KDN+dpgauTxHAyR8W7MNR8xTZ6jML25dNanv/pIUovVWL7whFEX1t3c/d18h9r5
f8Nhqw6MV0v3skVUcuF/5Z5DGmICF3irRwMyvxTjyb/EwDo73MWCJegxsMRyxLB8
qON8DrhvIS4mq2BXgIhSyZ+gW/9rZMHDOhLFOWkHcSpiGTwhlQfVJA3Kb+jjWd8c
U4BHbPKnnDFKVC04JgROMvROFb9MdP2WULILHD1FSWX+CydPxYRA109hTMPAxBpe
FYVAgbrr7JgyiYJJ8GyaZ8Zz2Erfu7qm/CGhJ8hXzUClmwOwPSjmiaIW2Em8fs5/
VGKaLnZDlbRgovMcUfPTGafkFJDLZRRt2u2gzvQb70VGxDF07mbysLAgPymZckV2
zHpq6JAocAHpc2Mqq40DV6vVzdJL8q8sdXXRPvAUyFVMjxQIr6j5U9vmxQn/nq9y
3EeWadWtxzwZJLSBlARSpC56L2zUAI6z8uoUXsDdbUHOCW8G+9ogEZf5WbyJ6G6l
jtp05xddnXPKwEQNdA8N/Vr79wUuEF5WM+SynLS1MY51kzeP/gj77azfv25T878R
KFUXjso/2vbU9TKq/7t/cAkDd/Cf1RmzpmulIwYEPQUGdVu02N0gZ7E5hHhKq+ZS
Wzlk+uBJQYlyI97GEz6rH8HjhmgOW6C9v6UGY75Xsa2+pJkoMbBV9TJ18HiM/cmq
Jx9nl58F9rIMD2YNHTqJmN7VH4FuaTtuQfvI3AdEa/sqKtIFv8z/NE1Eiu7Y/0yj
95ZAaf73NtrT31TUu/c5FN7fD60hFnkMFFnn2rE4EXAqMmQceh1v1xrCeF8Z//4b
gNyCEi2bdTZgFKkBSrZ4gMnu8tqbE1gNw5vmwS6nyMmLcCmheeq1biev4f1RJ72T
5gtmRVToLtCvZbY+ZdffQZMm9MH46sExCnFmGZYdX3ZljUiLmX3IlX5eveeg0mLu
hVCM620ImP+3I0so+5k0RS01BCXGtQr35yBPiNlkQCn1R/KNa04TKQczsrLj8nxH
1p09bbXxIGt6ElMkjdG0YtudgnMMPFf3yIraRQbfTEvtyXPgNTiOoxmJBaAVl/QR
t46A5C+wG1r6RHG+oZGYLgZfnghwNwKKCSAZKlpHLG23Ut4cVmKHQrM8PSIEiYqQ
TDN7Ua322sCSfec+TZf0ETmHbB03lfECRUI9b75SBdX3Rrw1KiPMHz0s2det0WvO
M2SkXLHmDQS6iSOHu4ISFOQqCVl+9e7/hofb11HcyQAaoq1b8GgreKwa3Rdg0dNb
xReGIGwJa4ENtGoJxWCcFLsTkuaSYBIDM2vEP9kxRT0iXj1/tcJLrSmt3DfkfDmO
HI4i3Kbf60fvHiczQj+hkjKwRtQrRhRvwjOWNACUbcIIA2J1FAQJIlRE2jfiFioW
xThFG2GJ8N8CzdntgEqEhg1tU48J6vfMx3Y1ptiiK35A8MhBYDLRTKY1a+qcSJSx
Qj+wd2xn5O7UztcPyYxhpRTH22l9Gz79VeD0vQFtB9W620xD6XZo3mhXiSbFeM9i
Ffc3uXWBr5CG4odxte+Vn1NX/MJ0lFE7iqKWCxOVKKUKnFYwapmQLp2n+h2G3w4X
wVLuPYpSr0Eh/l8H+So5mws1twEv9Ue/p6YhWSvo2Ss0LGb/TC/ZVOuQSEuYl5s5
AEn24T5UGXIOKhTjCh7EC9KE8HG4AGGQsBTPNukb04tRdnvbFgGvC9SNrVRmCvS/
qi7D/4rvwYVMTnlcw8SD4XllSOZIEsteVmP2NUOeoVZhVWRoeWfkIE3TNHrZigK6
+yDXP43X44NyUdLklwAN2OIDdaXHxqvey8/aDOIXWrdK7xO4D/hCfNp4Eblu2PSQ
vfsm+XEsd3PCeo8XYtGt85SY+n2L2v9H7Hl+p0mjLLPOYVTCDfAO65cxFWd3qVce
LnpLyzI/cUOZj1GqeJWpv+sytG/6qV/JN4SGcl4PXvs/B0lsDFG5Hx+WA94E0nmi
OE5BP26yeiUFOM235Cis4GDfI8A0bPKxezpp6DpyChbBQJLIvQikb0b1qy0iFYGO
rPZlUd2IA7g7PAdERgWGvHGXlNVTNLbSmPgU6sImJzyS+Ggp50f7zuD/1FzYhgnw
sra6d7YX/GS+m3w+2kEdFwsv7vLPeCwKvv5zXkEcm6FWRcyhJIa4WmWDtZTXDHfW
Oytg5Ch3XorNE2xKR2ImD8oEahiCifwgQjmouUSOxoDCispTwVPhmLCgeN8SSQRf
9ytKacbq7zt+VnQv3MHplqICDIUgbNio9wZlqJ+ZbBgC7v8KeK0Sdru94wpcasEN
CdyX7/YGd844aknyNAPceKdUmNH/hsMo5Z7WYRY0WpN4QVP4CTfr3zsgHEYmLNOT
74tqJGJsHqgZ0aimfNWo+MfHze4K9kRz2owVnt+B0cs6LYnPpkhdPfxy6U0I25ue
bAFapaD0NWMMbRTL3u3IUMed/VJg94WRfKuNai3UDwb4yozwisnmHJPLuSLpLeBE
swntsRaT6jqYl2ctHFcVg6psSU7bPxahOlSXeTumU74U3Uy9cvITn/CQXiCCEFLr
8NQ0RJ35eSYM3PXW+k3XQlL8C/x8FqBFEiuQNLeQWwXLEEleyFO8LWwvcuLmVh6m
jTNivQfyNdEot6MWx5LYoPvlj5SLLD0mecKDVKSuDtErQtRclG9KIMFj6rHpJ/ij
mzTvmYoqQoHQHOdYu+sluskBeEmEYBRHzak3J/satfcN9GjjncQgQuqd7WuGrno1
zJQ02HOqgQF5c8Z2Dpvh6/N9+RIhQ6aBJveQWBTyQNU5AKytmxPxy6GTbigWVU62
X3SvG4MjOioWyzUfylKcnx+BNsEQ331Ot/QzaUkLy3UPnK0QkOLyNMLsOQyQ9Jtl
ixXbAkNkcS9MTL/vzEqPwbBqgJ4DJ7l8AsMqx+HJ/bwS5h/GQFFg6oLtIzew2v59
4Lfes0/L6FJYhnCEbe2REft5XagcNynEiXHXppV7UVuCqngTVok28RHyW0l7kmZE
QhDyBv5fFLCE/g/5OVVwo6DXlyQ+hQXNCf5gNUYlLMRFulvdGZDtwlsv5Zr+iTB0
dynCCI/ruvaCSuEgqNtFM/9oMdZhw1be1ivr0z7dgmDkgdNCmC18+0CebSXDem8A
K78Lfb23/aNUuMaqUnfXDei/OIkzR7r1ojh5JD7Zz3vciOAvMKuZjUy7/Z3h6QrK
CWYDAuRmMjh0ZjM22Ypd5aVgQUeAA6+33TuywGoDqpsgrJLdFoLQfau0LjsZy+Gj
R/cU8ULstrcI/VfN8ZWpIhcO6mF7vqvQa5gk1jN7kWPsJ0CbOOtFI1Cz/VKsMlr6
g/aqg7YJKZjDDaza5vzKSlQ0Qp5QKApJbuZowOwa1gCZ/UJB+FB+lTt/ma3Yb8ed
ipkr/7c4eczabp4BQ/61a5SvkkFsHt14M1do+nuIIFkQGfAiM/Ud5ev3am+WxkGL
LaBP5M2HqVNp16I7C14X4glr7lf2hhD7lZAxbqoXmCfV0m3GHnLFXrpaZQu1cIDg
uDm0e4bYxfVzh+VrigqFGLvRntI7Tvc+3jagiE7QERT5Y99thdnjCDUXL4Uqo+z6
2FVi4r5CezC68nAYZ/8Bp/GRt9BcKnA3zfrnQKTjzSMilmHOnOFKNK/m/yeOTLJM
ev8Hhe+pGta+J/bjJbZ8RSUP9AeufDvkoJI1gW47RqioNxk00r6RAn0bxGsyf05D
UeLCcYtPtlmIoMU8orczbhuSyETxD+mKD0HCqCDLh5w91EwYjSQYZl/C+lo5J191
/Tf/s7IMkjvg3F1qk/ifXoaFHBMNdJdIiVGBgLrNDiAcf1Jj1Ons/zACN9IMpZTa
YAAc1403BcnMGbzNVZla89+mXbcSybVVPDKu/VdQ+fY8QycE4S8bCgPt4i1XoqNt
E2GSyZsef0NVZYyP64jUlAUJoRyJ+tKF8ufRFVazmXi27LhdLFpDJZMvX7Ab7MpS
eCa1yQ2WXBfq18aNccJErJe9WE47KYL4FIQy8o7TyVhoGlT5mDRAW3x8PH1kJzlc
JwzH/oPJXoZJpMHG7mMR2Pd6q7fsljR235k+XbYKUdlbD72uoT3wnlvAP0O2dFa5
g/masB/dzRbSwQWjQctvb6VOWgqONgKbYKO598MtirIWXUJbxlQYV8OuJOLhmhxW
Tq5395HKFYgxucHIXKD1c7kJsuStlkgjk76EmxEDPSyNvCU9F7mA6qd8kq7bJUwx
pqRTFZA5GQYYkbYjFpbp6fTYzbrr4U0F4MbO9gGxlLs2gj78NeWZWQQnW9YbetMl
DSmaOz38GACeF1gSvC/B3tQjcKAPmgJSqa+2ODACc72lx+s9Q/PZJuF6Ejxb8GA+
ZAcT8A3Qp8TAXIAnPCE1z2+cqYRcP11sBl94zI3cmUyciT7VQFVl2sR43YhcDUCm
GzRGcZdRp2mzHVLjuju9z9My05h/aZxYNP2RgZEscypLeCW+kP+ujQts+ghCt4bn
m8Zn9v0F/KabxXnVRdWE7JZKiAFqYrZrkURSCWhMvQuJMMB+WUjmM3jM3OJTUKZh
JRxj+F/iEOK1x+1VO9X3pOFQ1VlU+GXgVgzzzwh37f5+mudeeZ8KN1zs5TX9ObFO
x/invdnDCR2Av6NlzqFXmXSLjyTjEMZkYFDiBjEcIPVDHf+f4ecG1FpHtR03e/PE
ROOMQEs48afrXip0AnYSqUR/WX6OuWcKcwQqRFk5/uYy5KcOg0PA25ysT7P6522C
wEwPpwVGs0jZR7NLSMoGv0tRY7iMht+lsr/bhWqZQzcZcfYMboePhzegvN4f/Jhz
IL7geYLBPdnd/LDr/I69EBag5tfOSUSZ+t3SSG+Tpx/0BNlLrLCbMLaMcmNc7pSm
+hI2XV2GxOZZzt5CRRyYlIlnzwM5TlOC8lrkIuuSa/tqd15vTUqYs6l1RlRybcAl
KsbNVRqAsUPCeWTvkzO0yO1iVN8UEKyEu8Ds0NG0EGfip87v6vxhuETMmGxtlj1n
CtcohcFmRosjmAeQd/T22hvS9/eHRl2QAX5doCp3ykerzhwymSean4ButOymlIJw
G0vejw+Bxq2nzb0Lvvmug1sc5eloZkhQRzrDLnwIvhKpsXYjOH49YufCuZwB84/N
sAE9QuKYnyNDYxlRPyy8Z6x+QtCJKsPHXVCiYqcvePvRxegVC88ALRJFq2p/+BN2
wt3t/ZajXcZWFiuOROexOGVRDVjUFygFAw38RQDOjZLe8zUUe/HIYVEHt5wiPz/6
DDYGNSAqkt+0pP3cVS410z24gKYT9bnVAwcpgJish0mOfbpYqn+J4sa8nd/ZHiCl
BUbHQVrZrXckpLkpf5fW/f3aqliwnq3EwsdAgWXqf22KO2fc4njhD4FjX3+IMM/v
Lgd+jRACw5EXaHDWzLohWMLLPV3FPQv9guWcVuUC5hz5LXoY0YQWPeoJNRehJZd0
WEMgJ3szLZ7qajSQM7Om1YM2VTXdv8gCybWgN7njloKZ7vdcFhZGERgazPkufhdZ
pn0VoBuxneaFhIK6UepwQq+IpzG0CyhsToq9lj0QF7yVDejEpx/Z0z8PsCL/OxjO
9mRBRKWdiQxsBGVjW9AobdyQ+59oHzXKkhBc4pbX5jSsw4uBeqUe15yDIAmPsmZL
L9LiH+5hBSQvSMq+ncUcDBBGmFF54HMSzyMzO6zaVvxgcVF5MxKeO85ePa6v690H
WydCY9OSFY6cAzSqwIxX1atRNn/AIwP79dgbzeJhK9zRiTNkaf5ItHVvzMPDoDu3
0CaE9bs9Cgm20pRzLQ7RhsOpF3e5HzHW8lyG/QOLMKO93mDyjqnpW8jtF9LXcqAo
JSOM6b2YhFeYD97OBr9AtLcM2NpimdFE9YlOxh0SzkUJENScNGiYlB2c3aNqVLAF
UU70yj2/eRlO1Xlq6gCxLcNjk2SzUrjeaMCakYtRz4DbyAhGEIRyht6lO6Yl+aSN
9zAZdqeCe/rWeCs5zFQHVyfisVN+9fAMrAWYODy/ASwL9po26sYzxLRc7zbOtomR
gdOIVeJMMove0qjIKRCBZET2L25y914uEOYFjXqLBT7NjJH7GFhsDhq2SepCYpfH
5BzXnVEaKEIwfJ50oNKgiSB7zok54p90g/NY+zhdalHKwcKhQUgL4iIAznO0TbWc
OzVCslSXDR1f3K/iRwcXr+DW89/LmQSKgGDbXPpE2Y6FoDARBYpeMA5t8PhrMjxV
cf0uSx079MdPhehzTA6QDDwlSWva0gcjbtKowGwHClorRHyYFQKZvphPGWwiTLe6
MCLLVPGVsKF30t/b/XQ84ZfTMWkSDHve4xKP2eEuE8fQQmdd0dkk+/6/SQhOA+d5
pLaDbf55Mr+CcUbZcqSI7YQs59A9X2kUb4lLHsKjYnJ3AARtHjaf0nk6h9EDSjl2
gJTcVb6E3U4YGShcYWE0PNcrVDXm2qAab5Wm1BTUEGN5t+fvb0UORd7tr76x1Uoq
xSfYN7bvvwgB78BbxiE0/wxDZVBmf3qWLw2rkqLOw96G8ppXsyHObFAfH231+EdH
GQ71xxGhRibmdVgQimPPRx3WUhZxMShdbQ1yeGqKyFo7kQBJHL3qXkKMze+Gh6PZ
/LEpPvHrwlH7ElIHr8Vz+zREplOtI+QdJrPyOUD0ORxIeoeEJ6W2bdBtw3FcO8Y7
1IX7Kt98b0n/zWycANplg6kMdpQFARGagZ6TgToi9nkOJ9mXWjd2batfUURzEEry
cJu0W7s9iRdNIffwKeB3zCBkaJ9N7W/N0AfIeNaxRswvG1NZZ7AOpc6kuqk5MLe7
nrTYsyDUanYVtmy6WPIuTTIStrgfMEb0e2XSaRQGvwh2o2cQdgJz4779w662kFc8
MhPsv20meJLZ/KAdzzo4hHzBsDw6oI/MyIwy7mnSWzip39nn1LogCfzYImG1h638
xGMmOJ3LFKcAPAQAEOL4SkpihXZWedIZNVQnLyZQbd1sRl2YFSpd4TDJ44duFZSu
UlfSBigYGYWrLPjCMqsUPcuvSJrn0TugntV5GDtJ0nxbNrJxmzee17VUxA5mEh8B
/rLSWu/eKTYjWfML9iRYzp4twLNOvw58U2nV2NDBIJHVh8Gt2v3SUvYUKBFDEyio
fWoNPNB2cbx8N4j9w2ed2ctwei2LZe6HJzERRzD7LsAlTetQ8JqIB9/jUVnKWTaN
klTM0lroZncCGfq1Dg0fnCATmAmZ8SxPdFP2SFo8mMKm0yP5dSGE1aIYEDKxMBds
5aZefDzx6L06x0aSoWWqJZgXJzPFO6tf/cgsJYAWQ7DhCc1aMHA7SvLBypxVTQGk
39cODCllDyjw0jZW3KMplrNyjNa1bu6weFqHku3Q3v8yUwJb2uiVYvAx89KfB0Jo
iShAyW3+3N76fwY8otiM7OYMSr4/RnwFe92p/bSkf/3e3fumbkFznIaG0SGZ2Lft
oqxdVt+FqnypB2JR/dvP3xkHRzUSlISAAudWPVWVTctOkoaqNjbhmeVnwRhBLbyE
pa4HRaGsd5bLGUO4xSNQNTTwzZOvZFQ4war7LOvCsMzXSnxGbGgXP/74sj5Y6FOM
qnYyBog7g6XVruP0ykuhHSyLYRYRTgN8hhCqTOqGIPwD2rsabn0rEMRtgQEUfNoy
fPtwOAOTohgT8Q1oLWCQ60011AHEsOYa22E5IOmNaMG7yylZcPsbZzlGBxGpgFDU
1KCvaeJMjg0Hn9pMmzJNyCAQq70OQhVYCSL2pVolk1P7xFudkDwpqXz7Rg8VKYvg
f9Q5sa6I22x3Ilq7EAPI/1BP38QFrnXsy4wAeDW49iqZHZEnXBBY+lweXcHaAJrB
Sj3T4hk0w73k2ul7U3ALbTyqD9xKMk0IVGNsOTFCzI4M3iL/8+4weCNTMcdS4KXd
wesIgGEV1/k2iLBVcKoLQ0mJsPiL5Jxrfsif1XhfmeMpQU40/gtweiV2EVM7TPDn
/kCe0dIcA5H6FaVaM4RdXYFk4NErofKrp65BSqX8G+hnYnmr3NDhoODU/n4EJDwZ
hpwQnTAJ+U+7IxlI+IACeUN61FF8YNtmxzk7izAE1oKf00GaOPtrjK4RUHeTbXLN
EVsp4fISzz8iIcE29vCsbdqebwfWvCnNacO/q0SZP5eYxu9C3RcPmB24qYFaj2CH
kUqa2ZLA+cAPFUfDQW9R6+c6wLT/rs6ff1cXLHjxiN8TYCso1Y4Qu6cK0vCPLFKU
Wa0eopqzURqmw+32pN78XkoJAh3VTTIQa862wQA7N8ygYyt5Ue3MOGIGGeqAZdoR
BULr+2Czdu3WIpicaCE312bVg0h8eQOvH6Lab0eM0gbI4UIidk1VN0Ur6j5vqDUN
XTS+cn8FEnPOK8zBuK1FMzuKfSk0M7b1BiNfnpuciEYYTBf2Z2ZbsjC3fBFRMB5/
6MTA7RRyrZm+ui2Fw5qbgVSrIs+SrQN81rbALV+mWCXu+4viY4p2ojTnM6OjfknE
7W66sqo4DpBo9ve+4WmagCrYFr9VCtcDHtdcesbTMwpuRYtqEyQjXqQKK0LjX1S2
xQa9vWwxFw2Zzrm/ecNwh7Id+ZlX3pVYLnCnym265A1QEf8Adep9+Z2DIq+LTdWV
OeBkwVUcr/59Nkea7zNlNPWFOBox6TJcFj7i7Har5peLmoXcJUMzfASBu9s86n+t
60IyC6LF2+eBhr+p8h1WfoPnlben8YPXQouVsgaJek6uRKgUY22wiOj2r+m05iaJ
n6smGxBPUUmuSd4+YNxPrWrHq38iZ6dSVm1GCgfZrlc8tNllGmqOok9QLa6H8Err
oaAEYP8bb5YtJ7uZqYnWAtpurP2pu+P6MJ1QBxbInnLHgtXFfjZtgLDz5aUNXkn+
oRXrIuIUEZv5n+KoiffqnvWF/mafO22mCCoS+B7p2vWlcxyitR/kZ3ETuTyG0Vrb
QwD1IURJkUz72tZAo8BkV1p7mWy9rbEJHiaxcyp2o2nenNkJHxmIgEV5PqRJmriu
8luHXAS/ZtGQ2P9BGLCtAMyPSdeNH4sjvcEXW03sumZjR8Xk8sA71NvHFq4+cYYR
eB7qev7b8HujAvXSLRPJ8I9PAq8pYwQ8wR0nePjRHUQFmFlEOOvJmOfIj77COM5a
91wbMxNtg+8UYMK1PpX871/ypFQ8E/WOCuiJVLmdJJXjrAeMa3CMGDfQJmUbSbD5
bd6YlwP02yx4NFVTWfFc4EQgHam0IlSNzDrb9ZgNq1AiDpi3XxUFkcKHWPlYKKbu
AZBD5met+XrLerg0vt1iK8AqOSsV4z+0lzk9mEMgAgympuQij/T7OccL07wU9jJI
06p6SP/NDBdoDR8oLAlNCbjam9prBo60K+IueiGoAovG4CYWsURg3+j2FLrFe6Zp
QgIlb6jVZeUOKs3Tiy2dnp2ZFM+nZ3pAZWdtvzhEN5Bm8ED7cfCmtpX1FUg9Z+FT
cvWzsjonIWgx2GxfkUF87qPXiCc3+e49TwG61lJMij2Uqj0aGWzVStJLyIQ7+0jE
FIE2O3JJs3dybth8iwit26i3LzUSXwfNfA5yMYjaYCIuyL6T7pJdA/chYZ8qFnOw
o02L3CipEmP/as7DZzEEZqGFTfsZtRyGx4fcxZtH8XYVoDAUhKt0i/sl+YlT+oLe
6kPLMgDpsLt3t3hLYrNShnDK8UNaJeoOejxjqqZuCmB7X3Q75utAKLDcFKz7lOS/
yJB8ciQDX9bRgHltuRE9FJXzmUHVlbFwK2rH+fXv2YODdHyjD2FWieiv7M897tnx
WYQCavruZDk3FSgjMqpfhM6uwoiqKmR5y8q2KP8dl+2aP9FTRZzVJ7lhAoPNiOc+
BhsIXYgKs333wIwiCsXHb/eQeCwo9OqJGLHOQsPjbAXR/maSSxweA5W0Wh82acqX
OgWEYX0/fXxmSkgkNIGr05y9UcmL3FLLCyXBlxY1ZweIzFPLgncPhDBqD0l+R0Ne
HUkYz+lH4w4nf06hcpJsU7VU3MGrS04AQ78W6aAC5me3Q34qvL6yOacqfjzwvI6z
9eucqMu/NJ5Am1Rb6EVXQXFs93SsEun3FWr9fbZbU/niVV69taMKRJ9+JoU5ZcoR
23pgHP+Q2/yhgBjWOyG5jAb259kDDqQklAlmJ/lEgSrly+/mue5yVumaKA/YHfKb
EWFTKdMKoitWR/ne9ZqVWiH3gPQHUSLdHI1sgseEAaYnTiqw1TFIkZEPsKyUupF4
RbMckVcD/CzsQNa+wJNQzdI9pZ/+mdgxaVYoCFyrR3W/6bNDzG3LD+j/rdqWqiib
ZuBhdaNkO0fvG/qNvT9LX8bunwWyMrGEioyERKbkd3tHwTscptsC5GHO2+9nEnJB
Za9A+6f2JGYsfFPLwQ7l5+ktv7q608fJ0T08ahffPv6w2VcDRoYD7qrMT6GtIbbZ
b96+ajy3sGY95oC9qAJxfIzjFqCE9cb5qG/24UTlY8Pz4pq0al0HByPsxjS+QsHW
rScaVXC9/YgifH+8M0+xMPt7cthMyT9whfJ+rInHnsuFkH84CNi+82x403gY4yy2
Bd+tVDQ9EMQ0lVPG+z2ukXRwA0L+EcKzTT0tEQnrIjugd7N3SLpgNVtNSbhJgFs4
diHEoxog3M47FdRWfDbq0ET7b+cyQCdOBSfq6ivhWibeCjL4isv3y71pV78haSRT
rDUjXgEWfSq2XUxznT2k/RhYu+1VRPyLZTmuPWvIyS11iiWqVnYr7HrvYtbBJhPW
fnA6T9NMpo9INizC2108kAQ2t9WRMtdAKwqDkNl8XPgLx+ycqehG83SOjOursIR+
7rkHQqJPQw+CgYBLcSf6dbl88gaP0C2qB0FSGSkhnd6mv+bPZcScHn9swxWoDo9o
pbzbupwMXfRAzdof0bk2MjV2vDVzXkx6pREN+fHIahlIft9ffpa4HsTO/2alXgr4
jDBoFTFINS/9QSeE51tnE3MdMekBdH0AMmW5D9dsfdga4g9B4mnRK2i5Fd97HWDv
f5LwNhGmxRrwLZFzPn1dKzjRohN053EpKH9s/6DzpeJA4YDPHDlMpX+d4XzckyYt
caLrGZNK92T51FU0nVhpd8CZCxkhe2yfCQzwoJzTzudOvdEIjsGt3pRUirpsdpk4
gZ4scy1cbVmHWVhc7pF85aSQ/Fo+x6Mc0uoRMUdiWEjhamZ8dhOnQX8+Lfv4qdoR
9Ip0InswiPR1mUKnBzhSvgqLd24kTN+PzhQkX/B7PLM/4pLdglaj4QIVMb3nq9pU
j9p7isyy+vU84DcweUL+iaEVmiCUnn9HR89fB7I60uh9MheBLR9Nf+Z+MYTgiXTt
t7zeYUEMhPUBf+2FgU3xA/r6ZQaaBTMvb0Daz8jyp4lGxdIYIysPqm7FExqmx3uy
Oc+gZdmMmgyGcC6GXgKtfVmN3YIZQfe2fAIDPLcS7u6kmwIbXvB+U4fKxFZpwOTW
aRGis1bmLxFz8UzcKiYyqvoTn/8sDG6A8NOsDaDFxrlmLsrmLs104rzHbng3TIZD
kmrrQ/KMDJBGtN6uCH+um2JoZNa4NEH0LKDM5AneqATCuDJtqvEZDEQn+e+JelIM
C5KaScujyInkQ6iqqF6pg6lDAd7OfuoxfiTiSerbhNil9BCyhbZZCBRuRDiF9HjH
2Tl+Tf1uQU1IlpDDXWUNYvu4YglI8v8BWVbZyCQA9cUkjkLjCXWRC3ZgPE+QPm1o
S7kD7mAoyVq4+iKD0li7OoRruJAX8mtq6wLyB5RTkmMgSGPTj0c6oTGVjud1BXZi
6p4sFnZBy7xZgzIuz9dV9BZ/nga6HhpuOuky1gSCu+N5GguC27wVb/SPBclgyflZ
qWt9zWEqQ+GCEsIqpXm1vXJBMtZorj6a9rT6RjGlXpj8uIT+jV28Ra2rouNPIKI0
pmHpU13UNPhva1L3Ky3shjl1g+H9mPIeUAXad8LOIXIru+zfJawW0NZsDbBOeh4q
KqF6ywcasWh+Abq8vhH15dTlyYEBPujRBtot558HA/tJanHK5p+G0ZRToCjCmpOv
YxTFRveWjM4CsQW2r/BOzahiUivUc01n7in+wip7jt9dN2zSYar0Fs+7PZoLtxA5
ZrYUnF42LkZ+67OI8M4jubGQEmsyc4G3xEP3vl23/ftcYhVzmTDIOg8c8c/H85xX
SsYQLK7KbVE5uxPFCUHi68qNqYRAJkzn+ThBqpue8jVxd6Q0OCj6HjX1YLufgl0n
a80Qd0d7YMKm3fed3AsxS+6AING/oavKKDtmOfCSTU072id+EsA8TPN8CAyCCbk5
mSPud1NrVO3TDwzepnAIuSdlTQRgejALErbAnrCLN2sv7kbM3UFQlbGTUlNeRMgv
yYVajtX+GNZQTESoeGPp3dSAtzZ/KITkXzxroM3pQa7gE40Yl9wTeXef9RqfeuwQ
Y324R+WeBGjIvW9ZfKuN6dox/UMNwIq7K0yV/2QzXl1eT/VixoMGiIxyVyIfi3nv
WrZwIH4GbgXU9BluGPIiXmd20nihJy1VAOT0f8/8Mz+3nVwbg+fR9RXZjFK1nE4S
EzgbQbzy+KEBu3303jIYvH+eF92fAp2WkKu6I6AmUPVSU0SJLXrhxthvmv4L/EPS
u8lml6zmfRunNJFl0GZ5948MCrkOcP9pnmy/yXAqC8D0LGM9evl6um6SHYsjP9zS
L9XUYtPyQaH3mSXecmYr4q6ddygoWd0RqwvPID4wHayHzn1L6GfXP16rv/W2ElCQ
nisj8lHIhkTcmNc3FMC24WEF3DQbSlJ8aGkN6eZU4BASVMTgmv9aeSLtwwJvyztj
X3xkLTqNONcm5a2pG5gX/wWR6Jr8jMEbxfgBgyiIwnh9CmEa7dW8b5wLfsPNQkOm
M4Wi/QWkOE2y0NJHQpCBeExpEn8OPyCz4kRXhjrhOIp7xCyYGNl26Y+JEiRcR+mJ
BpQVC//pmpKZenfymMK3QCqUf8O4j4PIwAT9blCFNjt9m9D0TTba68Z9W6KskBsH
fphqCL9mU80oJKxeXAoKbxFKsR8VNFiQv07XJ76kvMwkJFzkwR+5p2/42T4o3o9x
H+RbAsMSFl72rOnnU46nlNe3BHuR0gClfupqqys3xAOCSVmywVuvrc/IQzsSJVw9
oiLXbHOtN8VtSok9bOn9XygZRLUhF+xNZmYYpRNuM2Siu2jloCnQ/ydOnLlA33FV
WVFPB28+4zrt7uDoLaDSAujSDq2JBqiVq0y8cypR9OMe7AzXFF6ne2NYE0tEVdbP
xitrQ2tZ/vRCgG9PME6pzBx9QkRyAmxjyzVKWnxYkxzwB7y12/VNDnZmFv6/EPar
XNr9PmbiGkfZhE2iTXasyE/bJMSwbDOSA0utWKMeIeUAArgbJEA8ABtto2wQMy4O
WJaZblu1mN+3g1gsj2VbSAS/L96YxJdf9j1VfdlIz8LQsQx7oX3tk4Cbd1wlUiK8
6IvXt/TqznHDz2FyHWZ4E9L7Y1aa1fylx3yXxywspISHoRRA44WWy5uJCiwLfevN
/QtVJ7z3bNDpUbgl9dnEEYGlW+fyGgaDz8DhVPwOD1T8Zg8FxvThuIb4HX3keQQI
DWc2bwDsyh/+3cMjsVphAEGFKkr+Swb0VqnAauraifBADbSPcZJ0c6Uyfiqj3foi
I/nIMJMCzZ0QchBLBp+LZOuIBUkY36xGAMR1Kb7Zve6sVRH40WKarxCjkY/4vBY/
sQa/XiwNr22jZQXWHCLQtywDKClPGqDUfXguPOpmG1cGV3y1pIwJIneRkEOqig68
RAR/pl6tK3gXnDKwdWUX3ETnpxtv1IssitCVTSL6+Zinhy7ob1lr6DgZAw8q8t1E
UA9HPmk4DOfabKr7ASwV0s+kLc4QAgzwbHU/97R6vdDLd27/21obkwwKo9GQhDbX
MVMCIel40h7yaNbAvHqmOgE7LGkaV/WRkJigbh50Wni9C3gQaCVY4wcKPyZIDDCn
NR9G4dw4uxY9Q3MXxp3DKlUg6QFEVuSVZWXfHKzOyyJfyjRTXvWoWqKGldrgTsAQ
c/IAFO8XQixjMAr8V4m6Cz8i+DeVSLxW2Gr8xOYLfPFbN9iLO3SQnKQ+vahAl+iX
S8xT4Ha+LIHlcOxShpIO4HQMJSlQTWym4x5S8g2ZbIktgdwuirzFUIMTHGD9HwEy
yZL/TptBarz9JMfT700cqnw4IyrWofRkz99KKmeSUf5Z47LVPFDL+yMVuA7GqyEI
wS+OngaVFizjTN6HJR4+VuBMVohM9Wl330bOnzjOXzeyV60AoGaTS52ukBaZCAx0
fvnVBpmKSEqrDfmiHkNvGWC1rDu0UOltSCsMsHbcKGh6RKZe+ukDA8Y+qi4VT/ZU
dJV8yhpDdWwBjqAb4Wq2mx3YY273B3mZVOQbiX1NPOsM7NK/5KPfu4vxfdM1YhU9
Deh2B7CZClFrFfGE8n4jBulQncP+oTRlUDUe4XdKQaw8y3+jpYrLi+1gDKt2zGui
/Ic2JfM6h0FOEgfCrF/uavtmBVifcjY8OIuPlwv9YW5wDYXRJCLncyvyRKY24lvb
hrKy9KloGhiFS8CI3RCVeWcVHupDiLYr/JZDDntzUnT9qA7YvEFd68C+eNZ4vXfy
FkWJZbbcd4csHO4n9p4qO6q91TFc5LpOix9wuUhTKz+Hv8PwSv0G8Qmh97wYtK6t
s5ievCRrOZ8ZHYKBSTeEIZkA/2obKU1VZbx4S3mIawbDGW/ejYFo/ot70zTqwVYC
JQqYsbSEpfH5FmmAFda2VpYzUc2SUymkqCe5HicxfwMXMUjLJbkkAGZlzGUXZlJe
jjxZDNU+iN4MK3+BlTjHkhEvoISvWIPOmXYfk6VnWKkDmqlocpyomoLw5NFcbRqK
2RiUFZhxGdTWnSvYntusFeBhaKwWWgpS+eRjkdOA5JxWU6fAKMwvhdyBj0hcL41A
HoOQ+2jo0YPz5v7/TEeT37JViC/ID/MHZKl7iBsRzqHTfSJ9557nIDlIV7Fae8oY
63vjDt/tWkF1Q/WqhyBwOjMiq5xtPeXW3HvAecCcMJNPY5xVJYEC2nt2w5Lwgegy
tGVEkaECgpnGOzTd09AntP4e0uRMuRCvfLLakQ/FFppNHz5RDQ/eCYvV+qJ3tjDa
IGKUYlanNa7hYcuRSU/Whe1hpLcI1/vah8gVP35JacBOlu9it6hmyOTamf4TwKut
7VDnH3VBycUizDeMVCLjuj/NJ/rRspq9ZqeHkrCEGycCfgb+2eJkxohEFVPjMd5H
JNu1emy+y6/Akeb6kVP1lDOC34IVtlb86W/cX4G9cbDOqopzxzkond9IrIxFjZ/6
uIR8ZKYhRGMGw07OOb1XOqV9ebmnylCpJ0R1sdNVE1mfZ1xyLsbu0DmjW1tfriJD
JUx8KFtYANpFAsWXwISJuMf6LNhNrFrVVjHJDMzRRdU234LulwyNjhWR2Wtw0MN/
G+qPA8/xCDOGuSFhRS7euaiHcK7LiORY0qM8yM0KcznQYqRYLvcjDXQ2Sv+kbDkP
r9e54MknkI9t2v6v69ByWSfHcOO3QQ5zGQO7jyIeaC0SGkMRlXDNZ9rrATdTtf8t
HwrJjpF60OCoQJonD1EmoZQkg/ZSgramMt/vw+1DiLkZe1PHNvyQtfdudGqA74Ie
tKdsQ3n7q2/ycJci4XGYLCNdPF4V3weYewWKtnh5I2G0o6DOb0U3dSB5zgmRN1AG
n09rSBrTd8fc+DoIZEJZpsO1IXygjFFzbEKSLRn6bm7n3xjchheSd371MR4+CKeN
pd060wWa6v2afruMr9gPsqCfuJhYTeyD6CCp2e7XVUryNNVGA591YQIjfsDb7JUj
U9BJkC7P/x/M+pzxHeEaX9q4ythN4vBezzsiGsiLTUlz6VX6AvrYmgTc8ExIBvAP
s91mJlOfMWIjwQK7GRqYOVhXs9MPztSBsjZyp6UY3+tJaHRhdeG9H0cNcR6RLZtP
z23oXboVbe3aTXg/JL1a+OyqsTw60+xHgZqAhDrqZ/s6a8cQJu4lFcaaWpwZRV0V
+IfuN0eAtWZLjAtVu1MHhQYKjtwS+H9JbQeAIVxwh3b9HKKoqLQQjkKYj23yG+no
Xuu1Vkg0oVXImG+i4O+xxThMmwh0Fnpw0ZUkiJwsYw9cf0KLDZdg32CtngQI7ATl
13VJ59ez8txarAL1DuaEQngiVPo4FcNdqvbV6Hxu1Y3bd8u6IPNGQNzjidahlj4T
KsnsBQiLkbhHGv0Ye3NIvbz5QooSpZc51iJ0wP5MsMBsPL8aRRRDO/YKZiKYG9Px
iXL3cf+QzW44kyv0XbBMBMDYPwtR2SBW+T9I4QCB/NyQrMjbYSKP5IXC+h5SROd/
nRM73yB6E8b6/9sBvIvJjrsAwydJqbKFjv+/sSx2ykYT58JUGzmI+xxRqueemhck
hwThNgD7k+KeUNJk1egLB2YdH6zpeyQJJZ6I/yO5l6FdYs3dl1MMxjPMjd3VxS5E
arlPlum4hmx2CcThJJvReGmBu69SIbszj1B9GV4ZiAay37AFdEHh0munuSqXA68Q
RRUvGEVDNh89JNkZ4GRr0l2SXxDUKEJoAh5HgWUdhGeJerJaqBzRMzPd9gNaxH+b
nhTwySHvXkhYJGqwL6UjFNMdyXRzfTTZP0INY1ksh3w1Nsx1yNl1W5Yr7du0Qrza
qx6fAmYh0PdRgcgq8v2Hmfy/YEJNBYUsmEY2RIagXkHNN0eqv8itG3UAVD8D6dSd
4dkHWlszChoh0WqtsPR6PlxfHJzkRFLWqXes1QBjc2GEH+ciupw9w6Qey9Pn8A3v
Za509BhqbTLx6a5wTdmLClUFYzWxUJKqktiH3nO0zbjoeJit59M/mPytPyob/JOS
1UsmW4/bR11RUCr8743NM/B/XdbHh2IhljBLZODLyuvR6p0inX2/U4Zqt8ju3uIb
gmAg+39vu3y02lhwDkBbXBZg5wRG7cHpwhCWRLDEg52mso5aL7y4jzof+Qj9/2kT
lX45JQV8rfdUIvzP5ggIk8FO7Isr4sCGAQz7+++tAU4EZcOMkaNZr2LPdeOi46Gy
yMHKUqorP6dtJWlIpmM21luQsShoWqoRqMe/abHQ1PLx6Zx7dCj4oCZAhDcFLByR
3CZ1M6wRA2O38XAXYkHVHNEi9NGwI5sJIi3kZFo5qzTBytTNdYJ0ROpgr4Z3iaHy
i1/FgYzRwt5mCecn3icZFruEYR6oKfmpxhyZphmbEky98cWSeyn8BMu8Msy9oM3Q
C0kzm1MgfyCQCtg6TEjHG8nY6Xsx3o5g0JMio19y0aYD8rfT6C6pEch7pvrNiPso
gPU8wFpTUb5ymXn7dgykZbe51jgXfq/AiU3pLH09RyyiYYGRVwUIxdhtBWJPfmpI
LOXZ7sTay20e/EU6JAKUh+gDAlUsTPWUS1ZIOFlkOwzfBwWTYMPIgDiKPoJ+dSjt
o3zSUr4WInwDZQQ6qBut6VSWxIyIyzK7VepWuMWfCQEz/GqP+8qngG5n7Iv4PmNj
x/AubFcC4zOjnPdTj4umycxpL3Hj9OFCnRNrOlYz0b6suHGYUfVdyrpuiqf6puyc
Ks0MU/ONlDUtMArVr9425I/cyYR6IAFxXsNFDagCsxqZo+pQXIBHo5nKeqdgmcus
HcD0toojiAj8iujKpBPMsNzRdVIa6uYO7QBYZqngNq+ZvzqoiEKcxFhPN1z20hfx
RvmqQSPv5V2mdAHOYRDrvqC2IPbE7N1OBLNIBYl8DwSGD1U31ql3BZ/buZKDHCZ5
GyfXqm6fGqIKTNJaPyAdtqpI6cGrx790bIpwFg/jJab49KFTF+FIT5ydNggXkhT8
RORWNv2NreJhceSwuji9DEW1Wi944MAAtFvsdvApR3woL7YjShNL7DDAVrZscFM0
Y4C6BDC7opAdN6pwqdDCXKG/w394cwE0uvSuayry60qMG34YCMqLe8zZmZ7lD0eN
z8ulkPklxzVV2Z4Okx7rSAoUWcuGlOhi4vkoDzcqrNgVwzvZOlkflUaIWCQBIDyg
dKPDlvascbTz8p0ISa98gtCf4lPWSp1liME/FBrmvCsjc3r+7JVf6WfUyCBkNDA8
uDXee4M1XgdQbZQ9RzlhlfJr1SnV3AF9Swj22FcyrYway2KFO4QG2K3KEKXiH81s
7VAoVdGXda0zwHyTdZm43PVnAbbgI9Udj5DHOlkvrRUCHKkLaBSk7Rsb9FSfa1AK
YdURdYysVWnOPSfSkEyuISl9ya9lbndBQ+MkbIBtjnV2WtX1otdTHGlTlnDWZZFD
FHk1ZlF7KPglpS80Ab2Wgegio1i/F3gTcxU2QNnWk96F1u/pkdwnahQ2Gx160kfY
98oZea9RSBylyVn5HclfydCJJgFBckx7+N5EMwswxitYIiUqUchYpOZ0ST6yzmnG
OAj32IPoYBzU4QRSxQHt1uA8+OYYwEK9g04Ka4k/LOKRWww9JE8v1K0u5PsJ3ZC5
8FZjq12Nyw1WjLg8218bkP08gbyQ9Gl3D8plcR+NJ+zVwsTVD/UWxm7/+vEO9FVk
V87NRPpTT6+B7kAODMy1AJSslLMVz5rogy9XkQ9CFYcfx9ood6PnI5hjCti91gkQ
q+DveDSkACycY7QW2zYWoj83LhtpTeNRs8NSND/HYcIiKGYgfgP86X4L7mvyLcP7
d7qFVWxKODrR9CW83HVM4cJ5It/Lf3PCySIHrJJzxFBEYhhxS8qXwG12Q+yOTTL9
J8e1/O+XCjQxysM9q1O86zkGlI8ZUoSAgPXdBvEquVW4GwLF2g9SHpCPmmnMjxOz
hwd3kh9QUtV8SoX8UtcXdArSa11p1/v0euBBkI3yXK28obV0VSLKNIjD/UG+Y2WS
bE3gXAdGh40BZqWCV3YPBfGlF2Uxu49RGthkXF26BgNNhcZLDFcP/UxJCO4HTCtZ
w/bSV5JWWNZqfUyVwoJBMWDBof3Ceqn12kCNymcNoPHEZm4Q1iUBYTJYOsk3iOSm
Kx+Vn5q84kfGDcqEeqlZP4kQBGcVwm+0f4DVCx2bzW4t4GGmBQtkxweK64Gbn4YK
2QhnlulE8ju2yxyCCJ2eDn6IQiHm08ElqJxA0OXJqEoGc7TVBA/wAlAVw8Sdh2EN
4jVRwohwHcd1NmGcA2cVUe5Co9ks6ZnDXxUTZmNC7fBg/MWoyOiOuMEL6U+WELj3
HZ8nPyLsioupxql4SvCFHl7nEFzwIuiMkUnTFxsNlV15k0cSuUwm3dNHTjVgvEee
ic+QKcbU7Yy9MIl/RLnZW00lgyWHoOQz/FX7LFXWlC4QouwhpFPg5vH9/Wc6DWPV
fHEtgpsPoIVPlfSaQq4rwP7eDPxDPo8Fk8AqZSx5frSDSXi30iKbGD24/uzSvC/E
a9aux4XUE3cLA7B6t3Uj0ALljz22vUdNEMO0/PGjiJQ3XiiM7DVE0kASuwN1xghf
aKo3r2nWOnzz/uI/47Wh6fjU6B5f/VlsTerak220m2WpDwl6dfe5+5+DHdRnmvNS
LH+BEcgpZMeWCu82+tKk1QI6d2ZgyrhdA4J34OCv5C39wWBYV/G7rF+8UN7FOtB7
kXkzWDJRlO4sOTqJyD/UISbIkLiwHWGpTV5emxU6wSn5FGtD9derAD2Ctm98zVaj
jCw8//BmmStGrGAptQedAjdFzB2VsXq9c7hBrQ5VCvAsA86jZNGTZ7NwlMFJj+WV
QANdqflDzTVaId+2T7RAWH/C78DGSAG6+3Fufsi4efBwyU/ZYv99vw1ZS/0jTo6i
AEjolZ0koU5Dv2AgQgNKbwdflfEePcf8V5jxyjOi1VUabjsFnTVz0iZ9umFVLwZ+
ov3trDpyZiw/5Zxq5ur2w4WhvvgmOdZ8fOJkOQ0E/116vufpo3VXXKnM0+zvcpL8
l7oztdGzPPhDQF9U2xrtuaubKToIrNpD8Uc/BjUXaatgsl0T44aDmwlC7qgWX+hH
iET8gjG6zkOqI6Va+QXdtkEJLjRsOfOFn7HkZd3klNT/8m9MiupaTT/Bzv75JZrl
lwqljYc2T/hSthIUPt8G9QVS2CZ/XOrKbOV4HQ9u8E2V9zu1Hf3tE/hli6ZIenRY
Stj0yRzzYRySB5Yt/P/Q+nyf005JDnrkEVRkyhPkXMXfjOYDkScM+YbTm8cqz6iS
q3XYIOqTAuESUdL6p/RUXudIY1Ey9uLzqP4MVahJ6KpbR33UY+5kGOT3GVaVr02u
SYCA+zBiC2/AsI4KhOtOyNPSkyUYfpywY6y8pZTG1UwyUfgPodMnY639iiYHC+4U
l63pDSGFWp6/24jYcGSZlJ87MFufhV72DuJ3BeMNugLpCSg1emOpJvKesW1NAp6k
7tRyIrTAnBDm9DdU0Rh+ekCOYxnMOc37VHtv+KmBORug2nyhu1tQ+C7WnHVw355V
eOJlHR8GrA7aJj9YKj1qE+ejWGnPmGXOpGfDo/NBm1r276qrK42PnZibrKcGB82k
avTfv3iuDcK7vHVNc3qT26omAghEMT+Jqpzv7gjub8INPk6kj7vjo9Evkzwomecu
BZYVcG9iFj+BmMka8ZoRfRYjxzfWXtSG7g40+7qXGBzBkeqE4v7RmIRO/Z2MjF3l
7QroomCiYs1xjQFLP8NQCSOpUlmEwid7pGqesO9BBObRPzFX85pPpsA8jdumrdwZ
fjKq18kQbC52zii/UJcqA/gHjrcDYRRbLX1lWrea/l6fusPzPF392ZBBd6OBd+jA
uCUKiNaNTwsphxI/jWYyFJWhF+hW2KTL8dDiPkdQHLvO73m8/ncIITH2vtjkvL/A
VZ8MUY5/9WyFqB3429eO1jO5hYjNZJFPZPbu4QsAj6xaEik1EiDZsQbTtWm0NQFP
6iviMmsWd2ZqbzVHTcQ5d+SK4EY8KfSVagqGRf82M11vWGE9UWNdv9vHk9IALWGG
uvUXEPQ4/xGLYu4wkq/v3LUU3kDNNnF5E5LGy4x8EIT37d7HgU8MUeGegg9+LN4D
lOU1XKD+nXVPpcWlrLTZhmlDjkm14OFQdehaGYc/CEtz/ypXkDsJXnr1K9HH+w0/
bYg619gVaxD++OdkPYAraSo1AVH9LT54AHuHNuiOiKn6aP3M0DAj2i9J+Q3bK7MO
4cyQ96Ll4OwLomviOhbVflGC3DXLPSxjIE8fAOX6+vxY9Dw/rhJFrA0EqceJtBrh
/QxMN48lzERUi94etclbpdvt/qHK8zJ2ysy08OQBfQmVU2T18IVvXGQ2H7pgScEH
JECt/s1jbYB8wkqy4OCG13Dmi+YXCAzXJ6ziiIyPxkWApX9HB8feJ0kNk7Ou5NAO
hK/LfKOieo9MbQf3mtaj5YsKMbBaHZyuwILoW50Npvz6xmE5FEz6FWL5oiEafeHx
KUYBqJmh/IpsTT0ZyA2vmMbQp6+1gju0DI1bE7tbZhyg8MF/CZe3bJzga6nfoHXY
2vCt7WPI5YeGoi/CzE4ccZr9ktTKH5TOoWW9MK9shFGFHSqGXPBYQ0FXAcQogN/M
KWNCh57jjsnTbpjUkq8YtmiLSTs/6ZhB4YwTutjQrRabAM+Ndv33dUkYj5vYZDFd
vtC71mFf2VfJfPFjY/InuWAg0CYM8DXJJ7gIL6p4eGIkzNXEO9K2qsSbyvh/QRSu
pBkuESoJpuGQobbXJ3T5H42BEIRk+SPznktldpmNnbY7nb0hacsa7SStTg8WbxrY
G2wpcy/qKg59YbuIjYMdF/Q3DI7o84Vk9zgmdc22WqyQvUYR9ska7vjtutqkTQ0w
VOnVFxMEPoJj/L7PebBSb9+7usGdTc6tQvCI+bery2t8pz6AyugyocTHgayFSrN/
lHjdTlj8c4rOovRNuXw7GCIWsTFZ71+GwNuska28Q2aGzfdIvGp69TVnR28r6ZIB
LnG5xUQAQz+z1yJTCzNQn72S0LyCGg4MExWjc8sZpLi4Bt69TfssdwF5fOrZNvQf
WlJ8PhdV3iM2T7vNm02p5ZjyCYINYswuIEzdVxm3xp2Tkq12JivG6e1yq5Pkmbeu
C1bxGlREB8V1NxuVflphuqJ+iXHL52l6OWg0nWp2pmDyZQIKAYHmfz7G0x00leLZ
uOWCJRKQm9IuWo30LXPXC5fiThxn91E1873IxIVTrTMU5hivREnbYQ+lZJX8UT1D
mdaBqAtInVtLiVrafUWzBKKH7eCCkp0bxuYcbmhUNtpNh+Z2XYT/qGUze8o1YKb1
nCLO9bNIfTfUjIw3ZkGad9i4GDS9WbW9gwXYGLbmTOoCw5sphZRjgsknSHrh2cs5
+vlMkiIwGNcFCdE3gN9EUH0dIy6/gkMprWtMUH/4lm8cidIj0wczPv2CgS73yzHm
1h7Mf8twLPloTx5Js6QP2EUh2afqW7aOHzDmEd3G38QQjzI2IHoyHu++qxcMfOED
3j0TZ/GVykJewnBUPUmSRNUoiFnCe+M3NpkogY5sHESleK2JN0ikE/GdwPXJx/Sg
n+/LOvZB44Y+P0U9GMtronuej3lLipAPhpE6yCkyOMcT+tXqsRMQVi1adEh9/lD/
A9MUUwUahK0FYbxxyRhnhFn8G1rjgwc8rj2x1N0m9ceV2VUXiVRcauTMb273vxGF
hi/UuWbseyrooaT1EbbPPsj0P8NQM88fCPE3tGdlmMqvxBC/6i/RdrD2M8W+KwJk
wI5Q/tUZoi0Hqr0DNt/kQuYibJWdfnxBQgtQw8jgNNNd/D/KNZHDdi225a9nDH1G
Uq7LYODgsNokINYpm+/J3APT5CDxfNbJJvIaRaXoiyf+W+xMiWNfGoxNTiO07ukf
8VV+HDymEMjNTLIptWxKzQ5WX+2DwkGc240whFp8DOTo3MTt5Gk8ZaAZYp/2o1s3
b6s7bVcH8E/xanyl7GYMo/66t5mf4COzDYsXJkPTIZB30Ohr7J3qgfFc1tniZtaL
yFInVgm8nioXOPgGNVlI7Zbm2Qw3tP7itOASbXpxlQ3g/GhAe/oMf7Ps37xpRh8q
esV2zprzhqcY8kG3LR4+qus+ifwQ/w2M81BzNudZYh21z5/5vAfkkMW/njCaOmNR
JW3b37nNJlACJmM6qsm4dxD0F5eigdXckg5zDou1Qge8ony/3mkX15YcIP9NMAzf
FHYE2lbedT4kKU7rwdoNLfsOQ0kEG3HxNhSbGttG/G706kN5btpiVdrM+Z06Fh9+
ZsVTjMAB+T7fAZhAAOtZHp1EjWGrhaxqDMG519asT6AtBbPW4N319KwZEPcBtfun
AFSprYK5sgnIv9LRygNNQrxZlduCYf8DJ8h53LzHQNYetlha7nMNMDgFyjJb9k9o
eMSYd2mrzIr0XIKTbPCRL3vDO/JfU44DYjP6Ht57YxIsul3eDZl3ZXuwI8AiUneS
yZX8p/McdoTbM8j792ZL2YJA7CZCzwg60jIqkqklHbsh6LEz2sKXB5TCkbBh7+kr
LOB5WpaTejLO0ZoHx21Tll8RgJWrsnuIeAYWBpSS/PUZ+o96r3EjeEaaA7aj3SVV
x8oUFzpinlSq97KdCsiO6OtofYzuONvl/7PDmFM+VE8WVwrE+lu8GqS+99UMwumR
h8kYxYtAeMZ8HhBSgQxObPiZYtqvBRlCztNvl9VXRrKRLWCSSS6AtyAOAagRxoOZ
HJlXanSHLGZlRAED8MmuPT8OF7sSnqe/cTm8HLPqflBx/A65Rd2jhTLhOI5P9Aw4
7Q/aHbCeNXEc2gyNvc+pwyv3OneXWbYn+6/Bp/M0GtdflbVf7EivvCJxDpwBtkmv
WJp84A+zA+zIvvEE0hsZEHV6r9o4FXGkxsGQtgxOXvXYAsqNb0emX373SlD2M2T4
DcoTmc5TKL/odke7UyMNmrpeklu7lzpShpzH7241Z3d9ZndatEGZfqB+606LLVAa
pILIUseDVNojnAaUzo8fR0FGz7MqKxKKhW6X6yf8STogzxnEoeRCg/QxNSLhBWCB
5+GTmf9jAHh9cCw6KYO0Uu2Zul+PVhpxx0gzHKc5HJXiWtfImYGZJ433TTRmD2Cq
euBURQvNEW6u+epZ+g3vL7uFxscVtdBKiCWlCexQMpg+Fd1GFAYNGbw5OywEM22I
yNI2MCbe3TNi47Ly7pE81hZBuLQOLNWEQG6z4KlZN1tmrsTLDmHRs0hzR+PWFsOj
sT7Jh1Pg2ZgjuKIrRRy0LTIoqGxlbEgoWLztrjfra3wNxmy4qOVl/bic/F7UpLt3
SUlnjjr7qSvBOTD4YULegRfjwojosvqXF47alMIayNIfEAxZUZngKWCN6LMRU2ET
JIK/XUXtS8L0NlDgldwjn6iAJVtnBqrJc5gs/s4BENKNziUqMlPGHyzuc+iahdLL
vxVtV5RdlaedFlwtv0BKM7Uk4jgFHq0UAGhGpdksYKuj6TwsrnJAZotHvGqkvdUb
lYoQR9dRQQ/dZwFiPyvEjuiQ1/ZheqY1NI2SaTVum8khQjk8rsfvOurWwCcWsZZ5
rvIeNyVvdXDy6ujguqOsvYPFwYg9/EZ6OQdhKxLp+IICpULR8TqvUpNHVoOV9uNP
okzu4Ium5s2Td6Pbeq4ZctE6EWGjVXlhHTat+9b92GCnMXAF6zerhFtAZ1ZCGmC1
DCW2a5apl/BngB86n/JbwkKyGtOXm5TiDuQ99f2aGxFUeFJs9RWBw75el3mIiFB1
rUCSjOvQW3dJpHmF62Nxq5b0jB838cuJirEdSubZcHl8JQv53nLlB7axZVuo3f9O
gjchx0EAXRcSoNmnrt/iwzSTP1ccreuz4c32tR6fJs401/mDxnsca/2qKp++3TsJ
+dSvnD764Gk+eri79IeohMn92dFGoaeyIo+UExhe+I9ouBU69LrZxqS9KljqdEsV
AZj/+xHUEKtySLCF3PFCXs1jDTNiFM4w7FYTZqaLkTtzrCRC95ZZUy1+LjgV33tp
Q76BcEyGs9LUWR4mthb5q0aP5iasOPtLPVtgKa8EOwgVBvs7RHJFP6jxC51/UbVI
0HpLdByk69IRngPqxgoeQR5cLS9Sz6r29DxxdwsElwAv4fU4FpdSYZeW/Pw1qNSZ
4dAd/cIP2g0cNUomKBN81RX23sxQkJJOOUlx1YkPTh2OtYn9yHGI/RQr2xTSQ3O+
taBM6F6cDqRtL8+/W/nVxz9h9o+Kr0iCfmdjgda0XSBlBg23ciIzRMD/IXF3ZRSw
zjUCgNloQPN+Z2kWgvfQZ7apfOm3v5YWQRkoAmmgM2IJk80Dal48sD++KHtfUC+o
ARkv+gk16kry5n1qm7v6gF7KMC2QMZj0z1WySvfCZ58FXd+CsJ+++s/rX8VnJEZ1
z8tBi7nSn/9tEk2JfB9WX5qccrJ01yAXqQpYSrQX9rYeYMTZjekZdENEggijb8Ef
BzrjougrfIftfjWWqC7xheNQCxkDYhjCpI1/ksHQrGp7fN7uliE1OQ2GOlBzGxjf
E5bzGKIPgUWsEA0taCOW3V6iPBF2suSE2L8/6CeiBYGEIDpRaZwmXhsM7hD9cGa9
EOH6bYao51yIxK1UBRr8DJjj6AeAkkq/IsTFQD89206ekT9WRGB+QTAhpwmkdy9K
jESSnxzL8d0PR4Fv/Rbsw8AmedFFl51dq8AaU9YN02by8+0pqhoQ/uVBFjRRmJgf
BhXuBBZKH2grU3vY83EhE8GO8vSfuvXmQh0fvHRZPpt/sb6elwWx08/AtofgGWhM
1QHhGl1j9hzw/ll+GHzqrSBfcXDrRHx8VrLg7KHNTNj3mE4OY0dHHx0cHevApY9c
ui5TQ9Z2S1ZDShQrBHvmjj9zJpCPNXI9G/q8ki/IkNlUnhMK++EXYT7qT9/sov4B
6GHGa+xoolF3OoAQkeEzxMTRTc5fxTAZ9h8E2rcdS4O2kdiMzYCG0NlXoerAmJU9
Wt4kDVQ1hJIHuoQCMVe7tGZLPYkcKjxGPEPitoxfOTAKFo5anYZJaEIsqki6ekbz
YN7MLN33AKc9qu3u9Fda1hFBQGqWa+DlAo8deZ9v6OTIcAr/qTQiLgN0sD9WdcT3
e2GA7Cqdux7Ion/yUPAMJlK3rsEpW3ocYz+nSRDdItkhS9ux2mgm9VxSc4kcgthP
05iXXXUuNTVWctUL0UuMh0PobjyIpWdlZb08N6gIxrzgEN7v7/lyXMJQ7sf2G77b
ZMCrfChf8cSJGrmNJMbdGXVrJ9PNPpPj3Q0DFxiQjV0NMPlB90fYtJHIhzQw1o9n
bWMtwYTYIYg0fZj2JwxavMA0+c6ET9OaaIhMSaUoMsECfEw8B6+QN6pEvuNkSxoc
Lx8xjUIEE77e2hYoLPSe0Yq+768NPHM1v9NXcVqp5B5Ec89lhvE5WujLdlXeeOMM
KgoYY3OCO6I+rLAOP1Y9y7gFDedzBv8DMpNARiwMDlIDdyqUEjh62Gx1OUeAg3kQ
5fGgVe36IYADKHmNKpZkvlgvOP/XUKBkUtZmn8CgUZjw8BOdsz3z2UbtqJ7fTdHr
xS60rA6qmWBTejkAeaOy8fZtCNUoTUj/Vev+gHDC2Uw6mhqUFc9mFiDd1lEpHQW5
kaMB7bXwnLS4Ly3oOOsX8fwv9DZmgWX0lUBgIQqjyKi4cir+o8SM4zH+I9Vexh82
UvJf1S/iBImBNZiMbZwzuqga8d5jmzDpyrINaKzhYGTscKOubyre4k+59Z0EgFzF
7wzuwNmzRDUFavLZ9CcUjNWZDol9XffwosGJN1ICLft7FDc5JmIJA/EaUnkXbGQL
NVaRNvcBYBvTbpC4hgslwQy+ckY4r+vhHD1GeG1rFmRJTUil3wHqBYV80Q1KS+Tn
uoo0E7fz0yuBhZRJkcp19uvdinZdQTQEmAZwR0caLpXFFeQcQ8gQs1qY1EpO8rBk
qTQNkXPjvrtfsYQce6qVg4UVxqsYxq+hSGd8IL8dCAQPSv1JvSYzruCEH6NnEYab
vCm1eIls0jRXt9vUvbbIjGH5VlIh90mi2QdZ8Cs/8rH1D5EJeYzlPj6XcRu383fn
yNTLEdj4gtFbM+ily2N+zzEfMQzTJIhyBUlwV003Lt/06f5zAeO5SkcNf/838XjZ
/4/WhYxZ/tLvqY0xy5fV7wwW4/ojCHAVXRcqWr00zTEUJqXTcIZr0/UVArFyWquT
C5evfjGLg1JDhznetP6Zq7GTCUL/bcyc/MyHVRn1mqHndt+PKCwXwGWLCsmaO177
rGSAiKMqZhSfS6ypLriRwfgbAEFtK1UB1gcoUqsV1Fc0qIwIgBIHrThMGPJ36NMa
r4SNsRafYClKYMz18SDakF4opVaOab3KjDQEQEHaCmtxywGEgOCT5C32mxJ46FCO
1A2TWwhkjnwZMoyjCiSbOh8+NRKgov1PugdLF7g7705vd8zIldJzYV6+ZahxWXnz
2oagHIBYwVS0jBgh5zJEAKqd7c2FpVWChlbPeco8G2g4tZIBHR3AeY/s7O/1CcbF
rWHC4G+6UkNBf4ds1BzNFQyFRdlwIUI6KrAWjipzNU8mJfD+hptfVGfctJtgPhDw
i7/ulGMpSmJqBAqqZOa17JQdSdtimyOxLZVeNFl7RNv+5MiRL+K+fOiX6U4DWLWp
CJ16nA5BM7iu4cX262PMZYIgEWCWZxg888XHUCiR00iMn7yoMSlDBa+QOf2fmF5p
XUccr0AkYTlxLFyCAKDYWa0vZo9T7d3Eag3U7961ZG5EIRZoLdubkTefCRoLrSqe
YoRW2Xj5F8dAsW+rHMMphSZkghUOzZGGfxBbCBzXI2M+ZhZqCwJo8mV7VnAqRRwM
f6kKbJ4G5FXUBHvhkSlShUNO9bZd84Do1Uop7CrTKFqtHhIXfTpdtLfA1dOjD4Lx
hNiuHDZiLBC5QSrZyREybJXvQoWWNiDSS7yq2cV8zd8k3D7lcfD/MIya8w+QqZpC
dhLKJZkumVTKpCLF8V6DxRb2JdXsFNgJYBsppPUVEC/ugp1ypVhhjc7iQf+u34ES
3SygqAotN7m3nQz5rYs3Fre1d4eDtbBQM81wY6ckN9MYqOil3X9lyHVYKEFh+lTQ
pjZjuCbF8CT0aXG0MQJD9ejvr61ebZkgbR0W0aRgeabv6d8Cz0rWzCEFGmJLPMVX
SUuYmyMSiuUVNWIDHhMmUh8Xv9fwlyKU2e0z7EygNFGLYUtQetlZmLW71YHzqUXy
tnLUNHPwHAMXVaRWvR3Ji8/uHjfAbs6M/Cdtbo5Tq2JNhobLiiFZNmupF+s1zYte
vUSDpaQfRb78MJq9/i/XodMEknRnXBJtKDxrGrX8RMP0+h6UAJX9j+NQmb2Zc9rL
7s7vRZXTr+wGzsLyAs4Haua2qMHLKP2MQfOTICdBMivUAo4uDaEir8WXE2aJqPLl
KJ7XCfa8v11CGa4i52DqQ21Wtpyb9rJls0w2rpLhP3GA5pFIYMFlX98jsXlpab7v
GQkUfMiiyw5LRlrWYqJBlmLQPZyVwqs4kPtTx1wO3CnkLHZPvKh+yjnsb+ZLFp/X
59wcWdoS1JWnAh2BSk0ZAPnXcUQwmbsyI+Y/yyV4i2oI8OxtrGCjMUsG80n/bSZ3
nuxQC1+QKJTOR7O/fVOp1CsbbHZEIGfcdwM+bK5R/XCAvKUrWvYwtXXI5sqqAVfc
VmydRlI69qKY0tVmwT/MxD3hj4qiemV0orVBPnx6Q8GggsZJuCobIWgEt+n2/JEX
1Y2COrPdaLA1wHdtfzhgtK+xDhKvPz6GNO9q2ONXViNGD+62HF4xbYVwIkXzPMKs
mcMSHR/0wNFac7jKmAqomuQDXYsPhTQxyoH9UVEGDt0AYwknMhxjsFn26ea8yO59
iuGqGnQppt8JbpKtWTwbT6HUX3idhRBwNg+wALvccMWLT+nVB99TYsGjLiJH/yq/
3XD8zpqFP77wENeBAWjLeaaO/mSmgZ631Zwz6djC75ZoiRDoIjzk1W+hVbrPHCoN
2WdcxJuCHPuIQwDbArtYfkQPzEshvEQeKNlO9wG8y3ZoqXvuhg7xzyhXVGWsysZB
yWZvUnckriIlpx+bslseeZhS08iGUZYEM10UGDgYY0eXWQM3/1wWJ/U5H/bS1v8p
bwt4FVGyGLnbSc182PGYNaGDjKwUUHl4Jhmha8jF8ZcEW0RBbPECOdTxULW99e0n
T1Trb6QQj466W24AG+Pg6PojUsi8+Huol1By+J/mnNaVX93lC6k60kJsaO9WaMEu
AGG1DVNClnWQgA3bb8IH82re09YFDtoC4/404rmQwJKv6SLbAzO0ePEiXc1DopzN
IJW88b4/sua0Sn2/vMIN/Ev/qIu4+yzLJDayMsRStBu2l2vPmLGl5/nXPb8a8OaZ
jPWrE0xXxdSRzBZ7qZ5EM53hZyuKSDFxkhu4SBTyHeVgoy3Zya/cxdexq4/SkZIP
ChOUwDQkpgImkKXaBjVZfhcSbpeOW9tjX7JlPhDHohLAJNKQoFxV2vieEPhHCepG
SB+J/j3ep68/XNI5jqExRlxm3+gnvF1PQmoakLV6J54L8/4zW3KCAhg7psjnHaaV
1GlzguL2wIOcMqnwlCjkWkEOqvuAtJSYrjW069dBMUv8yN/zApMADjvKHiEX1JQf
+6Lhi+EMmk4zqR+N6F2SHcHt0TgOfucXe7k0eJ5Upoqh6VPyIQ+HoSQ31HFQoi+U
aWQzzV+IqEG2ztEiFJlfi+dqsRhI+n6ywZ+i+T3912Gmaj0zw2qjXa4LkuiaHPlH
XUH3+IQQbAGbLXx8UAauNWUrkWBGpT9H/wVcgqQSfsexrdIIO7l+DHXzpDPnxDIr
0unnzPUm8meaEGVXh0I/CvYiC4UJZmFUO4W152EWLWp44RgjBdP8VhUWSMsmmXAK
FcJrO/i1+nNn/UdN+hPtD8GCGuRHnzxepwwf/IvyWDqqkArsCl/H5SNZnoLSj4sB
+uV219CTVKtvsW2AQx65Nu5Nd+z3IHTf3WrjKHLlLlj1rR1MVvK3m3mMkBwICAoT
YOiZObSLloNy5CRd9Me8BbU5Lk3wKRKH0jV1t43QcWjtmJCO4REltI6EVY7ue8/D
2teoZHMrfPO5RIAFW5m7VWjjFsAezCu3Ugld0l0SBPf4g+8+GPhfMXumPd8mBv7F
uxAnJJhccYFu1xXmA1wYtDqS9V/pvlTwY4ig9/yfSJDlwmuDEAtOKmki0Hs5gSlt
e8sxgTwiEDlZ4t4PsZik/RVAouxQFTPPZOugxB83vCxq2hmoIjT0xoHbtrcHiDCo
38/+0QqKK8mZJLG1/oO3hxNUGFSnZWk7rHt+N/RNNAaQf36s8Q0O9YzJ1dMbYqdy
08fbvPgT5+8g51kaf7kQ84jxCxDp3GrMP+Igdqzihj3ckcg2EKMN+RTCcrd0UK/3
QIS2wct5ZI3ZhSlGa4OpEWsIJSXDyJKxNKHS9TK6rY8Lo/B3d3df58HPMqMcjI1v
qE+iWVI4UTj5Tn+A235P4Aszunc9pefw9ttZMH56R71viGktcB+afkXFDwB8uFmu
BE/eCnNXIBcmTuyxmuBohWf3dsccOgin0AssqpcOt5hEpGzmtX3NiXMbwmcgeEVe
hyrtA1WufmwkbPydvQrXhrFczQxU08C98XLC6NaqMnQm372ChaOPqM2YVqMDDMvp
YHr2BxdFE9jCCJUIugPFPD/9r+jYoIQIQRN7dY8VzFUMukZiP1MBBgCrk8ZOtxg4
St4HYsR4rq8WeWRfuWuiXEzitLeUxZ+fxzgz7PLb5aY1AnWAybVnRvA3wnDvm+d+
jTsM0kfxRK8tys6SP8pP5Imdctc2ZnKDqUiIsJc4uxwHHyJqIv/LOpvq1Y6qbngm
+oBQF70JLCAKKVKQxqJDH6bQ88ILeKaIqrH3gxnDzQffs/UOMmviWxYsz329dXFs
0dhTZCsRqu6s8kIwT80Z5DPv4pGBjVi30K8WJw2y7w55Mcih138Y5P286iWznFOc
eP/K2Da1sw5jUyaxhiDPNVJCMqjeOmbmLE25w1CphJZS+dDdqlGamgertdJ6v64k
6EWA/JgFix75sddfgATokbw3k52eigQT+tM1DEbkAu6He98EHAr9h7ameQVeBNHf
QCkbskSZq2YmQqBbzlPzPZ8vUMa+BrukE1abgN4wwNv/ZiQHvvdAVzQ5LjnV/nuc
EXSy+cXYk5yVIdK62UEoz2ojLgAQOkPuzI0JHj4miLVYayXKrgid0HaUx2vcqWdP
30aFFfWzWOPDX1F/VDl7tlT5gh5RI6QOtW9pe0WOjKJYodylEB/vLN6sm6Fdkaui
9OTNrZzX9Yt15QjCjpB3oMDWQUDWTE4lfdPW84nPnXCzF4WCg9WI17MFHZh2oTIy
XN1iTHYxC7SeZU9H0KfolYx1NDAMJWecP1uBFIp4nGAVrHVkwNJCpsi1ftH2Mk3T
e6QdgmGO+17/LfUhUzY8Eu9cz6cHs8x8KjCNp4fIj3OEQlz73D0oYQeua/mYOBtF
SXmBK3J2OyFEOwshDdJ+L8+RpMR4q+YJVTjD3oAq711FaKPwkxoPBqz8vUrFiUjK
0EhVhzruP/MGTsPL5uhTpzfOq6wgB0BbAII3Ydwv611bXXM7atKSgn3VRH2ZMmXi
9TNcd/vNTCBiM83QFAJpZwZesrDlqa357DGqX4NEDZUIoq57EVlL8/ffawreoZzN
AEtCaWT8F1tj4ezbw2vQpCCBTFV7plgWhZGLZsAVxHjFMb8qrpPm5phUE73yFga2
wjZ3vuUqmCA/cRRVkUKU34VMt09vZTocnnm8BUyEarDNRMFcVYBBEgVmjlhr18Q9
uiLiQnupZR4ASie/dXCfVaRMyy4xME1hv8Sr0hpJRtWRKvFsZi0PpKEesqv19NAy
umxySTKoBK3tCGpiMBUE0UBty+oC6h2w1MagO/XC7bfmAGRf2jXwXoqA6v+0K8uR
ss5+Tmj6WsFr8g5g7GhHsxGLZXu6bFIhrdnvzinEeIOsI7bOfHvH+9xr77I3Vrfu
3nEyKIu7lonFJyNn210jAaDNcTOoiBzRSihcOIEKztxWfKJqB7uDUH/urZABFflD
lqPoTj5GysJ8qpnvtTSWmokXryRic3+VjmUJk40N+G6CMC//EnbPjBjIv+0lpIRM
sBAJAsSR+jQBG0IWPyYJcsxg0ZHxiaQR4wllOquKjhNht+9I2zWVak2B3MI4C0CG
jArNrBsxNkWtTRyNnmFLNSh1TQdpFOtG8QSppfQ2yJ60BrP3BPm72SVQRG3h29NO
jFxi6ySStaWfQxxIErbTm+vnonhZ+zbDoCF/76WRTFqiVt4Z9dL+NnW5ghjAgjfl
DFycbMoH05RIZ6oyh6iF0oGc+aY69T0IhQi2eeKi1DvIc6TJW49UznVs2BmfqtiB
/I3Tt2OzERzO/JJ/SZcWfM4ZTLoi+4b9W06e4jAZaenfP3KHLyvWzkjLAmL+BLxi
rHW7h5rjfUuNpZ5dDIrZ6jDt8jPwGEvB53RHb7MoJqQYHfSv75hJP/spAcn/q6Jc
gy2+IqOXgk6HXzFqTk73sPZL38DN7vaXoqcshhwieOqnXs3UgiJdT2IX2MXujVV6
HTOwfF7sUH8j0kuoLybim9QWhEeogpQlcCSA71Bw/gLlvEVIYa+LIqwhrzp0eM/b
vVj+Vc8qcOPG9QfsO1f3QhDazUhKTg3gzIhQBJylaEFpoJcwbOT+Uxueo7Rnksin
D35ip7t+iNaUkNh/Npfy0UHVSB2XQBFqcAGyKujeLwxkajLBrvcamMF0L3dz0B/O
Yz3oGGrH+w+rJwPQZHiNNgaliZizEBo7wXE5ybDA7wnL1CxscBvDL33ter62XSIw
fWVFfWM0kevP/ieMEjBjO9wZFkYxyPAp9F6w8UJT8wE+/4rhc4hNftddwOWujkxs
behB0WEfT0UdvkGhT49/V+fy1m5StoYgoPaTxn4kygIhxm6mLa/ZUjctZHLaL07h
xnI62KvF9mpIhBWE2IYoAqEewLCSIJTBRWAaIhwQgghwvlJ9THMAX0Tb3lgu9VU+
+f5dQ/msp/FSLLTypu/kslCGWz//saxlfjOljddhxtmhihh04tpGwnKmWC8USIjk
O05Km6qclzqVtFrdme0BN55r2QfgGoOqCkJZkYVFOlZtzCV5luI2l6c2MzObJVdl
kCmEUY1KqPPHbTSudVAE5eBUK1bsqzzCCjOwYhi2Dx0leVZpLR74axIH1xS776mb
YLLCS/TDgmY6MeRPmPoOsPzHpB/lA+1P06I1+q0g2DAM6n3dNlAynjpg5ATq7WQz
Kuq8GCpU9uHEBj4T57V1sF+0eWFQNtgMsL5E0BeD+ost68P79++RzAP1idveEtNg
KFhOqZiWqEkb4prqlPaQw5jeeXVxpp+8PyGtHRP1T63BxLgJN2NgRBqsw9xPjiFi
u9lkr1XfLLQd5QE4+9RpDD1kU+NijYf6gFdyE3x5NynQeXhLG4NGhovkveyQT1kB
q+K3T2ew3nriILqZW2tbBI+/He94A/wgeAgNy3Df+yPdKFPb+BRhVQGh/RP35SY2
nY4U8l1BVpML0w2ZocG0bF90RgR+VCEJevVXlomTQmH6it/ek8ocsM2B5i0SsV89
FbfB0XnfaXVVgnBwXSyvqH7MGVFsmFNX1P9mBFOA/y43VTMo2NiNzUgKZ2SCGdVA
cOC7MagOexsgrI6g6IvZ4Sm4jFszmm43cMS+WRHjsjsG8EuTUYh93nWWyKwW23Q3
0CbKKGGaCeA7dpEyPCX2MXMZOQ8c/90tcR5WgiAolaz8WZJ4ICCygMB0OZIALhw+
L2tkU9gDEY0Dt+7G7BJQYJt+H7+Ok5A1LjW7Ur5DVtyKXDALeq+HaV4hXQHViq1D
Kpe2SbanRgjjlzfyfLzejBza7HC64YPOcxRG1hYzNo8q1tgkMSq1CzO6wraATMsJ
mKsYkIcebOEvfWzZu4w3LiE9NMk45Fd8LqlsVktRpBl+yjec1l0w+4Z2AlNJxAYc
p26ywrfs1HkrM8zqLx/Ra/waqUWHd9k/bxR6IcLOH0c+1wDhpuUXk8Ub4vxrZ+z/
KCuRBvzHkd2QFMWwo33nltCaUov7pGZKejLwQ6cg6Iz8T4+g6FRoa3d48j4cD5EA
QuHnatRFnmq3sdhmlm+mGE/KwtDYIo+dR8Zi54WY5YowR+wV6epmQd9qvBrq8anp
adRjFIHSDKFrj40n6X9iZPCxc6GnSta94Pm9Ut8BRzq+5F/fsOSbGLwprYtJ6dsR
UYmjKjhbQyyrl25GD1RMsykm2HWoatlcWp8IHIhYAwv+TZZF29OjKpFSkov+a69B
KGwHb6L3Qv/lxDjCxN19vDPQhYkjV6ZiHeCdAJE03myQTrL3hNroglZhSB9/OQTl
ebM2M0GtrX2JW9TOgGORw0ORyrfrJOV40jaGpJIAGxIyl9py6wZrfDPLmjCnzXYq
vqN5I21AxwauzJtldp48U9ivdZju8J4CBMRUPSrL8raWxd95C1LUywMsI79Hp39o
VgR3AU7/df7Z4XwEpKABflq4YdrkLnYFTcJatW7fLvmkFh57e84zphw3U2senErW
tY/sKmGHTxEW9qAUxB9t1AzIVDzjzgLsso29Gztv3XY9eeIDJNEUOoVUx6pj+U5W
X34T3iaSXtSECUHQkkfozaggo5gdo+clliFyclM+kjkXcjSHP91DmetvEWay2IJb
J41lduzWMYttJhLfOWI2OcqeJriXPLaKC92a7b8wypMpUr4Ey+5FDUjBCZ8K4BSZ
uDU163+3zA5217Y+NNCZJiyq6WxYU0bgyaHtLLbpNTQvPPPHqPasAXYw+mKv53A8
EPeFqjtm+4TN+lUYbygfVkrloyit6p7heRu2mZ2SY+MryUSO+h6HT+gv/QJaTClL
osWrhd+aKeoFUQD2bcNSAkM2ZGH2rD8MB9/9iTteUfgiask75ije6zJWyEKawbym
XKY2agWBnZIFGjsZjxzqkZcVPHKuVz1uatoCkhLla9eXPkphTAL3ZyM+YqOpGRnd
O+Rs2BDC096KHFThvbkS+njFoCFLszXLpWJY86A6hcebfiC0Jm+50ECvTPgT+9pm
u3NG+gB/igvbDBPzsxKMXQXRKUVvKDD8hgVmAcEZpnCx4ghPuZiSOHB0/q8TbNzi
Qk8nr0MocQ9X7iL7dVTPj5mbgSJCnPAymQrvbR2ncRTO7W9Skz5Y76DzvSYZi07G
LcS30CqUPsiUwArDP3o0CrG9lsdvHJN674SgfvR8B3gqa97j5nMg4kaJJLXUwly7
gfZNquUzPGqfOISWUxg6iu3SiRf3bf48hD/w5O50sNzspU5U2MY65u8OgRkoUZZ7
ZJGn17vrCT3ibzCAWQOMmho7W9nzjKiXdrATj8VU7PzS1t7jzNiGn6LeADRtmBTp
sSd6lVQAwJ7T9hXzlxQO9hgISwGzYKFhFNrgs+Q86iD5MqBWcI6j8vpHaJ9xD+py
WZyHr8cGXFlMyir4jkjnDVcs5pMY3vWMt6gQ2CTL/IPh+qxFchuW4KIEfI39jXdX
zUQEULswcxaklJNE/5X9ZES961pYquLQXctZW9SOEHt7FJbOTGjvxCSukpEQ9CAP
SYO6Ot4HVzzOM4+wDbPn4KvXRv3fdYYfSD43xDquZmSymEH42tW7XoySLtkjR3tv
3rh7L9TLpZ7ViLQBvB6UJMr/p526g9wJ2J6xJ+xdRvnkKPRLSLNHqLkCXpO6iX0H
Xcd+PwS8M0UD1mlRz4ef3rbystnC+8UM9TUvt8h+m0slVIOHF6efEcBaddvxZ04M
+xSRUWgZTj4kSolBjiou6+GiHRcjEUpuFA4y77h6A4VKCn7pWRuMG4lEBL3cS0Yj
FMkPhEqRjhuq8usI8fJ+I9a6lnQYdlMg4fdAXpR9gJl49Y7pWQgzdUWO6E+ZEwcH
z6kooB4iIf9AimDSS9IOYdW+MgjWkSJ/p//AZWIVQ0zLJcXMH9tpcXz1dESe4dAq
ym2ZPKDIVzI6rT2EkvF4XK7Vm0uw0rlCFIqAxqgI5qa3vv/BD1hFs195rgLq0efz
z44vyzeAODT3sz3QuligsVyhoTrNqKtlvRjw5XgDLjYB8rRSNsECGWjfr4XTvdUv
cdO09D0htRR1EsiUQhY1FFsP3LmEtGjUKkMkYy/EvX6Ov2J+YR5xnCQK1tvAUWaN
TKT/CjQglX1jMj8Ucp/RS6LGtUKnwBDfqKBqpLwYk0LHjlkp135NAm6u36UwOrIP
jguvMH9JXY5S5x3+MmoL2OsiacMEghwmkUIiXT5SOvvO3lbVhD/BQOVUS+2CJVJa
Z4NGk8+orBMSbDcv3+ZUWQNXrIj+wPM3kLmGj1tvieEqkSmA1X1xOEnCnY9JNC4I
t6IDRpLosLDo/5Q0UpzdUJn6A3SgyiuV5Rcq4OO7yKmWvhB0mT706EYldTSGk8DQ
XJT3zpY58gubXyX2hlt1wNPQf9r2/hA/BVrVgNp9hNaTmOAv9ieFI8Lp0tR/O0pn
Sjy2ie0bUn3FDOymITo7UBcTS+oidWO9gxLc3nZqWXrxObtUK6J+z+HSypwAPYMu
RdhCyBJE/G3UyCalIA5MbYhpg51+Qwd31iteeNVaSTpFL/BNmbprriQI5NjCEAw8
3qc2FUfj+nly3goV0K0FHqb2/jffd0M4jriYrza+MHONeBkwqZJHAsumK4VgBRCL
tgbZjQkSd1CHvv1LX2sZyijlzBSHjrGoy31dr6kUwaaEwiBzQmo+pvCTUMycIDPw
orUZPOTtw9pxFrZdnmiv8QA1c1F5ona1YgrJW8mdmEd7d+EgUd9rlceBhBvr4C1Q
LFCWFhW40tOCjRgtBRAiWue/KY0bbxQH+u+Mkg0hxMVDPR4XLSK5mlMgySod8gna
cUmCv2Bh7STwdHcS6YqRb1XoNH7IZqm3LtW9cTRNQoUQ9JL5QQzxH5ZvXcTNb8Mv
MwVtRnQ2EZ+LLurBHR80xnOAb94LyIui34caOOZRP2r0kYKuYw8UtA//qQTY7gMW
IUTcqE83aVKbU82/RREBNDJpAKAUB5gnmamllJX34AkDWUQqrFM8QpajLZRbTWzT
aYxNWDQkFAUaHyKCiZFmhjqHjkwckkBEliUOja3RU6kXET7AxpOIyvJx8/DpxXzd
qFuA7sfTDjNm9QmWugiyCNI82j0zmttwZo9gIxgIXpTE7C88TGX+C3nvDrpzI/nt
GwymtnoRLkIArldjqDr8uZkJ+XjJ/xzCsoCo6XfWDQw6O3JYNaoupatwk/l60uJz
g2CRyI803bASItkoEGTEH53fOidy963Zy6+on0cM9N2nFcQsShiKIwbwy3CBfLw/
HbomuR7F2LzhNrsCrtdk1gPPheugJY8MFoA22IS8c6O4O+YU21PMwJYgmnFlXPNK
SenU5BQntcj/uHjK2L4Xm5bi0dgRevRB7HQZzF5HursMRF3jz2BfrU7HcqTCjnyE
lyIcss9vayMOFn+OsQE7zHcp53iHjiQGMMS9cUAKwONX9IV/fJzNUVDDL8IFkIEh
6jAxAmvOJ6DHZRYP4YkYP6tQnWFecpNGy2GAljMcfrsdwUr1rYdPgjCkgnilfJXc
tEmcwQuKDoUP934zV6nECSYgaOKp//YSh0ZuaTRiwmaoVc6tNIWgbJTvZe/49BcY
Ub9n3BxdRyjcY/Qgwsc7OiffOmbQQ9X96Yjv78AKnFSbMvO2/+mrcdEyQs5+2Pnn
2Mb36E1G8EzBsdR5xcyatWsuStn3cBPdS4BDtFGOe1W+EQkJGz8H7pI8uLKppEBn
rcjrZeLNsICMl/V/Tra8Y07MrAiXdiMzIStDm9nbbQDxwK9PB7arED/yPkmroD5m
FbffgKABFLwIhdSCqOHFtzOr8T6dNmU7rVZ8jH2JPGBAyBGIOguqjjOib7tRIWMC
1Gwg1Yn5ItTmp0W396VAppqO4xdTaKFX9gf6AGzQfGPr8hsj5TmeVh4XmNKOkXbz
m1g9rCB/wAGNWjfVd2Nni6ViBOwvC4m5p1FL2IOIVpUcOrbEpzIEAkG0GbqTBChN
YFn2r0KabCMqlREzGrY8C9vi0Ci3xiRCmzRPHy6i6PcII0DpFmRikvEZvtlaunYo
FaBGaiLtOMJLeGen/ydxo4l/eo3m+tlzYiomoMJBYPO/B/l6HcvSEhZyRBTfLFVN
6uP5q5kjSmLsTdfuxYa43X9fBk/YwTEqqk7y6oh99mOzj84N9+wY2Ht6b2n6eAZM
rzS9UbR9o2RGJO7ubpBLTtuG0EPqvyyf7A1aPfVNn757XZJd1w1cbhnlnqDbos5Z
wBGTYa6Djbcpe8zQQkNIe5XKLZKxnQKr7YcNflOxgaPwmFEJT7/Ivx9+n9M6fr1m
lNlbuWfzpAz31i1fuur64RdU557wg3tpsfeAXvYpZAOZ8gg4eSXR0YDQg22e8VTo
n2XrmYgmiGzhTHDAPgJIyAtosWslRzMMHCbkiFqtM0iZjjuWAJJqScecDevTz4ie
6B04blZ/M6SODwikFAxBbsRQV9Xtjg+z1Wkp3APp/J90oIYUBdw4kPhB4aEbnEJM
szbbtfwL5n7O6mcK9FaBdjALbtk0Tx30MAsHXaSLF9xr0PBEP9AJTeJzc+4GCicz
tB5aNjrdVT9MNotGo4KKtS+T7EmYgUQnUpDxp5HYFdOgbOKPmyKL2g6BTIGiE8vG
iVl4r0tjGWElxAwgngVoNLlkIaX4cP2QElkx2VGve9NWBYg+c2oxhwsSY866P9nP
b4mn4aW8UvRYp6IyHXVAsEAFXB4jZCNAy8fB3iKVjUw4Doj5lZ/u3icokf2anwf0
IXFFTEUs/zdA6PB2uPmquNh24FP8GOVyKQsAZ+mNRA4ZsvbdonzG7XLD79zACo9O
enwYtvYjybn+jV827LWSO1QoQSuUTSwRUQTWGWDSSGjdC8k6RGnBwPsv2mrgH+MJ
hJEI7KLXhaPnw9YdebKnJBeHppXRIKlVV3oE7UKIZVEKsz/Q9Ql70fY6UNYhfGSs
HKfs2kenQPo1r4n46wTPOlEbOhU3BiX+942jEr+GqRd0YiN5qp1apjnbKRcMSotM
3qPDcSLEAepF1y17grRI2dWoYIPF84mAuJKOdvOOoYeMJqIsh2yNnS4ryR1s3TUC
3cHEseA7Ix1R1sHmTR+TcqfunX0AzquqB/0fHzfGVfgAHKdQM8ZRkTc0hqb7AEFq
fWDOCR1FE8Dhg3/W9ZgQC1agfeOOSpo9jxBjuo6QJE5JzKPV4iELBaNzVkPf6Iki
PHtCjQWyZe+SFAbo+hpyFK+4PZRTzSUp2B5IJE7Wd8LrkeTNY2yFfupmcEOVupN8
1JwA3Ckk5MU41ZtX+eBY1t+sD4qgkUp52CEUHg4RRfoKuHp8RvRQYHU+5oG8mBZm
xvKJWcjpRGA1hJLf60/OK/mA5FNsJ04tRxPAWnwcFbhcLOE6SijMBg46q7ZwSJfs
ZnWNcDk/M47H7QSJWswe1H6zgRVQ+jv9DwKcUld8zQHrfZ2d3xEzU3uQW7vQ4LiT
T/LqEfixomi4djlA8ox4hpDdbBKpTX//AL/KPJ3zVu7EvLAyR2tDNO6l4+5skJnq
fkMJ+Xq3FK93AiuxZDG4NuKkHOtRxy9irccCctERDdrgH7rlBcg1PO5tS8paaZIo
yMoBZK79CV21FQbjiLtOpdhYzi5bOXgrFksilTalv5WaIEnBlAPixmX8MnpQEKaR
JyIqPUoj08cWIJr3l6fp2HOgLedxUppBWJKIYtn0fudRDuippH1Xx4+6kvJsoRNV
HHJuy5Vj5VvFZ9Ln65IyH/ymFlfTqBGawP3DLHtvMgYxaB/j0roEljFs2vBTokRY
aHWjWkdFnFv8XkhbBnxUWq0iIAJKDOyKFtjsLGjdlfqg6Jz0Z0MhrL0dlXbaIDdv
a5esv/l/jKm05QfanaFEr1b/ejBLEoVrgmLvKuCZuCZGa8GKo1tSfXdEhLMaUhyb
JjsumxirCAgezXF86YY3NsdeAHm7R5/+j+hrXAKhYpQDvszATHaIg9585Gpcyx+q
8GoYSwupqNy52P9E/6kDv2bO93z4QUaAydn6yviggJJmMJ7beQdbIBcR6c9a4ww8
JhVIKt+IlA4gUpK7uK9T84VXeAR4tyaGRzlw6+TRhmBmxraSq0wuo8qVvAvTA1OX
1rvZ6C5oJleIIst1BKoFP0oPzLiP/rsY2oHmI+tXwlvCYmPWh6D0vNQgXG4K6f74
zf9ndgYdxj+9isjy4ynz1mkTDN456AfYrPRN05TnchGx66gRnSjxb5qYZQR8MaqX
u8Tt7C4qowx5qz8aaSLHChg2L5lp/ATpY6sCnyta6VlRVO/qD/DPQXNpqPjfzLml
DtZ+zh+6e1DdMq8I/lPt+cL3WDwVl3DTc6D12/QhTb311Pz9aSLi3r0RIuh7R8oj
RppBy9rgGRUPAmareJZp8TPOYZWfKLOuR1Z3qLzRlf2NZkPzjenOa4paPYwFGBCV
uagad7xz7xgOqdn7x8vUobgBGSuNT9Zx4CjkS/ofCGy30VlS0pJVrQLXPOYi4tjR
QqPKDZQwigAjE8x+ub053iHLrY9aEeCImPcnczM+cmzFPyAHB1D90s9MlU7p6xd/
7P7EBhokzdqEklLpojxbmjWJJrCoYnEWBC8JrPpaZdmGTwmbe+y8GROa49LXhDAG
Yfenv0CuBhDcYahCuYr7iDdExxP4pqinmOE9lw8gQx5TLIcNPe4VaEnvZvDITbTp
Iur2xF2Vd5KDkybvDp1WYTc4q49Rd5HOFUDmWvzHodVkQo2gMA0+JTnLki9Op2d2
R/hrJg5mtam45JMnn7ETYhtkV2SYRWhKn7jtT0Vq7ztGIDXWKSXoHaHBzZhvm07m
NMyLvZm6EaXWvsTA69wF2WmhswYyQOOe1p6Enx15i9ryQAITOBGEwvEBpHI4HRA4
4puFP2X02vnydhsDR8uHMIka4E8yW0UpASUlgi2T2urtQWU213wOdK+Z5W0pOgR5
RuAtf4ZsPmV7vhzfELmye5QTr3ovRK6LNgn2oIyU59GjMiV17827o0MZv9lTydOr
wYl5YQkH4wTtweupSQrJjsTTs5xDsSEvu8NLv1wUK6IYGrfOvKb0i6C6hSMX0P9h
aK1S8F0bbWOgjxAi9IljOaHbwfmG1E/kyr33xeGqsyKS1pAxcwbDpL/qaOqoc6+z
dVspd5sN+OiCaRArZu7rDN5wSRoh5vlyQLEf8tvFyrMr2lHspwEHTNZDljZKdsDI
yAExRxPAKprh1x4pEAZQwxjAz0HmIR87xMtEc+I0+ZK1HTP0nQRM4bIgbqN/csrq
/MkkFiEkePyGFvtotD39+IMmRxvWot813EACsxVlf2wkMhdtsGHn9mL6R6P1KlVO
S89WwgB2opRiltxC6c2/pTMfr4CxUiPJnGvPGBDe/3Qj2yamJ5aK2poO+h5eEx9/
xhc4B4yJ/PNs5ASx/TanqQjNVa7Y4LMflLG+SncYNYhyT2exnT8dwRnKaL5AX7bw
KDRQ96rN1iS1jpRTUmj7k6adyl+zmW5hYYTO0jlqGH2fa2Xqd3MZgqenjjSNcnof
L+Gqq1eiolHm9Pk9aLKxWubG4AaKBP008o+1hS44tKMuxIgsZ/OUz/N+7cD5ucJ3
hPx1036zlIXxPH8ibxzMpwKyzG5B/EqsBcfnMISvs/NnRL9mmip46/KnXaS8xCnM
W/69n2tarzAR/ANeN5rJDHoZFBuKlSx+CCiFsyAL1kfZPQJh+htrEpPu/cphGtHz
UyxLNW4TXifbtFewkuHWbrM7LvYx87Vmp0GjlqbDU26BYMP+U/vXHxJiBcFKIH3c
xWJenKh7F4vLf2QksMVPSq99inQ/KcZiFuc4wXERUO5vlcto9rSCLrzWsOXVcB/4
axNi+tgiQ12bReh4XRdjP1jG4qUoLiWjq+kqIIrLU6vlwO9vZtQdZA2QNw4pj+m7
/1PAsarf80iC89VLIjKnTDujY/VXLDTWgutzXNsXre+tDU9QFiKtPJSMJ+EMQyWw
93ZFjI8WlWoaSy4qC2ghaJZdH4BSfgqPEq80h8Ik5szX9/gGroA3xUR4Wcpk3PKp
60g8e66wk7Kr/6g3fzc7Wgsckl7kMNX0s3m0KVyQrvT0sWAKoeloUdtwF652qZUH
t4GcWDfFGrS6ffFN37xxaSRbmbIne1ZT1TOwdpnL9FwUPcdLB6GCrRtS/PqYpL6i
xdHuOvYdRczxbzQEZOLv0OfiMyR5bI7DP9CSl6yP0v0peOrjizdKZyFQc3QkZQO8
c1Utco7DJ+XN2d+25GrCRdtREFE15PFpjiIc55+u/2ej+k5aQEKUrtwiEPJ1L2WL
xHN/u5YOMwx6luN4Zg9Fw0Tw+ssqLaTCvjQPKDN0g1Lg6UK7F9F8V24B+yn+UtTj
ih5KK3P9pMcKgNkBfR3o2bbIRP9foARuTF2GAbssdzgOjo49ONN0/DaTnDVsqNsG
E2Gvl67DdwsI2HL1K2r3JdSssYQFc710Dqb0mNL2gcZwz5aQ8P+jFUsdfK2RfHNK
UR8XuPGLWE2+3ygrBAGg161qTs4Dyj+ZVRPopAGGSiQMvs/XFV7GaY39xx1+d3wD
9gVkpb7ziwUxoLro6A2cLhNut+80QgHhCQ0kpQGaOc+z+3uIYwz/IRFfwftYdnsz
/cBUKqA+5LSvh1va1/FL02ARgUBFXp6ZkMKBDuzf1tONzZjoDjrtxwzO5RQcbNsn
FwBYBpYnIpO4AJbI/wo42dyIrjyLTzYsRf8ne0GYyTXn3j49Im2xVcoCRpx9YlTl
HpP5ay5eEbPTKAEb/qtpdP83bk/rfLos4UhUgXKbc9Kov1kNciJIMDf2tS4MOb4J
NcLKZxB0IZYUxWSBaMTY7JX01CFUgC+b2XYYRBUynSCEhNpQs3Rlp0NeJIuKs/op
yo1wVFZsrjCdwvjet8g2Bvufp1nnmTLsz+15IDVBY9/+qoMszNNy35BFriUj9f/x
bkZfZInAZRtUl2LWYtD1Dl0w5QOpE4t1T0dg0BXMt6uhUysV++gpKO19IpNZREW6
GpRAG2jAy2XKRDFm+XSiXa2O5rQMxTEgCuwPDxvJ7tcXmg+lPcoP4V7eSYHBxR/4
fJVbmh5bPQKuCprvvC49xXbZOArKatoqKOsM0025Dn5ZIyErQuZb3tX+HGySoZI2
lkIpt1d5JFiNBUrJ2Z8WTwT09Yc+87IKJziY+BXTZX09wVypjZV99pwLR3k15jqE
y63qB5Ie5Ja8wz5jeHRElr+pg7Sn49jS3WPzWTI/D3cRtx6FqH0qFX19J38VZwHo
YP8MEZmNYFwSy7OioCUv1ApHZ28weEc48j0nGrLUVTORidii/n9ZiyWr+fLpXkvR
SJIaDJKOmzWj/wxYnZvw2q7ibIMrd8aBFY5N1AYzpmHBdDAPKL46lq+ZMBH/6DY0
UEPAJ7jAmaoIm/ksVjlvTJ0r2Oerf+0Fxp7A4RS6NnKE3HxRONhLWDeYvzBCqUzz
nAIcZdMnjvyo7sA08+LuJjN9cCD5W0KOMrEIciyBo0rVUiiCwt/MIYvw5izsnTkC
QMrmkt20zGDENVH0pKV1bCQawTAhHU1O1o0aKEcT5cENEIZgpq3UTssUSM+mCjET
citVzSfRj1uJHB1e/9AULiV0BYuBDrLUvE1NDWfKqFvBspQAfbN18ZGhcRBX1/Wr
KuhofoN5WcqcHkBd6olis2v6GUE26glOdwazKROj0wuWtenj0yb1M9FxvqhpV6qj
LgJp8hUWKC5kpFfHdTwyUfdqvouoWagwRNR50u8GXY9Fq2Vmqrb7rx6y3GZgK1hJ
AXQbEgFoE2QNdGHDRir2khG491sqn4BFl0xyZd5BV/KovLd/v2gFui04JbfPAKu6
d3o+1c+1Te4R/EXfH+YYj3kZOUxH3h4wtXuduLG8HAP0POvP7ogEN1gkxiXtHBT4
RTY7uqlbvv8OGjP7cvQdyO34tdmc9PkwRcfa5hGS6MG3Ds3pl+aVU+Q6v5Z5YklR
uY6A8OyaT0d8bcfmxPEby4kqTUQz96GQnzNcs2m8HrY6ChTXh0GxLItVNtLIt/G6
9qzuLYuPmEErbnTl59rnwdYJ/Efokvw5vYBrs4FNa2eUvLqbk94AAjxZGt8Stp1x
bPGDneOZ4Ru6rU2KKTeRYlyrxuC2aPhWIv1h8ukOY1ylyBht6ly9pRBlfrSwkYbi
jqjQCwL3bLdicNvVrvdqEG78P0BMRj7+CC1vmKAuunyaEVexIZahT3H0/Lf846rI
Qz/wVZ6LAUH7hSKgwaC9N2BN/tdC4MD7q0Qozwx+yL66LyClmKYApxukHQDkkEgN
A42KwNZj60EcX40pKdZOH6dv+1A8EQchIRFyvuhFYxUWvmsq0RpFfGp2xXCxpWsP
EEc9Kbh1SMLyneqIrMalR9c4yUW9ayMB3XMxCCLmWT7xuWsti65ZaonOuN8nzadw
Cs8dRqhmM7Zo+vzTIOQpHDOc1nHrHxOwaySeXS1b6+6xT6bzLHB4H8YBpWBPEbOh
TnhsxKo1q92R45CiLrTWFI9KoG/DDLrm3Q9wHKp7SH9HHck5/qzzNcNTOry9BmxF
0BO0SBRi6R6xiyEkm7El7OlCCubV5j+5DJa6LvqTeYqRtsI121yRBE8YykG8BC+f
zWszddfKqmVNYuv2VLeDPg5IZkR0r1QujQbXDiec/IhjgKHfl34AnQOdSC0vnlWu
qxjRPTS1ogo3G5oBfiV1AAnGgYz7Sq3i3rbMt6BBtl51znihxcTiHyXIsz//8x7w
jbEeg8KOBUc7MvPtiCPOZiatR+57qY36ktVdxWmt2zIJNfZ6uatRcLpG3uLU6e/e
R45qAChgdAnsP2lms9KaK8SfSSV/CCovUVqssSK15mmlCfGhPTVT0TyR9PN3R9kJ
144YgSD3mPt653LZNRmli2WiTs1r0q12CR4WrkceRS0UjhQHbVqs/62obzEvwht5
ZsiJ4RmHt77mO22FtnkPCCk6yEZvQOAImxbNKUF7QKLyPscE+tKWKVguBasqoTRE
KLMGduwBZWNx5f59ryNvXZaVQ+lK2PEm993u0BalLsgRfYox4+EpFIGMg4N6tVBD
sxgbrHc/Elgwxtxy8AgjWXNirVlAq+OpSaH6AorfyWGPX1XkpUpnrhxTqLLDgmn0
Tu76xcOF5ChfBAF6DSBDsuHTIqSAm42HtC9bdClBrUZLAfvJ8WHDrPwhljZkXLqh
0XHJZ8fVswMHNlum2NISPNuEQa/OaVX+coQWnddox3ojygVX2uFd6EPzFKB9UZZM
1TVBw53QA7Ky4Qx8NqMga60+HovSAB8lXEjULKMuOYyAigAb+fy9kruy+XRnCVgV
oEoLUXEa7QQQTB+XhulAyuVOTrjmtu5oAP9aixzXnO3rVTxbax7Im1QaVUi10ALI
dlTVnHScXrJCi+Hp/Q2O0U1OfoHj7fnjifNewM0LC45pjjpgdhn1bIFeKr4dx04Z
4VEswao/U21fUdg9pOm4Ex3rZQ1FASlNeK7mcD6kiBcFd50P6OI3dQs+stEV3Fh0
k4QaofJ6dblE0YYuyh+I06y3HMUk7kYIJODb7VdVgAaeLiXdCYjsAObb8wYUjimA
6hfoC3LTHINxxw0DGBr/Ruza0FTW1uzYWoZGw3mrilw4TBZfpf96vOAJ1Xq4gWzW
oNhJOgtlvznu6o4DQt3PcBhmgCyT0VHlWltR2/LCy2Ofs2zyQgVuqqoLMW0EdVTp
8PQumWN6Tz8dfsxJa8BcNXz9ZFcGJRiTvNk73RKSR6unfS5Jji+yNkpvHqc1bpAn
VCvURVd2ey9Hxu7rzXv8Nb28WpZ5uVzUaUAyvbOZU+BfBa2UJi0nFVb5tFcTSMyi
gH94W3yzYOq4rz1Hm+NyOptAmnPhqHSio8t/V/jpcf9Q7JsiPNcjo7IpAYDsnQ7m
fHG7MaYL67TZg3W65tVynzzRVLIGEv+U6M0k4F3X54ZFj6NfmdNL+ZWnTK7ZG7bq
XUpg1uJDQ4jf7qC0wVdSrU88Olw7jv+LGQs8PBMYNOZ4NZx5C/UY1PE8Md/+AckP
1PkSy7RGE/SJUEKJoSiA7F1ynQoU6mFfTw2MEHqd4krOUhlNtojMcXSKwGYwQHY9
mWXJKiYgdiHa9dZW0wrpoq9pSKn1MvmjmqFyNE4TGjZPiZurtePQWtKKnJ5RKMos
pvYyQEXYsfm7oMY3KCikzDg+WcyFvsy2hqLFmUUkEwMCBmuJMXqrm2F3oXvzsFRC
YVhZazo5u/AHCTA+DIVd0lVa2I0kFCAQaozzk0cNy+bOeUMe7CQxk1+AETHXDBhH
ueehpqQA7z3avPuQqfaGwQ9EnDA2zUhVmfhu7hZ/WUdNQxANqUEqrk9yo3L8XTLh
F1I3/9/T1pgfvqGP3Mvkgykch1ZjlSytVGD50lDXG96xwOQm+NR9Fr3zRN3i8Bns
rCHCT0T/m83F1sIQsIWtJrzxnbzywCo0QH5Mtpcs6TLV/LaqmAnzuUeyJz/kZOzd
JnrwI6M53RloTcAcad45U/LukhNMZQo3ijjdKOeTH796j5AhFFaVSBFxR9aB/m6T
HcO6j2CJtSCY0CItFli4Kt2WYa4oNDAWKfJSqsnD1ktz+dNYLJogObWdrNyYwXNZ
JINBulxAf8Tpg++IDjpGwkYB3JK+iQ0dqzVFOViklV4WdEAuQhNFfebrMLFY4e7g
xIK6eu7U1SriGj4HUwhv5+9X9K91/2hpMUbhQutUPS9Gg+Ts1V+L4dC2tlvRTNb4
JSCHVsjRrp6fBYS+j+HsLjAtfTqJTltPqm0oibSYomVamcA25XVNb3AA5L1Jd67X
C3yK3K0Hp73OQuFWcq3DQhG1MM+8INx9jJFYObb2IfGqe50JGS7N3huERglS+3Zb
6ZjKFud5VQubun90ThF5O+yMDeQIi8eSeue/xWJpCXsUCR+4jRcB2IAHqjSrObxT
cjygShc++g8/RKHJUDKPKHKp5+qg/+cxDL+KWamf0Y2FRhKbGD90Ts/NG+mLZnf3
f+0TmjuaVf+vn0G/26SC+K/+qINM2VFVAbHzfV/PgGr9R9Ltm94Js0iVn9m3wvkE
jk6oqo/9Om1DwInxOuNyonb3sxjomrnlfRpEAVUaqdBoGRkw7c7cAJr4bFZk1zoT
kKwYdnd+PLW6GfIrYqttnMQ1yPc7Zm1D5XgWwAKv5/G3ATmDgKKihNu4ljpeBxGF
nObDshzqRfZfwedWRSzAcdzfy4ltGQnehukcyN15nTePmrgOEMu/2SIitfyKrVhc
ISmbPqaMPSsJFKTeZ6z0TaJ2dia1SyOg6AFkSZiF8MimaSRRyaUxVutNPT7e1pVy
WAaXMv0tdNLB/KOLcNoji7Yue6/l0KsklBNPp/WUNyZYD3dlwqI681y1kt38/oQo
v+s7nckcGE/xsAuuVv4ZXUdYNEKKIG2UOD0iIu05zrGmuG6ytMdDrmeZEpGuAVLk
9+bFIN5yXkwKBtsgOLXRRAfMlDoryvUJZwZOSEvd1Qm9DSiOTk9a7aIaO0G2lDdM
0cmaHhe/ftIdrQIsq100l9uzZ3Gm6KQxiAFNAoURSpAg4cL7r8RTZRslnDdErmVs
de5AxztENOT43TG7v2DlkjmlJzQZtQvbqRh/hAKIvgFBK6mxq64yh1YwVCdeCTqV
ikk9zcgUfQCE78MFh83XxCGIgrBILf9RPuuxHbQbSeQUSAG/iQYqKw0Q+pI//rXq
mICvn9xe2VwauTaSt6LURNMVK6ONiOklg/n+Ep18cfNklphntLB8DFyaJBzvG67r
xg7Tnfj8Drq9ROoAaCsyJxu0NuLgsJ/K92GE6GKa9DTgIPWXGDFNVLJCXGqq/MD4
qLurm28V4RMUiVq3JubJUU8vau9LiAJKiihIBNvYHPu8cYQBKnS11CKvhN/eZUmC
X9YhflZWOBjzqL+4CiRBkhlIEthwCCztUvMBWkDMnP6ia6+FhbQvPYEd1lFIUanb
E0KfqLClcA5W2Yq+ByYb+jUGmEbQ0bmmITi4htEt3rkYCeGtSy94eU0XJooEX+yT
c1TsiZx2/EpFscUojMEmKxP4Hs13WDTQBxMiKlsY1tYm4rM8Osp6m2rK2ya/dADe
TxF2RVpP2ZOghe7oUX73ned1Tri8Rz6RoQIF0nSjBL1CbwFpD5a+vC1kKcfRw1i4
NYdgoK0xrHh824XVFwIT++qVzjzm1ZH7zZP50uuVztFWGlJr6FlHJKmFIV9DxlQy
3YY72hVH2Z2LMMxMCPN1vRl8AqK5yvoVV+QcNy5Bfc0HzeZ+UqSKH0SIJTTUqmfj
gIyF1VYYXAkazVUzlIsfKAZ5RtiDsXJX5/lJ2qZViLMPujVHQmdBbJ1jrdAGGQpo
kumwBqZZlal9byto6mLUQf1IGP/tPtdnQN+mSWG2VbVXZuICjuzhzI+/wYBXnJ7N
OGUnIyErbM1zRYYYUrGnQI/HVD7VGKp10uxHZfJXfIuvvKogpBGb6sDtLSQIT7z5
wBNpCj76toE1mWiIJ3CSpSKFGZiuaZSGEx/5gowZcsfx57VJJAgNHWmlWoTs2F31
lqHDcHoB5bkxd/6UwWIfRlEZmSKowzjb3qRKaHlceHUBZ3DhghRdWartSpqwKHqe
Pf+OEFmX3exNfZGlHKVlCjKWCCrKtXoxET9/DeTbDTka236yZRFub/NJQRizhDu3
c7Zp9BRUsRqPeqWwqn2yUP6zCJzoCRPDoC2XhQZ30yqno1KBuGnbEzy2tTH26pDe
kIH/+H74ccztDdfA6qotZ4X0btm4hnOFgGW24eIzg+aSbhvRVNgJ+IokaBe4HDaF
P2/+euoO/KjVZP0dIrpLTLogBMJ9Iwg4qzNm86CTz5e8kfxo+wAZP51ptOkxYFcC
MdFr3Y6oyIrcj1M4LqCtiFuLDnK+tqtdmUNh3NegJbICvcsKs6tCOAc4rWlnWDMO
tJib4SK+eCB28GdTV9HqSAKoXFQENA83ucJULZCIRMCJCkQlbcnLvwJIwFyzjrQT
SCapETFH2SrBA6kQIOHHfCD7Pj4FNM3MlnKYboQAy+Bza+DibgJV0LomUYg37fo/
LziN7AwGNATn7CX9aJdcG7qzCz5RZqs1h6GqWqabpSJubgM03CGrRQ9SCQEszmN+
RTR+EWh7LZRkQv06abqo9tWiQhnZ8ngotSNYRPVs01cucSua050cb6lvM8KqSO7r
rTdbx9CTxlHwrowGv6E63tlaxUIcYtOohmBsvgk5MtBX+tRC6yLmIiCmWGJrcOeD
+dqSOe8RE+pMLUNzJhWzVohag88+NcAfCr9Zn76zhQgITS7V0mDfpm+DJ6SUlq3P
pJaU+JrQA9rI/R0vl9rf3CvtfMe+09oVUNJRB01SXsEDHP+zawIPUAtsybs7dZyW
4zk8TldFr8QxPDnfE0wVNQeyARviFBUECQ4RC9HmvcId9m5nOtjpJOWcLFdIKLi2
eEkj5/Sf6p8tFQ6mQHh8Q1A/hPL6OF4vTgNknQErhT3W7jHwNPEiLQ39JbKrPTSY
JMHySVtTW0+rNTDp2lS2fR6iGWzDD6mIYsE4gbuAeaBkp6EYkQgm7Doj5E8jXUBU
S1eV4AoD8z0EIY412uLo2ose6frINflI0vYbVgLdkk1poHJxtPtG3c51UMPNkzGJ
fqH4E3NV95xSOciBmBF10rkDWvTS8yv7/fpoFHSI1n1Q82qBvFLDmoAuFe2bWG79
GIlnJACZaPPGwoXM7TNyEKU8wLuTToBLa1poQIZCeyAbujqrTvGc5J3/iEFdWsjJ
vJ9Z1tDneSh4ta1SDeQN2Is4g2Tf7EXjxOwuC0EBiLu3zp0iLR6cJaE6K7QlXy0m
vANAvdLocDBY+5n8X5sV1TqhMiTwst8Bl8uYrv3c2cw++a81EC4bOf7EhTNA+s8O
XiEN2tRmLieClpqyP4yDIH55FFs5q1MGf1q27ZgUMyIrd3uyuKzAcyU4Tv0kmWiH
LJIADo9RBbT12cwKavLnyT5vMlToraL09BtQ2O/J31D8vNSakWDnmn8UKJd1BJwH
8OnzH1a2gH+HMeGm+Lk5iHWGZl07upHTGKF3DE3EvBIcpamnxJhlREU9HCCR4Z9t
3HXE/HNwzvo3zZWQQNy2xablOnkLdvatEr4UqCS0hm7MyrNQIiROWFPPi7v+keDE
TuuniGnGC3YnVnmWWhJgJAVxiTmEv1iPFf8ZBdb3ReeJ2QMQ3I7ZLp60ysdNoaOF
HJ3gxVpz4TW8XuwVOq4G/2ygPSdmZeqMUlXUU6Gi9VlDw+sP885R7/KUEkepdoLK
OlnXNMnhrh2znrofD1lvrtlrtp8XiGa2S3NQG0t36Vbi9ikSZ/rKojbrw+j5dH4s
/Ygxz7Ujke26S676c4dfVXS512Y8duSfldscySL2NBIgsBRvUMd0f2RAAsyvSGib
K9+SWplEI9uPvBfSO+6kkT43/xJNyX0ZZbGA2q/7UalREKvVGuezbn/4ScNRrPxp
o2LB8lLi/vQNinICRq0vtnnxETOd9gO7NdsdlHONraUg2rygtUQKgHgN+cvpUtZS
lTEVHXjqOoSimuG69mCwMgv+BpmHuDbtrtUH81gbNXKA+Ww6gfkcFPF+vXg7GUhP
q2l/LZzZBvpEQnihEWcwb3nXv2ZY+6g07emvtlT1Yn+JxgrxWf7khAKXwmgFgSdJ
5oqI9sa+k7g3+YOfyZLJZEVZHo4XIchuQeQHThnhExzXmUsw3zO23Z/2s/2Jr+nb
hLuGyxr8AjFV8c6uZ2LDLMqT8V2Ol5EgH0/uDvC3cjvC7ydUtSW63wHqIVJH2uaM
6uZqmbQbLHVSUwSSMxI+LZE7ItPifLrat+VuN0waxAXXTWFW4tGz9muMlrqpjPhp
ZvX5aOf6JLfhBN3tChFJkWHx7fQKQJCpXZa6GuvedFoTrC9J8ilDbbbFo41gqOH2
ye9CY1N4s0zksCJd3AphLRh9TWazF3aB1bGqWNYyCBLpdGawhKvV137Ts6giYT5L
ttA86QFE6jLs27btcKmCSGGTLzABm2mS/AxCum5oucEDrfMOin1qOBiPMQwB0FnO
5tgF9w5D66A+GxBebdJbw92Jl9ufxTXftVSizpRhptWUIPTNCSFJWgmr8vZuiqJp
WatIMkbAy53WHa3mICJotz74UyUrVxMSt+J0jJCS7oMPxiNEqcEw1DGvhtSSOrMO
8RuaU1lduOSm/LlyojL7Ik00oIgfRuge9qJR/mJof3grWTpJTxTnvk+bHBioZKq/
wIAPIh3cpiqrNScCC6Qsv1390giqOnMevtaXVS2bb1LlmfV58+a1fS6o8KyEdFSU
cqEVgu7Yh3z8VggeSGv1LNaZ/G9UpNmOdmlK0Y8ssxsV1I33EdOmXZP/sKmgzXTr
vOz7ds7287Z9h6ZC4D8A+48xs4DfqTjynOGpEvZbI5xTacNmiDYARIarILXQ9A/J
uHfNajDVDL2yCx9JbRZMJaKS2JvMkIya9t+c5s8+YmqWIha+sDQaPEjhDMasK2VS
2yYeGvrASP+CxoJz6qQlN4wKBY8AqEwr3gEbYOHbIOqIqm/TED8VeT+Qk87O7M4h
EOmA/wi2vyaybaPrZw/7jt8JLHO8pyU1vOZFuxbWQyonbqpTFdj5qeS87j+Z0+w4
NX/Tj8HtR3R7nE0XPABq9udxa9kBTNoJmfFoi/zLk6BPy3pKqe5gLYLl7vfAynKS
E6AjaWBIjnAer2S0HTIgMY4jf9lKqe3n8M6gBHo3ae9yJGGLxqES8r7EPU58XOJI
m3jH1zpWzq7U9PuYYDNEksvqywVQ8bzLl+1bmO8FGv3JTWc2xW9QEvo0OubcNTKd
MRgKxlfNE44XOhAU8tMw/aldMGkm9E+gXzcc/gorZV5YxRmjbqyeon2cySi82PK3
6qw6EehZBaOp6D/K3WsCn5zdQEWcbjGyH/JZniu1GeuSmalbEM7pOVeQXA+zlw6n
8IE45OrXH0fUaazTKQNzMDlIhl3FZ1j0pZas8Fz8nKR3XmDsl2Y7W2ju+izZmELm
6OnvB0YaUKTYzYbqN3IC2pqFeDUm8E/KcUmOGnNA5t5zwEnTSAv6x+17I0TGUYF0
0OSJO8wktm+ys9CP84VZASiZ8Hymfzvpo3mftpCO10jJRLjTs6XW+QIUGiWt4/11
Nr40hjzhXzToGT72DM6IlfPWCbdyEg4DSznFWzezAdXuevzLKatfxcoLhZiPeX7s
7DDTeMy9hrSvNZQO8sX60q2wmLBlUAGH5aUekv9ZDnYB7pkhJfv8ZmrOipobkAud
DRqYXHb3FdPuKh665DhOx4Cf4dQ1EJl18UNxpAg0mZjfdxOVkbw1k+Pkg7Q5hcGT
YFK41vHtUwzliVaNSCKtv8hNunIehlhpo29z0aUeLhGWhVtRsXlisbnp3w2JI0DV
euJ8RSlzP4OndAWlEo/yPlIU/yPxd7g/IsWXnLiY4ky4kTKC6BfPLW1BCtRKx52b
QLkECz6VFP2hvvmzZKpjC5rbS8nSWndTCkKFDUlxeVQtNmkBGCTfjV2aKQ/j5Cbi
KIz+zFMKfqiEquX0GwkWZk/ERjhP237/JSzWWtsVLJLsfkef7Y6ekugK4++v1JTm
lQTqXA8w4jrjvwCYDJmX2cVkdwZvXiIIoitduZdb0rQjaj4PjV0EuIR6FUtHR2Gv
94CjiNIdTUe8ZY+7zeQQqn+rt3xWHIN5IgaWEBZvr/mrQ8zTxzuGl+Yd5HVf3aFD
DS1+ZEVO3ghlT+V/O3s/I8E7F7wyLbNSJ8wb/OEEDPmGEF79vhocuIshPvWcIXrb
pOdqJhL1ocWxSdVKG0aSP7jFO/9ikASdxCM10eJ+zwC3LrVkw08vV4GOXrInuTJL
H3keL3cy6mfUJk0KT7pX+Ko0CGS2HONI9bw1ylnEjL/WtwsvU1B8KLjrFGgVm8WG
f7l6KwhWGnFZrO8ckIkt7asg7uUW5xRck3+Vz0pxToKl360VYQ3Cusd7PM19P6A2
uZsaYKbUvqrO4SGjdL56M3Nd2r7WnnlYWYPvmeAw2x7+21Ism62wewGOfR75Nxhn
QamVGcUx3hu3gxFIeIwzoW7eZVAdmx7T6k5GGl4NyzDdMiLq2jgYsc6+YkEW1b3R
RcbV441J4Ij+5ctMkcSiTOndPmx3jXcywkXM+6rbD1TRrb5o+9J/+atJShhJjjUf
MoMhIgRhW8T4jKujGvOXhWI9q2NhZT+J0/ddQ0K8Cm00zUj+KUB79LBmEWeVI6k/
GtLg5CCIrfA6nwP1q/SDSfY/FGr61cEIF69lw7LCWf9e+RSej+n9T6I9cvxjjjL+
pwZqf78XnLzS5aQSkWYWY1SbDsWnSTi/ELCUHfmRuqnvPrgX5bpLb6jsEPlca8ru
/D96h/2HJ3DnHbnZh68KjLvPdZbfHLzvg+ASw9RIKiXMjeCOeFxuy226EdYeAWYs
du5CgDT6iWnU8PRYvs3K/t1znFNpGkb5AxeGBm5OuThTRePyUcDhYZk6er9U3e+9
F0UexMQT6ECzWHThnfLmPNZdHZnKpUZpDS5hY9UjZMDIvwaFdMwfri9LEBQybXbE
d8p/+rdLNWHdYyVTbZIgNbFoWe/vDWeUAlIZ8V2w5Pj58Id3BMtSgdM2FwwYxk4S
piNEP/N3llqot/q0q7AdKDpTpFBsgTacu9V/9tPSsD66iB+cEZT1ZfzfNlKluyCz
MWNpHvR8u4jdRq1Ou+DbXsGfazIpNYJHOSUiPCXivMZvUltezcUMu5DpMA9Z00cr
4fIQchXtxo7FJSFZfdoCwvSxYsvhsJquFwO/CNp/YoYem8KBf9c74+COu7rHtZag
IkTs7U8CpIYl0Eu4ZlFmlDC2G1Dq/MG4huen7FiQrBVfKeMl04XtgA/3Cb7LPfIo
/TN4gtKbnxStXQziOcvaNDouT4qrShmydBfRVuThbfhFQ5/TuF7uDcu0GYYVMCMV
QuHWub0pF9BSv0WCNkIvsnwrH/8fmGpJvaMt8B24nh72ygOm5XlqDbfN6FJxi/3x
lXftlKhJAvxwTzY80je2aZ7In3m1hW6IPUdM1UcjWqfJP4OMX9MuQobTN8AZ3uk2
zTqmoWCovnw/k9AxtKPQUxA+1oj6U/Z+oAv/CzuqZ06fmlI4lROE7E6dMlLXwwWT
wZ2HSfX3c9RtuhFsavmHkaz1BHe1OUnOkNwfTKfdqDTB8RM+HAxA8phhD3AnkU1w
Nu/6BNTyFpPb0iR6ewvL0f+nRRVFZOJyUhkFCB9pgyIPDC1MVx6aURYiwGmBL56Q
tXiVxAYm7ylqisNJusHZp0gQz1Qo6QXfdfN7OvbhrEjjY/Bza+FiutD3DPsLtU8L
krG9qZXpih6cR4Ja2Y3RG7btg3b7e8w2qC4YtBWhKQAFO/bYy10UrK0QqScSL50Q
cUwqd3fcRaj8cnCcX1S4HJ1bjQxBB2kUSMJ4x0WEvyojWzfvU9T6g2M4VFWXRNla
4UVx5+1jjzz0Tf2iqjaQ+UuNwB3rJx5O3KKWi4s5/tg70gD5f7I4sD/teGeNxUQe
MTMv5eZQm8TziFRubgEuVzuGIrD3SEt55D1qa9ffohrSo9VHMLolHM6kZ06jPY0l
6pXeXd3u1Tuu9W0QjIMp3xTe2ojBzBPUtmu7/zkgImp9NODmUA7+uKYxHrc35xWr
RMb5Vxv0nwMZQ1Z5kdSPDF2FdwbJYl2f8IZzVIBcIDFNsAfR6XFstrxMdvi6+QnU
bJZLLKBrTGQmmM4J8eEv0dq8+IIkDj8Q2yRjiPiemzmFdDmrIonZr+W2Ho4q8Xlw
xeR9FLEk+Lx0EMGTOLxBydQjo7tA2fTDh62+1pTxBjFhcuImG1EBCLk50XWWI8kS
55MpXEoFHRMcaXIJKXRvHyD1aOl2VZPo8Keie2bOn1kIkYzsyU5DJTUX73hEk278
PAvzzNx5lssS83fd/HPh2xZ9Qw1yv0gKtKXnZln4vGySg4qqrWtqlBKkqqfPF/+f
4ObYhsCWDZYyv+beZceOV7hFI2Pnwix9oX8EuMr0Uod2bgr19xcTKhVjPPe1QnYV
EDB65JwR0yAWRA1SpaiyjUxf/CdxbBMna8B1qij9/NyOsTuCy6SBxc5ZAG56ytpy
gFE+S+4hTcOJVa/NhT78oeeiqDjWrbv4cSScJa1HGXP1MEA8Q/RL5GTFARH+Byio
zcXGMYQwQS+Yq5gNS4RvE79M6bWHWItirXRg4FIbeecxUDeFIXCcQ9Pfr8yaGRhA
rgf+d1U2mChBsL23WYFqbLR7i9RYrJo6Lx50FIB6dC9MGGs81jt79cHcaNph4+pF
WGHMQtnl3G5Z4FgR5n3cxAJe6pHMFyZXa3RHDr+tVxoKrLdHKW+J3Bg77YnWVK7G
NGX9uGmkIZPY7XNL5+hmVgELVRnCD3+4vZHoZc4F1h/T9O7YUghvoSdJY7bUNJyA
dS3X2tFQ4UsUrTP/Q5XiBcWZYpKOO5rzKxUwR/QYMZXgZje2rX7n7p0CjdAamrYm
94OgRfJH4Qxowi39JwpQ73pFphBqhabHMJSxHXVYs7L/QFM2CA1fPeoOAqOk1sxi
11fJYjJ9I7Fo+VhYd6U78Xt/nLj9DMv+qU+ZuUHX3xHyCQinKIhxB/bhdP5BT2Ja
kAtG8r8FqfdrGpYrnon0vtRIYDyB/htnMhukov1wmRGWAX/aejOwc4FiuMY9us68
UToN/VRNbJkJo61C/Yt/5podPtwJ4jZ8g+ogNPM18gA7HCapN7ld/g9WyqRs7Sbt
gQOaRvgPltxPZUdDvpzscwhGtqXgRh0LEsYFrhTAJR/OjqbZeuSR513LIh9VkCJk
DmRN8v6whsKLDx2cv0k/jEiq/I0BjtCY/omv4t+572CgKzk2twIZre2Qu3E9xovA
vYuW5GDJrVqP+rCUXu2VPj7O+tawRON+wVMiyT5T9D6ODFQZJu3MnH5M4fRpPqfg
5x0ub1DYF8Z/8zNVm259EVOVDYcchmY6GiXopiNrTMbZQulIDb0jI7hi2EFNDaUg
mhUiiUx/bKVulbLYPrwooJCK5psdP09sp5iL/inj7LO03w4+Br3fimy39QFydNpK
V5GDzyouDJxDU6u8w+QLc/RNdBweBH1XZNO7l7E9s5Sg0r5rn0fJUTzX9rWYMymy
CgSHSvimgvxKM2Naj7kJqSJV7Qujx1ldwpoJJmTeSffNHWtVmc+t5i0BDWJOlZja
Wbq3ikWykSZctvmbGdLyfuhff1wUGzliJ+kDYtzZvnEUXqh30UGGMrM4oBT6qUvP
8u98V6usVzzoF/fENI2ru58jbpmvdYVTNcfBpWT/A+WrmTYPKutnWb0st54B+K93
uJQhyrsUf2kZvWnN9wDkttC2iEC/GgKMk1nuo/gUDxRcknxjtIFconD6OavvOnTQ
sNT2xC44BbQB68B7zbmLAYw2CpgrMGD8pPpHJGrHJrTDHw8tQErhTRI3hN+UQChc
tL/l7kSxNjm+yn2j71c1Eskov6zz9xora3Zdmi4FM6wL9chV3Wos6wEdyDaQ12Yi
YjQErTWM0em4fw7GkH5e4AGzBJ5viOtu57SCno6Sl9i/uAeksEskG6MURHIcen3w
iCZXrA0o4b7X1jHlE60/1F7NOLpC6uXDomr401qZwgjMExWXye+dmXz/fQycm8eU
+6sft6l11X3ITvvPwyw9iAe2BimlA4+zEHm4v1FAsAZCI1T5Cw2JzZXa6K4x+uNT
ff4zeC2/8tpRgT81hO5rtbBQ+bQedP86VT6xdZv7w0SZIkyTCD7VmKGQJihlwKbR
C8PspcEXqgSaM9iBhY0LUfTb74WEYAUsUgdx78RQU8tMW7gP2R6LhdjAioe0Gni6
DM8A2uAdCI1Fx13Ew2QtmL4geHc+2RWAPvfZkl0renYDX1J4qOI/cKTDPKssYcfd
EtAAQUENVt2tvtu/rjndU9HSY8Ye+x2qj5x7q40zIPxEQKRYbDo1LvV8vkS0wV0T
jtp/tRxmTAsb8RwmgTFW87lLF7waVzqYlokAjw8Qb5obgL+QmV/tumDICoTzV3LL
3/CvUCagBodWqBv06dMN08nmdkpfStlHSmyIcc/uXujjK8VUrovCedrmb2jf0IRb
PKwQOogM92x8g0cPyLVdB/qli9Eb2YLuM0qOEBo1xkZ6XbOZMmYqlLuGguvit+HP
v2LCAW8DxuD2R8YXFil4nolHmuY14hdy4+G6pN3S5ExKh/JYWrYskSOJ/K7hbYbB
EftsOnqgrZFrJ7dr2vmuXcRevgmZk7n0zuSEo0ibh1lDEWC+pP78klzGINSliVzT
HzJ0UdhWTVK6t1HtkBr+ZpwFqOp/qk55iWSCahjmVzEh68atdIwKOjGkISgG0qCS
AKvgPgpooNyf3bcHHKuyu8jL4YQLnifV/5LV7zjZVnoi7PV/B5WVg1x7RK3jWX2J
dg/xO0lT/UQAhzmsU5AvilERgqQM+3RryS+ppF/YX7B6f/YD/RYLOTrRwDuWN1kr
vPo4zei9CzAtnA7ZreJ9c5qQJzvA+RYh6hpaYBjh5y5EVw8NL+T1Dky48b/yXJRB
Kt8hr9p2e4ZZp+Ci7TGnmOmqIYPnDnFGyHRNaVAmTxXCV6DUgHc+uk15qQTKnQPM
byqsqtFogLNxhhTSal6JrdkuMJMnqeA3pkrMdpytcaehxieftJjGrBKm3Pxw1rkA
cfwcOMP6ZH75PQVBscqLKfjinnBRTV8Coqff4UF3JMi4ruNJTd+IpLdMqPeZqiwS
VkvmZ9OtNBgshrvSniBh6SWhuNAjT6PmTHcfl5tBQcN6L/XP8NzQSLagOt7J2avh
Trd4bz9FBzQYoLUXyuuN9tMcQ1cHhwovlUlnPNvA9ylLBFXlvXFCbuC7V/8CBA8C
ELXO3lxWnZXrJ3CeRZ71PyD4w3C8Iu7/vO2Ai3bg+mOnTkCOsbVWqi/gFWlLch4F
rFIebZYqcu2nF+8SuMGD20yJ4DpEv/dw0YrBIVOTCPwekYrMt8OUS9OJ4r7WgcRn
9qTLCdTvyzZDyTEPUyEC+3mwU6rVqcXq6xGmRCkmhLBO7tXQioHczCLvxsR8/yxQ
YoYkxl3P2ZdaBz1ZRzxMyQP8fXOOhj0La9+90c9ujgouY23ma2xV5Hl6PdAwpVpC
eotMAg5pQTRk8Nf/IoBDAS+pJagWnBWAR1y2SlV52qk+g6Vak4TBKizd2JOFp7sP
mSHohgWlZxTKygGCv4mqLGY3tkCFFM87OJLksba9vdUFft2twQG+TBB0Igt56N1l
g4MYi/UjTjvt5bdXuedyM266IlGlPEsZuBeDFd8kFE6B2n3hVxssxwidjsbDcZ11
kGwt6IP3yBAaZ4fn77TU1pfyj+H6XWZA0c8evWyuPhqVCNVJ6HRB7znHZWM9oyu2
p0+JEMKzU+usBRVq0JgJjljlAl3JfY8GZnGxc0NsiK9CSy7IWnCVe+aDqC0T3uHP
a4kv03pgJ0EVpjbeBUulpAt+qsUJnGYoefhigmYjXS1oSEZE1Juc34fwpHL5W6wX
XfFEwVl4EGACBdFyjwfdjxkGSd07D/oWay7zNB1rJBJo0XlFRY4wSq7QfUl72/47
sTUgdDTvoMxv0oG4fzwFe/lihuqoXsUOBdaCoIXGW7oDudj40CxdLCZyAtJMlWhf
ViC7a6a5nkTRJCVB6o76Z9dCuaIr5jAHTnOwtK8KgNluruXsvsLWWVIVSw6WOq5d
BaP47mrB/rsMku5JQTMtUBFte2WrQzMk8vsmRS4HYZwppjDGTNfrWpZp4H5KEBm1
4HZZksIk2aqMMWZc/a97a8YO+omwHodJSfvG5VYNMqvnqig0y9yHltr7z4vXTMuM
VVy/Fn3ZuqBwv2TLL33K3lSrwEdO74C6Xiq0KIku9Fk3LKOHb/cyAeBPl6r/xC9P
rUo/T5tO8ZMc6u0yoWhg8MIaao6Hfddql1LOptvV3eBjcI5JiuqDbgFqDbVT9Hlm
igrb35jExKbsUceLZJSEv/yVx1OZmEyDg0FxiNGlCp7fnA+IMKjRLQjHRjgg3pfV
H1lewo3M3XfiKyrsTLjqWoT682wYbSpmVaMDz5EZ9fKafOhL+8X9zfdUsCzOA+HW
09DEMLRuuLJyN9t+WTG9ExOgvgpQUVIBoAFZISRO9KRI+zzWzlzu4BBpGs/C3kOG
YCYu4hYfcIKh9CrCNAjz2TVZoaF5ZpQ2kBTQuF5R9pBNIYcgijYaImUth9vbC1G0
oyk6RitCH84+ZQcCtOFW5rcNpVmHZLE87lHjJsnakyPQ5zunnlAWWG7CtXBFNN2h
9VgGW5MOM0PizhMRch9hPGPd/FAaJcUKuaw6BuRcde/jWp49jwWSedebBu88uE00
ilYQWrjjl26cXCAWgbA5dV3x3YIe7DonLzDeFpH2/Mfcv/X6+7UF4TsBALwsrYTw
TSoBS0XIXxdIk6R2BYTz6EkYzDQuQWcfzLKn9njoGyu7wMUwOWm4AwRTWNX0yyVX
wBH9sT803J65x55MUcGyoJCUo5kNa3GYjpP026qc5FqItY7RynpLSee1uakDmokj
BKfK1UF23BQ3nAYkGbSvmZiUVhwMfkd4Fpxjbc1/InBPYMGjPgEzuzE/P9WnSASF
Eaj4hWhR0/JDNoJUb/wtCc//Tx6XDY2cT4Fmv7efLooMo180XoUiBtzQ8iGGIj6P
rh4C4v06Qw9fA8kuoZGYOLzXsiYZ/aMfubT8RxltOFyMfMFSPoyfjJFivSDUsD8E
qXvFbhId8xY/DqszIl9jzvgIbN5EPYUdv+BYqV0G/zbNo1wMord72/CDo2+1Us1/
jk4SsT5a1VCOmjuWBzpzgRPnFIzgVV8GBmarJ441tgDEltJfljd8xqTqwAwE1E0f
4O1eENm3lMOzp7ziBpW1OSsG2nOGCJ/hngbUuIPRji82vR34Ej/JbXHo5+Q0/bdW
NR3J4ezfBT13qJZxZH45lMv3o1fEHNxhSozy3+09zMKo6rQLD7iyEDmeRa8kMPnx
Q0veuuZpOGkvvcjUv5kFFZu5iH+A3fHwvfcgfqjcZTwif31v+lY2Kki4eFcjBWB/
jHvTkS8kJ5k4NC/Y9Hq3O4DMrz6tGS7jzWt0nrPfXN/1pDrilZsLBOr4YB+ivtSz
tZVqiaQ9AERiLrt2wsOPiZIkhh4mY/+g7WZXsfi4RXWe4k/IRrssGCZrNYNN7n87
tkwtNWMOu38odN/C5y46TYf/mXCwU85Ug7OFj8kF5b+AuyHOftdNvf5MvutZ+KEi
uPRAAHW/eu6EnuUwoZ5ULlKWRB9/O5T1DoXpQ8ngW2rXCq70Nd1tagOpiBWf095D
8iawjx2ejFZnw2hZCEq4TxfgZRzK0ex11WR66KOdlCMPyKkLOOIoGCVowP2s7Cnf
hlXTi40HUSEe80FGEE5/VpWSBvcADh3qDxru11kKBPhSGVblVXjOEKNP1AW8jh8t
VdTtrvrcmbHU8nQfYQ6ov/Zl6b6qTNNK4hzMJN8VWlZwes+j2wK6YzcIZ2wSs9OC
U5i1MfZ0vE/xpJ01e9zSvj0pHO9Atz6VniZAuG208FPfedl1xkXuHO17w74/ZpKY
PV2LaGUmfiVrM9JTHtHNPDg94RT1yaY5jI4BVIC0VwdHV3a16KTwipTgw5cychUE
DfkiBajYfxEWqY5ObqQOh8tIu1Y9W+lgVv0ooDp3VLXM/s95iQbISkptUmDqFVnr
PstZcHQFSwcV+Tjb35YDg4Ja7SBTUd5v0NXDmaR5ghztzAZrCjmRWEW0D8ze+wdh
Y5wN2884sXCgxYzsGp+xAY7anE5j91Ip+iEgDw2YrImFdMBo+OyUQwLzdadUYld0
N2DY7JwOViHSYsRvrQI1+Bq9o9B6d8WHj7tRwagAITJL/7BOwr7LYUag+hBCoJUY
eqes4b5n03q2tZ94XjyRk3hm6KbNn+8GgucHNaspleoSe1tvpM6P1FzK0iLXmzT6
UqfkW+s//7MnUVcQVLB4w0fjbRjsJE21b7sQafocuLNyn9FqpsdbbIt0MHCS0nLW
Zca7fekaYKSUY4Z1ynL1UkAGWwVw2W62unoIaXrNFeJ+jKdHdHjXLdlGH1X7NXBH
bdm7WuzRgkMKNxgB3S9cseqHazfbsdovyda9l8t/7AzE4lUKeeG10ZSX8ITiAysP
HfBCA8mPA31dKqBbOlCS3fOUdRNnCSg6F2yPxA3k0AONiaf/+pFL1aRBmvMt+ZgX
4SCTytMORJF2+4GTS+YHDVmgyZFRDf77cYoYzT7XEza/UhNtcrrYzcqzs6Lzb/+V
MHSMEx17hHfpVHOSa64jkY2LjKA8mzbj7HJCV4qjN29AuJDR+MKO9V8rXu77imsV
4r0ZJLEQRNWS211QMJjdr1ivcIcZEMvx7qAhsjEE5gk/BeWwt6tt8iWxzOdWAPSP
prpL6XZLphjecd8VR+0Qj5OpCDF7wPAyiz8wMgdxzmZiE+HoxulEzpPQi4hFIX/C
dIfwAxdcuj+vRHJ2kRv36oKypcaCpC/ORwxZttATJqPnswzQ407sWLiL+LRGqSnH
0rtsgeWLGlmbWhcKN5zUYnPZGW/9JgJvBLPU8ddvxxRolpHEz87dBoVuOUH5TnN8
vn0EGEo/GmsKgKJOb9L4rsUmO1MERoXC5Kd6xmUzpr8MEXN6L3DskrM7pP/BgNpb
DXWQ5z/axM7W6bw1NBwVERGz5yze737z1tdzhuUntBoyDXtFpzCFJYXwazurX6B9
gPhAPNqgSGmkT0DuoRtmE0M2fRCbeTWoPL+ArpF/ta9Tto2mgwLDzz8HGVZlMfjs
wKroSs1eRHLLk5xCphWNT55NRA/LiHWym6nw+qsNsrE0gUVSieWmX+5WVpHtndiR
NDM/it6ReDKilIYvjR57f9ge6NtIQEj+LEkWd/NCxPIQ5uXvqL+zSPbIdlL0lrEL
sbWOyNMmi6FgAYLuD2tk3ipuhHKJEmuQZVNWz2j/j5nwev0mXYbadttgAGYasayk
9M31XOisSDJGpRAiNH3DHiRRmSI9ruYpHVvBVBZpLK0S6OppzOpfGCViyobOC55N
2l9SIx2wj4dJjiDYI8VnFkcd4ZbFrhYM4pmI7ikTsJLze0+HphJEhwJaSyuKoP7Z
YG7z+oFbw+VoWssyDwrKjtcgYtUkUNuA7F1rtXse84D8QJ2mmNyIXVeQfTqJxwRS
PqxeWjrHCW+b93EGLrXTlBJQ0P/OKpquXemSN79ahjqBAOCm4UDiCeW0QmXNyGWD
KX14lU7lGZ6FgTQFpNDzZ8UW/CXzk4vT0M323QCaSAGf5+YOpf81Vyc6T9ozDHxt
7cQPqp26+CBKCNTCoQwvfHul1xGZ/yc7fM5uU31Tr+1+M7dASsYfEF+chlCSSe/e
U62uqhnK2E801xsJj5SghuSKINL/NXwHuJ2zHRQg1YDEHqHphCqF+zUYdqOOFNK1
h6eNWyeCPFn19DkQV/unR7chMb7zwwWheiz8xlU7wrHig0kCu4Qi/AhwL0ZfWA3j
bRLtzOncahek3OfAQ9nk4cZK4ZWtPTlxrFZ6UdpnjQMRtrTmNzxMgaJNrFmgAS0y
REymV54QMGtWhVxJ3SVoI02pr9PsKHlKiy0Cx0h/1xsE1Yps6RkVshylFg6TndEB
z2N84eDvkQOGxYGALLKWlIjB7RF2oZKOjaKtnGBAQXdvdD6pZ7PbFpLgxUWXNUQl
E8w+7eY3IPL7cVFML5S8XxLkKThoGKFADScZ5Uxgf1gCkxKlPvXedJOzlYi5qNxn
S86VQzgbuoGTOrax8b1MqvhuVTPQfPMYsl0nfiKC3rCPnAoxnZtdh+Zme5U95XtO
OY8J3ofHI7lCuOdjpNxTI72r8pvO/KUdJwzZhZocQZPTEzpgWahO9rdsuFuqPK1T
75KgwpaIudJBFJEURHFJ2XKSjhgkKKnRwqlOihnGtksk6FJeNDA11psY9H+9x9xP
bEVG4WrgUwI9TnOyuLwY/ZdmbidV4eCyTf3w7jpAYsmLMcTOI/8DE6Y60IS6IYrq
vjFFoVeINyF99qryzUpuKCouTMcWLMnOrySIgPz7QpxJDURte5L/tyTfLL0sixd5
y2ZQ+5zVb3OWvmiiLZn1EK9U4mYY+4/VAbUo038gsSfnx4X7UOSWcWijI/yBy5Bl
wFDUzFHeexfbEI3BtHsdAkKn8yEsEzwxhukL/WT3j4UNpmiCZwJhQhHWL19h51sW
rhwDjj547vyjrSZGQoXRyimiovDSC9iBdBG0SPdbImnYsBDASnSgX8smFTVgzvxS
9y/Q5Hr8gDx9T51Ak0jz+bPJ5RCJt1kqEp6JGQclfa0ezy4Uc7Fp1OldDaEu5BXw
CpEV7XhSgto70JEVM6iwRU0nXk/k2QEW5pBJxC4wGPYpM6eohtKCJ5CnhsmxeMio
gWxIGIvibZTw/YNKWsRVKaBda4cIECl8pIx/SLWNLfTvbM/N8eaL5Z3e523mWPFr
hludXRlhZ6fAxwaaASo00YK76v+yP5WYZNLZD7jfIG/90Z9KcHVBzVJqNU0qPFNc
mObqtpjuBdkohiqnu/4w7dgQzO/PbNa5nULHlkmi5tNqRyp/vg01q+U1Nnwkr4Hu
h0Ga3AVueCCLiMRwVOHHEX9pbSFzlzgnRRwuAcPp3hm7YgUYvo1/y1t8fbTzwNRD
iMQvzOZsZz0lQbBgX3iGZBLSxD8lqQ6VNNWyq3gOEC1JhzqUlmdv28/vkAN/R/73
Ob2APiQKVY5hJBGzclDnLe1k2QO+Nkjd1BflNV0PitCYL1Nb8lTkAlGiGChDfcWe
Y3zomjF4/760EY1mzuvd8WsPo4f/3miBp3GPDJ4wzUrW5YD2sB6lN8RTHWEf3Toc
WOQLqZXK4lJ6DMWEV58UE1po1VfGtpvtxpCy0JxDXRUex0EAmrRIedDGCCtefKju
N6v7XDqbyt1j9tf8kpcRtV1fzcwEgWndOLS873EW0CBPuotGkDI35Kho+0CDzP6P
/Gjb9kq0VWhusLaVuNOYys3UHVgI+84EIPoIQaRn6bW2lms6GuFXw170I28yVQgk
ti1+IA4JswruIF2WDXXzYmvL1bAFsUetfZFB5EnOSGxuB9iBXl5hu3OaqTbKtm4p
by0qsS82WJeAiI8Hg//3DCFz1u9s1oCE1z2FT52Rx2F9FmcjdVMg6AtRxAHBK+7r
aA3sy6/Snp4AHeJWr90hsW+uPpftAiRV6ql/DOXtoH1w+ntfoB1yVMEHEJ5YdMiJ
m7LgcimDQ0WWtyiZj+seqQEw8tzxP+BhCRvMn0H8y/lkou5FVOg4IIfeVM1YQnCB
otbO6peNTByKTBKDOeEV6AyZLV8/jo+/6vZErnVuLa/v9OSkyOw4iL/njT9kq+cT
ZwHJxbUVg9Vo1TyT90JNADb4/qeFOonbUGS/c1GrHAniaqLF0f7KYIK73kUz+JgM
n2uVCSpFF6J3GLPnPXEfCcNtz6QhPr1fnr1eSGLs9JUKTdhewPchQriGq3m8wY9x
mtWKAJ4hVviW7jA8J2o2HuBCzods8fXgWQb22YfUHQSbDFROMysr+xiLzBj696f8
FWsn4dgHznx4afx/RzymntWW8vedcFurINtLUnh17UP5za4Z/bz+4KO+hvGMQEWH
9/9d8nIYa3INLnJ6lAN5vCPUDO09+NsVz0uD4BYGPi+hqyUE4lWShUXYVkIl5hng
HkYaI7EOVJ1GCYiG2FPKhtQ/BVNsVljjIurpfZJvvJH/DU2M1MK8+sO1b8l8e7Lw
xjBoeoIb/I4SP73kj3/9R6euDrh0v1G3AlVRLZMs6GcNFOFBstJ70qCE+HKgcrSd
WsWG9CHBV7x0AeAyjOfcP+7KYTz1KDuEsLE2e7xvgiG99aZOkJEBGCMHEpI9yYU4
XVsNyS7UdHyoQi/BokCL+qCrhYy05Wm1dPcY0GveManwgOQr/bSQUm17bTMivg4B
JMGfU++FRX0yADiblJPDQsgnIpI+e+KJA1SYnIZtiSaENFDupMksP2abodubnf9w
9AowYlZD7SYdUlCcnQGTryJ7mrMN9S0S2x6DFJ0QuQxPV6tO82eNFnYGilvGSFJB
X3/F2aScWDYSkVnJ621dT0xq/7TvtEi2xpiZaGxjI4PJQlHVYNeelieEhGnGl9O2
hyELipukb3Y5N2+n3WQxFjcHnEBZ9Z2IgzV4wXYEhiUnuZjJmNmoPu0RCUbMqTXw
cV+VnIWCaOhgh8/Ruj9Ca8ratgU98oRbABTd0Efjxk9LzOgz7jJefkP7bH4q4HkZ
XA4Gj3md2HovcPzFV77Pma1m2TC5b1PPsaN3Ld6MhNsf9o+O0aO6NqbSmIGa36+G
aGwhAP2zL4u1IMtHsXgPqnBCahccFFGfhUw6vAv5wDh8/kt6a6ujg3JUM8RrJXC9
N91m+A6ngj87bsXqlzH0TIrirNKQUnrPjOAdv8hFmS9pozoQR/QPi/jcVlFlrENc
iqJOsgNZORUeOgTXfLYQqhty/Ue5Hdz5M0YSv3iY/9/CkzWV+B3Mj4tUe5jJM8mI
gVBmZiGYMwerdp5D3/ZUdEeBMgsko2tWh8c8OfuFwGnHMRAEcVRsQ3WUOn6Jlc5G
gusOa7D5lg6sm71eCZ1uJIm0e1Fs6f8Qf8m5CnN2n9gXdN1+yV8qds62Hr2tXWO8
ZhqOP7gyPoxNaTuUFGcp9ER3LZXuFeKR3/tV/tj2hYyvHUHLYdSBH50BJ1XBiqHH
H1TFa7sOsKwxvhYLu0hd9O/SC00E3XmdBgp8STMAMKR60yydixYZWO2jlaW6Or9J
hticR7NVYk3949wL/5K4O0Kad3dpaxjBuj1dO5wCfdV4slER0JBPfbz1g17AEcIg
pyEtNbiwYQ64/HMC+QSUqe1wLaK+SaDexRtquJ1cUtCx+nGtypocj594JiTzEAx/
dBJxDgcT5zdUoPdW2oyuxR21q1qMXWWjzDycwdxlGyiF3+xCHWcfGrACJA9hi3nC
gFzseuTCmDaMYO0rFEYqkcAAIZ3C165uun8TvB8jVHLiggoITpU0g6/cDDOAJDej
c1vU+CfsF+TI0MU1jneKqk183E3T0M4geYcF44dAi4K8mM6Qnyf+dzcmO42uJX5v
HkUpUAhydkwXVtSbwVeM6NPouTI2t8gAIrZfYKMcmIEUYQY6I7XR+m64rD2FO7mZ
092sERbrFf3zWhnc34QS0rLJkEDFp8pXMsN4cg6wzN9nb0+fTIGxUppFjaKHqX0K
c1RkHgBu8dH8ZC/CtzIYVoec4WOMePSAIQhH2jvTysENP9/Nl1VRwbdis8ebL26j
BZqqeIboFXef6o+BxFAqyYqWwLpP1/iBmzDew6HhzZDJRLm7ApbSg6A0p4l0qaHy
CK/2/Xlv+WCjPZ1/gQOqivG97whe7qam0/3DWAr+CG5Ypfi28/Q6CFpqj75rxtFg
Al0qB5NCcm0LnsxZQK6bCfTj9phwzwcy/j/SH9xjV6DbtjSvt7hzj5s9cAMnkjqf
azIzs2j+bGSnU7HmNihZVg8HYrr53/4NeuOFOxQAU45dVt/lCoqGWp915Ww2wpxN
SpzKNl/UZP2Smo0IUJh/4KhEpsDEdJb3gN9QAkjae1w3CQC1lu1jyVjmEboxphi/
C9HP0e3xK8J9nj+O0mEazDPPHyMNM+vWG7GF+m/yh/nkWPjPPaQ0cfzzHQ2h0Gsv
qLpiwCPcbboZESFn9JGXwzBUmviVKJV0njIUQ6Ok3U4mvpK/SdGw8P6a69EMheQl
m+/Z0aFlrGrMN1XSe6eFxfZ9btexo6P6CjgcaiqJsAqYLfZYzX0Z67kaN3shmWNN
R8WY56NkC5wjsEja9EeKX6HwPU85XLBSpfK6BcX/6pdJSiStCTrZhHlwRj+QrnCz
CY2DBYACLtiAO2dDXbddzl0K8PBKoEp4xigygOLUYBxcgltj1annhHbQ8mMWGCnv
38gclYk3qa4OZH8YHUHCCm46xpJEGt34VU/6qGnMjTGyWGhGp+eVms2YHBHOrnqT
smqEnBftH/mx29ZJ4MOX+WPtbFwYOnW/Iz4D0sY7DG01G959mLEc4JIb+76zF4Oq
HDe9hcJKTPUmM+ppVGo11zhAGdUKN/7AIf4GmW9BasUylh42PX0r/O4RXhkGFCk8
73AXoelGGUTsxiCfT3d7u2SMppSykLeCROpLsk+pcAeI5owqrgTQrOk2rH4uqUGJ
nPOCXPwV3oRjdB6QjpmY72JtVWzoeWAoA6ZzLxAS6jVkp2kGTH2f/WaGF5pTT1qb
iYryg/YBxgSmfwkba4MJxGTVlnUKPsStMJ2Cpw1QWSlY79tKm/hgRf2y7TrheRyq
4MVGSrecv1omzRwHSzq9Yr1vNxyrPgkDtQq0eDSHUVKHPP2eZ/7Z4YUxFZM7WYmQ
ifeuWm/eJNDVVL9DALFs786PP+6udoPUD2GnI7x8m1zwqQ2emwtgq7TUDtHWNNa6
fmBVtGXO87NUFAM0fxGe9lDW2w3LOLTVcMtJWSuEdfSTo/m75HBejK6HE5A6PSmu
xXeybZth/j7zT+0qsgZhW6a6dvfVutGMlj29qMmekVtl/dP4YSixfj1ltvUtonY/
VXdqO1kdjPY8hK3L3rSV9EE3GqxAforEzvSYxkDvhceLOXXEqvJVBhVyrYlWdi/x
ffCzLhN0LG9o0JdAYGytMEUiFfdhqLysekB9M2e9b49g7oP7/OlFzcmylmUcPsvQ
vHkw5knWv9w0m8qLDb3nn10bMzWQOkNn06T40PzvCm+f3SJCgl+LRLrUx9NxayuB
YWUL7ZL7g8yMvKMt044nOHk5FsizU/jGmhscSaYg52a51+OQtrMbCmiy910q6eOq
4ncwFFbivMu426YlCVdDDSq1+uBmBPsUxIZXA4TTnnfm9Rriiu8YqBrv3p68CLoT
1LaPmQnTNXyPt4LZEEdrPI5kXgyWLQcLBRhY/OU6iotiQK7yFoGrcZ1e5S9N9kRG
X/BBvN666P/z02Q9J4Guaa2CRr00fkEs8/EJEhf9AdO2k8CP+P+GFzVBjYMRqTaz
EoRfA4iQQN4bDS2aR/hCzTQFHng19Rwa6+pPC597UIwlpaDAldFGpDGsm3OEBZZm
azTZ9ZsByx+sFKAGrp3SpWXdJONaQc3xVDKn1D+goqDeAIHLFBKtSi4PCW6oD819
/JbKl+yqGMggTsXuXlUwNpXsXV+6Vb1a734+a7vxbMT2LjaAkzQXtV1vCwH3clnf
NAVUr+cTI8zwd4L7Dp/Xl3eU8lLUoIzwJKrEMsoafWhVGslbJXhOoA2Y0IhvegMh
bb1aJXrZmhC8TxJnh4SSPZCumXT7KMtpAW519f5pAVdTDtwtneWSCgDHBEPyEPXW
aQaUUonMhkPJqqfRUxQ5vSeO88IT2eGhLWXhoVSxcRQzSXDUlbKOLD7ttD5fufyT
zHcOcpPzjLZzzXNcy4IIBvQq+yewt0sy8ssou+/caa2/k7rv4/zIi8vKwhoetSFk
ArpRES5hY86sx6W0LHEHPoVPN0c1GFxCvdcWIZrJh/S1MiHeiytmQ9raXZ+0uzvf
Tnp95Bei3s4UgO3KyXaSNbZYgT9n8N7OlvvAuGosKkILkFQ0pLeI4S6tfAnXfrh9
8VXeXFXQTLQDoiX2W6iz5Femhk3q4//EXK82kHOoo8dB5hVsjN6saNGr4s04c+Rf
YrFbGS8Yg+ZXPRyBaBBIb9mIvf25SgtPUgkGveYTd9d2NKuIfOzk58E/K3UhoOBm
krqIyq90tfPM+eoV0htnnJTv5QJ+epm92QNDefSw8fpAQN6Pcd9sVLPfqKpQxW3R
4mmVHeceNN3rvvFZvdh4+FDpl5Eth+b67UVomWv+cs/f3s/EVKhMZxpeYdkUPJyz
XQQXtTlFtcnLZYkmOk/JK8Rl04fWMQQJbkJ0MwPPpaRFezOZjj96fr3Pwa4lRVDS
+WxrdBrM1/0SWGwJ1eVr7AyuiKhfRg9SyALwccZYVZ1vxQbyDJ7guVg/xyR6SLoG
Jw75i0ZesuRPWqACT+04NoTPmZPslwPpvqpr6XrCSrMdr9mrkqk9FE7CX6P86mlj
PXdLrisrjQMF5mzOV9zDflfk+Wsi8i+QyH0a9u5/QeCiW9EjhUFxMqwG1akE1gvk
PlTRFHDojbXYA254LjrVIQOsgEzJlSbQZ4ZM8Q2eFbvRovYzkVN3EO7/AKeoEfQ0
nfpT4QJop/vNZVlB4agqA5mRoJs9e/gxCKfUCTspcl7Wwe9Vq53vXjsrjuP91F2h
FL8M3kDsx93YgQz1hg35ofJbifi05s3CDx7vQDxEbUS04DYl8I9rgCVPBDDGVoiT
rLDq/iy/UFu7ByZ7WVh6HdRqas0gfg6PJ6SzjvM08ws3cq0NEG9pecfK6H/Fr5lp
96xYNC3vhoFGCCfE9FxFTuOjTDgdhGsIy+r2qQDK/RXIYUIX0epnaYW1w2eJYjQb
efvyz5NdyZgiRdLXCorxTvEeUzbfaJqMFAHOKoWnnbLPg1RyImkGsSePwmoWrt9Q
S0n+IE8X1C5taY2Yk2tCw7FZg2XJvnYhfsCXL/0444WMPnBJTo7+CNvocr2rU/AI
ln34EHQm+7j+tigbWTAoWLdU2OSJIBA08lMClyzk+DBbcEG1JKWUWN581SzEo5OV
sXK1myIGn/nSsSOEFItRndj25G51k0QI9/z83rlNROlG1z9qCMwwQoUISuFPxU2r
WTg/GO/f8qKkx9yNv4XN8oLCRoxxJzxUEPuNcmAOu2CFYenIHWpXIZC7xdPOmZyn
aEky+snLf6JWVgW/MMgCotXe/xUdJ32F5u65tkwrOR0JcEp+lYX+Ylcxhwwd94sB
u0wy5S+UK1jGzpTP7nV5ENCl5Sw0pZ7LLXROUVu3faWmfbdE64hQtTa+Jnfv3Wxn
5kWlmsqgX8F16rw+wWI94rC7xOnOGcdL9jhsW8I8ihhV0xy4hfHQtZ9OZwcrv4pQ
Ys3nLh9RYnY9J24zsWJZTbhUAOwoZDOa7tp9cjgNQGIH20CtfZETGv74dOqNbXuk
GLjXiobxzPRrZ85+8c3ZQcNtbn8V0V9dPIZtbvOgn8/ltrubQp3HXxx1cWL2P0tf
YNIZsfiJQl84NKVYrG3ymosr5ndTCoGHBTUctKZMEyP/A89DETtM79pbQtUvT/JP
xZ5DwolQ5oFsdDcV94LwS6O+mDp8mbleHyDhwwE3svNjNIW6XJX67pouvJVSfL5t
YQ+X58PXaFmczsu2SmPMAkz7JPh4KZwscK6PfAjjB1Yh39kOAubTrjVwKzggBe8q
w4WWYWoeRcRXtGfQG/jVsmRsmXQ95Z75LTcB4zuFiQTCsR7VnLy9p6hfoYSRQrdC
E4Dyni8iAa2iz4gQzEYyFhTNcXYuKFUhNtSOCQOLmazBVlVJmt9e8TwM8Sl1iPvk
hOJQCUj2NOhufZOsAtSod02p9UNZyVQZQed7LmCKflFx1Cey0sCRO5zqxL5rW5eZ
6YFcuGg8I6uu+klm9Z5Bg8X53UDEtwcuSgRGUosAL/T3nwa0DGtPxoxW6y4Jm2pC
KIWW0r36uMjhV7j14SnmKJvtsGR9It2+e5hqEeK0Dn1o0l4LrHw9I1YhtSCBQaA7
ZjEWIaipxB0Be82aUH49UusY5i6O+rdViE3LKLa1FWC+5Ko3IDx0iAj/JMMwJ5jE
Szukfl9hNCqY8YGd6d+f950tlgzpaqHvSZIsejRcJMt5ISyWHl+Ic63wt0DhGgjv
p7jm3SXp3QzmSY7e089qz9LQ/O0y9MWaH6dmpa5rjMKXZK6LCNoxoqBqdNQ6aYnN
IIlhUJjamNQBfYV3kd9Osb0QL959KgQDGCv+YvmTiE5VP5WMs7NJruHaa4Hvr9D9
/0jnaslNGN9RVukGRywLUHaDqXgsNNWclrX86vQqGc9iANY6Kgcpu7AbRkuxvZMl
NMe4XnRuW3Y9E0LIJwpobyJ6eiSWlj4pOU02FN3/3l2uBUV2+Eu7//Ws7nAVkIOd
NXdykpAQWBx4+1uuXgBeHh/a+b0hPFYIFbTglWJnm/5lnupiqC1PO5EWDq969nue
WhFLk/42DGkiMnRbngtC1rPq79hppSNC71aw+UWKrWHmDgM/hlZ3tU+Wy9aqZFmt
kQZOFtV5UQzrV9BEwOgmF8abw9PBlOHLjSbWC8mW+KJkEMIQIXSlkw4UgIMqnXet
28VzAtZlMfAKLFcmXfbYssrsMAMziPEt0NRN9jCel7okXPbqwJdOIUU+lPL9EU01
Rx2UpWIRhswQp4XCeu3T0lHD64OWVwx604tyGSXSEaQeiRRcHI0KumaEeWYtAfEw
Lnwl0go/6zPeXT07fE+nM1KOL4cguAKu0zFxZSlwIeqkviz3zKHSJ3Wk9NG6rsYn
ed+3FL/TU56H+o5fSmVqj+U2pPVX2eST79lN/M/Bz7sSqK74llFaZE8wMs8Hrnei
fXlgNhks+TwQ1iUnO3Cmo7ikjWEdeRNmtvZRCisLCaSwZYLtSPx7saGQykj3MVnv
MtKWBic56KxgoRLcUpQ5e5dDS1dx/ha6Ag+TZy1W7mPUIBjCjSe4b3f4YKNrEitt
rmny7o44s/eDKyhWmQBY3e7Cne4+IZ4ZD//AWmAA+ZpcwUFkUqBiLj40UeQ102aE
ptYnNQK9e9/CgefJwE3EOEWanfowrbJPBiKAAIJPpt7nPNnstpkgqUwOmNbt56QE
FcKd5dMRaY7vWgAyphKT4wUDRpmqkCHCCH1hdMK5Ygit/HxOoWLTrxpj9kK1bn1A
kVXVjCYne8IsafdKqDeLUM5+TJK+QGcfxO7etKZoVGgOTftZJtwINjXh1eyNd0aC
R560dpsWEVqumSBKM0g1dJiOrc+3SPMpxOSVvHWFK9pt5m5fi8OqHm1KZ7OENbMJ
AedCc1ePLMXJzw2TFFjatijf9gTS1vMFx6FQi39HYz67KnDrmBB3GiQuOaRC5gic
bqDaAzdWcKwwicyEolPXcC33hrm+/cMw2X/oPo7VR7pTMF/cAgKwnKRv9LQgpzP5
IUIsGTn72D7AjMJTiH56RE8yoo8FtJ4/leoSuprlC1Jy9g9xAtEeJpPclwGH/3bb
HmaPn1kdMvpr9PJ+G1n46Vzmrp4sdFxDvilOdjEhCh8FFQmKYzFKsb5Xk2FAlsr7
3Obn4pzt9T916z+iZQsCg1DlbRHM9lraT1j4FKqBipqu7kdOpVGpb7ClIRWcE+0O
4KUWXu+lUmsXsDPqNRdzK7M00HFFEhSND0OMlfxt2Ry8CFOFHUNIy2YddDCJcHIu
VxrsrNMt4GgzOVP1IfgK80hOmtnhcAZLlkLBV68aZigE6U4vCcEm277DoyBqJA83
z9p4LvPN0EF4JfjWI3p992ensgTqHm5EOOpKYUb/cHJb2EgOR3BTSTdwOFsYymG6
T3mX9ZdGjkl2MB/FmUuHmHMEkNGCVFtRsUDFJD89Viyt5g5IDwehUNTymyaGLsLs
HX+qNLcdqVNaOBVXm5S5xUxGFKLDFu2hWVr0/bPtuzDoRU7rKb6zqb0cPz5oNJHb
NqIpw2J7REloAi78hAqsLAWLVdPica/ChKF1lgEWg26WQhNQUTjQAuymrAfpQ3Q+
zHknuww1TpFQtpW1ZwiffmFdcVkgrJR2RtgMnQ/YoJ8rTbsuObYBZ4kEA6Ae47Wg
hO412ttFKGGgp3ZyvTibyvubs7V3v0O4MHEk+zT0OXXjOxz6je+PdTYwPp8ULvqn
DI6C3yoFGYFYkBHVIqWmdnHaBy2VwmIx0ak0ma9nnd0S2UIwS7cFa0pJs+P5wxQL
8xzf/Vfl5B5jE4jNRx7Bq0efhvlx94MKGlW8Rt2HWybsr+b04BAB0WaIlQZ6v1KR
O5PrjY/fDkKxieB3VTLNnIUW81i8mWn9wlVfM0oW06qrBqGTnAgYc6S3qbypOYGp
WI5T4h7BHVH8PMWLT8Bxtd3+uuvUEG3GWOY3LA6RUfeOA4GuQsUToZRQpj6csMHL
5Sd2/QWLZ9ahiZHT0P5gW6aMfcaQG9C0a5RfZSP9pWPz8T78A08frgrqBz69HSPb
2/3x5shjfwkjmmYScGXKUJuNNT5F6MkayYtJ8CmD4eDs99pF1HOA+DaXUjjBR1pi
iwACybtmrySmHhRdqXe5xkeG7MP1c77u4NaSrD02+fKmB9GR9MxNULk0UPlKitz6
2FpwLiAjl7Uc8puuB/zRFUW3IQ2iHyFdqe+gOjZViE7vMkqcXcw+CxnrbHLbUHPS
po2PLpiHX1+bh9ETN/SG+0F1SOv8+IXgU41j9KN0TxxZC2dV/2vSSx63AUPelHvB
T8LftazcFgjGFp2DhhE9ahSMq10K5MWsaxLhEG70k3a/jjRqKn/onsWS+43Jh6tL
5gpnAL8a9dQDh9w4SNk1p6R7FI87Uuf8E/SYHuBKJSrazc7YkOgRBj39BWnGUhdH
IG1Ryo8sgi3q5DDGLrc8DMrL52fp2YmbTBUEu+seg+/ynJMk1HkfHuNp3u8/jLss
WOeoZUSoAUJgk1/pBTZaT3jOZstfAmiVDnmM5vk8uGaElw1jkSXXbBs2hVd4Eda2
c5B+4GVJyzynHofL/qP5D+97T+oi8GaHk0k5Riee/+wo0KhHKMYWIUj6vF332dgc
puLhSfljN0/UeedAyxeb+sM+fTpeGWG1VN/pPs20cxLF5ivfw+4tjOSG5LzseO0d
smBpsHRrs8sm4pYoWr+eM8EF4jgno5EQ/2nfN/vNtsDnVPX5YztNMP0b9+UE5OEF
Rt0g1cUzGn424cchsd5H8/7bKKiSAJKPsvUazq4OWClG3xi89s1zJ/cdNBszFM+E
YoKjL3HEtsstONkOhWtMpV5Uu/4O5nOzjjjVDy3BkEMVTshEOYg0qkNOIvA1q08d
fTvKnckzzAzLQvjI1yGGZNZxy/9VXRHHYJXi9D37kPekYBeqWlMctHOBwgdwB1HG
j8jC1UMGXPRjXdpdwzStH7590Byn8ZBxXSYIkXvlF62NvJmqTR0BdBZoWN4/EYz5
U+r1AGmZXWLXZwpdLkjVqnuKHDDOfqH788aV2S067rLnPpPHM1sZOwZKTY1cMIO5
pV71ILdwflCfIW+PPD0st6KdmkxQ+/gzDt+g+s5Gc8VSMrlnTuAqlwY2rkGKNgFf
3dAGHZSdNNHb8Yrf3VLwlidzt9fErzuxzIsmmh/rkh0tkquOLn0tE1P1W3mni4TV
MCa/LHkNrCJLtH1sB7wibllLq6HUAMDNb7bT+zZTtZpY5Y1GOJops7MMtig7fnzR
8q76CnyaML84oXgv15t8XDOHLLiHq+2hUxKfg5o+tQjY5jA3WEwO6SfpMFbL7gzU
Bakfwu1glJn5Oozszqil8dNrhIFPr1EiCdzR6qztz1z11L/30AReSJK3LL/eJ0hU
ewqWUmQK+zgr5gasy72bA3MFqprhLSauXeRhtdZbMESITjrvwV3chi8yu8ov51mS
ZDR9Vw8Q9en3o+LowvmijHbXUkCjvRd/ELLnpwQqIUXh/PeI05OIlmxlnI5JEn6X
UsDeMcMmd2724o5jo26WjeS0G4CY0CXvmBVK5AHuLCCCXkkFcwkObOZ+bTuzof7O
CifJoBXjAE9ItLmH+WFTShRQCTEAOfzelQGYk3NJK05wSEn+M/wgARWIz44g72mk
aqXsJtVlPsg2S+cvUxvvQ/NF5iczdCQhr8teUzfduvycWHFT0Xh+ONY5inVbLD7+
vQUzmyKPerjtrkMvGnhFtklgAUr8qTf7XBH+Yy9oWkSIlieN7lf6U2KSi1q5ACIP
i5WntYOEfKVCYlGcGq64TInJ7Nqj43YuoPZMt9hhBPy94GTLe5DeQzz0uDVbJ3iH
3zBToFZieZK1gWA8HIi+3X8skN2z8Nhy920pJwKMouBbW8B/vTDYt+XlJ1+U3dSX
yS4vzuWzf2WCOiimF04+X8mwENJwWKV2ccZY47/SDa6Mf/C+/e9rjsVjdkXLA0/L
cubLmx7WXeKO0DcdZ+OWgeh+h1kufRqUwPqbKMNqQj7Z+RC99IkgAa0+e5fkae1k
N7dO2r2vNSZVLqpFbQHIaoDPOiyQe0zyUWfOqk1OuTx0aWhvVsjL531I06P5Q1b4
0n41NYaUDKR526UE5ZZPUv1/L2FYCOycgXBRTcHoHscd9bg8stTG5bUltOel2uwo
Fdol6tS8uh058f1P3wmth6bHxRUdFJrff/CXOLUgGf1qYrPStEOC/GGGBDiVZvq0
tvfvoNPATJB41Yy7TV+bV6j/uET1nBe9GHiUj84yOVKYuYSlnsFx3L8YocmS0tt+
59lhg3IUsSAvhO51zXyXIdQ4iZh6PpbHtQEmM7NyE4awsu4lFXd/osyV5qy40b0t
YqXr6CmS3W3McMruJ16yOLFMqS00ECmysYku0hOG4Xbe0bYeUzgFWtEhAcs1MwGT
tWeTBmEaatLxTDlMRTCuNnAStIcs8k7l82MwW8Icm4e7awPoZ6EdORC7GTp8L0gV
oME6RUt0/PgFF0TEAc9hoiV0cVQZONsqDEdALrs31wqnu+GGAK8OCiMvTddTeNs1
fwWz8ZrXzzPwhVl+9wEm7uS+sKeWqriL04ggYhwMXStomRWpJV3/hHstRkznqq6a
KlnlrknWRXbblkiKc2/QasJZqUduluJXnz+VL4kDbg1DqHVlWBS31bNDEMCLe2gJ
g21l0K3fTSttwdGyhKjqtXTyLlwAUF3C7Z1RE1uSxb6PTiCbu/6vcujFz/P8A2Ui
cfDwICLqkOUhDVxK6RCscGIny+7jP0q2vWymhHP6Vv5F1FDjk/YhwUBwr0OiwzrX
CwC3QsgvvPhaM+sSx/TuvfPGh6ADUsEkpSvRVTFAokKyYZmNVqkyILPLg75Lf/Mj
9pTo6UDiSmh/HnfIjeDaGHwxVg5HA8ahaYfrwtqEsr7+FdIxNBHkZOc3O8dKA9uv
kCNHs77DyCYbvxBW9FP8ohw23EbO+gkl0pk1lmyrMWGRBpRo+5JQz2H7+ZTL/WC/
fe3+a4paLodfnf13RXoTyriB7IfBs5S/PCD0gEd537XTJKcvRxNhGkI0T5GDfsYU
IhaJ1087Aktg9Gzg39VPpdRUOJc2WnFX0IcC7V1J2leoTAsOS0oqIqDgRYeuaiz2
n/PYdPxOMukpYtxJNwmzCK6dOIbRlR9j8vGuIE5BiI6228aIwoRBHOo+w23S7czg
eT5uqAE0MbBfq8OwMqqNjwaj0RzNnmI1V45VWPF4gQCfwrs3Esbw/O8gK2IBKObM
y8BBrgY6bSfX0SS9vD0BLKme6MqF6D15OSB4YKi6Ao+v5tbVqCe5KKC1lw7oSepG
mcxYry6vY2tzXIXnGnqUNFE/mHgPQwRV/btM6UavdFXMetoTEd89PPH1O7lGcR5w
DFLG96Txru1jE9bJR8V2VWKBcwo24Ep3CJPkc9DBRpVrQyHh40cmcB+Ib/lUnUpj
PEpRgrMqIalPTx4NGUtKx5vWk7KZyWpA1QqcyuM76Uj4THBZ86LjaTFhn55cLwlM
/ZR1x/mUFUfcrxcLahZ9i157qdmgbH7yTDtNygoOIB84w9+b+iUxCJB3m8sUty2X
OWeNe4VDjtCPm2SeX6SMWEoHay56NKo6Xlw/ahzZg5377O/ivBZe8Z52wB3QdV/K
qUGPGk3ZCLzVtbgIcww9q0+Aw1b5m0MelBAykJ5xfo23fMUzhBmSdtj9Iu+BXieS
PWGSlkhFbJOlNOrLfufVrkbU/MBRfOz82bn2vskpbGuYMAgeQ89VUcC7pvSVTvqX
8LvlUWYZppRX6Hf3aXEH/eN0FksNaHclt82Vlm/ZzvUMDN9oXsvI6ItRR3CSbeM1
2pGzov1WB53LqgGEO9bBcLb7qMWl4R9BxXMnhkqXAc+7qmyVoWABu0uIztLRjjpF
0MFpJYy2sMtn1tdFiSvku7+IsL82s6s13MUxA5jssAdUFB0Kn8z2bt5g3RxpzK5U
CDUlUN1iQ6jl/7n79jh8+W/rNt6LdQHqAP3zdvzdvl/1MZONWHJIKzt/062D82vY
KdfD4QGJrNR6E3Z7W/o+wZquX3la3y9WM/zNavYxZ5940ZEjt0KHrva18ok4uFHg
tvRUDcI6U93SrmX+/K9Y23h9X6/UNez9M+snJFtZNqGUGp5+MauNIk+K7QfbQ0EI
FddMNNHBfLchEoqXYAo4CoUSR4lz4u+fwgv/XcbywC4M+/YYOQ+0nUFWmOcqli/k
33Z7nDZZ5EhIFTAYT/n3gXOrGGiPkycrTlMxZ3mftOkTLAVvEsbqoy0kzsbAiEum
Z7xa5weczYArbAI+Hx6HouNJhK5OjWgVYdxLjNLBXUk5vvo1JTaFyoTcteuW4u8X
vvxf02yFsuLKPyZAeK5P9le9PPn/rzGUG/1qlG+VBcEZVE5IovtHnSgETLQlbCrD
66jMYv7QptOm7L1JfUQ/FDXx8y+YXd7OKAZtqDcxGMtLTj9pV+lZusjZJsq2/Zl3
AFEsDJyMEyw59pL2SyPmmXeeP0Ux5Yt+ULSimuqenBW/NDM+jI39SMOc5UwFfrGe
pKC7HTI+Gi7JBcWQs5sx0u6L6MPFGDogSDoWT0Z0DjG632H/GoLBcGaQIt1hSacE
rRj75mxAjeI7fld1vKrzbUfrz6oYpIwIcGeVjxTurGKcFinAEkCcc24LD8xy8Jxw
guVoaMtLrKEb36WC0UIY/xL7xyM85ZqgMwb7RG0c7YQSxtjXkCbR+5mDKXuRKUsc
2gUGUDd5QiJDBEEdG+Tn4X2LIKMQhmSYG42OeexyR4PUb1Gce9tc4zc7TDy0iGCJ
0g1LGbflMy+twM0S50WwoWOLLGQ7jnXSZd6JDn+bTHTgxuuu+kAC5ffPGiWC1Npv
07ffBHkwA5cxTKK54FVAhL2o2ndiruEtcWR3Py84lNwXqf6A0LF0FD8ffakV2RBG
oYlcod0hq96nuHMZYriMCuiI4mnBtTGfbDO/33dNqihKiG51LSAmNoCQIptiOYTR
rhyK4budtGlKpRz49ljMdNJc6057pEqXHtuKx1sjTVjRPrqW50UvJ1dmxi+IShOb
WJoWwZKKXFg9ZVhEU2URurJKCyPrKHd/Q+p5TmYP5ZZ6Nm8SoozjpqJml8zkood8
964I+akbK2QN/fsT3kJhtpRu2xHkuYMDAThTxdwAqofstPcWwk38CxU9IFBrptBS
jplVGCumavIUugVsQchqNWu4t/gWUMHxCJtiyfOYExbt2uee1yRxZ5EObJT+kamO
ypRrJqbCrprxjwpwMXiINOhiTqnjWMfmrz0MQz4V4gzS2Ej1iJGzsjzXt8WCHXOJ
Jklpv3xCwc3Va8Ka749KFE0aQNqkOmo3YaEpm5av/zMgZDKNaUFB96/w/6NWcQ/J
3u8CsJIjv3zDCBa8Bj0CCaxcJoAcn4Jfs//3/cKTpjKwTTBfns+B9A3LA9zsD23K
mGaSI6OBG1UuBHDON6WF26H8bZXNwHCyq3woP2JV6Tnn1Chw99vEEaKYEXoybpc3
DHsCtLS2z65qHcUbjW/uyrpsOazc5TG8TiD5Fbk2+DiUZ89OoKDzUT6rQuU+YlfT
b8Iyuxr3w4Eb06bs0vg2wdofdL6NGjbDxCEjO9g+LJmvL71H0ZK2PZi33/E+91US
zUynbhOtndiEU1d0/CFk7s8rgeUISw2/tCDT5Qv4/BLeNjrtV630vBUp0gz3rOx/
8RWTI1g2QaeJx5Bat7egcADRqJu7pJZ2xYUXRuYZWFDVzZrY32AUxFgqH3+ZTbAo
caEJGOcqJgrpxzyZ3t/XkaDqCXXCiWNDKtVWNhHvCX4bgkWSyPsTdJOxpf7ESmXH
B/n8hHAUyjlmIZFaruJ71uqwb8QMAdCKlqsWE5Zu61AQQUmw4CP+3K4Hr5dXDQtE
Cjb2hpYh5pCihgsGp4H+Lp1jr0Qr9B1S2stHmFFG51INnEBF8OLv+83wW7SobZQx
i/5ZM0GwBaXKVwi6d+cptfxq60ZC9jfPivjDIr9Ik6upFqPSoCoCBOHsZUAzgdVH
lHhNTMtQvxpKb9PcTSOeJ02kKbYmpH2SSyZjtvXoi+fPT8AG9zjfPf4PeJ2JIuxH
UinyA5cEeW5nSR5DgtWUu4xXJF04NiDgubKfKyzcxQfni1RO/FDTcHPneCK3cI2g
y6YTQpYGc89sTsS+wLHVZCkt1RTvNgrcdxf+JL7ceIvRTR6R2clN43pTew4RSu6V
iEGb0Da2Ep9UWMtenuQQEOCU+AMCi8dkvLt8kt9UlvWqyR8RYIOkB/8YIDj9OYsn
if5L83N0AKSiFXbJ/Tycxh+Dor18WkSMGKQavXxSBBH+EY+b/2B0BBzxPlOMZ3Le
JqrwC+LV40y7ZaxWVUl/W2IsaR4NRkgy2O73R/9t7ewWmP1AklFBPTq9igPXyfCW
qwcCiTRYnJPqT8S6ODVKK55Z2zNlJE2Kk6csOR5cdjdolsJCHyLt4kk/7YFNsjxF
lgtECERTW9N+LnKOgh87VJUIlmEs+4SHeWBFezwjXB2xcb+Mu4AIL67SFX6zGzDb
y9bT0afoP/4UFrq9ovao+0+MpQtJiA/lA+p6W84dWGb2gpQH2uqg17S/nhFeLq3e
hVCEnp73RIn2oOr4oOtiSIFWnMrfeIk+n/BfeqmvuzXVPyrHBZofXJCw61mj1JG6
0/5RqLEVe2/TCMbNg/a4QiKhY20wKMYhll3q6RTebY7128SF1TMbm++Hd0j5IdO9
1K/8ySqdhcXh+BQA8ZY9yls/bbJFLjTYhPNHrSBxqPtihET/WB7EuLdOmEATkbok
h3X7o5KcU2L4kBwFB6JyzTlEMVer6+bhRFh0bFfqDhnCa0YPFvS1icxKwflhbYt1
Ve1ROoXMQQlUSM1qkVTBhh0Nq+uYvX6bOKEF0UgMFVLgNt7NmPsAMPzBawhKpuzy
0BVOApibjylD6XxfPxqabuquKJpgD+WIMBAJvZTkXYbdy1Hl/cWXBa7W09rBw62c
n3vSm/oAJE4kTHfZvoA/MGoClnYly/BQeJeEGaiXrVa5tdnGFo2CyYsoh+/DB0dF
Psci1AHscJ/ZPXqlevuZWGTVEiRicxBcvdRghXLcGz8CJqgk3PfQT6ie+/EmmwfW
/2SLOuiiFwn8JmhuoTY7RPlf9oqygfAhASR6UjYe9TZaLuaHXk7TJBirzlWWo0+5
kzk1w/78MpTIACdzTzy4m2afp1JBUBBAaXMrPvzb5CrxGq0c4h/6eMFbnaGeUr7L
IWL0NcuYx/NlSfvYmzZUxz5FnCWi3aa8eqrUEQIWV+dDb1l8D0UINNw9WN6NT59T
QhxiB1Kylc2KxLgBfGFN11sZzzICML4GIArb8ZKZsxvnB6slQtcpR1JZY8ks96YG
RHNpxoCMBvgYJCg1QonylbHLJ/rtt657FOde0oq+c8b7dDH3QEH4WOaYslGiCwqZ
HhjZuP/B6xV+uYt4tSQCGGxGJ+cKAW5rL7NcmIa3z0UG2nV1qwpg5Kw+l9rGbSoy
2FmwyPLuXYItmJ5na2MP83OKyGBN/R+F5BChPcaxmK0i7m9hx+2YeRYWTavuOte7
EcxIixv7SxCUFBqBPfeMKG3VTQk+IjNJGsWHBCUHGWPOlKcoHgJJ+WjZsdESriDT
zFXAjqrrgsCsWEIcKi/D8/ZjYRAeu10VhjcTDbzU/zBz72IdLnDbiXINPNu3nYmv
0ZLqcxcyRZNicosemqK8uBigS22eR/cjVavGsXJ0jozPAZI27dY5/kc5cIanTIB7
2aOa1Wh64MTwO1aaunZovjtAfzdBnGU6FTENLv0k2Re/YrUpFhYQRd0+rYRcbHbu
CedrsGmrh2LBWxELo/smQnEM+EXZ6MIiYBv7Szas7uI6o/yRS6w1yoEP+W4PpSM+
f5JOv/DlfbTXGiBUH9DAqmonbyswhMTA93GoaCWFu5SVF1uE7dtn92D5BQBBSrEz
tjegfRj+cd//pfTobm+MIe1PQNrHgMv/lsJbP1khJtSa45PM+33ZdI5ghTg6eQ8/
vz8Tpe1mKEnUq/emLnkm8iPuRx5dn4cDMF19WKbdAijvwzQV68WaUDNM01Gsf3/q
2CYdVXjtnZlX+TRtl0iwAn8LAMrjA2fZ6kfpPD+r0XpumAMY10p0x7aJroc+SXYW
rcJWw0kxe31Iywfhxn/BKN6Wy4uw1Ab2Kw1FvEUXVJExNd2MkR17T8rJZYzdKI4m
/ECu4j15cUyzWdI/T5rIRhiP1tkPVtX80ZuS160BSA2MehKc736RoHX6dZqwk2EM
WgiAeIQ6iPXSUle+YixpXRBauvwLFxYo2MZ/p9lTJCHjcian5S/aQTBTO7Rvp3Xi
Bf1k91BPZp4cq7jvG7941J+8S/W9Ps4b7qbtcOslaW8vNmzdtrZQh8JAqhBFEgjR
nNt1PWg2ew5Cqk1pVS9Ob4AxkcPPWSbSFg52mLUPoUGFxPWU+lSK6XHzuPGcukRI
l5/8ynQP60qY1Q0CIgFYwkHHl/axy73/3P/E/2sQjWGCZ/8vUGwvMk9YCuX0Emmk
HcYy2DiEMm8s5yflkF0bJO0JUdgq3nC4L/LBHeULIBiHdkgtenfONrQjQ/kNOjnH
3nRlnGXOpHpNvkn6RhRqHGj1vN3JA+KlM4osDakBNHanOk2qkK5C1jLUofDj52wG
XcYj1w8jUuRGHqIOUdhWKM7fv47dtR1mkgzQcD8QHdgviRTn9U7S4ZZiJyDtFRsj
aokpAiAHcvAhZPBhbxW93m5vDli9QWAhUmPWorQQScBRM5rSz6pVlYBm6+z5byOu
hYpqEDrV4JftYOX2uzhI6exMKT1CCIxfsd7B2imWJ19NExl8n9DyY9Kr+n4JkpU3
rJzqTSAbU2aZQagQ9e8TUruhzZgCHtei9c5VKvFrC3R5IV/i63TmhFPuuypsD65O
oLxr/Bs0TWNLhfpwK4Uz3+AsIqiLPwJSXBhfiCqFJyy1ArhIKi/Z1f/gFsez+/fy
EeAKPn9iP9UNP5mO6Vs+4IfLHJtwzEqtSHX+WhcWecbFFEHSEEOO3QkM62Hl4PLp
ZZQ2//aXtUC48Ak6xNoPvLMKRV2FW4b5T91YHJ3eD61oQSPTsI9EADFFDBhPfE9J
4RzUvPrE4lCI4CvhR2seTiRsV5wPpumdiNC/jhqFYOV0F8KObKjQ58WaFTgU+yBc
kPhm3rorB+jLLtY6y36c7dj7LPsPsoh/boLUPGp5YMzO69iBz9oxV15YnakirlSp
C4V7voq9B9jrBvQVRmRPKc8dTNsKtOZAvvqNmp5r5aK1mH8ryFMqhO5WAN3w4EN2
7fd8piBBpNtTzpz1MshQOxFBu20IBbmWhajlfc0YHTUUlcnFUO2+eCLyUo1Msz9M
8fnq9CLhHe0iuaSA/EJXuLXosyRE+SIFutUbNbE8aT2fqIC9hzhgZ1IuHPK+LRPV
s6bce3azoushS0+cG/kMMu6ahdi/+817zhT0E2KFZ4rkjO24sfsQ5caxM8+T3Vyi
l9V9tinxUvc3vRszPFszXRQJj7JL14K3ndyGD786AZqh32qwWVTIJdA3oSE5yo1M
v3LhxSpX2UVdV9nhOWGMdIRkFaBuNzH4EGad/SUV5ix9kOu6VLp83Zg20JhRStoW
ECNk6v58cZCVCj5nyaqLt1FA0xDruBlVxA5nqhIWYanbCF1rgk5losLPTFUng33t
0lS9r+tJUzAPw2+hQWuYUwFfFOoFGOjuOZq0G/pQEwFfXpp7SSNOirH38eUts39V
wbAoMZZjExj6IPtT6+uZIhJc2qp9VuLQi5bOr3a54OBgF7SUvVIUMtTvJNYBMTt7
nyKr/a3FsasQkgm7ki2f5g4+8qgPHXkUjQ6RifxtyoJ9owb+kcnA3TGLvIXbWt2N
mT14vTbkv9hDgB9vy/2ukuuO0xS9fLligM6XpRWujVBkVUzCfArhhkB9sxkOWDvj
gbRUF2V+yMjnNqM9Pc3sQQ0vfmAOX69+A5+QKQKkosIbLp1/nQuyFDYP0CUog9Du
yGGad3hYsy7MdWkvauSXHBOBKbXNvZU+fM1QkHKJ4edgIgDcXV9JxYjRunSRgjoS
V6CMDoYRSsI2g3OFY72fBSoxiMExaAU6W+ze1tMLICUEK33g/zwrPlzITsF3l8xn
vATBkyKGpdz9bvlJUn7iHFNrJJqb9SvbbSdgERsfAl7BGPNrlzvlGwpgbxcFDIOW
74p99ALVyyLinqtSdGRMvpJ1m9/dEJRcKOfFTHnWi2khFgKnEYRIhQQdrU+NEucw
tLzkZkTdRt5igHxstWwiehZ8NzI3zo2us41ITJx8An3hj63bC+BnUP2JEroQlgUB
snLIdErMMLWKMA0IMz7hLc6PmSHvCn0VyE2Xl4/8aFwsiwl5Y28Q43DBiV0CCHKG
d3rVjJP7Fkbg24qHPhRvcTyV+INplCn0AR2eBeLwNbLuVOqxrz+9uQl2sHc/j2Lz
McN+pyDZ/vBYP9YfOTlfW7HZBc4UWl2fs+fTNzPzKPfbR0QRtzjdHxaYPrkUnq2e
mxT1iKSpyqk8LQ+fopMnm0MDtvwW2gId3f7qF20WofkV+nxH60bDqI6xQ7v8jmO3
Du4UcXzgqei2WN22ysxqXlWd5NjB0FdqWnZRqs1FZLnqLrttA1HoPOVV3wbrHWic
klXbGVvgk29zIYYsje26suUvjq5IxIPrkDtJiiT19zYbdgi10HXzApfBJZ+4YJvG
IZlyJINRuF8EU5zt3+WSoEj0SHwMzqkvG59h3tUwMbJRvEyD61fD6y8cw+rkTRYr
m/wnpB8bQocFmb99xy8vqCYBvmg5FLMLoL4GNqp5YxBF8xs72vpb0P9Dtt2Ir2Pr
2sVceNFYDvxFg0/6fN+nI2+igDml25YA7ouXmUJIVCvwS6xLVbu8IDLdcenqPE4G
SxtCqwhh9KtVTFUXWxoPrYPGkDqqudc2Fq4DcBv+GaS4XAi4RC41EUa02iiuUEhc
Tz84ugcS15Foko993CmgYr/ecUWFgf/g/YSvqzUt6zy1j07p238rjsd8AneMBVdu
xJW+zUr5TfBU1c6nmiJ74SSVmZOcuIJQcwGIn877PdJcGZ83a2ZzgpjH7ylq1SOh
5/A4LOJLATMKYSyx5OvwiBDIVVc8ndxSWB+AoWwxKqigLH3GfXXGKibsnpLGDqAY
6qKFyOof7bEg4+SrPSWG/lzcpIuirzNhL8oIEFKMLQW4leqEBSoz8sF8fvH1cvbF
qKGcXMbWKjISk9D4IXwc5qu23nelFx6J60+d+sEs6+vxIwlM0YCOQRD43KmGxtlC
dpl+Av0PqNBL4quS/rbxf2qLoCpF2Pp7GJuCaedt9PdwUdXVNn1/y9vumK/2sLZ3
K65wXYprfVoIPrae0jzUME+Lr6FlhyniR2R/+EAtotWg2srf/IqqkgVE04WWiw/i
WcOhkHTSP4hfNIABwIOcR4oO2Z+/IeMYjyJ8/ZgxevPW4s2BcohETrU9dHMbCkmQ
Cox6XsXVEEtnZGncSnnrTp0Ayb+9OmZHXMR2ZRHyjk0u6NMmM7oWtS4Gehifett/
HzoVhc6CehwqNpgJdXE6rL6X4jzG5N6Pl4lcVjkZxzPI4GfuX6Ame+8bs5zhgvMX
trLJ2+M9UFM4AjnCYumwwifAHH5PPLpsK4p0aJS8+sdBMi2UOgmTfNdj7JTrIfTD
Lvf3ECd8cPeqecbI7U+RXbB+7UX/GN+U+t+zfB2B4EMW5kLVjli9vLzxqyisYuMv
DIdJF7LGqsoLosTTGu3DFf+7NBg8kvVEQSs1QA91BYZ8Oh+mFHHxPvMmS5qcfaiA
s+7enNnONIyo3lonS2XCZ/PzUhIPMX3hvRybX42LCwFQaN52u//A8kXQqWfprSgO
lxRqevFSGNC9ITJbvewh7OQqKjSGqvk6m8a7WBdte95+jMYtK62S0hQE+rvQkfz0
g91XuPf79kwFnRvaRgmXvY5XvQbC3q7SvN0dyz/xJyX5d+CkMX7l5CxQqDy/8hPi
teonc4a7llE0cTFYSz0AHeOhVgr2mC/uRsiU9mKm7sbJm6jTzwgLjK+47WxBW2oG
3Hx/RvOmYRadbW7dCH+Wru4382UuO92dQNMziNnUxlUmjMcn+prsOS4+hPpHQzPb
JRr2sVvjV9uLksOkF/lg3tKcWSyeuiJV1f87GuvUjfBwX/MXWJ3g0qL1gGo27MOp
h6eNxT70+81N23LVE771lHIZcwdd8EVjWNMukEFOyD673w+G7FXdDBuYa0ncM8DA
Tv6NG6+mQxakXh9xTdI8Qbv9YvZOm94AQQixj/8zDDlLkNSqCOjl91Y61lXX4z4k
hXoCWeP7hYzmPneJE6oCCS83Xmps8v91LU8O/Uu4BoagD5BVZtxaJ3UCn6L640yu
JbVLN59dRrvAm1+0RkRsAFeJc8NOmJ43MMY/COTQqWR9bIdoQJywOSDJQuaq1723
aoUU3j8Mer95zP1LIs2bvEmvwhFAhlu5mqnLsDqF+Gv57DlHnLSjvq+sWQBAtFxv
QqHGwPO2xJqzxcJZAA4/Fpjtkj6Jg6IO39KQQksdDLddp/Pr9SSEmyWVBfV18q5C
VRrYPpEAOwsDHkUw5hTM0GuIS7p4xj3sErcWRavcGrOyMbXrLVuaVurv8sM2t/cs
jhpC6lADsppWNf+xN0uENIy43PGvBm5StCrM4p3zAhr5ZS/z69NRdChXXkt5zFCe
CdTAXQGwaJfhN5Etja38oq0FC0JjIiOtseF7eGmioop+izUKl4l2JGPD8Z98wDf+
zlStzpqd80rjUHVnC8reiKn6rg43tzabo31JYeEPYPndnOo9v0yQmzqvpxL625lo
m9eRmkihmczKOa7acIyUWLX8EcsTYtGDrLeeFmn8fgMw5jIPlBs+jmBVbf6zCZ67
7DJX7kZYR+ioFTaUufdh6z3m2jtZxJGgMyImfbs0Ttj+GgUjZCtqGjQB3FRTKImw
hbAVmuukC5n6hXTxfpWYKPiODZ+tySA8HK+PTBHGEYHFKhJrEIQD41oFAnel8GUP
aPXzr/aN9CZGxa8FE1X8ntY4i42HSCj/UvkXIINmCCrGHPQCRwh1S+jla74rZM6t
D1VEqDvxxhxKs3wMdIWTszCqTQmAjKgpU7oTJ1Ax26A7Dn/vfGpfHJFmoFi30LgZ
knHtFNPwFFotiRAEDP8Rp/PTwXC/HNdUOjvpg8f9yJQGFVHzy03L02mQGqkfxccz
VBi5iHLYCLc4gF2MFHRW/X+BtFqJ02wLxrZwE31LmUj3Zd3PdH3dJeWVaN1Ls5jl
M2KRZot0j7Z5d5UwjuJq4LHdjEa7XYIZbUcbBJ2t2eAyjIP4xbrs0PfXfXp7A7Ee
mwHc93F1hbZrHjiPWuGSi/0P82uxf6pWeSqhtVW2VDETL7xB7Q37b2/p0UeJyM5j
StzhDxf+o4j6WkzMCWGcxy6e9RhU2lhQW/CsDqs8uytLLn1DAziILjWcJdBETvDJ
Tx5sYSULaJdbci/0ZVeV2huRqaw4Yk0NAdMpY/KCA3EyGzF+qzaLBgihw2jNehqO
0nz10zPRcMEjCj5meuzh2aQxIK0kRkVIKTRmUMOMQzRFjTvzYRnztxbvsb/vcaBE
695iz2gFG3iXHAH23ixDPfms+wbr88bjl7yADaKffGP0XQHvi8r8Nxh/tNGd8u0m
G1YwJn4ht7Xvj+DUhdZqiT7hTi/hIMsCZVCMjzvkdiLJY5g9wecb6bXpP+IeMTOW
vUl3nOc3ikvirADuqj6x2E603o+xrs2UDBW6SAJrprb8RCgnNYxPiXAu15124ItP
thlDoO55efovTUIGUmn4u+9ShO2ybKIQv2ol3xZvmx2q34vjO87nKnN03+8GYYSL
YsdAnJicM7DHbw0djIBgVv2WiS2jBwNyHxazOKAhUVvT1hQQP7iMqscHRRTwVS16
jk3uGZ6aXejEb+1AEup2CYQl1ZY51EqRheJghJK2crJ6Bs1rXFQ13I3HPpX9U6H0
iG5wZS8jcS1nbbLWDHNW9/QwoE4sdpP5cWO4Vo2KDEPW6gqDgX5+XCpuQeTzSI7H
kPO+PViLXEzoGn6PdvqsaIP6TzCOg1nvTqDtaMV+LVNRufKNEHhPW1CjII7GP7SD
sqhkxattWJHxkvwpNIigwJMBA9MTbnOOKje/FZis08XjDLQ6e4ltsXuqY5lIBVxw
rzwibfZkvA4ceAIgT6UruhvMoP1S0CO7zOO/Uqz1uKIGHCGFhOsfQtOT278NiGeU
+m681eKP+cQuLYVwDH/hyXNOOZlWe+e9biLrL1aKD2KLG6Mj6B5GYTVqef1eVxfB
kMLCfeXD+888EgJXR2GpZOtsdKf78TeoDRvAx/jUj45dWIsAuXIaXt53mAha01nw
5waknLGPwpR3et3NcBbnY1RW36729/RV8jjnOEFJhnL21JZSYUMwNbDfWl8DzFW6
3xZ9J0wS9kn0uJ/tr+XZhEd+IDGKKuQQvm7efy0DmuU6O4Xw+D2DURmEf59XnFRG
LpWOwEZ0Q6nY23c/d/dL+yqeNkRDKEhgQ0kepfhi3DdZKvf0xf2VECMUjvAFpHrQ
AmCBU1zaIjoebewwssDsQWaMJD/3EqYZ1RChL6OdwQzlOEY7mCPBIiMjU998ujhr
yIeAsvltfp2BG9h7Hs7m0hQNmv/wh9Th/v9vOmGm6o7NQOqnFFfmGCs03KNg2ZxY
twlwt9g/SfHhHJlIvAUbV0B84y0fKGU6ZbRUSFdkL1wmHDpovYciGVtEDckuxpL4
tmCjy63LvQaLsftHWI4iwbD873G2ivGNnLPxc/aqE8lcBx7pwtWrhOZZxBV4IWGD
x9IyhMSsL9Rhrdo5ePMzdukCIm8VKieFGaQCv/Yku94J6P3iupXENi8Mk2+9T6Ob
D/ZWaubNmYqKPNmygH6NYbJC8BcoqgPEgGbFwLfMD9d+tNCLerMv8qNUAyXF0ldY
rMJCk0p2bBDcKLdZ+EMYs/o7263h/D1zqK+A3fA6JWBI7LkaVFGN8gpAM5LUGmm8
p45ZR/4vip+O5qGkZTckkYsnxsQZpzjHhHDM84XF1uqXoSh2bRMBp9GyCr/kVMjs
0BFJ8SgKf/5Jf65bYN9nLekhfx9CnYAIivDr4/nM4S3WTSkDH4dttJ1X1D5jkSxn
nMj/mWgMww35HfSLRINcm+mu4qfweBgk2hYUGhvA6RtjviqVbcecIG7nmbWyKD40
BOGzNDrL0QAwH3IZYYrkICEiZWyV7J1dQ1xwdKqa4WIX+PPSvvbwmYadBIWjWjou
38ACaBml0yGbkfunfCpHxNATrgO4rCdspDUqxD941fjRJ2r2tkf47li6KBEKiUBs
HvsMDbKV+sOjiccoc+7e50K9qNGDDt7PIzj47kQmMQFvl+9/mb3bDiK1+1o8Eta5
G8HkiUuVhlII8x+2etNfb2lphyam7Om+tHkmlHcgGXLMoFuhQFmg14hD5BqOxdp7
k5QFV6MTxpO4yYq2+5qCMt4zoprmq761Ixb6xNylOyeyUV/F775se3XQAPOJ4iLN
E96g2L2abY9KEef2WL9AS/cTygP0wjQrF6gHGcN12tNIPkc3udbacSd4zgKQ0OOE
qlCzt9+Zm4tfv/m96RpUfPYcem1LwNZkn3mL/qnGLHahc9Mp7ZOj4U63u4vVF3lz
sY/MfHN2VWE9B2HLcARIj+3m4OSrZj6ssINqTFcqWANQYVFm+TavNr74Es12/hEJ
MxDsJw5JqPTHCWwVgfVnCvavoNDPLQyMNylgvteDf+23JwKQm2/+CRZb5qerD9MP
8cHxjA/g4YGRHScksxmBOcOoFojZ438xoPtARzqQBQvHiQHbhMKaUslFCauUisBi
r+NKHi2gg8NKcEVyLomWQuBr/WnLX2eOlVyUuTgaZkKnmMHOuOG5xBxBQ6Nw21pZ
+8kiV8Db+zKcQT1wJnSH8OXDjV9hqenTj/rELlvKGlHjEsvjlqEpG3bnx/wWv6SY
lbZRGHQ9slXR34ru2CXEJKPJacBX+mHVsLsV7Btm4YWQ3e7ZaUkeYtDGXKGrA9uh
FLNg0yd3Zops4jQ7jFG76egCuSvFxcznLQWW9okopE2x6ovxi7jrEr0zbuQiDPlu
tm5bharV/oefCDn9mJ3THMB28ZRhX1j+SFa9xCDrThYso6HK4di/SaDtpgBpNzuN
+rgwcReaTz7by/nLjyp4zh4n3x1FcPEU9S5Eu7r8j2779yTFA0j+osVwLZuoMlvj
F2lrOlowFvTu0LHyZeWF243/mdBM/Cy8IHBsPLzgwJNDWQ+LA6bfF7ih78S6sbXG
MpTgo+KUDOpSUYffI9lLjvT5SdkSMLPoMloE0M39JYsuuty6DODG1+gR4bnmUJkp
nsKZYcRxFjcZejH2sTSXNIiIxAXSQrsTwYVaYqjUuPg7x7q3+xbr6Vz+a2aKJ8rT
t7AVTNVf+jU3opO01GQob4v846LS9Is5K0jZSEZxrfauV1tmwQ+GRQM2tEK7+Qf4
GoD6D66VEaleujKxI+xevQzGFeULUjvSwzCxSY41HG0nq4Ohb7ulLCZdfT/YNihp
eEFj2i2De+RyknB6RwiSFb+mq7kfXfvgvW4z0Dz2FELSdCkMSn4FXpW7AqDQCEkI
yZfW0daq5NlHDFYBWUnmMS0Ji5wE3DPTRmkg9xyy3bsqjE+GH086dzLr26UtAnPy
Ye52nGUINJB/6zrx8g2MZEw/szfcuoaoKvP9r3eQYCX4/fktB8TrSqsvxHPEWp+o
+TrhYldknWfDvKyPS6ufRg2RT2FYU7pVAWeHQ5rDonEUHKzKGK9NKNqNsPdYeL+s
Z/Ihc5cDKUCNwEywhyXCm6Kqn/uYmFDqBGBtynKOvrnmXK/W8Y12R73JGsBOT6fW
0jX/Br8NEn6BnapYrddxLWE03IFyF0b02re/rdZKqUBz/ZHcmJsvJY4GKNN/kjSJ
5UtPJQnUf1tqY3Q5IArPlhZcShonNKcSxJlp7kJq7SP/z7ip+ucKAdKLE66Pu74+
p2C7iZsJnqoIcuUxNyHULHR59TzIPf1NwfidfU59gQMV/om4sjn3BKpOB9NOOufq
QO4XMM79YS93dmwjkeRts7ZEHyICyULXMveiQP2WcEJzDJtUowsotcSosJsGbM7b
quSji7d902MmQNJKkBCk/4mluwbPJVl3fp/NziEdIoVxXoXxvgaYxei+M1XgEwOe
fCw8pRGNOuKupwDPVjpZD+MxzmsP56JpDv7i4Jm7lwVARSDi3tshlU/uhUEGFApj
QhH8Fw1Oqr1xeDADKuoJ7k9pVgvU6Xgkb4T8o7/a0cZhfdbj4NgNi60EwEusKdff
6Ugzl1blE2pXuxZKe+7UUIDtK+gp1Ife7VMpzZqXs9qhbPk/aDMa1wH79PYYeqB7
Nh0LoFoQftWGOdlNvEeys+7w5ltlkRfYv1UHqd4HFDJ7iElpDadeUbQI8f+Dit5p
I64pBBWb1u67z3DO3MpZEIc9D+fYs0rYnrdMO7G9XJWXPa1fsNXtFBxOoxGH1R/W
pSHqtKfmFzbOYL71131Fk+NpTwEMF/08dS0f/HRpUiWIzVzmgfoNowTKlqwgJIze
o2VQegGnEsZ1vIzksJnl+uSOHixhjCGPcbj4Bxtv4NDa6eEm20d7kchMIxpYdPmz
QO1OOq8CicfoB3bHwg+Yd1BwcERDvKgVLPzWaZSkpF08aOvaPHzFq3RYcXqgGgwF
nmrM9fSrgAXhxNmLaNBDnflSKm0PQ+CPYJ678YpBTN6MyHKKregelXcJDuiozOSB
fTgTR85VX0f6/si8oo8eDfN1KYA2cxLEQieV8X4d9WxVJS+rKwRw/WtTvW/HzGYE
imFhG68fS+A0rT45tNg2STU9mjBf67EWejHhNCQZRnWYjkEyFwyXs0i59pKV79yr
Ur9/smOiZCmV1gMLUmb4bXaTw/r/Kc3UmLFSByWJMXWDXPaUyue+vuedvQfGHIEv
Z6AiOoNC7SJxcJ0BJ3cUlw6IME2EoAgbyfLAVZZEJZAPS+tYxPAJMynIeUk0m0aF
40inO6oVArBqelTfSfSHBLhRrPWTXuIHTq/V1JEafGfB7Z2QqaHV/Eqob8HHEebn
pf9MMQ6ZCHeIaXgSqssX2rnzU1K4VkHbCmAgt71H1JeMZj3xHc/slf/5IxQ6WK5p
dpjWFZUDjOfbluptx3x9+XGG1Jjk7pKi6Jum98KWBuXeDzb0Q/voYNUjfr8l29SH
LuldCrAWOnJkt9by5hvfk4PZFrH5LXf69gcehkCNWN5iU8C1r6PDy5/ORj7LI0dA
YpY8vEUeQj7ZxrPSGxN+nZBOPXuJbMYtlYtiKwM+a67EwHD7BTQh0Xwswry2Mokt
aA9pb2rl5Fo1ow/UOD6GsWooPBWHYbK8B77MVtXm9/QFy/0KAWkG94kD7avWp6mV
jtw182X8c+mQFVFadQHKvVp5MWR33c5dGS8vjlg13WYWiFEBeIQvGPq0+tfCjXKt
OcCTrFGipCjo2H97iVKmmAuzT1HX9o9WgtQCyHt95MXpMkgnjwIKmwiYRNsMPOr+
7yradn/fQWw82sQqpOYb2UtQRwG3IsPBuwxJIw0Vc88HDfV5muxrPHQIniYzGTmF
JfkOPNPruVzr7uIfeD+841mFxARIKOGb03nDKmkDXMeBeRvu1kIXmxomHh+WvDlr
c0198pv3lulrT5do5xf8kbmY8N2O3HmpsOSM8/gtU+R7Sdy+WIl4FlJiNMiWZlYG
Yq2qOXzn7cXW/V3HPCXqtGIspZls5juGVDY65FjEVv3OZG2iZeYti7jRTKZ6v8sv
+7tzeezmQealqIuXKsraNwkHRCtbLRUk8mg+BsEo4tfnWp5oW0FzW1Nx7UiuHmFK
1FQ7fBJOn1Y+KJd4hI18qKdcd/c8A1RLviq3fH1adXHlp9yq6XKkwCkLFtpYibDn
U4kCexRAQUY0VmcsLUe5Sw6MZZ8XFPIA9jkUJ3NLuKKl+JvdzXKtIFWvQRKxI0Tc
rZg7MmR3ZF3cPlKOUQq4vBnkCJQiOo4FRy+R0DEioVMYis7Lo7Eg4w3OuTAr5J4x
CW4tp7/hrWpP4OE3zKnDo9jkFMRK8TcTBdDpR0lxYEFc0ik3a8Gc889WTH6Xy66K
cxXuPypPN1tkucAa1dR65C4WUEtbo/M/X63muJNTj9lGd1jzcYlEzRp8U46Xl/Eh
53DfRteO3RDg3YggEOhbzjTyglc2OEVf0qPZclPL7a6VL4jih7TQElSsg9LrW0E7
4hOx6KOwLxvm1Nni0c5A0saPuK663kiF/51VAOZhOL0lkD7MsOUCsvHl63amGOoo
jlkqEYmY3ZDoX5vGWZBSoJA2nJXs92jbaO/N4+ErBTel4G8rLeojscn5LKuztSE0
xskOD0o5nBFDSyFM8uOYhdD6wRUhlWjLIThkJhWsr3oPIMCVlJZYVjlV+5ACJWYy
qAHZBQJ7C5IR9K24Blbd9Hayy62Nu+XgVmVirJo1NGpuBnTq9lG9UFBjwnhtq1Sl
zocid2++zZrGeHlblqs3JX6BQ3FOY/730pjHe5QUe3IRG2V4FaH0mdgSB21CKqsa
cBLoXXujcZhx1qz8cx2IXtuXmK9uSl6iau4SJSzJtVchgouzbk6M5X5GCfR2sFY3
b2pKrgM1RHzYk/QaCaZa5IHWbhws41OAzcfnDyXn46Hd5MoUK6USsgpOXmCteg1S
AaSOjfIJGzLu913Febp3SPXKPQfewsW4SEz+W9g8bMCeqP1jyBGzNMCSKC8dVqQn
go3iIoxetB/70wbbx2O79loINLR1QmzuCWpzLiKjFup+afgzGwNSRVd55KC+B5hm
5L8h6NqwydllREkcKcXcQmCTu619gM/b62Ow95invD+oO0ex4AHnG3idaBAdAEzG
hniYPcA03FVaHr98fEgiRBP/IAK+TOYWlNkNMUtYdBba+VjtdvRac2x8O0RbR1E8
oWtgBfPs1InSAxkYQvogyorE1dTP7wWV8V24l2XJC/c8KWtKRz43wviJr6Q6Zicd
YJ/x9bGOBeN5Vq2LJWigynftNrNauX1RJbv6URXEeqvcInD0QWc2epbkExPxU+w5
dsYnavXiroUHN7R85iBHcUYxe+omoBJxCdLjf9Gz0T0LmQHpyIPtgjEJtivuTOv7
aeaKPm0cNmR9y6C2gL7BcLi7qbkKK5HtMB6Pgr21UFmfRTcWtAlY3vIK0g/KYT6A
+b0+use2yn2QFi2SaEHC5/yG1SXZIOubzbhtaTtCo/JRgeM5emSzgmOftnnU0H+s
3Xmj2SAnVWIBuhERbW5ncNaqUu1lILjB3/zHMVULQ0JYo/NJEicqPpJsvAn/+6NM
Gw68bnF88JEbsh2bOmnbqSPYRdqtoSHdUAZNFY9c8bO5voNFYxEp3Ed0QHilnpSL
+sSyyOq0/Ge8W3FoVwMYDI5VQq6MvL7xbTGXMMVMhrcuLVozoH2tlt47B5CWIBlm
jkTD6sKu60sHCQeou4VHWoUzYvbkm0oDUKkAgxLLlIVSvAaIV0UR90KaHCbxpvOw
kx5twErWafEJ6pGbfwPPqbL1yLOwJtRnqtcJ9hspzRDp11Bgw11yT5Gsh3BWwrYw
IQ+ASkpmjez7Za8PCbgWIUEnzxg1/eaMDeLsA9kPsqVFcQkLemKWVDbKSqTWSTeE
hqtBURiQ0CCBs+hCVja3g/Lk8NmVUL9yFfKH8alot7Dn4CxFO8zRYc2cELiWgbXb
slqd7Z+WXluQe38qy56z+StomyKe0FrfwGLhEBj1n7HTZc59/x4ocUXx9PRwOHaW
lnQtcKn1i87mubhEPIXFBhDvuawHKz0XIdV77W19ADXlTYrc7nFlti3w3touHcvc
naFa+05ey+oe/PgsRdTCzPKBRTn2IwC/rxzYH/3tjlRs5ruAhI7FVcuQu5ESXjEU
e9LYS0g71ZCTu2xDFTmAvg59T9X15y8zZirAM5cpP6sQAlEU6WtV8FU78jU6IOw0
hPvKPBfy73AYOJYcrNu7D7uJY/DPDLew6yb4hru/CUrD0JGvkbDdFDG0a75lyoRD
LPwfF7Y8FvR7TrAzT4CfO1rZiyeL9Pb1PCtax0kp2u2o9Sqhpby7Ddl+CzgVk09I
QhzvAQbgQUv0PSLZ3avw5SlYm/SxLtoT7j/JzspxKKjdMDA87VQHXzRAZdMcIvpX
/xcSvuF+UPpl//XcRUCPwddn34iGuY6zuU/kBcUOlG7V3BpMO+/iDCmUdxlRyvyl
1gJkifcB46m3pFUelj9QyQDzjCbkgPUV8pG4lK0zc9LcQieejdFzvK0gJZFXqX+D
HsR7VByGLRObYxYHhknyR6xeSAuPpaUY0ZIRctLl0Ke49e1wjA4I9giN8QmWQxO9
odZQ3qzn2vGAHQFdvzpk0AcOYpakkjfNe2s46c9YKbnwzOXEhUowAe9haFKF1Q43
zXgkhSYVYeAe5/zvZNDT7EnDafZluGJrJYxm/WM2k/j2R4Xwwh6N/GBTZmxJ0YBi
IH7ukiZY6VGz3GJ17NlrKsC9bgwBp4E2HpIjtS5JLh1BGsvzVbdLAXiO2xOvrW+h
KHo2cALxgj01Y8iiNkU/OFCNgXatV10Ze4f2kqfXbyClugAJ8FZGhRdFsOClrbnd
voxbZTExltU50MKhCKliYhjPFKjBWKLZNUMdC7clTLZhpMuPyf6WNsYUjYEIFjpq
a9lk1HMmnfoSBAgcKJF4JCoQK8uJTqiSop/lMoJF3bAPCxtwY5PM/EkCGT4Y1NPZ
BGfIs4dIboBv26sK6hcze+50Cq/xaiE/hDcEsGKRdLRbdGqMnjPJaPnSmbOITKFF
zhKHdonJ0YWrfxYf5fFL+E8TcLeWgHyStKTpAw4Hh8kCQwgon+xACKdNoP0y+Cp0
Pqx+ts3M2lBHz2Sy0BDII3KOlnJj5wTTjri5AB0UmzRXPtQh09FT1DV0DfwHiMW4
9DEZIRi8IyRfrSPnlbRxQq8jTKd3Jr2VCjtR+KsGV28VQDvTVa2v6NmfDjhuSckP
7F1k/UINQM27c3BFxkQyhgxkvyrI5wqjnwY7+ZjJ3DYbU0LrTt6OoB/U/RLrAk44
6/xlOB0cHeTbkrUS+z6LVkM24NvGjrYke0GAbXmSpxktLCm5ajIWNQWSeU/MLYo5
/ecs1aOucdZgysEzBOt/Mb2eASFzFx3nEhHT2YwD19msW0zskv5AvbHg1r4sp6wH
ecqtclx1FtdQsd+IHc0igd72x+9GV9aOptRtLYUTEffvkf3eyG513tFoC1h1beIi
tG0XJVHf6ldJwpXKdMJOxtPNuCNYtBwvmJVwt70PqRO8t2iHV8uMAedD1evGaV0y
Dxfpl78kKwjbvCBheHJTUWBxSfesJD0URs6JR/3EsL64+YL0j6l/qlLPKLVGKcJi
GXdDHX5A451OgIYeJhBiEgxpOueQy2sPfxuRW4LcPyP0G7ioE+MLc08m+ZBEbnMy
7DNthodWlFKMwb+hx/sG1r3RK24rbJUN8CV0phaTIR2QJR+GaWZPt8ATV+3/QD9m
Shl91O0+l3tTcMFd0xfwcMSklmGjNymOJy2FfcABHQd7nT4TpmRr8GqfITDBNnfk
HERTlNJaytwt+65yP61XAF2UugLcM4l5pZJEFPrUz9YO5lG2L0tom5iuxTUBcwiY
YRlQ4BCORH8RjXWdvZo5KHzYZ2L8TnKQjMnZIkol1UZLpC4ifLW1QBiWqiCN8Vo7
px1sawb7LJOLah74rKZwj0ks670NRksnjcSOU9SMznvR/+F0W/6xE4mGbZoSCFAm
O3sTYTHjZM3RJuzTh/S2uj6JweweYGTYYws4fx+JqdAx16HPU45Ge68lLh4MwFjR
dEZyW0slALf/W38d4HkVNVaY5c3XmjO8ht0JyU8sl6f5Fpcc68QM8k9HFJKDmn1c
AUPS8Za9FsWzpAYfMovNc2XDONilXOL4JH35mezKGzqVp0cXnGeR+yopzw70kdw/
/GyY4B6nwvqJGpjRZpHSgn4VBwl0dSwC8lYKd/hUHd1aCEmSGl96fE32PJy2C7QX
OEU8JbanO8QLvsuXV2I4x3cQz8jjKG+nRSdzuWs79MbcfO4heedhMLGKU8smrEv7
jcXLxGivkzimUDNbNQI9tiHUm7cYiE/Yazwlt+rltQKyTzAmS1ZbPCMd5QwwgkiR
u62XdKFpGUPmUWTqk/k6ZOczvtTb3yzLbZJBkADlid8OMReBcLssHkSxBFnvY/W0
DvVTRPdo39pc6W3Q2pWk90DYk8qzaDbipnkyF7SncKbCNiSQd5qqhaq7QenqrJmX
No0MTHzByTdqO78JMzXAouvamr9hCQHjUWxLeiKjOE3lMlUZAP+uOKx4V/cdLR39
xKysbP3RPMrrr3xolXjks8qNvH9YjR9MaWl7cn0euTEDh9gDp9HuQDzm9So0rWef
DbCj1TylY+p929rMNGRauEnCGuvAt73pQ4xVD7BT0dZXyIjmyFNqYuFn6NDDBZh4
Izn5AuNdhKCWYD10b5QhD1vM2gjI+JRUQG4baIFhlOHmYMYGNphBQDW6LMtFtB2n
5oPx9tAVEEGHftMoP4g57vheDLjdpxL5A25Nf8k8K4D8EIzKDzDZNEDg9xAPkTSM
AP8ir9byDSYQN76NOrl4SlPjOsGOkSHP1J+pDh7ZG+O98zuUrGbS0/EetTbvvPt2
EAoDeTEz6HS+rfGspwnHn96A/URNVE+Aa9eECnn+AjtZkLuPz+AwOWxwMbkknUOQ
JSCKJJpLHMIigQLDAAMPhDmRzrE7+EH5bfTXNmNbyq+ssDPT9EN4ot7fSo4uEbNm
79aEn7bkBM4BIJpHL/K9IAjJ4EjFOmx3ErydvVXbFET9OwQ3bv3AIuxP5qnbUv6L
2m/yxoX/sm+nbb7/E3VZmXd3LGyeQc4dgMLF3iXJqiPrHC25OIns26gJD4sDR2KQ
bn80beJha0XCUvzdw1jff4bCK9aUWziEs3JaaQfSMEOFdlHEdWZmKBzn/bQniC0w
zM9MH3HBmcBtw82JD0aWveJai72Imy1s3KUPxFjxCic6xu1zFn2g7vBcN5dUf3oF
YFVZIGfbcGiGwTaTCXK67mcXyYBV/vsIJ0FvqSTZtgtyUC2NtrOD/xyx2rDE0Hcc
l/Nam08jwzFDuQ63rkPUWD3mSVRCosKT0iTJghGUm5qQHiuzS+kijtYXMSUhQn+G
XruEh+nwxTo1V7MuKgpYYsm6SaViUgnPodVyCAsdlq+srasP5odJzSEjyvLq32Uc
1QasnMu99U+PSElDDA+23IY2s7Gi6E1o52ao8D0V/S9fVDHMOAhSy3pnBWmShTjD
SmwFzREh5PbK1udQSdnM3Ozm5TuOzSJMgU9SjRlcAR85ZcqSfskklpGO+oZNQc0u
iJFy43uA1z/oW+qV8Am1H7ny05jhDlKPGy+CCIVx/DNMI4Ugghfnwqoy0hWvsUJo
C9NB+vKSu3fCIjEgGQfIp0hwM2ef2TB8iws1+oJiDCYnqAQb+EgKdO3zDQocnlYr
xo96mvG4Fh42e81xLr1zB4k0qzLGAckmG7koAQ4iZtMVCcSUcPdidZO6xmkL/rGv
iXIcoqrXTFRhuESV4buSWNSdRqzCwxe0y1dWo0YVTkyi7PPtgZH/u1PjjFetjl2o
9oGgUDeSbEJoinDz7S1XNQ53buACXPnR4aAS1Oe7wlbtvByySMMATax+svncLb0S
ISmr6fM0X+4gleS9ucZ6PhacKmB5q8M/wFLlVg97FvoT3ARRFVj2jQ0Noyah64R4
NKbmSKq/GVCNUjJ8BhBN8LvK+Dx5hb2O6LDHRvccF9kpUtnq6Y0DX+57Zo+CNlah
K2lj9Go4/CjhcCYDFmFbj3++EaH1p2CARbt2Plh8nTGEasUOxq6ktPesilRbaENJ
jKGvcomUTSoXF6XsG0ak4YVtgtiGmXM6/APM4GJyfmh8A6l1hXkjKcMAoPbsMQF+
vmuAs3cSFINILUhn6xOjWgHvyjyZauJ+xGfMxGeafOd0Z5Mop75RGUTAbq0B/3mA
4sy/9Bm1k/Mn31Fkf2IPtcQpZH53GMdeQnZ17BDPDLHPKGdmARTNX7VcWeHI7vI0
H+jg949JnUt8REL9eNR4KmHQZwFoRhS13RKey473HTHypzpgd9ssnsezZmqPAzxn
0p0DKFKLfgOEIVT2GGlAytBI6XPpwJOhArMrG43nVLNfsvWTDHHs+bWHIjfO0diI
+Zeq+u3wh9EvX8nLfdOIItUxM4yv2zgfrY2oO3PaDJVqMs5OcYwYBRrsCvozyAj3
0DnBjuJfwgJso5Mbk8JFgxJebP4K9KE1ZS1hk3V2txxNWlyRty8inj9X9vTf/z8y
O8ZDhc2Q93d35u8thDlfktgb1VNFk+dcO4uUCCSnvbwzGPs67EuYR1qMh5vBnAz4
SHZuRc2NMiooTImlNkig+eJt4b/pRLpF3lfsCgt3Zu+ed0mklyVnwiXvmAtSHn1D
WFXXYF8MY/4cd6casKpZD6QNzRsWczdq21S9o7EqnPbGBqjR2sXTKWgJKu1wYcHI
mwX/UxTMRfQ3uu9vIzOe1jAIYZtNGeky8wNly3ErTunsd7J/V4Uenxt3oioawR39
GalayPxaOBmEEzg7IAbMz8A3hxbbAc9Fi8jX5quk/C6X/iMp0faZzrDHN0+nlLii
glCWnTHcwvEPB4iKW92v7a0WCpj6hPl3g0MwFccuI2FYY0fCnorI8ZCGyyotNBTW
RuGz22/S1nCuunhv8OtUjKcmDtlFlhDHkN/fjaPj0yHl8NYuWP+AckPFdzYS7uFG
21jKOT5SDlv+Aglzvl8AekqNDfvRkER5bzwJMm1pSdhFWA36/5KEsB+K3riG4aZF
cansV/XJUEkExRgG+WH5kgwJnLSwc0X7RXOHoPbFoMA4/b705KzUhcFc0ogWTJD6
Ke0L9C3PwS7X2iX8jaVFhnCgsXOAt/T/ZUGkCa/nJQoTgUJ8oVYAzKjisbcAGdFS
WUj7J+6xIgck3XQpCyL75RiWnJvMoGqrlo0Gtdo75p+lNy/C2ND7m3HSi7L57uzg
5UtFatcRjfiVZM1r9o4L5FOTCwrvk1MRrHhY//URjLr/DrrSjDDrNkoibk3vwCtV
W71GCPkJGq1KgQTe6ktTtI60bdRX6uoa9T5ItBgPtMyt9d8gInJ1QdBVBKbfBYar
ar8s8EmimU+5FrheMWvnu1JvKlgGkA/dvKzLifU1Psc+z+yqYTaI/UMPfjdayaxX
krag5cU5EJGrloSZm9/o/pcSq05namUPz1RkOYKfm9DRcHFIwgzfFYl5D6iiL6mX
tsIfoMUY3Gvs91cDDHyNGQp6IoskokMTLZtZ8mkpf2x4D2raZXXJ7p+AK/mWoZ6Y
bk96duahY/Sb8Ge9oGRIBCXdSMgsDyBaLD/oMXXSA+79opjtA7o8HCJWQz6eZZuA
ppXenaKvw7KB4RwIB1ZKTNBLkRxRO5rWIpXudn13Mf07YPi3vUA13WVZjj7X3OfK
oPvUs2AhCSveKJPOH/cKFZ7hn/Hd1aY0Tb/MMdSaOkcsCV/w4zB4ZUQAPAmcpBbA
qmPxrd+hwXQy19eAfpoywxvjv4ow22rF6SZDegdM4kyKARLQdIV8m0JNUaj3lDkS
hJ/nlf9lqJhOBi1Wgro41DkGl34oXh6EVCV55dBaObYcTI+pQ5y3LTMWiDGZpiEC
71w+T3C02GiPs7mphNG36SKRjms4fUUQ/ezRIe/yuHaVvTeMIYGGa2rn1ptCLOd5
oDcHWXGDVhOy3AZLisXZYW7lOZceqXVXrdDIWk0cxHwo1lHWeRmuWDUdQOXRXvDi
z+cb3AC9kS1tTjk7E7TKI8xKjG4YSBWtoq72AZrwGO+PcnHqwe1fDjdq3TKFuaHq
QHfbZdZ/dyLwuUHOMtzy8sUsCI6tNCkzzNmom0bWYRx76I4ul9sX/JhOrYPyKh3+
yPfSGJLAISNfmSBln4Jsod6/iLmxepyQnygPpvUIdac1wChMKl5p3Jact3gbUqXV
oKS72QBZiNXwsA1LfB480l7CmP6CXX8hwCZbIn1sJOY+drNwrwDwU2KDra5liQsd
Phyes2bn5x6013RB0KHIi6tj2iZe+HQ1qyd2UYiFmGqU/HSlUh29FU9nolcLWDcO
rXgFLMDw57aBoV6A3cJ7VTW8FuLAxxPgE1b5+7s8MCkK/vVo20d01gjojOWmriOG
BSxfIqhRrLsvEzTMtqikOnk8aQjnWtYLNEHGF4TkFnyb9T0I9/5AUA9ddbIlwWDe
+rySd50RY+TsKUw2zP/y/2jYQjNrjWI10xlOO/T8Lom3z5AV07Dxysqt9rzVAc0w
9CuR3FW6RsK5gJJzQtBPu7mEBAsT1ukO985hTmMrJPUrpIbZJLGwBmku7EOUTzcy
QF1NFHS5CQqvqcIsbi9mzTQ1rLrW4lflgt7imWkapGfk6Q6MxZalEa3y0YW9feWM
Dw5YAoFu9kV31S3YV5Fdz0FCCVl/3fNN9jNVuRDu/knlNdQdS980X8/9QhoXoPFx
9VsHC9a7iVm5CfO7PtKBNZm/jYGObGizynr7jqTjGDxJGTFzLdVlD/1Y7UOtOhX7
9hj4M9EaZtBBC1Ubf/BSmMo9338uG9rNhErzg8rZJ+W2LKgE8jiA/wG6iFkYtf+u
n4B+OFO+gmhGm8jXJgQVXeSeGud2jQb1zvv4jsT4AUqGb7SsjtHmK/Kdf3VP/084
tQfj9LhP1Zm4XonY6h5YT1PZb+p+5I9uAqpbRrb1465mUUmMUsQfnxJ96+Bx7bJ7
w/6HC+jA4qstGvjmsm8Ef/jNjafvhSp29++/5fyZSJYIYe/l9X7hbMI40HutXYmT
f8AvGDFlJg+9u0HcqdDr0cTdiWHOVfBxMB57OEZFgohqsZvwdVHaj4Cjvl35oSif
bY0ylPyi53htS/xjALhdmTTbCIktVH68KrzbDfsl1Kau6GmiqAlOahOg8bd+jTGl
uzII/O505HJQTUyGi1Qn3uKdGNKcYak7EWWY+6biUj5aEsMkgX3u3mT/KMdj48JK
1nyafO2u3XHEcA4oa4tomBZSnQFd/q2Yhu6NBJrZKaC4us2NGHWpxTvN623QOYAY
ojVQuBNjM+q/ykUj1fsawB0yRbUW8MyC/duQPRk4SPcRRfwv8l7fopSdzf6fQDXZ
AI4q908rsAVIdZ76L99kVMmN6Z17nHYcC9JlX80xqJ6T8e9tyzb/w6HXOI/jAeJM
us2cHkJitMbmxqKaCjfdP9ww44s7guGTpdIZZA30ApMYpzKBLh67VMSm8WG42Cqe
Ec0P95oy/DTV4oGsfZvX8BAhgEuv+ZLlMXzag9mGMRmCBcKF6eP2hHYuR1+HSA2p
t1teb4DhOmtNBU76wCKr1ZaG77dVZmXlncD3fDmzw6V5kZLhcg0ou/QgMfzbdPDQ
VCxSUKLg/9mLRid1o06KIt8oJJLJ2EcOZkYQASOqRA/lD7RDUNoKYGtSHHWW2LoS
7CweEOrHUS+IhsqJLNf0yu/GDluaV77TC8//bYVqh1Kf1amVz1fEL8ELcOZ0rS/v
M0zhkZv5van7bOwG5IsL1KdsuPR+gjQO6dXOmrkLH1f4Qf3WmML/TgvixgEO+s20
/V2pTHU6r+kJHodd+tZYYQHmos9P0xs4q9iEViEJICIyc+Lq+POQZWQyrDtjtjM6
idb/44uRJ1NeTcGd63nG+6bNkoxuwCIbsZ3V910rGcGSN5GIPBzkziH+nNjKH54D
IZtAMCfZdB+/fO2PNcV6ozxfL/uXh1FBOHd9xL0299EYrvbPoaRwpne46SD/cX/1
Pdfur7wVeEqZ9esCJGJHWz//aBtI0u18NnCtywBwP6dmAX1CFquh5Je+Er+RX6Kt
OxlVaZGyTuHBP/5aSAKbr0l7cX4IRET8TmllbMoGaZJWzApdiDfBfZjIiSJMvQVS
xaQhDcB1wLxVGL75LEA3ZIJUDEAYVGSAp3YhBpvYWXab8E7R5o8TgxmxTI41pU2P
hJfovKJrnSgTIw+oTf8tIz06RTKjgSSooEa8IwCTuJzQrtv4XtUBUzp7eHF1NQkK
hRWmKnC7527oYUDQHap5ZFwhAVlsdROf1/gU7nxvBMqP9ZZQOjj2pvkh529Q/l0e
QAcmM/2/wUB3FzIFrW+LIUS79YcYVfPibNn2oDRTmOmAzCr4RXuPdaJt3akqKmLJ
9+YkTVPsb9+X1rk4WQUYJEsa0mrdPornhJ+2pIJRM0O7dR/BtALETZpoAQVDGQvv
7pP093G/uwd9btsrv7OBQ9TV82zC0tQ2k7LSzzVkM7Iw3k4lYYzgd9KwUyn3nSav
KMsWpUvJN/kClVrGo4kIuFbk+k0ErsoDAlpeNQ8ZNX2/Y41cnA+rhuDQcFUDmrH/
zh9GaVsqk1SZgeJfpGHUJ5OU5sIuzRyrhxhwqB/6wwxPFdgZHTUqX4aV1le9+dvb
7jZkvJMAWMlXouIkG4rjvHUCP6q8fFfO2UmEyJwOhNHk9N6opd1aRmih3yfQpody
pbRzhsh/S/n5b+jetSFgmCkiBhwmMwi5MCrrLjiFbxEiadQr2VmfGef/PuaYG7AO
XNHPoPpufeoIcT6wTtkOsrbVYrrOGrfPzn3pzMx50EvZ0BGqbhoN/GloQCH586hU
ocVBTORAN3q8D1XqjnhjuU7Kx20eaPXhVUQtzufBrjb2jNcdwmO4TmC4fEteV0Sp
tTeiak5FifPUDZSU00pgJTZuv1M1mS0ZBUvgvCLOYzzgpJe6RBX7ER9cz8b9JfT3
UDQ8P8L+VGJORhkrwamojICi6J2ryP1xBpuEmO7Kv0LjHeqewI2LiKvqHNEpFXkI
4HciY81P/J4bOaDZrzHLHG1ERINBzOy8SAOlOCmyxf7wjPp5k1tTBUvudekldR2k
17oXDi4gaWOu2i8+KIo2MiodTEaGjI9S6aM2fYKopEWEIDvp1zhFhgwhoXnn5nzg
ElfIVT7DdvOhDPlT9I4/qDatb2IOO7uNxbOt+DHIFUGe92KO5bW90mSzqxLFTBeB
5ka3QzMxAyJOg5aRbsUHXT7I0jmLelZtkajsr+wFC9q/l8DlkDmuWRs7DqHzmdBQ
RH8rdwKNVyQJ+6NV9J2H0UcNwKM5QDus7peRK/HoaXt5+l37I9Zci1nP9FCNcus+
6TuC1oADcgFA5f2/Z7eMa7oWySl0kk8/9MXJHUDGt9/mdwUGEYSBwkbFFabI0Tpl
HB+w2V5RzCh/1ycdWlwxY9PKtNOrj/od8Yw9GqTdYuAQC/LTo+zDjfbKETQK+WCk
ExuRSMYGXbJKgUo6DikMiTX+Nh9UaMdJHtwg5nGtFsQpEqdFePUCjvM1UIQSPC+s
zZNrJOJmJ/+YDIzcmxsirMX5+6m/qngz0wr+NQV8xxNRP/RhM9pAhsAA6lleVd4D
FO2pFXRGwcGpRZqNJ2YxbrJLcNQ7nAXuj8clIoUK3vKQYtWJZ65sntcdGiBqv2vu
hHTHbf3jBA8MOs5U10a2HB/2BRcJzBu5rfV6iAyZmT21DdUw7CAfobG0lnfKYgVG
juC8qGBusQIkI1OQhzf2rHsD/bJwQ2gxU7oGPGyDAMghF6Jp9Z1XCNpUmL30guQ7
azvsPu7l9IEvCowG2XHmMx5aCqvjyWFDEYZGulYQ3EMCWzCvHjt7Bq9Su8xq/5Z1
j/jmXso7TbAfJZC3mAyUMzB+ZtCY8qJN5fCrR9uaieck4K10R7wBvrs9ZC6HPGzp
seMfxGCP9Q9IDaggwfBluaMiC3vMFcKePU0iFBOIut7fJcHt1RXH/2RM7IfRtMQV
JVMILoFdCmuaMPSte0/BxNkXo/PtKv25qxSFML3z75bMcLzp4RPsSgaD8ehjmYtx
ytDlSuecZ0a2DfiLjc0l9yyRzH7+YOxb6Sksafyw7hJ2BTp425O9J3AO9j0r/6Qo
c860dO9sMc0jdguM3+e/ahBtShsSczJcDJzwqfC0WQG4AT9Z693xCHNlfOTphszI
7ihKpwhWP6eoj5Gxsb/kAlBQWt06f74f4iSExCYbJ6vmnIfMcFThDDzL4G3N2pjK
tjHp0l5wCzWIwmt2v5WptljdeZQL+zZSvsewefeSX0B77DtEUtklRvbTMqoPm5/6
E2nW3KbLNWADRPeVvWj8ccl6YiNPWcSTMbC8gkbrKNAzaADPeFRXbiRxkyMVXG/F
WFND5RNHjZTDfchNAfsltjnpcjvB7uTHwYTt4XSJsYfIEyiRVb13+1jfeOy7RpfY
YYR3aQtOJlMV45n9kEn2yh1sIWx1scwU5iIh+oLaqe3/6WoC4SEBOVkOEjLDxEPA
0GPpnDi6koXCorhpiOCnUZ9QZxR+UtGgM55/VzX7UuliYw37bHl4w8ab2calWdWv
9ojGf+8UgHjTR81d5V/3mC8tWVCQY3rw+ryrpYb3QzNx1wM0SBvd7JiZfHcL2pjD
RhNRaA3Y5b63sD3NmjlzOPRYLw+vMAG/VsRHhQNUnmns9yW70eOT+2VOJcjvtAj7
98GGKy6i25Cv06g0L1yl6CJcAxqhIOAelOY6ot4JGwUXbeuODzBydUTVMb4qoGkO
29v9HmCXmOFxA4Jl7s5CS9lekfn8FAKRUsRViUxt8o7hdSgVSB6bT87F0+Lc56h8
tVi7Fiw26MudmWIg/KNO+WusHenGoPlWIQJn58ck67IXi45ORAFqKG7xjmTz6B09
qj1Tlp8mluwnJhRYi4IT84FqgyBycoN44RkrSwoMtfCd0nYx4WYMp31G8HR0lmxs
SIcRWg5ky1rZsDvhxSolBJbbbuh50hBeuHRAEJmjlnPxemcmz/dGq7QqcOmGfrld
XE3fM2uRMJr1jXjfL00MsNH4Yq4KccrsDAojXGPE8Rw88iV7OShSh9NkVWszRpw8
zyB6xxTRrq+C2BKtFAp+k2D6/WaPMz1ZxG1Qarj/bESQOk2G31/Hz5071L/3ddgT
LPMgFApnb6SARbfdcD8bDcJF/KTsFvDamwxWTZYToPx1ePKc8sm265l1jd4edy+f
Pwd1bIAZCOaQ1scL9Dd/pe6GyqQoLLJ1GwPyEAmhkB3Wh23PfCAjHNwxqW98gv/i
B1jkWCDbi8AnJWRyOO7LM0OqShYCKTOquclOrhOAk0c7YXvsopOGBnLaUXdbhsq5
Rx1QRjWndG5Z6BGdGw13Gn6zyk26dwL9I45cB/5re0YzPqiMJnKFBcJ7kI6NFUfI
Fp0Te4tTwOLA5jW5Ft/on7nXkbcsOiJPPuDKCgovJlV+twFW5v28yuYYN8SLVhmg
Q3dbuZ8plwQc1FqxHZ5+P16WQx9tnvj4LinLxlOZACM3M0skJ6eezFDRDLJuSATq
+tOC/mzy1fosCxb9VdeAOZA7Ey4ajSAz/qZqFUhe3XpALv2edsnUmNP3QxjvmW15
Uz2sCukZCUVK4fb85pvzoUGeA0uvpFZiYT5y8MU/z+8IlIetIi/pYgMrL++/AqlL
ryW0duGi9w87LJrrvYZj4MfZW3FVuf5OSV38QW2HAODjJDn+wgxLELIZNxSjcnCL
QJMppQtVAM62YyGrKtHyMIddwXyFu/ikkuLnHac4o95dpIioqGHofDrl7cnprtSu
iCnJKCxLP4wkb7e61mQpsnJCA+gyzDJwVN5De2KHteDyAQOgGpeELd5T3oIRCx/I
RisDgmyq0AHmBxbBK3FoAxfhuCmxPxZPbmgqFBRpevhKusZ6j7w65LBTY2kXdqQX
WXkvsvh4lqu3KLSwxvcCoCSrpOdzbdnuz+j4Bm9emGW84a+hW/j/VfKji16POOFQ
xMzWQhrpoWp66UH8yFmoYxQYZhoxKFcV5+8SiJYPWEPuuDyABLuGcRJsKKI82zOY
prL1oTmlKTTPHdB+qNCASTYPTK8Lcj4JtOm+CjcdadEYTCPRmEykvJWGXZtb6bf7
u2EDLhaXlNlBtSZeQXFP2JRFoS1lW/pPzhOhzql712fIFwtqVmvQNllqKj6Lw4g/
Rl+mHnUTeF+lxA+OpcP3BQ0Ma5qZtz/gkEW22mguJ+IlwPC9TfKgEeHTs7UbI1Qh
P4n+8CXWw8hzDULxj2Yt97LrcigG5WvDIOJiSuC3E5qjYL0KAc+Os06itGEWQFcs
zDIWCCUoZZ3P8yO6Z6oDHnGqlrjMx9W7AlmtPuok8RWRYXZGrYYoz2ooyvkRY0E+
kIiMXAqT9f7yfS1IPzuv5OkO0TdCcm3ffzmIH1LAmU6AsYEbHs2Qklt9CLQ4SwNO
20JTpYH5onASVGEsjbySUryUCi6T1nWl+I8cVS9/1xt9cuW5jQVYIMJ4mVpYhRF3
WAZxUYXeCGa7hJXZSXJwg5gtJrxZaTTZ9E6kftAYPjeCUE2cUJZc9dTREq/Cq8X9
mbDFfkLzXOYEKwbiHhVkEzx7WdwurEf/wZ6mauzf6fCYcVRcNklx93DiPbt8FXjD
HWOGxtLJq7FxUucl3Cwl02C2ohmFbGLtF+HWsO3rTTMDAEhrB2zBIgsuzBzDxyDW
XpNhG0nCOeJ/FXfX4QnPU/23KGt8b9J1Mpx32Ll94ZhAUZrbhH6XMz9B088Y+8g1
F+iQ1B896dwTXdm9HXYJ9dqTAOd0kDzx2MEK5aOPySDZfCPXDMUFaoRRAyTDAXah
/YaA1fmKXLTmO4qJKgKa5iHPD/ME1LoFehcEPtIU66M5op/eM05xWOWbFVmqC+kK
fqTyS1m+8m0/iBGPkvAl2w9j3W5IQN7es5+q2yRuSvw/uUSdiTmZPQyQj/qzTnrZ
1fCMF5s9IE1y2T9CyrhWoNmpHrFmk303Goj+X469RrZ/ql3wgv0nBj+Z5jlBPkdN
+DfliMGBRlGJMiJq6Lr479B+vVw6dgIZWQ9XORoI7dWshYf3HDeedrYQBDkdHT9f
HX6siKsmLyLl9to5gA2kK7f7wnm/KNoT1Ia1+EgxpcXFnrH6JisYRFD1B4hePkMB
sir6Ihsz1Blfe+wqouX1HRcF2MsYwjhZ5XUVv1I9DxZtSals2xcArfCjht4cRJzS
qCtq6abolFlb/YaeAt7iVU8+OUnWZlf//zWypAaDxsPHmt3usqzdnlsVec674HhA
Jbk343rXrQyaMTVkpBAdRZ7uNky7DPByjEPl5Vu3F7ZO+QMp3lGaleVuKl9l7ucV
2JXWtjSlzVH+l22CN105VwMMnYISBZw8fuhY6oyyk4nzkzJ+1fz1OE4zsOwsC31R
4Il7MENxaFF9juyzU/YT30GzziZuznNcRK1J8fFIbnFv+JNYjLaqTDXZLr9Ez50+
VY1nVp94i+8EpWCOIop3/2l7izXgzMHez6KV3h9WeG+lLraihPajG5QxGLs4VBJb
TSH8ezIXB6r5hwekYlBy8gMidReC+b1bfEp/2r0yXjAkCabqdnLrRz9NtTHC8ubV
Z3h7vn0PwuNW0GWyQ++oth4gStfISfDYReZGZEx0DrGLe/3x34EvWi5+Aaw/Ekp4
v7ZTJPx1gQZSQaeJarEtTg6A1xlGIPVfzuLXFACp3G2HX0BhT2L7L1139tWhVcEv
+P8Mhxkai1DK6aJ4txO3cGq24/iq9OVsLuTLLWjZ12fJFhaUcHf6K3WXDg7bKoer
0NNV5JxqUTRaBt+VBpYDIuLjMiwVQnuyVmv0xmTioY+mVyKhO4KbImbq+VnVs9Ac
occxAuedzH1klweGGb/JT7yOLJM2nytKP/aXng1aV8CPajeX/HjBoSW88oB+iE6e
bjS9CIvKu620TMSkuYQuLSzelhMY8IuTIEgrQSV5OvJhYRoHirBpj42uGV4HSOGl
Ozra6qv5L9bwYY2LrSdWoVZEtaaxUUtu75gHoKjzXGhhezazUcPf9rOnoAH+1Gee
rWL+xP2peC+iRf1uOb5cWiTs31AdDWzCqL9cZ9UDYcZY6PyvzGbJGZFTE+B/b135
Wxnmrl56fzjy/2D90iBd/XcYip/JmkOcdyONTpzpG4Yj4mZ1wLKMOHRwYJUN1ja4
owCr6KWhGczsaDCrDJmuvHrEEXgh7g2Sglm9nBA2gn/uswAgcx1qp4Qwvb8c7nag
Ac4UM94AiLKn0uz+1kk75UNXy/egDzBHgp6UfRJPPgaz0iJE4vcXf/C23w31VlRy
giupf0TiVhDzzsx11x9ljMx9DEnjTlaGmfZYHrIH+36TorNrodToodpmQ85I4W8l
00/PwgAToqVgSh8RgTs31xPFrHIkxVKV2N/MHC89hgf9s5sUmZRj7vGkHR8lAut5
VT8EiNgpsqBooDMqSOfNFSIsWEXQho7Y6kg6xtMmKR3+m7yN7n0Tr6QXQlsR873N
pARuVNjxfJxokIFiZU7qLtOkg8tNRymj4UJZGZaeuugTNBjZJhHUoLZAj/yFGJtb
CPs0nV9Ey5nCh1VGmeoOqeyJRdpnP9vKO3paHG8AXYTU9xMAdomvhZKOdWU7eNlD
2HKhGWcWlPuVUSmozMMHbP906uEiYMopuFFixnAV+ydR/v98BwNty9piOq2tFN44
ra0vPOnUNV5H5kfl9GQAqwPSnElzmzz9ERv2Vzg5H8ViedFaCc1sbV2BXJo0V52p
QG/xTFHKEiz8mJOkkf80SEFPlERnjFBekUR/uOWsbP4cuRBqy1V8kR18vOwoUjKh
KolnZmvDVgzwvBvn9aB8/Is8Y3L0dWHs2M98y57MffqmysdeOiG1pO8s/VL3BXKe
1tDQ/W0eNCkdgvFN/fPJed2Mz17Gja3gRmsqSZl/H3zK3tqCjzXTd358vRfxW/0Q
ZrGggKDM8QRBrHB3legpL+2dep7DGeAdus1JtWvfqfTk09t/mPbeulUr7MLP+oUN
Z1mdr4D4+XNHOCVbhm7RNcr0cv12vB3K+LP9ekNDS7MsNeH183STusIpiHCGIAsI
rXFqHzpiHTgYwNz/hGz5TvkKf8OICLI86BrAwY465xN1b1X4QOFIygkLARj26rAj
YJC6qBda4j84P3HTCtKoasStUafLWacLqhBLIRgUSwq//XzwC75cBQ5qsksL9wkr
ViBisAd5w06LVDafZIaaLT1UMomrOh/cfHAGMV8iwZW9FhFylLVchNiLdzKDVkcg
5V0cSL4ITtd4kSRkkqRRQ4zdhl2nobhQxKY3wlcoHoiTljJX3BJnhTZX2lwLX2wp
pgeqegeMLqPG/WL72vehylLlrXeRoM+E1fibalXtEqLIwzyXc/EbVtYTXHEzFPwr
LD/H4k8so31TJT4x4GgpNAVWCHqUJU+kyfcWxoIS6jzNyCU8YOGh9O+DengU/B+K
dwsURQ1EDPAj5J0ffVOtcrbGxOXZ44wyb00dJu4asybDjISIiHjxW8SbtNNwcH76
YgF/pgZuXaQGKbS6zL5Sij6jDXjFsFCiaQqnAeiNMgLllPkyQTUkcobeYqIN9Osu
f8/ZuzstS/BDkdHHgCKSQSFx/TAOkoEQy3IGEg1eMblCt2PCs4WCDylvkVRhst1f
GdqkZWHQgHbn2ZoEReV2QxXjUC4uQ9LSiyDQElZNoWGTZMnzt+EbdnH/MCNKEzCM
iI5HUMI4YRCSW3EbqVWxu0CF5MeOIauw2EPIKITko/raMvQrGCSbYomxUiLbJrWl
PxPeqHsOPjh1f8eeA/FzwlkPo4BMZ/bSkuL/sMqBOueyb02PMNrSMG+zTRYAHaDf
e9xQYjqd1KhCiWWW5AMnltebDWvIZLER5GEvPCgNCkgpIIP0Hjyy7/dy+vm2Mnc5
u6CAxRcO4RNZxMQa8PsICUNys2BFFGmUDdTS+FX44Zn+Pc5nmMykcp2qtb6dRJEw
Da6p2eYvC9apTDRPd3iCRVgN6V8kBDX6tJsIQ6eA34oQ1o0XC+gSFCmwmbWSezYF
vLZTNy6Jnbg/n82A86Y462n0QHQYffW8wTtUmkoBvQTUrkI2MDFrK3mR8e5UJPEw
znfHS6yGJuogc/rZ9fBwizIM0cqKfXfK4G0CBDN4P2iKMGBsuPkBI9CN8kmclO0O
etMu9rOCaZeT749YGgGsQ/kPOKhww96ZqQyJ2zM4QkhwvhQxTsV107v/9LoLb/OP
GTIEj4+pDhkM+42430RIx6lEEk/qVVgAhXstL5m0VtJg00AtNUKbO1D+qVRWFYYr
XiI+AGGbf8XPQO9SGeqoOCQ59m64MRMS4Iuj5XVOkFJ7tTccbJM8kqXe+kUH+GAZ
X4qIFSSpSOdvnTBPWTh3lj/ptq8TkXA6LCntmhE82dPVXMmGWWl+gKXEWGpuQbOC
R8yi1ox6eiU7b/0nlHZBEBQef+W6RciJxf8nTVXYv0AVVIb8EOE3FaVQwC8D6xRH
7CCvlf+FdQW4AcHN2BCAmYWnolpUsDuMQGe1AgqyATRv9vuHoPbOpNlNGsZe/3P+
zv2vKQDIA57CAMEYt8Bf6xLsSR8lLSZVuu6IplqpWOLH/jRzLOzfRFQfijuKPXs3
0H5jrAIvD2OKNb0RhG7MLxSa+EgKgjkoWeGA7uUICjzNXsPyLalMuhwAbL3KjEYB
/2XUWH69wFp66TYr4IwwzxWf2xiq3Zdmtp2Ex9a7y0xM54OZMdG+jtdlYgsf1Mse
fkFZs4W+mFfC838wNlsLlp0uINrxljfMXE/JDx99yBWByY/cG9d7KqEqkwajegIa
zAFJDDdP3e/ywsiWiZpZBsrMhLIFcQ3nRnnvdg8VM3wsnBW+yts+eaPAd1cHdmeu
LTpfc7Ros8kwVlFJzxviwFnOMJaIIjMRGAt+kFnzSDSopheeWnGgEHwaspyupqZb
n71QVNIAreFQcxdZXo923LBxy90hrXPoqTY7yrPsyEYPOETcXyli9Pvy/JmUH38I
pZXTDq4LfNtQUrduw6WmmyTQHnapRMUo5VreJXITg4QctKGx2PNTrdxGQgWMnAeI
CYx5fQBkEZkFqUn7121RNSfZfhD4YQSt0llC4mevQrXmU7mn9e/bT1OBoR7xC7vI
V8qarTro0k7W9MY8MHUNsSs2+/4iRGGLsW/XtWNsYs+nd2xIlOQnY7P5R+Vhl/ac
si/MXhTQntcDbF/mmz2jzzjdZucnuCdogFB6N0+EcVFne1ocT79+D2HcebV3HpKE
AKGfw8bubAi1T9XhSjSdGwlDF9HXWWcIs8HVGeadSisgR+IFssfUGjjZjPXj27rr
zW8N/e+Kc/RE4NFmFUaJUby4HTCLEmIHaZK5qDHavO9d7WF8wCKXO29PxwIsW2rB
nkQPbjEYAscf1Q5/zjCvr3O0YZNzV7mujRvHGg77Cf3HR0GNQkLpxfakfWh80SF8
1kYgxrTS5jbNnRbJoDbeEiMBVNPJNAKPG4p2x4kkA1e7qeFMV56NpkpLRFDaPARg
esazrGKT5l/YcFIX8h9AmbZKfA09iC/a1reGePKlJ1B2BJuikFBqfDiFSvpqsj5l
pDdvCWznS+awhLvX7ZQa5fEcENPB2HHS+tSuZUt4SY2YP20R0HkTaAWCW4BR92Ht
8+VFwmpgsFw8vOe5sjlNf51RnVuPb9mYM19q87v1bmdAWOWmrEYrtRhAyhRRdKii
LsWrSYZvEZrPzJfw6GDQTJE5+cJPipoSCc0LQPmWJTX3tEp8/YwDyX8s08UoebaG
BU0hRwBkJ18zm90zuzof3ZfRDJ3bZf6NT0rBtXVaAHFhFPxy0nhNNKCjAAfM9YYI
WBK7cV1zCby54fDOYwBmQFhJB0HyWjlm7p0RbEEyJV1N/BJFBR1iL5Yxv5OC55ck
7GJ3mZfM3Tu4/dBUVUIqQ0Su0Dd4BS5bj8WtQky9PSPTypGWcTSNmWjCcYwvRGiK
DUy5XsOBRnTWZmEbaWKkcZopJhnhLjztGNA/37RcX7+X15BpQnHqMptEjMiCSAc6
BdYSrwV0ao4k8R0HJ86J298V8bCad1qfie4PLQvSXHl5bhV6+kcvUd8y0Fc13Uj0
kM37wRFQ6aGCKmrymzy1nXj7tESksDEKmuml5BOQL2PqMMay4R46EQD+vv9aS8Lb
+s5EPQTgtHH3jJjoL7v+q3Mxf6UhpXMwNVUc9477rpSHYUmI7YkRZCt7bUbljSVj
P4T2gCmroubXXuEqSpGqFUpngPiRRKd/i3HZXFl73VcCoZmmW1fwwaqdvjFi+J24
RtaGJoz9H037b3ZFtnOc/DQ1qsUP27Lof5ISDVJCi+iTX5kEFTSQvrS6z02oZ1fp
IaY5hw3NQxBDW2cGNSep8K/Rrm+ggNsWebEiPouDKDtzLK5NsDl45gswJqPsA02W
N3nL90igKRSBcHzpDbuCRZ1p0sfLQXpSqOh0SDMuXvMut0e8EwstvK3wjRz5zTvE
rkTN80o7yVNCSvKTxwfIgyJMfHQRcb92ku8Y7tmmI+IeO0afnuLGFYhFfWtxcVTL
QlrNHp4WT1zcFgKpcjpUIkqTLHdXz+wC7PFz/JrgUiFlUqqozQsYR0HFiciRwkPC
RIh3jjOQ3ywLe2wN69k11M/koXadVcvqZJ8cQrtqLGFBxikxA5ymS7qj0rmqvO0T
xkpogy/FroTefuLkZyGQnGrGMnU0DRoKuhdRZZPokJfU1PoO18jsYlZcA5tw9g3J
rbUUOnKBGRl+6v379PdBinnWsOAhndzDOGBDNTWDtjc8O1Du3GyPcIuTcEjjWZIn
YZy7F1DcroIEQr8iHN8WNAMFaFCUetKvipFcdCM9gCjA9MaSfREoAqHdpn+HUK/u
BrALnBaMw7qBQXGtemb6RH81LywIGtJ6zMcBkoVFefDzQQRaYg/FR+OjaUOcADiV
yvBDoLGNnNILnoOL7gCXcp8oB5kDWOBLZk+eR+95wLKLcTYce8Eglmh0xEd6cTVZ
XIqzoxOMwtvGHXTdusQ5xuD0UFzE+CgdwqKrGTOFoBV8J7ozK/KWkAT7xExnitEz
0qKp9irPoYDqsWG7+KtIXDVWlo8DLgPeR/wS6PaVC5A5AiWCPInPzV0mEgJwClEc
wMVqLsIgHMzHOeSWy6GJlInysxI6sRETElcmgJkQEXrg7IOARWYikk2wMQVUd4HN
mPqPTqQLSS8pp9BTmP1UlmOC28wBmpVLZPIzoZIuWYwmDnaDfzXlzVqMKSbrNAoa
fAwGDvnm9WxnETSGJ9llh3ktCkbuUvXf7IJZ10TWkFFLx96OQEXfw10f/k40qvx0
0YbofQ1qENKbK5oAqGDOzli1io/pxVRsimdqEqFke6woGawhhB5gYhgWZiUwhTsj
evhH7Km42HpLd6dWvrE6KO05mwqvUmEm1GiEpakFGeNWYmKeiVSQT+D/dPCN5bMq
9AwJLKwhWMuE2DXQ9KunevGvZHy8B9jrb1UFIyHpi2M+yrN5XY+et+EJEpXg5GBF
n/j1B2DVNWARDurxNobSenDJ3YeaD1TgXZQg1tATcO3/irOGor99btuuwzbOaTSu
Bi4ywO7cy2i9cNZxKyfpV7A7G4B2XYaJu4BQgoDsbGFuSAxTO8OCK0kUHGmKuQhw
yZQFRSEbqCi5j8IbWLo6wAV7/Eqog4ys5iUuDHlihBlntHm4XiFlDlrnWZSPnFqm
AgWGyhi78diElyOsGTkxhwzBTQ5BpiCsY/8/ClSepiscYrbwoEx4KsHtOPSJb8oY
jzVU3JlnFmaMiV3uGWd3o4PekWHD+J0/R9jNPqgb33v8XvWsbsmKWRhETCGzFZBY
D02icctGd5DL9wZeI2GNcgF6vftOGQBLW99iY6Xu32li6abifAA066hm/K1+lQQE
ZP086+Wz0M3hb2l/iXY5q+52tSbJchgjErMetunqPL1yEDkRKiNKcAsS0zBQxXAU
yShy6/U27rNpNubxCUopgGPb0r1QV8wJP26/9fzpsPEg0sZo3GbJAmT35s1MVHMc
rF4jKBV16nQ61slOsPQKzGCJEO/MbyJNvPjM3Gm+RUkxuYjw1FYW0sJnvFS1JoEP
Wf/qZlDp4knsxm6/VE9YlYGNFljf+HakPj45pY72UudvWAUCWi/hVtOXdDmP/iL1
joboFKXDIgufli3NL9d6eovicVojWUkqgKBaXeO6CRMSFygze7msmV/VvZ61JKhZ
uAKv6iDKvR2PQiv8ToNeRyPvEQqfiWIvN7VZaEbhrSxrQ0Gh3hBn/DcOJvBFCy5J
bdyLnI6hTLXWBK+UrnTmNVMWJoAOgMwtk+ov7GBeMeaM8HQE/S9r2FhzW82133F9
veV5yT3LaAXx8FAEDYbnC61cK5cjX8rzPc/opS2RX8v9HjKuk049nluc+nFVBWMm
WSkdcYbIj0X5qcVQnkG4NBIfaLBXtRddH9sFZ7p43fyA5/VuCnw2CIq+oC8AFlZ7
UIVpEIZfLWl9eiEFI1nrAYn7UPkejxTgYtKjaq7nZo9IhS/A+WgO01WjGkeQD9RX
7nF98MsbNqRAW04xhyHrLAVZGe5My3UwUAHR7h2Q9D48easvzNBmsi+01xYTtZwv
8b70TSU2fqZlaUSbj4Uw5JVsJJW+qgqz8gThL0oP8O3Wopirsvh9m20XnFKRbugz
3PehrDhn/rWxoazLGTeMWMldzPGEWbVSj80tmm7Her9XpCY8qSJXH4DAGMgpg6OD
h1CW/Th9tba/rTSBpSXHR5gCJvFm2OMBMnWn+UJI6IwP/O5fZOXGHb08C3XFJXKc
CG7byTb0sF1PHnQShomeuM7wo0uzPLG3vaDRIUb2hOCej/IyrpFbCAXOhu2yjlQj
+/gzO0BsTWDnKTxh0OnRiMVUEGE5dnMhCArAsf7Q0okzFckLiLlSrAI+gIwE4EiJ
zMlRLIYkN0V8O1DxA/3gtSWnUJ9y5x9JpCqkOGeYQvEEkmigG6bqewPupkKsuEOR
AEd4ESxacNA2qIhuejV7TtyxJu1ADJwAppzIxemIYqdjuvhbM2Q+Wfy1EKlsgS3F
2US0/an0lW3CxKf/UoUn2cks/A7JSno43Nt6jzN31A5bQRK+xHuV0v35MStiLskW
Xig4kQuBbJJjmuE/OvQhhg0bOxsH6rzPIMFv82HwsW/4RIxULMm7rV+JZ2n4XeCb
97/Qc53NORjV8E0jvAIB3P5avWleGMw6DT6qW9PHS9Y6OTELdBAdjYy0cgngV5Ls
a3s42Kn1k9fhbpyAXZa6jO34YxVPhxzJZubPGK6u5Uv+fkQAGZorEkykPbaa8khS
4JlDakcX6MSKnZLVLV0meQFcjsdC7BwIgna0HJDRdfAzePP8Slt2O3FivDkYv7wH
EDl/pxDjWYrzU8BFA0uip3CHumMUAY1QGHPb0B1u+FFZLK5vSgXx/KqIOWvtm2tz
/TxA61NHKEw0C+6nmdKN71ANFTaJQlBejh29e8qfM3UftXO2R0WMNHdwrUA/BtJe
darCRwlCFNQYjPYu/O9CeDYCyeRrCOdMUE5K/RuQ4IANL12o7n8MH3ffXzmUuCLc
7m0k6yC9y4G74Lc8sviBn8LJEqVX9qTj6VEgRnL9dB4/FjsRuy083z3WEl5vEXrQ
0XOOv7Z6aoovKm5sFf/khCEjk1ogBtQQRnhPWdBF67S2gbfe+jEadsFG6lFilm3h
lzUTTSozL9GVc9YuUW/irNj1wJ+n+bvgNbCnD2a+4Xfqrz6xGpPjOJVec61hidV3
7dktrMj3czVo2H9AS4fkT+PaLy70kPtk9goNPLxxteS6YOaBByFV+AIt8Wr0/m+l
rc3P2ekqgK2pY6TyUdtb6SsgxjTpa8WICWmzlvL+djp78VATvooG2YsjR5luNJ/4
pvJUU93hQZwXJB0SvKNyLIjQbeMTR6cvu836VWFOtSa4StvSjJtRejSGI52yYtUe
vC64u1CGk8ip+0oSNe/xCmMHWkkiOJyYmaFUXrahqwJIrMpHa3LQCDLkt6ViFdIY
Ymhoy0NSjAioHUwOLuh7fHYFlcykcOKnlhz1G0IgvSd/3VHBQoCVimYX+sP8GewP
BaMZBzS6DEuQhx55WQzKLDZFxLdzScyTUbd0XPr3tWmfsNSHXFMOXr6593HbPVi0
hg7GJsxgSGHNvSqqeiV82DMIxB/uhLjunXl6kSlBxwgSIOcdgA3oXrsc95sJX7SX
vORqQPBRm7G9wvFG8ZQAGSypcxdYHlWT/24+yIH48ikJuBrgulkhfeJJwR/f2FlZ
Cxm0Fb2FaETOACqqMYhe5Hnlg4hmIzKqWU7ZX0D9q9Qo9TbF74pUZVIMzs+aDIt6
bhObpXYfEgl4GDJtdITpIgIqzx8qZHqI2Zfg0irZM04Aus9csDaJGzffNi+29nGQ
cGE7lRUuQdZi5yuvwQCl+ykmGftzOvUeHeaU0fYfQrV1vyulYJMd3I/hCxd+5aHo
seyDxXQH+okzV4qRVuyk1Hg9j7EoBbkT+rk3qgNpEjax4p3Kc6h7WyeVxhJdSgY+
xBLDI1aCrE5RxyhbXkDC/P6lCQsbESYEC6SguhMhpQyz5Um4llEVyv9gfgBvoC4V
qUo1oxR2PxJWRmEp9AR3P91FdvFgQQwINabdf4NDf9HCG9JdMzfhFmgVlwi7OhW/
/iLZQssSrdQs0J1UQ288Y3RbOjLT+VbQqcuj8sKrFZkH+Ns0z6065CU2fhvwjevg
XSGhoz7jtFiNjXcZoLtfGzt+AYEmAEmtHV4vPf7e7GzZdrY/ScxHAAUibWKJv527
ZDhOHZ/yKYhfP/jmvAFmq6C6JHWNe2kkH6isd7kHDXIuehKI9eXOOHsG+RNy+OW+
okuXBL/glcNhJZDYT1o7AwmUpCvlXfmJMF/f9FCKEjP5zyCCBmmLmB+WHNc223Hy
569D8DS83+oQGc9L93i9OF0vUN2OhjUNDQfPMwNiuBpn34syB7aYfLqsjiuuVNrB
oRdQBE/cSjC7wa2xBPXCnX864egSXAvjutA2iEkvo07tw8XbOcHw9hLGw8V/ZJ8x
GunMCBfKzKB4WffNKWgINbK9dKj0nF7+uESlgRmoqvJqQd0vQzsd3EvYHqTIIpLO
bix2CGzJFX5rYAHKsqsLC26qKHYef5+nSnooOqAF57ayAaFqbrSWJs076XHHim2U
xaimB6Br4H5FsGXTdAy45uTW2SsU9Kp+DLr8Zhi+yUssGCLKOhUxGpcbf5S0UeBY
KGOZRdRWpqsgBUuCk7i7RDn8No46IeVC7mgLza6YJxDeCgxU7uVTemR8FqeRDH0m
XfzYlvuoQU882FdQWZ902KiSkA9WQYGX1IxtAiWlmS9alX96cV1n7SzSXmakqA/m
zTyrPn7V/iTmD4nHnpEulltGS3Ez0Ifa3+XdxCouDNIHzApT9kvczo49UCNBN5kk
C52m0wm/myGBT+2NPFoNSdDReIoUE3BVwZvD5Ys2xlHvv8w0kmvogIZdrhMUi4gP
Mzs0bsruEBYb0sUBG4GY30ooDm4KIxZNSlXcLzQ1CiqpF9UQFOIjkQy4iwNYDC7Y
b5WNRwLKir4j3fhoa03J4LDL6XtdX04eh5Zheszp+i4Vta6N6DfmG5IEhWDnpZd5
BJZqeUvjcIDRi5t64z/bjE2sfReL9FybBnanDasOqkmKTmYAVFZ65vk430UsXIYn
w67+3IIS0kvqFoiDGO7OBmL6GjHMWmswFp9qibty/I6g7m85eTHaqnfBiBd6SWBZ
LvJbzTBa4hHWuZ+yTEdiF/8hYc4SfS8huWDzdByB0s+Q5DQLBSrLofR04gimDqhd
IaAsvVuF6B/Rz6JIzsnsagvl2uLeLI08glQ7RZdKxWwNX+f6c2clfVE+0kMSKzN7
2i8FOY20RC1sCG8ie1K7B08kcyVYFDGOSjXTyOoba5AHO8oqVfpatReXbnGAB5ID
Dlo8ImmmQKaF1erkt8xvkeGJS/utSSlngzbv6WrUzawkNinPEuIXaUqs3T6mrEBO
XtnIIs/4MqYpKhg59VqoTLJC0AxEqWE6v+9y0N7s0H8e4XrWZ7dvG/3IDsPLOZuH
PzT2Uxc2+EXheqUnxVkP6ftfN/x1jekaXpzqSJO00GVcX2eABepDsM59mZN6qrXs
I1/FLqjtZZtKy6vgeO2EocoIA6nSb+28LOBCdj2fBp/ZKJIFQCTEES8j1qTrZ89g
ODcaxJISDYyMKQ0gVt8PRv7x0OsD1QRP/ysTIQ97aEVYGEd+cmy4aGs6C8HaToP8
kMGJ0jB2X1b++0IQTwMg7f/VAPBMdO10V+1BeuVGlTT1FPBx91+6OpzPJaKrCqKR
fFsyN7WgS42R2V6wAKzMh4Ae/23xLyDAnfgqtMpMv3RMNoRlyZxJQA8Zai7/wx5J
QnjKNOxUYAqNZWXuV6/FgTVgf9OBr01hMj2tTs8RUGsCH87VGI0+/TdqUed9vvcC
r7evU9wwk5Ob10rljShOETyJwD2S19xcGqKKh4C8RCYXqfhm1FaYyPy8/xIVI2eK
Z64I020HYBQcFLsXkjF9PxxamUbHI12AblkmVpssl/oh980aHN6AJq61n3W0267E
4ybqSkfsy0Sxr6sz6faJAq7QCzWyqqjbRxGT48MiA64NU8z1+yb9RCJ1Dl6o/cvu
V7MkiOtGk1aE5Pv2Y1f2Xe7I2fiacol5lqZ2mwHKXksVRfXAR6cMd3q9Y7JpzLi4
SaQlOlORfFbkd0BqALTOJ4hXhCJb1VCkl8AHINVml61XgN8/if6XN01W4H1/VZEC
iG7lGas3zmMq4ECr8Nm5qVaBVaEvkGQo+0PD9TxiJzQinqxXvKn8avTYL50Iurg9
6+N+MBgShKJmQX45lfgoIOBodji0bCJmx5Vvk1IjmMgC4EubQ8+M9kVauUVp/Gch
3DRK5Gs14jBGgMjkdLPWay3eXfNTiDGeQ5u9Kkjp1hpHU5xnA0kjRUJgNW1Nsi4E
kubrC0YMkU+PrYLQB2Ly8jtED/bXg0kxCQZu7Bo2HHuUZx4z7vamxjgU3UdrgzTq
LWDG2W6/KHX+vFoILG65BVeAGyAVm/ARfaXFaRYUiRWIB45ue7pKEgfBCH36fift
PGWsOe9V8KD/11jslhoDT3RwvwJBwiPSa5J9Txy5m8Wvs6Z4uQbaRS2a98gdmI3g
GyYTuZ1MTnrEHuyIrg1l6l6BIx7tm1K0GbvmXzwzokpaJkAhIytAwgFmIho6I9z/
viELCl9/XLZ1FvSUn33LIXLsc5ycd8phWmtMbBqUj8KJ+6fOQArLueW6ZEIL5hZw
wS5+hiKUuI2nOYGmJpCWx+UMxkO0xLiBtbImiC6GEsGadeIlKr2/t+gy8IA9JJPh
6tkeKPrMG+zjJb05opdrDhhxgCsNbaiRISk7zvBA9uv1zFWY5UQb/95wy1SM548E
qby3bujCrObSueBBc9d5fvQQZp4IBS4DnstlCYT6r1h6cKk014x3h6U8N73anyau
wPFlm50EDPxS8PxudmuwZQEXTBcicx9XowwthSNQCjpGZDEhV6b5XvecrVviGJgo
9GZDPbDgCc3ne4P4hKPe4suKQJ9ar9eox54qylfH4jzT5s+Z8dg9A9Jc205tERoj
DSWBp5O3q+ntyTazAEmiRGBFD5+U8nW08+1kX9UNTGzCEOGnwnG2693ddla335Ph
NCeQg3On/Vjggv5v12i99g3l72sIOJX0zUd2sZlxdYw97hwpoNhSzLVf/4a83oZ8
hzOa1zWdMlUxvbNiLVhhVWMCGX3N7Ks+OWrtpooVk0/BDXaBqCm2aS143u3DMw6b
2WschrCArCkUjL9yWKQ0Hkke/Jbr3FNfSu697ou10hLKc1eJ/G5xRlGTHMTEpF//
ZLOD2a/Bd07+QQ8PapCyFHtSXw0N3Tpf1h/oAUFRWA/+fWxMZPzCKzoAQG5GGTFk
Mm7DjY22B996KpUd7UQt28dVHwXPhlHpzmNIKL4ih4Xc2LzXErDpuxJzlckY7UYS
WKwhGXnds4LCZrRPWaGdBlUKyUNe28aIiBfi7pkyGLWELLkFEiBloSLrIkFEeiy+
pC05W21c7nHllZFV4xffRUzIAtGMm0L+bQLmDboCr5obMXURvDoRohPCXOHCKiER
6m0vvmwDJ7pnWTpg0oOs4cz1pndCg7KFD+2oUSIMgRfAqODbJkYIjkb5AVh63OJD
6DxN0e1PyeWhvCINsON+GnS04ukuFl3iEiAfqZXsHUJFXzEEfSVWd4dNJq/y5IzA
n2lKeicE5Ccc3JGeMmlr8yAiQ8dMER0Ar28Q1f6tRgcMlVYrewoBxLp7geHa2MdD
5RODOOYampsWbQd9Cj3O0nX1X+VQEbQRM7ZU3rvj0q06hSBuqiT9+Sxv5nfh7zoE
+k+jUlT1FuZ09+rFj6ZBU4D+j2jBVxlnguRJDpUhHrMIbsx7elF2iGluKwE6jy8s
8E7D19I9FrXAPaq+2NnnOFuyRNqzMpfpjYQ0PgFPgIG2znKhhdv1qgUm/nEEQBlJ
KkLe8y+WpCDPt9CUazXoGJZb3pLpnhGrnNoaDn+C4XfZcCPhfrcgTGzGtf0B4396
J1zxdjlDp4mw1qNzZHiOUj+LWXjZLO/supqWFyy/nBxiBLLlfbVQV5soqCudHN5K
HrEhqM3iKGTEmsWs16NinuCeC7aspwkuxjbBX+7f+ztv0ywXcH/ZRWZOoRNgMSgH
NzsZfNGhEtXUh65dM/NcFbgRLZpVCkgBKgB2ETNPF0t6DcZvPbE1KIbXhmHVy9MO
ZR/ti0gNzpFE7C+Uc9e7E9WxzVY0zjWuio4QpUC5mCdsgeafr2aQA3PW0/EC5yrN
el7wgD8yeuX8cPyZ2VdyTVcmF9d2iq0ERSXRLkkzvd3iv3fyB+KPWp2N5wCfXj4y
ZRqsGMsW3cQ5aJL0vCrP8G0cI506nquVAg7bEy8MU8A5T40PnWH5TOYh7ixlkZTl
xWrpiFwCk1hIfpllqwpY3lwUQc4c3Xz/QzdvsHs3usuiqdUMWiiFa6n7+Z7qrvFH
zPqdCQqJ+X8xdDdI+jDf0FcygI3ULNJ/swcFRZjKqLZ1J8Jc6kLYRlDlUB1Gh90z
e1zTtRam6e+MbK9F7TC5noSgZEaBP4jUkKRa/3E0PTTAwgYb3OsqzpuQJ0COgXF/
jyvsrVZ+sIQmZycn2wLO6p+O1uR4LvH7ZvjSHKkdKAXVbSBdunfEgEqiyS7fxUzy
MlPprDyg84B/eQ3VACoYmEzk9NX8guP3+1Bo7tYmfLoK+/ZQb97BrieftTKuYupN
VV+VheyEtgbyoIv6mnNAgeFLUm/YwceRp424VrlFvJduwyisOJxzibRLL/LDBWCa
hIN5Q8ZU98ZQxPBJTzl073cBYe8XQgHZuQTejCDwBi1I+jfkRlw6AtYWrN6bY2mu
qjQWyn4oxBVK4y27N+0+C/7vZ+1PLYN+qNvhBz+1jULrURg3jGl1v54YBhBm0xw2
lgU1hOEf1z59hfo/dr656rk/EcNTGs6VhuVNMm8zjesTbk/Smne8fiQjE+fEm/BB
vBpUE634r8xC69L8MuUGoeFPcmODosahekhyR0KMkP0pDAno9yzKQhuCJZfnojgM
sNGMazqUasx9Mb1ysJCnYOeIljP2SWFVooSJ3yYDoTZvaS/1a1qUtEBTYDyQPwKN
tLcH6AYMdymF24FSeq6PSEKRr5QKXV+VN6aGDodCaDAIkil/a3xHyS9MShjY8j5I
5demhuxCC+Xv3XJRMYu7JA8gaT6MDaxxQSOHlYEmheGzwbpMvW+pO5lRe3Ve0PJI
97V37gAWUTCBZDy4HhIObHxeEJuobhrfRPsfMkbJb4d+qNv0nTg7GcNXMAKM/v8c
TvoepbOEyW8b8+MkX8Xaec1DRZpRxwCP+UF0JueoNYU15K2rRc3TEnhjxczvfkBd
QpE4eeSGTNQXV1wnjq9pqa+UYMRJcQsm6FNe7yOy115EXzBd4ciidn3IcReDeaP3
64P40uA69hhMaWNJHFEKMqsQ6mejn1zDFpBQuLAmmp6kFYzd5yi3MQ+tq1/KTcJD
Nsw9WiR+2AjHKGHvQhIAGlREgsuuT8i6gcdH+Oz7hIT1T9kWe1rHFF2gn1Yn8r81
KR4tWh5kJFJZnCtbZ+Ib5GKf5XPaX6x+9YNvSklWMD1e0YM8/cFHmLrgv2rETKD1
JH8Js2vflxhvdb4SxcjoV2MOAW4ciFvy10YbaJgn0XWvQS2bJsDDw/TT9Dghzg7B
fVU6OXlgjGvmSybiLGEKKnnaB+g2ZaPdqI0D2Yz7seJn0xeZwMad1QbaVQrrJfgL
ylR2ifBluEgpdJi07JH8NhAZjWjCRkStfxABDkhVlNUx0c+OYroNm6CRx3D60QI/
YAIQWz0WxBRC/6Z6xp/nuqxpUm7egpVmu9x2Z1LuMjdWleTz5UkhB/ahM2cgNX5B
tGWsT0gtJH+VhcJNp/dbUDl1s28UwOHzKiOG33p4+CxTwBu5mbHwV5dplT579Ajl
HUXDS1GvI0lSuCbc5klrjDT0Q5gckr0udpe9TpkBspBZhHTQFN50Kinx6xxHPM53
FrkFfcmbdOR/7jYsoaWhFFawsMd4EqhnVIkwytBYUCwLScrhSV6kThrWJzgMYpSc
XymC6VD/XVipNwBJg9YBXh3MwyBsWy1U/vs82uB68SdVafhxjiZLti5yLUJDEjoA
Ujk1leQhzLSjHb5ztf6H1IVVTVNuvVubAVvWZcCkyoZxf/a2shL6HTGOH+G734x9
6NOdPuz2efwq3vL3ep899oIcpJni+FBPcHnnBVTfuVTgzP31c1nRbMAzBXFZKi0/
u1gsJVddj0yQo3w5/lIT1l0Zc+nWkNEizZBljCI7X14sp2ivuNFdQqBxAq1Ok2LM
YotLvZkFkh3swdDERPiyFFCUazYoUFub9o8ZSTJeA/gJBEHE0XcH7VcPZD4IfU+J
aIu17vkqC4KxWDeUszwdamPxO47G+niAOQHJkgIBxidrHsr7V8++Bk10x1+lYrbZ
jzdpMwWppiLASpx4b0I8TNp8/nQjbbGt7RPu5/J24hiedSrpX0ngyZanOSLEP5ha
hzT4aXxR6YrKBY7VitOffmvWYBGH7GrwmTFXthsytM4JP+a9mYKkXF0QNhbnOK31
YQ9tAt+/niQ6VkBfKiGkZJqBE4oAeK5uG2sdEie0GtOqZxBFT/ms2nDVszU0HWs6
9/nJp5BlsZ0BpX4fhK4lVwBOmWQczBc/ux5wLIbJH1RbD12BlBUxzHfLJe0BvBBw
tb4l6E7Kzk84xxiCnMjwcDotXWtA5xoVKIIRcNXOS+7AjAfGVOrWXAQ6e3xTfDiB
2YVivzBZaRlleLyo/RzQ5eOjnjY7BRMP5grePTqrtcY+RiPSyfpfceKvU2sEaB3A
bmrG/H2JB3sTWz6/WJitkJ/u7urrbBDi970LZyNCBGGjWTmDlCHL/pV47JileV3d
c+I7sM4ggns8pkueXd3yICoxMcns5tg2f0EUeuLlSWqICgK9dVpxS2ned11Fyt+I
x+QEo8p9pVtxjgvr4Usw/85YplTI811UqSIj6NY4NvnmUHu+L5sjHj51XzA5pERk
JSPEe9z18gPRTg0CDzGvSOD0u6PYiFdrmZCszyh7Lpk4sI447UADktjELFBC/M7o
24sZIDT7oPLVm9PuJnbC3eqDaxUsm/Pv58s4rNfGxXJXJNcclpuqFE64kbUi44fu
73pqZ412fkjTlVKdC/PxHrZyGp9nfpeDaSS2vKb0kx1OghzEql+3pzA/YCXtLWcQ
u1BZ/xu7imWOCkmR5Bj5QEv9zgxe3J0F5vog0/9PpL7APGns+Y3TWxnhgKO7P9kq
EP+kEuSaIt8EVJsC4WbqgTZ8sv5Pa5Sea8VQJd9NWhu6lKHmDn259Q0KFAQLdiL/
JlglVlgtmkBbjjKqiZRzltcjbje7loyLH6cCzl3/T7HOiJJoregN6qMxZk/f1rxx
Ve1gaaLZ8OHOk1hYlQjr+8XZtbMONHfOgx94ZKhemkU4PmVqyoR8DO+J3hYeUfFD
+YDHbv4/Yuo8+WHxhfN4uN+ltQr0+I79IjkXR5rx7bC4GNIedfQIPdoKSC+k5y5q
HUmROqJFdcxzmUcOMhQh68VNznwSbZ5mCc7oneVf7NQCjpLKhYHL617GJJv/hHX6
3YEewk0qd+wqqoh0PbqrVXZYuhrdJRPrVmXZE+Ks9UNaZqh4joz5HN+JX0NMs9Ha
xVunGdhQNr9eGieXVeF9XlUHaupLd0K8Ps+gCx+Ai7sWU0kJ9X0BwxAr28wdX60X
ccaOkgO14RPLPrFmUe2MHSbMTpzECAunzE9LsjZI3txugFGywqycn9QS+DCf6/5Z
xxpg5+jR0VarE4RJ1lW/i6mlHe1esgb0TATYpmzTsKA0MBe/4H/cgqeIyaER7ghD
O61VQY95mV3LBROOxfAZDdgwERQ9b7rFqdggaKtf8IorTAo6l7zMnI+ogH0LPPO9
ONp7y4A+fAScUL3pgXvr834yLbstmFw0mYGPVU/bV+LWiQ222h6iV7Fa2CPbAQA2
jYZkwG8WQeDKUmggE9lubE5EMB+VTXOE9EyYEIB8lmXmUhFYIHJdiDHB5KYAjC5N
M6f2NjG5Td51yWIifO1dDZWgDg6nmcqq7J119Ra1KEgXnFOphdmYtSQ71mpbDBCJ
+PonoWLi6FfYJurgZF7JcdZi+Q6bR47BdWFJJlHN32H+PcwEOYtWRD3wJpM5D+9z
AWbb+iBNIhFTUa3CQg0ge/RFN2Fp5Ksd7IWNTxfeNzKovYGKozWJfl3jjnPDkU7U
vgNxbkWzHO7B89Bx+gAshMxKdJ6RWEMhtvZ+cgakIW/RBsTL8UP0rUZOYSkAVqx4
osHAAZCNG7Hqx+ZEznlvsAaqr57qQm10DVaj4VQMmCGY8jft3TyaBBO+J4yNFBUM
TL6vdZZJGKjJlIFfZBc7bSG0BNNd7UMm9nG6epZGl5+78RyuqAaOe22qEp3L7znQ
63xGtQyo0q2vaAtPCXL2lG7NHNbjZVvVAFwvSTmvWpDqa9pa+s+jqbqz3bhP7Gsy
4GeESSwCRi8PVGRxLz1wR+Bu0prImia/y8t/dylTRkcNlVE8q/hDUj1YSzIKwZbO
iR8GNJfUD3CmaYlCqZjut4TrVdgYGaRGRGiVtNzZ+SywzwmvnQK62Un3RjhU+lJw
fQlKco53h6OCJopoFOjwfvkxXxl65RtWtpC13/ZHXE7E2nkxPi2n/ZTz0saVKaKX
S39R5DhxvJlZthCVdkaN2nf7e/QoCLwngXuPaKLJnQcCzEoJTCgVzs1dqv2/9rUn
8+6G61eE7oHgKNI23zqI34wMQRjH+y9Z2BMH40voYcmPypCawhCI0q42zx7CwKY+
0KBsPBqfxVFwcftKDt3GaydCdbXNXFeFRR68hNV6nnfuueUbbTrEThKOnNcdl7YW
9RDrZ8BTiixf5jfJ+NbPFkI0GUjyrbEtJfDS0u/Z+InZuLij6+VGd8nRjQsKJk00
++b4+no6R9mzBcEbTYC5qIbWOLByXF/8Q4kRo8AGx+kMvrfNITGfBYsy+vLZIizW
s6+MBoJdMh+6X7cCBJpl+0dPVJYaHAYv8F0zmnQftctKAHqA3FM02OmdoLKuSr1s
pPGgSrjgtkjZ+IqHUEHMy4iE87DqMKZ2BJbY+ix9hfKfenzukEbEixPEnWrFeRkh
JjbQij+BrFjsxC4xSOWP7fQytof6ENluWHrsclPvKWq29DWM4pAVgtoljonVeHTQ
AU9goUw4kYC7WPenX5F9PHJHT5TWIjRPumrCdcW1oUcfkYYRkcYeYeqF0rm/3N/K
614FCTW0GxouB3sAmR0hcLRnV7v+k4BvAwcvAuS4+a5r1NKxtXdYe8qclv3erO6S
yfoVu2kufqkboYjdCFxJ4S8j0bnaPnUkbVqCZiUeCa2EWPDnnMHxM7WXv2y/s0GR
XzPIoqSkd2CWJnY7OnTipfxfO22PleXs1ei5Vwfq6dmWVRbBFTORPIog3jdy5MTs
+cmx+0QLyZvmamh5PpASTYQEUn/krJkQi0hFZ6V0WQ3tQZMH7sULu9b42Y1Hf5mf
JgP991UM81yb1qVfBG6ygsasQdwnVB1FKrx7iXS1v7k0n9Nn2XA2nArGQ3mnrNNa
t2O87cmfb974rB9/3jntTleYmv2ztTWj7T2FPFDg7DhX3lqpdX0/zUZMsNwbVsg6
GqCma2BS2RwhTEOubViXs+g/7UyPNqF6ebnUK6aj9aPgB0upheeiQZokm+qHwXtU
M2GW44blz1glmRxdKDp2i9OifxYuqbCPypYhx3vd/oHRtDXuVg2aPuiCCyOVr1N+
jxCigM/Vze4HSElJPLeZgAQw1O/sb5eXPguPBKHftyF54utjG+vjWTLhOKJ/34/u
sIBoq9nMwEqcQMGJXJpFUx/D50HsneLd/kwjyZhr8R7Q/zY5vR0yzC4lGRx3g7/I
w+eOSrNNmxzgLX9NCcH/4O5oROquBL9AC6zkc5PyVY70SN0bBFHecLI4EftcUHel
lIKmYA8ALBNQYLMzARGeOIAX5pklyuoZDdERsaCd9Gb4cgBC1j4Sj8tPIfCxuZcx
uTe8FG6WMi0aYiwn6245oMGVmoa9/lv6tyATir4+4WWmdYo6IOvANg1JtnItysJX
awk95dxYa4r9BkE+aXAmwQOSMqPXjmkH1PqLDXuCo/WGv05SE1J2cL93RxHJdla3
E9X+H/Mlj3ZtRRrIvvU7NABgva3D4yiTYX4G9LO+unCgz3lF3nzQ8EPm6MtdxDMw
SaUsGENZeZDRGu549/guyBzIevry9xlrl9IJCpnb9+b73+4tkcOaDIUMQkVKrTk5
CnqekNyWyz6OWnixT99xmeKwgK7IrBy3E9PISttBvN020aNqwCqNX5YpYcgg022H
vE58+v17SoxkiJ/I+RGWGJPHKK2KS8gRp8BZkhglO9SWMbxL5qsbV//cSMKJTkS+
jmHFYyYKYgYsWcCvkWuUbd67MpIhMRXJogMs1yosRl4ongcVK/g26zFD7INURYtH
fM3Tqz0cw4Ml5UvNF6CPBl4izJnUkc2ADa26kBLwjKWY7r9tjbGqNVMH0JHxZKDs
br/vVFTrhWB3xGGir1Vuwu3vJA7auB6SDSaO6kSb/aXCp7lBwTEoozwlvFi9gmgp
bCGVKlHhIIST6SUjkV/4UWh0SudvpXacJa3rljVok41NGwAmNCKqnfTwCuld0GJN
sbuPOZch1cj3vE2aDWKTYY9KtM4R2j+AYHMo5NjnW/6MAurL1eN+kEyI3jQmIftF
nbWs6BqCFnBgP1C4TjxblOaMz7kjyN7/ElayUtkhmVkddJWbDCdrwBN3wlgJhgy1
sjHcWvQtq7To6J1XLP5Cs+BsMeihcy8+LZ5QeFFAi3EvzeTXfQ8Yb7IY/Fduj9wx
gy5nHGouhshYA2WNrG/Nb0k6UZf5bdI4U4niXHWLiD2A6d6lTeIjSspnq8ungHFs
7xe7DGqrUQ6IPTT/bCYatnjZxjznGQU2Z1XcHb4hmiOlXdyYYrsFonGyeZTEVFv7
cSisD3jh8BzC3BJERmPMxWiycWMM+7gTQBZm5tmatXxGBqTt4ghrc1UjM0gy4MUD
aLR5vvCxb9bDmQdqjSIPmJ7T05PyJBxdWeILf1P1tUPwKDTu7o7sQWd17L90rZdj
eBNmYjOuVlk82sfvvJkKga+ofSsmF8NOvGul67WVXYdikHG8L9660pKgjT0gdFT6
pqXQGWoH2YZPIdx6ojMNjbAACunr+eMGXgqWi0IOmT0L/+iLf7jG3Va/tDUsWsMm
XDlejm5GFQYz6U4dfli+/z8DofFJjnkK3C6sfdI3TChg3P/G5lnpem7hUsEZCK+p
+VoZLMskm1/3jAosj+bTyaXGg0RKBzeJME585uTqa00LHHTtlxPSBy6O4vqmnA+2
2YrR+W+TujID3IQcxluUHsL2ovZ3n+0tfxxYQh4GqqEQp8qiz5g3dUx6SNylpu+u
wY+m0aLwyHFcINCAXMteH+h6odSWsc+43pprgviqaaqC704Na9cyRFlvhEBWDwO9
tz2l/Br6CN9ZH+KL6UGD3choBfj0EjsHvdtlDGd4SbHk1qIuFgFDqIHUFRTSsmwT
Ed80/6Sk9G3oKowXlczSB+vgqZr3dMqAaI2TCYOcVjGQd7pBzAxlOzjzBKHC5bYW
TC3C7g+Lj0DELeZy+ZRDTUnWZkDQeQLw6Mf5nX2U1L/gDENwsVnS6HL5u2N2xzid
fLdC4sp75rlabQXg9lnReNGoAyfysizVhmdajBJ6xgZGnSI91YicgrD40fqz691F
HCAvXi2huMnyhlizAIH0Jz4ebW4s5eXF0yfCeapdc2F+t4Ha5Ss0JZgJ9rlXYdvy
zgIBF4Wg0RThJDgA71VD2qgMMVRL7pJ7Zm9XDe6jgeHcCxY0WoMfEwaEEhZmW3WO
KbHedbu6OtIMuswG7nhr7nC/Fi8Q/vCWM4kbB8Oxd73/avmrBjFoiDNzeZmxHexg
60Me1Ub+62hxB2KS3CL9Z6rBt8xLsByc9nxCQrKwJh+1uYmYjGA0JcxnYEAfOAsK
xXOlNgqQDPswhhjbx9mTqHE53ONlQn2lqhhlYzuEI3Fy9s1pADstPXz/TO6pYyRE
xAIerwpmse137ZuXBsUqpnnjL5wV3pxBZI5CAEGDjZctz3TNtwiiimYh/GktMtKG
HmueL9AKaSrRS2QY9MGzjKvRq8zfPi2trKoiX9KI4nwrj114kYZKKHNq01jbmPm8
99iixHu9sHLcrwlorhiJVA23ypb3hQpU+mxCsXclxQWkcFwakobLv46Hyd7WNZFo
BRCQU8jkkGQWZE4Br5J6P1scPFWXKEOL+svkEkfAcgJpRxralNd12fWYKQ9/K07N
E1cifrjbu0U1tQaTxL875A5gAfH3UnG85XNczTVsHbvGLvTUnmnEUtOTWjuIRCaA
q+aNmAJL7pYNlNlGISxyaUpoc31L3SD3EGG5I7aq1o3L4LwBIzV/TqYUd2kLccIn
dA2bN+M9YQrbMlzKxGwK1Z/gM8ZOGczstMicrqmPrXC7NYhlhAprtXRN61BuLj0m
u/AEj5tS+pk+rtyibk9DBSDjrE2YBMrnUib55kusLp01sFOVebjQaehWCx0lSsaX
0qgRnPHCMaVNrQEXnAAwF2iOA8+d7pRsE5M3GIw/lm4GXR89q0eTlpl34+MO1+bX
iWNpbb7sdnTChcS6IiiMA8WJduNCE2GGWnLv/QeEwD1ka65kPZ9wq26uO9ifiLs8
9aqgdq2VuBUfXmnTYYDGbmnH/dSd4NJmYWC60Vkfm3YdTbP4281YO9V+VoWhrWtk
3jeNPxq9Uk9XnA1A3zJZUmr4Z9Y08zCvqNnTwbLYstlJAmSGSR+42z3I7f2N8Ukm
RwJazKrXdfXwylDVO4bXNQOQiL0VRQXdzw+1vNo1l5npY122/JXngUJCxvO76LeG
te8x9cRfx8JmhRIZKWzkpcWLi4K10/hik03Jo72VA2R48xqJKYINMsvf1kOcEk7E
bCqgq4PUMsEdAO7Y8gSuT5Ro7oJMvy7EkgcqJG31LZOO4dIiKbXi02zO9+paMJA0
zD8QZkb4cGPFfdLcqZegnzBwPJXj5iOHPVku9AyGqtdOdJP1WRXcW9O4Zcsbw6ZV
XNyGEnRtvJUhPOB74QcJtjG+fu6P2BFnDIyRWMwQjrYXcEl/d7T4ARgQEIRWytHY
r/3QYLsmuQ08Rhr39tIVW6IIDBPS6S6amk0lxWPVRF4l6GrcEW6s+W4ksL57Pkd8
wveFy8ZBujUMv3Jzd1MopqA/4Npb9e8Yian6dFPmUGWLC6XkmmNmjKd6n5UgQM05
Mye0cSiHD0vutliTg/9RrY3lEFUmINHSWD5rqXfMrvQueWytjoqSoGnA57EyH9fe
7OV0W/Lvtk4emJD29nm+eSVbnkPRY4QmYnqWLIdFZKpp63Al/2aKda3fk/mPA/Wo
C7Rl4Smzqa03dxV/z1Nq3UkjJP4VdOZBYi6UJvjz+Esn9rBied0DtJ2WVYTJR6aU
D0BN6GPpjemTwI6hDhFiCtwb9vXFElsb31N7MM48Ep3Pf9kOuWjWlZtFJSrv3eed
tQkvOKIJGyVapQ92/zmCA9aRgdkolEBSo7pmcreBUJr189SteqwYj9Vu3x0Ulw4t
/B//Gcgl/zZdC/zpEyD7KXri0oNtSXGSXTzu98ayUgxnm2+1aX1GrrWB8mr20FDn
tjGMj2TK5QTH24R8eR3PK+sPmtEmT6ApHz+tcbHpUuvMWOo9pHNU1JMGcUBUqMrC
5ZV2pMWWV2EuP7ZUIYDi7yH/sg+AvyMa5VNGbVx5PM89psRxXfNq6/XiJILghMNM
LPblnUK5XusoWk5ZvmcjwVXVYgFZ0ZxvR1jNhAqXPB7HSdEkhsRJj1bJtLZ2rxxn
wrHsHcO9VV0x6qFGAbSjwE2L4QrzYfrPa6zVwNtxF7lQm55FyuH95HoIPBsf9TFt
EDdfIRCeTS1F0+8Otq9JcV4jiW4Z6zoXijfBCXyIzRfnMFycePfxNttPVq5oG51I
Wv+qc046iTgElSA4a7/HDjJIpKi48WV4rDsfT+LxJ28P94WGeCf3/DpwQ+AWsOy6
zC7Ktv/aPhf52nWfwT+WX44sEiPq/IXGE+gg5aobEU2OXxnpf40LemfBajmcQlJX
UHIBB+BIMQRwTpHRLFtqjBbcqRz99OVAddjkUxW/5GnSC7fW7HuLezgGzI+l5B66
H8/rnjRTmrNnyjSK4wVu1x/maMtJE6JTYyJoXbTNXZiwjkxIhFuCi65jS+X4gtx2
gSaaX8PyYgwl8qHzb7d9ejuQgo16/T5MwFpqLfsPaXM9tqvfZFLrFMMAPahECgth
W06YUEO7MPr1UBeAqyBioa4mHo3Qafq1FYQqhuk9GM7URb9JyYu0GtAwXPU/zREV
fM+bC3GBfitBIdIh40+OhYMJOuzl8AfsLWi4lamUwKUMVj1J9zsvWnxUiFI/7J1s
vfog5Ig4fTdQkxL5BJbjHN875n4XEv1F4AnKwPU/BKXX5v8DCEymflgXRUhn3Bpw
2MCeC9pKZj5kwLheGr0o6XBrAMTjBtxR5RbwNdaRE9Xrrgr5LKH2pMe1JghK/1KF
s8achI9mDJlusx8s+gnlSNr1LFsQZMZ2d5FrQ9gmzsmXdGoXwMUrf+wZcllrc4LA
Wg7NEGMu4lTZe8Ol0Ol4hxTWIW4mSrm3O+RitjQDpYLUAGayQ7Utla4k8iQ6keFS
sGdpdVUxcrMnU3f34fi2hS9kVB4M2SmpgG/l2Pu1O6I6CLGBY50gHQNbOZvFczNC
IAyPXhAdWpwxJ+YlpUpwTx5XIh2wnV+RsfmzPRgMJh8dcZaVcdv6CGPZa1TouyMx
0AqjW3tBO1GiWfOOzvLM9SLdwOdfWEW9e2Jl7VxAI0xodLlskdA7AdD6gNen7xX9
xLn0KDgpa0T2GJGce7binuVNyUO/RGnsV22zOymw1xUN0fobD7DbKuLXiP4lMCSb
NlZdv0JtNlqUsV8htwVkXOT9KD4QXqcN0CcIytNVQ1dkwQtXgT2pilCQihucy5ll
mW/HunlWBfmAFmX4ToQYCTdgQ+gWztQ1ywl3O99peo5s/FQhzPeGtJa2bFE8LuwI
amJd9Fo7OltEgfIwXZSkZ42Bj0Kz77u+Lv3qmKP1EA7lLDQ/W4xaKag1dblQ+GPa
labDndkSPINwYf6nt+lgDbJDkcGOa/1PcghaiOoL3894RiswGElUtqCnNxxK18dU
brpbzD/m1mAk8rA5/192htX+XF44zZqZK0ZaqEZdG8c1sYQP5Nla6ZCw/qTZw7tL
2lHTKS+20pExwxPyKxRmS0fZOwiLbaglWC+HTw0HO9M3Or+mGPEEko/GQd8SeNLd
5pc0xkf2FExNsy5KtHV3Tmf+Yvl4mnNsDUO8I76bKtKqsCVHemfUslH2A+IH99iP
674vqzc9FFxz5nncUwU2WQLicAiv1u+8WglCbsvU+bdXQ726rrojtcHkSzjiU2gm
67Rtn5kb+wIGhrjyvPnHx8rAjiExmr+yFV5IkCZXr30TyxEsA2a8Eq8Da5o4Km8/
fQEQ7/ZnZw9mBNHihe43n5msmDQ63JaninDOYFUazmJ1OnxpemmOQs4S6rzz9+dV
2dPdGIKRobL8rie+SAZuNEv5oa0PN+LHVV1JsaYZNGlsg9q4lEC1I2lTAYy5ezj5
FlQSAwKLo2X/05CHTx9k/dl8SjJL5HpDb79WZ2f1taIO+CKyZK97bnHnfb91JOuT
4mPuC+u7dDijxC6MUIv7JCTtpUMlGJ5KXTXkhUoys3KRgT2GvBbNqHtaXdZXoQMo
YpGh+IAQeD3o3WWs4IUKEQKJTA/DJ5EmVhK749Ybj5EUL8bvVupiIVHJTbpp0M8T
BR1Zsel5kbYHYykWpHJ6XS5xU2EBwCrN4+eUJUiI78Qhn5/Qo21Y2N5M5ITU8ir4
t7uV0Y3uPCM1xFxece3kqaOTJxhU85zM2/gIPv3D2Q3SefnoNGIjAJXjFyiIKqef
f4qTBd6Ous6+gib4yzZEfqObWK8Kp4ey9MBLIzdGbtU7wDsjb1pP0jFZSoPtc9n/
c9Ap+msKMmPd14GHQuvTJ7LB+FbhzzHvLvs75EPFVJX29+WkSLJHDtUJIpB2Y/PB
QLFMAvNxGZkMFJ29jy2gQPIa9vhtAy+ieg8eM3RG3dFSa3RirNopAVCezmlbQO8z
SW1f6YCijqMShgp4N/kvsr+9hPfyKPHV6Z6D86WBJAT5cORe7v5LQTiUE861uZ3Z
7Y/+olCUaTY4cl1VvF/niscSZEgWUVoSxl7GIma3GQvjCLCJ1pq/7ze0oaLymvF5
i4+CcUI7WVbQuEKEEdSxs3Iott2wRQLf/hB16BVKpt/4dFHRIXFfKO0dFfjuzx/K
YED4nka+cJkt8/BOgZfjXT0IH8yjd5rruGbIXlKkfEmHUxdqiEZlO4fxsFtsarsG
5CrxP9EYN2EIV9e45IyegiJYkWqAFMJWlWJYd1qB+b3kzOZ7FNC8Z37jq7f9VL7x
h2QVbCm3wA+rnmVmXO5Z1IAREpAnxYe+H+vtgubGjC+QUUZMv9Ff/XNZq6P/jODb
YAIW7HRrENlVlIBPmKzCe5KqZ+k1WJimAVIuBAU4iFNqd/PTsjwkUv1TDZXCGcn6
UI2wROvg/Xmh2O9RpiMdELOpOL9R8wOiJ9L0L5luoS0w4Qw6xnHxuxeCEUNMkaWq
VY0ewxFq2HvRcYtAvP3X5gfDRrjogGDxuI3w8XrNlNAMAjwZWjMs8V0O+Z6X7Ew9
4ZYhnpjb31HrKPDDvynXhf339Ne2bBhH1ExEzlRaSFBqt380Z+6MSrcq5P9VTl3/
JdrdN3z4g9XyLYRxdGwgzH/Vd+AdbfArBWHZc0l63G2EQiBWapgmo2IDiH1R5tQ+
hIU62/qvodgSk5YioJEdnOl4FUf5PazhhphDf3Txra0FfMssJl15ioVEeryFuLnq
Ar8B/Eoa7f8UCH9QOEpvIbUzpDChYrqpPmCq6LqLgG8S8GcwLlrBXuhjsPkjVY6D
2TECtK9UKOGqE5zbq3o3FeMLHVgsvQl2C2LgOZzLQB7rtxHs2hhAD6sgk9HJWHKf
XFVqBChqLPXsCwsGdwLdOJsVl53YikZ5WwrIp5ijvTnq2NAlVWXMg8jzFBJOp8MA
twlpVGtBdAaMq5NS76zWc4SiTD4VsJJP3MD/3YxQlyzlQ2MV/S4P2VB4IOnOb7+k
NEca8cCFvs2+fbyWzXOiTcfljuCCFD6CKtOnRvn5zttzg+nOjqWTp8G/hAv3KjUU
4wXKOlDJSMmeFUveqMJC7vjn4rDYELIcjt3etzUmDSY66UZ2cu6b+HwS2vqZQhj3
jaMeAUdwKHqBFCgEXqKOibfb2hWgrRUh49fgf37xNL/xfYJZc0F0nWxnwlfkLBqc
qA6jul3qAQ3iuOiDwm8TSkK+iyVMudPooxsqzJ3egsxLGwkPqWXBU+Xi4rbdhbBt
qVE4NpJC+BWVwPAITQ1iCSmTJc1qTo26dpClLtEpCyCIDH/U40MnwIGTcoOKZFcR
FF2FaYgRQfVeL8PmlE+OEW1uQCzU9/rYE/VxitftsJpmf1PFtITXp/cE11PVRB90
58etWxPKcez5pH2EBQimM4DjUv59XVxh0hFXD2NerwdtCOggxv7Js97DS0hhTbFC
cT4tNs6Z4LssRYeq9DxIfgu5oRieAiREjDGuDC4dTZ/QH5jRYOWU9sgxu540D/4v
k0/ztyVar5njAju+pbzrYIZ38OWkX7L3Me+e+Uy+Vvwx2EF+AujerhmcBFi6j+Ie
bBOXpPBWH76ILoHNGHb4M7hldTZ6BPhsOc9E+5Z03U08eWJfLQCkJ5IOnVrRV7/s
VMwmMVZg79Sj1bcWOhw04T5ZaxsEnHmpRjsBoNNgQ3bHEEZOHV0z564YeH4/8d80
JMGETKjWZYrHaPcVScdorH4WbP9jLy81rWuyWyvJd7Z5JUoDUeSAGsWcyJVIwbOu
qSY81I8L5eoAejVzRXQXpeeNDjHe2mWtgrLoAEqveyg7z7iYJY33XNn7XONuakSs
235LLo5j/NgOU7M4Jx2ZTe/EHUA/cIraab1x3GAyJgVEAFTAcbAGVsgwwjWsYNmk
+qy/7rGoh6sTpzwKV45g4IykuU9TFJZmeV+C8ZI2TlDuXzbuq/OdSYbUZ4ZvZmDj
z288b5Vb8fmVfOACW7S65socoOkmYNT6GtQ9w8Fm2Ts4gh7udMc2i7TED9su183I
VhfFIzjUmvNL/+xXeb4nVQJ5RiUF5OCC1TFpCT0zs13wRza5lYCbmSSWMk3L7fsU
9eJQD8tCd/4hIou8MS0EvQ0DspWbsRkGLAybNzp3GFvFrZ6kMDR9M6PEuhK+nU1z
8ijWsIvhG+K8k1Nov/OK6AULTlpzoEyFQ+D4rO/u3YBKWsNl4r5Hc078+D0RPjIO
5L29fCEe1Fs0c2MCj/50Eb6SMupREtobV22RiBJ9m0yk2u2UVRuhdWNbtEyqOA5H
O0ykxbtMx3QdeSoznvZLohEFnL9f3ZtmD4u4MnMK2f3rNj78GAV1WxpbuNn9sqSc
KhUcZiUG1YXHj9wnx/6r6r/vpuWvedmZGhOzHeUeNT5KhvGzqr3XTGV3joqy7fZb
r+YhGDyN8QrFjEgJBc5v5cwqfSaSHZ2HSwzucqNGQ8F/3zKEXEnHplkHLn6vteji
fb4CCKjCQaTLHLFns02YOFFlGanrVpo6/LG7/UoTqAXd2hWdrdkQAQ6s3OCKjp1W
nyicFOsGkcP65jULqtqjmCJeWmkgYacZxNudbWhrrX7Y79BoeP00sCKfCDZwJorY
lU47ttz88Hs3oofZjAEQ0cFSRuhNPpDNy9m1R8jXVTbURXk5DJCdxfzAoeaek2TU
9uuO9jK98wLYlqAJzXxIkJubaFDsXscUHbRe8TJIrqQHzy5M7rivBn/e0QlQssxa
wQgXNTxEApSqvL2uqrXOAPVSPamUNbcuSRWkaLoej49lUpnajDMrhXeUgW7PAyop
smjKAIeLzfTQ4DimxLFPhbLvdv19kBhSyaN5cqMUF9izzx4ek581ccD0wpcdNUTz
5jWjxtfbIpKjGlx09DJzf1i3cq7rqG+SKhO3OPqhwVR0YyysiANHJOIAjp1ZX53+
ZFoJ6zAfWZ5B+zeL0kh5B0wHEMts7fizzh5BdpOtZBoY/P/RbdojAkODntcATKFm
RlIOjWVibVShMlTQQjxAt/kZeu0C/0Alj3sjDxrlIiUvJv6+6eC/PEFHF3SLXUWU
JvoaeP0vqlpN0oYdlSr5woR+Ryvy+kNRWz+pNzYqGSkjAj7XacHjaNfM2dd8KHxo
QhCUR6il1TAqYHkTI4fXYP1IVBiyXSYtcgTiuSfvdD/LhoGS5c4Pzk2MeuZEsXP+
H25zvu9oPP2VXxkqOsIztKstAQ79r8mrggHRoh3zGwbEgBrpQ/5cbw5Jqf/0BbAQ
vCD52ElX13IjW3iB6CxryPWVAzr84GqFW7qBEfBxcTwZp04VBpnkgkMSvh6fRYAO
FO5iKMV8LMU9QVEfilj09BWh4PjBgL9i5AieLRITo3XPgsYW336SJr0jEYx07Wxa
3xT+xYXqW4oMMzUPlVUPESwdtirjBqUGkdgmaEcL2C0sDGjITxmycwZ3wymSuie+
a4L2O2jGfXUGjHVmhsSIg7y1cPIXn+GUBCsMxolyf/emoaFSbJ0rr+Rql+nzqAw9
wpKfkH0hUOuUMe4eZUJ/iU74y4O6ChESZ1xB5PyWQ2/4LxHIm7VWfP/Xtc+B92b4
TjTCOtVdkxtH7vEp//E3eB8HWUo8sR5phkXdk8Iqm98wzbLVglo4t75SJKE+IRZN
MISOkX9lUuDFUi3H9yLvVKwvcXXqJ3J5ERDCxkjUp5rDx+s0ijh2tfGZnZx/LqwE
hexkYcCJkTQeWJZ9qpBNTdLOgTWqK4E1tRPiJL5N6DoV7E7ocmaithbJDA6Qijol
Nq/dVtsAiOANLjbWnMIV6YU46VXKIq/FLvsOI4J0kzho09JHtXGsHOJBhjoS34pI
pJH/4grWFqNWF/t3RJw1bqLd07bJ0KzNEtKpIZTrIDDYDJAIxhnT9GvGWRf1G3gd
M+Cp7Cw6d7NUHfsplEyrieBYF8ejkflIVl1FXjdss+uh9pi7gIReaJsD1S7jdg2M
8tzD546vDAwC3Ix6JC4EJ5cC6GnGWGj49/AsnXslU+AhCdhY3n/NQab6hPEVzzF+
f6LBcR4DcSIoNa/1FKVeDUdtnY/Lmk7Zo0YWCOUq+LeEOXB0pVFLusiYaIFhfa9J
YGyo3r0xxiS72p2io8r7MOgz9T8unBHWQciXKFRMn0ag5mt7E5wvOh2tNPfd9kSk
mIUFcASUcR92mw5FJxcTrpXvqgi8N5z10kTs+DiZtfUz+cpgck2TP3GIL80pwn02
Hz1zu7AzBftMZIyEMk8BPNYDYlO2gohLvV4WSYj4dXJ6Rn7bBJZ8qe+E8Rha6k/X
1JxAWUHlg65P5IGt/zlOlKd0pIFf9cpWNW70m0RW417r8bLGgbjBrjP4FWpK3klI
0+HPOWuF8abMVY1xMR2ibm6nXQ4iLD/OB9f4IsrDq6719elFp+koXjsqjCwUpKqn
jVgfmT23LS1Q8BpMoHozmXu+tuckhHrajNSVdN8EdvS+uH4R94TrLpfAawZPBTJ5
bEM2XbmzlqioEUMzthyxDV5yKw30WVfNeTuF/6d3WmarFy8M7KHGGx1cMA5JdBgH
e/ClMAwarR6IlQkOqSUowVBdhFzZoZqUT7T/nctqIb6xG+s/B7+1IyRHrpFxt0+E
jNKbvniVIY/EcZvwx9/foBU0+zzjBQ8iyXdV62QnKzTt0u6+4PBK7Pp8QCM52Llt
10CdCMZPeFrOV4OIjxA533kM1w1LCD02bXfTyAuoDKcLKb5EqgChIe/UFU+l849u
ZH7t3S98YTuh0RajHuf9Gt4c99RWQ+FyN+H/1yRELoID6UgKl6OMqDeUzKW+cAln
zpQ/cWPUCRb0z24szYAtL3DCnACOW4mFT3hdDrnjtjYzYzXhou6dm+/WbFULNsZk
6jEkcIwmfmqnX2EsiHzdaHSPKxjH+FOQylc3lhpYdnPInB9cVOmVYH6RTGL7aeFi
JoImyL2Pznznp4zn4mkbhsx4wZaOKn/v+QVuDN5i4m9l/N/A7ZEQKqbt2HQMzGxK
vQ7nShV0lDJQzU0cCJB5mmmO9kSH6ahC0g9tIhirkj1WjFc6f91oSEjPAXw0Qas/
otCwvwHf9qzKsD6O/aAQoXx4m2gVDxL788a4vjn6uSmVdwDbhVlpIzu0lE5EaxXG
b1BrS/pYkTYZdG+s4R22xve0+eDg4DhrBuTDHUMK8Upn1gR8pMAoamoTa8wph7gq
tMPFkfeYDDNAuHcxXQJCpfRqXsmUz07nzPLkU1MDN9QzUgKZUJYLbWr1Bvt0q9uo
Nap7s/txDlRnPWm39nPszhlG5uF15+iiGQJhVzUKkXrkIn3bfawg2NDhbaWF+kRr
/wJ/Duw+t6iRwrGLnlpGxbVOGgWwXy90n++NUEFO/73Slrd93TETzBv/SosSCiis
LRH7PEEsfTzeAQTTP+U1PlKEgTd2iVleclq2Q5qnSKNJ76LIWVZ3ZCis41MAyBqu
c4Q+tJTi5aUBfKVp1cEAyaTaj3XzGJPILmuw/tpdPEFGHGqFXoxbD15rpGQG09iT
d4nvBTqC3JlPxz4Ap/RMLNuOw/jMVrobC2iQs+yTbrORc/PjjCUaLAeUx6PYZE+Y
2hdNQaccJW2Do0wraLQTM/d08jzOqNdYeZNezfW0VA0HB52cMD3Mu8j861f2CeRy
HszzMo/S1WWROO8UZfFyujKrBCEbcoyMO/ubEg5T2nD8LXxpx2WTl+/lyyTEgbax
3zUO0s8E+7toebIVIDByvKroPfNBW/bOGjqc01YiQo338Bv/vbtWupMQSz/R5ul+
NjpWKV088gegxL4FfU9lhObNDFiFC3qCP0DIY+OxpGbGEilK5ShWarh9BfqxK2Ib
REfrjGg0y2P6FN4ef6zwKND14svkCeQ8PBMb1Tj3LAjF+oxT6lSyu14GXctdQCfh
xadqnvLe82pqtfpDyeT5Vu6S0znd+6UpcikLZULINfJ16DEeRMQTDUZFnHqwkjeV
T712dwvytgDr0l61ExN+G+ZhDJV+D5GJq7RSxXHB9EW0rdOQHP2UcwK8PX2XzQ+l
mYGsvhnLwbVCzcAfIGI2iGzvKFnpNmHNMZa0G6h8xY0EmuoEuXI/qzlubLAJLKkR
/YqSfQSXmmeb0cGKuhV1Q+Y/ou7/s+chGjYAf3FUYhYVocExXfSTXeu/toqQCXrQ
56Xb3/jJBFP4zQs564qo99Qh/V+3ed/qfu+x9e/11NE8gxN2DZNfkHQWkRwZY4vQ
WDEiChG1f77lDVpb7844BNldLZmsfhSK4ESuiTKs9koLViaL85PNaEh8mRFRapIO
gkqwwBUlVfUY6+NFCi2oLpuFZPLWuqALEoFV/MFfOpCyftwjbZn0eXjuy39VW9v4
9C3grtBKzF+GmljKyK6T3wkT5IG1mboI0YQtihKk//912DtTe33hkDSoBJ32c2IQ
hfXFRkQd01zlecaB128T5YnxqLOGRiijfZhjcxaF1qqgMNZW/mthbVqwgHunYocO
a2AYDq5tsQSZe5UOVV0vg7x1KWk4nSoPJdIUhIHYfzX66zSwoQHKi1O8W2p5yO8x
6Zi79HcI94Vc3Rki9BmQuuC8Ob09PG2+vlbsq4t8QBk0D6dI+inX3VVazX2I+5+A
OGLECR9PbbU7BdcOSnyoxpPAdIdBUdWrUPt6uLyFDeXUzGagfI6Mc2sloeG3GFBi
rqT7Oywr5vBJwFSljynlOtxyqaMrDEK+jARURANF+gWTz6QNfMco/ltgo66+3E5V
HFQncWSXVQd9Xfi7OxpsSplt6ZwTV6NQHcLnAJYHZHEgrjjKX8Q9pYked+4cXu6E
+/dDkpxmCaOL4bQHnY34hYzG9zln1dQd4UF+mvWlmsGDULhM3r30xuGe1w0ezAmD
mN1er4Eek+VJwmVJY+aZ+D5QI8/n2VxmzPwrvGuwkFSYnzDU0aZ0CDm8sUxPN83C
rsHr9BObUOoSrlQ8cssaDLcuKgG0PzaAGPhzi4LisX19s67jWLQrG5mSfiZ9nIBv
qD7SriFwpvVqHSBx8pHr/cLaEjtmMlrRayrTTy0N3yc3NMjrXM1kMHrRQKVpjPHR
2RKFvMiKEINP+lLEpv0xN8bUj0VwQa4bMnuPeMFLrkpp9X9zu8T/QaIKRfIEIejY
QDXThnm9O6BOi25voCet3ZVi64VMxtuHaKgcrh7QALEI0jAEi5lzjuBqvVyjfJnU
sPTSgEfq8exZIs8ODxxtLBJAc9MRf4RnSzdzU3lRTF2IC284DufH4UNxvK3uAlno
+CF4W/V2sUeGU7SS3Ikte8GQXlungrwawVs74lLHdyUsRArJ0ddS3QTFaa6AmpX3
2l4nGQUoc1MSvqaq6889S96XEhi4wGrQFoBG7xGZFlIlN7GtS7px/+SHQS6OIiFQ
RQCT9XU8Z/TkOb0ACyH9d1OR9FX4HebKEPvZrCOALKzAxxfMyNx1uaj/TK/aC5Ak
A3rXBw162U0BI4Y6CgHV0xAdvX/rX0lY7IHpNQyI8Zx92jD9nza1wvjJW5G0ovHt
WM1mcRnNzSJzYJeHvvj5hAhB5jtqoYRPZc7poExTnAtsE24+ygWtKmDxGycUfKth
Ed8JIhdJiAlu70l327dEehukeN0hVVgUhWjm8wKMPRV2u6yhUE5lRrGM38Qe1lFi
9pja1Dq90ay6ua71S2qspwSLvDAT8pz0jIM63DnSkBKwqfV9376+KrFDYnr2Mf5U
DANvZLh5qPuI9Az+vV/mkdbpM6RNpoBeM2eBHF50Jnzhjdkfgkxfk9eEmqyDlRz/
7n08PEwf5A9VFUMFmtWsJ6pHCBoq9i3wVj4batX2I83w/CYaOErpu1+Lyc9ZP2+V
86INaidaqCwYqd7Z53W0saMBIYo9Zr4Vv0jKXZCDQn06yPTG04f/bwdkYVVfZaMa
mxYR/MynUq++d9yPzRRffRTr5VwYS/ZrzBBZnGB7JgQO/CAsOvKw4NfUwODXWHD0
3FCshGu6rk90XlE6R6B/eIcM2N5xlMO78/KUgItncUDRpk65ovUNKSY9Cj++QV3R
qTiRPE6T3NlKZlNNPJpQo2DsW1PKR71uimLVVY24T73TI7U3xJI+i0Mob2m82rAu
Gpfbe2gVFEFYOR7MfWg/uLEC3BJbktRSCNwxFE2ldShd0Xbb1uPFtPqPRrysWMO4
EpyV9Nn3nr+oB/2Zkf8AMN83SEazlkOHBWGbOCl9RXSY1vUkFhAfc9ol+atTlprJ
Tu/MsNDlulhjSH/wFb/0X6jyUQJH9hzH6keWPo2kWoAvCbW8doJuC2FKQaaEQiP0
niCV2IVvrAondrZvHCw5WPKFj8s1uDht0wPv5i5agpFcenivm6ELmVD/TVSI/Xjy
lBIMukbCF1cD+2ra2ihmZtQTQ++n9xpQhpplRJYhFUJVrKuSQ82zhJKiotUVS2wz
T4Vezc+rY8iESGSf2SObTX69VqZNSy848UO2NRa+6ezFsvKIGkU4ZuhFp5pDJijI
3qLFbYbx37uNHnAWAps5XwLrIyxHqlnxlMiWjs+Vm5WVJLKWQ9JptdhbqYoe63QQ
sK/k8KfmZBOGE2uCiz/yMWnlm2gHN1WDIdnmpgmxb9lz0zJEdbcB5NfIsbbxxqwg
262ig8cqdDPtjSoE7Gno4WQV35MMJmBQwb94h+rj57RBSDbBb2H4zJC1iDxKJsNw
XDs7WT2ZSNe7rPc929wkeEzKf387F8ic2sUYZxf3yqZutHyWsUJ5yl2e8Fa+xLsD
eKRWOPl1hhVtkPSfeeqRZohByr0swLqwAkk7Soxl0jtlNwk1TTgIpudPElgsPCSa
DydYNTQgs/ANQqr0/SAPz/vlf9MK/VelEQM2Bnj5x7HDR/nhxYzgptqCatALGy4u
PDP6mXi9MQkiadPfyAPvddz8c2LJ6AMxtu9T0uLzDiPsKuO9ogBjMEW0E0B4j7/U
OSkEn4VP3mPUzSzetBOsyi6gHhS8lyKnSaxl5EPf2lzKF4Cp/MIhzSuoWa1IEeiE
bJvR1drbLOHPuDoahFFGD3vFxF0jum6JYmNXgOz+XzXrywKXcPNHDyIOhUmQqSZ7
r2K02j6J6/d4pd8W/Q16HZLFl04L5wuLC3fpEHtPY3pHF4MZ68VjrXDoIhBi1kxC
Q4naXvd6CiFrJnG+or1ay+Nm/04uyK69YOtdMj6RkBmvTE9TOsNYNQg0bKVV4ZHY
6rW0OZqR6MK1XBD7DrBqQlhJGIRyWmxuUTqlbjy4mH7tQMgvTCfu99zlF8NdDuOq
FlSv9NNbHzn0rWo8HGifn0lmviszs7nPayEsGuPxC0HkR7xHCyBQotIeVpD8OsXF
Hve49+k8Aft80U6vcgpqW57q12jNHo8MsskuLbJ6ARor3sZnlMMgsnejTgMk/9Ig
jPGYHdFqI9UX/HW2GAIkWhpawWvsTT5S6yETmMMX55vdK7Suj5zairBdNiqFxf71
D+Gj5UYvC7gMZg0CywiJc6gfc8Conj6h+DCi4n/YvnEAs/cVVI9qJwj81skr1y5d
XQe/rDPwtI3WpX0NBR23Et6d0anmUQj0MB/Z0Yiw3PvHUa5w99JuvwoTv4H5NeI2
6UQP7po2sR0zxNFzWLqaM0eR7XytCT73YJHd9jsuPxhtvR6AyO9zBVpsowTMitvd
Os7bhPAn3reJYdeWtvYFU/yzGUXzh8QMluulG1irXccC/zL2KPR5ZgJn3LvmtL/6
HPrUhlsQjqhDQTB1pkSRaa9I2rajwgZFtUKGrhfzWt+844juZyTLOhM7WidgZFWq
pelVgpEtHlD1w/XzVDXDT9dVSOCPTRYZfTMd8/Kjn3tRwghEPZaASLLI7ORno2gX
YOBSuQ/x/p4lwuXYR4PXJR5wzyZAr58PCdV2WissIA6/1Yxk5gTCOxdpoeMcsIDt
MWi3FYSaV5kcg2Z8hLgFWOdDrSstZeiLOWuOj3w5Vc2+AUUyTkJrX5PWJ4RMyMx/
l36DVX6VtbuKePQW5+GYmWNivgSSFGg0h2Lz+2yvsNhKGbCTNgCwbbh3VOD0tAYU
dVo+NSR2A4e22p1Ar+/L9Rhu5qAZVUMBIniCFSOrYJkVKjDdFR/7dyHUFJUGoODH
W729Hvw8ws6kadsubU5/cJWR8fOzk6oB3aqnUMRLzI6LeQhwHDD18XB49kOQMR09
YVtflGN2x1nSlJcQSgSA0WyJiIkRb4871YpMa3J3WA8RFqpT+Q0RGBs3FCbyKyEa
4UjE6V6V/4F9EptiKz0YJVl7ypgixXkusgCiaebiVtJRB06BEtEeKgwIClq4FxAX
b3HOOP7uFZhjJS75/gGEJXReog/r44SQoOKc6E1LsuOPXqlj7FjEfxELN3vFPIFz
D8QZSYgIRRPNVRo8OHPgpY492vpSCHXuCklIqDf7AIrQMISurch4TCNlKf2HKpii
/6wuh63I0qEO/+XMje37+7zkc39sS7C/jQhbbjcgy7Pl6I/eg58/zAFJekkYo29d
uwYguhb2F5ONAWwaBFU3TIlEC1I0sqsDnoB7L3qy2i4wgYL1DOMDjRusjSFovpnq
yGjaUaf+KxxGETYZq2yKAZmNeVPTX36D0dWX3vJLPUFLnAjnuPUzUKE0z0lWT7OX
r7ewp4D2mpnXa6ZmzcspFkUb2OJdU7mJnYBMyV1ghnkg/I6vBxWqWarsCH5ad7FN
bN0qSoXE68fdndCGQwKzQL0rW8mCfxMUE2/R+1U2ZMwjyXLNdhRHQA3sX73yJucz
u8J1kg7bEWImXR4SwDAHyJb2niFiNDhCSLuMuVVhF98JPFUwQ/uDpnM7A6ZUZQ7h
EvEV4/AxtwCMTLu5yhEcgrT1aWna+f31A9M5r21Zvr0fIQeT68xoQ06ln05JTOLc
NgguLSGVomN7RvJEys6o/lC0KNGSCS3q3/PIFKPreoJoHbz5sipXQjo9NjeieeX1
brqQD/+B/ZTQGb8eVxj1GK+IsJjVwuXUQOJsIHa7ystw+FapKGrN42Fp8F0Evial
Tv/1t7N3uYOMaXBBL/Me++KHyLlErmPucIVP7hnF3o2LFCajFzRSRI2lU4lVWhtC
MEF2xR93PMp95nHMmfw4/UE4PyOOeUGs5mt6seW+0B0q+032RKLJN/ZukYI+J9d4
z/cR+0UM2xEFpjACIQGNCpJwoGNw7NJak87Eu+w0P64FeWRXKsG4Nh87AKlcu3BF
DZClsJkIvdGxkbyV1EP2UKGdAT2SNKWI0377QXsO647zLxosL1YcIdD7WazhumvV
TRpIn3M4egR4YlFneBaYKiHHMcQsbi5E0Mncf8EGn8jOgjosmemIJJyIP4nFhrn0
V5PzhRZ+6SL+9bpKg4HABPQjTeHQwNgm9tbaAFbPk+BqgJrqbwkni92h3C0UuyD0
GOlxQ2ga3nL9izReBHVKLd1fSgJ5LM6mQAWTxNKzsFqMDRR0i3+rbqJ6vWrCZMyO
YE13RZTPOqBkWdoFiINa46GsBkVT6Kl5ZieOr/ttneUuMS0z9mpiTNXByOZWUG+q
v8nNwMTXYXotTaKVzPR8yEQftOIOILTAkaxIrMPQe5oNLboAC9k6/XwNYF+DsQMn
Sgl5bpH/XIQt5Zz57YnDF3zudVcnN3in/jQIUdPTk1ytDUYgiYesf3Kcf2Vm4VA1
B4d0tBiwEv4mw4PqDBWeZpTkBoQYk+HmH/NSL4UYNRmm4SnJ+ONavT4AvT+HwFuH
hOl39fKBihOIAfG7k3OsMUAbYTbo5e71s+SjjSzzsew6Jr6TvQT2Qs05bPuiuZW6
VfueiM/7bLKwU0dNn2hP2lpynXSM1P0rBVydY+u+WH1Gi9uDgwCYzLPo8GVPkYgD
N+014RKaMVLZH1bOPthUk/5eHcVp+tnztLmECetxF6mhrobhBlYxR6dlcOJcIcIZ
nCWztSQSFKCApLGZb81p+V/ihR8C6zWtgoh27bc8Sh+7Ko+9eVzmYG6SnGn+2Bin
n7gsT0QeShbdD8ubmLXLlLl/nPWY65WrLa+IW05P2l0ytI4EwIfjyB4wCoF4YHTC
8Z0JcZk8mOwpBnA4FH6PwwfLRUqvF0AivV2SgFQ4OnMy+19ra7iNLSTw1/LYDFGJ
KitoOhGiZpjD8UYzC4UE/DlQqWbMB9POIul52jjhEa96e1fct61uxQEzFXrJXkFn
lLx+GICox1xuKjzhP9PdM2C5zi90pOfqIHydxwT3BExffpe+0qapaGMzW1zGbIX9
w36UuePFY4JueYPBr8psOHBWuMtMdWhA9Lvp42TwFT9HBoB2rHtuj5K0KiKzhOXQ
Fwds/XyeDfDD6ajYeSQj8CKdNrSYTlznv1UEPqpzTajN120feb0diKlEvAnU8rdQ
/Nl5AZ7IQOnfTGsvjQuhjuF8b97ccCB4YqdUpAgdEB5UcsBGN5rglrudIkw2mym5
MKlipSnSm518B8L5DVbqdvhagVH4l+lwy2tD4DIyUpWnohtCQFlFxikOwlwM5S74
DkgJj9qQy+CfgArA6gAKRNGkSqlEVIcKkMTIKHPmDC5HzkZ8AttQ0mLIS9qRD1v0
r/BznF+490Kly0XRTmUS3mH8PQHuU5FuCNUcSAGvm0wQiUUAAqDzcpSyKWfMDWg+
tP3ZLHIevL+EdxdPfnpHn+gJCAdleUHUTDoTv6LbCqCYTtJN99i7i10FudVdtX/V
R5CmWAHh1uMLseJFWcuFgCKfg7foErbzHH14PysYoA2Lpza9rtbWg6JgZtMGJA6q
PUsz8IrhTZ46TROEqykeR9l/j561CDzJrTDsxtgyvIYPn/L3QyIGIMK62wbCVk8T
tdmgXBaVaXrwlyf4OfTHIZb2QE+pAhZeaayoVaX7Bzqx6W+BJlYxQQWnDq4ioQz7
e2YcCLWf6xrhE3LusHjQgw/XHiN6PHZBCDDTmPY4AnrCuuqsUNwQXdTzdLzZQOFK
EmFmdiFLnPywp6OSpRHrfQSTdcodtE5Zf8frf6hlGeIBQcWsd8eGfSgMlquRpv1p
tDi4yDvVRNaiiTtcvh7T6/QB8+AVaX/iTAf4lMppGp0HuLhOusvI6XD5Rg/pKL1P
+7bF28WIpdwXtmxok3y1EJ1DXZ8sOTzwIpJRLNLgyDbc3SbLhKgWABqaoWoin35B
mBckedV/+JpZypXVogFRTKaKWEpUyPRLeee5KsOnZYuiL2HMi3MYoJB4YNfQGgTE
NQkoHhyJ9LOFkxvEuUdlkCP0avMyY1v+b605dAnq5OunxF//9wV9zTG7jv+0GHSF
gLoyoCqxwuKevXN5ln13lgKCmQK9ADvY5C60GJ+8211FoqAR96P2t/UlOmJg6oVa
Q7SBGjT1frBXMFqEEsJbbnGmVq/3OBZ8Vi74rKVrGxFSYfLPsLReIzBwnfaTINwP
fV+edmpN+aKOIOvO05bIVSzaoxK48lvYuH7r9UBeLtbFgIaG81oDbnmPtOZ2ALC4
ZjZPRfvFWcLx2uhd/ngK+szvdLZ7Sy328SyqRmBJIU9gd3Ag3IpJQuSMU56Oqxtv
/uUgDBMmckbKpnkfbmYlt5SbExSg6UQ+lP09X1t+MWM2PtXejzQwjGSCH8f8pvW3
17V7/seaA5COI77GdJCwF4VIsGTxkaSVUgo5XHR6IvkvKRB6h5xTFlEQG68gjD56
qw+u7ehVzjXQQovT/+pVloAlqSEjn05lHFrmbvRT20vP0GSwIeXx0o90Liat2x5U
9Kshj1yEzAF18AYMIx8f22dWgCh6NerHKgVrPE7q5gEPNzhjv+P6t1vARUfbaUPy
BTGrc1TiBUeqAASBeiYMXQk0b2pEbimwNlH1reIMrTtOyBmcLZQVjhL8oV+86XX8
oYosB5JAq7NmsQ4Uyel2Kn7rFvX+BdXLlqVpbsmKm6t5sMuGIctLsfMoFaI7zs/C
IJKZhaiJtlWxEx72qNDqhUNAyGwrjhcYaZPNJUrMUbbXeUl5KaT10Ny+QfQWcJaJ
j2yOngIkOvLs5goJtURO7YNMjIVyuBjD4z2pIsM/4SpRWoKKPi8Z+SwRNmc84228
+tswujkLIt3UcooNTetdk7/adk2ZAjaY03jt3v3zGz79MRQ559qKTnjaPf60LWqc
PnjGsIXha+DDI3G52U/CUPgTcVPo0hcq90RWH0mQrpbfBPi6q1wTGPU3Y6qpava/
7LwcUSIBVWLTkqLZ8JIkncUJjZTe2Ln/3Af7GU65SKyp1jUpvQXQfw7gii+Yd1Jd
hegbB2XtCIu3sHw7DVqw34NFZ7eflBVOi+fe5E8X/NP0ng9vGPLU0odgr8A4HRmY
FRa98ggJ2cj3k9P578+la1SEPBE4ZG42zWfmVxR8Y0MA1P0X9NyqK0W6XSfzn/05
vdDM3C5iei6culFqoPiarmuazkh+AmNqavCZE1IoQspqwyVgTDWInaFvy9/Aawpz
8VMOa6OPqYVrub4PxuT9oUKYDmCSFlbRS3SDiwYrEeZEpAH0GQZ+7HMg2MmyifI7
KOVaOXkJGjqmMgQVgWbJxyhYYhQdKUOIvJ9Ek5x6qBNoCeEzz0jfAYODEQ/LCpF9
2FFm3iNOQJfzeO/1Wy77McQniXNMMvk+ILdTgeP6m47yRu045u9F/mFzybt4gpZL
Z7R7IxgiJ9xf7wqriyakvELQF4n/CMWGDkoHo/W2OlZsR1OHjc4fKkyvFMZSWJgu
gmWX1dNKNIYnCY8IqQP+0SYtqLnOD3LunljmhS2SUvFnUauGR+3v0lgXrl9duuPL
/QK5p8PMVdkJbxnKkHjWFcltYcoNHff274ZpdXkY0QaMMWSkCgiPI91qgy5aLjjp
r/fYTCwC5Sz0rA9ONh7ZPaqQsqdm15+OeulDu5A9oqqyex2wmjYjQOzVc2ch54eM
QDZ6W8KPGcYkKAuST1H0RwvxYmz7QbqIQexAp7aA1+S9BPB44OfXv8KS1mB2L97j
J1ONCfmHYBRIGr45q3NQ5aw3jYcl1vjKEef9rwy6dav/MveLZVeCcHblVDRwS59k
udGJUQU9iQhWmYFIXBDjrasADWMIsbEfxAqzinghokho/lVyHhJjZIizKkiPiv8x
HpcBcM64+TZTUfOed/HhScGx6zz07hmLM1+78S5pwx1fnicyLO0GNdLScMmXSse8
c9068pWua+Yywt4YAQdlgYn5m6ytpVetbiUDSTaq07ZwYg5i1FfoO9TuS7qh7Obd
SY6v/FBGvdt4l+CfNX0loOEZUWSpcPU7qEnpdDJhlGThD8o4GeCfx0Y2PEHy6JUS
qlW6KZSWKIHIHBCPbHd/k5C958bnFEWJ9afPuGQz2WBGNtoAwcmWbjzo2OofcO7P
U4tgip71dvoJ2s2XSQELZ8+TwMgN/8JnjJ+KKO9oqfkPO8hI0SXXNryuO1nYcQmy
MrROQoXhctH0cZ8yPEMV86AHUfWkOUC24xfsw7u0YRgULyKcyC+eLuYc5Q5Mma1+
t5LPSMsHQaaf3Dc3+Gq3T6FgQ4urYwBFBhxMBz11nhx+b+AS9MAHkOosDXBCwYVa
73AsgkI2oSUoMf3a+Ix6r3p08qJvwFoim2MYBeEu5vvPHcsba6aD/IPCTWbKStMe
9mWT50To95mzgJn5bY+WdPFJvOFRrrXN5g4jndd1c39nM3M+XXx65JVue5SRPl0/
i+KcOj34pLOcwCGvvoPnPxGMJ91ouD7+UAPqp9m+8Oavb+EBeOgUoKIbFytN9fQS
926o3vc6aNYSuWHhEVyGDcOmkcgUYjtJLQLhV69YzcZ7vEtp0ksy1dS9BkKUBBiX
uZsMXyE5G/NluUMKjX+jNQ0fjFvpDVt4bmcreXOZlH+RaOHVJ6457osH+dclQEHA
L2pDzdSFGIsiKRUAuqTjxtRwOzb0dbjS6jfxsb4t0GPsq6LT8EOR71Eq/XXUwv1u
TKNIe0q/nWppR+WEBSPCzEeSVBe8yvqXeE3f83GP8lXPsEAjMWeNshi+EiXpiZTs
eUzgE42djjNLPfHu6csIt4QgyLsgLjidJf6TQSgkA25agrBweFzeOrHYpNJ8jp7w
w+Jn+BpyXVd8Lme1K0eVAWxgmI10yuj4HF/kyMrE9rxYe5jOvKDHdeG7nWNKzpaQ
pa1ymnhZjd8XC7h6VkYi1GjVOK4RjR9SNU/8McvggpgvHMFwM5B9VPCBsIymrcR2
7jqT9fH9EwMv8+Bx8rF15d7LYeRtmYtArcuyWy5k1g7ZtINk8lrW7Feecq1BQfUY
W36Pz7iv+9dTHPfVTeMNFX8tonZ29X7wlXdOcRnXN44JKju3M5qid348+JFT51Q+
PoRy2CJmbKV/iKixGC3XnqUFFG6AzhoHp33lyHrzLSNVGvezRc62gfm97HIyHdvr
3TwSnt/zVPqoNJyrEQeme36Xzi5WSsQljEhRu0F4BWuv84pAvsApifAqyqQNxXBx
QDdFl99cfUPurqZ1GQo1jS5euyKkj2WgpdqG1SM7pq0eUEoddSv/yt1qgQkTGqPn
KOQYRF1P9q5A2VQ9THNnMuR73H7eb70kxCIZd3ALJ/RUmuBYuUVCrhlI5Bx6sZ+W
USRw65i+CWG4Gvvq4jb5LGg6IhInAOve9Rp5NHSUjvF6fcp4c+l3CqrRtgGSXnzw
hfKN0Y92eZx0WjX/E/AhW7dolO8YpROtfwS8du9zaECMdg5FvPBvW3PAaqW9sGQc
h7Sb9ZmjxYdVc6NIzHFA99N2c93tnXqZolRgrdHgcgMc2aw7SPDjoQTzLp7pSMHE
jVdMDAs5pXDDfzyVdFVcJXBHdY+bnK3xm/16E9fE+UVNwfNFA71pSuBYOTVBT589
HvcNtkK2ZK1vOxEuaLa9oJSinFJlKFKmxEPvmhH+rehBrfZMmxwaMP8I8uRibrfF
LlpO1SJxncI2pMYmtGkLJtAEZ7HZYTRaE72JUX/PHFnVO4pOlSkAGyIMEIfeDXqt
9EBDiWIq4RcPSpuEFvkzrJ9mOxtRcPH/stgBCWkadL2CeNH1iDOZvy9vqE7UhCUi
jMW2rL5nQzWSNaHM7Vcznt+ER6iwiEyYdrMi+zK8RAd9ccC388OBR9kLuuxF1sq4
XW9hTQEjS/6WDL11nYHbNLBDw7rzUD30Cd5DNvyYfayiKymU4aPOp9ATqkwcYN1C
mlX95RF+gb2YWQkWRsD5j0//dmrjskg8AEI7wOf5D2Ff6edczAiRe+uDuAXKkB9U
pNsm5uRjBt84etMhv6ARB1kpYXE2NsQdPM1KDuC/NDQ0p67Yd0JEzGRaFfoZeM6X
R7JaBR7KyMttrmagbDT27vtNU6XEaO1hiMj+lmUoX6ZLL2/acLv4C41tL82FrOEm
9KfouukjlpIzMNTtEMUEemfK1NftnUz/Mws8V3Qd949B0t+geBA6Y/WbKbJRsZiy
zOWY4FxQqOgo+e/1x7tozaxpZejTVkpdKAKjyHok9oYuMmdmqratcMSJwI6FT1PG
Wo6/GrKW2UZb8G89p8yryqKpw9zR/7IGlceNvCYEZnF+bXDsqaGZLKD++kh2oTNe
dHFs1GDB7ouni7Nsb+I05+4S4CEEaHZTsWe6Hc+4b9m/SJ2UIaM7Adlhl4aRoIMw
k4ek+1+KjEGJUqEHbJSjpY0CdUmVcSPoNIb/bNhMnnuOwRkl2SyWr2HtvH3+/C79
8I5OyItvKW2MBvmUzD1JkduPLqVdhJBg6a7RzP3KZjWlWxbuedfTmeFk+Q2WcvIX
YV7m/qWq0z7IXx+WE0VHSZ6rEV7MsoZj/f1XgYfp0a/cF5Es2zyi5tHuRRKsNOeo
UIIoVZTanAuS5ALGKNuVUmRUypo7aviiROWYrkzF8zbU3WZu1a69U6y8r9gnGLq2
XEImp+qXgPzoCe+m3lQ/sT1UiMPGRQavLQkFvG/1u8N5a//ETTmSPr7kHz9dNO2x
rCRwPg0La0QCElHV0hfIk/OaDwwa/5st0KiiTudzyyb4QwHxhQO4ChOJ3SlmkyGH
WMQVSObiY+B67XqEVkCbUgpGtLpdLRWtmOBZjliFpkqvZ0mLcqXO9HXuORJn5HXm
R1w28JCVURwzpgQokLD+Ip6fgqwOCYUlfAzi4k0fa5cxdvv/Wh+V+KvfcI6tPzlH
vtfrZLPwLEzV/FcIIlNJerPopJqaQ/A6GtONdhFYWgL5aHu0LD1pQEe1A18cuMku
2wXgoWiWjGrxmRa/jREoni9XWa6aerIpr1Qfw+jhwmYPQyOe1Qo0jwkiYJJS7bMb
wOP1wQVI2C1ZMpjGSW0dysG/ZtWO/DAZF0V5i72FhLxDax4vxcBR7uUVu7stwlqZ
9WTTRKNNhWh4C/LrvgYgSqylrq4CQxtlm8oHcl51qMyHulWb6wQzM6dAJiBBsOHM
W7nY4tJpeZMSHbtnX9k3WiTUmguDBbkp/OHYdxAu/sXVjaEUDg2OLI1iXoH2+sFB
DoUNexuTXMM0nJQXL9V15nHAHfc91Xtx1EPM/5p4j/GDdY5KpP6gmbuGugqUW8fR
q0HHXtWmfy0dSzxP9idiJB1LLwFL/kNrhdLLb9KPnGZa20Gfhv4dxH5nInwQigNZ
vOrkCrUyQeYI7iOc7FP6dhb5/oonjreB4uVsDB7BjLSSiawyv0lu67CE1vKRkhst
RjOWpmA/4yK6uR+k6AG2Glok3fA8wsWqhAS5Gc+w895JqZBmOPO8AASPucKld3dF
cszEZrAoR7eAxWCJU8ZTxNqFPRcDKaD+N9CVKHbXrpGKkgPgmINYkfMHrFNP6JBu
iMFIeRB/byISQEqNM2SPQfzJUw6ecCht2YKrGhga3m6CRzfHJ4ZlWiZxbUWlK3wY
UP7q8HoJWmlk7+wwE/BudTq9Jf5e9HMH9ZDogdC0r+v/uDgrn3BS99/coNTXnpqZ
B/EZWjWvOsIO/mJszH/KHtBpOb4MosGR36Zr7ddun2am8LxtOIt9yuzgwoTX03ws
77nfN0o0gJsut7IH+SwEz756LxRYZFbt6WdhLuZnIp+IG8mCCrtnvOhqU9NV1kM2
RQvfHsdGtDUbUKyrQN9+OIRD1PGOOBgEGCDyqI/oC2c40HGPS6LfblEQLpYSO48Z
rN6HwWMdvEwAokz5WBpndOXpoJ/KiB67qWaNtWwXk/GxAiVfr/mN/tpSzuBjug3k
Ge7k5I2rW8CgP1SitpVLAh2EFDWBe5ICJnXZ2g4IRiHn4UEV/tnBEpTWABHir+uK
7pAuxNoGUgImso2VcFJH4o61KPNHgyl9Scv516EkRM1EHtdj4YRbaVB9OOkrSgoc
KSHo7RoPQSbY5CM/rn/DcYlfYW5OccdmHqq3lqOKlaJQ078sVdoWgegzb1StljFL
GyYIpiP6X7bwrFy6MC07pd6I8fF9+WtvBJNGBnVVvl70xHbG5ZTYBu0ZNxy1hHVm
8fiSYPcvW0qzGlsLwntRejEMGbYX5kluZj7mNZmgxClrcgHs+CFjKbhc/NL7/fSd
eR81KMDwuakSoch98jMRwUlxOJlHCackErTnIUVLBW7Qa6WKhXZ9a14/3YtXqPdH
GdK8XQ7TriN6NXMnKTqn7GOuK53gpvwM9dAahzAa2BJF6mIzt9FqZ7GgCeghAiqS
+PIC5Iie3bPeNGh3Pu2U9CluvoTA7zmFf+JLCLoSBdTl/sBjmSJnv0tGZ2M5gtEj
VqpbiKEgHwvuvSME/Q6uvxufPojA+3DF9p5yKPv7Gm+jVFoVK828pKg/MaXwi1bQ
vmpHMPxnPxhMaA1I2hulJ7E50+OER6DKsXilPeqyb00pVz5hE46eHaQohLC4Uzaf
zNJIBNzAXIBXpdSI85bF/gIjfHlAy+CnMcrexOeGls5NYEEa0EQjBTRW4QwADk9f
iHK9skmWHCsnRoYQqv+wGwCs+zZwTnkA+UVtc/VelL9NVmLiVsgrfvZ6U+88BOdY
VrDeYCYj3lKuEsq8tueJzRrFdvOC92PXbi6IQhUGts3VW2qXt2pdBO/jCfmcY+CW
ynerKIyWnZ6DIszR7UcUy+QxD5+pKNd4HVY5IHupMx6MgHgU4iJtQA6/edyefmTU
kjCWXzhvnxSmVMU10U1GcW0w0kYZJRwXiR8kiPbJTu8mbUOU0998yh84y3SKjWVh
AJ1SrabGr2XugnKR0nL+mj+kcpMtCgB6bOOTuSZWJark3ZKSBs1n5aK7VAniDxPN
tP6a+IQsWs2TsENmEQKU6s4OJDuyNdsXCGLeSPHB7VHXaOmPKrCROG8SGwO8hDQE
MVOHwV+pFFV/LdU+5fW4e+Kt5s8F5DlpZkxApN5I+oCBW1w9zXUlkGPuraVR5Rwx
d8pQ7W6qT07rGl//VYfB+MtYUejOMFIT+oj6QUFmUxySEew0dZiayB45SE4lmmnc
KaWygFyie4gpegBhDmbhBQ2GL1YNYfNxCg3fnDX/8uf9wSauDT5RXSmxbxdBRULP
FoupByx+yS54IOeAX4Nr0OgIg91vME0B94tmfoOWZx97BhR3S4x5V2Wn59pAQ4wN
Klnrv6e8hX0nS7Cedcd2mK47d1iWhohAczqBfZqPy1nExLquPkcwODWwzoCwotBd
1WLxcCm1vkgL9388rZikG/+MYKD7VLfiylt0Iy/lM6u/CoiwgtmCP/T2c/K0iZ4p
IXIeJLGfzovBZ+XZ77C1b6uwe84gu05ee7lmjDpwQe+lDIAl2/4QKC4DZbHzYzfc
QEGmvvCBlNmgQTZBe1J/w3uw83G9t8+CnhFngD2pBdDCE8LADNDit5iPEW7eYLb0
+dKVRCop29dFkHrXdsl8M7Hqnt8M0H6C3YqGv9Ari6cTJPpFKHtoe3JpfcGGxWy5
GGO7OPkgC5srXhg8Z0K8p6yectbsa214c7NxQma8RGdhUHMP1K8p5sFbX/OGnPmk
oQOx+hWGwtE8usMZb7mxfBjM5dzuLYiC7rGkuzFBvL8vFuPrr29UwCRK7gJJe1fY
ObjOJC53PsI99EkPeS6c4RDbJseSLx524Qj5l5kp7xx7VbNMf2iOXbA3zer3tWfr
0wRpmjuPqQ/S/9V2daZXclilIyiLgsglMPztbrqOleuisZtRUF2yx5juGJopvh8W
DLybef5Qaown7+mNfgTomnspR3KG7S+W4x+ILs6aU/j3z8gcOtEuL3CWCvxxb51d
wEU0D2zZySP+hEJ0ux+ZU7jtIzkonixyjRMM4RM1XzrkIn6xPkO8IIVkcYcPTN9y
f6MmBsUuZbQE43y6H4mTmYA6w7lutgdZXjO46eex+yI0jB4LhyqAWp33fsoa0S2v
nK6pkcEtmmxBF+s12crVjxAHKD4jLT1NjyCL3SlHwVLqCGGhQMyO1HHx+JmblNFj
ZL3qf8YFVFz2ufQRFuR0eHRM/GFrSbPHlmKN+NR0UfPXOR45s+KalPFKyXTq9chu
50OIAkdiuXIuERh9PViiI5/nZMMIxYIWOxA8j2PGezN4h8kCkAZG/FcOgDy7ppmh
OAM/ebH3lISu20B+pe8X1AxHODW5vvBXry5i19UY4TTxKIVBDAUshkoANohnNwbV
WRsADHHJ9q9cbUtjQbnSL8PsO0yEtosS2vKu7fNEL64NV95+5BpAP257XPJotLCL
NqZTufLVPhZwKBEGVtplH82B542uu32lHFse9uwl71JIvZvh4HQSX9ews14abccE
yqJe96PaE+m+Eclg60uY53jHcxylkySDMjBfRicUqRgLFlCk6KVEGWd+NxBizDo9
vZ+eSG2PUz+iw6REaJJv1X+haRGYQt7BmgAnnT5C33mI6uo7+2RVxlTk0LodiW5r
8+j2JWPT/rdF4NQEMvAcO/lgBujEJkePjw1phAHzY8Biqgnhb+FhJEnTeiHK3bKY
dPKLZaUdqf1q2CllYACkZVPHdNKzE0CWlJ24XHXwgDm0p/aXGu9jy6Df/xOGf1Ri
LAoKs27LdLbp8Nqf2yeki49t3NmcQTx27IlefSdq99HQeUijTYbIrj1Lnqcz6Yq1
KuaO3P1+rVmAIoKXAD1z7jCCgRbvmrp+ZwKPuBPWwMHZLXA6Bu22CQYLap6OD0K5
hLbfhsxmpjH/hXpv+cGd9suzBJEtAbnvXDnPPB3CcG253czVZcxMDIYV0VhTP9o2
HjdZC/vblYiHEGUNcdcLxp2ZQygiOtYnEMT0UHtsCMYHyI91PP0pA2tt8M7lwy0I
EBAcMpNb49gvSUzDNYfLf549NPL/eQRGxEpz3bnbDpxK4158Uu/QMCPhMFjrXDCr
U8PRZ16PKHfK46/b1qw1GWFKQLFg2p2zZH50pK6/rFpfPM6H/Xu6AbdUmB/M4LPm
yc9UQiDgzgeN/2lpWbfEPMV8gXs8YxwAAW4wHL48kp7z0wg47Rb31u0yeaTXzdk6
NrkuyWJqDqU18i2zwX7FnEDbG7CEv9kRsxVFg98q6IbkucbZEsRUtLmHSvuruz57
YqeCFaLsluLThjdytYrdVzvRf1PjqOZfPUJztDtDIhvjqnObkjdvP4Zwi6LAQdMB
20zqoM4/3Yhhh2kg/3HGGnlgZpwS3gNxkl3h+o9wNY2bRHn2fmbsHLX6FI5l9nOP
Kb4MiPd9zS61exRcnlbLTnsS/RqOJe8vMMdlb+MXyxefewF/GakfAB9lHflHSOha
qIdB6nE9LGoObtJtntjKdPCmcOWPcpQegy8Ztl8Byrm3uSWH5oGx7rEknI7r+5GQ
YuxqPvFX4X9g4DvAJbp8cVVsVnTsuradr6J1DUF+qnh+ftky7m95YI/O8/u8YMeq
nvS0SaZZE4+hINySLQxFnFodIiFG7HRPP3ha1I5yVe3WdT8q7zJeRCPRso40H3zY
7061JQ0Fa0JcAaiygsboA39YzM2LiPz07ZaObswPRHQBWBHE4vztIEgd6DWycgs8
ejiMDDr81v7IBheaQFcD7NZDr3KEgrVLkvrpTYRR05BcnDtAV1FPz+Y6SbEzOO8r
CWzOTI39uCC0T3mQXjsASoMRzV/uoaudSZqv/xv/l5lIwSpvvV1Xotod6C5aC1re
AM6wrJbNAu93B9Ca98e1ficyeMI+mo5J2Kpuo2hqgfsvm8p54U3QqtdrdoorFJXA
w1YJaj4pSwI5FN68A5I+0E5BWrJC+v4gISnXbt07htvS1Z7FfQ8rT0YUUKyDYAep
ZyDsqAA1+vjWLNIQg2L0ie+zVsBH04hnJ5lX2edaxfEhy/KzbeypESgPqo4+tRRw
E1E0HnrV13jQiM1UdWIzgTo/AadYQmL+Lcmc6G7vQKU5xf/6OuSGLpmaFlskvtin
CQTAwDjIJA5ny8Mt0Tz7Lgz+icihBnXKg55t0AXXkT+FTvpr7Z7kyTcs5PdxwCBw
/WG+k0riwxSNl0odA7nkzamYHKBsuVKkIDa9kvRA/qSOYt4BoewI0jbODMdGTwv0
fhQdy5a5DCvgkn4YtMWt3ri5aFM1e3vtt4yUFBh+DbPWlm0L+m6Jnys8IcTwEExB
vn4Yjc9bJA1ljLL3tbdlXQYZSu7kO6lTOonB9Fy5hfAKgVqMOhmM8b5BMtUcRSdo
DdjeXJwodfHMZ2IhBwLKqiSX9a5lnonPNsfX0VpNg6QHXHcEqwU63lSGu3px1MyP
zMkJ/cgpBIAevlOqCBfDfaDM7n06oDRx2pUI1RchfgnUgBnBqHC60ZvLtnFckauE
HDrUGlhtQ/tgt/m5PmjEJ7eud42W7B3csTNgOxATqKOkzy80T3mxFtTZLg6OCGzc
JAqPuzoY5iscUcnI/+/Tl6tR0o5ONlkVxydqE2OceBuMTcf22ll7xL3yg3jgDC9N
5/3HI+THQrOAEAqf2LZtC7kHCTTbzVKZkWghF69RKtwr/ymT/bV55V5bEnyNm6Mi
6NYJXUBKxv5C+ndYJfboCDAhDrUlQlhQ7LWNDV+oCMEoGVNnSBmawHfVB/uEqzQi
LM3fvK9UflgMdlM/GZorKWcWRC7tGf6s53vSi3O6WfG93zpV/baZxGwxLqMjaLaS
graEg+NHRJvkpPcWgVI/jkCYfVTOldZN+Rnp8zU2/Vm7v6LE0YzfXZgkqTC7PNWE
syEWHgZFMQnyqf5BcEA1pi0h75rTgp/xteFhlwqd8Wd8UwkRvhFAgZZ/kMSadymN
K7HAvzLhebd5fYtSmilLe+xE/oOg9EDHHvexv3HS1GGfNUX7Z2klO1QLq2lKjTlg
0MUWVrLwQleCTGQn8nzMCYgyoW5AAPOOWJaxYxYI+2l712dvU7bfBxVP8FL6TFiK
dBoDrVyl5B0Nk/fz7bBIuHfMt0HZNvmE9/GkewqP7C80bVM1pYQZ6C14OyoXDsuJ
3imdK10X/7Hu4Zzn6ucxeaQwzbkFR8rNPvFH692RK8iPuQ1OFulgULxypXCjv1yx
Y455y0aT+mO85NfHGyjXi6oNyGyzUHYOl4IFvRKRg8kbG4M2FZnappOSf8UxrdHa
wgmJhMw/Ya2Op2du8KYRHm7AfUGxWZ9HPSnN9WtW9NKNk3SfmbjlaMTzQGYZdVfO
450O17UyMAHuG02eWPAqUrGPp9zAPK3hfUU5I1RZawfgDKtw1K7Yz7bJ6LliNh1p
vyBNaCMPAUSuUsPjWubnuLaK3eb8Yb2i8mVv1mmrXXxn4au0Xa1U0R9TZyqDt3+x
fEknFrkMHihmFfFcbDvVue6ciIGhndx7d5BOr8C/U2kSdKyUg25rdnmWiCPZJfdc
S6iGtlfh4aKaAUb4R8XgLYtggjpx4VMyv5DsmUWO9ZCWMBiuI/l4p86xeNobc/HZ
LC8nZCNP/Ye6rn5zBlvSwHtCupRTH5PFCO/2ouadA+k8eFztkg/vED4rbC2zKnkX
ZQ3IdgcCVmlnFXYO98Ya8D877Jzs+gfZXlese59+RawGjk1teExykHBq9Pp5OFaa
KlXVd50gBdfPXlgxRrEI8aGl7sg2M8Jo8xg1sUQuNN9z9cIGVZAWXrrlLrX/pHfj
Sm15j7iUBpRwk2ieJKtPx9QP/gXi80NkFK9k7gAZ2xBOlTgo0lOnIM7sfeO+VLuB
17LAZznrbAyHlkd0ch7tyUsvO+KY3RuzQECj+f9qDijgWS2FjkNBnX33qRgjLIqa
8Zy4moU7Pkr3MOVM2xnVCRFCmyU2x2Haw4g1VaPqAdz0HIK8ErWwKNpSHOD0S3lR
jZs96sCqXKTd4CP1DVZ1721UkhvNSBmHDowTCttv0cA0/sRz+52zDGSnv0i/f4RF
BxKMb9Q/iL39hW1LZ9WX/L61JNJv2Vkkf2kqOKYJ/Y8RsAy6N8LICNvVw/+Bx0cR
zbuLP7Yo4+zd/qcakAbGtdniTr9TjXPcSKesj4kgNbzcOhpfZJEF60x9RcUAhrh+
w+JwkQTtRNtnR4qRGv0Lnb3cPzLS/eKllw5btrwLt2ZmPsFA6EEukt9KJQE8ZeMA
e/5kXdtjunPRXJNBgUn+2O/UOlaGmGDIHdBvH48IM25wJCFHNF2Zy1UrkuAUBXE2
dDVAzxn/vtd7e++dC2Sa+U3DQ4BpKKR7sI3xMSqwZ1BKfRSLGMHd4nE8OYLMc6i7
IiaNUuRq6OKdYH+2m2TtcsSCeeVzIFDLUQ8pZzkYvD4PmKuAYdTOoeiMZ9jTZaRR
CuHWzljBPHRCQygilS0ht2JNl7pXhEsuUF8B7QVHADYQd8+pIa1fCVS0diGf9j6b
gf7b341446xKkUmP3z7taZmFn5nN8RiIv4sKqTD9tIeND4jio3wvITNcFZokMWJk
njxAK5yN6pox0DrvEtrYAN3GXsnSk4YvKbjJq6LZbIJIdkrH6dmsfRvAdEh/fDV2
ig5teSGDqAm7AHQTCXBBI9JnaFHbcij9EwAzhMVIIqlh6he1psCLllVDAYJOT78K
MkmVoofZk2UXodx0txb/YCsl6+5Q3HoQbrem9mW2Bwd5F082mO8I1WhOBjuL/5be
J3b42xoUbQiGRpgPRNc4FCEOZjtV/sJ12oD2ByQAWg4ffX4HN9YpjeZsmg50yXGj
E7U8Wn4KG9WmwC89UsqmemmO2k62wW6P3JCpYnskNd6wHdUwI0Nib73nxw0AOnTT
ifPZVxV7qZEdo+LyCvrFpbKzuzT5Uu/hkwicG+l4K5LZRsZxdZh6k4XdhI8i+68C
I54DN75yHyDoKIimi62lAXmfxtTNDuM+QmoMlg0dA+EcFThk2gO2gBoiM1O/8j4y
WJVXzQW9llbw3is1/kBMLbhtaU1fL4L+l5DO4lNNDMVOSkOnqlB0zJaywpJOcbIH
4fmopaDAWC2VyhB/Z123RrF7XKaUSFZlWenn7OSnhyjiLj81xOF3U272fbupKSz7
kUWOajtOmVE+C5AIj9n1ULv+B6fkV8+TKg5Jyoc9h0EueQxseYU8BMiRXdBIYW+d
o8ECPWxrH4d4LFUIFd+1JE49Lf/++YzUUfrgDhtlun5X3r6XgyyFYIGrhPb5ZL7E
s6Bgl0HUgyku3zwngA8RwxBfAtbeaPtflHlAX/SNHa012Rd8Gi4nPIHPYIy9kyjJ
+9eOHb2ekex50O/5qRuAc7xtpvT7nF8vJNeWywYw2qgMsdGBS6FT0Us4PKqSY9TO
N+jWoPpXfg065ABCsZkxFj1ZXtOSiQS98b0XtIROO2Z0uAOx/izC+efbrs4OQ7Xq
4VtjPraSJfF/PZJCln7qGBSAnDccSYAB+NBMj5NwMXatkXG3tzQXZVa5Ueb45mIY
4SvbAzLi+QbEkrBffje9vyV7u6STm5rlPkzu8jqsqKztkCerzMyLQyoJRaDFclmg
s3RyEJaw/2DMl8o0FJoCVjZI4gAm/WKpwYPfnziX0uLieUZTHbAW1rk7IoMz7Li0
LhSmwKirmRAgQcAZ1ksGand9IiyPrhZIgxWKH4r1i4OoFwjxX7HfygrGPuW+whf3
pgz0FhKPzDcb4AsNIhy2hIKhKGdBWf6pkERVRYqq1sjN6+f9pGGz5XqercoBSUxK
zFHi7Br3OWERajTJuiQEt2rs/o6dvfvTtPp5FX7j+71GmjZdYBLz0gTJQlKa8sDa
33hhmS/qkFHFpgYLB+GHPCTU4K/kzSDSVpt+iVlV5cMFk5TKLM9o24aZZRHtkZ3H
sTDjxcGy0bsQA6J9gpbCpow3TZNiUfAPGwFJNJhQviAQdPx22TJBJUoknZ1+Ejkt
DLXNm5OHfcCWTUhMf+xG56T9RIDSI1Bx49G47PCA60+aMLOCelplPBddR6b9V3da
Ffih9zrk0G8njp0IErr2TwsXXoqAkYpvXBm03icZZFLz7yVeQXPcCrHyX42ztYOL
IS5GlSLrna4trv2hL+R8k6p4j63E/uCu5X4hvbDh5xz6r1Y6XAIlATpWss329xao
ziHWzw96DkxJ0pe1l45F/HAhxisU9DkNFvuOPCS+1XoBlDzi5EQXbOaylZIgS0WS
jkMCYqE/Mma+y0gCT9Hoglel/7dgA2c8PkeYnOd5xWT3NtZYNZ36gRLOagJVc9aM
81c0+ykgVEeNpE7IKu9+I7hTj/nFhYHA2aUaHrKRNwSlzKGsoB+EQ/3bY9cENats
DrXnsZvtADgOeUWtsmTT36ypJNhbCdrTZO5GNgzJm7prlHn9Oc83NPOF6WSxxwtm
hX74j0s8NYZz3GkwZj+rERtVknp6OorOpbiC9bdRN+Lsz2PDaMQG6yBjpJovg0Ty
3R70SVcvz6Os9+pUz6bIYoNvsRJXr2XlzXcdLR5+vs15cZYNPIE0HVevqnOMTwLZ
51Wre8X5wVbqROGu7k8mRWMgtrYOXmfTibd+MHnQuPu+puqoWkzwkAt6Uzi+FOE8
XGAv238ImrrJ44vsZTP8YBCPzBo0bAavuGya6xnZB+dHX+JUjCnYad3YFOLcIjE3
gsKwHrcub8LJKbtTND7jL++E75T8i2nycYhclinJoVfEfJ5spuI08WvOKpRD6vow
hMD+baCgKZXUYFPJGNpPjuIoLhGEleJLzX9UZl6dkmfBw7jo5Rk1VPzhs+74G71X
rJ7+7yIRYgJbVlGTg/c0YzWPwfZXXc260Tml2fetNuENOZwkENReh5zUGv5I7vO5
cA3KcOna3r7nBVjYA2idVEV2eBuVDygRvju6WE4alouNuF3yCJ0mJpJqkWY+o7oB
gWBKVoxMGkx9RA3aBGWphC8ukt54N9TzEDi3TD3Nrz/arVcbzevUFtMBmw9A/aGR
ioE2Y9hd26OnghwEABxk6U7oIex/rlUH+OG1yg27TAy1lBLFGisUldHnIoB779av
3CTv6nEMqbyNaWSIxJQI3q6+TFuEMXhGvWz4lT1MOX87H1gEhVOsJKxBmkYMCbAs
DMYIo/ZRl2cm8tI3K9WpJ3XL6goNS66W+ktnWqfNkL5AI3ZHdZlRIkWMa0w73GaF
8JhdJAU5fiJjF4UL8pV+HrZK6M1qeLuAnWamS3GM2eO17o38b0ytqKjqUtU4C6wI
+ID3Br0yeOO423wvyWEbF34jWoJ788call+qbhmOSzXzREf7hiGVFzX8gL8+NlLF
KPzI6TumTEGGXEw9S9TII/zBcKZ0K8GPTrwo25Tcpbs43NIdmZaDUyswlH+17CG6
YnKf1fMGI/jd9XRTf9sSCMpNgw7uZq6odIFHZAvwY7A1NkFRWPuryhbYBuQDsVl2
w6W5EU4fSlO3F8n+HhYHy332/6biJLX//C0+ZeDmSmYRcvBHApl0/T/PHRY9WM+E
uKl+W/O1menpa/uWC+9syeNq81oariiVpNseAkwRhAtJqVLNOwPhAPSwOCWK5lKU
t2xnT/cPKm/OeosUOzRes9dcY/tJuRBV5h6lP/ITN2DKC1dhiM4RqeoqQyZDqLjy
0vcO2UcZaGbhIDaLaWVYdWr1R+K8iXkv2b+bhYcj1MXbTfvFdf7jWlGO0jh4X2QV
5fzGBnxqd+7PRN3WWKs5WaX/avtM5kSWrtSKDkFRqf6w1AvkN7OPBLxNo8Nc8qdd
5IaqXQ/ifgQo6N3z1Maq0z++199lJ+QiD+EwH0Q+ro6uuNr2ooOx24zwDTWEwjmF
OrazXiw8rpsLdGxjSyZss7+Hq0xTqms/Qpu2eu0gXEnkdhdfexCuHtrLKTvdpfQi
pRrjZ/mDSUocqox2T7Ns7OA3k/5EcwcUqjqOTijjV1V1UgVtelhvvNcMP6HYu9Od
pYfWUzGs6cgzdUsfBxYFebxd+h1g59b4ZfXltQnw+vJyPrLFFF0apVPqf/c7B3Og
FJCn+HSjxKnZDhttVYc95FpXdaPk/SDn42Px5YM7qbpk+j44qhDq/apb7Z8LeC6X
8naWQLmItisoidpSGyUkYct2MGdu1E7F9DAtZ8qFQAQ9WM5UWJHYqrzY+x/NWVde
OQA0GYzkG85FlcSRMHf9HC3S4c5dcIz9GUW/TRgazkfIxSyaIaSt/JnJxtx0qpJg
EAtaQnXnjFTwngd4IBvn/yKE3NfAhdEW3TOt0CqwlkpoiNS6cr5EOPV61TuqsDQU
1zEU0/DBbnCLucriK7RR6NutDI4fCVdR+S8dHxSHWVID6Dn4luUlL0k3El6Rk52u
IaAZ5Px7Pspq21S7q6r1oH3LgUuV0Q/x5EiOqu1WWOHLcIpS9QM5PNowYYkFbHWq
s/1CJlfgBjGWGrXPP3DQQQTRlyoe/Hnda76l1uiuZZJZLxVBKuXr0F3ur1XvTael
0KEKjkMNV8ZY/OcqWP2Ptnt+swG2WsKqhS/xzsUAue6OTwbJJ50aq8m6RIXLU/Q8
QM0XxUE5Sq9dyOgDX+qK10QE8OpLXAiEfEiZht8sO0gYHqrAsjiqc9j0MdQcyoqe
OPfth1onTepnVccrhwYbzAG1x6YKVaiqk0pBHgo4Jfn7a40kn/t4A1UVqaEtMDF3
P46koBROmyimm/fR7CVxUyo2xs15ErLFMXw0H3mO/bbarxGX9bUslrXut/p4FfX4
DuPjKGBctTlUM7ph6GvQyq2p+r61B6GgHNM0ZqKdsmuauHn7tdEh7bwT7wddLIe+
C+v1nE4cEZenhi2V8KzqmHoj+c6QONVnTfNsl6B0Yrw/szZ8bLEVoZkayiMvZrFP
oS+WdpHTZDBOg1j1mHpZtlgCN509gFk6Nbq2rrFPgRz6ncm9dfwBXTJ8Fmn8bp5V
xCuGbT09JhM3aRFyv+a71FS4jExdiQy5KbRXqt52oVRPjL668tErEkhrFdMCyQE/
nYRVMTArLL66wiC2BwWe2O9u2u7Ml9AzAv4Q4FyA01CK+Ru7BaAi5bMsxWsyah0V
C2EZxrjrXVlLzjq1nv/7jsfVj5QALhJ8HNpmqKGOWxgVIqINhOBYjChyvlf3yTx/
x7lMN7EL2shBWoCNObIhZLFTKh1fSsN46zziC6foVjeM4+abrM7s86tSaj/F7yvx
MMlwXWsaNi1kCvF3QEU3SLqi1AS3bPp6VIMYcZFWAH6iAVTj89Y3dlA3i7ZGTcDS
rixmMPf7EwRiACc1GZzMNp5bb3T+p7VChXor9+x5F1pCG4edM/uFaEtMC6bsiK94
bferWKxbHLCm6hl3p+6qAxL1G37aAFsNboNoCJLMZbT6ZhA/RG7CJl0Wzovx2uSS
AZjRgFzY6iGqkpEEOjKQVc6epADPtQZU7yLpDe06fwgXwC7X9S20fMh8K0OpsrJN
HxnOdtTYsKz3OYtwsb6p3EhT4Rrlg+2Zp0JLt9yH65Pw57qe8Cxo+8vYpLBjtNe0
SHQrOMw+0ycJ/0l2eSvxF8Sn2082uSv8PqvCqma2pt/jdf/Ui7iCt5NnWLY6u88y
zMUSpVZHDroESZfbTecjq3NTCXCNrM3c7S4GJV41DbSoIh4C7OnfoZ2jyuLVLxqh
zbHhEsANVKg6+S72s6hBuITJ2Sh5WkloAro1T4SaKtNgFZrdKivzQIiJViWo12wA
s33ywWzAKQCIhlWMpJ8ZC9TwbydMJGgv8JCBxHOVqQAJCPHxvYXYTCV4A9yxs33c
2QDYulP0hE2Vik6ag30RfARfLmPkn303fomqX38WxcwGizs5VLWZSw3RxssjjkI7
R0N46ddKhcxuRp4gzJSJKRBdM/4JdjVCUWXQUPG4WMgbK0Szpwhtw94EcaY1L6e7
geTZMxGM+33nvMEhh89OQixTkChtuRELWdAH+FqEPw2xf2nd2zAmnvGz9XB0GR+E
u2w1vecosVDtm4z4Mddw4l0SY0yzhvfMFdRRoGbVUWsJp/2LBOieBCh7FKyCyy2e
CehPMHyitxyxamK4ilHJcbMjaI4kx0Fs5cuHsuWnbXmieok0zYsNS7cR1trIbONA
LtwL7drrK+nGoGUkCeRqTrrga632pdMkdYtNnPq3z4WdwtII2QDZQsY25ntHv3hx
DlaretHMAbTnKybSp+ldLAPpnD2GSeNpn5BcN2VLY6/JgwG4FFLXZzf3ckv8YTOw
b0bumZr3riAuaMtum+Fg23REPztCrHQq2+8cusnjkhje/3XElNsFd/yEN2LfR4/b
MNtm1r+C4Sm4ZntbMsFpsEDWRJFUU68BoTErD8CWMsoQlJljPXjFG1v6tH1MbjXo
RN3YQrtB0kB6tvL5fwzH1ZtVAs/9f4iVGdQ3w0S/SrKQE+12V4Dtcl58DwPDRM/l
A2GHmee4Rb4wvLE/sSDJPD+cWS5yDdpLYnCV9NveyiNtJnOodRIZ/7DV+XHddvE+
sZHl1yoJNjIfYFIkzVYelnIrdDj0kfSsAm2eSS1N8OWYfKH6jMvQGGi8yVC6xnhV
pL5CZkuvUMMQ5xa9oLQmM8pQTR/Cgz5WsVOorMZvqBQz554Dc5zt/7RZDlayGjkK
aoXyI6i3Vd0SUlulvZnmVr/YVuRu3+1lTs03Cr7KngAzdRR5baRt4Fsf9rDNixkn
3l+B6YDfYqzlMsekEAPVVbLH8Es/ntXr2cX8gWWMXSmVlaTrym/H5xxoc8MRdWxF
1b22PT0V0qHxSnvtKLMXxWNBsOlkDknPKd0BQlfkwzrF07tl1yzbwt0uI9wskOSC
PZTVYMJ8BAkwR/7eULg6VoACJRLZkzB3b39ouQZI60PtbsWgw5lvDv3Ho5HH+7vw
dqLKVh3qs1QZ2TnYqipOwkEQAnkoDGeJ0ebprBm0sh6QSBnwtzcneFkkSnSRfhVF
qurw8i6MbBuMOLcTjFIMXnTe1lXYYb4JymKHTLrO0bDlb3WLQD6y7f1EYbVWv66C
N4CfQRf//0kRyxm34j6eyDHgedsR19kqTy6e7/mfsJwobzxAlQm/kqAdiBtLNCXW
2/lcofJYLEFza4A6hRwNKItJTNbqOeX1rXYBLEkhoLgL78b/6M4/lbxNHE0YPs6N
LSxIMR+JA4x2Ma3LVtvXjmJKY7QbklAC2SsRBVlvDetNKvrh9xInu8zEKzGhgQkx
8oTfwXyCgIaM+OCW3YdTG+t/XXfSma8PjCT5bGqt+FNFLjs/YhmL73+ReJR4q/z5
HHV7NZCIJXsUQ2UkzfxIrRCGN9BStEMI+PfSSYp4m1+bHwSM/lnRrwtwEh04KVDR
mAtNlIoqFi5aaEt57xf+sCMdCqlCMEied2M/wYO85/8P7uH34XVKRSf6EsZGjyzE
2HtPwZBKrPr8hfGkOVMwhc1BAKGIHpoloResVObq5DW6S5dEntiVq4EQzYAb8vV4
f8SKjjM9zhcBnv2/uhJTaV8JVVjOP9b6nlR0ph/6t5W7ChAK8ig5Qw6H+FgiDihw
1tgFE5TxbU2Rb4P6czItVASozALpOv01AL45L82AKFQwAQ8zaBsH8mUzEJYArLnG
8tT5gmdCtmUZTtQ6X/X2Ce3+3BuQfmvz9x09F3+cM8IlOYIBMEMA6mQkut0NnGjD
SjjHTS/b6gpvKLDsXFp/baAXNwEqurO1PqPx+Endrz5oc9XBut1D3Jky/72jPlB/
fch8mdsnEhNk4L2QnnUPhj1XG1BajuVc+y5T9qVntGAM+ba+70AkWzW6D8HffJbW
i6FNtKhxdQQ//Sx9jwPPRQ5tXOJeyVMHLyqZ6otP54f9HImpmo8eYEYCQJrHAhMs
oit8t9+dB0Z1rE6l/uK8SMe3FdLygx15KmsJuAs42bTcbJDHbIMAeBD4zX9AMaES
8U05e754b+GJazmMUJJCnHAvwyRsd4wL8wrIjVoXV+qwKKZR3UhwESK2lAS3ckdX
yLKb9vaBUI3trPMYcVdfnZiIebEj3JCXee0H/DNswsyC8Lw55p5Zi0Lvq1DNMbU6
qXPhgAWrKRdwaQXMD+I+n+ivHG4QnBpPFMJTPm74qHG03U4SXZxPf2NbzSrKDhUx
ncxWQMjpTFL6dvZH5sDzjYPN6loTFVk617YNKaYoE59kE51huv/RM+b5jpDFNaQh
nZ5vCMXNlag7gYW6kBs+vFK2E14u0dG2ak5QNSCEzrqzO9Gp9atdTadf+DaQ83uF
/wLegOMjTgrRYedxF0X1bn4bs2Mt0kdU1GurOxrgdrYe2NE461S+q40Kkf7TX14J
+KwhU+KhxOZyBXm02i9Cwu0+R6kEHxnBTA1hfr0CLex9T2+LJx/V/SBZZAg+TPiQ
TOGyy5CySfQN65BB24+dta0n/LNWsS2tERBxVStfpKgu/8z1VLfkCuZ9V9uOGYqo
jFaUpKn03vh4qi5pNxQYXC8Xtqu0TdXNXn2oD2F7/n6wRrHPgroTFCHEaZU6Livl
H8Ui4h///s9AAEemPEwDjdkmI0ujVT7wiVXWOXC/hYLn3UCI3NC1PU3oWNvGBm9e
6qnQTWUIvwzwJvPLY16ACAhz9esp9QYC8W2JSJeAOrsSXQnuVvMfOPgsSa8/PFCb
SIZdTWNDN+MRM38fiGXdp0Nh26gyVUPvUfQ0/rbSbNIjQgbqu7GDG95qyexqHZp/
/Kr+/5K4OEk6rXXFCL/PVP0KqwxchishRErVkTieQJZViQDcLFAkqMuZ4l8doPPP
pK3gPXW29NAH2srvk0mPEFv3doijTMYa0pU+yCOAk0g2QOJFjf2vwNCNS+zbdkwa
O8Ycnlw29xWkCLhinj5+jraVeR2tF2GYj7TDTIim/d7Txo7vQ/SzQplLluCA7H6b
LE5flZXtyptFJcQppXiZT2ERzhbratv4yN75OEkmcHFSNIhyw84+K1FCrcwIMdN7
GLr9WQfSyP7zfjwLWuEOj928kb4qF3gXltZozNHadCyXRpmInH4g0iexd9cXCQdN
cZsk5kYLDwhrjFJRiCfmA26YrdRuW95vPx9T2zmNq5KNZZZPO7eNYGN4qFNp3vyv
LkYop9m/4cdlgfKYJF+6gYc56ic9h0cmhuQMAFCyixOOyhnj8NEF2YixMLTFfmT+
vHSAZXXsgMU0jP49ci3/oGXXLp2EC8g7/LXgv2VlUmD2j5a9MNXo70tqWizC3sEn
i0UIr8VU4KrX2nztDxcpfh49SQJx3EpdXppjEyU00TLuqAHjHklGdN3EFK7/hzLd
FX4bAeT6L5OQROxzi6TtWP0yM1VpxlG/cOKvMStYqdOgRL+FNSkVnjdfhBpR8ptc
WBU549NoErA6qrF2RiuUvhty1pGdxxleouB3PI9PzKMLGl+yYDrQiLXVib6kgYET
v9CfqYXD5h78Df8jFzegJiQHN0YpT6536RLlW6wo8OTXyidHE9wxKmrXWycCdxtF
/vPBTg9bLlfoQfxnxLx4LzplOiC1gZKG7ZwJDJq3qtbYaaweLYxDPx5wtQQ4OCMB
wYkkDTBw5pyceQK0Dwrt2IEVEjUpw4xF/xPeHg2SOUtZOUm/EOm96QTfascwRB2L
4MIG8JjnLcavJlNoIoUD6Ca5J2Hjg0zctp1Ei+HDoIvUIpXHi0bKs5+WKWtm6ZH8
DpUhqYmZR9aKpgu+YVbmztFnYsidH4MMCT2B3W4EYNFAxk25I9gnM+5O4Ni+7dPN
EX/ohAHCvc4EIWPcbUELRNXmJNCvN0zs/IKtDWCMqiURJIsghbxjD+ZVm4TWKM8Y
yD5BtK72m5zE6l2ednLenQ5sBiH0aproDwa7BTuSrrOoRr3EZymFiiz45bHdrXvG
pqBcF8gp7JPVUVJ/lvoc3PkvNiHsysYmYT34E8JKKrLWKeYNu2Jw4OtcHnwWDTc7
xTjZkkNGTCXhRhG8Gwrgn+MthJrcU2YjAgrbx8cLuzpMowXOvm2SsqpQpnBreITB
B85gayYm33zho5//GumZlK1aEPI/RgX87W71dQcAOA+jVOXmaLzKrFb/SjpYxBR1
8qSPGpTrA0hfFYXHPJzNsmz97ZPbk7xOsMWD6h+MBx4ByJBGUYhDDmVrh6F7ZsR3
guGjsA2yit/JHetfvLxDMzYCUFiOPQapbqe9+D4Dd3yg1SfzZTSIw0Yk5yeTTyWL
JuasnVNi0MTtYztKfA4iyRQob7pZHvh1U8mqu5KhzBJ3kz+v5tlVjj2+CDdSxI8o
YZtx8Id1kdI3l1SLTRJcNjrXYykKuV0rvL+q1rUKSlHQiaUq5P/TW4jNfIHkLPG3
8JbyOs6NL6v5D+Rzyw7MU/9e6jzmXElgMv4NQmC0zudSu3n8RO1n8vnZvSuu0/QI
w5ZD+GHdD2Oq4cpGT1d8QH88/GTRVlW8UBvUn+NSADJ519lwb09mcRI8BtFUYbvC
BAphCmZXXqd7tDAimwKjoeqI50jrbjdcqZf/qAnuvqOqQf90nqWtZVfOe4JQKueb
v2SOrgG9hj3isy7GFybDjbPQZcCMJUfstomkO93DGp9NxgG5C08iEL9uRIV+ToQB
CyghuLZqvInFjTiX0Owisi/YmNt4HTZtfADn5esFStc1uv9PDsjkrvJ2d24eSfbN
q/Ao894yK4A6pgGQXL9r7zvVg5rWmEpfoc40xXn791M52gLrZzk6NWviLyBxuqVV
Mk2h5Lkimi70cf7o2dT6scFOdVp8I0BjrFynbzm0Mg6c0uBxEj67QXIa/PB5OdbI
1x46tnJd9nsRCX3a+ybqvl1Hq/5qFIFS6nQk42DOLCtBqT3p+hw+4DxrqyQFYkiw
0FXrql3uhWGAsnsFy8oJQBrZ/S/lQjTSbXtW8k3ARPtKggKytXygDB9t6jibXG/E
92qQpRiv6P0Zzzc+P3pekROL3iSqIcrWw0pKiottwUZsJCDwi1xVq+RWg+RL8ZTn
76j5bh6aBrrg2H6xXYuNfMY5pSD/gWXsXgPj16dq00EoId0yDkpbv7eRfFymduMK
OVmDnXV+IQ8nsYEwAZuDPAkkfR+N34zIfRVWXD8vlatAtXC/jm3fKRHix/KnuCtJ
+FvC9EvfalG1ps0PoRyTtGvlGzSZmP0E9VYdsGoq5wVmMvzMZaSwzhXgOUrfDOVn
O6eyJ3BtYtCe3LRnhQkYQNhtYZltEnwvac7Hz+uxp9T3bTHFN9E55009lhM4wEiX
HtHkMChNOAYu7zvSgpIV1DDc1j//MGcxbgtVoepxfQVvYl9c9re6ipHIdBiHB83v
GWlHDD2kvi9DkYMMsbzVDxdvabAEIZ0DzZtW0Zzgi/TqVKil8kPbpT/duNKiFLi+
F8ZgcGX40kNXe5oh+wvlQaUBDhTe4+0Kyiqkm0Gf9sQso86Vwkt0kqv4W9foCWGG
tmdMxTzXFqaLxj+usYe0+jRXakkXczD5qKQKhYKeKtoPTX/F9tjomgULK3Ja/uXd
EUtSH7spfoLZ8RpLAWcGRiw4jFwnx0qSRvXbo1miwO1JtAjv4lz88dn7VaQNoSyw
KNdHjDeix53DQxcTQMd7Qy+QIMrdpv0coEkxygA13+C/O6BlJxKEwoFsmhvQAQKs
uTQJhr+zd/rlrH5NKMQ5trwajkx2VrPRd+OGjKmP3wDLmPtHZjRl4o/nP/+AFyq9
53hQqxCUiN/xYl0TjnTsfx5l6yV8Q61nvoNEpbFvEUoqkbp/9Rg3uGRS6O1Krv40
qanfbyOj01i+KHxLGDqUhumpRXxqIYozK3W/AvJm2YjKycy6mOU8aQNFTjxl1Lf/
LknUwLqQd70xBcLDzHVChDbigyGKCc2M+Q6qECYekIgID9Z9gdkW8tjQT/eSXi0v
YH21o6bzwsZabR44ZkD2NhLES2QvYJ7zKpAOKfD9r1hOPrRmaM2deUhBNMUtv2eW
zzZFRJGwpkiSNHaW2ZuBI8T83vs6RCiH5ybN/tj0H2XkBKRBseEYTzppv2rb+iCA
DMDdI7/T1QtowfcMjj3ohUB7D77wcdrvUdLZdFsdckqR7LkPMYmOAliLBgN7tmZA
tHaOjeWsjD/tQP6Xv7cdMLiJk1LeAy+ruHcxyxK2xLWBq8hte8MLy/Q1SGoRukMd
AAngN218b03YbVcDsjQqUIbA+OZKl4BRJ9LqyMbMBNjqAOeCOY0PkNoqimQ1tu1T
n+3TCCf30RcMgKg2PTAwdcAJ+jdyekDb6epzKJwsHHhx+OGyZ08bLzVjqPL3JuV4
sgCHiBEpDYa3ojFCDTJ8We5tptvidn6MBkw8PYFG5Joi4JZbf6xawEaNn6I+sTJG
nxgkOV5LsPb90pnvQUQK5ugwzvpNuduhZiSgadgb8Tgi2ej8gIZSQM4exTKdspyc
jNsaMA95TWbl7TBtYGHl0L/YcYF8yF8sJisTpeF+e9E3DsiIkvasiksJJxkQaCD4
gbbL1ZiEv+5wFUqQeCw2geGt3UnBXLh1/ZQzisuX4y8e/R7b4NEaUiKGDg5pSv5s
9rzTLtCMV0IaaZbdVUV61cm6g5l+z2UcxAeZtcymdjIX2hemxDcyT2peJi55GqPx
WTWYBzSw3Wq4y3TpwB93SCjduKh92l8pCxQ166prWOVcgXvO7aFtSEPHLgx3gEDm
sAen4r1hTYwfeSgho6sOStRx6xI9iTFgbxrbeLlGJ1HvAorQkmfKhAqCx0y3Lytv
0oNaywlPmWfP51Spn21AClthRyMG1wP0ad4CYZVTAh7TvoHHlt3g25/ZVzbmkJbU
OQpu4FTTGGAs+DQbFGqDZLSE7T8FJ8mOrTMSmItHT++B1lD46/cgT+cLyqUKadKg
WCs4WI7qci5cnmc212mzAWh/HJ9m+dgja0NJicz2gm9MvHN5FSGXDNiaBx72oCvc
9FJDjz3qVJzzHRMJUEFAuI05AyfEwxmKs6XDL6HBYQCbzUHGLN/9oefnENojCdkR
xeFx2YFp/V5Wre9AWpZZIEEwkBARClacBryUTGKdneiwfOm3uM91OYLwdrD+uYXy
/EkRS/Q/DiIKsN/u3lrzwVg3tmu/ekU8u52Y+nE7j70FTjRJrA9SsWMCS/MHgOH6
uQRJbgggw9nEM/BMPnvI5+/Trt8ilpyaxiRXlw3iBM2N8YsMuKGshm0VEz5YVFS5
rkbWVqdZqVzz8OfyyZzhJCYc6hqhNmECQ1iFM1wOgFWgNzbRiM+VRBRIzr1h1Qsl
lmyv/BgjTgxqKAJTF32LkySZCuAdz/ELuu08ThNEVp6HWbgcptw+IDtiX/WceMfg
ul67xLc4t81PJ6NiC7c9/p2MjAZCDph5ePll8ujwRChOQ7G2TzoJh3OMOO/k25HV
EAuGv81Mn3kip6cE2We0cuvjLVfXyfuZWdJi4FOZVY4zMoYvx/72JuoUnAQF2i3d
3pAqxWNVb6M/eOzGHXvxsZDw378RxaiNJbgYmuVezLJR/gMWgaKKOYu5g8sA+WPZ
U8q1zVGRm3uqAIMZq4/s69j8L6GUVTDmtgEOgjO1Q8rcnT0jFfEWvoIRiYmTqmLh
wbKs0+9XTfCUTww8qruUELfroHMT3kcpzx0oJ7jcrly8P1kJdXCmnS4d4DNmpEWJ
v1BSEmCOcT9cOdTembUq1HzAP3G9nXWa4kfFtX6HCXSTqJgDyYuWLjQHw5e2B69A
lBnngnQM0oqM4g6/nURjOtJGcHhJjhMhrsOz8sgHUPF2fXwzkB1sNBd26IYrA10G
rwvCDl0ZbtZiGPioKoU0MveMSI+apiDKKAFgxKpt/IQJZPRN6CDyd7OuJdxEiy3G
hxo+xlhBDI5m1tfrqwTMC2lml0nskUhiW4/1zksHB/U6g0WzfLyv1r5K87U0WCtX
WizVJFWiV0MbnlxeJXMHu+RJQwyusKCfXsRtw1Z8w8z9n1lNGlqEMCuFnyJp/1B3
GoF2rssKOqhS3/iVzGfu4KVr7v3V9Z9Ud5xIKie+tSZzpEXPEI+eTN/tcRSUY23y
4MDK9Wwbl6FXYcfJ2RwdwSI6OmhDJf5Q32ICbGdtfKXSl1l+S3Y2cumh9RnaoXhe
Aoh+2//oKsJ5WsUa5u03oCwkAftBvF9oNzl/VWfp9TAQWrK/YFIVJs+CoKhJlhtd
MLsJddqQwEQARqncdQhDwcPTM/Um0xvHgKh9W6w8x4ZeoKlN/lUYhOxWBaiuewBI
TWPMibQmcUsdsEDCqLbBgsyPdLPOrptzMmkB17Xc6jDswIFVh+MXy3PMzXVUB8Sh
bK+opZeLe/iYleqY+7i3j/dPCwuMmWTkEhhkmrO0pg91J1dVIAklLHQtJwC/6vOX
fhPc+/PFw/GY2/Wz+fCUDbpnpCEGKKRtQwTZPbofKLU92O8dCm2rUpiUgEwK9C+o
BMkLsDK20KZrdgBu0h8L5brXU6zpaZQE2UsqKJSydqSsoiyeJFXt0eB6ZbGnJPJc
bw5tmDviW3bnNAhoy5PJdtk4Ho/TKYkEXf090AH0rH7xC53+M5UcA3SH/Jw0GGtB
7/T4RKhpGIZZjRqrQ3l6gimcsoJbZrLoEJH1n+SrTJi/FrcBdayJAQ9mRJqa4GYW
F3ey7Dcvy1oUaozL3CsQ3m/0dWtsw2lEY6i5NuhS7PJ1EFZRWHdsOwO/sC1HLcwU
AE+RFuDH9AOSc05mhTznsaeECDtzO4am615gWE1y7TlggTs8cCRbw3hbuhBTfY6+
cJ0lLDwJjMc5ieh7kO7LIQPcvUbQIaK5CHaGgsDvRWrjDmTj5Lwsezd8YLqeyjaD
pupI2IBZ41yOrGvxtE6+MJo2sz1G1jirjKka38YsTK//PWki8mu0KSpLwJR5l0v4
TlhbBszhTzXJxndLnnVSrcAwLMdEom6+JXuyLC2+sYsNqmcaDC1W1zp7ZIcZQRmc
wzHZoujs8Mg8kPiJDvp0SbcxZ9h/BXovrBsp6IR3esK4ET72bE2Y03JJG6qdab9O
BsQbpzNKbLJdIIXa5gKKkP9WG81h6IRV4rTYOcj56Y5LM+DgyFs58BEELt+DRr1q
QPeqMGVJpYyFHC/edDWcbqcrBLTTcsywkk465QOUB7ASn8PsHwGhkBxjQmDgYk7C
yP6zAlVnjzaAv52wfhDYTScaTlJAxqE+k1olr2CSOxLViFnZHkAJojbL0LlnrmXz
nv0rjuYDvdm850ODf6ByYWGn441LNVgKRLH7v2IQqin3L1lf1eSsrdsU8JUzcrYG
CQ23QWgQioKfLDnmSwEsrLZ4ryOsFEXeGQFu7wxS9lxEP+iw0jYYJ4I+r7BiWkHg
BOy9TpA0sZV8U+qnqmJlHQ6GgRFym2lZ7ueZKzo9TLrIZhPs+fh6Lrvmq7Wlj+Om
hjITeRvmeWBMtR4/1HJy7Ol+bjOTud3hNQU75A9K8JqGXABNTQtvnCeZbrV0I+NE
1ebXoDWmHG3oY/mSDOxagdALsE8zXkN6uxNpJ5PWMivMbtMOawWne7CyZdLBe14x
mwvXG4XGhVaw8jcIOx9TV60/f3t0wOXtIbWm0/f2uCl1s5gBiNwZQPyLfQXfzJUW
s628OWimsZhtyav5XwhKMF7YTaCmAD/fXe88U6y63S0NNfW4FtGfSibO9KIexwlF
jj1WTsdCdgpmmtQWca7ZjOAovj/dW9OuGtoCAqgth7V4nmMZpSTiBU+tNPM4hxfz
3DA4sOm9a1v+hnHzy+2iu0ovPssfLhVCUIco6+2MmP/1IA9jVXZnz8K2TanK+K4T
pn59hBZFx57l3dZLOtPmwUFx1lC1l68LiG6hUaEQG5kmT0FkqRhimCJf4owNMxf0
p8RUHacOx4wqSkGasgtMFnroO0ps6v/YcS/aYVFIh77pyYmSbDeEhhoOBzEGWW4J
oFZTsm/iaMwu519AaOPQIC+qoEf4GuwGOh/i8iZ0FYMm+cXMmMYu9A2zuVlIb47C
s8fGRbZVAVVZQRirWIjq/5ihpboIh6MRUUUy6UzTd4QI8rNAg5IxNP7MBdtFkuIj
dMr5H1qZ+ZRgCMNe9dbzonS0qs7L8YTWLWmAUkZQZl3bjKhxRpshnE/qhB5DQwG4
pf6qOHDZj3DOKXx6b0I2mnCQafhv6Nt/pk+urtxZvw52i9bt3BngpTZrLVxnCokS
iyK/On11foJGmeiaxUEylS9DY3vdlSDeousnD/Bkr5pReNBiEZ0r12BS6oSNOmiR
70nvzUfEt72mljiU6pNDQFrVHvCX798lbyWo5+W6VYz8I8x2RXt34BmPqmowYMxX
tuIku1xHcpcn+nNpYc2wQd2IC1yMPAsPz2Ys82qBat9SHexbRKKxxs0rv5cw0kL2
shAAAr8itv3YPTq6Jg64nd3CIaZkBSKDc0WxhsNYPoYj8pqBOtqU+MnlaynXC/1y
j16SHOBQiC7rkVwsGY3jRhXAWwKwj9YW0GMmkaQceZ1SKnDDMKTN3nwhAWRI4hnw
y1LxRp3Q7zFf5h9LLp4gnvA7hirihrMbl9NqX69/K3ScgXJM0L5D6zs/XJ7E2T+y
Ike5mZM5FhFZ2dhBKjaVCjJ9TJXCREiGE+dxLq+jgiBCXzFcfD5e5sr/nFu6s9i1
NNHaiNAwn2mEdZmcXQPEJI0YHEG2hxp0bMd/MyhYC4eztQxR5Xrwt1wmS+02tXWL
NVhM9aJAcyOH2EQt26assyCuSdI56KyoGWjslFhqz/WDx8zoavdm+/vrGKkyUScE
hRpHxJphhtmVGbU8XRn9LOxMm3KX88g8tpUuf+CAwTn6Kv7B4a1qbrDuhh2tjSv1
1hK0yB43Vip/yywhr5PrWdLBl51b8cCWb1czQk6JdRAoZU7ZZ9yrrkqZyrj8D0iV
AugmKTsXdrxeqASG0fobyXD3emvcr4ohIbcNzBnYe5hoL4qPE7el41dojUXMpKJg
vF1fzl5Ay+cImUe9v1+5dU54XTrK6DMpFR8J1Mv2IuX9PipexODmzlfyU8zhis1S
n6JNaYcoqm0bmQQY0iTgPpNUjExrjf1WfoZLX+XB7hBYfEA13Ja1wmg2Xivwr/M/
Xm7fbm0BrTRfVZ8Hg5FEeUR5czl61LjVxHRofbYZJQSTpro52ais4wQWWqhoQeWC
K5YtbKZAsnZd1ss2tak/QXV3QjcnJB8rMZGZZdd7VlrsNwwei9PnKfif1UmEyn8O
m4NavREkaA3hIOJkDTqJ3aSKf8MBWxWXWmATX20Y1iUJW/HvKqql8kn0uOYWpeIW
74Fv0Vxd8uZGmDKpsFPnePSXj251wv8+ffAaretFGJC+Zr/qlQMhf1blgIU9TWGt
LT8XBK5dyVf0CiIlSQW19/9RhNfpTmbHTt8ymrd6ABLXQ5p9G/LT7IM54qy1WRfl
sUmOyZCI5QoUopFcWyc7hw/OvtCc6ENie3sV6aQpvtBx2IvqgAg7BELubVp4F9pN
z1stFalWvir1xFQ9RyicFxwHuCnvxv+VFHPW0bb8jTsQtae7ut+BgPDwhHVVIMa+
mCBzh7aTWxbCWErxkOG1OnD9OTcjREyiX7BgwWXmJPb1B3jXt9ARHetbDXW0cvtZ
ANW3AQcMSRXMLL4ndrvCRxyWvOLFVx7INYziqayZJ44kMi734+XTj5AMv5GXMjyc
ZkOjh527U2P9JI63reeZ1sF0mjwihM2FaqcChU1/ZHE7EIAzJqyPTEs1B0ZqgJ60
oIrT86ehK7d3D2JC2K0N+V81nfmJ/j+xeXaqBEXvjcgSdFjvyzQqRfsB03Cc1ZuT
vFzIl2LKhwBP8BiOT6wlM9AzIuT2xHTLIS7yXzIfLtY6B0YjMge12rlrU35f3iF8
gpeE2dXs+ou2kZZazdRk7nTlUpJwWuF+pq6BTdtJyWtxjrZpIykMLM1o9yVxpkDR
fh0MkvkY57SshWofdmR3nwPwsi/NRE2PZp5kX/qDgKmLFRS9kUbCEBztdfWhd1jp
mBct0t4qUQU980wHXoBQmcRdu6FDYIlVMbaXsT5jYBb7zGGkcvf4UOdy4XBYJUxC
/FhUmTdQjj9TwUlMFGB0/8PUB1aO7eSeW3Y3QkzOTeexUiqrExB1PArkQcL3Nd2S
aUV2ipeHerGqpUECoCoHAjZoxzt2nCaTXg2T0si4IxLIgfT7MxvV5v2/Ens+AOmQ
gDC5EPtfOTmqquaglrCo3oAjnNCU20CYSgGDd/brzvRMzcM7lhQcPA8j39DTrScJ
etIZTkTYMdsctiLz4g8ET39FTtXEVvzGTR45WtFkisHR0kUsHuTGMxbPaP6Xgr2d
VTcNf6ThH+74RhdoNtJHRDGGfSPBEy6iSbDuYTtxZtwF1I8FvEXCpfOliJPrH1Y3
WJYjiFV5ih7SC0o6/j897loW6MPtL/kk2oviJCFv3ZTusorwvdpwel2PlFIQgVPo
p2w/FTgV4kA79yrHU7zRAOzttVuYKzLebeJPdzEY1xxM2/lfkYVtKHgvA+KlYlLL
0eDpAFg3VDlZaSYkz4qNExuI2uYDmGkuyL4pmaI+rI2cMmIWGWSr/ADZ4Ws8ANse
WT7GJlbTpXhm2xj2JNG5idL9KiI4GqDwdCDE7KLsaY97ElTz99VDCNWIITEloCKO
/h5e+WT0yvZE35UWp7eU7tu+E7qVSVaDycFzjXeeVz9diVpdLGCv8QBx49AuEngj
8oAuZWusr+5guNPOvL8M3abbWO9+Y35XUe2uXrvxIuFL2881N8keL8Cu45pu6FHX
CHSOXAayP4mAdJDFKoj3qVak+1PbO0bQz/j2h2E6JekSksxJ/FCcGfQKUv6vPFq0
sBrNhEHrTppJGeDHp2FjskmzHKc6EpUQ7OFk1fBNGOMnvi6J/ffxPnYbEXHZc9Tj
lUudEZ1ytSLJQxRRhcoEUiRf3AxVdTtnCEcHljff4cToNi5EQ/K/HNlD1yKBN9Zd
ReA9wbSwdpo/thNAG44noBC7Nl+JFAjIBm2Nv/9rpPTWGHmhUvZh4X+G8nVWl8ms
KiH0YarPbpLjXvJWSJ87pTiPDwcvdMSM15K+HYIcEP4z7g3VrBuPt2T8RVgmg3O2
w+tM6TqECTpg9bjLzgiRW58mQwjnGeY8UWII6NGTjsy/VxX97dk6o6U/hHRuIgdv
4qzet8sPXIGXPcFVdsHRavjX5Xez3SbYNMQY89xwIyWpNhpgvzcheduKGwZ43vkw
Cl8EELw+/SkJvwfVLTZMF+sVR1x0f84X1UT8jgS/B+bNRXzKzot1uWmYdW9HfFfm
BGxiL4N6i0ZrlgF20kcFviSYXBtpX1qmW5y2xaVbLNorj0RnCHIbYID6NKRS/l9q
RRmHAtZGqeNkvd9uDzPhV/vE94j89TgEXfhbNIhQAL+P4Q5gFOqsy1Qxnf1tVD5X
pv5Mxt7ZzwVynt12VQwgTyXqJ3ZaNaZN6sULRXVSGaO1BZgaX+GXekk241tkVA9d
CoFMmOy91BNTT/pf/xurCpKs2nagpeIIwOhe68AhVF6c1cu1gO/qgWy0/jB907ny
QNl7ped+zAqxehWFSMYQTQ7BaFz4gJ983WQOkTV9GegeMTqPfgnmvyNWF+g6yF/s
acFMFDhyP6mMAmulGylMA/kmhrdo7+9UKIDHJiQuV+pDD9J97lpMmDLNGgvWc1OY
hNnwl9R+0T/EiVX3w/uuHcPFDm9LZ5EF2xpqOn4JEeYAXqMeq9zQNrDTOtRXUGJ1
OXQm3b3lzlj047+67qEHZIx0JGPGIHHrY7mlAwtd1/pOy6sgvOAuaLm7RqSopeEj
B87X7noQ3QPWPRnJIC+iWSmXbp/sT6W12lLZjWXaxWXZ7iuqu/33AAoavCH9LNKf
rOeZuZuvt8fxQlM0PdKX17d0p97CU+16NmXnEGv50cjPAAyP4agjgk29j8xXgcPC
dwB7cJbq17DkjbTSZTfI132ogkZ7SaqwpC1dbqoIVW2ev8N9bc3NqDCQqk7KXCNT
wisTuiT9WVS8GU/O+3S0wAqxN9pHMoyfviqJq4Qxu9WHLDnF3CoNhbPaq6VRCQ70
Ju7umngZk5I4Zsst3a1yqA6nY79+gkV7KUHmd/zg7AY6zhmTNoY4riH4AcmyFhAr
qXQa51C2N5a0xmkLkFngLeizC/xoExmYmMAlI+K8zvsa8za3HBFbH1Hz3Ap0lMdf
dBMTk8WAdP0+4kTPhbgS3LSOzC3rNXJlM19isTZCMd5291U6MMYOWu0CpJR4UZal
IPj0JQ5bf+IPAlUA25ojF7eci3JforCHKpSperMmWD3dOOPIN3jszxqOsMVpCOyK
HyRqoL7OZYO+ynhrKZJLj91fT4BORPrtej7JzWDWYiZeWbRUe4BZWow3sBqh1uh5
3IODp177PoFHfMyDBe1GDd/N4QRgiP4NGK2H2gRQJSqZgV97NagFMCtOE8O4O/9f
Z/rfr+JHkaNsFrr4CDKm33aPcUhuggLh6EW13JIIr2UA/hfdSXj4gvMOoUzpOht2
B/IYyvQyhm2wHIR+PJmeFoWi1E94R3AJigt98WVlbjrBwH6F5VJWZjUaiKZH8Aqp
Xd0UPGtMmAsQ9FpfMeCzJfbKl7wuhjnn7/XzdjlATmSc/nKdc6ufmpH7Fi5/v2lC
hEgdcuKGIg+1WvtwSohgLGkEsPMThr2P71VtG00mrt70hFAo85/WdywLIRG8wCYN
Iz/nB9nmHGjn+qzCDDvDw0nwPb7058Bd2xcqi4Gdfta4v79lk9hHXwPOlrCCPHb+
3KOfG/lPRjyq+/p4fuGfmUF8FNXlyr7p9N8sitXyruWnfXqzANOIW2wLjrK/fXhX
3V9mFnAi0LGQ8EMlZsDgCD7tvKJ6TEEFkXlPOcPhcAlKXBvkqDhuCAeGPTeo9Nb4
hRF7ALieJzmou+ylWp5iaxWN+qH3uQbrNzsXtgPF/9ZbVu4XP+zkFHPiANbuwUFT
0PZaIpNhnNcI7hYBBdOrQuFYyLwv4Do5/4BjRMZonNy2MWsjSz2kIfvQTDQNIXRl
W3mrQrKXz0K45n/S4x/xH2+aP8j1AgVSn9pfnTKCBOxtrrEUQGRh/AVkt0jhC6Bq
noLckPONLoww7m97BmmiDUMcVvZ9Gbdt7JXn+D476fTBABPWmEdZ1irNaT9tyoOY
RvZVTXYDUdk2Jb54Td4nz89ReKlTx9kfwg0Ib8HkT/gEw/E0mgnX9tRTwjaPsJA7
A+jxs/PMO9bTI+zgZuWD0NiGsXrXq9JmH/LcJ7c19YVl0URl9SB9iYX7gEMCyH04
wim3JNojG9Xl6CDRA2Q0dK5y4ysPC6JM9a/rmxshBmR5U3pKeR/y1oBnO85qPfL9
+kUNzxImn8a/fM0zC/CIRQ8u/0eI+bCUH2QM5Vot2UWVplvDgxvtw21qNas76zRy
VVsNBZZfJaw3HH2Xg2kzXMha8VH8QG8g2cu1MrhVtYMsnOvJIa8Qrgaa0LaVL4dB
kJOL9IjXkf9HqXlxA6BdeodbSmU5yi3UeCBlWsVef8gq6SYpdXFpkqefz3S/l9sN
tDI6B3jGVq/znsqN2woTaH6zQsWN30i6tx8ZMpNvnaARcmwDZ4cQfPW/RCJiXqss
H7zbzkwUbYK1gCu4uqa0sb6iIaNMSS4eoRbqutIbMhJWrdBVvhUapwLBQOhEzvFW
ANaK/hiPnL6Agn7bhEcGf/nAjqwRG9J4zuYcTjWp0LWpRn839de2KE2RURNBhNis
ODpCCUSyF1fmtsVbuewYyXWPw6mVyJ2wLB8PElfzemvgFAPzvfF1/1mKdn3VldN4
2v9MhN+tveMBxvW2ZDmSbUwz6ynA7lLphWljtDg3hzWJIPjiqd17690Ur965jeO6
b/HcNgbaFcfqktjFt5SIY8cFFEDTFu87wv7/RTBKCrt150st1Yu5a4v0+QtwhOXC
+bAiZQgkqcdh7VYMO4JAFkiSuvxqQNqwZkQOcu3n2ovwW95H2npFXqg40CBKzKpx
qUpVgPb1Oggp5JYCQhs7rRprp+yQsaRgx+B+PTFipgYwmph2/U3yvunJvG761yMt
X7I7Je6TgXUyeIh4FCe8UvcVVC2fGg3jA9HxjlkqNSmTbUz3Cthh9SHOkSq9yUtT
dbX6YqNChmnVBO282jDsTEktDD3GgzlHd1+qaaXQQWEuC8RKcNfBYEWT7xZLXEiX
JgN0XiNW+h/0rnlWNWwN1lWT9sEkmRCdy5lp4gy7NLD/TI1Wg35itpPc2WdEeXWd
gNWAZenaU6ogt/5NUOzsGfPhQMPjxp4FEVuCrJD+AfDYy+QdSuFtS3HdJuVyceDP
IBsr3vIaxQv4O9/Qs+5CXOTW+IS5sk8tke/+ns2wghv85YKJnB7Th5i/t8toXmW0
TRbkMGHjQ4lw9vM3K984ex0VvZO5i9uMToCVeDXm+t+nhAnWDqx5Ijj8ZI82n7wv
ZLXUhwBhib85TZEVE2x/pDluZE4JWXxT+OoTYIt60tYSiGjBy6AtgOpNiwafpJ/p
+ipgsgIbpx57c/CALO66jy6S3TfoWxp6rS7yVvRDIVjzvffFn1MGMy0pG0h+4BB3
bzQnZCvXxaFl56kqIcsZhN+e3DtKxOAb/m54r7ZcPt7TKMb6asGv5waukJsR82TF
Sv+03j3pi8c2eFQBp7q+HLhbhz9o2xckhuAH/l2o8VlB5R3QY3OYg99/rggDyXue
6h4UfMq19fM2O7SOVGBd3gOXni6AZWIqMpB9ciBCSMuckw6L2hVswSGpPRT1cNb/
/Z+tlESIGOZviY5yO6CIdoz//GSEVgzck8+iI4y7bqHJZCc9fHFTW25I9tGniQUE
HyqfD1i+7mq17wkmjqnFD7+icTaO7Ia4zW2iByZ/k6SQ/poYS/fv8DGf7crLMZGY
aBnRBZ/LNgD/OhRt5AkrLjQpswD9Q1amosSO/+1jky5jISdlBHsNi15eH4yPD8ta
0aJoB3CWg1y9cqN4nHs14EJzev7JD0O2Tk5rLNMVvFhVQiCLGQCrQEp2QmQm51si
IPnBDzkk5Id+mXU3S5FJgK5xoL05L0/c8lzNyTFIkMpQYFLt9UAqsbeT1BYp49rF
jU5JMy/y3/Z76sS7cjEfwloyQbnykt+9tPAtVhiDNIaX0fYg9rfoKLw3zDTcpPEM
5CK3NNt0Nc4y6J4bxlZtTRRqWEKZwgOmJSkhQnxEIaTlgCxMwwYChsjzUAFMZ+6i
ktnQv3bJo9945u632wahzISxZy5tiDzSOCRJkqUNP1VuWJwBOT/0+wwg6J0ZKiaS
d36TL83zi7w87kKQdRUhu/ekf7PKAohcL/TM/jbAb0g/JiAsvztM2yR69ed6hUzm
ABAS85mb7KkLjccIjbmGB3pWgoAqMWQPG5dTiJdEjpM3FTM+GDMZH1iDlH7OL4sn
UQMPZbpuEb1KW7dSJCNEWNwbvS5UDh4UV8qAdCR7zbrJ3TT0p5x+uHMPmtffk5fC
86f2dxOq1yO5YUteAwdX09Mc6WveNRHTkKGCRP8Y48QuBX6EIyooF3u7d8gUDaBh
EnvgiIfDot+j/wkx/5Bxb2CrvepXU31pQzXlrcTqmtzmIcrfOms75JLHA1VZHVrY
mT3AnSFfVS36Wy4T5SDcq/MTyNewdlvaGP7XcDQukYamim+cbKFzdBAFNOX/Iucm
bM89qQ7G+efc+pLgF6v+n6Fdqkn9qEIGSjAszi7oylXlmHvJHTYzOKzV46Epx/1M
3MVenLXMyKOzxxLp5wMCMewgYJv+aFO5oOGCCxsM83P4GHqIxIdr2zHGHOEncKBy
PGXzntLAbV9O+KVhauGf8pS1zOjmORGqW0VK2sqlpGAs+hNU2pAhWxn00ghXVfMj
m0ar0yWMW5RnwH/XDFPLPbYF5Pp8E76oLDdjz0MbMQQyk+Quff8jh5b+1/lAEuXu
9+/OESee6hNYAL8kgE0qfAKQLgpVZSMYppXOUy/Xg8LcqE43CE/1DDMrjRYNki76
JGW9Z+e+MTmccj8TWtFc5qxDbQN98bUIL46eqnuWXqD2mP7bmHWdLrn1iah+jLUH
YvnJ6q4LHMQyZxV7weXe8WiTsJyoiQDwctClvaCMK6ZOnYQKfj6GfsmeHdw4Wdfg
CZIaR5XnPoznMJ4Wba1LbScRHy+A8C/ZWbxhTargIGxRnyuCoIz+UgaAPP80Oolu
qI1fIXxOr4lAGXX5pFvIipcxeb237SAzCbgdQItIz0gAWYb4c5SuaRP4s3jX7aZX
O1gwiey4BBiQ/S5FVC3jHUunrM9mPr9pwqKtP4E9SuoRJLCC9jwJb4yPO2s9t744
ODw7JGyI/Csa/cHzVnF6yKoAWEvFX1pYc39OcnjPryy/YawBttvXzPBCe8kert3i
JGoHzu41fku/I9PPwOSF8a0IBmy1M1ZiwJrFv2e1KILqGPo3/S9SALjV0TvCVJAb
G4b13acN4LEXb0oW6aU7QhAtK8FoluFU941Mc9LDs8m3v0soehxWZsqmWKfC/ALC
tUElw+2tFDPt9xSfXdrztjg3M93rJhLbZmNdIc7mRNDlqrGn14lK4oIvuY20lQKr
bRikWSit9vAR7WBoPmiHpdnQNNxq8tuaFjrYvEy3bB1Tlhmotlnfwl1Wew48EIZc
Rxa2T5RDo+I2M7jPv1MwyG63kf04FJHv/sDebhXmMZtgr/WnvFrHYEUFIlEuaBRw
dRd25nuhmTCwV4cKs85srTMR32ktDLkg00G2zfJIkpDkPSvt+rPFF0qebAYgx5wT
M8Z8n4KRD9PVmU9/EL/QinlVBY81TkCiAeL0stNWJ4HFaX2cIj5MJyaZVJH5Wr46
g5/BXZIlIsP0OeLe3BM5zz9DsAbxjSpdWWI5Iv1S+y3nWCqIzCXShnHmmDx9FkkR
VedYVNjKgaXx0TPXlVVgOzLOYCsanPT3IsvHqRwef4TdXlpdbxIdVKqcLtdwXXoz
3i4tBEJ7jePl1xFWZ+XuEyA8klr2lSmRZh/7lCmny4RrrdMlOtp8u5sOMfCT0Z98
z1u2V/JTqsKNQzvy0SDLg3Qxn3vRlM7dfO6e8icTZDuBbCSc/ZU2MuXMYnPVJQRn
jShXZCAQFPkkYFFBHqx8p7PsRnZMXhA8iAyJW/y8AUxYdyMxl1A0Jqv1zvxovqVY
O6QFbKoq+iXFvqCbvZZRjEe2sPf1iG3uz7HND8dMDN6b65cw3vZplGQPo/GYbRGs
yxU+sx0r7emK7+Wf9qAJJs2dJ8d8lTCv2SFIZ44pEj+ptJP8GH5O+R8grq5VtBXY
lY3J/yhdB93UNfgqFVaNDVIZQ+LMX5Tj25tET5FZwZQujMei0SrhKKIkuCbQjwwg
grt4B+tUrHr856TcQk6oX12YyYrtQLsF9rk1d2KzFOxa7utjDKWvpGFBQmt52sPy
dSgjH+yEPgQBNcHV17ODyhEh9JpSAGiyANekd6U/s3Pot8FizsWHMn5HSqmLdpGU
j7vU7hQls42E4LljfsofDUfDNT0ZVsjsLKW1KSBCg33XbRg+LjuSavSmqvACzu9f
/ER6fvissjkYQo9aCNeMYy1I+cYbyhhDJlupkFOsAHSZrrP8NMYGpNgObc9gFFQu
tjK0BlLw6atQcnTX8B2JCvd7MLrTPer6vcaBtLNgJlxX59w7I5Ww/sb7uTKSCtZO
g0NjsVAgZc01IM2wOmqHFpkjthUPFVW8Ep9ufra0gfiWiNr5jQN1slnX4bEDnp47
Bg/asJzEuhllhADSuVRMgtVxh45MC7Mpya2JhsqRDu25vRq17HnfI8lzMtwHPmzQ
ghvugLvwK34b1Y0R+hBFi+R8oq6nSPZWbEx6Fn3sStz62OCUsM+7BFq42pOSsETZ
rXBQ9r/HLlCrfsXUJeuhEzmxeFgirZ7ncGA41Snme4bPoz8qvPptZGTyLyF+Jhpp
Q4D+dszJRZ0wBtzkGoekj4ru0ADhMtlyNF87mN/rXC3sAKGxCHXY8HjKkex2CrVg
HAE0lst1MRAPZ3UVDhFFlnKu1RFTK/OTDF8jffCtM9tRP8ACDRKy0Dp1bfXTknkP
VGwrVbXa0tbO+KDXY67QJ9QR1kdNmbEPOUt0dHaZt3IbSca5M7EeUc4P42Bs3JuU
atKMWHVEOyABgVw2pSVF9TCL+LfMWU/6oCII3jS13rKPVw/Mr+odJrjjCUm3Dnyv
2iLl/o1CjViTqhcROj6lL290J6CCtxONxmlkMvNBZpsgEv/FWpFCIPE5o+ehr8fr
nrmDoP7VPf6xgH9frusShHhHZr5YjLM2iIrxBFJq4LlafZkafTp2aAsoeDxJ0k3d
A4r5eU4dpCGEx54irG+ktPn/sGRgkrp3w9uG3jrGZoMeCX42kHwdinn9fu/Frn5/
spSot8pW+pGbw+fbdkAUBIEU3kDAquz+FPoOOkCj5VsJfjNG0oY/2eZZ3abmfbmS
JPjm7N2RQrQou0cBJCgZVgbfRuUm1NmpQk6segCSCZI1DWJ02X8tkH2v9mEItwRa
PBW+x25qd5vCrKvOhYWbYewX080ZDrzl3ZujiZMDAIawBzPKCCUCHOkMkIWaITAU
3Qr5TE7Px0ILUeVdm0Af6IBZcSzuxjkY9/fHsVUwEWVneAc9ilnTkFLtmMQCx+UN
ntpS6xejl3PjeRquSUNcIz1W59TnmhhNCA4d+YD0BEPbyG+j3AkUooriTi+1XueL
l8012RIfKB+Qa1acYBsRJx7mbu68ltrrDzU53rGvwHdhv9vdk/Ow4sWX3sx1PA1/
lvDHTVSYk8oI423rqvisieEc2EWr8vcLdiRMxq+fvCNbP6ONbnGvrtcYQx7IVWr2
GvMU3pIP9TApQTus1ZrmxAPSR7TYTgLJApcWoZzfq47wbOKgAgzidaXY95814JzZ
SIoY+3jnMkl4SE1UsjPWenr6b//XKwyWTqYGa+fhymT7xYGTrI8kwpenGtpYXyNx
Hv7dsUAvQ5oaL+T1QFSJqhhcHkoIYLaxBh8AbgmZqKgtXKpNGe6hkDx35ev0V6u3
VTtGbkprP6WT0uIsIqxYVJNw9+CNXsVUzGLsy021zEeqD37n6wh48JukHLshYhTi
XZ8p/eE+/GSjt9pRFwhSVFfj+Ft5f0yogIw9Mi7BOqOw3UzbwSTp30mPzMs6C+vO
E7SV4y8g+bWzgCVlnb0EGxUsnjvYRv2ribvjzB8RANrUDS8ghMiVCCrEEyQHd/iL
Y4sSQkr71giSDhBsUUdAQfDIsOv9xfOpWNkETyicLfK6W9HleRD0wWrRB/31HJg/
KhAFqGgNz2eBZz9mdwAkBfyeI32UO9P0dRytRxd5YjOcviXYfOUQSzZb3fGX5Tca
NNwbSUKFvIYd4dmC+Gndn3iflo9+aSqAcXtoMgQ3U4DkTksQRB2tBacwMr71kmLH
ciFhK/pBzPxxm7ClIjIyS50rYEiNEkBXfFq/PCMZtCYX44QWX8UaUWJVFZCpZugP
l39WskmbxBDZKEm+NYhN4XxF6QxTWNBYq+15EzfB3phmc6kXtKHKFy5QcY0AxyPK
ihDJvPHo8c1o7FnM9WkmmsdXZtjIjDYYLSvFpejWZQ/Sfkxnj5dkg2nJ/s9pYlSp
23+w5w4RdsLay3p3Llgc1nhFy+mByGjJOarFxbh52/wLLxp/LthUYOAdYH0ytrx+
z4IC1m6x8fYbvfg9cu6hL6snF0buWIqsa7equ2Aj28gotXbtG+zOMnnMjSm8A6Sz
/e8l4iil6I7KM6Vl/+CBijkpkEXQ63bXP65iLUMr7gEUGlnN5TnU2FiVASDdzxun
kN6JVJ4f0jDZ/HFYZPEHua37Q0VGbxukUN3a+gd6fVUXypdRU221L7q4hOgD2VZy
M46qal+4RjlUOLUUpaCN03AXgyoCvYlpwOo4OQybWETY0Vv6jW+Vb7uq0SJWDdss
c0yl1hks6EiJd5NojvIFw6+I7chH7Ki/b1dzX5uRBo1W/7lSCkoVRlPoXE9cKKJd
sxPxNYLpfeLquvd+//0wWNT1Rl1NQXplHXNnSDqEMU9jJtxMJz1lmVC/WrL/L5XZ
rTJwerZgZk8jHgYhK/OkzdlM7nnxkHwC2N0fv7wCHoMx37e+eiwLUHqI1nadkJgP
AIoGSST50+MrLiw8PXuZh+HVtdUFtCTZksifhzH0G/miHpAaTd1R6voc8RVkv+9m
mAzNynz4JR42kOx7ThsvX/B99+TH/Obrjalij36WrW+ZBX0ofGDMSuHKOOmjJNrs
hiZ4CZ842eRA2g4n9UL9x//LMhXiVtNnThqFz25oc7ZVvJCyI+x7Kz2Ys3Krw800
DT3LzUrEgSr1fLL/kNf6cqL5iTUv5vXWN6uMZ/ss+7ublpyF9wBxPcPG0DXDJ/DR
x/4K2qU4fWhkpKg6LAHOLhHG6U0+RVQ1Y6jYN5Fymk2cZV5W/MWZ1ZKdFq4FUhxi
AHYz0G601x4xnHG2iPz5cK6LzPa8TOyZxWixJEwm2Q2Yh9tZf2pTjEdbk8ulT/PA
yfPSl3y8FrFq/vyLsEq7qxVVNPRS2uVatZD+LLbpjl1k2CVH6CIKJ3hOqZg89REv
gEqVzL2JrfYcKRWFx6R1dI2aSoV386G1mKIPnUks0auTHZYcg0xfcvJ30zNaN7Zr
omV1wEQ9aQx+SJyEUE7ZpYKRDbDsrYRVp2yeOACQKw22za2jvlb3pusa5Llbc7Xc
2NA8xoTQM3En14tzoMtzZb1GLt6KD55v2lIjYEuyltcW1jQmTeoB6LT7GQHX9mqa
pWBfk97TB98Pn/QZ1i1fZCNck4l1JTpzkNS3nkkhAv1pC9zKjz4oqxhLyR7kzQwP
1EkYx3j89ffZfTRpjqOqSmDVuODElsSRwNFQcbUupdCIdZXJ0qBYIwcfZJlLzTzH
rj66kU3jMVKKDnIj4HNIMxRB6/tx2rfrI+LIeHCLqy71CDB0XqFSpQDr4kuTGGYp
Xmt0sXMGYyJv3CHad8yrxw7krWh21auRDfBjsViKYYnruq213nQ3OeNQ/RxYz/nI
yDn5tHoIvOrC2RzXLPn6RoVwtvab037zdBEIrETgHJCk2hLaUq4cCR1Bg2ZOIrHZ
e/1EQtLOl0cLNsMphFCZF7ZLzihfAPjZeC8M4mxiO2zJOsxDlC+kNEElJq64XAUl
sR0QSazb4hnfWnhr05EfYDHsg7CPiOibOtVvKeVfIsSaVEc3eS83Sgq9+Y0Icwd8
krfHj5f5dH2vgpbZdVQ0QH4fIbZtdu+RA65M8oS3QKe9nyJ8IXYwdZmHb6V6r5wi
pq/ctSYgkmfgHBjrIgU8mEQAVXWrT11nUExm/9M9eLMdlKm7wOl1oPUYzpYIzEF8
s08pHIr5fHdJ0Fk1sPpv7g1xQJeh/DPcG8xTZSot3IYTpARBFuy23vK28ANrCxiX
oJfwZ7IrE+OTt1pGAhWHplmKUlxasoKYWtADvuZ9YCo5LDMRtSTxbiS+X5AIz3Z8
l5kV+FJ80j4gByDy8+Mg1dfJ059BIPEINAj3em+3QYki3Ze0Ym1K4xh44qLn5Wii
rklLzf/P28ZdTJ0L9Vw/GHj/qnRZBZpjUiK0rAfCA4PiaGgXTTcHZewAT0mpAmCZ
TjaApMfLgq0BzFZgoSluECwWv2scKu1oTgdJKXFEx4NxATv2g7qXZSGhtaShEZUB
N13j11Zb9Nc1YxMiqGQ45k/km0CApcS7cbThKGhfpAvu5ijTNg6iUBjMUbnYP23T
Yt8ER2UpMdHNI/MO9Q6F1LZS4WYYay2ECy7Qjascw4mQxgPcdGMKSQM/oKeryKjp
qaM94+6dcdxj5r62E26a/Xp41l7I5L35lIgQYf5GWuBii8pPZ4ravuLOLBl8vmjt
ktIkG70Wk54w5Zr97p//7wD8k1nsmbuWUfpLgp1b+3uJtYD8oCfXMOZbZiQEzyHj
kZVVn+IWDFjW2rZLT46RfxS0gsQok6nPuZ92+Ui++kXx9LhhBW426xrIHdK3diBk
8y1xPRC1uahYT2ffJA1WvFPKDDlbhGdJHXYOT8+36ikGCdXeuoWCxpgsMQFF6WiX
ldfXDLe4y9xVw29DlTazrioX5f1juophWYZy+w/xKM6+KrO6r7F2MyVl4NgjiVIK
bBNyS4ZIeSljto0sq6I3pPvRe4do6lZeAGEFxgQ+LDIxwNKfniM0OiasaznnUleM
2C/q0oQC0nIIsnLMywtzwFUBwj/QO6HujuhBzmSBRiditjSP+8auu4OkZ7b2VNV5
1pTiqPGgGc61KWrSThQ1D8AzGkvqL4wL+frsb7W/Dytkvyny5uJpZJQAWLbSTLz5
DvbRoKbaP10bcvlWHHNMKk3csSHgg7Soxtzq+NWPltiM47h6zYmW9V3JhSeDNCa2
VJtL+6aFWWbbF4jKoJ4ZMlOYbgXNPDPGXEqxzVQnBjs1DeWmZ0xIEHtswb5R+LdP
pOF/7VivCtaBQSmSuqmYENVTwzZqP+kbNNog5KQL6PFxP37a5ffaGiBIH/SXMwi7
7i+0Z8AD/n0pgUDK3OKbNfnm3529Az8MY56rBwGpTRxAW3YpiieuETHGCOLZa3Qn
LmZznIPm/OBEgfCMVEPw47mKFYrRpN535hOAQlKRjK/FnOcvinqaDd2Wur2Qqma3
fo0UhnqHBSRv2AkFwuNBCpL1HzHDrnpJoqGAD93M1OvmNBM4u9zY5iZaksjESce3
jQClvnCIpvyxJF9l4eYD2XkotJD9WuGjLQus00w9u4Sc9HZc6+LMj37AFSxcMbJc
J04YTE/Yh5V+BPgmlotiUSnddbsTZ+V+VLxoJd5hM3cjJS0jekuuelo49PpSpW6s
Gv9SPrueZKSDA2go6rpuJ+gnprm/xDR/S26xLfki33frsVpQE2UtyrKCEGTOAdW8
yz+y6TSNe2+mBzXyq2wqAySTnfWMfo0MQtVVob+cTTS46vt7eQC/Xc319r3rlKBb
Mu2Q5R1q5Gf91Of5uFgfa7F8JHjtQmpDZRvPnJmux0HloAQOs6p9ioIdtkeDU0Eu
WPuFh7+rYbP3jEA55HGX0hT9RC7P+uqAVGN9ThDYf+K7782paQCMOvhWOoTMdjJI
BkZ4HQDKBijwpICUd2Z4GxYipUBcs/5v79FbCKZWhdO5mXAkwRW0DtC/3GivFNN0
j4Irjv/HAU/8FgdQItJnY66hhiEIKNcbX38bTQmcX9hQOud7vpNq+qDokzvO+xVs
wfiaEqjQ8VbWZTuoSHp2ahTTO+rUMC9mD42Z/3eGEk9PWNe1DIoMg8KfodSFOBJQ
Ys896MaSTlnLaTP+F4Bx9c9eXqCkfTFWxUw5s9saKgwfJP9t33U9YNDXWc6vUnAZ
Z1Z6NouGUeCt7ksroRl/suWQu1z3kmz7nWefApnijy25qM2yaXF96Um/EIhFLRwY
CZks2DplAHSjopGClAr7fpnS0h/XKODYL4o+yU/L9YUnn6QIg/0Gqqh/+7uSEeX7
UblLHJr/YqCD2tnDOPhrhU7yTjsmiZkkr3fiYviFnv6Nvw0pGf0MURMfZMvf2/zq
JaKAoJ84OQKGcgvQnMWJHkrWJXT/ieOJbhvoLEdDXgp2LVwTp9dSsaJlUZkcNskg
k7SA7kKwUcrO7G07qk40Bb0p1eCYsSz0xD7y8NqliogTJtoPUV7faxoDSoF4AIJv
LYXJi3wZ4ritzS1LGyH+PuXE02xRfs39szpnG5FzP0JWyKq3kPTbkLZ2DFukmcDs
X6PPk0eS5jbVmUlr/ct0sbGGf7VIc0OMly1R6jqs0jgrshOMzlhwItrUQaJi9Y8q
9i1DoV/MsiYiyuQvBzqbqJQG7+bdP83vFkUZUu3qXBW0kcrw+sZxPZnPOot9sQuk
8LpAh1961JhJBZumBvIRQlEXA554h6vOafIJQrcGNO/a53CJ3PfTXz+cFeXHAFwS
/uS4l79caU4w8SB+NB6i6ne4LtdZAeEctz9z/x0BzXvtWZQfZD/XHtr03e1BI5lY
AmUqj15EoHH66aQnYa711JW5UTvMWPfl73r/a0vwaFoM2MrH62g1GmvH4B1bu+BH
V8YvhgjVmPIoUC9FalKaGlMy5389T5odzrvw+5Ko81ZUu/K1vq/049tpptaSz8y+
AtvPhhrdTpAApwjiXDn+GXeb2i55GgiSTU5SP1E77TedYXX7xZLhmVEofMP/PsMh
t0VBjs4T/1NmKrlDDSSSYNWyDIKgVXZMoPQWkhdRaCuavpW1AnFW8PRmLv4tplzR
saDdIaVRrPcV0v1+s+m5hJ6p/dV1lToz58VGz9nP7yistug9xeBjHwDz+eTBZyL6
P3qijSvFOB+rmclLFiqBaWBcSP4X0Lfa9QHD1N+MorJa5fOX9MFcP5wxtiu7kfK2
ee1qnDm967eRP21kdgapM77Oul9B2vvsNPZCsWgFR71zHx5uqzVtT0D2h1LibBhM
fEcB9wRKWdWtSWMFYeXYu3JNc9s9gWORb5LGP4TCAmkPQLWoSSjvG9SZgtxUVfSa
GzsidTNJ7e84trJb6YYbe4OtiQLS9Gg8yKp7ic6YNzBiaxNbc0Y5RNDNoKZu7Zfr
ZP967AZsrWZ4Pywvm3ZubH04Jl7zJlxRFJdKEWJuRlg97VqgRADdU2MNfuUFMKxq
IcjXbLFG+rWYf+8N6cyMw6btxRSHKPtVuD4S1oIahZWKBgk/HKTitSCdmuYK64R2
AwTHqL43r3wD6ipTP/qv+oTbJN1SwOZ9+n+XqbEyLB2VQsXIHboacX+qkdKa1RiX
uwfIbarNFW7q+sHUItWUHFSPf8TAyTXY3xfqFLLIHM3XUvTV9JwxFAoGgQzXjCk7
4EWmHTQ8tsAyxCJiPxOSZua/aVbcQwEMieSY39XKY65OUcpU9wzJjEybcoBsQHKJ
E1t2BvgG69qCdn/Nqo7PF3v7fpg1YrxZhRmAd/WUGw4EVscpy5drlA0aj4cOOvqz
WyODCHCtO3w+6r5/4hdYfxAqUwCGBpsW5hoYNSoTZ3fKAFyzsER19fK8XSbCxbrl
sM5NSZnhOyMdV4uEaKct6xwZn5+3scdt6a9tDdsYBOwS7DBYDxWeQCvWqZUxVOIZ
CXBi6NBWNd+5mIhHZtnevrbrL3fo9AxbWMgtvEY82tMw9KQNsVxuH51E65J1r9eX
PgC7n+VxQrIjWtoLRvjFrk+Y11zsXR9ZOgzA5LUF2stmUu1ghEzctDt7/MSsBtC9
ONPifu4S1lAaLHbNiWXSlLtyCeUCtDoPHjh55oGQQ6anYk0J2w67WCgXvBps8PKF
d6upeJkcSGQ90iQ5RBJFqIAoweuOjM28SDR7QEa0dI3JNv3l4S4aDDtQpDHiUZGZ
aZTwRCcIx0pMlhccf/iAKzIFlPvUFh8uHAhY+Fkmzq3lFL/l2hcEe6Pc5i4LJcnn
JcUxwfDolZFtStU6ic902V/1NRYv+PGz+8qxTkP1Cb3twcHNGr2mCSoEVeON+GQp
UjDEB/owxnC8gUr2oXWjhpvz2xNxz7gKqyVGv7Nofwuo8SjMSSTh2TPyto8nsaSQ
jhBXb/VNmgl7kubxW7aeP+vWm0DSfEUpU+XrOvb4Mv4jVHXUY2e7XxVwBM65DqCS
FtVdvgy5QOthdWvZujllBLpb9E9vD/MPI0Y+cCqDzxRcdZi2OP6BfRZsps5rEyR7
62HkWls2G0T32Jfn0ZuraK8CTtpD4VO24vfCl8K1X5NEWjBWRY9xnxMF0W/YlDoI
nGB74GjQVtyJedLL4A8A5L4jKWrStXaWzKTSCQ9Si3JNMEy743YhvYFFRYwk0y72
lQhLXpy0p6j2J0JEBWW9xpOb2KUDy31DzthHuDV6AY0I4nRh9ReoLVetXfRLmj6z
zcMjljiYtOJXPS6ygiLkNHVXmyE14fsCBDK0ceASBV4wBtHWFxpnmOpYQumqHp7F
4jEtx3NWj9g8KlKHvoiNsbDkeagUMuf6Y1Mxg14Q/SF1qNPi4tkqTuF8tWPfZX7N
D8K6MMUJkrw8KMrog5h7fjZDzQ1GCasONbEyLmv8SiPSeHP4rr9fwZxA2xchYG9R
43Y5BECVMs64zGNyBM9m/z4XafxUYYFUKwO+vCVEkh4f+ljLTUlyoHo12nU1oI1k
OAb6JdeEysK0ATGWB4VsO5m991hxx3r2UqAbtpJKRh5TgX2K6N5iSu2gY3QWVSaa
HjaMhTkzHhNwXgcKvIOy9Rooa1dDgryKifbj49ush/3GJJ0Z4ex4Awbx+0pP2Tsg
zfl5xLyWDpNQqqkhTbt7o/8hSe//m/D4+z2SvTLvXMmNXlPZrOZHfzX5qyGgeyqj
N++uvQuXrc5PFR/aiu+jBiYH9g76lpHrehWrnuRMR+u0Sh25Gamg6WexPLeDqGKM
/ANjT5bpsQEeIdt2kWireNHYIwUWSKBCyIGBjCens9Dgd5rDyFEVQc9nauABJWWB
LtbVo1Rqqr0QfDnUn4NQImhBDNZSlTTw11Ryn1QajbDJBO8nPfc9evZuC7RhcsqB
YB/WTNtQoPd/UMAcS2iL4LbMM4rZ1NWEv+VHxAy2JkCvF4M+eyjFK0IlsCVffZq6
/zRV3kE0RwZB1fgB9bNlyzbqguQcNWyYUk0JDYs5YU2p0OYvmDYw8MfccWKAk8Nl
bfLesGRxa0wQFt6Q6PGGQ5BCKR2oaO4zs5OrCfv3Hy4eO2Et2RY5uhjpMgsM5w8p
CCKTGOASRBZbOdriqOD1JrjjoNzP6iCtK2IcnYhir4Ms7hxkZ11L7d47RqgvXiNN
EFqRK6LMPP7MkyzRck3qtiLAuOCua19qBkLSfVBc1KPbKrBcxl4RyV6yN5xKiQgd
Y98B0i5p1tde47xiRlOPvwQFLxXltsVgDVBl5wAt4/qxv+zOUaiwtqs+W2pIJ2oU
Z/mGByaxw2snPFveLqWbVDXWqJZO3YaIWFKoRjAYDMnXyCnzdB2ZmTKddTFbncNt
rRR2fk0L55P8fHWrj2wKGfo6cgPtZiPBWt/nM/07D3hUCebXoSPhmH+ntmshKS+x
iKU48X2dr5LHye1GyiYDsHFdrsiUXbT1AlYfEHgILdOAB+bU37P0ZfNexw5y9OBb
SeqJm1Ox7vy03/5W29mTqKVzvt4jwRj0/LhrF98GGWExZCcRgeTmzHamvk0lnfZ/
7+XrrqMszNJ5zmtYr4zYoK3T/Pwce1Hf4RFrSBEVPRNBA760vYVOKr0wBr73b0Ii
38AvPi4mL0tmA4KxJMJt2eAwgKUuzhq0hHQlZo0xaRyiqJSEg8+ia3ncxcZLO5Ip
TCuxlfU1ll+i8XZiStqMO03Ebr1xcBubSujCXDmqBajSwXifeCc/rVNLbHcxHdre
wbmr+JNnQa24KW7Eb1C/8vycLkKifFNkn2NfIxNqzHEZqc13Fp5COzrqlf8VtJxF
2jfC3sPcdF7GOOApi6LSjogOXVfV8Ezhhmuvc5qS6R4/X/fvs0JeDcef4iK9neyC
BLGV5Y9evZhS0yGNbdfbZhr85wRtojEq9UWBGvEv2TrfUkFKzvDs5XdUI83ovtzM
DG3i+of9hjgAJzplTz2YIyOrOWlO5jJw4YnKGD0SMuh+7Y9SSm/eqE+0Dc5qDuCK
XzZoOI5fW1tao4OY9WNVCyUgS1I7Ek7Z7S/ebXsbwhDJOeeOtwHkkHrfwfqfF3G6
kBzOEDkpAn0rbaCN9TGM6ggabFjmdKrt7uM0z+xFCDogDSd84I9FrC+ur/el+UmN
XJl0znbvGjy1uuqOUbQqGBwYZmcFYEu7lBgCSjjuThjowiqwiugJgrstrdoZYHLS
miwyKcco8zwHD6e+bANVLKYh3MhuuWeLb4BRPvI+xkO3nrK092wIiyY7lz/J2HZs
J0j/H3hsnvHSK+tKWnflmaKZLoXOf6WUy6h46ykQMPBq4CZRxP/Eta3R/m2ndqll
PYd6gR+Sw4lilHGtfwtqWU5HBrFB5yfWPUuHCC+/mfQ6Ecy4TC0gW8hw/aTYEwRb
97ZE7tpAA5SHYHLUWKc2L/j4f2shnHiPD6ToR34guO83msMJf02ado3zi5P3anTz
UEILQYEwe/FQG58aVJwJZIPSBZFJLq4CV384452vnGI3BMytUI0CUDmlsV2LC2Ob
xD4mgzhXdDds/YHOVU9rsaNRFe5JfQyPBBbP8z7OwbX/RKNZwXk/RXzzIjiZ9FYp
ukLcdVhIJzykNym2EWugXrj7/zQ6lUMVHnNqUwLWPTEofLHRhpvynUPIynWWDnNa
UR0b1j9Ijc9AEhss+bBQApEIA181JIJqQ2rZj5SCdW0pd2rMOzOWjiO+ig9jIA2J
ARB/BoM/04MU7M3qpcVew2GmPJZi+em+O+QZAWw8KMZGUqCcaw9Kv63noDyqYyQM
jGMFpcCc88+kLZgVsSAW1IQccu+4roMC1WKfQX/Sl+Vpjum1RSy1PQhWHgq+JO63
p3dugPprAXfbzDSYP4uBB7Lcd8Va89cM8h1k6KVKNAtpYXnkxiPeGej2TKgjWsjM
9Sid5ThgPTvGV4+VL9LcaZ0BuTyRGinJ9Z4/ccSRVV53p0oZULQ9K/wlGDNecEBj
OaSSrFS+pouSq//NKSZy7ywQsp3hJSoSx5yVRj7thI0Qir5+W5Ij+9urY7eCj3LV
nIQ7hCzJcE/mqyZ96cHzzwYUNQDKXI5XG7sp7wvigRTW6muMm//f4a6jKfwKU2vP
MUEde95XaaWpDJKZD/OjDUhlckHUWg9q5quGa0W6G8YCBtVkFk1Zbv8f0IPWanz4
XNbA0idad3rc+Q/eLIXTqU55t/3fYO51QQpl8NLpHiqTh0xBrdrVr6G/CEh+vI7w
iHsl7Bm5ACqp0bCtMGyXkAIN3O75hH8HMGpBvG4SwNLoc40He+ECYwPok9B9mb7f
XIizENbMuziYdguQIk8H8mLb1CGo3j8Z1cekqYA8x2xS3iVitPlSD3TRjx+Hx/BE
FXtM5CS5yvXa4bgHkfYVmIGyFm42F1o8rdjww9bVBSuYiEdCyuRTqNNo5QdexV4g
gU0M0FT7q8s3wvXWtvslZi0zEnAw+CQ47jLEIaeLuIyGU1W+nBBAflpHIN5NJrfy
4565cyqTsnMv4K9X/3P1nyNyhn+5aOdtZD6G5S3ZEi5pLW1RcbCOyvDXiEpM9mK/
NCJT7rFbezoE98Wxak0WEosLpLRGM3fIOhlGQ7fYWDfVwV0k6qWp/Huzw7pRZfjG
UbbI9EOCWMkeO9OmEH2ZFQkBHpOOx5es+iZeWFPqm1P4gwn3SRTEJPYPU41TSxpC
A2+dhqYgceOo14rGhVErF6NriPtKxrr3ZFbqMEcT6VVLG6TJpSmACQme6VkaPtvW
UhCBAnfgBQYKYogyQNId3bZsTZEeAoEc1sXpuLSQNP66e9m1h2BhrcW3V1SN8j9i
k+KjuhwZyNknjWaNzB5oBJsdntGdeqRnS/veK/Yg2Pk9MVAAvW5i8NGfCpIfipV2
ED2LmQbLzF0/h7PRi2PnzGtqQNA/y8qt+oeyynDN7m9fIfKwhC9MeASB1mHO57Ai
kmFqGyx+Ot+JSDYGwG//9et+054dF4OYBvAfKOIyYQPdHwCQvUnErsNuys0c2yQ3
PZP8QWpzfkCpByHYHQXGS2j7I5q3bqA9MDCnw5z9d93kYIdeil56IvKND2wFa0O2
cp8nOJSbN1a18jO7lcSf2dI9TfUD2ZiU5SVfzjsV09nsDzbwYMev32qcg4C211YB
g/jhCeaZj+0UjKk1dtGRetPm49o1xLIe9llnQQntkylqtjBvZeh3Ddy0iLnHRl54
WvWrERKmzodDhN6tnHS+OnZBIidyA//PLlVeUjV1RV7wkAp+bdTfaxSL0CuzNObH
iOwuDhr1Maho9tgzlS5a2077u0UsegoITM/CrhG6hbRAYTg+Y/2qOZIU3Ncgwznn
CKMkPpItTA+lvPvQchu3YyLmenxUKwAoKfDlwZYIOEwdJv7irlxGr0TgomdAmGrk
n7gdBpI6rg5jRG2cD/fd/6tonnfboxSfGvrfAwpHXXSDg2oreBAUm3wJ756sWbVE
mDbI2LAPhy6dZRvXcnfeSKW191EbdY+rCp8KDGQcmLrNFxuZ6qJe0LPbvRc7fzRh
W3B/hqTKUP+byqzWpHPJM32jQqqHXrPyACNasLl3yRfmw6bAi59Chfea6xJV9Nvj
jq6sNUlE4k1rP2YgWvF7AfqC4XXKPr9DmcKXU04NvvlXAXpgfAasw4Ge1q8GoSL/
VKZuiP+b5/cDo+LQXmpK8JQievVsXmGqwqRBKQimLvTJNGBF4e+sCyeeK6CGvsTl
xu3jTqpIzU/TBqBACQ5A2JY257q6AQBfZ03pUTlwdqFuTzUVZqN4+1JD5XnMXnYS
87mQ9kUAGNgedgzkjPeAQPIIxH9rZH2rk3fEvP4rB7Ewv1tp/byaUFIyFTB0Wx4s
C9WeQwuWHQ3OqRrGKAr6p9JTlgizqsZ3/zbT+ZyJsGiOfM0W+Nz/bAzZsWZ8AQnn
kRh5UjTJVof1SiZgAiBEPQKhSv/AZa7CLeaPse1WbwOxhOzRTzTlSLG1PmQ7MCsS
hRb6UOvRYYvAVv7g9M6fYrSQlpkOVs4LwFngO1TTT2kONFEG1M1djXmjcbI6N93u
I7HcldYJ4meLCBgBExvc2wGfBMh0RBDnygeddVZ9ZIEp3zfjkhow6o7fRlvfppoY
LgeivwAf3zC8yz9pRz8W3nvlL6E5LVDRU1FcnP4GPWZp1KtZKI97USMFKe/jq6oK
b7Vj3G+tiWET39QQX9HV2XN3rekvDvpmG7qAyZFitbCMH4f+tQXNlj091v+qU1Tq
CYM+CPrkM3aGPdxOV6z/kLIDZnlqVKn/R/psJIdpoynNViSnt9e7nVkPSoV6s0u/
2+fpyc1LvfnfZjlc2ZK7xrVxBLID4XWfoP+gquWpFNaLQAX+WN6MVDNVPY7BkP3o
FNw4TieUH9pJcI+5mQLSo+8B2c135z1cW4nFeOLooPPqpVEmiSbjtdWv0BgoBKcU
+53WlrsWJk/LwMNtQP2zvWau+TetetqdOfGz1ohltRmBJa3xO9b4pPsTkDPlmdDV
X7kLPKzMRN2DI0gSxp3RzPe/t1xXOVtsJTs5Lb0FE5hO/0fxbffde/vimDY2ZiFu
KuHpB+zMaE6D4ZJ2i2Y3S1QbuHOlnBgcjc6BOWsy4SXmY0StoEIVnMaeaO1UPegZ
wC2aqNBu+Bs5s1RJwS9+k26K1XLczJpe2/hyzjzzsnfPWYu41vvtdyMIiEVlIkZs
ORBzUG3AsF2JE34I4A2TF3ogoS7JHk4oZ39W6/t08RfLgVtLvv8KgUpQICPJ5vO0
acNpCnKEJAgc87inYvnXXlk8RitaaDIc9hHptKLp2d3rKCgntM1zdWCiGi8JSjQL
kZvD7l0XafvIVPS6DYxsAW0nG5iHZv2jq0hULasGAqKPQ1D0Ifwevkk87e8ecmtf
psTTG9wGGpTX5IMRa/NkNPWmQMvyuTLrMkaGbofQaxr9JN/DD0LDm8+sbv7UpPDN
9EdlfnQUQO9zfR+E/VRHcV3gJNkU8h5uQzfc0/PcpYdF/LNEx7TZK1tX3dzyh+BX
um0XhY0sFjg/74TkPNDYGxo1Db0MX4tFUehXvtDcsIjPRqlcjEGAUzY9VX9ZuYM/
iuyWS9HiR1ARIkeRm8H4wPKXo9NpyzRtdQ8pipE+qhUdzyFK9Z98eiTAjX5ZtAT4
yoOlKvo4SyJbE/pefx+7osE03T9wgv6iXrtRiuCCJcUJYZja+EIEOmXTXDuYEVNp
5Uy3IdkSl+VV9QUrdo+hB+ksVWAYiTehMAFhbQqcazhZVNnxwFY9UHxpIvaug3GG
mkixs37sT9COP8K1U7Dq52tEDwgPq5L1uOunpPXRGaWo7Icijtgin/RjP3/Z7/Aw
2pj3x0xKO/EotRtq6Zu4YJDRc6Pd8ALLr/tQmAEkpxyPMMHXWM1lHBLfaAoPwipX
pMVKrc4BtJ8kHEXSa8GVLgIXS0Q+FKFP0xa6zMDgYCGIZYMsNCoUeAwtK3ENUf/V
CQzMWgsy9RhyKIZBia3NcjwxQUtLI+o1QHngbBWBqI1utIgECLmB3p7be2vqoeOu
hr0fXFj95MnssKAlewtsAqfinEUFr4eg1Am2OVSUm249aMe3x0MjOmiuYNXzV3Ft
bY74ITad+H+giVsxScS8Lacll49ymT+BYTq6N3O2DQR/7JCnOqUbn6FswBDVzrGw
dSFV5LUEpQwwtvAon+Iia6K/mpCGKdu+Gl2riLY6xLcYdBFRIw9vsjFCqPEwOpXl
6S2w6A+cmD3TIIvcu4r51X5mXJCv73F7HXt5rZm4Eh1ZfuGGF5pu9GDT2s1Gjnh8
9syeOMIRzBWV9kNTrskB4bh6ryQMXIk1l0d0I28P0guWUoKyTQ9Kk6nzZvzSWGh/
RhNwR+1SU4T74Amk5OtWSOUioY/Y2UVaw6sKYQu6TofSlrYaxCl+MsiZcSrkLJMf
tUkl0phfAiyMcF9hlRRL/V2n+P7VixRTcnjDc6uDiw9SGD7uHsi+4TaNSojdtxF1
s7JbtuJa1gA1sLUbhzY+m/mSWvQ5SjgSTRa8K/DxKf4PXIwrOZNg4JxTIKT8eqnv
Ew4DmsX5lVUWF/lsrha8L7n/e+IO1x9Syz0LadRuKdCcEIah2/oDZqRjPg/pLOpr
dLfbdY2qoIQ/3A6ljOF4WQjIPwbBLby0D14q0S6nn11a1oPTgXGZyrwjxsPivwNe
6V8Fe8Nz3jiuXCFqfBAPGNET9wHK54vpxpGl4CNEpUoYYCMBhcULPS7GpSLs/aRH
QzBhMvOkM97NCKpJHYeDUERSX/hkwcJlMjJZBLRObtMzcqXw/cdj/7Qny01xFXiF
G9vXptOz7UFsiPs//EpTcTpL8UXWx9PXpNWtNYDYB55HaF/PhdILVY60jnFqV4sZ
M2f/MlUU9QLYW/Sm1IT1kvf281N86ZhhvESSA9uANmjemce9qBeNH6poJkmst0PP
qO7pf1qlrkWkFwoczSwISGoHiC+YWhbBT3+S+fpDKBd8sEsD76IL3IkFXEPQav8j
RLRhfWovqNx/hPzs5/NDe6xcihk8oMb7Q3BED6KoV4D1sA3LJAPgRDexSs1CufIp
U92IgPXTvQYMzGuS1fuzx1cM06SMNmSNUNpKPAF8vrEWmZDagOthHBNDVACFBiRj
SmqDDXzdGR+BKIvXPcpYGsskm48UI33hzeMqtt339hDmgiiZvOUTngOwLTDvumcp
duanVmwmdP5Mria/eT8Zd990nVSd6vw6DHqkKSQZFyB3HfEGDOdlDIbBW/2gPaVt
Uz6ytffQKiWcDGw/VLVi81qebGjAMtiy9KHiBeip8s+PkFzWs55CoxPJ6ZSQnXJe
MgXz4Pb/UohPFJFbVfyloaK+8LBPqyDI2pJBHBf1ywwZT8MPhCqgo9RuLsHmUXyR
E2FXhWJJpIraDq/4E9rrU3G/Upgd1TQdJiYvZ+1uS6ZZgOUoxQLZ+S3KMBQlAHku
9sxuq52AnFvgc8l65kTwCohTscnAgNILqjw6Dy2+LU4jGRnv6amPKXJdn4vsz2d9
RylAghMYyTuCNGa7iiCjXvDpRSGnaSAmHU/fYxmtRBB4e5GeBHOBeu82gS5yZmaZ
i+8KOhGQ9wplDnVphm0RxI1d1lhvYC04upeJv2PfBWqqkkLVOgKBWHIRU2D1vB55
7qL4Bj42kqXzxEQf8uP/eLFpA+InGf5go57VVNBcVUykHSWU/thsGL/wpoHbf9cm
mBWIQhbmthChvPSv8oS6LporttYOMSxPSxg3GW4tUEhXjcb98U3mS4nAlmLAVfOt
rE8efat50njMjDSKrmDonLIsZR2IlRn2sWr+x3uss0O8lZb3uMv9GPDRfNcJTGCF
j9mhIyqEF5oiQCuvgXViBjNfbqGMNtxcqc9PBaUJFq3vc1YtY6lQUTJzM5eDc+Sf
drPaElZS8F5SpQhmCGVgdWDjUtvs3Bt5ptbWMRKsp9IKk58ZiQi5ehBNjQSL9LeU
uOkI/eig4vNFdnkYYi5D9f/+nbkJHbEiGb2V21gjMQzG5h5NMTgp1TrjN3pv0nsz
VzeDsLULeirXdRsQJXPmarkpPDyGrWghdnqiiNkthUFLPc2JHeCM37lQmO9rBAyg
vjBzgYsvX/1eWjQWJZr/lw1qHWp0D3mtwRuCJBIfXQbxQqx4lOa5Po9YhKhqFw6Y
Eax0RFlw77wM3UbwAtxjIZb3LV/7JL/2P562IUaSuHo+BfCUFG+4xWXk1EnWLnNi
isb/ZjuHAjvpPjxK/E4gXzSoIgbONWYczoNdL0bsTQIQIa4JDVYhfAB1EY5EnBuF
LRhioNTSu6t8JAaDXviVIVgJVHhoKpQMtL7+nEpDfm9e1mOGCltyl4hw+Yj8/8bg
/ZYo2B8IUk/kAFcC0tTRTc+wYDparpFc2lDMThfbORcagjVZY2fBbt8Xm6mbTLOO
TmS8SDLgL0Aibqb3PrjlwwBTW+RniZFrpD/TBYe5wsPao9Bnuz5DAAShkrJcyj0k
jUDScQ/k6KcrVlLkap3BEo+hxAW8aSD8WQIixgcqVyLIUO0nsX8OEZTJqtN7v+/A
DqUDXWmDEwZyg2v6E0tFgh2vNkESTP1eMUrqps7FTBe9clxg14MPIi0QexEtZgrO
czszMoxVFn828nd+G6RO1SZwtpA/jKpwbtK/0FLIFBOF7twAk7UMTBpuxOxZvKa0
00BpF8Ud+LFZA9aukAVG/2bqdfT7vPulOuLlLHFm+Y0+hLeuZPxclRlxONpr8mAM
2d4Smppe5cjjReWwFJFgTqM4CQhppgTvVgXyXPZRVfVhzwP9jwZ1QFu7MAwGjSXq
EK6X+1XDnZQM9v01c3bPEcixAVCSLOvWYqx4itShTd771k0J1NpO73FwypMhBeuR
q9ViIxMrx8XE0o+2dZfYW1hvisFZbR+NIavzGRL1eKBxHX57dFzHW+Uk7pmRL11v
WSiDZffO5TUh9PpbyP8Td25qkFTbRZI3f1a2o/wWcshstWxZA6kjYBsBJP4VoDBJ
FiVQkSAwvJcvOi4VhNFNQZuh9nR/1qCb43LWSSRuvSzsfhIdZOR0wRNcDagWi8Ez
l+xx40UfU4v6l5H/+RhWsZQMmE2+VK/uz10Qw1UOXcldPZZpFOmH9jdJjFZhQOgE
/RZwKssVT+HACBKytBV/+PSSQKz9VVLyW38V+mN8AVZFNEC5NWNb2v6qFEILHkze
rGp6Fz1iVIk5YX6juEpR3h+ioyu5/NPj6zHtPi+oOaIICZNtvhlHx65M7TSvZyeU
dnpghMH1W5nr3SIUcXvIxn9k/YbtchuL4yiLSV1KDn43y8Mj4jAGewE69Alkx0jd
/bq5EoSY5BCv19bxxkqo8ApWynsGigoO2aocLyrf17J4fUdaZpoxOCLBTNlDlXUj
pLGa/Ad+LEup55xFZ6SiR5xlAbbOfqNuNJHkHofZAPXOIZhLJCcrcPJpqLp6IE/5
81owcBwzCuktVQkpiIgDXxKkiiF52K7t2JMOfOiTH4nQFJDTlUioXT6id3XfPqTX
qXnYWilH3gV2OEQ14zWPT0LgL7McaEZa+KTU0qaKFxXHw3ADx3Rn7g+jKMh+yFBW
q6ZEeDnYRdDx/f2IVw1QTsbE+vSoPFeMKQN7rf19CUF33tu4wa3CS+Fg1FKk9kZb
eo2jPK/3556ytvguJekLzVaBnkJA/iXli7eGAx42tszYDKWD5gpJeHOEbDxZn0oz
S/+WK7tvJ5W+Jx+VxxXzs5guoZHSMrM04ExGh8dhWOb0hsmNQq14eYblXhymLa7Z
xyK9OfsDDqrafZvUi5/A8Y4Hay+T+mCILGUoVXHmwIGhGpWHbj4F5QQ519bSOSOD
hvelL1NDmX09obu20AbbPBf1iWVU5O4Xz1IL8F1Cu2oFcIWB3lhSYTvKQHWJE382
ZL7YcieOpnkIV5h6C6loD6ih45s+qi4ya45Y5MZvj+VMnp2CaTgS/fnjOeeGkFgw
StGKf8fin0FyOc3PYMjECQWwSkJIN5aONlhKp6EtGHxY8sY1FBIg7e0deLk1jdJM
D//K4YYEWq2An4gQZi2RP7CllFVJW15WHkNm1IavXOH1QjFsWBYLoyN/WZn3vulC
l9FK+7mmccMovfmAfmfKzQ7ViuDdWRY7Yktt/m9tqx7TmT7Oc6CcSAu2j7tqVbmE
0CPSemK6QyIPEUjlwt1zG837A8LSYyFCpiBrshEeDLukcxH1hZVj9ipTDeYHcvgV
wLl7sAe8rw65gWbwKnG84nU0iRS5I+lbVvFwc7fNJfVe8Dxmqp2iPSVkB7NvCqJn
sgfdkfA/HQVrkYEm3xz7BZYQw1gWENvMBcqKiBHaxwKF7FGKGjiYzEt1MgV5a72u
2IkDpYTLE5DK7YgJxdhwkwNM8vyDeCsKtwreGZ5iq7V2NFNk8SaNPs7PoaRe9ahg
d0hjJ3GyU7bro/dJqKunzhdrZ4l3zgi8vWXuah7f3U1UpFL2h/KL9MiAU/34E9Yn
30MfQ+g60bUcdot1FDL4NcM6lxOWoCclQECN39n9HGYlUWABCMqVK9e991GRL3zz
2T9ov1+eF58pK29F6ttYx8s9mg6W7iOCn7Q7GymqFIDhrid5VjrONLPiWX/B0PxH
OzRQQmGV37bOK08KHWNYIeYUxR1gPX5iEabu7YJOSyXAHUyke2BQJ6WpQb+aAogc
aOGwWdAeLV+ADRpPLmy1odFn5wHqiIQPizfrZSG6ZQ+8JA6TXiFvvu7Ul/U59a0f
5zpYDwXHKJbu14WSKigIjMzvPBYSC2qiONEQEdwAkCdXfGtWrTxqbaHdB9l7597u
hZwDnR1hnbFam5mA2W6QU2hHy9D4RScuuv39uzPcSIz6XyCZNXuC2aW88HNBnrhl
pOhSaQd+M5FXieYTATcHU+MUevCIyjsWyozf807ooaj2zGNXUBYWvxH2ZYET4p6a
vAi0gVOvG8OxRclA57DaKt5plY5tWUTF8Lcec82qEiblVBE8T5Kbkt5aMPJjcbTh
vHOvfFyHduszD6dUIwpq1F3POkmg9ABVnIE43rOykqWIU2icJnTNmDNlDYFmohC+
m/BzoN0lW3ou/dQaSGdh+GtUT/zIafx/KU9BA7GcwbZ9HR2siIzPd7jxYtkgHBDu
rKyJ/m+cSwgdf/9aZyvGZTyDKW5Bl2udFBlho28vipiO+cuSVpB3KciuATVxnhqN
HdURa3XZRBeDLWHcxD/7N2TIlqzMkostFe37yFv+GAn7XwSepl/uxi1sTycrOtBI
1xAppkvqRcUcia8Z0N6E9flX56D26KD6EYxEpKYrHLvD1M+h8CN7d+zwp/rd6vrH
fDsxUOnpeJ5woVCqyNo990bVLPVVttsLwldCmC0x36jlSf71dlxaac6ARQHGdm98
ftiM2j1Xs7AYaPvULemutgkADj2v0Ehrh5hPJrJOBDF/c4Ap8cWd/yTitrBFS1Xj
Rrk6eyV1yXhwijyPrMNDRxgAJIH7dUk2/qwt+qpa6Q1S8vCICIweDcqtSNhw0D7h
dzB+pvy0OUrUx9KgR+CRYZ5yhIVdwwo6ggmJnpZfjhWJjxwmWRaKOLNgnTNo6vpg
OXKzpMMAxPSdM3tuS867GKMlrIcqv0ilePLSWzfd0JhuaSosJMIdfYUQidnLWFzM
Hy3yyHnqTNNNsN0/Pu3GO37Z2gkEqm0qyFkqBeJ888xWrAReBDz+Kn/tAhK4b8zJ
R/wfRfMT2OpqDwGZ1qBRpbWDKbZU67PvTRvZ6X4u1/YNxYehNB6x/gdb2jY3cGqA
oB0eNF80F9DMoXWvAELtOfSzVhpHSCc7I4FeaRG1EfP/kBtJaOaklVg5cmItJU4d
60UT5OF9xGKlWzfsn4Mea93Q+913E1rTvH/rITYghYTQl2KvPfmqMLms57kXCGbl
otOPHSf9gz8t2VNFCxcECTsjkszj8yVwvVoon5tPGXULzArydR5ldUy5ZYX1WmBm
wfk2Sxgm03JSz83iDqg3MEtS3M6kO4FkDSkD5Rj4AQwf+YIr9L5Q0xkdV29ThXZr
n68cX9xqZH6J8fhnVQ8bxkxPXjsGKt4qapkOfZBKO0ZH6mP1x5SaPRqOZJb3Vxat
8D1KDZcenltGcD7ab24528I0REROepn/FU+iBKskFaiEA94eA7FKnNl/Z/Q3kujy
WG7xLAVFoLGqFAtmI9Za+rNcIoEDEYHkbxa5wCvtjwvA7meX9d4mFbuMM9hTj7fs
T6K1ilCBekQ3g7p0ztVhWV1Iltvat55Tg3p6OTl1ENhkDLWwrbdRMUCL6+RkCFeQ
V1QqLp+c4sfsmq/a4ZSWsNCtxqOQ6YwGDnlHLaCgiIfGq0vVNahozSdHk2U7jxeX
4H9wSjtHqBMr/1Z1NMmNE5KwwM0HSIR5PFF4VzewfLTgTGjKdCZStbXIGL6P1yFj
P9nHCuRAr4O84UWAEa7SLOTf5+SV6FKGL+RyDEW/hLVRIBgEq0806DVz6oRJILKh
AAIaelkojVA0fTU3THkVhnBXLPM/uK7/vuIAoYxIT9tV3xqpvNGhkPo6Cyt1rHM7
/+KLlEBf15G3pZHk410zbkmZP2dJqoR+K2mIhf4YzLvOiiTCUsmK0kSRZLqUBKCX
c7HY3A+J0os417xQGvMtA/k+V4OISS/Zj8evra4HS4y43TFV/utvWrwqL2xuUv0G
g9MPlYYtCNwD5UmLmNcjcionNpqjGEkbpFD3k28kwv5VUHwSG97U9SWsCpHEJLtT
bR/NXHOpHYhD+Ny3oYT7rEQMniWfbbDpcwiiIyeT3YzBhnsTZywcoPWc6cuJQpGC
8aoHqIWIC8gzx1yO1DOYUa/Ui/TVrVS/0SQxIIvBFFgmXnDIBXF5wlntrRte/zL0
wTcUjMzaNJ6hs8AqoAdCD+XWbQuhejw7b1LABZVGtwBrANC6dUDrO8o1WhDxeQXI
upolm7WAa+UHUfkJNlPp1VugL/vouQGb8K5u/5zYYXFRNYxdhOBBAXBBjBfS8Qmr
PWOhinRNlvsap+ES6R+T0SVS/ZwSC5qVg++imP/L6xdYJAW0wugBYpIZdFgqyk5M
c5SLHhjohCSq/opyvuuX9rkV2MKhVb2YUvoq8VFHtidV+N+X2smPfI80kzn9BLEK
j9IEkaCwOeEk2B6qhPgqL5Qc54ucQOdu5cygzjvgoeJQwHK3Tft7WwHZdcWw9Hdp
fqFcQnHagxgitNRJDS6JrWmU4U16gpD2euDvZYtrEONvDnkYDRmDYOkYgpVwc04Q
uJdNxdV4cK8GXTeR46WIwgMDVEJs1//cS9oGNe083O18bbsVaQDd9jCAAkXnEl02
qW+AaapHdZho5WWkZUjG2jXp00fu1ffHc5ZUSlza2H5I4tlLQ/S7ZvRTLCi9dIfh
yI+L898pqX8OuNam+1oUhFo/qbb3flFFKVd/OxhbPe8StKOZH82G8cuDL14bhx8F
8FYD1YqgtqP1u0t5QpI/JS1ycOcAXFW58EXte8pa+KnJZrqIhuFNp7dCUBT+EpKd
5bjbSLLCchKxCrqTdm7XILF5yee08UWWX5vUAiVXDGj93SEJ3TaV2XY/VVDKEkHr
0um6+0cHS9k9SUEI9XGYOlthaII6NEOzI/FBRaJChWRgL444voqsN3UpgXvgY2ig
atCgRmQpxtE3fFGplX05DlXAyNX6bz5VF2MdhSxqIxbTZiIfpDULHf5fzLzgwbc+
nwRI9hADtwFLex4MCgSDwCPSEhR/xaQx3ZkTwOJPftgCG7j30sqL4Vwzdk8d/cB0
ivDDVVxjDCLE57TkB1++27/ILNehgVmfyJJum4RovWuZAKF7/AN/J7OdSp5uJQc3
/LEcHKc6f+/RBIvty9FzKw1owXpwpz04nUAoAJqxJ5zYzapaOnzew4gL2r+kbplY
B2HDzcsVXpV6kFHSMctcBtQRNPN7isAYxr6aIl228GdmxLyeqzu0Ul4fHDSrEJE2
I2l2en1vf3nMFqYnqRmmPXFXa8CeuekJxra1x1fPSt5mhWJa+3gHSfMKTaSjL0sp
UUtxQ0RloxtLCNPMBJNyxuHIS9axw91lA2dlBEGRSvkzBZCHBjnrv0DkF7R39p7r
l1G9aL1C4DwMQE/Z9DevjqnEk5uh/anXvwNl4DJNoCYpNo/rAeSQDR88SaZd4NAl
lQNZ8Hdq+qD/M0Ol/tpmtXP2LAva7VfGXLs7Rq3nxlAfM0uWf5B00dBPlDf61Cwk
klSQOvJ74h/kMh/wF3+Qzo7LrXYMG/7ghQrk94I096P5qLVIbWnt/5HYLjr9slI+
hghsFlfbj9/ndjbqONGb6OJHM5CXR6o+9arYZ7oWO9H8jTgSC3YenBgeENpsuWZ8
Gy27sUuDkCEy0ny8/74iNEa7Pqps3s0gb9EJU0VgTaliUp5OOSJX0uFMBSBW8PyH
x1+roxpWqWAiy6OXVV5CZpjtxtgNgTJ9mKyq070fvQqOlbBvye0kdZOqBrVsofRB
5CkSwnylcnqbJ68mcZd8DhCPtJc9LSKKM8SrCBgVgV28FvekpVzfGJ/taFGlBJVX
wLpIRLsYSHbE+AuifIbE8Fnpi8VEgHcvaqeLO6nI1vUZefTJ+IdGicO0aDauPYQj
M98VS2+6BMXEErS5EoQu5frw/fO03I4WE1aclAYPP5bfnP4Mmunaf8m9jT65ocIC
w+E7g07soxaVgXB06ZJfbWWQWH7Nu0INbURl4L0uQv3Pyr0ZsrG5PmChamXIWoef
nL10dYP10Y1FguqD8n5FA6jduHKVqNKEpIYH0NClMDmvKLSPSIkpnAMPfY8tase5
8R2sglOtbjHNfeTA02ddr7skQDGURCrzYyAXudCKUBW8oERGq+BUll02pRilclK1
+VNIsTQGK8Zqwc7jbmnXeQ0JHD/V9P8yKAKfPItZVNed2OLsR3uJ9vyrHweZX7MQ
GjY32uXuk502DHHX6b80dQ7ewT7m70Oa6KY+cs5zgwhHgcC7WC2nOfMlf5Z9/Iad
g7d1ifP7toOEnN3OD4dRKZ2ZBBwQxV609kGaEU2eNKUFY0Soild5K20Y+NvHz0Nb
2w7XU4zgH2QXazrHghMa+gUf1kkRC+L7iZecZSE5Z3q7ORWYD+3SviEcQBrWAYjB
aAG9ZQY/08szNXBKpgLQBGX6kH/TO+AAQg64en3rGcr4rzhD8Ycm8TWLshE/rqBa
ojDElpEbMO1E3J6r87THaPJHUjWo512fyQ1EKQ8N48/UVv7myMcXFItg5R3YI6MF
PX0qXRce5eSjR5cM1E+2j1CMEaOFVKUe0xCNhxpqtIYy/2JRYFTR6kQlCSm6K2ok
Vs81fWYooFC96gTbBVO9+afjzdbX7DvO3MJKpF+yC1sMf8Fn2GzB+uQkccD6Y6z7
yuMwhP3UuuqPqloFAYqBGNpJAX19ZyWW42P9js4/m9iasK2u/kh4vOsHhCaR4pQ1
mVfwdQpSd0CCB+pU4MuuMfcNx1+0sRv/62eH1Sm0MS6qwxE2RQFHFLTb/o2Be9bA
wEO3ZQvKQR60VjM3hCpMhVFutqgVokIcRJLI81weT4IzjyGPeAZsfEjtrk8B3Lp4
CiSZvacT0cfyLQiaXZwCpFZlekvcaHFSjErkFGYU18YBY44HcEiRU3Qn5KA2MoxX
4cEI7yvhQEU/2AdR6Yd+GKT/l+QCewrAdVzYrdxzBQH0WVSphJhFZee/eyYpdp+9
G3neffXAyU0ejFtSe5ig+a9/UbqRCZlrhrt5FmSWHEknHV/PEHhaDUGPBjYVVJUL
PSyFKPWWv512T1uYaC33vCwKOgSg4zCvDo/wdHQUVg3bMMQosCBZIzl9ClWu8qK2
Tbou9nkgsV0pHxMl9lnKgvY/KPSXiKhj1qTWa4ntw52mVL/TUB9X6nGTrbAxYw0j
6a+A//qy+lqImvkq8+/g5Y0h8lgykAwV6bX918LT2LHG7jGiLbbNFCWJSKvajDE/
BFNc6CUvIm9tr1+7P0RhOxnpv8wC2WQhcrdhi9xXDA3NCwmS+DxY8kIz1aiLgy7w
LYcGb6mIVBqQv8s1nlK+sz8BFuVcgCefJ9juvQfyj60o+Wf95mfJFQiPr/VaFo2b
AkTgFaAvQJfBtjT2qrAFfZ2jYAQv1bdov00UJXEdInw70HBaAS9V4bUw96UrTLaP
qIluLIcP7KH38GvVq8srQCewA9s0q7h5oDyeuwbtEihqynq57nlqtpViJVVNDMub
N+PFaddfDIYAPgKEOZY8x4rsB35JJpHd/ZkDSkcAdUIIDTeCWybtOd2ypy0HbSYU
zoOUTGh95GDAIJSkTHquil0nNFPgPno9588QU7ttWwzaxIMEl/mufmCeHAFwTgkC
gubdyAHrTyntKDmTcrR7p3ATXLCg0swzgiE3Y/vjxPjS+t6ZTf0OvhhneM7JM/xJ
onm7dM76njNioxPvwg+nK0XNgL2uDEJvD611fY5nWnV2LVKLBQmgWeBbkpaM2Y+c
XCYSGClUZ/STt5G437fOGeorpJIuptaTVKGcwuDImqzf49fETJBSKXov496ecrP3
X7Ab/aWVIHb5oQEhLfgmkttF6LZ1D/NBd4ztHxUQTopOg+2TLjRJMJ5ChswegeTh
Jc0kVQdsv2DxF88W9fM3+seONkY8+JKMCDszaXjJi5k/Hwjh1hwBLPnYbEO7GsW/
AVuZ3XmRG6dRbBTOZjinXBDhkRoLVUgekcQ4SpMnxAl970HnPgd2MJACxevgbQPG
/rU0bdcTa2ieDBNZ/+dNcPxmiU05Q6lSOccBgqBU8eVWWxgDc0M2OUlqymX2pi9w
kA1XRAcCKf9OPDuWWzUcF4/HuJNrOsC9R79XgJGsIl2meyeRp90PhcewbotrzXVa
eAcbs6VlU91yNcQHS31hWXy/1kvgCL4p654n/YW6l/BlAStWvJR4r4Fjl5PFNVdw
cgSA31DADIxy9YCMRXp57wS6PL36FZX6BjkBMZcGzk+QSjn/Hzz8Q6np095LHGBV
WZ9lc0YF36WNyDnOmBs1FBDW17Xtl5tktwyw7KwibkFR+qmSLn/YR55L0Vp3WCoR
zLFqHqZTtg1W2rH1Qa3kawRKhZ6sHqVcB2rFJkIfivrykKSI3UuYlojs9rNIwwUE
teGbANA5HoOdoTYRWwB/s94hOGpih96JmdpPxilw2TpNg68ISAJtODOJUscDCmtg
1BDH7EFQkbVlTEqHsB3Q198QIll6sLyfWlHrhjCT4PEkxCcQGeP8s4Wq9Z0pn4UZ
XTsyTMCHYyX7t1ZP94yS4zOT01oi/LC0qaeJQCfhtwdlFHBtJYlbwOtQZS+Yafpj
PbxdFVsuYMJvem9E0sL+e8wIyk9Ao4yIS07IGAnc1SrRJLMZKUkB1xyKBloYnKk0
GX19etlJhcsyajbGn3qlOGNzHqY9VWIXUvu44UM9CSu8Bx0vkzw6thA78mFJU7l5
TqnBQXzvYwfnTvavtPFM2OJVZ4aaYjenQF8twYA14cO6tKwlgwDtI/CYQ+kA3IPB
a49H3+apzIGVW6M5aEnqCEY6hrlcWWp3X7mM8gQc8igsQBU20bzYJ3dFSn39MdYG
R7R+T7vc9IdhDodY96TymDMUsyad452yZOtqBPy7B9Sy76k1IqtDJ+HhRXfYp0Cr
xF0JVn3v4bgPz0WiD/CpjcsdP08F+jt9YdXnnu6EjUpannDITTkOPMw4luXpV74O
OTn16PbgpIdnJLLGhsM0gGjAvulEh78j15rZ+diqsN5XiDIhCIExuW9CGuVy1eJe
xcmCzqyh2EddfA95u1Gm3/GV1PZRShehviIIrWA8KmolwR0YY8LO9dGOhok8WuhL
OZeM2TSDJcJne2h92mHCZJaAUAFB4iocUpc1LhxaovV9c3pqtfKPKfP0B75/nVoV
WHXCFSE2VtBv+ULkKccZKo2pRCVPMX6eGtXVEm8VqbKJknp5J8N74bYeU0fa3O7S
yhvSIejIMhtucxYwVuurkCY3B7no99UIFWfi7cUKsdr36bA7NdyS2386e5UIQ5Jk
0mzrl8XAU5GPtmEP7gOCActjpZIQju/1nt7EylyBtTih0GLasz3SHy/kdjToWRza
Nw4GHg003MKMlI0YHukeMEBEuNRQQFlsyHAavWDtMXJULGccD0Lfw1d5eeaQQmrD
A25gWw/yoENFdMt6pQ7Ii7DB0fwp/y7axOVM4kqNJ8djRWQywE98iAebYzCs6fZm
3ZynKDsIIadCfqegG0Iv+rqP/Kx0eaPMmzhmpho0kkEewI8VHNjiPZead687v4Cy
r8UQ5zvgmBf3zTagNjsHVMuqDPGWkNSxzgFiR+gApAd/SJcBMXy6+GbPDIflzygx
nvCeWVC+pr04nzPuD2eVuuNlaogzUD8XGUVJ973Us/6Oe+8pfJ67YGsjSuTDMOZw
1onAEo7ag33M7F0mRE6QpfxqqhvRXCGXWF/ZCAJhX1UQfVyu0VK5/GsNn6rfWafv
iPsbKTuBk62xaJOj/D+qRifCQHrVW7cZjnTVyMwTabCe5VQlBZ8p9xXvgg1nXzpu
qmUDUirAlsXEiih4bJGic8aqKT7X6vfqo1Q+S/qHX881q8G+AfWtuq9FsXh62AqA
PRgMxpazBpyqI3SOao18PA1D5RPaM6sfvA6l1h9Y8u5D4zdLrlhypoBUCq47tPLI
bHf3tFVKFsO466H7KHGdxx19/u1FzU/V/Qy+2JmMU+Y8tmFFviYBw+aGBod0waq5
VzZ0bxFvmDE0H46eMyMhiS3anP8hTAPqIxj8tb8GjHUReNXIXnLbiPe9B+DWMrMS
A3met3SNg0uSYuqhGbG0GXZ0eAEkLqIyBWYt1UblhcZzOTgwRDJJNcESB5eS8C4h
K2FZdw01KI7AwsY/pGlJ0u2z+JShj7eXMgOgnQaAXsPevd6HHmZ7uKNcDqjX2SMl
rSOhzssKTcrmhbKc/d610IRgmX0kqxIXEYhMnO5QJfWqEtGSFtRGrXaNAD9n6Dn3
1Akqz+Qd75D3VA7U4C6Zgv0Jr4f+EfDdyRYSSRKBk+700SHwV/PPE0Jv5zBvdjIh
rS13uGMtHTgAj3Men6q75iJzi/3UbV3FRozQuKuD5qwtBMOycmk8Z5sK3QKbCRIb
6ENvYUzUKivlrQUzbf82wAGIyw7Utg/NLSWcSEyUaDvdcUiWMnhq6dHUpZIOHZGV
V5h0wOYmIbQ45bYGMiOCBNNCYRzwR5sFBOvudykXkEGyxSkSp4YDCFVwmfBCOmQ1
Un9uDrsiPOii9iX4fb0GRcYEl9DKqvH0As4oeHU5Upe+pxvH28OYDJ5JfhfJSfLO
gTWKE7kuBYirJRMNGMzD9byWeRSS9roAjmJa4qh85Y6EYVnAqUBey46yunIU6eEz
K+n1rS7g0EA2murNWxXwTdcS9ilIEacjTZaGvmZ9FLffwk5Bb+3sub/L8QtmnVKU
rdselQggN8NT83yefStT87h56tkIAIE9fKNgDqc165D3I8a6zNYjC2rnKQIMjX9l
shTv337/nqTUeeNStoNGP+VZSeqhWuBgfhEh+VG/hOhpz6JnGRoajw+zI/TMaqYD
OkqyshJkAKwsviE173ORYLjFtJcmD6hUmMhd7/DYQdcLWVcmcRFc6xO8Ns9qbzG6
LHPP0DQ9+B0DiHYLsH0AkrCckTt7tEGa0284C2fc4nk5AQFy6A7ouBicXmsbJ6nq
dybwOF8RW+HipKF/XFn0mFvTLfNetfqfGfgZu0pTRC4kD8oc82e/Gur3AhUQ7lPO
/+uwAdnccfhf2ZYOgxxBs4kOIVpeSpTSoj+aqpZjUSBcJ+dLAQ4uNT9jFGcsLFir
AXle191mpcEGPsfb1XgcXWJG/4+JKgSW6NmKUif+K/dTzS5ewrtcYQyiajMtYEUA
f6NQOyRc8ohGcTIurggX0yeJoc07RUbNZzmm3m+6tw/GubeuZ+/fLMCEc6u7eEMr
JrfNTVJPP/USrP3xb8VnkHupBVloA9F6VRfimD1iJWg9/VPbnvDSBo0pF/3mHoBz
C7M8snWPtaPv+KNVinBI5roWlMh1SNBfffFmA04Mm3i3WkQ1zcU3M32a6LjgvNk7
35laauO+LTJgzaaLZK1XvUDEbnDxYQB71TjmqsNrVgkw5HTkqR30QgwzuNLopADL
h4kx/TVgRGXI0JIt6TcGz/Zkk/Y89JL5G/ujVYjUJYC/I5Dmi76yMxwU4mF/TPS/
6ZSq9rtGurxyqisYKVpEfFR+S7VWRV7R1qtifbfBOJXma/cpXvjNZf5hI3Glrrlf
PaY5T9i6ZTROd0lJe5uBNleW4VJCI/qUx6mNLbJNhvk1kRQuAE8bE5IaEHboJjwF
6lAzv0R5NNHBSgQFS8qP+POVZBvE1q1e8wBaKn0FpL/0+wRlgzY2BD4qk5pO9b/O
/MrESir8RH7qFO/d2fLqFYWzJagElN0a5X5nIF1DZu4OYjVKFeWnATlRZkidjIRN
IUD0jd5dVezEnC7zt5sCIawJmoTsm1BtqtgNyAYoyplmO5ZRXrDkYrTWli+scdhy
Ib48wFfeUPe640TV5DQij1IdBYEN44SfEnEUImT9fr3/jkClCX0xngvDeQZlJQSE
GeXsBi8hBv3cbPuRIAt1D3+HvPljzk+8gqdxu40t0uKAP6Ol1TV8UHqv+2yB7SWG
xNbesQXAFK7l2UAkti3xPPsVZLEpTIVNy9GQZXENTq79oE3/iKhE+XOmmlzW0xfG
jIxsYRdRHsmV0uIYip1J61gakDoj1lTckFgzN+QP4+SsBQfJeQ/00vHZY2vYzopT
jg8/Z8G43JSnKtvb8GOo6BdgrZrPuobF0wtQChjwskWS5txIqmvPiw6BR22WYK/P
knyzxEFjmDSogwCeuf3reytNrLGfZmC78EcccRe0KMMwWdkSUIRxXRuTys2qQaXQ
yUYPtEbHyJkpjTePilW3gK6lIoMu5S4TL1DSJ+ZTOPtdSXIKGo6UNXgXIMN+51NH
A3lNAQrmHhrwvoWpQSn3dtmmc48P2b29XJG3w5eQyBGkNULjvDsLN807Jynnkfdu
akBoFtd2AZHzDYHo5Olvt4v3JUa+u8hJvRoszFmwjEyvHl90a2hKSmyKu8hCDEmf
GyOcDED4lF9kz5Jp6FzbP/gGU6ZAuv7i+gCN/x1uucywlfxsii0MfGzK+UMEsNgX
ejKLbJrLzPx7hf8Z2LsGOIofbef1ydZSEgtcLRYOXROxW7nUkJrthujhZYzT4Jr9
NYx/Y9LUxXe+6yXRciyAMyqwbdL5YOXEvPQ4DhulCvzzRKVA5Z8UPCSD3JsOcXjm
aXUSUfB0yUQnk9UY5rmvM9ZoZx23E/nKNmuBVV3lHZedlhUjD5IaPbGmZ2ebfqsQ
MzUAUteWUVZ5E7g0dR2e6k+ngWDHaYTWkg5kv7dxHbmGRoHZRFLrdfvVBLjvu8qj
53q1pmC3a59EY9uhGe41PX/M6qvSWUiyRbCKbozUHlVSF5iUOklMiyEJbV9uW+jn
viySwmpVM/MsaMTLPTTBighfxq8ViKUm6TiZZDGZn8+D7d+yHV9sDGFriSxDuUNF
Xn6Jitnyw5r87kqtKD4pxqHFo3gF1iKVb60iIjVoeC5vb/iZBH7aSttEqZMulRve
1KYijNZ8/ZKGAlCRKHXV0/aWZ3T6sGBq7BTpGIFeRWvmYZv/XewYXc4xKG3Q/YLr
yl3Xmi6LQwqfa+2XRi2e10ZVV8devmKUjnJSIF4NF7Trtj2NejKAujZfPo0IYmXs
0gkRRqwJIBkDzQwe672r50STNZHLn1+D0ORJCJJ+Sispd/6f5J84oWk26JF/T+F8
FuyyAAayCJVXe2UyWs0AuUAQV7BdybOicIZv0fyTfHaoiaTpFPjO2zvHla7FtQEk
x2nwLRB7/7xTU1HBnORPnPGyC6V1Wiz9jgYSZZS2aaDl64xwavtc/TqUIgdr8mVa
gosgaH43JRAnBeShZhqJy0WQOjiFb55AKDrJJsPV+rq7XOdAHC07OP6r+uu/nos4
HxpuTlRKTprHV6b2Id1MEKi5BK6kIWp8tQGUlIOeU84kumEFoZRSalMe5rL7EflA
ML6yV4wPBi3X8+sC3ukAcBlJcXtuoAH5DpwaENDOaK7DhEtsq2V396L8LA/PNsrV
ow8VUBxFgOTwPRzcGwAy7PgQyEzD9lTIkWp719AZHYm7gyE55MHtNTMoCdkYPPI3
j/Yh8By2vpLkQZkXU18g1sPTIFLD/TcURzlPyQP2QbOPJt07YW9ZwaaOx5eIlSNl
yMeHGSVQcEIGZmjShOzLGBaB2kkRn2Zeofm8fZmMb2C20ON0mSrJM1vMYnHZgS+0
2rF5qagDluJtDSOjEqwfc+WHiw51ikYHEOU3DSPO8+W9v/8UxHuqGsK60An1ZxRS
3LTLVfwOhd1TrXPJFg4302Gnjz6U8+08ss1ywUB0DOz+QYfzCzzciKRntKyIdK+1
4MVzmA3MniVNjNW9PzIB/6zhNbszpzxI8mzh0s7VYspYXzjSViYek9gTlxTIZ1Ll
LxCEFQcZxBiI2zfWcyop+XGL68DAph/NLfWQm9xp05Jx8ZT3WbYvX1UC25jZYwTS
CEHAt9k9UplSbNsO/GRD4v5Cyef8bzVWsJh7zRR8h7ae2rURSv9A8MCq20fUwF3I
rLGCn0u//aElN7KWxghfAbUz2jAkcbD3x0aaV7fEt7c8kCBQpUAuOf/kAxNWkEBl
bM58DUaUA6nnYGWiqsTeP4PHnySE3C1aufPOoJdNYPQhzqwcyezuuDYl9mju0u6b
T7+wnzTLjo/wM2ZkASZh2QySQrqdKkAY+KBLLhD4c5in7i0QiMXEOwWTGCUAVhO/
Q8j7LK0phL9lRuLIdnMaBhJh35wod9rMvvKy8aDQq9XhSWYrXv8U0tn54LTiKazP
8qwWOQhEypdNP8PDek0uUQogSzKrTaQOQsv6ImJtqkbt+gwQv7XlIh25m/fxAkdZ
rRt3/8WV14A+/v57Hd7mAP0ERmMhyulLu6sJuTithrIBDe/hBbJiAaI6UPu/Zc/L
2iUv8sdkJC3Cvvmf1Lb0vNXQU48GPPYw55XGfUpHanEIeqbw0dCeveQRz6GFUEPS
3Qge3x/qNcgEOAaGCQ5wWhJwmV0iW+0Z2gvflHKy/KMtulvjwiz9UgPANnXRYYFz
RVrzC5cvpVgh8OGSyBIhjACSEQIts90hPWvRMJRKuaV5TQYHT8p6vN8w7IM5ucu8
P9jL1tq+7GZXp51zA8FqGxM+uRksu1KSC85ViyVgZSxYAWzUzeyw2iIEDpQQO4ev
D72iYoo+1r++CtUWuKCgLRAeu1Tz7SkrvrGEQ23ylcwBX1aBMDhhJEMfH0yoe4t/
tH3SfHOQYoQLbLDJB06L9YUwtD4QvDgtTIOq8EqBLvt4fVWyqYRxq+SlYSA9/kb7
wUZeADfvygWzryVnjnl8WQD1GCWgy0XNswio+Vzvfdqma5WftS7iniFPrHmMfwNL
hMD321rYTj0IMI8SuAhfgOGt3s1cXDZowlJYX/OMTQe49tp5qd2/fNHCBIEwx3dJ
R9BSq3IraiUKUklAowSX3VncjnFxiGhO3CCNndK0SVPOXXM+GF/jK0PrcvTSCRsf
MsaiYLkkiRU0SvzWT5tHQVGVwr7Gp9+J3RSOse+IRHpYy91gcYkBonK4VHoUnrs/
5N3bNbfIB+LI0wKlqW6ZEAT9eUdUZvpfDcE47cbpXq9VdL/+chLoVtVu+1Jq04te
n+0g2fyn4QnvSh8ydV8t9wiG1cK3/4C5Zv0B0G43ucDSqw6Yty25bammDrdTNOLR
PeBnpc7EyqApvX7mhTSM/NV2MpdDNdheW/9zw3VMy9lkmLnc3BFplkzF2WRU2rJm
17LxeRLDh/WR5CD/pc/rX5wRrupw4DxAq/dRxPZex/KZo0Imkw9irTzLCuS2jPXd
5oZUXRM5Vc4Bc1XTAm1zEWU7ApsB4zKLcXNZ8mKzh1QMw7OTEhhHwwUfYOiFpaee
oehJ5fMdMtmzkUA64jWGn3aFWdOlQPeGg5zGyBMiXbQ+efoJzAsBlbkgYCpz3sR+
tTo2aLNj1J5jYGggqJUxVVi3qofNSfWxIBAwLmO6HOEca+ri5SxyNoyOCGunfv46
vZuWE9VP4gCjg014VMhGeivYyHrvWBW49BBHjkfkRVMfqvrcBkZ20q0C7SzxKI0D
4FJSAoEl1jvJgcGE2s169Gi6DUHKo2+BgrH7LyWU4+oMO6dAPanXUfa2cmr10Eg+
M2h53acRZDZnsTpsBogh7pdHAU7ikpDYojQ8+9vCr0fs9xGN15JYauwY6vX0Heed
byfRGeUScqRLJHOGKQ56/YXwdOQrB04N+ebD335n/HoEm+6TbEIDKzmU9q8tJiiq
yOqUEAzKORa/cJN34QedeDt6duSqGeLrOEXmQ+J4Vnmuqb6mUR/d+S4nKe+RPBYn
YicVu/3fmYCZ73/a9CqOsGqGFVp2uJcJ9kMJYS/efID54EzxIWOkaAdTF66ITJ2s
IwfjgOoGNO9dZscx4cAhbOdZ1GlbeSTX6DHCOCCXsN+cHvuxJDcGFdfZH2GAUkEq
8TGTK8W0h92rCOLPmeuBS864MIzlYBPQmkrDTczT5TcDIG3db6proPUesNsi/uCi
r6zMH1ceJJFjQe431H8LhIJflgti2I8uM7wQkJ+weIOpZJ+ES5UuF0C7PeF+ZVWw
rbGG8Odd18PesbFq2fCRc74y6q0/zqw5zxf9IGjWmu+lO6IS3vKdmwPNxTYNVMFF
jbKXOOIaGKWlKx8Vrzj9KXLE4vS1SpOR86ks8HcGFRTZiTcX9yjKttY5JNgZ4WOQ
1FqBtAona3wdDjy35tW7DGoiK7hbCUkpPtEa3jAGJZW/L1C9gN8Sd6XOjWM7USHU
W0ZwlbYhhQlI23CE0VHcOz2yP9+LBZ7TCBfG+zUPzX3gQE1FQcLB4m/UT0FonJpP
YtS1iqP+2RqVkgEW585HVzMwlbHrovv2rHkaNckI+bZU7rn3OQ1bRnKL07DxjU2C
YdbRiTJgrQspIcMroUxszG3Oqq1lX7C587etkQUhzObfxQyXdoPly7VqKmP8hweR
0Pq7KJiQG20oJ/exISVUI8m+9ec3Ik3CEivQN1NRYpup+1PXSqx6rs1Kf4eGD2Kk
H20TmPV7COq3rmWS6/uhgOMMfvgF2M00A6KoOLat1z6Gff6eXoAyq2NbN4iSKSqp
+qsb20yGeYNJNOOfn6B8IUTmpN2ckT8O/657fp0MrNhX0X6kD1Il6T+df8KaImnO
bk/55ZAr0/IvzZm963tOHek+SbsM8XbbHMM3zqCtYUgriwirBro3hs8PtmGAz93v
OGIna4pTxBp8ah849dL64cuRMkBkIflpvAgTrHoTssQ1V3mlQ5J/r8PFHtwzvaIr
tSigQB4fHAVmymQOqet0CT+eXq53RXkwuG8+wwPcqRQBEHA9hdrExa1wmVibYuya
eQ/ml/35jq3gZvY4rvTbDWmVl1SUekngUXZToLn/3dpo/8xybC1CzY2grJ5hXGxi
oZG2I0ZaHcFMoSaRZi8AZPiWrzPfHz6TZ6/T+1r0rdF8428mpdV0Yjz8LkH0OrXY
7QUPaoyl2VQWCtKAkS9V3ZcmMsOyb1ozz0SxpoKIQSc6j+i4XJALKeLIfHm9P9U9
kR7gcCqGPvho6VxLePBhXadS5FPjXdsISOfSW4QcD5rm44yooa9sRNGXXccNqYq0
OL6h6othm18oGrtbcJ13L++Pms1bw9zDCE38MJjgWWBMNcSFRQRgitAphpY06r42
t4LXjLCGeDLlRW6ZRsd0C2HRF/U1n8lVLyzmx6pCAPuBKyjOk62LLEE8rS31kToE
L2Z8mDF9n8LB+7rFCjzjX15uxWvEeL26uX9YyddB9SW5RvxTh9sMUR2FPlLTQYlN
252cX2oCyYoEkp4Drv9en3nUW/9tQlu+ldRagP17Mb+Vh/Lids7yCVueZIksJ8z5
V5nY0mRsa1sfrn0kou2rHtSQg2a6kRvnwlmLBgGr7ZZsMaGpbuGMct1DcRLkE/gY
VKJdmWrk6N0LoE6rBQUpmyZXTw65ejr5hhkobzDYMdwShiwXGZNoo1DXbBGHEtil
7eb+SCq/Tj6ZWk24VoGwUyYbVBKKmFwQx3Tg+Q2GTU3oOay8YYsl1tDiYaxORFb+
o/tYZ/9rccQAd2rDlM0i2vK4WNJZ/kQeELugLXVmvWDsp+NauUS/qKAdqfOUygt9
xEerqAbMYPetsCwSNsRMRdTvip3h50jxnfiVKU3bffXZsjzV/5t9U8zP/FskHgao
k9D4JPjqgNEmM09BCLOO+1vT+R0zBLQvsbYgyvOSWzp74yDAhxnj+WeA4Cka6nXe
/latp23aQD46Hv2MLFEIBa6KQEIrWGFoiMeYe410HGt06QLLswaTM7/lVRwz3KXl
Ib/P9sE6ecwuvIJQRuiv/tiRA5wFUCaOrchnAU0+MKmeaouNaEcDC8MTsGP8DLHP
PcfSeEhbL7zzK8Yf/PlaNCOWZ6uieHRIFn/js3NIBmIaPxmGQ2HWGcvw4/WOyEoN
3UcRokWtjEjMgVs42iRmxtFdmimKWTdNv+aPTCXFDqnbXmeQP2ptper8mnz1Jgf5
rZ2nxVXwqRJRjlSUeAqnLR0hQcklGC/CUpDm3p7XpVHghckSlw6Boioy3OijLX3d
gfg12O4ISmebgq5MUid9uA4QhYaZRHYZBTOXInrgM3Ou+FF62uSNkRU4BIOsddtM
2yeq3DsgzW9DXOtSNxCx6NxBkCCu8AHiKFw8Vbsh3oU6f+CJaJdWIE+8HuWPSc+N
T/iDwEnbHlmuDcic8rBwJi5TMAEOOWhaxemP6+HGy0SzUsBItDDwmc4ZwoRaRvqN
2x9zyVt8WJMqLj00cHP1HFg7k/erDN0t46alCto/f7fbATcqyStWaWgx+XzD+dOP
ERUSyZl8t4a2nhWUZHEAW/iGDqnm8QjFxrDIaS6uROMViGiAigZXxhJhYSEjfoak
ubArrbiooPh8L7W206kUEozWMPwOno8CjwBaCvwGgkCY9UaWR9PXdtwU1oEDb10O
+tdmtBT8lUtdXg4Fl7Fo5wNtWUuEw0X7vMBCMNmKW/LyjfQPFvwqGdvGy35Fl28Y
TFh0XxhvO2Urb30OrsgKZ8iQvir91jC3OnWA8S/tqTIwgqbLpIMnfyx+wuQeEUla
x2jlDBlRdES6RQKWJhFvyqPNN1TkcoBT+6f64YrnZh2d21pqT7TWwySgL/oHaP2P
x5x1vX1nvYoofjHovOusLYoZtM72J/xMQxSpSgCi9j6vDHixb2dfH6SYrv0cA21/
VxjKaWyHGl2BrA7TwT6CMQsQyAbM3li7Abxa6Ww7GTWDtTFn3NRZcdX3dqpFTUOq
wfU1k/QtaCqUOyZ9pX8KdxTzFGLtfm9f/JNdds2iYl9aajRbnsdJF6B6FTbhbSTY
q6c7JML/mpGbK+m/FP109BIh8QpGf0/3VaS/isfvK9+2wunjKMw4BJflAikkEOpF
fq4FLstPdojJjO8D5g8rBVrwB9rpQjChYu23Btfccf4JWnajICxOmNuJ2K3KV+Mw
WAE2ACxamcHTuXId4t9aD9v73bRkxa6RbE15xicd4m74rMhmKrXdLx09r51KiRNp
nY9Gf2woUfbLi9GeBiaT0vjN12Fhr4w+txbKUHWQOpF6PYyrZV374mDBTDqIwxP/
mAsUitgpFdeA4jN0yyDJYLhpIDSDJHZ0anMVHC6tzU9wo9HhZf6iF664szOPMFSx
bqwpFBp9pmyhTy0a1g5hsOgugJWooT2wGgnbY3WJ0I52xFKyO6xzACu4kv6y/W6g
ZYa2Lm3CPmGwcf9557qnrw3tcOv3ApLVs0aeAcEh3eM2CPZ/oQAzRXH+Dmk7uKUg
Znw9Tl26byqnfESa/hWtIPi21yWBp3B0zWGilRbL6o6DixSsFULNQJwilRoemFe6
hytTtS03cpc76ch88aBghIiDZitY2r2ck65R4yJBBUdbEmzr5ITY0j3E30JOean6
AG9llAnt+uWsKHq0gKq6Qgb9BBEbGqm67TvEyJBwr9fuQvjLN1EmgzEG1mOHAm9j
2SDxFC1t/e0bcnXsifp7Imnj+jgInDWn+rPUhVRbVadNELzvsQJpFTrni4mE1Fk4
uUDRJIpC8ScyPxEonRbsrBojojrjWvPcuFGpkEwmeRtv89judHoGeujdLBRuOCTh
or9JUKN1gnOswEkFZo/o44DsICROaSBxFkwBUgeVNucaWMWY6vD6if/ryx0OWtxK
pkf7P0Lyj78HeO4aPrcGl12APQAk9huR2MBhnOM7fTrhZuQrAYcsHdPQREonu+I/
D3TE01rFMTE4Zu1LD/aRGI0x6TnAqwHHGXrcP+UCrao/nvfRjWNcGG0He3oKNYg1
QUXbssj2Xsz0+iLIVShpEpE6Ie99IF6niYG+qZ88x77jWo+gdxtRKGAihjQTim1O
nZd1mXUN4wCD3s4hh7CTjgtgYUeIzBGxY+QTqUKNTbsSOBbwnfL23Xf+IExot9G2
OL0ZwUWtwjcIWfFBQBMy9RhWLKbYABRTKWAIghExtdYLWYH8dbbvYzW+vbWlRSLn
N5uG2uBNhv29WMePcHfDHk5PJfAeRilXpIH6mlEknV3Sm214gsRGCYkhiKk/kbWX
AEtTuHI++jddpdIpI4lA/nOu7nUyVJG5tez75HU9N2fsA4sHNVwiD+YhBePM6VsR
41Fl24Tr04B1/f51mkXJhj0CYJXQNmwMAXytejF6a+OWp3hoB8JFGbTvnPtfM8UU
SMEz6Uq8xxYk2ooAlqDr5HMFSHmOE7atjlL42TNrUvoD6FrS+aaXTpr2jqvjEKJp
6v+7vUxlWDEul3XilgJetYXHKCat3607jDbqpyGUV07+24Vvp5r571+XNc59Plr5
gMR5++VYLCAForvvEzJ7n1mnZOy8JxM5R17evpeH7GAZ90AtkTRWYBxZ59ufhObZ
15T25zSaPkWGNCdQnJQxTOjN+78OBFEInjBuckRSsUpO+QA+XqQX9/nOwMY/UJsc
GKdaJ5F82lqXdpmr/dzp1Nw2NWMSqS5IIdKUznlBERlUS960kI+Zlr1DWn6qptPd
8uKunAuJAXFMFn86Vz9jJkcw0BF7k8Jc7FoOZTU2Xhv9q72/jK0Tdl6pzx33z0Jx
dQBF0Lp6vKNjiX76Dau2Aemmmf6ylHw8Z5gZE9t+eSi9Kxa5jtPxHtBxFdGDgycZ
zrEGaAWpKXoxMxaILqfNt3JVTNr0zJQ933/rF4Nt30FNtaFRmVKh0GyQ9S0+ZZz0
F+GkttZ6aCETQOrFFVhGE7+ttUzYa0QRQC+NS7yAg5qUl+7NEsJ+TRtKHSKn7D1R
CEiao+y0QUq2+lMvVF67Td5pSlO8nTqO9omPJcRe3Kke8wJzy6cUQKEwewMStA05
DoCi+toT4rc3uG12XB0AocRr4ZkAbjUkRCskElOThsWOntxLD/0rvXoLWO93THDu
J8zrg1putESUjOTS15tLtKJ1kbUs78OlKTOlSzrQkiotCXwzgJmq5qtve3CuUrbq
RS0VPj8QFlNxEzddp/2XWIb8RH0uEw7SA54ggErC7TDO4FYTgZUZnUxLaQqszJ2w
3fmY6uQIOAnXwzmaptFtwiiaGgIqxScaHJErAefCAnzGoX1RBSXfnO0gBslLLu5j
CjJrqPXh9s8VbGWm5mbYIonV/kjJB4ySPODXoP9TjDQno/TQT6nRK5N6GBc7C+Uo
37eq2mN2hNCZYEOMFfXS37+imQdmZ9ui4bHWjbENANui6D6YdHVrnfcGLRxb9Lnj
7jcDXT6gtFGqjsIFQEpeMlpG1JdY3t57cw3vnB7571uWD6CTjDSPCUBEY3c4xlp2
rTrk6nTOG/QDKo099daJV2kO7IgLRFHD8XGgxc9hY7pSMZBzIpptncyJu46MIt0b
G654bDPe+NT5tBF9xL3zlcyWXBid6D9PNnDjHXFqeIGDMxABrstmDUQIede8BHWQ
uyvxJYYJnmyDF8adQP9KceM6fQ7xltCteOMNvaUbduXfKujVRBYxOEoyJnI8Pj3j
Y/L25Zv6pK7hJYbZeBtN1dHIB/j+42y1n8rKBC71y9RX6PIMuncw7Orr44PcW09p
yM1/R1B/4Z+Sc9Aj6QogcUwbTXm7lSHWDtQd6mG5fhp9ppHspaWi7ziVfClrGNOc
Ix7NPLMG7/40yrEsd4hp8fLD+Pj97oF9ujKokqkWCSzfEU6neLS/jHJBgfYxXh3U
lMSNXrEq3SsSeirgtg+GcE3Ht2MQG+51/4QVVb7XA+mmEwxlfFNqufAhh7xcTLSn
kBj+8dgsFycaVaCkq/ZD8gBdANGxqv8QSopTSPJ28+efVuDq21D+gIQlcWf1XcXD
lhEYOldHhHfpAFe27UyZnJ23qihuD5VWohQW0Qfy99imQ0HrAiyiXl7pER6yhNqD
9CyeNCz67du01Qw9QJA99MRGrozDC6nZ7nLmwL53csj5Z2MFK4h2Q9KykW3gIWsv
akaWQTzTY1lb/TUP8tVfuVNu2Ml9Md9bNc4eSzrjh+2pghfhc9UnkO0nBOGmpDmB
HxivQ2n5TJTXXQ5W87VUQ+hCtHIxHkyg75gOsUcglyuga7yr8xZb88JYWEHrOo0W
sXQcMSfiww9bDtXMVg0KycmyYgeDCGiUVayYplh0tcMThqqaqRESJys8FYDxOrPf
TiYRvOtpGMfK+AoDck8WeXcM+WjHQG7+z/ZZ5fXqtOJTMb+YEMPUlwOTsi9O8NSi
0IZJDpwRpp5XMfJkkoQAgU40MMLrVWYXnjDxd+7fF0FdP68WG8OlCsOP027ckRMC
DC12IGaSguG8/5QvD6AOkwp9iO8fNQ1gDEE1S0g6BvN/5xMwbzCwLtb2wNydGyaD
Qj+uw5rvi7DtYQvI6Rm4YQPEXhbr5ADp4vZeoRVbYBeQ4BxcEZ8wmhOZGB7DCSOm
CBDhZekIdGpFHCc4HDF+8TDH10hFhJXwix5qWXP2njPFPrMehelTfLcJ5PD1FUpj
kTpsqrZoOvUkEzdU3u1sH9rQswIfzGOITnAGD828q6pOBP7BXrhkQf0inUv2+5g6
oytTQHHBNeVd0RiCrM70QcHQRxzbRNE14WPwDSchHHlxWsQ2nYWivLBGaOnb1bvw
RjlRW0RVrA4le+u2h8gCcVdwdkT8qThEfCp3yBjo+OaptDqGrO59aR9i7aq/qV0v
x07ECGQicSXH7Y4DZJaCQTZfeld7zSBAcWfLVXlfQU3W+Uhb2e+jdmMgn+ii64wf
XxtC9V1RWkPOFrFjV82cBkw5i47VgBj/UXIUaC0T9loK5iLRCIpRb5fBhDwmqrZc
yOr9JqoUEuGCLFS+FlF1bcdQq+z/CzTVdZKxb4hvI+0MZOhDnJpYusPJpWjvCpfn
jANLn36iNFJGgIyMZkS61nrGWKQlo9tbgHd19P13C+7oKCntGgy+AdhCLFU0Fl1v
JLNqGfZ9A0Umclo+1O6rj+yWlXRdb0gbqtvHe7l4OCGYjDqqr79thgowR1vJNATa
KioXWT7OWWr4y2O4B2WQ0w5TqIugpVSdjRMiteHaQXxL4ty3R9xWFxa1g149Z+Uh
8ltxkN84AfdyAvVQjfx3noI3Ok/G3BGkbly5Q1Bnp3L2PGvjGffv/SyWCCR3C5Nq
VY4ojujOppeSUwCdkPS6mttxutNkfFrRQdAGGOCYlHuHetS3rLquMBC+/aoaVcLV
6WCFGxlgF244E+TMqCu6XFzHXWCP2YWjp+O+FhHZ4QtfMgFu3NJHOTQ3XKR9TcHg
skYZi62YoTMBw62dUPLFUDbCHSb4vmts4Nr9DnXxvLmDuaW/TdVzd6ZcdgVeI+/X
LWf393/AgxRYNYvtWyQlp6mrOPLY7NiBEYksP8tdivfiY07lhMhvFtNn/eHjt2pA
Z4O2Xxb16y+f49zmFtXxpc2WFKPFctROMUimf2ozrfWuvcjeFAsE2Fa/v9cGQLNj
mVPi6uRPgDccH5VaMpJreuGeWAMK3kVn9HJUVnH/oPtKC3YOXrAbKxYCAgU+PPwe
XVvKMOkuHzk+Qx1VSEgQ0sjbmEStnOtQ3/lIrmhtrnPWPZZlqXmsYH/alm8mqFAX
st61rKN+g4A6FzOhfnS7bTJ9MCQF3nADlxuBgbNI9+/StLmcHcvzbqCMVIzeqO20
Ab2t5J0k2hLyxKkjQwOpt/i13JkDQuBuDpnB0TbcwAApeG+2kRyfcmAg0MOHj54x
wowhBFzDG9VxXiczx/sta7rWIfWJ8eXrhMK7l2CsMGk3iCpifpDGY1fM6YktOTnM
cHTokCqjKy4VYZA2uRyVSFBy5AxULhWtfa4ODayooqN+UW52eknNqp8yqkHajNVm
kTw3s7vvCmLxBK+s9FYWDtWRpbQEjda194sQHCxL0J8TMFhOwbSZVwtedPzh2dBK
fzDEsFr7ag2eZlTXdpFqjQsoBf2LUmx5OB5dqbEKh1bSzkpr7zaIELIM12RtnLkl
THlosiUETfLzeurpJJlAHlM9daKFCBT2BUvEJKl3s90jeRZ40LlUZoJNjPdyOdsR
y2+uLRJwEk0tG+a4P3s0mQDecnplRWnS77MeaTf1EqoSaCo9UxE0kx5kOr254zv/
5qVUcT0OZyRy6M61IdGIAyeLS053UYPDfzci7Im436RzM4zBAaJd39v8lPwcvUMx
yALn6xpDbk8xmOXyeItOfC+0IZg0Q9o1xISSzIXhzrP5aGAPK8rTh4eEEsnE3gm0
iwyA/Fnk5xti1/cOEzDFYk7dHDkU4ulaKFHkbevUW+cjS2i3BOvar4Y4r4SRnSjR
MpHkJrDBAHeGQstCRAUCNajN9t6VyDajo+E05yYeWdVyrKFUB5rOVHNbaId31Rk8
RylIYbmGjq1+124weFvNc/7cm+qDfm2y1YVE2mA+s3ye9jmJ1fqsethPlfQd1MgJ
75HHUy62qspxHvvRr1JCLT8LR16sARlaIG3Qy+OR9qN/AVYK/tTdQDjoW4a3RF/O
xFxScfdLlbnHFy6QiYD2wmmKD4j0mP+AN9ddOeH4vljTfBbNRoAB7gwhdjbYSEUG
hDCSU/cNNgSPvaAqrW74b2/2qOc5jkWAekvS+hvzk7pHGOT/5xFoZ5Ghys35wdhb
pr6J1h482M5dC0MsIch8AGOstyO0+kRVB5hi6arsZU0xvsaSM/WLmSf6+Ka13y6X
QofAIwPwDvBJdQkMWFchcbsEeJRGaaCH5ztH0Bq7CRizfUY/E4piXbNLYOWxPXM2
gZb14sAJiuLflfWmS5KZGMeDFDwy9qR9EmDhfGIkGFAHzBY/1pRL+QRafuv0UGnz
h1hVLtCNfyDzcyhtv93mb2OgE2Sd1HaxgUuuNABpbae9xdA8XDH8IWDpTLGGZwJk
xMM4Bai6u+J9YDshEMh6b0ZdkoVgQOAgX/O+hFwjNwEjhMgCSI6nhDQVnriLmunD
oecchCq2YYbfZ4Z2u/31ONKlCQXuhURND+x000Kj93hJmpzCdXgIXtqK2rDqiH/R
p73v28LuzWXRavb3hgwpLg/EP8JuzqJucxRo6rEyzqtQMuxJFmrUUsTKA33sZwOJ
zblEhOGm+AYNYcgDeFwaos3HFsnmA2Uxj7ACkWoHYy7E1HKyY5Brdrpp652WDSEE
Np9TQHVCW8xx/2X1XTvfBbhgn9MWbH5knJcLZC+ghxLAlELP6B1MVq71OQtlsbxQ
5zAwrwu8aYX+opBs6aUHP24Zo0X4+oq3s8BSdHhvIUiLvgaUZjac3ajieZjq3pkN
9pKidj9/9HJVL7mBjiXVNyUZgIl0/m7lv9q5/XVcrVObELBPsLhhJZd7AIIYSFhD
6pdaiovA1GeObu48W295ccmgTDXmw0I0g00mjuvv4UlZJLVGv0BDai96MGoBjlhT
OL1CZRCMBpbI2/x67IWxEeq4V9UXMI+1ytQs1gCaipcMbgYEojGxP5Q+0uTwHioh
LhwWixLu5xmPY/Biay9VLrPebWzDVCisO2GCxuF8nPle1ds8Bea3r4/i+PSz7v0i
ciAMGXWqchNjEfI0oAkYSRTPpHd190xrjwtyEoLZfxx8ApOeDIW9jqybnwlnB2zW
Q4egPejywIc8E+L/zxyjfDPpKftZz4L4d15N7RekFshC3RETQv8+vdgn4DA+aNaW
QWVTJhLfZPqkPu4q5YMYPGBE1Il6IHAM2BqL3M0Wbp3GnrYQ6h78mfnagh2Dz3yl
rTIgspD2FCjg2WX8o1jG2y1ox0l9/ErXxjbl81IszD/lvH7vvjPFy490SW4pwZsb
KKfruy+H7BY8cUjwSXDOvs9X+2di7rDeQPaZj8Y9bTAjWUfKkf2qmCh8JU+GDSnQ
CHxDvaN9o8+x3c65kYvYeEzbv8b+IW/71OypWitIATuTSmXo9srgSgtkBQyePThz
oL9eStDTfCgonZfUV+e1hEo4i6TQG8v+bJII9EsRYFNpu6U8/4p86Vm7KDYOJZoh
Z6L/sQ3F2U6LrJJGtiA84Rn8csytN7duHYPG0WmzKrf23mZL0fcE9xZpSBYvKjRZ
uTcYdjU2PBxhGPlOkU8CtY0JZIhu4uGRjYxjbkbCogrzgy0AqA6MnWvYLdJqNpuk
Q7GrFibY7dQPjW3CVRfw0vijZif3XzGWbwFjeTaA+lPPqzIeck3eRuxoF5DlQ96n
aksusarLyYnlKIqf1xDe6GUuvm/ExtA6eBsXycs6rhbObKM0laFC0+wUfH1M6CfV
iEw166q7CSJwjdcxI9kRpLKpAJvCiNytRSrXHBYqnVSIdxI3VIa8f9gThj65awCP
x3yIs6IJ7yvDNfHk/rditnNctWjnxMUL1LrLjtWmUXGd7xZobkE30KXR830LMBOn
oyohsVbZl2hc+ChyCJNxKcwvpwIutnszatVXwthQXOIAodZTQ9DZR/Y0TxbioIqT
TeZR/QK8jWu0Ba71W4uduzylGUb8+88+2f0SMjDpytIzAU3E8vxKNjnRFXE6T/Lh
JuP90C8knwTlKDRnsOYY05/A6F5WbsfhZzq4pBRFlLOPyRhfDj7qMlIwZaJFRL4p
rg+Hh3aqlfn/82CDBXPSXZXMFZd8pZ+vxkP1R3oJDYC+Gasz5pGTtdyokkPGwDYe
JkkOufCCwJfVq+UCk2UN6V5rg7H4/ka6EVz8vdd/ZgOjNeh3uDIA2FSUescmdo6W
K3E+bLEsBCgKQwx7kNqu0lQIOscLbGeUKRwvtEMJ206rQtr/p0CP+ZRSCQu43f3j
i4YgCV9cXcLjD6SPU9LBW+RhCfRdROun71lM08j8Nuo04ULcDRHL24eg3IYxOU1N
LPI2d0ZmB4o3VzqPrZH3UVyivCvRvF9clxjjRH9vjldTRx46rhQ5GERo3VjWDL2h
qGlpe7Qa2NVnUWPCGfudIfvmpfzx4HM7n6kWnBlvHYDTF47X3T5qJVAO5Z/qnLFC
8Xav/jVu3qdQgSI+XsOLN3ps0dVZFfkkbHPW9Dtxqm8Yb2XEYnGZFVb0MYmz3l9L
YcP7YUjlFowm7Zjokh/fWaKaD2nwNAXAWZ6JkvfjvoWsmemQUONCdEaKq7NhvcHr
skK0L2y0khkjRje3/Kmf0PdG0Uj5wSwFoKMn5GwVML+fRTYGGEgPgyA9co+VKHeH
mvssjedHokAggd4DTl2i2Zj7S3smR/83wxDAna98U7oe+7b+Y1N/ziTBKZbfNCvW
gjiwQAZEr6v4bHfZT1306x95/NH1P2Y0YPdgB3nvLMARIu4MrO5NUQ5AAQ094NoF
dTKVxPSgVrDANEi9II2nS2UWsgYu2xrPhPoyCVlGk87ftpFmfteDFlgXb4cCdLvJ
6xFJZnuKYBdCf1r5iH8x7cXJd8yWIcEDTEaOGiEaa15bImbvF0ouVYLg27X2QJMi
fm0Dn8bGOYFwurss12d5KIe1VXUqTLMCLr0VIdk8DUafxlKFPgJFMNvMDLZM0U64
VZWo2Kf4jSSvmRrVukO522mczOzgyCg4Fwv6LzpQZHJ5M/2DAvihtrIyKOiL4Ot2
w/qn3Z5ALXQhO0+wEI95AXUnVk8fNiO/C3aojnCG0EiHWN2v6pbh0fsQWKTay65j
KLTHrt3m+KEJzj0v/fOiaCdrobhxYigcjpEnAk9gEm2pkC668vN5PWQIfVqQwv13
Ghn77p79wk1zbsLE95Nap1uFB2agnXV5VTjQ1pDT9pbOhnAFm+HQsOC2I8JZOwle
pyWWpCIOWXv14T916o+vtOrJFI1x2RedkCh5CrymlR20x0SRxuV0VIn+JCVEumv5
WFpguccmVlKE1rfEXj9FBXK0E1eeOT3AOv3jWa7ha7+eF3VTrcFjjqB4blXxCSY7
4ytFQ3KhJ5wRSlgY2f4oBVl8RW62hK/Crl8jSl7hzg9uaqMX7dvsDWG4GErUJYeP
6zb5T6i/cmHOvYZ16TAbBfT2y6tWRdOq104mL636UwohUmasqaLsLAdAWH9WqEMC
HaCDkD8ifdUHr8SNxtVPwzl6jSh+TA0YfE3kDE9uo6FqYO11EFMmwQCI9QvBtvRw
eDsn1Wib7F5iPSK3A0Sxa1XZLXo491VSVaZ7NRir6v1SjuS/UB0TuPneSntNvpaL
3tJ9d3rVN3etWZOXmy2v4fQSXtuaUIXqALalLY332n4eLFQct7SUJqpVxbCswmeR
b2xj/+AfwAooT/7ohvLophbksjpAsJ5dTg4ayLqAgv+uJaf0kpCDm2cxd7AGID6v
+4Mnd3u9AH/gzNVr0Fr5o6WX1nzdCYOPkmiiLAVDVAiKYAMEDBKHRq4elrbFqfCh
HhYHjQFM6WDLv40KeGcJIvsXbnYNKRtZl8hDZnNpjVFAW9bDIbHnm76TcW2th6u+
c5wPJj//frkIVVzWI2wGTcm9qWF8PgRlNpgvqdv0a8QdROyU0aoxMfAmUFPiIg+M
gz8wb+lv95eyM7PTlTarmjIU0uASp3dR/wBTSgD/BTmJVM97J5JbKviA4Ua0GEc1
Au3i5AsqwncKdW/6QtGq7hcfj1LQIuPlawvW3G3NUitV3H6MK0xt4vpq3nGo8x6U
M/wA0odPHwSWKquehPvEH2l6mXwHtBg1g1L+tF7JX8PMEaI+jTgUOvCn81l24os7
6bu8D8EH5b2XFpD7wjQsRxkLujZ5/YbF3jw/mEAFpv86lImvbhVhhYQ5AVPspPoj
D3NR0exI71EKMiQ+4PmvTW2vtLZAWT0aCvv1YWQOatwpJ33hb5Vqh24YTqUDty8K
izmRAk54ctL6va4H7pzFjxNho6tzHvxofDpKXIK+h4BhmzxfPdT6f4nhErxtgfKY
P/bUo8Sd6s9ny8PSwjqLjI/1tZpM16KnbFin49G23HtcRdH4jG+2AckNv2GkAIbh
MgsUYn84LfVZGHCvKtVXtm3yxJs4OlkYFsTZUh5yuzqYMtUXhNu4fJoiwusAk7gy
f+Anuok4D2hiOLKjqXypU698tQ3YmUvo4TCHZCAK/CbIWgZqGeyrUQdQV33jhKs4
ZWnQh+yyqO3Rl/gdZxty9OURJGFZ/MPulhNu23oofZBJ6JrXTZjRpJZFJ8d+Xc0s
arbzN2cVcIeXTyyjr888LNdDppjsm9rZSlUp4uB9livulHn0pQxos5DC4rEwGU3k
fAMxRiD0i77w6Yr4H+De2G1eclf0ZC2+HR+NY6M7kFCIPkRoC+djzn0nIFR0HSZh
hY3BdsF9vR70TJV40AkfV9yEZ0UNpEp6znh+tcxYiij/tY+UbK+xjyNybzESVvJO
DJFOXylX1IayZ0rk4N3hBerFn7N3pu9Dv5pa4rMeUD7kDCdLomqCHGVHXa73jR+r
d9vbSJJf21fomU9OyKzq8Lnm3yPbJ0rarRV10+AdrmJF6j1GJuzsmJhwT5E8Y8IN
e7Tp9Q+sqNZaVl8XcnGBzFiztHssUSqqW+e+ZjRH5IGGbojiXHiyYsCtJMnoA+vF
GsQOdS0K/vJu1tG05VGULvra1jHoSuOs+32j79VaWQ9waGzVWfJGvPfy5BFKpOXQ
xxsF/hwNePq78swuz8JAXLvr6Vtfpr+P28ngjAWxzXp0IOm2DV0ATgID+b9FObUh
kjjgi4nKRhoM1pb/ij2A+6DUNdMo4la5Gjfr72/AMJ7VHqGmqfRlYA2ZfpqckFRA
f0IA/sf/RXNaCdhkOYWYt9k58GSZQG50reoApYi3bahkKSOoY+0Nqyr/7JesUIhJ
7l5v7PF0U9oMLwJRd/gWIhZ8weY+ID1h9xe0NfzxV672T4y71JM1+ll2wUECb5Su
HDaskE3Q3O5a1BDUrujbm3O5LJza0ckp17CU6x9obEAN43N3Piy7StLD4jzzgtZM
aj84ajOpYfH91JULdiKfjLYOAcb88x0jHslIR75ifCqWTdDPmYr6Yz5KCAKHaJ+h
X1ei8F2Iqm5l/rUmJnUGTzmzdzfD+xjmkf0kewdaC5znoK9okc2p7aH1aGjJc0zA
XdZETQ4DN3sVl7w3NjKcyRhE7j0aFZzgepHLkUrlxVl002NM2r/wtD5jcPct0eH9
f31PDsVqdHRkSL87BmzL2y2yuxdk70YbhRiLpt1zGVmCmuS2Fg/EGWohqO02Ujws
RstBX8J/GyrGiIONkZfdZ+EOzj42KX8llGxKyVuE8/1B+RPK4SPL11VO64AF8lKB
1N7aB15XHz3yC0/i/E2g43v2IFPHL95jLlNmA9zE49jZ3PN4dXtmHoguYnmFWMQt
tqD+YY1hAUcytvD8nVUYSvsUrGf5rnejyCEa2uMSmrRYT5N0ZTE3hQZVbqAlJ95Q
89yk9sISbQ81Z0u4E+vmN29yjDCUDW8urr/y2WoAjQZAen9qmc0/joxdR4kUaDPP
WYOVZe0xTjepHal8Hb9y6lz81guOdLXvjDmvbv+9QmhlAgwbiUrechOPWb0bAd41
x4dnlAVbngQJZNQRfIh6NuMeMfGed1Yufjll7oIG/D5EKfQ3Y8I8wfaLHiiSWkKt
SLtmCXZBBECXvscsq2PJwpi+sgGKtu+dVRRd4DIXyE4U4FAEwII2ScMvlUuv/Oba
LNcQjsdQwCxuVyd+wN18ZB+6P5up1V5FxSLdwZiD3sWMQAf6cWyyMTEj6KRJaV5K
X4U7rfQvRYhYpbmbLC/9K6oVOGia7ULLSrCXoVSaIy/dII4BlIrfx94Dlj/Sgasl
G1ISRY1222Sr8C+4nVAkbKkiAJJWF7nDVum9Ni6Uk+O2Hid1VXr4SdzAyKbK7Fvr
D4H+XY2Xai46ppIJxFGws+uehNno2KHnJThMZkUh1AeJ8xxkN0Hc+b50Jj0BVrFp
xVAt3dqVvy8dd/DVL6R80djmy9OCNZOXPC7tzRFNWkl+rkCyV+VbJMXmupqgZe0y
76A8PUoes7YAoS7psLTYYDBIstiH2ZOlCLDnhSo5mcSu21186ld7e87VG0MEPwnr
nmExPTzpYYgARvuRmo+GZ8YgLQwGFd/0aVBVWCsdHu1weebnUmqybXni//+8K7+7
7ccdr7uc9OCzGkj06xqIYbJ5cQoJAM7kmAsqPbCFwtXd9/AMePxj5yax993Tk6BT
mESVeYrJAU78ElBUjMcsGdvntO3KggAuc1JQowo/9up2UPbnSDYelMob7BOLArqA
qlqpX8hTOeaUxSOincSQWGzS4kcnYuT6RQ7Xy5BKgQTQ6ePsIp4gDYgeZOBsldeo
MM4ZhaxJcX7nCiFAtfuqDVl4ue7lyEw6Gnfw1+hQ1XhiQQtDy3i9YsscuWNnx60G
cLZcLFtluhkxW8/rnvJe4xhpJafrDMDlNIh9KzLjGVPeHZxspKs1P9dy1IAjuw/J
qCtq+lIjvd7I8nqh2iosjZrRqRdfuF2upJ9IIjKmo3ZVc4ImAgTsQx1Lg+SMJ70l
/YPhqiK2ggZ3dSzBEm3T6QAUxiiOiacPQca7oONxUlNLimOpEw4HoZaEmx05g7yq
V4Yy4cx7lkXLREeJCKFStUnwHCnLZzroy0oJ597Zjo6qRiFjndkFFD250rLazgTB
a35GGbQ4E58+8RteUEHw9XExtNSvT9iVxFCD9u+4c9KYOpwiq4q6yNjMI95o1S5I
AL6b2cNG1p9pmvfBDciPU9GHydtM1Tz9cPs/VEwJh+I8KDyB7cHTaTKJYb/L7Ryu
XeQ219zPNRMBujKQ//0kPj0AVQbu2m0XfzrhFONUSBiL1L5FtTkSJTLN00JYiBLQ
dVHijDVoYi7kf9Kfs1aMGDW+r2144r5dxS/FYxYn3Nam6YZXhMfWKVvNv6mbIpWb
Sg+fGXgl4GrhSm2WfrSEqWulm4iSbyVLABZewQuYCgwITV+fTOE2u1V6wh2MRTq3
JEj6hk4of3q83M6+6rg+/mpTIhn31akSPiJ2Sym7FOFul78Hiw7RzRpzZnYfZC3J
sPdGmM0C1frTpgzjd0BjcDUlxwLOIN0PQKuZZXraJF8LZqZLm6KFV8IQbi+6fWiJ
8dbLUNSYTwMFLFPLfNkLp5chgUeBMQ4RstEdtnFbWswxL0JtCoBegeTmZf4cCuI3
eAnK9mhao8w7lwDut8iae5jReaZCVHQcV25OZMVrOknFD//RxIS/XI+NcYmAXdc0
gMACGI5fvolwwL27Eh4zzuLR4+7aLfDWvOJkFAbXF6CtjpezHfSxwiGQnoTsixw+
QcldO8Y/s43AowgWUnddjxNVxhgAqJDJxcnrbf74tbzw8okBZEvgXDzZ+J+6ONtf
ftXpo5Ms2bdy9zkM9L1l0/vSFVh9H6vHVs+HpvnaveqDkMPUd6cGAYk2VKrvvzKG
w1fJUCnFnj+0F5ZjVW+EgrHiisedK7CTp+ZpclRvO/7s2b9Ni2VSAYooSXOn+Rsd
sE18O/0EgGlR08zfsnGrPGEI4EfmwSNCX+JhkkBqEEFf+ahqgL8mWF8/cHp+c9MO
eBzL9j30ZX90LXueWowmSLEPMOCqRJtwNWgx3S/epQz2U351uBAyRpuKLQTn92lI
2I0WWSpZM55TibKqxwI1Lr3+JLVY+G+x4ibw3/pmfxdkYEtDmzCMSkvfB6Itt1MY
QyM1tZjHUtTw+2FvUjSrRJ8pkOCrAwZVohtKhMJtgrBJ2gHcOuZyAc+CpUmFihc/
f9psh6hMpq7e9bpECmTzJwOXuDt6leuPs4hHRkDZ5Dgl0p2KQcAx6EKEqaMLEo4X
K9lqqTQhObPpHya+66DFU44gBFRax91o/AvKm73XGTfj2fhM7pGodDui8R37LqtC
WHEIkZMteEJNqhz1V0sOC73uJh7EMTInuWUuRRsDR0FMWuBPP9kMiP9w2o1wZcbD
imEzpZa9JCSf3sEGcSx/D0X9hMvmMBk178xFB7ZoIWVSVdM5WA7BxUAxaTWp0ELq
Qg1NspbIu+7xhjBucBJScBEC2oIA5nNZBOncFNEVz2+fLThdrW0ap/r/HVpHgReC
jB67Zo4BDEVis/uWy2Ts2CEJVNSWmW8DJgxPA7fcjgJB3jKX6LtzXiyiwO9+97Mq
+KJlpHKj9Jre9FqJ2M0lJGwd8q+5trK04rrJgb3QqSPqIpQUB2ROV0AjOXUk3xiu
DKAOIDOC4oYtCuVKIb/z+evJJWt4+S1dv7B6W+q0RPRma+/ALThCADKFTMHr2kyn
1eH4Q7pQ4lqfBiUiD+Jd8MFcxmoLKPW8wN2ZA7z+cVauBFBS1rZILxc2qexxtoCu
pZerem/F43/NuRjAH+ezGHYYvdJ9emPw+56cwkCdFN5WVsvldkhjtcFy0K5mC7jl
ovIkPXQHz7WcEZ0iuDv1gmzPJEtNOPEqiOu6G9IzPW2j495K+tL+UJ2f3gBF9qRo
7FvgwcgZhDYxH8c5KsmXDgpWflguG3eTBe9to9ncA1QRDXcn0Yi4w8YB9mYjJUYb
z4LiQSrSlJ0qTGnSEtNWI71yKxFpe8bEnjt0f2sjT5fMmQTCgdagEHyWRE9kSlr/
TjNWlN4SNQEJMzCEf2nhUVNHLgRS6T1AoG1H7hCk/xy/m69o57UrDrC0BLMAavM5
lgIclcCdW/vTqkB30v5lbn0SgBw90lck/uWjsmaD4pu1jVihSXU2yj51I+p54Yuj
ULUdDu9PmY6wDjWwWkOIsj5tC/RBHelzPmD5hOaE07+pCT3xemNYL+XEZuIDIVZh
xMZ0E5/HAtYojg1GZgQMNjMD4nPfGD+ytdOh3TBl++NpOXIsZloNWBksBgpWpN28
eiJDqlH87wxWdhkuUMeObyy83eVSHbz4vw6ERGq0mSJ6M7wsrrgqYvW4NXb/QSiF
3NiEZ4Kic8h9NNfGsQSGkxurDTDFodzEq3th9ZNMpGmOWuClRB8+D5EnSoVoU1Yn
AdGYRrFWWzF62FrdqgvGH2RlXmpr2N+DGDgp2ul1xOVHNd1KlmawGmfkHRx28bGt
WrxKlW84X3jWmNE9z0sElFTSpP5JqzMQ8DzKl0VoiVFSESIphK8ug2AU4vRBuqp7
Shu3glQQxbJv+sdtxzsGy8zSJOg2pyFdcuBSMqYUxHCAaFCOFDG5rOx5xybv+fMj
GNdKl89s+/9q3YfKlOx7G2aP575mSNCdWHdFxEumnbc8shcEA/Rwiqak0/v3tmXm
mGlAmwQh6aPbrS3e3LqPofna4DtNYEh4qxY6uQf/HItOG8OHnRs2jERzbvmlwnNS
ETG6QSqcdrsPvOlCWjBaCQUGvQcmUkF9ZkFLS6uoLjtDvkDta+vtpBjX0bq0LUKb
oqJ9avl3Nvi7OeLmQqkaHhnI3ieEYUO1PsCorP3mXFELsqtWv2AB93poBlF8q8iI
XZkYYE8NdyPW8B+7+myj08L72YPh1rP4oQmazDuH8OOW3yczQS1ic/8ROftsG9xY
oJIFnv1qW5IrDyumY+bIzh24NvhKESsigLXR6sq8t5yalb/OQxp7D/WN3C87/aC6
lneIznjGldnzruP2dGVDL5l/r/BKnnxz+lrIo3G5yQ10brUao1+6Ps1u/5b8TwAi
QlgSUL+Vlaj6S6+U3PxEWB9qd/fV67nuN1E+UIebqxQymNTgSKERKFmpW7av4a44
pxD9imKYwRLqAl4R0bBowrl4XOXyYJEETecVYmX78vnzjZOetdeJjSSnrN2MW0/W
fgRlfWpxbBHl+P43IDMy5H7gxGgrAHop+2m+AeA/TtVHEL3wbnBvczf2qbuNshES
oP7gkMnRI6koI+DoXqX7mfjISKpl0GzFd8G3faUUGbKDUzeJ43vomToXM05kUP36
Ca6AzAREo+hMICjwEyuOgjLG7BgRTraqNXSgwavhKlLIM5oSMznZjjn84TB9D1TA
IBARsy+6AISszKRejNFUZyqbjFrm//svC03qm7lcW8g6rYhvq3MDT4BbN1rXho5v
YkGb6J/ACFVR1C7+a11w0ldx28Toe1w9L5N1RRmyEdeFbJrrgy3A1PDQ9YUTdimE
5BVpJVCd8yijexpvKop50QYpUH7NPxSufTBUylSo+uUJirOjUZcVEqbBZQ2Zzjoq
2Nn8jlpbPJ7ekxenBqV4gT9B6zn9GM6U0hqs4X1jvcRwn56DlXWHdCOmy91SZYgj
RGJM0rDMZ+aGBenC2nzw215/+ws/bzG0pccWMDlvTixpqNfR0IzWgQ8ajm6UXwGf
+Isk4soUuYK5zfnyivNrgrfllzesNr5C2xcQgqtXs+59y7Ghu2AF3/HAmr9eVS6f
W5BOiV7nuAYhHLAEocjyN4meU4U2dh3lY9m/rj+9qysJ8bh6fBeXYROER2t0LRHj
G4S7fNjmB8TBuGucmkaCZlEiYZ7ZO/i/8Tk0lQyTGV70KrjxTavP1MJQxjIAfc88
ARg1FZXwKX3+DzdW05yMXyVqpr+Wf59Zuwb4qDuHhBxypxFdvY4Fjcc2G+fl1+w+
gQaolBoctDxA/u8xsKBdcoR3GSQHCQmtfmlzdWTGrQJFC1SoR7I77MbJsCO4Sbsf
SJjf8ya9/aFdHNBOOpEIoj2tRbTOlI6UgG/PkKa8yC2Bo9rl2Rhg/QuU4c9zsWWv
0KAaJ3xXEPVk9t+f2LmJfQUukrAD0UBe7QODqELWb+U0GE85vUQmDfG/piVLLt+R
zi297f1jXi9rzaiTbFuq9DLs7ugsoelbM01DISmWSUHtf+RcEQo4wMiok3ElizVQ
+QTdkH8KN0qAZlkwnvBCTO5CU3DQykkSUKf5+oBj7gIyGb9qyImbES9tepq2MIIV
wtrv8IqPCcc5vW+yIcRftLRijqg2+zDurAvSbETF8rt3eO07OYiRj1XXo72crTX7
juj3GwpzZSjwUe22jd0a+TiCzZypjA4NUipYe8c5OVpUL1N8tjdhdRbJ2gEhMp+h
dE6T+AANlwjvzE/UTrE+un7rbeP4g6BHXVSBKLU2tzxlTKTHTlCVClOua/fSHW2w
8mGJGgMxgZUCsGtKRTikWsuC+32d+tNmxN5C8tCq2hLfY5Kgv4pi+L8Y7Dvwi6Fl
V6EvNKlZvVu0CKHqDgrazXjrfuvujOHS9VPwFddkBgSPbuBOxMgTSOQWlWL0Y8cz
asbX09wU9OEMAI6YilGWiNWAEbG4eSTtpIzr615id57O13S4w7+y11sE/MQJ4q9S
63DYPkWdLZkyVoAeiAEGQmsKvI6N6+29/i6jDSS7bFVKRewQDPNWPGEeYLuiNgaQ
LPYYHAU7zmWtSbRzz2KzTJFBEcXFaNTnifBbcDGQwy0WTi1zgl7/SYvF6alAeQ8s
b/AbYQgNXF8ixuAgGw8Xidtd03qvBshAOdUVe8Ulvmdp6XY4OLd5lkED8rJ9kq2y
ByZKURh6QSKKca4vgg7kn0WZpp/PV27H95xH5CFG4x3rGVmzCwCt2gQ6eHscxQ9T
LaWDMWRrnypvE5YPiaYPSNzkXxTPn7TnBMOn76knoi+ri/Dl3q7itiOmHvszrFDo
LjaLFlMAs02HCXSD9xTBEnEqNZlfUKmCTHR347GVD/BTZjn2v85F4OSMz0ygcPZx
cHPCB2oKK3f0jd8pNFdPphQxdtzlRQBquMilkOlpQqqvQHl7KANWJIYlP577dPf7
1UOvofDXpNydbulRAa2GVsuS4W25loOIehSoeIQrLF4n7OaDzCj1SXcq/JwnA6nt
yUeiIcr1iLTFiIBp5WOnX+hsUq0a8tXpjYMJY6JJy/27ogtWgfmbemkYvXcyowMe
LxoV9OUBWWGMeY9MG8qlt05GZRTVN2nh6RZYj7cjTKSrpKJxujD3+oykfxTFt4K7
hXqJHIDtErLIs2L1jkgmtBbSrbxR8jYkw4gZzo5PVoMMVMSdwiCg7+baF/lN+5ey
1fuiE89S1Yo42H0bpjZ5WOra3JuMe0JddWNq753U5+dTEOYFN3YmbIQd3N/lhCzY
YUNqjdW177A6EPM4Q1lqrUDPsfm9PjjLEf9vM72jy2I7zc4LbOyRSLp6uhmwEPON
gIi1doSslBFRwtgs9lzRqCzwqzR0k3rycDUZFg9cWHSZF4lFb8bog/9KOLld4SU3
jqwpChJ19uJIquDXmBlnk4la2E/LtFYGJHydfSDBcLIyZXR5SRO6a3wG7LuSL8UQ
UfRG6Wf/Ts0++YESno3yWKrGrsAb65MyFzOwFhyqaQ1fPL0rEOrKJlM4gPGAPADx
JiEg6Idg4wtn009zDmpbVig4AmteDznNr/9TpxBPNIxRrw/KAqmNrdJEnPi0hlwQ
fKsamhtfEh9Mn3SIeazjeaRX282Lz0w2Igy4aHTz8DaLUpsTV9n1/cY3Ddij8OuN
ILRVhGHP+Di3tOjIqxy8WtDxGTU1VLlKYtHuDyzfES9DdFKexqLstzjKroL4j4z4
Z+PLghh4AOLFLsjPGxxTYRGrzCwEZrchAn4puT5ZPcw61FXehbBOCZGKdmVmVgJY
NpFC92CR2I3c1psxUCgoPQoLr13ppEHYTdnWOKsVg8XocIcNeizgh0gaYhGqi2ri
BuORyoRdThYVuRHTv8fkZd0NfYfMRHTJufoYnPwSo5T26Z+LlYtBTZWHjqdVo83Q
SzyNOY8woDR541s1MZuWyPV62fxeHDdvkoqsFMHvpZiIWFEdjuccgI0N4t704UVG
KxBelYiILYV2YPA9edn0vhPwg/Qp8Qw8UZOaKPKFwHpdWGIP9DVwAzlrA+3Z+aKc
gbfboUYQsAPHi0ZyJn8Yq9C4asK4kPLYCR2NBRadTLDL+2jOymxPJf64i9Fevvk+
JWnWCR5rD3cQ5ZcVLxFlifJdogn6hf36L6IZoOyw0Oq+43VipMalFDS23n72XX7H
6gm7oxoKXNMABZf/saIoEUGh5B+KGibU+f3dlrwtjZdEdjRLsK5U1clwdNH6AoM3
mB/1SS289U+0768crUS7EY8bsc6wWwI+/klerJIlIW+enodFDcytMHW/byiBbgD0
Sk93cBWrFGpbazLJ6Ei8q3152nGFDE1Rk3KzOW06UGJqXxSMWxqBz+H5UeB1x/LO
LMP7Yc91WrDfpcEa68TZkNErPlyRFV4EHgCbgeQnFRySPjTKGypnUrEnrscspP7T
pMtxjDPAkKClfzeOjIvgyrs2X6tTMSpsPXyYFapLrCM97aBG+OWBKr5BMZBflUYF
lTTZ7l8N11U+6ymrhf3erJSiX3f0LG/kR/JgK407LDG2PdMbDsvIU+gI19GCNKBB
3py8i+DQMj0xfPw3dKizhGBIZ2zsDtALA1Q7AtrqWbmhVj3CJUeYs81v5QEQqxEe
O7DTohgV7gxltNGzQw+oNPC/G5MdIgndWP2TAe+JHUHD7daH0GjAsPX47lqmtcn3
bBJh4U+yzSlExpw4GboLpvL11vJZrVQ9QIYcnRqERwHeTmxqZMHLwTpKI2YEK0B6
EEDgk7LPPK8qIOxktc4SLe2+EJoC0odsGVp+h+y/eyO+SvPVothEj6a6KSFuxKYV
Cuzc6YkR9l87Z7s3IkwyDan737UakDfoNJr7sSwpOPaHBdt6DRKAuVazponZX5rd
tj/hb+q4nBBYie7xC2xOEmekqRwDkiDIoJWX/F1G/zg6Gzxim58s3MybtEpGzmO7
qkAigPlsLJW/m/Eu1Al31r9A+wtHf797xuJyd0v4Ij5tfLZbQu/mBOsJL1FZEVir
N0NIBhKsB880KjjS+ypEvXpxU0OKfGIHakPX6VWGr8Go1wk8U7AOcZVcWmDTO/eY
USE0OPLkVCUi9GlDV5O/GCFsNCbmAV5HSkfNb1QrN/ZKibG0poFGoCz/T6ZjKIFK
P+wJY3aEyOD1N5Kv2OK5LZ1jebufJR+pymV0LKvGiXUPLi90Rn1j5gkkmpvquk7m
9RI5i/nnKMlKdAfFa7z+xmmgyUwEXoJxFjIQBREzEGLTxHJwA/o6R8C/qYvbteLj
2ucsmSsG3AVg8EumHzgKCc0+hGQrvM+669qDtd833ic4Dsg9fo3fkcUzsaQ9r7Xb
9RmQj7Ke9i9aWhF8/GQ6nxvqoIC3ky1So3H1zwX38fEqt+OaQ7EtQlbPx9Bejbnt
th2H7hZfBMMf3678iKHCshZGJbajOxsaQWTsCGxZplhL2Z+KF2/6oqt5taaf+B4I
mRnVAO+m+z8Eh6MX5KbCnNHOfU6CfwQeXO4FZ3riytRwu1bbw5F8xFXt7x+xpFo2
LF05UjOFVphmVDjrI7/KKvMb/KdUNDUctDWOsp1cdm1xvpOyYUFL/YBp7XSiR5L3
G4ev52CH1OQwLWV/vnWV4Q/6ih1YPUroNX2/uXlvnJ9bA1+JqEpkvrmoJL0WCF9k
5/ELYaFQviPYmhlB+9iVNnoWcVIz78SATdYxKwh9Igr8WLcQrG01fN+RyrcP0NWX
4t2udqbY5R6rP/OY2Nba7H6FS5snheqlfmMOQsNtABqunZY6JpoRQbj62lKpAUBt
T6sLZwL+BBRRatakaAwC5yycR++Zbfms2RC9GvXZbvPjV6IF2me7OKNKHyRFtD+E
AbV2bOvr05NL99RJPBFT/ytkvNNN0v+Q4NrhduLmuRquw1RQqzjLx0nlrs6MQDDA
fRYqHQTztCFrHnejqhcHQCBfEW1uJUjIqgvw7DNvMhpLqSpQl48zLGOxn4HAsUwC
VGX8jcFFxc3jlffzw1zYXVD5cKjpx3FKi41aL7gj8QogIdG7DVTC6FkPaQ11/sKU
DfofEcc1NZpfO5Lbrm7x46ktjnxlpo54CM046fWC6Du77b9fkxpRGRU5WOmNIUAz
xm3mjy8/QvMJS8nBUlg5O+B9MqG9+/TKZM4sSRZWxziZ79zCB9cMP5PFsO3nsdYu
rANqVxwDPVpFwBKiBcGrxW7j8W3XjUqsLRSOg5Ph8bUEhs1EuWQpNRNkaGBXJnoE
FO7vSV+mHiijSQBFRZd87xRZjuf7qA/pMRKWA5yKtIxvM9PAyXTp0syd6QDrDfhz
KIRETewUQkRMuy/EfJ9KEhrQynCqpKRJrpLSAAl0VivciZXEOudSDVs7zq1evbBG
BNLNWP+FuVLuhNKToUbfnOH/fruy12T5MEO8JIZ08s2idGd46nGwAkc3EX1s4RPO
SwYScWWghNMLLbkZg4C5FeSll4+FoYIo5GkwtJjgyDuYkZmSPNhXtH9nGXHzhKy5
aqfNLmw3kBweOJel7rU0YmfneBnI5Q3LAh7CqTQHwWQpjZZk66maABiYKD2qebyY
UprvQAsueTSOWNouhwt2lYCcgEfI9b5rhV5UtGI6bUoK++l7fx0kjVTg1MSoVglK
AhRvxwtRYkwE1ch0OQ7c0v86fzJh++yA+C7mxDqFDQeNzeBo4OQenffoJZrYSSFI
GR4GEg+fHq7Ky1QUIFeapkqEODRfvbsRdx7uGOvSCSwCnQ749dWg67QA9k+9bEry
E++REjaKreRxN9xx2YpJ3HWyyF8xwsOcStNQ2F1vXr3bUSkxHuGhnmd+rtHW4SW8
tV+MwOm+Im0EdnIrrxtSU3Jit28GCvahkKUq3tdwgl+vBWOIsFh4EL8q0WJweFSG
ptvRhJVb1qLcSgLpohKrbNZLYCoxU7R+c6k7YLlfPwwZVPnkg91em7dAJHuL+LG0
rfZsc34u+uvuQJ9U1gJbaPLOSBxDDQBC9OBROl+iBlEbbXB3PTKs2mAwsiKxLzfD
NNEkGMeMGJLjfhiCMXGNoMZbxPxo+3n0Pl9IC32X9H1xkmHNCRrVijirKJt8Tp+L
iXhpWFF3aDUHIcWJ7KL4IxbfYzQzOxCmmtJPCpD9K9aLOdX9WC2QNbBFHBnQadui
/GXefsm4/ap6hB91Pwl80CIsO/alypSrgEDI8QTOunhOAtBlmZallVQc5gfLAERw
J/pIxwWszm8qTsSslxP7ZhjuJrYqqey6kiONL9VUjEmYPfk54vfOSTVgfTDL9RyY
6LOENg6AUmUQO60LQiMXYT5d+mkhO2L2eGej1RDLCeiTmAHFTgDBwqL6EpKT8lN0
abriwMY8B/fYVE4/zq2wGjOtktnBdiARclW5hnO78P4tVtqwIFEzWuGJxxIID66h
jBcGVIw7ZzulKWdqWMO09E+QJm28bmTgu+45IICp3wf4J5U7mo8MHxvubJNPaons
Dyeaz8/F+SpB1AZIhjawSM01xaD4YK5RLH0DO2la3p7ZVO4r9TNiW0zEuCi6MWlR
PU9SPZqN4lOYeOM7GTKXezu8eQRjW6xHnQzkMB8cXXTOswl16gpLVMvwAGYIT2b4
OhBlR+JiGGD0tfeixE90iSg3TO2tkHuOn8RJEY+HnQI8Yf4vUpxWzAFaxJCPCjks
V5WML4YebDHlbmaYtEmGHXPt44cdzBz0OR3CXQa9FlpBex97tAtOHom0EiqHx084
szn1kFnKQzb/qrdtGs9Rp+9ta+ee7+pT/COpMkEnADuBEDoRftJeVaFYyo/5QO7N
F5djOKxwm7RoZhO1cXm4HS0BxoNU7z0N421MKCxPDLWewjhKI6Ernk+eavAw7L/G
xYnhJk5eCQlXJJ2xwor/nQ0uTkAJjYzLWFgbsvMJ0YYM0ZDQsoa5/KO9sEyjxaFg
Q4e5ecrkx8BK+IKX8KjWZdL5lK3zDLDmjd2Iy8dN+qfEwOz1zt/VrMie2rx/cGuc
a/yFnuLCVhAJGVJoi8U75qdnjhaN3//BKf+oCdcwFaGuTT5domqPTQLQxgF4uvBC
xHVa6vrkSrji+j1NQzNiQiEsusX+cDwcZwFzAKC01yg67CZu37n7dmCwtQHJ2hkh
OmLYVKPoWo8axZieJtdpY1xANKzZyYNjdxIAQ68qneB853OJEWTAlgoinNO2ZPEh
jSxOolz4/s1+bHQYhIAj3a7k3/O1cSK1DPA3Io4qE5Xa4h/4gbg6LvHDo496VhL4
iPDSbrD/lemc+Yj6XIv/1a9ef3xAZikARhFcjqmrVKCMyFZcE001lAFfD1IO44t5
Y30yr0EYsvpZhV2+cjkEM3MpPA3534cWhb8uoYFsnBQB6QmFzE3XBvIOfqMA8JOo
8QqVB3JgeEzU/O+p/c82OeAK4UJLTnpPuY0LB3e5u4uQ7kOdn/3X6XZONYNaT+ke
80NBA5Ll0NkkUVnlL+C7EMMrszZ88x+/I2UtPnOeqp2zRBz6NAYKmupezFKR6gp9
prdwfNVXDko8+KyGPwcZfaXX3qlHNHFnSVnpC8yGhwsSLHkTEiRtwOqLPmrJKzPt
NZ4/NeChyRFUyIRbu0v9R7QG5nPSBKrJpxlC4HLUV3SUdjQI8BytfqZBRnmhsyVF
1Ot5lq4jXwI+DSQEJxhAW+eY4ZBFBfI/aAPJ1aAhGGzlY/mvCkqqccK3R3Dji8I+
ybyyhLuwClEMhgHPNnGnFga+kOBkce6SbatblmYAmzPH3K9hCY1N0UlB2vKSVY/t
w0hIiLVnP9RfxglsLuUzH5C/DCQqxfnFCW7CHR3y7RMAs/A2QIPUDmPgrR9devX5
bcSkzGFwZZrM7vw6/9M2IRsg+davicEyiny6cq90YpFloZgBev5xPJyt5D1Opvlm
MvsRI7Yk0zjPpWJFiJ0VCrdFdfPtt5fjaG4PlG2TL2lcNNnmC3jKjbZShhIVZ8q4
Dl9bgzwxxgW/JIzhoxqparJ13c3TWM0R2TPARihPh4lqEiE7T22zuKrWcjADfr5v
mEgJC0d+CqjVDbup5I6ZcLyGTCOUkvf/RAFcIQpeqiGb1CTn8qx/Vl6n9s30C1zD
vY9ok0X/GuCfsAQiSu/93g1kkfsG6QvSn036Oif66bR8gzkRVqKdiQXhWEOVMtY+
s21GSUuzKK/09t+gEg65IW+E9y6gDhoXiY4ZF2jL37W1ykqZaSf1uSVjMt0pFuOy
Lm4Ikb4SFL4CWpC/b5OLj+YSPlKG0ro4HyEEk6hZ6kMnGwi6Gi/EemaMumJY1gVM
DoWWXpKhuB2jrZ7qj2PNXMnN4E49fyZ7sPKqe9uv6pWsv/Gni8ObWLZDNQG40+Eh
wAw7UP9kIQkwpuLpVaRG9eRRGQq2YuYlXSneK3TQD9mZTKYp2ki66bYm988DD7on
EUcPWYDRhMlfrlGpcm06Tn3BVFlAOOHttO8zkQgoZ3hABU9TQPLq3KhzFynxtupO
MQ6ATmvXZCOtmLjX1e61h6WKQiUOZWuLyzc5dUFGI23nRzSZgz5KJNT44KjYIyLn
u1b3cTWBh94bvlMLCqmXDa9VIF58Sx0bPB4xGILesvHBDsli7Jjn7isK3HSRDMP2
u/6fhX+XMj46havjt8hkHKhrbZyoXv9RaH2GIqrQE7wioP8JEcrQK7SPYFAeo3ts
zLFSJkAo8XKCS/Hp85bDfFAYmbX6vMaawDScDylziVRU1RmdWiAM8pXqSGBlHEdJ
Qo3ttjbWixoPlHaPrX1DbDYu3dPpnOrj3OLMKfRAMDxWzRIztP6wwIAUwP6p2HE2
xwbHZkga8Z9S+v4X6efPgU6gUelGraSmIzhb3T2W0vVYNo8FvcNo/Vgd16hG79e4
Oc/N70VeumWidcjbtzRNk2vIBPeuY/smrWcI7Nw1dTT8zJZn1wDIOyRfEQMMvP90
c57JGuVfPvC6UxEpcxEVTa442VuEv+3xbrg2ZNaUtEozJidEo0pSLa1BWrhWsBDt
7/k4VedlsX5XBmRNZog+3iNOiAItBhLEh9Kj8167LV1OFdv2zRuP95xvVHDBU67c
/zWhusPQaCGkntRhOHDszI7SPaPcpj+5kHZYD7XyKGnxwPaXOdTHXvv7VqOtUySi
vUxKcWdzBwv9+SIC3nVo3NTnOGR5l0+WEOFG95OgYtSnnD9tNuXuAHhMswCvPCYz
lGnYg/gHb5cvIsgxPPmWjH92mPqpGtQDUcZ4g6Z8165GIbV1IE/jjNAfAWi8/28z
Di53vdj1WX5SPGetx3ml6Qq8Y81/2U62dctmEfinvwwhh7zIS18OEPOOvRHvZRW6
kcLpcCziGHGHIvr1A0vJdYnE0R/1fgKtgNnBHEbVhR0zg6G3HzFflG83akcqzrC2
NlNomjCAEo97w5LdGxGGb3RGkxiMwks2S2z9sYa24hhzGGL2x7jsGbCdnYPoqrqy
tIw1ZoBLiCcFVKD28o425POCxS68afjZajKgCcTIS1H9s/MX76siUWYQQKCesS6j
ngHwfqFSKY0mXDHguIhBP/39wtXhxG62y8bEKEnCWbszD7+ogYF3HpO9j3OTICJn
fwLLE2qLR2P7y5CEfqT792OsVC/FeJnfyaBwTU34oAwZ+ejfi7kWq/olEvkqJb16
1z8mExFGw6wJAuulwGUxxHfLjCZNus9fkqjfJOq6tRKMYgM6zQu6cQMzJu9JC8zu
xAoUeFAJP8Lxhek4QrNSfm64oISdm50xjKvSYMHe3kRNRCFJ9mVtjrFXNnypOWpX
eGS8CteZGM+zINbycFQPwsljsNW7wBQ7VCZYvMO3Qk786g2NZnhKFHtcytUUM6kn
/JxY8ASodA/HgHm3HJGWBseLQAfJOmFib4bpCxaSkQn3w5HQNqGYBaGce3PCszfj
wT/IKTcP36GwZ0DjvYIoEoyOLdBQuR+Xm73GoZUv64w2LNKGYi7z+f2MVb66i/YM
u5YdFbVWDyJ3u3e8LOOuWIzZz4IvuD2+OTxNLLZR1LI4x54BFUM0E5kO2fdQSXf+
ccIcbYs5SQix5qJ457tFJ3pHIUvyL/hzoxnkJASKpu2gNQjHXGTo7D2HNQrkPZB3
nH5wv9IYRL9UZk1jGHxasHtad5DvmtCDxV6HdpldJLGp8hszlSgCaopyHI9dIQoh
UHKZyCOZw2XVJ5Rv8MalC9gwqrzWY+QvQ3PbphsgsBxxc8u8XglN4AsVQs+3mly+
QoBpoPLr4xZbiGY77ws87+FeOqDOqnf1ntx3RYS3SByH71fAU//AnqFe0ZlxTFdS
ulgBVNaUfa4QlJN5v/pLydosf8uPzfbK6zmoG7r3htIzYkny5pakRh247N1556+b
AahJy/shFata0MdoO+REqM+uhO74MqQ9riBYu4Ef5XGRAuAX1l8eNAdLZsHfzPjU
nBewhaknEuJGklH0Edlvsq2D7vSRto18z7TforZzV40SkW2aEGyYA6pyVirKG5T7
2zDD+8NmJWh6YieooZCYh3qI+oK7ueQlG/3ypXBa+uJ7ZlKXw1s6idCrSaa/lI9+
Jnpx2mSUqRqCp8jxUc/t8hH7X0Vl9Fufim9/icVDNohaKKoPt6q4/STf7Lt/FE7Y
m+s7QZzrr+pUcpzG5KHL/pu/xfPHuk+C9mNKiJh6ziUGyn3uLXgpP8PNKeafP6MV
gcEmR/FvXE8xYolaE13rLy3LNGVZHsb9EgGwUYf9XUt6/GTjVOl5uJGnb4frlPpT
j0vst6lirzptlhpy6xqoRBVuE9jP+RImFGG7SK0M9hzm6fBPlKDHtNwZXZSfFuBj
tgZIcXtImhKiZ/eM1adD3TkeJsmA/VAt7TJ7iIELwUcPrTyzDV/BUhQEZmyC2ANP
ShC/Uoa8lmXgXfaELbR4nwWCS2DWIO17uM661bTxDr8zNxLGMjBwKOrxrYUgg0Bl
3jlpcSOVSNGoc2tu6a4Qx0qyJYBXjFGGwnE588MAz0bF8hTOpKWoJ1mAdoWS0T8i
jOLuXjCJ3wtuJeTkTFVEUQhTuowwfA38o8lvbFDLIBMP2KluWA82RXOz8o9CJrZd
/bPP2ldEH9ylzhlDE4RR8qPZWICcwTAge9kpzv2sESR80zD4dIkWX5eP3GjXhkTl
pee/dLaUAynUBbjB39VNvKTUvxAnjM0B3vvckoC7/WU0oCbXrL/BUSoiWEwrDCJZ
yqYDQfS4S9pYVCSDZmin3R46MzM/ANbgzDmJpt/BqPZNm7aXRB2dbcANj/Q1lf87
wUiPiRNnrhbU++HGVn0Xmc6fttqdt1EtBajq3ucRl5HFI0gKPG8zuHst4LwLQ31v
+VlR93bxb5EEY1PFXs5uNT83y9+ThVQaEHo1lZ9sQi5VYBTMfmwbrdCWM3Y3Epjp
UTx59KauE5p5pUDrZ73Q86b3DUV5KokibwY1Nt68wn4+0wgbfNp7xTx8yMXNCTiz
N+3OktLCBe/Cjmw/4hUh8LZfANezkFPwS30pV/nshlekavQjC/ecxr2JrDh2Lr09
/no2HiZJcOpL86sXn2P/T+W0hZLPRiTV8W9/e04jmBPBuhMrMfhOqOK3yUtK/t97
wgwtA5wbEpZsnnkDYhHRtkimCs1RH8neS5rnYTYR4u7cVqL/TJIHqUVLgCpNy3Mx
RLd9q8VRr1oYo7FbkCx+0xI3Bt4IRisVeqJY2ylh4ajkHyjRU6A/lQfKqO/h7XVf
rhEhif558Oq9u8q1sE8fV1++BcG5e+hdGYY/ZyC42qFq837olrXVXDpWkkgMizKu
DsPirT0eGVI085cVlkomRsYWtIMz3TRrR8dpVcnUqp/jei0qMqynvnOZKUNlJyp6
zmJ6iysYOZdYbU+Mr38R6Io4k0Zq0nW6YWBZ4Z3ucAkcIE79WBSebBLvwckkYK+p
1PZxJt4/nIzx+z0Cw0864ZK2FVxPXxKeXyCzYn0agHtkwvT0syNwYODBav0G7t7x
cCI9W7/MdOj+Zfgf1VPIh8YNCv3NPnXZFiEJUkz6wIVSx11L7FqWm7shJk33AqCb
X7UcKbah1PNVbDjpjc+MhEAZnEQny6nIxwaPAT3zoK2clCHfXKQYCwjD9OzBVs4x
+IF/Qy6eXo9rdn2Pn8fh/j9viyCapRqlIIN4iM5L0u/JkhChqxhk2EdU7XK6xv0M
NnIG/70UmlboUDpneGhGFqkCAc/45eY++ZaO3PFtEd5Y0ytdLFSVwquohgWqd6Wi
FrgV0YmW/uGSh4iqFP+GhGCH6SbkgoOE0FbINe6H1BVvRHB1SjOLp1E4cCw/m3X+
xtH3iTuJl6iodel0m8BzQmVNiXGgsScYd/nqYs0+aQhRvZBjT8rDj/wLphAYZNn7
GM8TZFLMOMxSqxjl2bCPw7MN1b3s0ojOmdBvpm/nGFoQLHVyYK/aYjnPdhGvDTfQ
X3fyxULvwB3+tBDOckMzqJb5wkn3K6WlC+Q1n9dItv8VJKW9au1SjcfETHBXwVOk
wOUVVft25QsTBn3O4ykQwivKG9nS2WRiww+4/Nk17rALtzC1VMkGb84TB3l1ainF
ug99AL7OlcS7wQscpA4i6XiHgE4B5HLhVnTJrrEYx8IryMwvOpX1yEnNz1WZEFhP
VBPGtRpOFkR8fUWKkom4f5loL4v8n9dzGsbAIuRfHbQyY/7P146yD4Ia21qMo851
Yggwe8Lj0+YNUgFKPXIbCg4j6wkg/8RPX1ZPVgT1t+grVwCMCeth37pVQSOFlJo1
o5ObYUk95DFzM8LfvLilROaWcaBcT10yrwoFSQXsHB+jIUYYBNu01ZaQjJtenxn/
8CEONm46IyunsIIUUtANG1E0StEsyEnp+C4vr7sN1qhKVtJT1bp9qItTMSBSDo8R
pBDQealmA6neCQRc4jWZPZLNwyrKN4He0xrjPwIgG0blZ/khf7XoK7/ET2LtChTa
9t7mA3jLXSIvDFlvvW8oV7oMJK9CkqIDKxi5yeXB5t3qb4xW7pM6xgxdfJXjlIcR
UMRkjK0EFeG8NPfXInq2Q0TM/herWgMyov9Ps/rSVqMeXuczP9jY8fhajPZ9hiB+
ucEFTq4hZgzbcJbAglhIL7n7Jf+XuaeA02WiWp674cqxK/UknJd1JDnJNc4tLdSq
oa1NxFzHw2rdibZajNGV4r8tKslqn5O90SeCICV1zOc5ps+gpeDSXFPdZFNVDH7Y
GsMcZAahsbQPVA2zdUCLmEuJT9JQBELITRJC0KQXIKJf+UkZnqpDZ0YUSwz1O1Yp
X4dS/ogZD3CH4oph94hOy8R0lDV/heN77pwwkkP5pWcrof+QgIQt1/+gnouBL5Mu
lBy+H934m9WWGxaXL3tc7C67iNUz56mLrS+JGszQric/We/1GI/JaTWcRPmSoYNO
47K0/3mjCfmDZ19VSCge0wU6chxsD8QcSFafmvKQsXG0dEsgDchOLtcQyTvtqD0M
Wy5uqduUc93ezQxJABtscfudyJX4ULoIVU97AhlaHls0Pt3q5Qj7V3RjPtypnYjI
iAk8yZqehjOfIvl4kK/g9qQLtV0ZYSWFtQJlYXJ4QPKLdb8QXET8KRL4C9HGltJz
kDTGFD9h1z2D1XyGYTQiTg4sofeS3ghRVBcS7j/faIs6eUdKYK8pFPuv2hLvPN8u
EQQaxCG+W/aWtpsVXDfpkTzJm7nBA0MtYmcKdck5KkIGx4izUauPiLh+4Tfs5mqw
Im5RLdI86gM2248rtRZb9QUJmZr8LqbR1h1lgluIaGJGRbgRhRL0VgTGh19FGgJx
a8PaclKkYFo7X/bOpGIIOW6fXDMiCo0iIZlqqUn+JZ5+Sko1wtQ2w7RVmoKRbf6s
797KVgMrDCRTpUa5JySPebU14R3gWQ/0gRSGHwBlvrMUidXoAtLTLCJDGQplYdAK
rwoGgnLvPsLkYyW4QsMSYHmolIxouj5jv30sTHOHIbSZLbSsErT+VQCJ4zVo4MvG
8Qwg/4bKiYpOKUrmGjv2oRtC3PmyISqQxjCdp4ZUMOTfs9zgptnICdFlygLJtTS4
PU4Xg2iexG6D4zLfKx6PdXFOSJ/Ok7e4ISfmI8Q1WUxVOpC+CWb/6PjhwBe3tfz8
eX4S24ZCb4e0jbb7VGkGBOniiSJpMvhGmhTRCAt4JjcA3LmTRoZbtD7FrATIjuPo
GSB30aPasceUR/7aI/ZA2LUi2l/IvgxrWurmx02F5xjfNdA3mFMvHE4R8yd7XMjm
ELztTthCfbn9+YBqumBySpXs+1iDtScwY5VD7Kt41sSOp8jMY5SK1WnFr1GSQCWT
Bjqzg4VJyoeNcRmpuo87vqlYTAWjxBeZO64k2cqTbsbqdS2o7xGT+0edmARpBK5j
zjd+el6KmCdpk15oJpDSHT6JOMEYH0VuVV53tXQ5+lLszinSddgLoEJJk/0dQFXx
TezPbvYetliWQWZDB9bu71k527aIIRbzk7/vgy19F5md6xOmup7n1ZREtsTdCXGf
24IJmEPWHqR1lkJsuOAWWTjVYqXPT4Ip0KM8N/KUDVi1zvz++p/URes5AeGctVFq
9OSlhHhJRbsMAER3ZCL1lsH0t3Qu/ziuG7+YFOdN8tvnFKMQmNZft91I3O7PmCTi
IqVTWoFEzqi0EGbj+jDksgoKR4rtEB1Ee1I0VQOadPQstvV4aGDQNVL4dpa2hfux
VeqNnN2NlNotzVmyS+PEOQdh9q77fgXVzpvGrLQxAklyZnC+lQa7X6LK/6X4JcT5
7UeQhHUcO7S8jgiXPghE+819y+iHMz9QZjfoxyqQKDJFS35zOG3i+2f2/64GkmgK
Kr7Nrsmbo8C1LEF+I8ruuUP2gb8m5U8FSXD8C9cOupIQteK/YDj4lYfdk8bvj64f
orI4yy/UqP1O/VYJGJQ0+2rSVJcS/foJhcNRfpfp3Me+4qlxe+i+2Np3a4cJESa1
RZVWdQqlimuKkjI+qGMrJ8Q5iZ5Pk1u9H9nXHI/D+j7AORWBB3Wk/mljdXuQMEKO
aZ+DjwHMQ4fPSdA6VddpVKMW8E0RuBstdLTGvC+Ll8n1dP5asn3KJ6pef9p6A/nL
ymLCGEgsJa374O5P4ubmr9kIpshTlylnM0Va1wGu0buSGu/tlie5ltmR3wLRBWno
zGVB9LjtNiHB+q8KIjshoLSZ4BSgIv9OoDNBHOs6lAW1UaR+XgSes6iOwqaB6EFt
E0cOhKa8cI97CcXXMqrr/Htze/V3pmmtoy2y3Ws9aja6BqEp/TGIgZyxuEUo44ly
7ut425xoLYGQcu29SlLLtrUFbF7LezN+p095G8CrvigMrdUEKMgDJAjighk0yW34
qOheX2+LeFNJI7y4T5/BMBcy+uc5WbkwlGo4WU3NcvOjvY3iAfHAHshyvFEFiGzo
Rl6Q9idECbCHqU7CG5cDnLEcjSB+jspugRZPVSpMXfnZ1/tk935IW8CMJRIQGsbk
4xRHJGmiTPyYlvtNFx4083gRE++XhX1YUjqngALeNOsCa5BepU0k5SGOaGdipgXT
h26KOtAoK508KKQDWIhWY56e268IIjU1SC53QeNlCAXCCw0TWjdwWgmrVie0CG70
+uJ1hEeFbkh5uexdIBZtRf3RiyBzGO3Oi98zh6tafswBXVZwUs78vJFA3rsknwTp
Op1ThTE7rpokx+sMmha6tYJypJNf+I7KJ4LxG8JlJD6HDqIErq7NoRQCNlk2hfKM
b8QYgYV2dujoiDjazj9kIc/a2SswRReraAlXDUUlq8crXlJ2aq3LzuqQb/OfMMSL
7kH5RP0Zry5HtXGM3t1f3wRTnOUU113XLRZo5L0UhlcGgvhUc4SklJs2z3sdoDIP
VhtcLtc45op5nPv4QIXUpnfdXi9y5j/ph9lBW18+ekLJ0mAEnzvwKx2831U80lCd
BLWF60UJLCiY8yyREOgcNFYqkJ+wQH6/JMauLQnbOZvsMoI6R4wDjorFajGGjMb4
AUALyCkkK+GNV30zciIJFbL++HDtif2nN8KWyXk/FH4B++94vGAU6qHbee6j8U5J
CQiTSGFYet/QtBk+2M5NZNy15LUpK1grOa+eiQ1ZIdZDHKirFuH/voUU8rmbP1C0
lK93fSmOQ3CK1TEJ/Yw30mPST2+HqlXueTuMZPHSjVkXCYB2DqAAn7ucrPrEtxG3
TiUfaooJb4LHQVuCG2SSNEcQnFpYqs+cKJhNXtfAH1FjwnX4BSZB8guGjqYWiBhZ
zOS3eLyvcQXKWRtclzWQYgsf6gAFaNVo8ajbLENfyG91TfsJDxTeNdescbbBupI5
0AU65NKjedZ4tQG24yRF2tviZftygeHetcysuMoQrkcrXk806gal0rQCxepIJ5DW
Qn4916lqfDxif4kcgEIfnbJ8TKK4MOy2es74S9BV9BOH7lVYe7fU4idp0hkELgxI
MkaiQOpvyJCQo8dcUjt1xHdbeTOSSsocL76GyfnI8wWfaKjPNlftyRpED8R9oMnm
wPwNVSEqcGjCH7oTb02o9Ap3VFJLAIGnGcnveVVzyGHKD2QmjkT8bdCJSsxDN2Z5
MsyjizRaqa3YW1QQd68dUmMf83rOFdqBdmNUyQUf1HWbQsvRz2puwrRm0mgPH23w
LqY6YLETd+uFcBtrPOcs9oWEsW/832OgB9WwYuyO6zD74lg6ZrwRcfAW1yuZJ5O2
VlRb0ZVNJNBtPhEcdVYu6Pie+tvqjMVAC5fWmnu+UDD8CbDmi/hlROeNiYfqBhYV
roIP5sHDyM727bW23henwA7ocY3x1tzhODVPJWfa3+HMElYSRAtBOCcnPDA5AsvK
ku7m3CEu6xD3u5QBrv6PhUqYh4b9YDSVEh9mWJtJDjLpz60gZ3C2qqqCreUtiOrs
o2l34Upo/KdIuUBxRBKWoxAv1WDzs9JmNGqziiDtkvW/iYPKchkrv96K6ZjTxxJA
dzZGX9l0PapOnZ8WIqvrnHXMaa2RVsatuBc6OiLhDdVCAl2acouCFv7DR2tafgj+
7Wc0lkelw5jvyNvdI3BxQL29xnJIeQpjYOkg1VzDf2Y/uU8/qsy2NBzRMuG2MWwy
wbmjCDXnUh94xII8iKYVsMBGX9AS4wiQxCtXLV022954eyY4IvIqiwusVKtRVgnV
WqOXS0aR4kmzIENOxouJe5YzUUaALrM5V+G1bT0kvJ7EuDGcYUcCoRxP+eHUF7j/
1b4pXpAh4W7woiTpPDgVLRJRtQ2hVaqPMCI2MaCNLHBGL32mADBSsW9FkrnCh8N9
+0ndlCuoFD9D/DowomRhme/9p1WhBqct1o3DLkhh2kfY8BsV50jHvMw2eoajtpzP
tBgB8WALTFxSu3XYMJ5jt0oXzosMNr4O+Y/dlHJAJQ4pewWthdJPMCZBJPCyqYJw
XfRfJ+4WZJ2r+TRTS5LaihnVKj7XWhU83Ya43sJLi8pNfIi8S8z0o7zRhhmpPkcG
Bdejy7GtB4EkB7OdrUar07QUqG7Hmddfe88d0M6fUbJCppW9lj8XcVpOutepcZc0
+GroS1+aLICbHY9USFN002gJYFaU/yhV7WZmkhkKt9iIjHbJr4yxSBhI8Hw5JEk2
lL84PshzLDyxhDYxUieyBjEZXLbm/FQFSiphkRErKHGHnWTEjJOpLevhqFd1HVbC
XIeh2U6gB+UZtfLfTOXI8KU09EIwdEF34V/4cAJp9joJrhzyvidyswHGu6wvSSpz
BKPAlTiAmgmnbJ/7mXKCkdwg9qroKmVxSXYlqeejkkhI+piE+nkOJMxTAjVPdZzb
DtCtgnOsUu/pwXJkmSRngZvtoY2PeB+5CfGGBXB3iJbNWzDSwKTR8a2rQXV+S0wZ
+pc/S7PWGGvJMv+GJavVws8EDaRjsedeWCGkaLDJs4FiQOYHWpZoDAOziaFkh5at
0otF6vKXZkQ01WDbCfIX7wNw3PGfvxhI2tioGoXELCLlcpX19Jz5dIjXok+jcq7l
WxLHonHW7WB/3sKDwIbpXUH8on8WWtS8WKf1w37VTM/6b+BzqXMt3Mmxz7CB5V10
lasVn8DF9knR6QycwiT2vYK13KiL6Jhsv/Xe/lzLBtd+hwgH+eA69BAoDKohtx2J
27WMIhZFhZg4UWwdq/7OsGs7ORwyKNfpwa1aSmGI64c2Paku2FM7KsnL8Yd3WrBD
wo+/5QrLTER8D7oeJp37+7gU8AfQ2p00i9guQLrIeh5ULBdHaBIJIm7rWZEB/Ycv
IuQ4/S1oT8DMM5gpwttY8xnJ7KU8NfJtrJi6XiTsguq4SYcAz+2DhfD1wTS7Fddr
fKBsI9gd1UPGTDmYFtEvUnBqPwJ0sgl0NbSx9/d7nYeIiHN8K2pE0ReDkAa4CD7m
ReLkEHaVJsczBH0ChfwzVNvGw4RFUidckvLeGmZ/Ww4uE/bzSOMPq6WT3+vGbTDD
k+g2eGj7dCqP0CMK4BDGNFuqVEwt0wNdVjPihXsCuU/XsafqLYhhqCZEfN+j7MLC
ibeKoNyOiImeYAZ7DGNt/MAOI50Sk9KssCpLR8yhTlppziEUd0ys+rS6Zix/aS/9
zp+uFtscgFOp3iqk1vUh+Bs6Ln8QGrRwr2yUiqfPpFeMDCfrSD6U87Bm6ZrEreIK
DCAXhxjTOdmXX1bTXo49pYq/hqUYlkWnl1an8LMPJ1kabxRbO5l5AuBAXCi0HZnr
mpPAlpvvAQG6nUcHC4tAiVjVKF+Jy1hM319jqRcgkbJDuHS/fl9XGrFe285UNnvI
gp4C5sU1AiRVJbpLphqDccwIOjKvQj2/n08UMaA6hJutzNWlIWpEUEC28qfpuJA8
5VFwCMm9oC2RkUwXsM1ePDsJ+44DdkU19nuOBaV0yZb/fWHLiqzZBMNy/muOz7IU
lDdKcuQT8AT9wMS/QGq+i+cbh7umjE4Mf16QKw+I83d7wQBAVorgi82DI8gDEHFx
lKkR4ktawovH78T4NocFXnkThRluusEqShXYHXJYUDi9A2KVyZJG5txbpjzwY1Fx
TB6/LYbsZ6p6Zuyb9/tmEIIfErVdT7fx5gGlmN2GZTvUUyetHDF6b9i944Tc5/rJ
gAMytd8+z6Mw9WIe0ztbI6QoDnaDcjDCMenhJgS1Zh0B7B7vrNqzAuItaCq7aOMo
dIwSkizvd5MfPHUz468eBVkgO10BOlrQEL2Ol9kQ61uy97NPYq+VVGfFu5dU6R2U
v3kn/sUfS2iTjrRYeVKkGriAlVGRo1ud+K0c/gX7C2jcCJFKctXq5XkZNKKdOuBS
+ImDjb9QNBNaN5RRgmOW8Ea+SIKkmn8AMV8Lc+1tJdx4Ff1N2kX9tZCiBLrr7KsO
F7G6mfNaxbKFCE2X1QiNm/MddRbOCuZtrHDUa+N7/ehoOAOmOaEeol3Cs1G1UvP5
kCtwWNaF9a1U9VcXNHJxD4JnRh3vhf7GIPk4QvLeILDqFl+rkVRHfqRMN3Q1MRrG
7iV2jqwDfq3mai6cyGHsMmV70lY6zWUxNWSezHABGAUJH58x7Sir6lPz4fyvAiUH
1oTzOH2C2Pd9pN/wv3YMcEVTfH1b1aORY+SJvRzeyHuMmCGKMbXZLlZ45g975/sk
meGzseUsZnbmVJBxczmM3pdv5a9po5NWy+Y+uQ7vUSwRM5PXS46xq1qVUBJ/JXFX
UGKPko5rQ70Wfu8HYOWz/87MZ0vCpTxn2q5pJswMc7vFzQhYx4gJGny4OhL7/eSB
64/u22wPaXpXN8mPHSUKBJbPYP5ns1Lnt3eJ1xxp1ClzhE5kRulAUF0S7mVDEewB
I54yXMcg0kuFxFmsLJ2DCywQE1AtohWMK832q2YXebPsynjWIfTC5hH0kpo7UmSG
3hqVLMX/CC5990usq2SocN91SXF7/pBeM+eXH3T9Rwf6kGmQ0MlzTJU/AsIEK6MB
hmSKmaxcgfpk+ar+zO2WqQgiYYG4zT1HY/XTrUiRnaFqlX4V/9Y6qcFZ8igc1Uxw
21svmywc43cbWoFfsdJInApc5Ut6p6tvXPrCsFnbzw1tG528xBImb1BEHTWFGkVQ
rkW+KRm1qghdf3PkclOc4sNElP2S1LGnEwqAINOZ3jjWXXI25TsTrgTCmoncAQl4
v7pmo0VcCmuFkZ2BqedFKUz+6NvmnndRo07DOmIiEWvSDC/LwYwKIiCwmyTF3w/6
Qcdk3sjH87iot9HmK/6a/2CqWbbYw5MDrcvFafz6gIDNsernXNQy2LN2XtfTnwOr
9xsJTohI8vJEaAZQWG35LF6nc38/kAbVdIHr+TbPN6DrH3s3c6GNBTVBKk8A8yFm
9pue3E8o0h1e+1DoSxW3W+Et/B/nrvcmIhE/8Zml55y6Egd7KAFsCwW2INEqKY8B
h0n6iCvv5v+tbkEhLQ3iZLHKHiUX7L7PO4lDKDUaTpC9JKg1Gj6BHkQ+EuoJgJhd
jcGBZb1NBQor8xSs7YFH/S1/N+3EGDRioFvT1Y/tb4uz/+PH3XBqZ+ESXCS9T9W4
bL8bY0swleUsI0j6z8dB343ZjE94lItOEnDbBMogPtjMh2XqNc0N87jfJzFZAn1C
bJndcuwx7qyi2VJxlqukCdqmlVz1cbyvl6g+954rwJhsc2Jpx7MulsWdCITKTm9F
KsQcQ2hGcq3svY6OQBmdVGm7S115GlqPcgg1YzN55NEUuiNClT7KO1MDzCbuXUg0
Q6ElzkgmnxehD7ZcHkSp5wKXIDgKaLpoKj4Bi1hqwx+Hb/NCazKPH67LCF8cR5zO
fy/5r3gdXJZcbZ7cA9bk57g9RUKSSrZYvzxYixgxFupdxi8fhb62KmBJAxP4MvEn
gYryC7VmG389d5l029x6iowEMIW/yutwVvDVD/N9STFjKYua9IVoxOgnso5+nhY0
y4YNbjB8OgyjM3CjwhuohxloRk6f/sVSAZ71lMif80ZT2hK7GdtfXYHx3dQ6pgZt
tZaz8zyNKO+tNDWNjBJNF6kiBReqh3MQdZ13orpqTNTZfr+nvLh3FEc8T1xbzlyN
fvORsH/0SGhZ7enSHFlO8ci76tdACbCOVgS9jVUa/UmmvOsB+wX5CHK7YQ8um2xS
LU+sEvbh24WNErBX6TEFnngrC+/kTb3pLkLs5QVEz+WonqWWk+UwSO753HJ0czRV
Sp+xB1GF7TG7VjPd7Q6I0K/DQsGyJ4kwMhadnB9MBhUKluR9Wcz0GdUzgIUJ2C8N
/CpKoWJR5weOOnee77SutGq2NaVK3CLvxpM3CaZA7M8RmOiSaPhPcCeRVZa0zBXO
YJDWPusrGzShgZ6OPmcCL9Zbxu1/xFrOBR46lNIhE7zulRd1vT7i15n34dKj9KLY
Z8ydVOPyuQwHg5DkEXG8MySfZF8k/yoIg4EFRMej2JhenAooBrjuTiMSwB4hvSJL
Ugi91habbL/xqiNyUi65qNmLladLEpysSx6lg1Bmc130fEVHV7WsGjv2WBTvtsVl
O5Xg1CbdlxqmoXE5igLplBtXkBukkDAiMYWUEmXPmgNu5Jo9TGU+hPY2xrgZbEIU
qLpno8K+r1wSCxLRNRAVVPVm0jIrXD+hHjNqheoFLsFidiptnDdYQK2/JbT884NE
vLDtdMxy1GzF9is8MoNxiSC/7GLaKIfyXEdYfdQKD8h4/GvI5d1G0KgLio0lWwKa
IlnaOZ9VbxfQoheROl7aGmF8pJEc/KyJifEy9MqJvJiR4Qw3dsP6RgiLpQjn+SIh
Eh2XbXVGnqga/Z8JC/6WauXRIRyprf24qNKtqOVLKI8ftAuC9QEGOfL66oVycI5z
YrR98YtDWqi40AEOXTxj6N6DmEPT/NK6g1R94AQJzpJqTRC/Ud0rAsvN+y+y4FxK
cmBv/ZCcl9xWxXWrhQ+lHXS5Nuswl8IgPR8hjVlgoTx7kucr1T3deB+gR5VnwWjq
EX6q9vW7ca/P4TeJzOnc/+S8LgQBeiNBY2fEuLrBzSu6llKHeO0D2hkKz1e18G6t
BFWELrhktWl0pZJ0tMyS0aBMvYEEg1LXcKQrDYaxy1r3Kcr5Nd+TcNUdPsePO7mZ
O5eNvVP3VwPYeH3yrw2AedPpy9M7lc9LPM+ZYpd6iHZuJjHA1q7LLf2C2rGlQ0BH
/cJkPP3jtiuTNGdrtJE+lU0KBVNiY41V0DLHttf6UAQFEaOLc4UljYJL12PXytMX
zZRm/LnJy5I6jI0XMKXeDBprwFuhM1aiEq0ig5fjqRVcQoKvz3fscstoaA6XKhtx
w9JxqXecsMvsooA6V3ciopRW+q7R4Apup6fVctG4caGEBGRQpFWqWkqFylC71YcU
g6mi3bb9BuIhy+rINzql4zvqlf2iE62+eneaYN0N0tR9wreUzmbnofTrHxf8aZqy
h4Dr6jZSr1SlW9VadmyFAHi4ltaxHcNwleg6hntekg3gteUSW82qR7kU2Gq3zCm2
PIph0tVsRykz7Xp5ff0knQOrXNiALbziEGOk+oUGPauKy7WKgIUD47phnv9jazE+
MnCz6vmwyok/4vpxvaiQw+YkMzM0YXcNQRBbuY4lzrXR0dEFDjfYS39vjTGNE9or
5ElL7W6YWtnby6EYyOw0UC8yit8LK/ccPEGKP7BcpmFXLTXX7lrcqZRX05KIe8qz
/DHXLT+Ak6p2be0Rs8PYwzyShRTCQYVbfUpQSb/NbgaZdy2WR4qIRZLTuXGbOBXi
n+6SWxtKyykpafGRhrVl5ciIK3O4b1xqvu5DP8PW7xtuqCkheKpc/A8POYWHXsmz
DWpFaYj1u7vt3B6sMarxOpqOkiPeg/TlLAtu1F6AwZGqT8m5huCVxnSWHBnTjbeD
ENYZBr1Y+6kcyu1r4ZOvdtSOSYwyfmuxk9cYDSaY8Zdv4ulPGsQpsFkQBA2qMVaJ
kYNGS45WltGpp+9MPHreixGxoJJLZI/FzKtFYR4EgFg3H9xZx7qmlAEBk/F8wXZB
qlSiwBi9rLj4RyoJTaNYBUc7tzUaAwKCudpPIONehOCKX2LnKrlnirCay3fqaE/A
s5X+WaN8m6KqwzQW7uBhHPi8kBjUv1XnbW+ag/W0ef2oIVIGLulgVYHZSNSgPdYH
0rbX0JJftuAbanhkAQbY6w3HMOmCfjTtVFCbdEjKlHM7/yw/9Ex9Yno7MNTHzWsh
VUz/N6gliEDrOIPROcfGND870UcagYYFyXjTJBtKzjoR1T5HCjkbteCH/zLhB9T3
4CjQ0dBNZR+MfOxiY2EFZlUKMl5ChvQae+ZdxhePZhhaeHzAWC9cYSqaCUs+QW8h
ktXrRNIoR72o5W0lC54W5pn9sck/kYHKtDBMWMY3Fw3wrm2uifEeBz+kWnsgP1c4
BNzDvVpc0q+pZ4Gqgk7VVBiyJ5JTer8nFgf10eVlDUXUXz9dwzn7aP4ttXefBMbc
o6uHV2pTqk3tMuUFg9uSn6Hr9RrnvCwfKoscghOl1xKyd/W0BndFCoo75av1fS/8
BOZkzmIB8KfQEs5pvdG9UL7exf0UYSkOpNKkv5FkND23akxE5A/0zvZ54YdAV/cj
QdoGW9fwZle+SlDCeonpbHaRA3NtlF2ggLpeNry7eXVtzQgIgDFIg9E/9kuA3WUf
BJvgZ1XmMvfG2wDZIn7/SCxmmco5ULyaa1t7I6hTCZWPkQGGTn6p65ys8UorGn2L
cPEozscNHWRRk6KlX7bd68XF/+lPdQM2D6fNLGgGyi5j7fTslko3I+VQaP5kxI2N
LFHpoa4bHgTekUkRVJZBRUjIXa2n+KCi7s6RuvA20gkff6Hg/68yzfOTW6yzF79v
/Aid/GlMBuKajG/xwnIJfNoNiQI7bcUbpUT9VkemFN4N7RtzgQjdnVMz6PHYsfpj
y8cYddDVQ3wkZiCnwT9AQ3HYwyq2gwSzMLyseGasevWODedriAwBt/ANoar366DE
oE+lwRzdHA3UTLb0UL6axAVkHVlXd9BZ6BiP0UbY83C5aBdfUCWc6rMdorwjt9M3
BeraS49Y/8hHXevi0/D8kyfA86zI1IxL1cBa+9MCsni6zB4y7Y01TOiNd3jklJsE
nyJ2sZkXGCwO0t1h9h0cbUIMTqn4oSAwIU+Pn9740rqzbkPjVJBatpZJJWOYqdrd
SIStxoHo78YOBEGbyFEclUkWZoBdAS8wle+IRAptVj9oVzTwa8SY5zXgjM+Q5EGx
FkVk3d71Y+TzVU9VxzCsiRlNO87Jh3Vodwgu3zE8xzqCK4ZUl1mNu9tPyWRXIaDh
DhpiLXYC3ND5Jye1FwVJW9arJIHYiiZl/l6NpXFGgKQ3Mn0naXJqRrzkNWgf2ADI
FEW20NHc3OORO0OdwdKMvKqKaAL+siju0CWjatpVeRAILJCnmWaZT2ET7SzdtyKi
d0iWxvW0JdWEMkweUbK08WqRtMGNJO+qdxWEqwHo3Nlqrnwm6noEryQP8RRgndMB
McmyXwSdWc9jLFb0UHaOZiPbUbQbsIOLnadUAOUy+XnUNC51tdMdlZUf+cUC2rgh
50YpAsEXoDDV6389AH4BY6zF65ennMp+W9n6rjd7bLjL43W0fO77jj+zJ+Ta+wKY
JfFgWJozoTOSgfk/GWMzgaaSO1/zIid/bCU18RHXSP3e6bva2GmyGBkiRkR0lLUv
ksHieJn8wiKLWag/S+3q5Fo0NB2jEbAlmYFwdMrl5a5ULrSR3Sr39+SZs/IiOPx6
8VWrERZnmlFUYNrAhMGRgAwTc3LLNOSXFeVrSpvkT1VJTaLlh6gKVaIIkp+pvdea
SRMqnTPQQspA33IQVTPPKmzB9xIjZWJqUXxO8zQM3RCwbee9miVjYnwAqCf5d2mL
Exnf6qnw8z+0TgR8KhO85kOfRiG/jS1U/gOAvm++cTU150YH5Ykdebma+mCVjJlS
u4LYCKK2oaJZNUwbUN8Q5Um9v07/7pk1DNaNSjIXVS9GLnB42gjN0lu5+D863Yp6
ID+z2C7rVOJ8rEPGGfHYC6qpCAx0Vw3Lq59AFXdUUlAJXk6Dn+l81F43GDTx7j/N
yyLEy/JBurRc511J3EuKaGTPykEM1MrJ7tnTU8iN62w8LQiwdFaAw4TtCoUqTLhI
M24xPtGKgoThVfmhUsCmDbm3T6xp4lxpgAM4z/unr0VUvUJkulbz7PIkPTPPHp7o
Fa7bipPoVLUMKuXIVRFw/DJFobPhTPiKMth5Qvj5oJn3CWE6fVGbE2vpWq50vCad
T40wj/kuE4xDj6CaVto2pLlsK2AMXWxdNgusH1Od/Njon+bF1ufHYNP2dQ4H5XJa
gYcT7NRQKbQJg6nVLNS61RUr7Qbh3RJ8HNiVTC7IZVyCVXXOVnAXqaXAc2mXthls
+Zl5qwvGhSpLAgnTfFPrY0SdG7mUw0bX6vg1BAaV0cCEf/GN6m8Zr224asc7eV+B
G3iZSkfDTDo93zocC0zETKCoika7plzQkSRf83IXYjvikuT5axwmW5NV5pVcacyu
cCxpoaIyGn0aNG+SBzIXQ+sxviSQYWvWaA4/5vseJnIsi1yKb01TZQ8P31+NEZOw
aK0n4mpddF4Bmi9ZD8s+hkBgrcy2hUCgGwQ0tfWXvVaoD8vSYOmxbMTbvcXLckAa
xH3OvAQ2QWk2knBHv1MaD0zJy6xpo7iS/R7SqTzXfh4im/HXo06Sp1UlNbm3v7aB
ton4E+R/5EaRTHnJVkEluXMBNiXkURLmra9/ptJfI8sON8ptjDI+8OZKNuAHJwOd
z/miehDpfOhGlnAf0MAw6cF1rPezxtPhB7gibrB8EiJbWihGr3rlI6x8dzib/kqM
8t/p+6JU6Z6D6gds6v2exrG8AlWdx7lZpAzNt35nZGvTtTuGOzUmvpoFv+1HubU6
/hM7wLoQhNoUq0h+tSSE+PILoohNBe6qIzWvnyPTojSRQB0auejxEioGo1R5jIby
Ro09d+rhNBJVY0Ke9tqPz7LdCQXXMAuIIVz6YUQ0KofaxSZiDbMWXtlGOj43ZelQ
gjULQ+8L5qMMkbbhx3Kiz3IfAx8UosKOfMrsTm5+amDGiEGimT/PwSisJM4eoPqG
c3pKFf+D8gSDt3z6WFmeaTMPGp2WbqD9q7DBTBYx/2LFKA4jrblWXImcTAW8THlW
uL+noULis1R7kjn7QibJrFXpv+ar6cJrTZccFp5rm21lapljE2dxgzpza6+Vnpkr
dGtVtCcs9VVP7LWe4Ystn+gWCIf/WLlbAfENoTrikM8wp97lle8suW9ASSlSqzZd
DLg+s2aWr+0WassDXByz07zVxzB2qyC8z+6O67Yqho/neX9n+qylZpX5lh9ujTqh
uq9TzYsNXw8XeFCawqLrpLhImFdUX8G+P9Don21Z5/GTANWocciGtRzsaPG5KRWy
wqg1lVQ1hCEo/CMg2+XpV7KSth+lGnMo/CEkYwQ9Lb08qgvq4a5vztJgV6PbuOGz
Mgg3OZcmEIRsxDmtMjn1hDLyE5yShfUbRNexR3o4vagRAtXndZoAbc+OssxryIBZ
Tg4QqiWkzLkxLPz7N5i94+1CUMuGO38JVmrHml31z4/nFTMcurql5g9nmtxqQHna
WW4LkeENJTrwU0qEigdECoHzOlo8ztSsmt0a+2J5dkrngiTSvpOyTFBCnVEy2m9e
grYtuFpXpwCZUwN+BXJvvLHjm+DMuCcGIXQSSpCkndrvLbqgFSk+0tq9p5cfsnNB
rYVs+25KoQ24IboVTykG2aOGPoM/Xb2lO2Evy2JBW3F2nEAsFLJfH0P+UP46NjNH
3rstvjSeJ92NWc3/SEjeMviJA/kxKZTaUCi4auC1yZcm3tnOKUK7jG3Z5qrpQ7Pr
vLQscNw36DX/xAHMvbbNHgHxyOeAicK/CPkU/o+uYDdNs//MmPPXO0DLYEG0z0hR
1hu+xIo7e8zy36fe2DNvhKuu4Bm4LKhS71eFB+EHhtsrK0anrg9pjXJWjG5Tx7RU
fEAQcwdB7STsBgngBFSzYIKw6ZwQ9wWPlnkjECNVadNGtEVbGlCgbFoe6aAoexRu
xanzBhwdD0wqCQw5cKkKZeY88Aj4Q4hqSUzmqHVyqkWpPXUX4A6zXwWOU/83QDNt
A5va0qYxYkwIy447Zq5DVh3SnJH3bPJ1DVMgssR0jU7kTWLhrv6rKMRaUoVatFbw
zq4nn5BhZfpZNLeFXPWDYKLU7QU5bwPT4d3ylK8FTVXuHNaIzR7i0CL7YaiS7s7o
5NfbfXCpKgalCpQmPoiKakAkrX+/6EsnyO6Qac4B8M/6FLSmokTzfyS0/TeZll/K
UFgTqWJC5+KeaJu8xIxK8VwhMvz41UEk+xtGNybjk0dTSNy89SOMA5hwKueYdb7N
kMtREeZdl/tiXBhPn1w4Y3oQuC7O8TpmwBu6xsV6kyePIzdqdlWDL5N1FMCQcQWF
Be9BzkgPxYyUKU6160YyHbqT28kpYM0stG9KV6ZLWELyratr2+gHf8yXjXb+dM9N
+BEl4bHVyOGd4MH6GEQqc6cnW/SrejqStKTLMSNPDZBB4hHPqKK2g0wOQ3FZK9fW
Jyl5oDYhrdyWeO3SkA5nLTFGRDZcP57Hv+gWRBPLi5pRhms3BhggjKNA4YEySih3
JwvSbg1nECUSeW0oMyD3DBitdmt+FyGnIjHtnbVaKKWhIw4t0Jrolu45jGlFBQ4T
wO5sPQFcARvncvDic4J4p1HtTfWW/Gig6J3QueHvwty1gaNmhp+GsRFAY4gbIpV1
qeJTfoyLV5pmi3ExLwEuBgf+KfMQgxDNN0v81ua8jcGIrg6NN/xwJDk02+zy3hg8
BvOsNknV3YCeD5JWnomA6mkxkw517lYaKERtn8vHMYBOfg0krjMiHyFbMhytz9SQ
2kiIT57UTW6SbQl334Btkx7H57ZdpH5Mp1LZcxGoUpKqkkqZes62Rjg93TxqjsJ+
M3KswhfDVY424FJPmJ1106soeSgpeoMpdHoOKKjyn/W2lJ87qzRqM+sE8eQ9z05U
e1WeAKxWf2ezFXKy8ZZTeETOOATYvgQsnUSQSjJRJJ5/syF6IkWEiyq9KPUmLmyG
A5tkS69pTo12P99kRPVLFYGfAbG8m/fDH9t+CAm9R4hwtLRuyaZd5Rn9C7ZBPlj5
0z3NkXvvwGs8dRJg2eKq82ijUkNpr4Z51LqKN52tgY1HTWmdOcrPEznCa0e3A1Tf
RnKH22Z6wPL5DhmkNkO0Ibk8IJ0LChSvJzTFJoHL2IodcjD+qF4KZI+3vpvkna2M
TWmTG3feWP+tMu4sC0qby/hXTQ0JwLl+oG5OvyGxE2kKiLJEKq+KowpHlbq90R5J
Ksv5BHWtNkSUg2OnxG3jJkmQZPuoPRzO0Uh3XlNFxsxO5195XN6ha+eD1Hp0bJe0
WPxSG5QW2AS3mVyqaq7q1nx0kpuaLaZmeff/EeyvCFEhfkqCDD70/74IdZLmW78Q
M884n9e7pW6gLkcPxlBKMo9IO7fOx+Y3MKpzeTKZOVwMukPr2LkNVrZVufgr6TfK
jQc9q94oZksiuk1WWzEak9w0FWktASZJVJ0ryFvW32dl6gjaRaB4Go/lGAuo5RNP
FXYjaDmlx5YY5ecBsxkSGewlEfdsVgHMaz7vxPcX27ek40FnwlcyklMCvk/ysUaE
tpq661it/edGUccBSOCBL+9GzDidFzlnfW2DsDCif2AqhUIgSlUvdCal+txAQhrG
14Ci4wFTMHrUZtvahhshAzAZin5lrxLKcb38TkHG6aAjnWoCr3P4ANFLndd4CLzu
sDwO38paSqGg3d5GS0gAcOSi+MLGVemYwK8oE3H6QMzMFtGslPMG+O8dxF17BJyR
D+2uOb3dLThftXZkMqqnbsxtIr6UPLgWV0cUZ1IZlDOV79mOOWmLxwd7ZVdSsHM0
B/6EBkBBDVoG6UQJZop7TwYgIIgxqTca8R7OnbuhoHEYfXQwvhYKK34VPo52/xol
I8Euv/+hRR2sfcl47+jAqgnzx3hD16RtGQAgoVWaqUUTsah7Yw+kQHC4UXLTO0fJ
EZUEfHwaQ+JDRZHUP6AHUGkNr4gdFQGxC68rCv5l0lYh2G/VsvChB+pTKYO5AMJC
Amwg+9fj5bSQsoCGUMeJY+tDbQLHg7eo32ZMXgbBo+uJC3jeRHaKv+ToWslZ2NLi
9+UlEDXqBNbZm54IQONS880pXPpPaE3g9zcQr3/Nvc2nvwEeAjBUp8/aZL9/MeMj
4Lsfg28kgz1HvQTN5I++xwrpRXwaZb6bor87e+oKAqKw2OQDdMLNvjIzx26fIGOP
XVuDedUZvQ79CO94e5o4kgT8fAnb8Uig3nOnuaXzN6NCcaTfAvxG6dcTl3DvrhPf
L4iqYNLmEspXDZTxa+AfY8cab3GCsRg3RdUNB9FgTacFs71LF+IJO1msxklwwzzi
mXoi07RMNBCuSJNoO5v0qu0EAvXkQ8uVJD+VDOHmmONaYbHc9phnW8b1F+Ie5PPF
wmXA37ddNxA6FDf8aYeW+9bM4qgz908Z+jyWbsa0jgPbLTJLTLjlaDV/s0jfa4Va
lTBQDV9c8JxTrhsbpEJphONWJefJQk0ls3crGH31FvFierOxqbUn9RrYlSXpNhQ6
m3fpYDZyfVugSTBmXyQyOQM2czjGAu8SHEO1iKQUrBIIGOuqgsoe64VdeBksHvjg
hI0ZFDkN0tLiEnAAXefDgpCeK4R2BhaKwVvh5hC5An4IHxEQ8nPYMsH/YCW/++MS
AmbBlfWXzdHOCdAdvtwwp7xePzhGZo/zNZueyjzMK/cYrri0ciCkpaVJBlSVfHr1
Om16fU+EqFeiHK1St9XZnZaEixyyaW+d4RAexv/RoRpJ8sIzoPhnC9K2TsoHN4D0
XZTD456GupAAJzt280r9MRWlvZNeKFcV6mCBlUT/VLyaxG4/SSGHyJGmF/Vn9/pw
UkBW5aJ8F28k6jpFrbTM/cETMbmgoDI6ixu8to6u/8Y6Db7MBoxg0fsTeLzwVPQ6
ok9cyKM1iIPlBJJE4qmOJi4W6ghQ1o+GLPhkGviCYHz+yEBOc3cjo6wQ1F7DrJWg
QkbNXEjzdS9azBIg/d8A7sPwFle/nMMVeXPH4LnSqb9Za9942yIS6cvwSaa5hVXm
JcjpAAwQIs/G5qw6Jrf3m6AQ+joKqTnfQQE2j3XjLK91W/mE4M9joM8r/8O2tKjo
A6UzQewlfkbToKpoDW9gPDwMfrkDo+jio84Afqk8eZcVOzkWhApbXsHDZgyqpPCf
RrJnl7dmZFnX/zN3yQ3XP5cMa3WZXQ4TSCwwPGArBp4o5tmO2LQLUwo2kwdlZqP5
iGAur/Exopzy4EycTbsomAhcWfieaI9ExP0MF+xK6dBLWyCQHGeserFFDcPPhmg0
xlpCrydLzvY/wD1UTASx4NDjOzLkO2wzkAcfs/4ZG4ryI6xE+yiDGTDemtcPp0bl
1oqyF8O7zI5rr69s3/FMtcdOUKIQYJP0H98v/wd9vsEWVXNE8T33gFgkf/pRF96w
2DAqYI6gimJZ59hqw+5nOhW2XUoDmgiB8iCH/VUuLKRW5KwicJaDwapb5yb8C56E
OETqI8eBvd0x/dCUJYjVkw/UU0MboxI7cDVvee0kHjIotmnZ1Yg8PBlxJX59sp8f
yXSbboLF0WcRXiLftj+1RZQO4uWYWwXqHE3mBrOm1jEw6+e1+M9TiF0/IBdZ42tz
vREHxZM2+iV8medIwd5nT61jM2LAyx9FshDidQOf/vUU3XjgUpqBf3oXYu0MH5+q
lpi7UfcF4M+9mc1VlZ8jKtzAnEyuJ/MW4kvgIF41Q1kl5SJUVEOiWNxAV38hlfNX
dz+IuW6WA7/HhWlGzHYvg3qboI2zfagOspSkgBLwkJXXomq9EewGmNVSJtGNmogg
A+5t2nvfEpaVNnIhYHaiZhKhtB5iBiv9Qm0hYxAskxx5dAEuBlxhL+oq1ya8Dl0h
HDnPERwBZMyMLzdUqS+QXW9uyBecpNtnvcRiw81AqaGzaCnqsZnLgM9bOvAl9/Tk
CLuswukdMPDVWPEwTixYBls/P9P6zYQhsRxsrW4ogZbNDFiKK0dGbrbY/2RSsqRC
7AympnnJxCmwkUiK3hVyRYtnTHj82lUANPPII3b2eVvHqB04Stbxa/FPZElGZXEl
y4qf5RghQtaRIYfKj4F1NlQW0cFWP86/giQbDsoQeRch5PPmzRPO8c2mqpWU0+Y9
83wsZxheeCzd5MnnJM0RM+mLXjLEWC5nWHd+gxE9lJEBQ8s+9gVJTbaTCCNk/Nmv
wJ++no7REJ2kzL5wLAMbZGLlZ+Zm2kw040OuDESTY5itmNJBChAus9hAiStCymW2
Yb6OvaSml2QE6HITFH6w+2nF2mz9E0tO7YivT9NcMqLxL6X0OtUFfNoFTchuCYtw
PKnu86TAXEZAemUXLm/i6aYZ/tmMVuoOtqIlA4CDsIU1jQDPCEwi2X+QZEQZnmtD
lizduZAsdxoYjv7snSCwfoWMiBlkIEhXKlZgo8cKqAxTAOHWDjEIf2VG0pgzHPfs
RLnvrt9SL5+9Bn+2L2EMzpy27JSFt1QOtYZ4690DyFeEIboKUdXIQ37EGijBEUBX
dSrrVqSN2UTGd0CS9Sx+p25AXSjDSmTgFIGgrWgbWlBI91+Dqdeiqoa4zfrm/zK/
AfPxvPNrkM1iPkG27WbynA+p9F1HnbmLv0geZVl+lbEV6DAfNNXY93IBYOXOqDmh
CRSTMJ42fVI6kfoBn3Wm4PLkwV2y5im9PBQuacojcmkNPSVn5xpI7lrF9gjclw8g
8p7JkYfwXn7s2xnyvNlN4s/rhdprwhdWnP/kN4pAAeBV1zBGphG9taQo5xXrqyO8
QSArO8oZz2sp09yy5Lz8D+67DOCPGXoN3Ir2Ix4r13MfTgx6p2iFeEeGHr47cDZi
EfGx+/GNLITr6wcJBEsvCLqt/uo7Jdo0POa7JEki0i+oQxXtPyZUtKgZ4RSUCt6e
prLp1WK0oDwzVqfo2IswY35eE6JE2ROnCgIw61rwG10td55711V21FNh2nTIccJ+
/zI0kfKgRSM0xEtIa3BS05vF2qJR+XkifJzwP7dKNXSyVofbOdHQC5GCn+r3kjnj
NDchlmlnx0/KWwhpUVzetkqv4ls3pV9scsCOPE9VIUgMcCBdCZIAL1fIvn75yzdH
LN++ho4RLitsh8wR0QLdj9RdYrSlwk3YlM0u8SaFI2DsmWCqn1Rk4d1W9UKUHIcF
CcD6V7QIPZwSHwBPey6aX4d5jIew/kiZQgp0360Z+XJ0/R2zkXjOKgkfRWsg/Aqu
fUixdI1EuPQxkkJHZwvtYQmAW0GYZL6edVOuDVKF5Q1IScUfGYpfNCSlUIfpzyNp
x3G6dMY5PZP4h7oEdbO1tIfyngzsmsWyfGNV1gbCq9UwFvpM5agNRgI33gd2iiH3
jZysgkL2gKU+TKQ7FChcNcR7RlclP+KjMMqIQ2KgBBQDpGLNm7JXZ9Hfle6FYPNh
9LnnC/XndEb27hVfTMkRs3VZ8MJohSqc0DpV4tfZdfPOSm47MaY7zToRRnZtA6VU
E0gvb9gd4OkwByPvesbuPyXf+HsUkQeQKPE5muak67eF5xZYJ3g9xz8Ylo/JrSZV
ZR9aoolKSaWvWp5pLXHIOKa7i/UlzWgQz9yd8Es6wgVxseVQLz3HfqPEKOTg6ZWn
ykKKslwe+r180CpDNK8Ylw4BxSyojk0fOw4fOpW5mh4sZZuoSokkXF1H/Sl/JbIH
Iyi+bhBbkbAyVwvFz9PmGiFy7xEQTCJWm4eP7iH6tL1h9dzEWgpNiiA9rSZw6vRr
k0YpkiuJX3iQ6ZYBvh2DVf/oq0wvEvDSquTjmrvhF6nURdsAocBDUZZMTBtnl5cz
AsFWvG9++DKoj3nheJXaGQR8/4e/EAVrZh+YRqDbIW7EDhmjLpyVPIALR4ILdMb9
M1Oz38feDLZUQtBAQ0+LTg0/cYrINFlB8xzym31C5FVqjA5WLS5grv+0wb/69sUX
9Y/g1kpE8VCFcXIlLtV7XgKiL+w5Z5Buqpu2J3pNv/huvyd1QuMqVEnUnYhXBIss
yDzCPb85xKEENohwJuJjG2m0TyWwPGi3eNR1KoLCPSqNaxqsylBewaUy4X4oksB3
D3xywNjT007BDyudk/zL4yjPB3skYUwwKmigQkSjDwCCxk1UXSLgFUrvF1SWuzxS
WMJXdGRbgFMfBPwlxoqOTjGzbUYFCm9grhmz7UYPSaGCNobOARmSGaJ+Hh7nuDby
pfa8g+gZK+fRKMyw5ikkOYRpku6PUxHmOc1YfqOQxdVfrXhnnXDH+9ID1scdDWGg
K706CBDViT2Ax+hyxfGA5mg33tNO9eXvq9Nb0Ntb+D5YB9c4RFeo8IY9SWIELjJe
0gu8bUccrjrCunv+FvtVtBsrkli66e/N4fALeGpKYfVf8aYcIfKwYDXjheHF+CZZ
0D9HTSo2OX+z5TsWj7b83PEW2OSG/v00nQpgCU1OHctxfEcxofYhnYqYobhkoxOG
Jb3nUcshfLqrN5MIeeZzq4Nd7VLiDs677EU0/Q2qzI85z9BbMNiikYIexwyeKmUG
U0000YCT7+Qaw+g9CDq+mlAroUbX4PJSvTUtNioHM9ngWKXJkOtSTz13OW+DYJtY
akuo4fH43GUvITutloFgW5zIOege13QF3g2ShSmuCrbfHTDYjdwrlvgHMp5hy6tN
Prgz94VjU8hIw4PflD8fIZQ0BX2poONoxs3YCV52D+6RmyZO+zFjgKcI3mJpBCIZ
HCYGRZ4MKWJ4H1gimN08YmPuK0L9s2UOtkJtkXFF01qhi8amweKOJLmSvmzf4jge
HlpJzOaumFZt6KE8IogitDF3xynSOQplNA9srEoDMiG1eji+oJViqljDrWwDBx8r
Ob8HqwSMb0JOA1qZOa197+cvB/W5Ui/9xgMsGGJHyKbczmwjJk4XLQXE9efQ6Gup
OQd/pX08JGHk5IgM6t+4iTJZnxtIh2fOyM9V+AO/gzJfRoYEDFrHpv09/oOOQA9L
Okyq0YxcgOSkB6kGmeNKDSqxAkDgBoh39WEhSrnaqTgLPZhUaWgLzkyLSE3Lyy7L
E7QeCRWBzDO0UXvsNvrGCgUWCfczt1zcpuRlCD2LAHvyf0lPoW22LdbFd77BVJfH
NS9Jg7lsv3IJjp8qkuLf5CvYF8UebtsfnzMX+uSAFbsThDsZpsC7E6UHv+zQtWfA
tUo3kHf6s2hyscxbR4rb91L5gxVAsgE81GFgGUQBoaNUafL3oQ0UbPg97rfruhN/
viDSB1TNKFz7U6VuWelNz57+X4BFnvm98h8/9SA4FbpmvR4Pl3pBt1XJoL9elBw/
VTG7VHKbZgQDUbqJysCqCbHxxfBH67gg/lBaT6JZwLWVBSHvGlNe6Ie+Uw+x3OC7
ppYxtoSRO7aPXPscNGAB4irWSk1N+Ki+4Tb7urcr6Mx2qssfoHyKkEc+WzDCSFjP
nPXn2OYPBysnK7sC7+N94bGEqrtwba3onD3evPnb/obf5jcYQaBYkpBvYVko7SQs
65bzfIjjBWkYuDMdcgmFggaBlGe6NGR/HBUIuTFCVg0liS1VLKRJMZA9xDG9mxqF
nkX6ftt0ii/+xOJGSF9KIGVf9MIVMb9Y44ybX8wwiFMhJgGzNRXnyAsV13pu9hEU
+4/FOG1i4+bfkq/ZuL+9vHXNLp4CngZvgM7QVtyHscdAGysSh+LJ9RTqTMbXcV0Z
RnOX3nsHXDiATlwOxXPhWNijZm0rLT3rDbB27Z8db5sBzDnyk1xLkKrI0bmCQDOD
ugmWhSfQYwq0MVi+CE+OkO3LTznAMPrTd0A5pGpBcHM7k8Q1lDfC1MBNdit1yviG
XZeQLHsX0foEmAXDTpdm2KjlaXs6mYXGU8ntLcFEzzss3gMR64MV0WLPgeAwrwEp
MVSxOqMlDCW4nVpZP04YDFmnGRk95nYxKCVLKFhi7/jDUo/E+hdlh+JL4GReOQ7H
i4HsoRJWuiaXTXmeUVUjQefLGnLnh6CLP0vhHZCzAq8ldw5Fg9Fo1nx+DkzQQa9I
ff4jFCSf98WPeT+0SvyrG2qF6DfsEFJaeCek84eNufa4BJo+I2mTYbYOulJF2vD4
DtSU87FgQHM4O/NmcWoOwS5aAKohVrD7shwj7WU/yyQOr8+Wt22Fu6yfX33gTOf5
60kHupn/AuAIZDHVY2dKNpDaoWDG1GyGAY9oJNXCnVRY8IXiBotlmwOrg+skkXky
sp8NtztP0D+nE7CCAliUShOvNauouhrHV9eosQ7Pg0GH8orJBprCRTlQyljnjh1N
STUe46w/GfUvarHUdQ6ZjK+LB99f9KaYMJQLYl34Con0+X/I7C4D2gr67IV4w2Kk
VFxncOZKYSGtc7wcJYEwbxDdUAhuXgdQGbJnp7QBYH9QSJQrywdpJYmz2yMmz11Y
m7FpsTU9xb1UagAbEQrHI4eivKMAWPYT9ihJVb7MJA9C3Jd3bqCletxWyJrWSHOr
IjpJv4E8z0FdWgG7LCrev4Ns/lKaAMQManMU9rqIMiyaiuDec3xrjM/sHVomFhqg
et5zkj1VYeC/IHGV5eVHhveuWlkY18IHBAXn1zUSXY4DWcbpkm49GIcShHGiK3Yl
BFYcQzTRmu6zexUTvZ1IB+YzN+FDACbGmc+AWoVsffGGJQck+0BBgrt3GOBj4/z/
hcyW4tZpshGuA8GQihjoKOgNjht4FK42maOUre/XrxUm8HgyvV37YWygue2ydzya
7NaJmr1aeD5SNKC6gfjcZ9qiV73Z81hWYcueOaVvbk6PTvLXJAj5NaQqegUKvjIs
7fIqSC9oi7Xmc9jpdah7yWNRSLIYBnL58xTDa8PZfwtkot2zEUmA1TWTPn2N+gWX
Uvzk6Y2E1JTAVsoGmn2MavF00WBe7hZInVTE8i0sfE6i8G5HelsFwzACQDxJHODv
3z0VdjRDtZYkyp3D28gUGTtQvxBHruF08+QcrJrUf2eZ8yUsGGHAqLRGdEJtiz9m
lYGGk/hW2BqpkpzfEKyl+qFsGvBqvVTTi2N3Be1DiazwxPYlHrsMtCTGOpqrL3HM
VwWQWDurheqj8B60j+Q3vCyOBjmV08eMvBNhmc8FfU3UM8tIZiTXaSAIN9eIfSXH
EdJuZ9TU9sUW/j8WDeFD9aLHG54K8vvSMf4don+MRFZtWm704ahcIQ/D+LjFsEsu
5rDi8F0qljkgF288iRBLrm1twbSYVn9+nZXAz4/wovEAHeDw7ZzqPAVmnCPddpgN
sCQ/KYNzlwvdCALs81YxNNy8fLVHk2Yc46O9C1uMtec3Iybvh3K2orkkJOXIMrwX
kGuaCZa78+MkM6WNQF0xuHQLHYrSSpKWo7FMsXOrU+U2NFBah/6PF+QIZk9+lr0h
W3rlBL7iW3ONtOoRnHPJPZlFFp/YuFo86As0Z7t6CYuPq7eTxF38LjJNZV5WR7H+
kYApG8uv/zS5G3xugUhTHJfNZxG+q4iEmaEIYmvNtvGXhDTWEjfGuXoRcjmDbD81
zQ1mPAE3jLcEehc8agRrQYHULkDDGRxnjq1Pj/C6urSIffeszhvVSy8FJeaOC1sG
ti7KXi7Y2Snb7WYd+rxRwqsIkrWZI64pY2lQDfJk/2IX8Ym5wZ25gjWlqNTC47fq
BuPJMhDY+gjD4MfACSHK+Xpc6dYjHYYWqQYcWVykkEExJp329b8vSrY8n8wAUJNK
ex0vxjfBo0zb339p06xC+TE7cv11WLE+O36Lgn/mjY+oKco2aEGo7uhUT5rYXGb8
4ulaQV/f0Rlp7rmgRY1aEQ+SS8a2RGaGh818ezYSCMl+qBLvF0/C4BZpZ95pjoUY
Nu5UaVLLZRhvRfn4Y5Z1jEk7LMj+555tlhWIlMtWCv2dAHxe774MDsjQe/fzZHfE
eboov3L0vYV/JfvYMNznPIugj+GLL2QZWJkPJLe+ZHqhiKdGWWHUA/rU/L0z09jx
1KU8W2hZdJOf5XdvfmdkUL6xvn50vzyo6X4oqf075vcXNvZ88ACmyhT1UDX9AlAZ
dhkwuWUYCln5REQuhBDUSJ5yFh8Dpxxh09E4mzT6EDBL9Qz31GydTbbjG3HGCu4g
H0NHdL8cFA/qxqVqvLGhaMAlzBsocDQjxV5Kuluht/7NQS7wqidRyJhLTl08Swex
4VY2/CkiqWQVIIZ2MYw2wRrZOyZeXvnQB+oqYaZHN9uDVNB3QXM0t6h1Z5XFMdRB
w5X3j+hNdqAxech4VDQrAV4srdUNGKhJ9g8xaoinCyNq/+aDa7T1xCry0RDCoGjo
sYeY9JiimE9OEQBHlCJnvptyUo5+DOZkG8UVcXgz70P4PVftA8nfyL+ln9eoYaSZ
ZP66ksFAr9kgmSrqi+IXwlqx3lnI5YAUVKaM6TPlqiICinkTIjNa5DH6gAlCVXhG
2DDbq53EI+a00ak/gUZ+f1Baa3igk1Hiq3aUIr2GaEKrxb/cACRnCoKaKsxfIlc0
R+Qy3ac7AMT8nzkOUU/16gmkPZ5McBe3cSRmYioYBODXx5jVqpsqH0mIpuOKRImW
pFV1uVjDDmVS+RDHOKLvtT4U3/ZFLvs04Jtv+TtH1NyxoxHPhT56neR2V7NZImnu
t2lexehpbZWcRjquMD1AExlaPBbTCau3AI9MTT4icP9nPTLanzrOu4lWlejYgaG+
84b3cSF0++p3lwO57V34WBF+ROr5SO6B0TThTxyx6LBjMoAn4M/HjI5xiyDgZqqj
6T12iSeJY58LNbvjzlzVHcK2XhpgtLxKodkHN/vQffnd1wwLGMW1psmxIQQFXm5x
1rR72fzBGyiFOx3Vw83z99inpH99qWDvEkqm4qZE8y8bOJsDnvsPZbg/qwWOcc5M
pFCKbLCZaDKB6Y7UCkQGSmx6T5dQHn/JtBOOs/eMric3mwIaiPWdzy/5oLepXvg/
3FVX9lGaGKwsSeOqcPaGcjbQcBhGZ2V6bqJRmxMHwxqSyAF3soh02NAKjJiiYpEN
OQMkzMwOAptRpS/3bgh4ftRgy35Y7Zm2e1QkHLjGmFJgFTaAm9ObuJbGkeMrP+gE
7McV/ofuRDpymRyWusVourqtWQmYZWLH86/sv+HQ9oESj9O+8bGtkbz9dja4gif/
qxSHbZV+poSi7F0Wblsz6c+t0pq94TCuqpe5OV6DOF8NlKZ3Z2UWrpyzZXNRT8eG
7bAqsaOgk+/bmexBd13c8s3S1JAgPWovBePSE+eY5jjwxe7onkGTYHCDaZnUr4e1
vO7RLPKyUvv2TjE/oG7MfQYPbluXxFf0nYFGi4gyvhjF+HTyc9iIZ+BHm09hGRPv
at85F0RgblYCB22/4HROUWfzIrrZaJMdfJ5EHuEHqRwTq+fOlffyHhdqDQ/WKrdy
lT9ui35k8P2I5vaMdOxLDY4D9CwslQFMuTLC/BEfhqc5F1Rzhf0C8OI4KkgRbweL
YGeAPaexsH0GSn252fCFwJXxcEtAMECACOm87qaDlCDDdZ9havFDc+MGgwjys6n/
LsaGvTrNQJiCeha7UJWfnmt7tWT60GE7EQq0Fbpgn3Ockzmniszg8hZfJtHTGTBT
76RsukJeEPSjSeObyvJfQnx3sdoJ2jSqvWVrCd5dQvjEMP+UVd2jnWxvdjggYUXd
ji3SADtQs9rG9QaTuh5Q0XhlFCIUCxCe8hNnw3Eh/LOtT/LXgFVu6aJfCxWgk8i1
uK+I4015/jWuUXwcK7RsZgZGgcOOLKKOsv3Lwl+DHydyBogDPA5maAFS+5AP/Xbk
IGWHEUHqnv340a2pKYYGati+35Y7bLsMUBuT1SfDGBZIasY4QMe5wbxjoAgQCjvc
LQbQPOqR/t5cJ/v/iKWrVj1w7rEjRHY5WIuQ9KTx5dhZoYHGCto2rYkRBbaad0qa
rfOmX2nFGeA0NCedxT5wV8wIAuvtprwQhi3fxyFjBCuGngy4zaWdp/sT096iix9R
vNbDbeY2inb5lTOJK+6RaFyQPd8KMoozXu4fKFIuzz2fv8do5nLz4wBSWPjCvrmU
gkhtxdW1AZ6DqPWAyetLiqHUUDB1Nw98L6uu/wnIoYhog4ejGz0N1nPl4PVyFAEx
uaVZadGHYAd4pFEunqpqkxSRZDhk0NLTeYLd7KwGDvcWFaxEyuNoSZwv0deQByHr
e5BEs9BsmqvBcUXEyjO58qY0Fc5JJdJ/NSBidYYGnMqla0fGdLukW6CxBVk2YJYi
jn1D9OERc7XsDRU3fuwRGtcxlMujw/eMP91SCspfdgPp7YSQcaZkIX1y0AD6qKfE
kPVVtaqEVIBNZAxVF7wWNyHa41DSkbPOMsbBxXkf63/LO6n1W1QBFUYIF+e6efJ9
hprXUYP2fV/jFxJ3lAchdF5LfJfioBlUprJNIszNwOVGCsn90CVm2TNNv2kvrEye
2N4BhrdLQiChQbs4lELNaTIQCuwDurMaQgxUMb/w5H4JvcOyvnKBGToCCfmTYx8i
QtlugjrhnU6yaE7Hq995SpXKiikr4UjH+hz6WrQrL+J1x2IJpuaZXPkcSg3SgATw
ETEI9+Khumh0YZ1eh+CLLn/flDJA2EdsPHUlhkPNnTLuzkBDR/AxTyUawfzYgke1
/ZUmDhGjaPN+JnhJRzdnkG6C6vLtFJoAwB9HOGlg/n7TtlOCEBM+RnHxeSWishdk
Y69chIQ+9f+09whYVTt17RlfHVUKQ6P/sy8YP3f3B055tSdVKj3dhbCkwyqEXcnb
Hr0Bazy6u1GU0osLoO0emdrLXE5m066RuhR8gqyMlcAz4W81cB+RumUH21WgWohb
8XTIAY1NJJhILiTKMahquqyWglLeXZXySqFhq4leih1eUKKcGHhpobV5TYfJbxy5
tjaq5Zhyf5J4h5ua5s8NazOehF9k8AxE0Zgk3QqkwFPUa7S4hcYsClE3yOAveNnV
9dFVG/bSepCzWxPXFNEH0QRIpCgQEHj4R0kpMQ3XfKX58nv6nFGcVM3yXtxL3bvh
+pgZQqPibr83yTUjUhblLI0eQ0711Px1tfnl3kSO4fDHg+DW6oFinfgk58HE4XnM
eH+Iyx2p7lZr4Pxngc6AngDWXg0i3QGPm+h+qFCEEmF3od2OmcvPTcKUvzULCm0R
6rmaoRfI+otnjp3qN7dZAqG8fueUkUAoBiMtJLKUr6CAeHD8SHAHDQaRdBnIZrmd
8BSHNbayaAeoYdSQlIwrB18hv4CAeeOjj8/iIsRVk3lvgkJB6TzNFshtKyY8CS6V
jpq+eUM3zGcI6K4YZs5J95wNk6Yu9VVgoPmu7wDu2BepAPl2ScsvenOjy4te7tGY
uvhQWTKumCfyIqUcPBHc0LJB1XBYusLyBK5ZQYOuUYMsrP3oU3y7rM3hk8jSMOy7
eRZ8kP9+8C27wYiDFS7v8JDWBKY+55O1S7hMtv97yDue/olSU8OLk7schECAJyMw
pw7+fJf55iACwspClC4OO/L6dKDVPtpNMC8Uis4dxmudBaeJQHtYEulwkGfmQufX
IUrbETIAyHWjaQ6lLoza72Ss9HCd/AFlrX5i06VgEsUYTHLod4a1kEpLAdTQ9+7D
KoMkRvcNSuPyiTMQeqm1axFCTf7j53Y/mZvnxDRS5BQIzZqlKj6BdNeg5V+qs2vK
CrbSeMn26VowZH4TS6jA9a/G6pY9ls4IRNrN5OaWcoLN0H//9KMp814nOlKQ7huF
l1kfAhtHDEX69Pvw2QI41wDWiwwMzhyG67r+WxMnjdjwaVS39vYMVqmqqZ9Gov/U
ZpgIjjzWg6hS1p3uEMzKZOEfTFom8ZApnP8U+bna5dtPBL+woWQ6qxrtse0zKH78
O4UJ9tnh6vC0IgfJGz1NcIitOb7rapKU/28YAJjGVvTBrisF5y9UDT9bwADveXtN
Khs4XLdIfZz/WQPjNBtESI1Alcl9kPotE5ASAUOhYJv3qIGWwIfl4y9lt8aSO99A
16wsdTsqZwbbnU+tqyeFs1/uZ3TzGjJ1+KLLhKt3ZZ1lgvBvvmp+SlTjGhCraXQz
1dxsvruRyCPb4kkasGICcAKTgZkkMjsgPkF1WSrhGUAH01l6PQ/FRc1rkf6HCnBx
BOsSvuFZJxMgRI6B4bBAMgHEyaOygNegVZSzhTeoBvvI7rPwEKpw+ge71rmrwk3c
OPDzicCnA4c3RYmDR46X6DwuCezkyinigHcEX8aRbDBlhEm0hCCSZ71Qumn20mec
GdTBYN7ebXdUcQ6z0m+dNIH10kFpVYhbKfTppQkPGFGn22fCd20Uu/Sg0EVmPkSx
pirhj2SIARNkR3PybPxGaQ0nqPwtPJohr85g8Ru6UpXQRnT3Whi8xlZTgl/KAHeT
NG4USwvr6E1NhkOOXv0KJpFmf3BEHwmY1qbcOjMMol4F4dA2LX8cYmcU1RLD3Od0
fB2YhXs48k8fSOwsoYnPnBhcuLvoy+UBM3mtVjAlJsNwXZLDqiS2tgSHLXml1NTu
GVc0DkP2BHN2w2EkyvObCyqfhUlkXZD1F0lZF65h7uPlnXVL+DtNcUoB4uyd4u2A
y5MGr2ExV2CtofzG6UkxM2gRVMhNm9hIDFpVyTk+nzKmQPbdmEyBiMrvbh3v7eHo
q00418u8ppn58IOdoSo9HnUREgjh2+idtdMkObMHsaAPV0lRsVhYywVA6WIah5t3
LHNp8PajjLZNMfB8YSUYh6wC0jW5KbMogXuupk8VVBTxUE33CqiD03UpKzTgtJfX
bRGfaazcvgHuP7JSLd2gSSopaNyFZm7anSdY0T6xaQ7JGYEdWsqk6OZ9HQT5J/uI
m4eNGBx3Ga1Kyy09VUr2Jjy8KcWP0MHSe1KrZREFY0SS9gU600cY8s6tl+vSyTFB
B0MwcZoFKfoCZ+mHxAO04Efu995cV+KVR559DY+c02GOK5m4BhPqx6LR2EW8Hsu5
Ml4LzXf6aWVffgmTcoG2ml66jQqmkWbm1UbIPE69kdBVs9DXsERi0aP6A1soau6K
uaXToKTi/BLHXMTif4YN5hBwk7/zeM1JNtTTVKj3M43Qn07tfOPBhSPB/1SYQHrn
UHUO64mb3TMEhfKt3eYdjW8vAo3dRw26GaHCtziv/CCJzwpOJ9voTQGMv93ppai9
de0Y83t7bKd/Ir06NGbdzF82ydC/10Q/p3aRMwqGRXO/lD1L5Qz6vbRGfkrg68k8
Atmi6FXNGWcosJhKWk04LZw0AFRNe8TByhb5jX+6fezZcKAK7LcowEY9DaUgpLKI
cVqiW6peKcgZhNlKomR401XeL9kQrm/b4xnf56/2eCC7Bgov08DbqdQ6xPYyCnhf
bvF2xHaEWFbFgTu3XIvWnrN1B0qr7X8q10O2AkCtM4nwveouX91QInyfzHKD93OG
QBE97lWDvW/vxfdefWJCNyR1ZIUipDWWSMlJCucEyu2dx+ah4WpIGnZkNIYbDfTN
k0ClZQfsvmk9vBvl2gpyKhmJM7yWWeoH1i0mY/Bnbi9aauU3U9fpYC5kB9cunHrj
wPXygumaCz0oGtItXyqAqueoktw5LkZmXagW+wxsfnpBpB/pBFGZsla6AuCfmNpI
i4CcRm36CRBy+6fd2LPj5oSAhbwvxDkpiZ64wJZaHdWlulA/X+a5ZzmhLkD+zbRZ
dTyevGoSetrj3mU88iNaSYnRD252JrX/398i1mWeD/zkugg4tm3HlW0d3HL/BNxb
ua32CCa5314cODq3SqOWAJZS8sM11dCyU2oyjAGCrT8bSTRcirUsi5ejyNas3HQ7
NyHzOMX5RC/uFY8q8cr53VLcYB4qEZZu/cCxLaq5Jq/O/8txeKMEhKWGKKbxvVV0
xZJ1cf74N2utt+MJvT1xnjrPR6POgMcnls7QAph1BeN1nf/G9ceL2nf/60ylrKnm
4Q2oeZ+ScL8UPDyxboCU21DwTlf6Hwh67oXwhdxeiNUTNiMKjNZdb4kEDQNms77W
eapy9ga4zhNiaXp5abzdSsVDEEMSoao6CRP6jK+IcDdAGEzKkVcBW237OFYSgUUb
vLVw8MXDo0LK/rSil+ydiow0euY856QAd9wIzVLqaKIJ+J9ulrO4MB8+tjWuBvLk
nKu27gGeeblZz1gogRmKL/fVpMycUDEWiD/IX6VEeXoSXJRbuMiS92jdatb3aDaN
KxC78KOHucLxcrUDrDzvpdNAC/Bi10HvdxxWyeD7TqGbUP1z9HFvmeaEctyGCd3h
9aiI2DI4YTbWwR2jwmdUfUN81FYQtKCphS2YIsI7Y+HqRVApGsMUrjHSoQOoVE4F
jxLr2Q1uGNMoHhY8T9DgRkuqcLP4CeUKJ4kJoPe6u+BllZx7pcjHgNiOgViIk1QF
lLULCzy7Y/55arkY9l6w1RnZJ4i1MyfP3zP4mfV8T7VKCCPMQ0+o6zRHvBKzDHX9
MkJ3ueIazuadizKvZFyfGxCD6z3D3B/ndgGC1W6BcvSbV1o4zUaepqdLQ4ZT4ubW
z/5w/BkCthmcN7RBrbiKJ29kaU2lgR69m54G+rnVW51tIDu1vFt9dRM+E0xFItrI
Dx/W+5AIlJl0qjCxBYU0i30G3ukJZRy9kAe1ruOcsNoPFZTerlxKgheh6zrgsHEy
tzmiOpB3P+37COthOyMSNZ2KFbG1tyVljFssr4uEBMbp+2EXt/kz9U3M1O1A219O
3/QtWG9pd1qGt1rrQufbt/sIoKmVccqeQmR85kX2Xvj5iWXqwUND+MUHYj1+0qDp
G4ZrB2Db1BCHvYU+XyiqPbP/um1+wk+uPmrU1finLJ1DRh8Xhqitz8OWBnLP/2/C
fUPLN6gW6EppAMnLXcZ52xnQ/9YWFcTsYSUn4Ilicy86nKXuJH09PC6HD/Hq2G4d
NNOKVDoW/LGCGbjV0iQzDhw8osbYLswJpFFkxRn8PbEx+m+T2bIq++wTHP0MiOyS
+HXspRTg664ebcsEWTIlf/zkjOWYJRnQX/WYIQr0V0yoaZFNJ3FZ1OiFdqvouVnV
iSussYt6bhlmFhC9O9CVClzDIKH2GSDILSN9LbfvIgB3INAP2BpOo59SWgmWaBUc
mSQzaPQNdfktu52XWQR+8nhwLtyDL6c7Edo72Xu53sBhkgmPwNWLzI4IpPP0C7WZ
2H1ju7+RkB2iuoadtEkmGqPGZfnFiYurG95o1N2+z7JVQCrOqVt4BqDLjEA/bJxY
0bkRD8H2vHASeQOMysIXH0PJIY8M7FJWFtxzV+j2VDvPD5TAfSPvxdGPLqDHW8pn
h0q0/3DSwlvWLODSRdRbRJAyFZUCW51lQu57mmcpgdDBOA60jj5FffVCX2CacbQC
ny5wY9h/iRN9wRJLRdOvfFXtlx1YWOVKf4Hxfe/Ys1aQCKjwKsxW0gNa06OIhYmX
mjiNLDqbKh7vUmRG/bHBNzy1XadhDsuzRKrj4EpDYuUVbMQkaacUgCcSbBVrVL2M
439b3by25xaUUqbMRerBuCQ4glMGq1DKaChG8uapNeyUQyJKFhRW7hy5LBAz00VA
OIguG6bOWwD8+z68Sw1mzYkU1W1vv8YtFni84mrKGrHMieKt8F/bqls/ytPjEwoX
uSG/sXexdMh0NMrWJgdQ+G8p7JI0ATZrfzFcp3OAsz7GZh2x89uUKK72OyhlNRPe
r/TdN/Cv55IaZE130zTv6HfDvgGiopxUr3Kdd0KJuMajPvmSQspc4PDAp1h3Uhil
K8Rj1XyE9yi9a+TfJpNfi4EBi/QbyclrO2LxYZirR1MUMEmmOfT9XnUY3qYCLcJ7
ttniZRtHgX0KQQUudyuHVWsMUovBN99hcJFIases1KnoCRdrgX8gplZZB0Ftn2PJ
GSMIchfkuYemRM66frGk18BQ+7swNtSczoYdjnZ41/CzcTpRom5npxqaf6IlFSt7
JL7xSckX9QVexkcVjBlaj5MhMRkVVpkTg3lgsirLMXy/AdZDJMTj+9501DwGW8lk
NHesQAmcXMSFxORmsSzbXhWuJgNKGrjx5yK+/ky8rakxTXz0n8HnNtg7CSG1jSW5
IandxpnZQELiqmmNoNolKBc4ZsMcYmJYFOrU1VBishFTX7XXT0Y9F0fH5AARiX9G
xjRV3JkckH4fSIbPjaf7b5+3WS8RwKMP4P9e/yni68EZUcZAvDwlzQBtKTE3qUNP
h+CrP73/Hsw0jPKWIH0tYtE2wN6tYf6NMFRwio9a+LjCdEmEopfg/apXVwtl5gd5
yHOHyAGI0hNsSbxE/33w5D/96jyLswE6CGWA549966ZF9DB+yQkhzWOrBMn9citz
CcWk6QdbiUaR9WAJzqMdQUqyIZjP6+wn8I6vER6TZX5JY0yzz14Ex1w++gc5hj+K
DBF1kfBNPuJmfFp1xVBKHiuSdldZesgrxCQqdkmgZdWBtu9iQOwVduSk9mPzMKgC
qmWAZA58OthlcEe/v5xSR1NcQYC9PsfL0qZ5zn+LrGPBZY+NxxRRfwpS7gZIoU2r
pYNU9ekX6I84WgGk8kmUpm4ns6+OO+CvOwTKev9mSntnqFZOwenZdVDQiZjaftx+
yUhLhmeBapTclnZt0kOuLtsiVpNXwRin83IVX+LgtWDx9IbN1GoQUXTtgRaMXUbv
SQB8WBZA9UuG0XqVXbxQ2feKYxA1S9cej7M9EDwrkrgjBK2FmLjnOjbjSkmLH07y
j5IrewZatDGDl8PaVE+H5mFEKdPErikOasnsPPVGbEBg/EEbBo24oSVhATvCXMhe
pcF1hDWLOkFG/LV0BLDNPHvfzvAt2J2sHFKrMIiNWaaBiH/LnmbI5M36gkxRhxgk
+7WXCpQ/QAX00dXM6chfR1TeZMTCRI0HURya5BVCCqQSsDkm5lpkd8uM5PPOW1B0
Jd/Go7PWk7QflEywhD/50KLJkw8pzaeEiKuR6jzCS8sX80U3/ohVYS7+93uhhuV3
hTW4NaoFgKyeiUhnHFyOOo5yJUX8LgrLNPbuQmx3mrWxGiQael9xX9dOPY8reca2
HxpoiSm5pCH0AaTA79cU++9EhUIg0GZRKqkGneeehFC9XuYZKwYswLldG2V07A6a
rFvoBPRlJOZE/fu69KM7CkDxC9WEDVObwo6LqsTPM2MLKbhwaNQOCyLyMK16GL7l
meBiGJk/9p7t9aRBexEpyi9FysJgAV/0tWYONsoAP1vlr4fNRJVO3AkI8DzIbmm1
Pfy4n3MAFlIANZKZlddIZ0vRjw7czVEnCiAuTX41xlIYmsndhT9XNM1HECPQqupl
emUhX8LIAQ5v5cMCmpPEr8UzY3YykQm+Bj7rdhKbQTa9fcI7WlfsMkon+GEjmJZB
0rE//ijyl8zBriQ28zRjVvizCa8YHFimwXXJSw1dEGymNaNo5Si4o3xvqSQkGxxS
kva1rrexQxlXs0//aCtmv6X7PRnfpInS8ml4wUJme/OpXV9nxhmfEbxMyqeRmqFz
4BTA1EnBwX3xS1Ukdd9gBUJNEUBko3nR8YyDgNZ6XN35kbWMrv9Gn0lDwMdLPd6r
+QlnuyN9qouH5fmsDwkDbo7f3/G8i9BHIMcFloowIhfq0qcIOcNRrz5XnLU6VIrp
dwU1djT4TBc7SZwrB2gaAOPw8w/LIYKlXL5ZX15GHo+EZ19Nzey7cHZu6dvkZIKE
eXY5OjKkCo3QfPJDL29jsc27o2HIhtohUP+vU3DJS6A//yxcDsOvwTbhktdFjJuF
PaN/STPgKHV/kblQTqf4FFggcM3b+MMGAWSkh49I/YTkv8/CjSbIhUaw79DrmlO0
iAhGEJsDprLqZZUKw6EI9oAviujdHKXdaGhteE9Y5qag8/Sftzgu0rzCK7jPNlww
Y4CCaI+l8on2GyMGS97TrsVa4FqqN8T4WfZG5h6MSSbPD5xUJgBjqkzRgEcFRehY
E1dmzNZ+DLCdA0CADhI0IK5I4bc8FQnREcemPaOnNyiC3ZVJ4OcNa3yjWi4Z58GO
ufqkhnELi00J7/g8XE0rxVCQoH6smT1cYTf0KYT0OtWRLe+seVsZXichUID3++nI
NHzdQuelkYv6wNU9BWrYMszfQQwFK5AD+gkg9LdiCBFhvuLVEyen1AylDLYWPIav
ASlBmC/Ju52sqHujZ7Xm3ijSCLu0r6Wu/IuJq0jog2wdQN4thOJCaqF5KNtJF0Ha
YnzW7+laUINu0FYFpCFx7qY+QnhNRFHNLxdpGCzswOFksQbvfiLK7MN6dCrWbgOf
eL8JnR1DwwZP6r847x2RXhhWeFmCE8ZS65PZK6Y9eWm0Feqs+7eWvq8mLXbjzb/D
11DQlpkG7+q8bHGbIeC5mLxXEgPa4IctBew7DMQjgSI8AMBeNNICAq7IGaEzF7Do
c4v5t1Al+fQ1L5VcNoewkA5W3gYy7nOfH/jWWU/opZpG1RMuVkPW/2xvHBdU471A
p1Kv1FxeAwkzLsl1plcBX3tVG6ITVfrK8jFaCqLluWta8IbUo/s0N5LTFuTGDVA6
HjIH1rR+S6DzTR+myyYyVV7Joph0wGFrxrEQ/NlZMYhzK9Z6R7MfXtUltANNVz23
fp1CyPG1JpNzEk0SjcdsVkDQj1K9qkUvigq75o6ZFPk2f0hEvPgA7Ih7JQsRq3qY
KcTR0DQgoUntuT31zbKO2lz0sS8F1QlS5wYdd+ZKgAFGiGvqTTMXgQ4qyVrpOUq9
SD2l5w7fZAr+nAtb1/hIJbKEGFTap1F5VTCJ2jgQhb3eGJXo5j9ZDAfOn+JTvCUi
O9pkh0+I8YacvoNgiFwvIQBu7W4+7YwFfROKedDsJJHov7LtYrMTvBfnDid0zrJ1
w1znUiK/m0HjCHu0dpBF9J8l5JfIT6yO68prCufu1nOWIHVD5xNs9DzhQqrHxZj5
dfu0IFiBpu/CSUshZqhPuhSzySV9xyFbcFLUszcohkC7g+yC6DKEwkjoDxE8fWs6
aYTzbXw5SqY1ZnRlOhqdnhZIdxF0nwfyLimjEyRGKQu7eM0Nd+l3psBeCNtE3F/z
lZasNSEwioZmaTm/SXKpLh7YskPp7y4ic2/G8bjHLz0loqW16MYMbyXFnQz3t5qw
D9uolXodzV5RvsFOGgW3Nt6vSBwOrXTWB1kbDqDtWmPZgtpttCNXVlGF+ZPMDHY2
SPQ54kEUNJtubUEyBGDNdhcrNhAcvUl57a1HUly8B8zyn7bv2I89jZj5qYQ9/QQi
TrwpuYnixu5RsCbSrdBc2ek8Q1TXgTa20o7DCcqdunFn1ppjFhMVMOInL5BbbmjN
z3T0BAM//bXm85SQCaXTURk4AHjNnSynBtAKj2Xhy00kRMndafINVHI+xEayZMXg
jfTipBLJuZDVzmES1mu4I6C+HIAv9EJOG4NSw8ChnfQKu5X5lGRf+svAUniHXK5Z
Ttd7iHlyMblHyvui4lm0yCsk0rclxjXvCJsH94KCYFuiduDcyrS/lbOCzy55k/Dg
f2+tepNsX8kUOjPeLdGC9AViyvQMuyhi4FS5V0pp1UYo/X2JGSYkkWiuUdCCPFfa
Ybb/jv58Rc/Bo8pvFilLiyCYreZAdAnn1iPY7S2NH9gI4ZRlJRHScBxDwCvH9EbB
J27fLHdloLjkoLQ6rcGBIPxinBIwo8Knpnw3i7JeFc4x8Yym+yp5LzowLiEDgBLw
CSNJdgLu8FkoJJaNhPIgdIU2hficOGynz1ps9GzzZbyf6EHK2OzngipKjCALOUfR
9UNdQ0kyzH+R8EPeUrUNLom7ncSrUiMMapuAAX08AC3NqCD7ExNh2DvqlGIXgaFg
U3d4Q0I2Py3y3AMS7HihOE7x5wF9gTehZeCVjg0wv3jazL2WuxlOQgsJxxr74sh/
+02jm7l2cuVTE404kPyGrCvqY333/a+M1oS1mvBOxkc9qnlefH7i/y38ifgBMUjd
F+P5Pg4vyzpCTFXJ4EpPAxuYyGBaI93SmcsUcKD77f+pVlShodxcqQT245Xtayn4
94TX9sPHxSsg5UuWkHcMpfj2EatcgTY8BQ11o85vNTLkLo8yVrEPl/o5nCj27NrY
mUmpFalDGic5paNmpsYJt9TLOKpOIa9ykTRmlRioYBJVQoq1GhrcQKpNIijCEMPN
F8Gj6xdkYHf6GKBXsxn/t3JTaYISVzT/9tPaQdgbjYnAQ6TX9wMDi1Px2BEsy5cg
/s4dAZm6wji1HSknqhTDEB8W7XZAT3Mu1yof8pHOC9O3MbQ7uOUcqpoNKIv3tX98
0Bwry1Q5Vs4UxfYTxqfHpf+STskTq9u3/9Wiss4lnYYHF6jg46gy3DR247TrNPk5
Pv90g4PdZugAEcj4qg6Aq5CYLem28perRqRF4QlbNCXEwY0nsBKkYLmxG6MD5l5C
+LUWmQfyE29d3xZl1qzLfybpAOJz1UMzJHcr5CF8OYKP1St33taXkP759tK7xqtb
Zkef9TUVhTZpbJWaixKTH+CcKTa6CicAjmOvuECv2vqcI2ckTBJbEA/9DGGlmX56
zh4Osoxd57MIAbjIfSZrkUSxTAoJCmv4C2WStd0sfdwxnvBf31oGETZj8HTg7XU3
0qBpI89QNiPpDsAuQewFUe0MJczwt1aV9k3Eww3jyMxM0m73irM03+bDBKVsPkNz
4XorCMgaPXC2KkF9Dap42MgQHDn6IJSk0CWe0TyopCJ/kpy2kw2gVHmSdEIOGMyJ
QmNBalEXxznwF94RkaEctraXWmQ+6+1uVm+eeXnFOgqLrgMcISNX/PtFlCj4ADAw
vYhhVEKNczrs5njDvQjsphu8vpPmp7rnANi7G8hwncpViuoIjwqM14u8SZG9PpoC
RTe6LO9S9PbQCin8vKEx+6sIK96HPvrdydyaSk4c1GznTm3yfZ8NNqzDsszinf32
05jwrUZd86oAayAB5mwLfDBjfX5qdHpAcGqDSeE8tDKO9yWVIR3Zk4MblwKBIFFn
oEd82Jb8UtSDq0EUrLfeIMVuLgEz4wZpS13dzP4EcSr2IwYGSWB+zhSNXDQEEbpN
WPti0mkDoQNPdhGqiAxmJLwQwoPHrfOXejnGWX2eBadI/+irIkoos/mY+CMFumFK
BbT+RkGiW3dhvvGBoDWdoU3lIyNOnU9b2ESotZn6lh7VMSpSV5p9fCPKLGqPeRbf
QJW3iZqeuOcC/6R5b6oOj/rUeF1RL97KV//Zv04usctdQS6F5GWL+CtzCH2bCgEB
eTSU7toF1SZLuyiJ8rlasyvHdTqjnMMPjM8ZZYYdUJ92jAIRBcpHlpDCVbB6L8ZY
uC9VjS4KMh95azSMO01ZgbrPkKP3iVTEUTENFYm0Kj6RJaQ1B5npUwF80hx6kdU7
lkBUI4oRNwOt/qViYsp+zC4b7RF3gJUN1unSamR/GsQZomNnMaiYrW/6tcnyD0LN
0GLFjRQoPj0ajnt26Gp6xx59gL6FNTE4OBDWrxTU0MwP7c62QoTJhu7u0bGESrCC
voVc9anXKbGeTLLslMqwrr6z66iKfaLBuVrbCEWJDEBTF5nZ6AUwpLve9RD75Kby
a9mD8ZHWmPyRjR/UoyFyQ+NRREPHvXgnFDbApxgB6q+LAZ54fvkroP0KhGLjyP1J
F/zycZoSXRunYM7sRhgTBL3dEtQz5plPmLH9YB7H0siuQ9tLsOqB8d0xuvqlil+8
ELlBi2yESZpSGB4xfrRSgF8fpgbR7QP2GyyvyJ+3mtdFROLuI8k67UCnK4jm37M3
xLSriKk6tSpmPqI3VIUbL6M0QTIeTLVc/p6ODLfrIpTSVKIA7jpaTe3ZirXkgWmg
gTm7c9dj9utcAZvfuGmYtysytAvW77cELg6hodC8iibB2lUamEreh9OSI3/iQvJC
3kyKjt0OWTe/b1ntO1YBGhL1SkAEDc9T9Xu/3nGvF4g6TKnACSVkfh/OX92A6b4g
k3rystRM2VjRT9U5wvtZqA3oEErNOxBeHKsGQikKwND45VLO5WwkX01yPjrpQRJf
2qzDTeGBUJB9l+XXMMn5E2/Za2AZzWaTmMyE22om1mX0pJQ5VI9MGQphB6vtwldc
irZ1ZXEyUIQs3Y9ftTbWv5iw7KSqHxXeIScc3bwLVQwGriujRWOWb2bChLTMXdsC
8okxksFrl1exK/z16lo1yR9JGlASZC4y4W1ULPX/npcyQi5RFrq7N16yLXnXX6Yv
xwkbdppqsUhxf9ts6scNMkBPfCXyy7zdZtoAt8zkUAeyOFM13JoxJnftn3w832Ww
z1aQHYnKXMVp/SqzZjuYTQQZwB4YJtuwDanT/LEO2SwiTkeYQtYmLags+GPbNrt8
v+dp/6x94h9ugxJpVGGIUrYHeXQnCLJzKIyNDBdYosWr+MqK38JmRw0mZgiEV8nN
0v0V+Xat/xJgnHq95El+3tFW/5v5Asbm+iELai9XoG+KTgXXgqmRbippMJuOXyJB
UwUpxdZuoff+8wFaWdN/A/0EA7Wh6xLgpolVFgePOALxUADtqaX2S2g2RYbAyMlT
emnOeiKqGiXjhxCF1bNkhJfeAycs4XxxNcIiFH7aO7teWSliHqYk9yVDOl5Z0F1F
VANkmmNkjA1xAM8VKrBPUMMv7qVerNkbDM+kN9LCm7ZSXsBUQiNa5b8QwvYTeVZ4
lAg+axd5E5VZvLeALU3vXzsLADLsUcBFB0OLrOpKovMWPz2CCye+nnYSb+mTncu5
8Y0d3BEJZ99gYjGWpAhdFqAGQx67p6QTqfzuqlZdbBwKKG0doCXYYi8LeFL7OybZ
5zD4FQlUYFQjIB84nsTFLdnKuCzOiHa81ouFc/lHP8zSXOa5PowqrEGOdp6SGfvz
4BqDZdp9LzrsRD6fyAyNq8HcYgwkBHIpVfBlCOhkGwqSUF789zTFPjMbJHN9gGXE
g5rJPeVJxvNro2NOTcuYtB+Q5oDTFd7gEO9PQZuoK0+q49y3V93MovFxk845v3A/
xxtEag0PxODa5XsRukkw2/+itWNFR+t0GiK2gvkZTxnHontocj6dcnn2vNg9Tzt8
3fIHRGIfxYMVQXmYkJcQf+QJsgATdsFQB5Vy6Cfv2zQKu46TJRUitUa+YTRGZBsc
En1wsQepyiNIeWicDMZ3ajwPXMNi7NV9jKDahbF917KOFOc4Kfwl8xaOs5eE0KsJ
kGfw9gUVieSEXbPcx/BYQoWQnHE2jzrmylnFADO5/zNAxJGMQDe2uugfA9V9Mwvn
yWPLciJT8EroiBjuYjanpAiwYBeJMVt8O8s2GOKaeoNUF9ip5DRUPHK+T2CgCFOR
KlF0vJm6XkuJyFM8RxD8B0CxMIecv4Tr8VWL8f+A3of1sdX8WRxeklknP4eqIP/C
i4rpIuW+ucKvr8LVMZTg54ohJgP9InpCaUILrmxmy/i6ri3rA+0c1+YRIs0aB8eQ
iXfmBavGpQNhmWAOEt3OH5m44M9DFOx49mJbIs9IQQYuoYFTELLPFFngWeKfXKNM
RMTmk8uWJm2smpZP0/fzWoeQ47NNa4O0m2NQBeJdtSlcLQ9/NB2qe3xrBJsmPm8u
dx54Slz/BGhlZnwJbd/KruKo0jclkHLshc90si2SITWPuu7hSIBA/4/pLy/BoJo+
Z1rButGC0Ap02Z5ICngX9g9hoeFWQhXTVlBgIfQYAXLWgNKfHLsi6URAjuGgmdsR
7vdn9eMcnP4GddrpxfsLjN1zTjyIEmBFJhjfApKpltkK/c2clVW0IUHM/RMYTPi0
Dq7FVwFnx6Tp2xaBDn5jbDC1y9rTFbCiVeFV027x7bw7oGVKYVyJiblxv4nxT834
L3kV3qqqiZ5rnBMrJWiV/1QLHx90+uINDTTTPqbkD9FyVPkeqwegp0nAWtFw2Yzn
JbGKZdy9uNduk4XtIDHmVHHY332b5p7B8DyUYLH3ackS9/2GPC7xKvndfwPh1Ub8
R86PFFt9h2inoPNI3yuSzDLmoO7iSSn5JsundnmKlWDOg6Drk26brvJpM9KgU/MC
Y4NoXmlpUu8wjbIdXaCYeCzTlhG5jT483Ny8xJnUPvNSBxdNYG1x02bjQuoXEnzr
TO6Tg3JQG9ymIQM0yWLQDZ0RBDb3F/M4rT71pwxUBWh48oocuzLa7S0gJ2su6wPS
RmHvYquTA6Y9fZX5BeIVxxtrFFOKLyt50NQXq3dL2Ms6GcudNgT0x5juNZGTMiYz
b5UHMxa/VQnaRnitiJGSTvtVszwkf45OMwdRz7EIfUD5kTeG+4qxmh+jwICv33NH
W/wEF0M94arNsRfkTfLo7Q5MF+IualoYAN+r3o7AoGNhqoKwlfkszVsGS7xSLNnY
U3tGj8n7X83lpgcTP8C4KWdOq2ZKluVGvj6OdtfIvlgDb4bmIn2KWrA8k68dmLEJ
tHVX61Azs/nhJvtAS5iyQm7Jxm6VQK5IS24yubJ9PE07OKaxBWoEZWUU7/0WxoPC
yVhVTCHs2t+cA6+fBz8qwZXZJMvAswCcajr3aVYh4zsbPChaScgUEIPrxmLxaIKJ
7O2Mt6uX2KuKQYXaGND7xznAT47EURj0+dm7nGRsLeXfPRRy8M4y36vPaYdxBSy5
V1qdhLqqdHAzE7jF+YZG/Nbkw0mMiV2tQzuLNxOOwyZSWm8c13KK3sLTzwjqtqQu
X7bBNKr6lGrMa7siH0A38hpoqfmun2Erg4+4aU3FBJVN3hZHkD6vEhOjX0vjRxhr
fO5HoQius0Zr9Y+b/GcGQB2eHKN4eXMo2vicb6RO8yApH/9ZMtmgMGfDpyYwW9zx
ifQ5G3JPbUrXweKBGb7o73d28WvcqZ6o+pD7IRbJPgnO1Z6goxCMQMEY2+g3P3MM
0Nh79Cy26A/dhrS0TrQ1rDS+jF6RAZoelbFGMGS4Ck2MvERoOTDAclstmzYBuRUu
Ef1xmwt2VgXr6qnjFeHdkJWZbElxcSJc2smwV4yN+VvrGgO5aXcfsfg99tp6bo7F
eW21ezzKLh30WZZS/TH/1Tle2e32wqR7tJaitmgmgE6W3BW0b9vNekn1SyyV5XbE
+MFuCOiHMl+PeRs/yGL6pkSS+9d5jTEnEP0uOCnxUCeOsA7jySy+0YUxDCgon0c/
fD3R8VHVifIdBJ4E7EtKpNevAOli0ICqjOdj5ZL4k+pmQbM8rTngxg0OfeoEuHQq
ftxDzQGf6mZE4LPak5ttycuzMXY4KXzeSUOSqTPW2CXZSnpENIDm9RjgIfAf7bKu
WdJ2eVA2CI2Q38MGcm32+K/FuxKMdKvAPOjd70qe8omXH86MYkD5sz0ApRHh+dm4
7XqZMBkOJ3SWDDG8ScJj9cFRIAYpq3BQpt0pQ+sMGeQS9WGuGHI3n5PL1cgsRTEV
QxKuKbsyx2G+arnPIXncVZx3/m+KvQRwlqhIRBMQPp+MwuOpnV1NyLeak3c0PYHq
q9OahbEEPgDqqyP8SgXerNDbaAZPRHsdoxb/80EaPpikO+zEx1B9UOJUzGbE/cb5
wWwg12tdZ/IwJ2UIe+3Zh22sdngdEOHfyY1CFIR5bZjx/JViSuVpPmKt13D87d7B
P1OaaS5+n+5W8/gy60029s3kJfWjSBOK6tFNzh7WAUHO5LRfOSIsBREdiTndVcp7
K/eZ6c5CDYVZ5OzgTexD7SBncdc0m5B6p88aOlceGl57NOhZtjszbM1MyaKeaUfF
UIuQjJZNQUvv7Y5TLSpN5wYeiCBm1l/DP4GMm3kltshOLBpPR8F7jt/yuPbiZNkk
3NM51V2EubJ0rCSTJ5SiKpkLF2asuKb9zY/s8qLGwsr1d5IofYu04APCFkJxPcwX
i/vn9/ApET78oLMOj/06YR/supSKU1SXUFcOGGUPd5JVzA6BuTY4OeBAUam7+Z2n
Py4lCVuZT+9N5caswlLx8PkDzMwNt28fJW/gnxA1eZijNvpofXGruCPnCIvTFeG7
LCyWsQzI6q/xUdekiezBHsXX/67+AKd5lGjE1ppT/3FENZfn8ZJGfEtXmFpkiE5S
Jbrc3kRm4xAqyGzAAs8euURtcs7Dsn4bPXAOmunmre3VkEWfxpO4aWsDXZrmzxMx
ewDsxx1LJv5BTMTzxnPnkwLMJtu0pW1CTpyWdXi8+ZvsLLBJ9iSb+SHTRsDSZAte
c4ruiANupsnPnf+QTCvpwTEYju0EmKrBVh+t4e7tCwo6WDx3fapYCZJKmmnIbYmi
nc4gUHiNGLIark+yEJqVhGmNIi7my0xuk5GkWLR/fjna1p++uZBWSwUf4t0Yb0cW
U5Kjs/jJWXy6MMKMC4QmK+DP7DO5cb6TPVCyHXftAFqoaOWCDXGQ2m/jBeGtbSBo
sygA60omwDtLIKWbIlE2XacZRfJRj/p7LYHZgqFbosryuPcNhgTvD3XNVJZYfRjz
bswr9f3qsjkBFA7SymrlsKEHyz19zkmhnRpeWYkBS2qSMXl/pyanxt0pySBpyrpP
LLhu5xS6wF0ifLZ1hFV3RzL25CSXpExY/DstG04Tha3m4AsF6ZWAaPwRDKunIMJL
cNwtQjzxCkxxNHp1OkKM3neUcrhNAo74IaSXDh0yQ//YxcfbGqH9L5KxaxFd9xbN
bsyL6UqAQ2Z35dEES5hyXRsgUMhbTg5FPSUDeanjxbIBM7Y8x5nZpZGtMC849NQ7
WaEpEjZ2Kp7ESCN4qA4WH0EbT2KQ4/5MBwEXACPsVYwx6NAhFSVNOL5Vpt66WJ+H
4i1QWelMlqfxcNBQlw4WTiN5qcQEeVBvtnUj+2AFBwORqGcs0r1D5brpm1K+e+ax
BU99D14SHC/Pj0RXtTPsuT9TyonCkDm/qqBmb7LSzxESursCDPNC916a9tcmgNEg
CBVaJRvpazdfpX8A7hZt9I3ARqoiyHezTdMtmqufStAa+Nb+/PfBEb+wMShZ2LZj
XhizWFRHEDxNTrWPTScRwM8IQuMTA6AecWiPnoIIMML4Xto1y8SFGZC+zdfuEViv
XmcXvwPvxzFw0lJG9/sO2tphODhlZKtsh8AY7bml9yFsU4ZoihNpdvkrCjElNHdI
10YoS/TJnkr6no1FwYGg0CPyiNhHv+zNgIARS2c9zPl1Vo1cHBEljbJb9WUxTq3s
RosxuNAK1lzA6beY9LlWw0tXQan4V62yp6ZmYxlD9h/TzP49X/qaqlxkHzRf5KVd
GfuXCZ64J6DbL9l7dI1Z/MOPuewd7lWhw7u9nl8FIOsjE0VsF3kpjW663n5pqUie
g/40TJUyKTjsY0W77LAUAL0ZSkMcPD5X38+pmRyWp3m97SDeldBHjuH59LgAdA+j
HiFVZ15F8CAojry5UnTKgzfZ8+MK/NVg08bnmTmwtV0hJxhglZjmlMGD+PAnwt/Y
uiRBQPbK3bht9FAfrxZ03BEypp98icjg61G4L2ZSKuJeUrbBCwsGZlpeMZgoTaCd
8ok4A+fDFs8JLUgWMg9SuV+LJk841Ccusw2BBNxMQRp7kLdwQoBjHr3dk+68Cnhb
aFEw5EL2ifJyqRHtk20b+ZEvUB779xuVOMrC7o1UCWHkSGeO7ZdxJdE2ddrVa4uL
kSs2SLHodF2G2gHsStNx/6NXCCYzv+QWq/LyB1mksODnLR5f3d/t5oVPP1DDJ9zy
+dah0Sp8cwSJK5JXHW0s139crdJoBO5iHJ35s00s4165thkVfqultkY+Ik9dvscD
B5E097lqfzZDB79mT0MKhxq5WjEOG/owjkfQIeTtTOnKuUPbKT7Xu6eP6TokoiAu
vSCSh+fyWGpSgW41pGHL4LjICzH5wws1215uQ7XQ4McQI2/GDpx8oQqCrftG52e4
oW5RvJNzeNmM//GDTaTvqqP0WABxtmgIoYktsvui+3a9a0t1/nOenkw7L6aXCEAH
Hw9MeRwWfjU76F97G14ndU2iASwKXiggQycnyt4J522icr6Xi3J8JG6rLfgCY2Wh
+woQKw9WXMCLCDvz5j3L+pkQmpAgC6VbZo2bQemaJ3hBk1DBxH79X58sK1xMn3ES
9REqFZCz9cJ5P9BrL1ifTIvQk6A/fXM5bl9g2Xw+MHiDuWRTWEgGNdJX4cKbVoDX
bg/TsDMZaqkdkQslsof9+TdlghSWBwFCU3MQSVfcwW9edbdeJO1ozRXJoqzvsFRZ
9EmmvKhiT2s+iX6qxRuydK5R11gJ2PX+UFDxvPGmIY+DW+kj7gPtvl+Jkeuz0qFo
+skNo1z4WzUkpLOb/h5KE7TIULYStUSXj6pTrbyFyVOIWb8u0EOjbIwR5feP+f2J
s6tGbyznDJ89N0uJQ96wC06k+l/Lk0TTMmv1MTfzodrKS1xjsRBtfQ01B+CIxd1j
hoLZmM7wNkIQgcZRljP07RzcbLZWRIXQ9Cp3V0+1AEdR8Kz92DBzVxNq9nspnzra
cr8tIykbwZS3e1CoFF1AreYcyYPgwYofd0+Octp3XOJxLtkW1W+HcaeN6JvWCN8Z
tBfVxpZJcFnjS409U97kVKTP/d7pKCJPESn2Ax8A0Euhq7nus1UAMdbIJyEwlSlN
XW17RwSNWvJs89oUFPTxw1uyibHbGnat4YE0ngn/Kee9tHNwdtEmd7rDe84Tw8Tb
c2I7x5hMNrPUkS+NZYjcFgfV4LmcajqE+dI4yBn/F2SqQiIZmFVOHbkJOmrvLTbj
h6OdkwO9OzanAY72Iw9CPQ8JHGK0GniDqzq2YZS4lp6vUAEnqgEf4Q6b+OWUbXRG
0Ylw+hxhGLWXxViW463vH6lL7T4cjdJCXw42k8bPN8tembd+ZWf9v2UFiWxQbB9t
uLiE7QG6DbRxKf/yg9E3TV2WH0NGRuXQsGjvPTgC7D0sovAjRaeEeLafgEmlCIYR
O+kP0/g8MySmVGomcIpcar1K3+pCW671WfqYn7OyRt8fmld8P28I2aH4/IuqiQ1l
JngScAB1hrR9qYl2k1nyczCXVlmRIxR/VkLTP/JcWJbiip9lP5GvzljmJKcXRQui
fxU/UTTq792sVa5W4fxH0G3EBLOM01Z5OcwOIBRajc/3TXahtMBdMAfxp/wjHimg
HiOWw2+tVkcY5qqK3uDqWtQUwGumlleuin+UcAkoyYVaAwQohhpWccRELtC5rRfB
tgOfwwuyk7pX0KnIJ68I0n1RIiPsHVwceX3UM52M63+klop0Naiedym8AcVxdjBM
PUg7q6QawquWaIQwYYmOuczhVOV5HRXoNTqD/Q1Tz7Gl96pnRGdaqw3yanxQbra4
DR91eE08NSWOtvLVQ+NQRzAXbR1/b5CmtjhblugDPPnXapvdmlSYWa8PleW3T+sL
Te6HPaiLWk0ZHoFOjtLGp70GMnFZoa0rWIy4QAGIqBRPYo3gdqSwMK7+1em46yoy
AVfzGyeFnPoBB6cLcNdOOjeSVvDk0UZhWtUPcjobFUJkz8WiBNpa5nwctopGGBEi
mk9qNMLcYOFRFBZd20OwE1pS35F48PDicscQVa3RNrmtewd12+7CiFE1e0J6XLUj
o+xag7HpTcbE+drfY1VGLfSr/eK6R/TXbjHJOXdPawhb+cmFvSfY8p+2ftsJS5ZH
jcJMg+OU5TjDwqqf1GFmJDRYj2ep/LangUe0Pl5M91CTxZWjF0XL/UxmBeJIpHRl
hkW3jo+npjqeMM05PD/Ib4uMKbDD4RO/VT5NS3NGsJbcqz/Q9pOREFiq16t6T7gR
NzdG1cmuheBc+ICwaAN+GBPm4QD3OEv8gbEbQsg+9UKAxAJtDoOeq1bEta4xKv9D
ZLsWRv0EbbvHFxZbT1I4Z60bCQxKttrYwm8BoNbf6CBYNniaTmW8uGXY7ZXseL+F
QducFWHB1Sq9tSY4QrJ2kR2aJvdDxMzEzy0v9DLLiamQcaV6a0OZJrUSmZvef4U8
mRm64SyVXUMl19MpFoh5KsP8jLYUwKcLjF34l11IQ4XVjtStkgsCUiK4skx+tuEk
P3AtKMnaLUd64Ab21tdFBnchGkSI/RhHOdWnEtfGtBXIT6wa4ruDit6e8D4lsWuV
YOTEVIhjnmUekmpYIXQUw+JnIXpmo3tCjMA1attaKzCz7QkWzJeghJ/Aqyu7CLJH
Sx9qOsdJrw1LrX3qPBjSGzeLqscna6l3CyRAff7ps5jT3iCKyGiJs9k5Ti6QwppZ
rVg2bjkvT1JhBTXYFXpnEAr4oY3hThJWuAuw6TrP1kiV+GNs3LplToVhDpZb+idz
xlaA9ZyIH2n6Zpb3M7GOXWeNeaf2vGwyWDEEL4wxTzUWzJVZ2SYq3dOnR0StWxgk
YZdhecUzy0/HaR41IbFxwyiKijgU7hXBV9S9qvohGJTW+Pu/DtClghH+jbHv6JrO
NxnJ8fQYYxUek9NZVWuBZJxLDt8TLvJQS33BQgXvF18VeHl0LWdHfjU0Qx4oH80A
FYjZY4sId49cNVwMZK9xyI3RGYDCxU08jTO/yV7poem9zs0tZiKW2ryf6XVeCHYV
uxPpXG0jkPkUiIpHPM0pptMNdN5WOgg4MLTot/ABbXOdII9+fDhmEPywY6xgL9uc
3IudsjLaQ9WDM1rFWp1GTPbPrvCcvH9a05Y100kgWBhslNJQEn1atoEgBZ/j7KTy
4cNl0efBpe8/PnH8LFmFaKkACAzliD6ETuICpDNguT2dNCtFeAN1/un8E9BRp2bT
yS2ae+7KOL/2+uO4h3+hE18Pk/0Es6TT3RsSPWV6iGPPNScVytLXfNs+0rmDCgZx
SnxBtAnmL1BCS2q/MWJdxM9ar/UdEt4ieDXE1MgpzkvPxlPKDfRRp/1nFo6hPDrI
ZZvixc/+ksb4Vg4EgbPNm1nGf86HQxTYIYpYpz4sIYOfVra77wdBCHK3uuCcaKC0
bJFA8GUDDkGZ7M+3jSlSx3m0ernc5i4OZiSni+QvyYbmts/ML6Hlcpx3OlcpEOq6
PwXF+nXQxzAOTmCATNSsmoO9FghX+k+2uYS9CstMJhcTd7kqF0g3HT1Z1S38GViY
Fix1uKTVp/dOEQtmu809L78H4CUzu7MWKT28UaPzokF9gDceq2155BSVwmwgwEjc
lQe9u0nZ2QGVe/ITRHOzNTlOcwE9Y42sxEg7RVu6tHimiCJKc+kSilsHibdw9BJR
1XX83TX+OmwQfnxYIVulzZUruWR6l8UhJlsnN95a7/moShaEk/id+zXAt9/IEdPr
U9nehWuU8FSWunnVZEERhJP4J0IyGc1un10qQMgfPh0FmSM0lt2j3t+0lKBqWl1m
K3Z7Epy+iZfJ8yT4wEcvFvu+gOJwVDetryGIBM55JeFZXFofFRYuBS3GRgrakHVw
y/XEgyPdR1f9CA4bFxaONys6wjLrFV/UDuoIwJhB9Yh9t/X58Ygyj9FYC3c7aGwx
nrccJBs1fLpqvfY1Z+YHhYUiXL/W3sbmeyn0MhxdmHamy2LEVj4IaExZFKkneCZO
gKcnN6tky0x/jclpwXj6f3LQyvBgNv4Iq6H/2MQbtVybOxJmE13MtgPMvjtAK1BW
+uRjhYYUoMpKSx2S2HmJhIZdHteTd13ub/Uqrf9C6GpoBw4fkaY8enfhkUgZaiG8
m5Pi9IeyMG88rBPfAHuO0Q/vUCa4Oa0Ns3x/E2cKapdcd6Yvs3gCErf710Kq2xcR
qcfED4oQAnRSp8jU+xChJPXqUyQxHEx7dU/lY+ihn6F2ixo1lE9rCWk7Qkb48SjK
8y6BYuAjfrf9b0plOfbVT024lXXCPuXcFwjwVYLHJtwdbdFhQZp0ynop9oOvBRnv
dCQuvrRkWoPSHJRyLZMcCRb1Yyvm45gP3e4amHRo3uJIk5qXWG+i2gFdcmQyjn1F
cD5jt7EGMhKnZ+XG5n7V2OtUN8xy+PgX6EpKDa7E32HshXiLUjo0o+DZ8W5B9iFW
h8ed4LwTx7l3zC4fXOaoNpVEWrIRNMeZFMuMneyzrzgCKJw6TNbLbaPA2SmoRppW
LEnrL6xTWtiDD5mTIuz6o/KU6L4/6Qgdxejgh6XFrnnxoGEQcwU0mhCDmrih3k3f
c7auNU1cOPjWc4zzXfJGTqVruioegISN9Gf/GsenMaIeXC+fIa0xq0zy+mw+ufAk
6jbwLFAt6+rWkngbqnOLj3sDi1k7PitaxKzGGZHzd/0zy7keo6Cx62795qWlkUqU
KB3MumHnh4l7tfqmPsLOnccUzTQ0duOtkhl5frf0a5VdotUhA1PqH6CubPKzk0C3
tjeV9ar2ByH8VJ+J5tDI4MlSostwX+RLbV4276c2V4b0Rbofx2tsbj4vrCYskwDr
vDwvSNE7fL/LcyUQEq7mn41yGFtkBhgPbYhJ8+p3HYcpPs/Rqfyy+g5lrY2KFDLF
UkoVgwb0pmRXsVS2qTDxD25dthQmaGDHtliqIy0ik5KYkDG0HzQUtSv4XvPZ3BZ/
DNo3y9U0nrx/dnGr2zEyxp7bM8NF4pk1RVZdcKlYxF06W5/rqccxtMEprf43w3Bk
0zIEg6ChaaMTQAdNC2HGKP2OAerOXi65kTVbrulaSQ7fxm8IXRQtILfJWUUiE4E4
N9y+36ieyexZsRGLsZ+FEemXlogLGwgNIMsexAb3Pye3rPreOl+5P3ZdSIeWaWuA
dzNr8H4TXfUIIJTFQXkz4tLnbXkmyhUxgKzj/2/oW5vNwWo5K2MRyCV+syziR11h
qhdDccXMOPVErYq2RDVcSApHUnbZGtACrfhGIGUVfoIUZacZZDjoAJGQCENmx+WT
PxO5mk3Xp5rO5HeQtRFp2fNdnHZLB1IfAbX6uwI+ouIwKi00yogcBSW4N1OxrXzy
JRIThCjYRKEqRhYd6FyYCyHR+Nr8fMMUD+LRdUrHasYDe7LWF/XLMPj7P9BXxdRT
ZzXvv9c1mWBZHdEpgdIHTI84PHbAgImKly/xa27tMK7yKRjZNjThIZTrsksQ0XkO
FnPSOP9HbkoJczjCMlFXvL5HHlPJpALGHPLEblKaEV8q7kYfxR6hookD0iGD9Adw
iUE13EqVGZMDAGJysBt1lsjyBfjjpBsdIu6tHEh7znI5d1Jw0XVPuZBEa12HuCad
xcOqvpTxmXRZM+bd6IC7laV/FkkCQYtbYEYeCKpZoje0dEDIV+S/P6ghzGpgYsSi
Cnk0csZDkAN9HKGL6RZ6WZvJh/z2XRculCeP0cdxDlt9iPoFxFVc8yyu5k9hdxW3
LYtONmfOy0zwVe2r6lMStD7maBVcQ0sxv731024tv8ZA/FxeaB+fELab44T7rZmz
5M3EZSagnGtamiAsEGG9jk7JOqEb6gARL+DqULMERaHrrIy1m+9zS51+ryb06oNP
pjroywzpIrXY3XjGiVyfGVCXR0xbjVicOx2+4nQq4SfHiuzRDH9e39g1SL9vdfIg
y195dmuQfdTL+36T3qdAFS9tQIOjRk44sbg4GUgRpFRZPuVWGVC66sVEXzhuo3Ix
ZBzYMRKeeJgPanse61YM6X7iazQ9cSj5k8V86GRqiD9KX1LPRWkyH6ziW5sWHN7p
eLk3o8Cp1tNJLYhMLVZ2qSWXkTFEcFW1jnVY9vLporgSbdDPDidFoqHMcHL10uJ9
jL4fFirmyuc85tqm9s1YZpLyxcK/5s9OuQF5LmfVngMBGhwyq7Yx7h/GSe2r5nAt
fhqfTgTNjRC9O0grzuqAlowcLNVzvzsui4sNlCazqnfA9MtB1IrcCjkmVYq2ddOr
gvyL1wswl/T8zMfbcwv991PrEnr5E7iq++Vj/7JM1Rid77Gj3sCAaTm49BSIG1wy
rxswk5MfKVxhxQ7eJ/pqzVamtdfm3UBdkm+oV4n8/izwhUcpCBNlpILwsGqBYSSl
fuYnGAn+DVbw1jLOt/NFnZeejnaVCt6N//2oZry15y0lIQWRV2E3aOKV4btFwe8T
l8TguuqTrQLqJS7dDhiodE1m3294PC/A18Fgo5Aymsq7zLI4ocMDMroPfaoiTPbL
GuZcX3/Sh5v5XAQzp2/9Z02XiHHD3TGuwBZqlrWNf+vuFMuIpbR1gVSBTyboCxhd
VoViDtgTM9aTOWNG5yhvlVH/GTxiw2dCpBCqFVxzclfoxYXW3Bm489YhtkdwWjU+
Gg/ULbgI6r/VtoUwnatmxjMx2gfmwhyP6C081GLJmN0VHeniwy3GdQ82mOHrrWoJ
hAfXzCkk/FwcHZEwHVHHMA9EK6xSWBsFt0tS1VNBPsz6ZneVgUdj7l9IvXNZ8goh
wka23lqE1GUlSZuDhI8wVxmqBsYcP6DUdp9P8vPyxXFkRiGxM7s57LvaqLSsinwD
XI8hQzOjzHKweo0bzPnX1ACDZSE/VhR1H/q7fl55nrvk3qbVaHcIDQfuTclX4poB
usRYYq8OWM04lLTjB1p497CEDWeztpd8RMGB99Dh9otsBSg/wIcRtUHgfTfTm6MD
eC8F99RQ+9H9XFgy4zaLM3azpB3LjtC22t7uO4Pm3ZkkADyuM1+baFbb0nw/K/Mf
vOOKUMpZ3DKpjdGAoTkgcX0sMeel1M8YkfRf1SCtlECOKiYtZyPrN97hkCeIc8vo
PNU+lTSItotBeF9iYYKGSo5tgZIGIhZnVKoh1ahcVWnP5uuAltLYfPHILP+comw7
3AJXM6AS8mSrk6tXf2s5cFS8ansS7lSDa4XjlUtmd8RpDkCD4I0OKeLaxkvZT0vE
18pi5lfA8sz6I34jzbEY8ywO9K1GmCXCGSFu05mMYEqHOoYcW/Ewk/2H9+LCQZ5L
MZLBRQHtT5X4HLsOKdJDoyoym0WiaGiW0Sbg2EB6ThiDQ49GH3M4kubVznUnlPKe
RhKKd9d3r1J+MG4VoVKlDQvrfXuPQ1E9r0I+2RXke9j7ZLo0gfDNnr0OwMPs32Ce
UimjMS055x/r0cwJqah5yy4jSAidFk4/Dxl+UlxAXuIYUbPYGNFh7n61fchJAOLG
SBZHUb3Ie+uU+6UHyygY2HeN3eQnrrv4GmM71oId03hmN33mJOPZzB4eh+tBE7CS
EuCRdBmNHi5fk4Cf5QQqJhpz/9TE60YgU2Idca+vTfD8afjUiVZgGU1nKir9G8mK
LiWC+R/NQOT7fueJWsQVoVOIv2AkZY31IPT19hHXYIGAN8sfLQSaJpzyL17UkxU2
vW2gh+Xp322ZKPEV2LviXq73lCNrcUxlrQwLKhd2obGxO4RYh17mb20bihzv7r6o
LyIrfiY1AFXb7AraqU3/OMuAHt7WnWCmP0FwfPrzF+wNZNllW9NEu895ECjT05AU
1FqrdCZW9afyvAv4MwqhF3thE03Iah9LIi7bRM5/x8vR+cmaH6LsGwkuSrDjmrXO
FgmzrZHi3oABLeGonPo5DsDqLFjkpzky9mPO9Bozi5t1NMFv1p0xv53VFOQZVJs8
lxMdo9sRPSGhdIvn7sHsT+RxgWcsobN33G08Fmwz8eaC5NgoJanTFxpqz9K7v+Dk
JJGIJ3GrH+IUiw0e1oCCJjkUvlN1dtlZnGv8FQRbu4U/mcm63k+TZM+zADScr+70
O9IyGjf/x5nBrquuLB2QE+hsqwivYzrVx9FBcodopveAQID/OAB8x27v3Ec+Ch1L
OMFbjFz0Z45rpD5QYJSiMgmEh9pl6VdseDsoJDC+7r03J7RGXgIOAliPL7i/Atrf
CTjaANLA4jMMMq+c/dY1np6o7u9eAi1nBv7sAMrHiy5uvr69JTqDqKEzXazUmcxR
+b6+s6+4mcpSRVVPWJQ12d0WERiIbMFS/rPic4V3TykSCXR0F5YTWg8PrQjJsEPS
EnMciRs+qbPEqXlRDwDW/dds4VlRIlufIIeNjQyAcQ8gPj6lL785OnM7oMD7ubiX
HwOZhWY/Iwa9r2PmuFHuJsDUcGJy7OllRbK9pZlqIr0eV8AutfGuLW2BeLLkibJB
zkT5xUYXdwMayK1x43X1Qdr26a6H8AOKhdh3CfwP7J8SDKPfUduSkOS+YlZ9AoVL
MMSjgHXX2rCBt/IJJ6jvRwcyzG5vKyoVmI9rDJOrlmYdqnSsRnkdmazYM2sVYv8d
Tg3C2r3AbaqHS5a8zZ/m0TUI7mtDbTL+xH8o0v9NWdaSuJnPOVhXxX/FUTZA3UJl
qRdeO5tEFyfjLxmowuYOObwKaO8VY5snlgtBoCnMnpObN9DmHzzZpStCHxBOLTDA
TllreHT5cjzXDko/Y8p6UsFC51AS57facKmOxmRxM2VAaDmGMNhe4ONy3Z49H+p+
fyKjhHxO7s+yyd0vySfAflW1qR8NWNiFt6sCFh2UhRHT1OWVSxKOX9G8Vurplm+E
BuLUS7gXLUmHtiGTqPmfRimgsk4Eon+E85qe8hutCCuOMuJtD23kguEMnulnpNEs
T8u+ZCUFNHPosMwA4HufjzM/ESHOTuWGJ0inQSgyRSonXA1SBXaGFEiUQWYGc3tz
rnHmt907FAec7Dwclcm+v2aiB92VU9iIu51S/rX87D9uev+8dZwZlh5c+6u1dVsh
N+ueTWmXdoW0bvKUOHloemBmijQHPlEKH5PmV/dHz5qQ2Qk9ddGer21E47We0He1
Q9Vu4NxAPPC8X71LkPqh4ds0E6XXWa4Ks9x2gszBJ7yldTeeg4nlTV8H1UjryE+Q
53TgR0x3eVh6G2NiELWtkY/VwgCMAPmnx1AjPkXca4u/bhFmhYnA5TlYhQ++gLFg
4lYZtMbpB07N+0ymtzyE/3D6Jg+zUB0zAC+j2Pv7ADt9LM4MbGhxpiUOjOS6mbGd
1tFENg9F1BYP/VL38UFy9Lx5nMKr7mANlG5FUHeW8n6Mr+40LdqsYVenfuNg2ARO
eoAmQKVY0nBL3bMzPSWeurj8spkQIj2AA52Ie9HaWuLPglmmYTU85aCSIRkTWhff
dEN6LsF+54wVCnw/M29Qe/cv0yyiwYqdEcYfM8Ny4SiFHG9pAkJWciO+5wqwlHkO
nH3DtixctiFub4f1x4H4xEPRjInW2TjZuRWxnaWE2K/vqEZFl/UzkvN5ZwbibK+f
JDku6SGAYKyHnY855n30AEoMQeuoi1/l/1Ulu9D855Vbgk22PJPydXxqp2OTXN+C
VPyC1mLwDfhp9tXQ0lWOwwrE2zcK3SbYm9/GNoPkaWq9/zS+og9DYSJoHTQ78Ozr
RinvJ1hyhJqatc7suQfLH8d8KdYHLuP9agPSXsmVQqzGFp7MEVOfWE6IcsiPnZim
XOyfWXUDYLBWyx+3+lHpOcsrxZuBY3zencNUz2KcNv1/T5F7aYupK14wT+vNw6VO
FrulIxopKgYGausL6I7c2v0C169ZI6vlw3mIIQcHptEI6uSHJiR1Ya+5/AzIGoaj
vhErvHItqYrCXZgJfd4I2LyWso1ojTEnQNmrutrFX4hCCqraFJk2BAsvi4HP+gQV
af8wC3yKtvEHc0lgYLcMuIPtCpnYvV5td82V7HxgiXAOXMcvLLimTrqumVbxF8Dn
3YAI4+6cY5xNzJz2DlN5CuaQWbFoWCjnDDDoqB7D5lV4UcdUAZ1c14WxI3vvcPHU
YJIjkj+jKlne0A3toEeAcBuVmG8pfjOQ8L4SgUqNBQePTmF7OS+bkmUiJWtc8Boy
Piy2kAKkelbi8ndygPl93ow5pdm+x1NPwqf7gavhlV1KVxiNZWIBTb9O8fvDVD09
ZqDfNQTc9ll1m1Mpof1+cqa6gRUJRWhPCokgmhafA+XvJP0SMz1SQjdHV69utKzF
+Mcrl/ndOiiM3srJeoRdOBEcr67Q/QdEZS7Qq5GCLQ/1U1DJW0fknV62PScq6zfO
Bc6LQBeOmPqGNV5+Isx2fR6TvMYkdRR5pjmv+K5I88rj/v0AchkaW4UyRj1K175l
FtOOXRPXnA5K1J+NxUs8mnP/DrUfIWN6jqUNjXFrR249IjTE1fKd606QZRkPLZhQ
/B6P5MZ1VOaK2oVqToXfa3fPxrE+j4ZcyVG8vxeIC4gC/B+yGpXHBWLBG7SFNB4l
YFx1Tt3GpCSAcZqaj/BIsmncoIFEs7mMo+c0VprELk6sWeinL1osbJDjaRtEJoRh
sURV7reTPBQm9BpYDewDdWk90dBja7w8fh4JC1UB3Rt3KMr5f5E2M2CDCFM96vRd
RnWS5pPTOh2DmzByzKMf+LbFLKusBwChyypRkQPgCEVJyvNRCuO6h+5xfBwa4+ih
/k4yw9YXyiLArDacCdAbiquKFqDcy5x89A7bYPVLb6v1zm/TP4s2xHGkBAlAhzax
cUQl7HQagx0vAhKjPRptdG5/rmoHKz3jNY9J8pBYi2OY2/D39wAChr8bPuIJicuu
UOX7HFRYShYXN9aRhuWzHnAB7DZgWV5MddVu0FID+Au0qL4cXIqXUmpKvzBs2j4h
ET6v4JGyxNkYJRGD1a23Y6KsXqpFwnDe9/T2M8D9jPvz8xbdIGQl4wwzvn0ljxvi
8nRZfXYVRHDkpAuo3e1v+VGN9u8T6tC/xpK3Vn3aXweiHSeCUAY9zLGB8WZ6TBIS
EYvAGb2E1e23FuacX6JPnGR/hNZS+HCpGqPjOmZbw66GzcQsvYhtyux+Qova6WKw
Wh8q5sVoSnzxh1WUbY8sKjDYynJS/uXBfsmXJXeD/0x5kSGd1dw2zvaAOb9An0vT
/Da6lF41Nt9kUxYWMfRQRlErLJtESmhUGw74PV6CIptJLS7D+j/O+aYqdZbGNSEq
CvkJCRzjo6nOvfkgTcN9NtODcomz+2VqGQ10oofc2o4XFFtqNiIXvdJGcmUj4r9N
kPt+GJ1vBRYCalop7cah66L2bHKE9bLJrwdAev6k4Pvt9DP6SeLC54NwCtgOfSxG
uBPUGxPcc+cDsoFgJ0geLso6TIRLl1RxJuVjD+3p5vdiEhAQC81qB1qz6mDU0REY
HRWfaFzQgapZvEX+s+H7gt2lCjo5tNnLtFqzHIZNNlivZL5TuYUOfH6yvDEDaUI6
MYWRo/23niAxSwCaEuKm63qdBO87Lf9t6zyqVflRXBdw6SCCOkaELdv5+0fQ/Oaf
HxCZpUENaiQv7uEp1J1NrqxTSCuVutM29w6/wXBTJw0Zy0i00k+BBv0zE9DLcBN3
t9SP8G6barIzSszmVvQnILCHVzUDeTViMTvwNsmDJ4QZp5JNE2iXvtAs74VUnFmy
eCCKroBU1Pkw0Ttg7rb6C+IUI09dO3kM9++NfZ7CksOcey6cWvtdxE9TxvLm9HXn
YgrcNXQjaAix9HRsEbKl+2zbWv0vnYQoac3aEIwCTxbohr2prxsG7iZ6gJOBYpFu
b7wpMoHUqX2m0ZLLkRtr3z4fOx9nBKHXXTIhyNk3fxY/mQSj2xydX8hVJlhrNk7A
KXg4hToFXYwQWj7fgEYjs5iQ1WMcaW7uwk+VoJMiYYMxq6GJ+CnSXd1WkBVLljPC
aMMvl6uY1eWcTpB9I9PsPGpzg2XHVR+IcwQ4KF4KiJ+RD3OX/lp+FaN+ZocJMNqg
4RHd06kh9cLqzQPymR5xJewZT0d7/4YByW4Y53Hvy/OnKWaHRgrj84Lp33VNx9Wu
mSokoXpIT5yxT++LhpGMsZm2YHG+BChZ3aRAnML0k0nqHXj00kFpWbrMAsoEGtNp
i6/694zQ9dn5pSXs1TLm9+Gt7QfMztuIVaeExFobhGsYYFEIGEAqZ4N0fuR6oDTv
NNgUGoPflZPOx4MlfSsigBjTyFekk/wRH5lhGPhUMFVptnah+NKZ5EnFjVff+3PC
56wPtr6O1mC58br8lBczhdOvWW6genuC+hHhfZKRj+QXc85wX/DA+/QK1LTyPyEf
oymSOBcP2UPy17Y4vMXDhcmk+zBRh1WVPf/jJlmZkdcBI7TwDV0kDGx+UWxbgwoU
eGjQFgzqVDVrVi+Ymxm1AO+2e9MpEcn3bV1c2uJDgKzdCFkhuX/VEoUmkV65O1yQ
9XzYW5BAlekHogko5zRX9R1z8C5FyKHTlKyG+A1/TQBRuh4JKfaeKb5Tyl9lY7Jk
pFnk19EHhrA7MpwHFOaCx2gC06Gu1MzDYNthBThoekjsNT6i18jjqv+ksv8h1G+N
9vkDFmfu+VznWk0FNg0H2VSD4hJ+zRqssw+f4zMCkj76mrI3YkIbTzWbM5pi867U
IygmEtEHdgxx7ik774RfSDx6oXF9E/lNJNREtXzy7o8z/9+c2ykBs0kT6Z3Hlb02
9y1Ts5ijx4CJImuWTduQx4UZav0Pm1R5ZOqDjdBLEY/kX7MuMqPkLjYm0eZJ+8ez
Lg2OWVNPiN65OohAgd/MXrB4SR/3ehLPsuCJ1SAVLeEL5rd60uTnVUeUiUekAkYD
Mkivg1ubMyjPQ+AiVpnUkKmjegfSn/FnlQyI3VZxyICSabb0F6lhx2IexVFI1r2v
avk8NBtRrknmTvd1TgYrdERy7lRv+hz1E9epUzwylOZ/iHdjIjmmH8ZvfLihabni
Pc6TgCIjJx+n8eAwCKJhkTgJI9bSqS3lNFi1mN9R1zufwU3e+QHIaieDsTSK4IBY
UZWM/SUWuspkSZWUEL/vOdOKu9aMsFZWrq7TSORFu0AuMpOkWDKway4jMp0nNggY
6GD/lhgRcsVQiQ0bQuuA4kVrvZ24xtobwd3Mk8HYYK3bPNBhSjEWyW/QctPKlZ08
OE/IQWRPM5YKHSwmqMuimSmkAuYBFRuH0n+5bV7L6IRCH3afeJfzrTVwe1PPIs7d
Ifh6Gf2DzQyOAjJeTRoJlnN8R0vEgApsrvw0J5i5i/rb9qNfiENI+yCzI9NFWtbM
yfkChOKGWqspQUco661uyO9ogT5WL4b7jjfrboTzhyvTDYajhBGsIVSUqSY5H8JT
7+9TJ3K0+A5WhrLMLjRrBgJ0rCRt4FlplThXXHP/UkJvjAqbkG2k3eOPN36N4/AD
YjXgToOU3MQSNBROfQ8obHX9ehPIqDH75Quz75mAT95XNXkI8GniaxbYTyNH7GB5
dtFqCzPGYYzWw0rZ6kR+Elvyv0sh4D/9lylz/XEhQV5bayISi94w2e5RvC5OpqAx
KVwptFuBmzidQ77aDJt+EgNd/jZ60J/8SvpoWUohu+2hXFxndgd1DD4zJ5Ez6mi5
HvdZ5HStkZo+6+6/XdvEm1oaCqr3M7kp4BUBfas0lCJVfGLucVGt5q33VjJ8c7UA
ILQB1d3DiGAiSBbfzC7aTgLUGu74Dy68N/sg3ZevXUL54a+kO0FOcseFx3qiie46
Vj+kMCsZJNkN05FrkauDdQZqleLLlY1CwKcm6nDarqNrl0r1giUseQ7KevH9Lj8Q
z2i3LgbLIxx6BW/wS6g6TCpySTwcNi9XviDlAMLx94hKUo9ORZtI7sZ4em+qE/ub
yj/sUetK+/zhkXME/95okJ3rUWcfuGhKElHXHhv1fAlSe1/ALYKybYLOzBBBLSbG
d0QIYqDMftnWfpIxoeiLob0hVvyOv1CnqvMG0enTh4m0LZaCIVeKC63JfAnVuYRs
6OdKtyRYyYdrd+H4SnKqiePsWH3cMPFRR5vyFSPJQPxWRAw8ZDRECXuLhoPheEpw
Qi1sLN5W8NP1CaOSQsHVncsrjVFKE7qnc1G9Vrnm44yl89QQOFmmTJOgFEt1fM2D
sbqhaVGSKTGwIMg+dCUJuebqdxvFQ2cMzmh2bgH8smIcIth7Epni6SBuUpyqIITQ
tiA8yOZQGDwKLo2nn8rEJWLlgJpLKjdn5YGA7waOnWOlbKo5pF7uRG+ZhMkSXWHi
FQoiEora53qmmZ+6mhqrtge8CZu6bR83htjJq/6jTgg2iMczQ6wrGHVaPgE3/vZ8
p8d66gp2yhTmCzxqaBHPZNEJRaKwgiTfsR+WEmFR+MjEpSgY0e++z7qvs1+1vBVS
uxDVe0Wr21Dw24Y2sweuwBCKRLnNMWfzSyDGpM8HmGtEkQHxgrNSKaDbMZsGL784
auy7vhE/l6X+A/3YMEWHBfQBlmwZyZqDleCaYOUM/VQTLvs3KZLz/j327Lqlf2hs
zgV1UB0x7mDDtDwv8/PG9CYijnb2sSVkuFE7RxUpw8eLysCbG2PXQfhz+X2nko5w
PIofjPuoK0ZVJ0miGT4oTJCc9dlBbSFscr6eDDQ/wTeJBu0eqdri5h6DVWiiKvic
nuxxdvnz9MtScfhXd3D+EZX7dyH3o2upJk8QWVSRZ5j6YlZItVTDgOBs/+ULc6Fq
Z9KHqDnMKHHS3XIUdI1BhCWBU0LxfEoc3N4LwoXSRZxabPhqFUnyPnJKn+yYARkR
XfE0lOeaBsV5Ze2F+GjIleczN3M79Px4cbWs7rE13LO6/yBfTJbcKH+5gUom1wtv
WlW247eyi7wR0nO+HL1nwVLKZRg8u/RGAbgT5h44icEKmcw3SaLb5BDYlKURBIam
BM2CByCcnEbgiwJYqvJTLfQm58v3+ZTYFnj2VRSRCmvDFZngmSIdSaLog25eRg9A
RAxukihPwMlIRS+TubMHlyRAbaabYHlTuyRJC7a9yDwjmtEpeZDvk0kkirpKBnhZ
R2bAWPjlP29N57Az6SWg0i7L5FQE1rHRGnbKu5lv5+dtE7jXGz0n4uAHOYxbxxqA
R4oxA6Eiy1VLY7U73OxBR/CkbmwQAnjVZN/vKhIHDjwTaOwYLmf1Nmt1Wybnj0MO
9JXpsdDmfPbdE2fI0TxFl6mOvW2ZmQrkwNdZeZeoEpZDT4G5EVUvir4crFcTxtek
dt4LwkhPdLRUwwnaqj8+20mI9tcTxMcPQfBvosEey4vR3ObW21hiEji8IGxcmQ8n
a6FHl/rS/Y23GBPqTa7rtokXU2DYGGSDwjWneT9/KFjbarPxRTpDpVQvg/agwg8k
sZs1lOFswKExY2eI84MLUNxn6ivOsxa0GJjMoebaNKPL13Yjm+0Ffjlj+PO6zJD5
iSqbYdGsXe3vyQLoZtEgoeKA2kwMDkMlNLUdeNOzBzuTM5tYGgNBWS+9ShJ3sINY
ySGWHAxlPhFD2qyu6UNQInVrrt0dxHcenRWlaUol+26Mp5jln5RViH+FFBw76nqr
fGZqcqm9jDg3rSCb5o9a1BK2KlEiWvX3qo8z1KS7MTJWu4BhYPymkM94puQ6qeJp
P/oEqP/wJGBf/xQS0rshK4IKWp3Hmt2JnT1aRrBe3IUMR//Unvct+uE8w4FKaq62
igjGYTvp5w8aN4jl8jXqG9BbOSrHB+/1vLLsngJ7m5qFhZ/u3aZKQ7wSnQKyXdMI
N5rRELmefwoyxuiifWaLAagpUVDEjL5OWuZicWInf0B4Cjsltyc5wi4n1OUo0e28
HxR9QpnVqJ8nhI/d54nuvwkkMqwyYyp9KUi2K4KAZugMBpUxDzkSdQJK6F/dRxKc
VCT5wnoeD2EKH9zLGA7Ms5DSgDsnPd8BHelRwEWomIvrfqGplPe5h3JTKqLhCnxY
iEl4UhiJYDRMcyBtLDt5xwM9V1xiuUirCNfyqeT3eH76CIdesOGZeNzVQrsjbGni
JTygUlr69NYZDNEqRqdcpWRq4fMwNkX3wlGGyUF71gd8Lxa7QpcAhceYq+BcoSM6
r2yxJsRpyBTTgGZYfiUR3dlTO3pBCztpyWzwcwi0eQ1vIKdlj/AdQAfcOC/cSU7c
pzjDPNyLlaS0xuFQHVF/NRf4KvsD5WiS8UPnjasYTsqbeNI9pCP8/Jk/MtuA5xjd
LE4/X66uLN/L8PLoHKkJFpzy/ssLaz/sXiPHDwIit2Q7NPsGnvNlBsl508lSuBi9
jpwJIysNjJ3j+48pR7DA8Uf//J6q4RGI5BvMBd8h+XXQQadQUVsuMjMvxKwW9Mxi
ZXomHUT/3bMIypjM8F+MDhv62BPIM/s/X8YC1H/lksvltXmdLReWILNSsH1HuSdR
HaYNRB9/WDTEsZfYCw+N/zKlAD8o64OQKasOw+KKYlcD9Kd2TKiib5lhQ8hPwiBh
cCaF0piheW26WWSFSEDdRYXgcH8aHS8Vlfo/eQsnm1s3lTOBg2RGn8p6fnSDfwqM
2Q8xT2filgm8crcQXGqXCDxGDpKk1DbYCX7XC/q0ienRZSQmUcg1d2ldRCjnH/yq
5VQz7L5SYFf8SeZRMh20ZLt8KfnKqGLWM4wK3wllO0QwG3cHJ43hG0EGSO4KBrJs
qJLl84K2gJuoiD8AbbdWJCNEx/SmF2BsO5IOFSOfV/WMM1nc6hXg8NqMTzmklb1f
dyvEYutvsT6FQAAXUXEaC4X73tq9p4m6z7MrvttI4j0aSl66D9+A5Pb+6LyOHTKQ
cPASKBGki/Xhsoty1Hx+Bin6P2tjnH2ZfHUq3w7pDddEsi/ALKKa339AWJUYx0+7
9nTAxlIKyGHUUv7ZQ8G1X0ud6F4vpiq6qnw8YXe9Ss5+YN53VOhLVRmG1Dr/P6HB
h+j+OJhrMP3lYxYKWtbi6Sz1N7hO3mf3tsoOgF0HnvhowB85174BwKVgyw6GHh9r
2oiKZcdz+He4mdLcNZmRVvtTcckm5FlJBM4sfHiGyis0Ji3/HtuCKDjG7gvB3E5I
pQ7MgfwrBVgWYov1NtXkCyZ47l8zxugR+Ek9xRJu8118XmWhRMmx+ZZtWKnyba/Z
JvOx/sa55QVlK/rICEgQSkjNBQFDLuRhaSwQ/QBAmA+ME4xUSctK+o5FhY9IiEr0
/sfftAxRgaCHxQTzF5Slh523BXkSyg6TtYpFRKI17e7JBynxXEC+vY6GS60ss6v4
lvAzl30viB+Rlv0vFnhjfkv8fO+yroyfaSJm02rivuuJV/HSojK0ImU9khppb1Rt
5v/NUGBa6IHsQIAbuDpqfA3sZJyMz7HnI86+Tr3Q0fWpboj8NGWyAjk521yZiKO2
UbHDwVx3cRu0N7q0b65lV/qHupeBFbycQSC7dK9Gf9MBbkXJUkK6lA6OxfMwQ44y
mgjbZ+65SRMUfzheiB3szTG95Y2YUKjpxlk3y3HeCU80/BisC5KnnrifD04U3mts
NcaGfuHTgrmV0N5IPsUmotTruEK0sxb0iZv5LsQnfy8bR7zi2FxQlgDHqS+V0517
N3xEG1EQnP5IB4GEqHr6dtIPwrljwo1Y2QysyEtxqFH+DbHOnvbe2QxUmjTp9xDt
islMmxyafnHOnXCAEfE1pe6JRuI6ses0MHXs9rUL42SfKvqIthSSBKKqin4D91y8
jKO4BVJ80TYEuHa1Yvsdn0uEUJwBYngx5OlDjHTse9NduVszbsbsqhGX3Y/5nnwp
7C3JzRd7yJxbCt3CZcfySJTfjCnBfRga9XxIwdEGN7fS6StZDcrA7m7OnI+NkXWW
5S5mJwWJ4MNPx7GWyTCAOFAjPuJ4ZJ8lk/cOwFV/g3cv3Jl/PY0NGzehMWGIkcI4
Q/zZsjAVy4G9J37ed0CWd4NypiQIjbNqpPSeVIMKZpFlvEWZnWXQwgIu36xalLiw
GNR6TMwjSJCNy2YQIdanTxwRODw358EyX48o2GLZihLuRMkXlVTpHharJMgc5N6r
IXZP/hY5WXMmzU5x0oV5vSgZKgg9OuU/fwliwFWi9ZKW6ZUJysl3AwQAmLXl4W6r
cbC4T/BT6CGwjVWXRE7bCPOYwXbHU9apQJWBUwagoIQeZRolpzDYJM8hWBgZjLDX
zWvAkPRZytz2TkyzgPLJ00FIvY3fey+LpjUio/6nBz0qgBsdjO+NWvBzt8667AIi
DkJK+UTF3bVh4PVaVaQ7kV5mzbaC18dlqMOlMPNd+vgSuX7XvO9yT+VmjAj/e53q
MYzY0SBWxT50cVilmxRZP0ECf+JLdiVvvFgFbu9JUSjDmJizTlHt7gQfEC+9m0B/
O5tP7QdbTdsXf9q1PsgcVVd7Sjwwu8egabRnykjh2pBxKLkzUMAaQVAdxFSBUZih
z4ktCed4OfnasGK0mP5lxYtMI2lJSOa5gUWsofBtzfYjqZbf5TNglDlamS0NC9rt
alRbKpSIdWk1l2+b2rSwBQNGnN62lzvXB0vDBiTyt3NeFne9LJZ6hyW/nPPfmg4x
JAJ2BmmP5fGHw4uUmmXSmfJsF2Jl5B7/I9AKlJNRSa9nUwLJrtyiCT5bsUTCLe3l
M8Kui7QzbtAPctoJl6TvqYUV0TdXYxyEjJZ1Y/Gjjnw6jmk32ijdFz+d2fMsNuBs
7Scdd8DHjweFiKJorPbC8m8zmuqy36HtfU9kDtJmJYCawas47rJ2eUlwlBCaaKmA
h9DFNw8GUjrBxOE6VyXCn6RufLBn/a66jaTmraAVXYtSTJ49H1i0erzQhqjzaQG3
rb9Z82PlU3fpxk8KJ4GYaszqlZ3MJGvlVnTMKkfjieKfbR33hSmrbcqKFQlmICIo
jG9D0AK8ePeT7YCEeZUHhmoOmDbzpixJK+jmFBw/OXDYjQfNZ/1LzHwKWnHqFL8x
KY9JMpJ2oFiFsIboQmT6a29/Ts6niB9qA6honaxQBOSzw93YwdjMXwFFCmzfGsaY
LCWZ2e6cPHRZ9mMdnHeiX/Epy/sVLjeg6vJ9rPi/SiBJf4bXr2gTQHMPFyLzrWy7
6qzMJNwLoEVNuwpdUiP3+8BHXykYqOQdTe18G5HCS0Hp5DO8as+qsSOX/ZCLBTW9
MtuLNssgYk5kBX4FQRohC/33/MVgzFY/KtPGMTXys+oj87DwJeOectxiWUf9LrAA
zRQbDiBSoX/oZpjdsS9lyWg6hNDzvh5gmZHXuJJNQbwlETLZw5UyQoA1ukH8D5i6
kJrAnzYDxo6LcHbSGkdQKfkbjFWuYFAgoHh+gMnvbj/xPQtoQLBtu8UtLe63liJg
mmRvy1iBoHOvdZMoGDFqTTqZ5ROS6sfSD7VPhS6eKXSvWgpUIzo3C7kJI3rFBtxY
67Xo9K6og9s19g6tt4NkXfzI3fut+JokbKXPkPr4l7M5BtssERB3wd9oVhVf7Hog
E6WeRJR3LS2a84JRiRngUzHcjYVLn6H3C34oVlVu+bVbkomAAmBX6A+1Q6l6QL2O
E8D7heIPB3/JNiIvbgSKa5jryHVpd5y9tUa7OqgtOrovExCpMO1i9+FW1xevmeVh
DA9HUmQ9wPaza1TI/+8wXhUY6vII+eZAG0vTsRFnYn5DuwWbPiQQ8OTnp4nVT92F
5QC8ao236vva/3+mxJJyPDNQOVMeuAOClrtq31EzhPANixWMf3vD8dSBl+UINHWY
eXT5zbq+rMUpN5U3/f7IXYrZKl14t2oKOAgrH4O60SP+43tSbHN6FUE3yyUelBgW
NhjRh4ykSYgyFJZu/5XTqFB0eKRJr3G08wWYTCW2KQkoIG8fXIZa949TzoIS/xYb
7e5HB/tNr/L8c3eDg68zlqD+Gn263YZFauGBIf2rTw2ZNJ0HiAZHOvuy0blDCLXh
FtgqlC1x9noaokNbUpqwxWcg244jCNZaQt0Ehjbhd0RrYWz3BZAi5O+D1JHP3Hzt
LKk95ECJcpZh3RrJYz4vhx/ormRPiimLP6pmvwtSrR711HoycLssuYn1Md7+XzCi
WR7diVT7novvXt72Crk1OcEe+ZKaqudyGxN8QibygGFg+dt/5hMb3ceib8F/B8o1
fGlSEZ7NSvN+VofKq6+PjC/E4A6JygYx+kcfCgkXU4psLD/Vbg7hw1c7W6CchcP3
XHQlsauOzsrbVL0vmfrEk1Bv9cjgg2X8wbrHYKaAMZsORHloxuArFWLuaLciGsbz
JcLmZcWivwJwwm71hwomDog0VPP0dLHRFYTCFp1MpkBHGYbSgTghj3IODbOaewDT
c8hMGrocCVmlZZbtOsL1CoThJVOpxqY0jvQOORdtBCWgmdxqFRk3JM5a3GarvQrL
FG5qju357/5UuJ9aWHISDETAcorY1QAezsnbw8+Yc+iBjysvezWsh4oTLnQiseHe
5byvzBXfXnWOq0MUG/BWJcMj4vQdhVSNRdKI+v7OXdARrIsNaKSNiby0pER5siM+
zQc7JHDZlxrCDj4Hp29K+XMDbL4Zm/j6B0e2AB6E5fiIz2DkVwMW3lLZXn5oRQe7
gkCq6Iv6D33CoBthAYQo0BoVabot4v/jTsvH3sSVWYktbrHRG1eOPkCwehYmfwcj
86PMdY4cF6jw5B6tzFH846Nmp4JZkguTvte7TaR92hl8YEcKVXl/2w3GV6uk0Ank
DrH8mL3ZbznPs9Lxc1B+eOjK2wd/tNJtbYo76QQPHpWmgzcvbfWravLAqPsyleAf
3GeK9Q93Oh3cUyBaKRjyTk7n8P73IEeOdbY/2dshZu5JNprAKDuQ7JI9wKt5hQr8
qjhyfSBIH/CkJvMThs9P1p7yYsnF3A/8+YtqNjIeCAJNwHugguhgx4Z9FJvk2FH5
uH2jB5uu/K5L0EcNbqM2FjchOXmISma6Wzc/WpvDdvTTctH9tXsO5c70+Zn2s42q
KvnkfAEwZgHeZS7Rv++KxnmFRXNkVw9g2M4T9qK2h1rJ9/OrRYX7Ph+/V4lg+/L/
rBJQgIOfUEoosZ2fP3UPzx6b9OVRvSzuuPZh0t8Ij+EHJndjU+Y73QzHdBx8AyfY
YRxLLPPRm/ZkeK7p2iQltFrge2kSkWnrf+Z4sRLOBvBj1NkAALNZ1Q0+BDv4HzcY
c/4AbZ0DZyFYraovWhQ7RGHleuIYlghGFHgqpw25vQS7VXdKTX1OW2AGKiikQp5b
0MdAfYvgVNyL9JGUD7G+UZBTWq8bejvDvGr5Nj2d9CInNefUlq8+RsNNo3ETbUuJ
qiajt9fMxrHjKLlz4C1Von0zhKIlMhI1XBz8vci2tTOeAux3gtPCPRcAb5yusjsD
2vSB0ft27AGAJvVjfIFLisvnqbP00fML603s3qfYanFzfT7XicztPIEEr+LqTzmu
bnMoBelJSE8RSaCKnzxCRclVnJo7VgZT+nKxLqBN9Gvtm1x7AUpu8GeIsRT0bJMW
N1FzMtnosxni4n2Iz7ndZd1bPRLe540aOJPttre6fu/yoovBg8elEffl46vXeZ9c
YN1dqrrhyhX8JMXeEdz9F2lXlxDFFCN7+/G0cJnhVHO/akzuwvpLjXtr/eGf45jl
glyCm0/l+kFT1oLr1dgX+x/J4+9WKEGPNdCW2uyCaDyxoQchJtO94pjAClkgxmly
VWbpEK1W+P2OQlU2WLw5antAtS8llRldOgTE0ASrjlwmTBImqWuUt8Y4lzt6Hply
F6aAnAfrwiPixd7za2cYTu7i0jLu5EBvkhxF7HQ0oMLHeT1BHN+VVHa8892O8Bvz
myKNdMf3UjAOVckf+9ug+SmaBwF6Xm2Ie8tMn52PTqQZ52DCltlDClP6HQ5zRBvE
EyR+U77S/IVj91d21kKHUXb5Qw7mHysf3CBZdnjVcbhw2/0kHa9Ve+HiWZbmAV4q
xmB3Lzh9/IgVFMulLwJEV4ifmvfZB/DOiTDWOswSpW0etlZOPtxA7S2xNAuzxwhd
NEftRR2OcXOVkNZozFBUSRsjHS9tpdcO7gy5RQeo1oSSomwsNwSyriotF3qyhxpB
JhCCBl4VHKDB+5WIPI7wRcyZCJdOYkN0QYOmVQPiCdB3RPW+ECjl1U4nWxNJea/m
jejExFBa0jVPwhrXUh3Hex1IlpBWSaxCL2vRUV2NbivleYDGO+lIYkxCGzxt4enh
UGQa2Hb+zFi+C4iw4LY7hXa4GX0LL1sKExrUJPidNCpCVWTAyySgtn1nPCwQaT1B
TM3N0bkfzk7xrORhhbwhth+l+qJRaeI4nV3JNEFNC86Y82+P83oJDH4jI3//QcCI
/DVjGtHSctWqGu24ze6UcUS6gbgXezwfc3+nBxcVOFVLiGfgsJgFdDfd919rdcHC
+Li9BR92H8a2Wx3WAorynRWcfoy4Q2o/bxd8XKOHasa5gww0WzPeTAIufo1CCNcc
ZXEa2JP9e50sG+48bOIgzWHOvnFjzYAOSrpXQ9AoOwdCRJcuu2wkyz2PCNTxmnmk
/adz9iEE04CR/LRtGZ5qow/ZOYqNTzymf2VgVogFQByP3x9VzM+7Jb+21soExtnN
p+mdvbk12xn2Zut9oIY74GXT8aYKm0jn7kzAhZENQk1ud3LRz/b/w+gJUQ/nqqXC
29HLb3RJTd3Wc1Xo/WHQs+9aH+KpwIPnb3SSIAmZo/NhHmxpEnlEf3sThDk2cKHz
h+R1F26L6JtUdnXogpyCyaLUCHJHDJkpEeuGx+ijbLL5PbgJ8qSSxdZVb2sOl0Xx
JrQsASlsL6bYeea0VK3/+5CgbnrdEcU1dtC/O1kaLtakp+kNbxOkhkn4kBfleEU5
jHIRJkt9CcIpzn4sMpKLr3tjfpBxb7TwHtwrsn1LFInjcch3fh4q7BNhCt5t40/0
OdjCZCMyDF29PhiPhx4vjaJ2ybIP0dkDaj4zQlifiFbz63KLcPQWp/wh3tU+4C0O
8Iqml/P1CTSphulOASCLLs9uCfoYxiu3HaM6SLOxG+20vEOFNNHlalyxIbwxAhcu
4Hnsn+SZlFwR/Um+nrWSdKeLPLVvttt8zQCKrfmSDQB0udZhtb2h8+tlDYLds/+G
cTY7eHEXvC3umtQMFxOdow0m1lEPXPHqENmac5hnXi5os9NzAtFoEp14KuDd41eu
BtvMY/VKTyktEvY4ayg4SdMNkQi8jQ+P+XoYBTb1uiP5Wwe9jdDeerIPd7SRm5Fi
WF9T4qXR6AvSg553GtBOQlI0kOxlBKFNUc0V8ILDRyqNoYKmm/3TF2hRHV21E6mh
nTrIITjgyegwb1ZP4jJeKHxF1sbzUDB/csTvOV4q1Be2yM2DPWTCdp/K+NiqrBJ+
qozb6gUWV+HB03LV7XRs0tmVJLdsyEmv+MlvUy0qQZDITPDAgdUybiRFKjxKJgUf
m7ew3HNy3DyNhy1e9hHHIz04hQqMPpwDn4R/I8BwgIb59j+5LArrrXJDl/N9nHqk
9pVRN4039vHDIM873mqHYN28Vt8l13QA2ehMb+lZHEz9u+BsBN1YHIK3iSTQTDPK
GBvFEVT3g/zmpNdrlKMv34cMv4B3nFY5rdRwzAvvBEaI0LJC/zU9R1m7mfFbDn8s
C1V3f9CLGkwdfDfOIYbce2woeaSFymCfVsINJTlhf7Lc5JTSEPuw8BkwGCoJw2Vv
NqKQpntrX2SpfxA2WNMJDmIKcevFypIXK0Bm6XTUOylsKG3boAAARl1WnIS4bFxJ
MDlmPH9VCr7+Veqxzd6BE2sPPw+mn/1CsA4sKYajOy/UbhDMPrU9glG3LLBTzN4x
wiLT6sJWrH2ycbu9jyY4rH9qlTczq6Ua5lYHSBI9IlgJfNlpdx5dtqaNssKCL4jW
Too7iXRg5MyFeltWV0gMDhrhN/TjkTqldxOHQNtefwGLPSUFkC2Ko3lHZxVVJDdX
OAthRCXKe6MtCRZCYbzWuSib2dXO8oty0RQfDJHtDKsw7VV32wOjfA8AeBsK5Bps
HZUwvS/fAgDVeXMMsJvDL9PqtgYGZae0laydr6e7DNkEhDH314WtXRZpRU5DBgSs
N61gnp15rLkAuKc7ZjsR3HlBHEFaO5x1xNPwRgL/DR12xbW4z++XWmBG1BNJN/8e
o1tu+pEnTryptXpBkdZf6L5Xo/asNhjKvjADaubPQBXeD+LjIVaE3klyLPOqWHJt
ckfsKURCeKCol7d2P4Q9DaVh5Msy/jg3FANioOuvNj5CEkP5MJ8EancpwM8nWfiw
9qN5GZ0j//OGinQOM+oPQO0R8v6OU1nduVAFh7Sg75iOAJZyVqyvQ6p39ZcvXf7d
rnXUueJ7Av17ZDnhzoz6rDn3Wy69Rz+7mQtmc1wYcD+13c/8mclYTF1N8cQeuF8S
TlGpCpGNtuj9p8LwV813qKby3ze5ppgR32BXGdmDzMGXO86l3FsLRkjNRnwQ2Aqq
jHofC9YbI18TW1faZeBNMcdHsvzxQEzgHZaoodMp0WxfpYxh+Q2ITEFyxN+QeoKH
Betxf38cbGY91fsakJGRg6AroUd0JA709cC+8PUM/2WTODc60Smq7psJm4TVqKCh
9z193ekEzcBLOSktrfc0micFtL/pBZbLX71UVTCplMp9ioysUF9LtcKTrnP1PlY0
WDAKrxjqnnppVtcTJLI78eSYabudjEUkvGs7n8x4ZeOhU5FeiTSvKNJ1WadzYZyS
8e64PdJQwxsN1GUTdAZVEbRSnt7ArkE3JCLKVwL5S/B43cOVkbSugYaSXmC/aqk0
b9/t3rscNIpMZB3akC90VmFU33DaLqFgDwkg6sVi4et3GTjZ11TOYQ5Tlp05DPep
/pmxdK0/Zn87CqHj2ps9Eu+SMhMUwgorQzewd5X3UiZXeBDRmZ/AzToe7IbXLQBA
whe1sTxiyNK4h0kUvmowKo1+T4XI5uceR5Ask3+dPldee8Wpw/V6PWO2tMEDMD0d
xgR+K+DB9FK/vjEpbrAiIJ08SuZwH2A1n31PqxP8nkSeSx2uzdw1FHVF64nilnIH
50JgHdRJcTfj/Eri7j1cY1R7LXHAv36krPMFbvHK2KQpsLyxi7Ry3p6nJqpoN76V
2pNDs+sY2VmkAdttP/4AVrPTOzPtHO2cUBm4S2HO1j21BIUuo7EjvDb/kHjk3eay
1LgWXd8pz/RAPmoJX/VnoUVZlAzX1XQadYST7w0UEEWdiWfFdWIWNCEhUTZSRlUQ
ahv0dOm1gcvzuR7g1MRqsl6/Tm4PXU5UQQca8P0EokluboQACxfJQE7zAk1K0zom
oKbsF5bLW+a2G/5Xd3hbbVVtgwg1czoZiMONwh8pFwLFdACVOOdCWnYgFb15JmdQ
09EPG3OHZx94c+g4R8LUim05L/6FPNRr7nH1/0hhS+R9MSz4JPJYtmjm2kVUHLVh
poi2W5qZIbq7gg1Alaq0GEQymPtzqy6mhzxRNwecJLwYW+9Ei9sTBRcfp261mCoI
CpFsldccM12TqNXTyu2bjZHyF2dCl5lOarIIgeSEq0RtKMqYYXDZzNPR9Ouf3NbV
3IwYExaG7PzAJ99ZRPc2cn3Hbf6fT17lvE/XaqrKA4ou26UqwykIfPsfi55nkqEO
6xZ0+3vxlVbMnisR0vljD2CyWcpXO6+DvOtnINZBZxKrYRSC/Vx/Cbf4yis38D7G
AmQCrEDls7S6WSCrzpP67xM5PnCRyyUQFiyDRR4/Xom/rkr5+AIHKC3uD+mVIey0
Pd5axYjni0pTt/mtK34G267h89a+9QCSRFb1ncjtOwMEMJX98aSmbkVBmuZC7ZMS
T6vwZK/5Vk7xoTilZjbs93rPdWD3IDgo64kpU+f9qlPsRIiBbfPyAXUatjMT7PUS
ucDVSbAuNS8a42wwzMjXDOc0/y/KnU5c4t/X4n3NiBQOg2PH1UnQJylKwmolwrIV
VSnCwtF5XQ7r27s8e/3TPTh5LhBLCdI2Uknxgs8BlOl7jf0UMxykGphjyIa7+nGw
Duh/B3Ipl3YxrzERAwV8TtaQmO4gra1d2YvU401sxqJVBCjjEizmcz0N4/36AyGj
/E12CbeOaqiG5QtO9XhGSr2a8er4bWni6o8hAXxh8b+E/vGfhJMUohsucb8gYzCX
c3Y56Uoc5uWUt3L4iIXf1qR2BDpS6XK8HdX6w6OHALEKNviG8bqYQoL2CjUNnLBi
+Mj2uHUMO1wv9hBm4URyMZP28wVkV2+GDaENmYB00FrK1rxYQHX7AZH2eBtCsvp4
er34tGsUDBUUKN2e/z4pgyb4hqtZox2I4KvfD1Gz9Z5BiwfHuduUS4kwoFK0DvJ/
Efu+bQohZfb5Li1I8lGQSSAFymycSfQvCqbbLKiVsllAOTXrdAJs0+VNtLWwKh1S
PnY7A/jgAuqwziZ/36Igp+49nMCGNsyS4xXscfHfZUV54yProCazAsTFjaJ+euGE
Ww/Gv/OGYwAjo8NLPRfIor8Fcu8VwhukfBrClDy2vdWRU391iC6Ou7uPjf3iZbUi
9FNElRgb/kufl2hGmtRArqGW8h+7u8Gxi4msw2mRKOJvt6QorMVP2cNTh7SMRBxU
l1H2zv2e9tHXV5R94jbscdsef++LFnAyM+F/cIy72JoHpelxTTo3Y60kZvUfradX
NNuhn1x7mvDGn5pmSShjxHbAI6GrRE34qvd5pwOUyy+Tr+G55YoeBnKQDVpe9jYA
7fnmMH3JZSx+w9QAw5RMXjRGKyUtdwvyw24frmd69c+VC0colyfFrul59BQVQavr
KCvDzH2B22r614Oay4DA/epKUHSIKT2rAlO5HGcHeOqqx7SbYLyrUYOB2DwwEicA
Zx4TOMtntzSGkiD71ISm21+qDd1TKT2rGK+XqrTbt6FlH+Cjxw7KwzZRpR1kxeG1
nraieI9jQdhfABpmOysJNy6hXM/gsSfXvWfJ9HgRlClU9UTuyZDmVEIfZKDO0nBm
TLJ8WohH3JzFQtyOnfL4dAT3aDPbmLVyX5FSwlpUZ/pk5NJ/1em0S9gQlPNU9lI3
C8BdaKNaH/m/MSnRshmNBLVqaTE1qDIw2xqw9gFKly9GTd+8m0Ap5j6gmnL9cn5j
5lpIArI98DPeFGZgZ6Y/DkB9lF0HHbee6PRMCGvY1WuvUwB8qPtuHF4mb+jbIzyX
SSGJTbuXxpPHsFWtqkxn+N/xcqruLhOj0gcJtSxQmQdTtHDsHFX6M6VobVtOFolE
ta5xUPTGYR2NPa0RYP3UVcQKLUUkre5dgjoL7o3B99s6XkPb0FS+85QC/FWZ8hoN
vNwzbp2Ije7wCopBd8N2uivZ6XprYsb38ivm+Kma6oACm4HM8/huAZzbv0lhnLHv
qG8ECp0vWv0ptC2ckHcEFM6k37ADLZtgVl/ya/a6NM35bQb8KFHNRBwV9vGZIm2y
0p4ns2hxxgG9K1XLUPEZ2iCI5mggQVBl9eVYQ1SPbvrgEH1gKTCBJKxSJdX9sL4F
7fKc7S7/1YOBhnKr6h+/duBpAxwyyegrvPVCxMZmoPXwwxaF88n/9TWg751WOnBx
Vbrj6ROESYPoB84mgV/GXhEflejJbDzPlc+BquOaTbWIgHILflkzaQ+3vgqr2Wx+
BYageswxGQ36PylW0LTGzGIBeZZWnttyiTkCMzun1fVx3HJOAyKewExTsibJaITe
YyCWwTvi9QADGLeeNVMnsFH5Tv+gST7cDriyVKLStxnW+XHBlfvyR3KZord2ZLBf
DNBEplUq0rxKXWE7E80iQdSPyu/l3rG8KDDMfzNJFT7EtY+18v5BAFp6ZTUJAXN1
td6Lf4O5uU2xpEc+ZyNGxWdt7FM9+9AgQWjjrVhAE1UemarKC8Se2KbLX9nIh9dP
e8WSJnB9OI8cjwLk7BFq1gabTV/LUMq53jpFCyGWxjOA/c1Bodk16JoPmFE4IurJ
zWYZzLBrYryL8i00zngHAN+qMIpYIRv4C1UkymFc9S/ltGy3vJMIhxAJT9fZrNQi
S+BGNStSKoH4DrkGuFLvuenE6EePF2qygdcDIqS1hWTqt4GIlSB3DvPDo1auitv0
e2tEH1Cgj9l5bVb2QOm7NWMs8vv1eInOG33q1ibqhieJJNva0lFiv6NMRv4UX6x2
/vGzm3FaE5dEBfDsaYzi7QsMnrzGR+axx+7BfZnt42Rsp9PuHVsmSvuVlMbIWxSL
qpVdapRrh6cQKZ2TBlOtY9vxyW2M1wjAEIdNkJf4Dy7kGWcOzD41a1sV8TqRxwbE
XuwBA9LIY8/TzjaReR5x76+Exldyy6hUyhUd+6a93wAL+32Ty1UKUBzZzjw+0bgo
CzVM+fBYOXvFL1JXgbUzckute5iho2b7qlcKDEIX6sJ+I6SgPX0B4GYQaJYnUPla
7fzGKoCr/7jXCnggQtLBuMgh0PD4KWnO+KhrKfxVBpDiTobxF6liHLR5DCmZbodL
14ILTCPFn1Q2i+N4IZm8cPZ12yNxMMV99xMcTbz2R3dFzfWUWJaEeoJEvVaMW+Db
NhGfozg6jZVSLtk2Lzfy0Zrl3fTkYGys0vCUYdeQ63ADvqBwFKwWpjWEA3ulgeSi
Dw5/BiVVmwrswgRvCW2gVCPX6yLphk4DZCLgZO2xJNg6xt6T/8ODwMb7jHyhQG8m
riaXS+MZUbjnV5GwN9BR+mDeL2UMUafaRp1jjnHFzA9e0xXiGOeeBv1TE3HQ3iYh
svWMEabz+ENaTRhZbMvR0NnTboPYjJ49ian1vAY/cUuM+r/vFK9WFqEQxdsH8WFS
onGTFau5f6NQZh8Z6AVe6v9JgMVH9uIP3IuOAnh+W4NDMgtVzNu01ACYKVE3FRgP
K8mWXjTEv6ZpuyUUl3YDC6gALhfBAn+rXeo3QwH/AAbtjA2TmmLdkHDw5xPYEmG8
oV6JpUgDijZsKEl0fZ+vqgutLONdUQB6RUZL4xnHE29PfuLg5HXC7o5ANmhsn6eF
xRq1GxQ7eB3Odi90K2wNEBCAk/bMDJVD06VVPwZdYXDckDYFA50Ut7X0AyCaHJVy
WNkOSmSh6KFz0dxWqEVIJf7LjZsTPyU/08tLO6e2O7bYSYXmmJMafsdmIvH5XxZ7
AgbT2ECRxqAmdFaI0RB2fjavJTXoDqwshyMJ6C7jynNV5p3VvRBlK0WWDtQUqZzs
auO8XDJhE4NrSN4uHIKTYOlt0dHA+uxneDII1zgfSbU7CRdxvVYnra1Au32h53Op
ycKRTEjjOs7uA2753SJopYnoLsEj+jYZNDUF3N5PRtYrdfMZQaL1hlrBQVbvl59I
F4OaWAbnmUBbWk+1FQz+HPFgT4a4K6Wbx2q4r+uXh7e7FozBGcjp3qJ3DxaU2F1p
9Q3qQJAY/yWrSIiwITiTdLsX8Lw259vo7lZ9val2grJNqkkD44M9JxyvOb2EmtmH
YAU5IBde8SKJITxgUtABjyY7n6z2I/MC1Xdf7ssWTCwd2L+fD3uqMLdaYozKKIvz
k7v+/T2BxB/FZcaGUJ/Ah0/WHUlQvFPj3EVYN8H5G5ydoR+B1hv8olwBLRoc4UNH
3zK3jUZs+ZQ5FVI/q9ls2o+FLOxpIwnyjX2gEgefDxbZ/VgGw7COOq7x0EILHNVx
EoZn+GK6bFmSpVXJtHxBdzlZ5FJRl9MDTq+OWoEuD+aUeqHq4Ms3RBwfTZQjwwld
VEgVWeELc6krpGJGUSZrDztgSglS1m00MTdQO9Uivl6iODrk/qb40CT3slWVJ4X+
bywyq74E0e7RNVR4Wb+lyqnOGRbWXy+Tx4C9fl77karseCscmItMkxERlF3JlHmi
0k7hG6liiVIjLayOLk67AFIwOOcl/OQApfmsWvO+O7i6i8SUnm8tWOtb4+v/Y8/U
uId8ADnSU0SgBvizYLP6StW50hadi35q5R+nmfWIeD7krbjqPKImacqVb966NX7V
G20nySLenoWpjXQAyBJhTqaFIda6FA40fPSx3/2KA6/0Qz4gbUsSn13U9dJGg6dJ
r6fTfHh6jHzUoo05heT9ChQGNTiDjYiIBQqi3/sh5WOs+Q3yTmmD07fl7gYkL2ZO
rlu20Fnp6Z0+LDffeK2E/u0Xflyfl739G8PBPeTuUxmOULsyUUSio6OdRahsa+2m
/SxLKgMetiV0c54ppvltESWeYomiYPRzx80uWU3eWTCVKgDr2hzPjjEZXvTi638P
qVViJeWEnMh5OfR9gnrZWbGjGAXZ//l+180T4ozXJnQKkcB8tKOr1/dRRsMzsLof
AaM46ylMuWH/PJp2HNql0nrDrVlQ1loorn1QUylYsC0BjeDU6xqqah2UKnqMlEMB
BjUxAo3rkQCYKA5MaddmQltPcUYkpgAvWkI5lmBMyTDWiHPTR1zLyel1R5sP/LWn
Kxb3EUPyujrpNt1juwmE3igt/MYLYwYdCD+TnNTq30WrYAXaLMgOqZ2wUM8Eb8i5
KooQwQAqYv4xw3xEvEYqT9mtrLm4T8I/qt5AeyoKWxIDJhTirHx35odhEeDK3unT
yjNRnNZp0c/n1DxScERxNrcMQcrzJZr5TRom+fgbB2IjKZTOWNnqqVfUDNdPeyyG
/KGeeWFDIJTect92e0GksvAKRCgGRnIjcQnXKdLQm4HNpP1KuwDEIkVMbmT1MAJz
vtSkY9+qs1WInjyW1hSGOntzCSF/MyxaxvC/X+8gy3SlBKIQXeim1V7MT6ETTgtA
QwnHp5IJxpUO/y/ODGYKy3RHdRcE90w22zxGHuhrLDj/Ru67zhvuagrLpjTkZBbm
BcFWbNdrl1PVIqedDdcsb+RYuWrh10Q32A6oC42NUgpyuGSdIgOu+GH8a877rSRR
5XIeFsYtkhZPsHh6X/QatyMe3kCAEC/j6nbqpkUiIYXocU4BxB2kojJI+EhGnL5K
ASWeCoZMzFfM4YN709ReNSFTK/71KYAUX6dL9ilEEiQGN/7QEl1phWT+SX8xHayY
LPWQDYeuGKcluGrFFwndIRHfT/tx4UIL/SXOr8V8pbcyfJmcQsebDl0RnA5W/Pzw
SdFovgELcCQdLrQp9wZ2taxitNnQuG1EyHjPb5dvvs5F0MB3IbZqZXy5LgUI1Vnj
NBQPrINffn0IBBnfmtPKPSSrP8rzETDYLzP4jnMcqW5mzMt9+eWskvyj4f+L4Gzq
i5/K7J66XQCa/HX0kgfGDgi9+MBCLzI3Spy64/5cnUd1vCBD5/kKFujVegCvfBDC
1i8NW0DwAQHsm9Z5cEe8ONZFJ0INd9Q2vHQ62tvDLFBgCPs+5dsxIbOUkGz7rPax
h4t9fON77EQUwEZpLIzv2WI2rv9Yey5u/0xaxX6vMbqaz8HWnv9e0Uk0JPPibXOF
bJfVTwJsOe2h0NkR2RVRQBwlFFL1Hj2fd61bzMr2+e82mo2bf0dfHH15d7t07Wbs
jiMAePn85WFEcFHo3CbYAzjLO3fK2Bbsas8IH5mC7Np8PJFYSET7DjPzMDwEw/te
xaIIUF2EIrQBLrz81/YBr1quEVSJl1gbeyNXuUtc6Y7wbhCP+kLA2VNQJJoyxQb2
oQIr6H7t3DBfvC+MVZZmIqItQWUqJfqs/5alWcTqsEq1TgCuo1MqzGL1PpSd/dBu
et4nSLGvcxLyCeMbc72zlr0c+8yhvYBMdla5VD9WolnOG8xfeLvaUqgr5qtxKWCw
DwaRK3FgoDVPnH75t1aykDJK1DMCmA5ghj9XHNVsKzItMQ5yDZEsl/Wy9Hqq1iqj
qF6tUVyTzcvCcICBPe2l7dT2nEVBk74wIwAbO9PhAw2vyRZ/1KHXTOjIhgiprnjw
YcR8+/kX7d9xqyoWSFxpDAumWEIeL3l8GXqhAlyEXfFuh0sY0DDv+oUk7+L0Q88F
E7t6tvNwJih7XYSiF2IjzTcEaFdmsjuIjZoRwTq8Mj5wQb4mIPKpj2bvLrMdA2vC
2QDt1t9DibGDuljk/mlq1rW4YKC0iAyCJhwZTrbpBLXnimoMzfwk07wyoz0HzAt4
NeIIdUEMXA5+e6D6JFRWFxL72idb02fSVelCo5w4sXfklMSDLlb43y5tI/Yizg+a
7hddgp73UG0d9g4szt3PUsBzwUl/ujVBgdtIc6NFT+10OdIqe0Cvk+OPYHIt3w2C
bAduk+sW4nYEu3JZRDJQQu3/iEyL0geOPI5XTT2s+htJMOTDSVMIhJlZIpcDKgl7
6vg8QIXG1i8y0yrS8gX915a/VBBRaD7r6jQSYc9BWVfhEUeGeeCUVXxQZzY4zo4q
6/O12s6JaCMcFKpN8NwiTM7J0aATDXRbT+Df8wHUplX8HscAFaE3jCc+02mM6vxD
W6C1po4cFCP5Q5F2S2N4xSAnpsQHOyJ+2T4+JT7mgZB46Q5HtzLTNYafK9JA3DEA
8/9sX3xrs+QGZRzZaO+Av3XYIGcha1Wfl2nekcBptUoWkJjkHx48SBz/4WrOi+BE
+g0ALjSdEmVNMLYiqdArEmbkcfYAFESVoK2We6p4zyWUO4FvrmKk1j2h9tqXuMsF
nijwXs72cueY6KUt4pFdWTtMVlOBpfVEGEbdkq+StUf/yoB6Yb0o6gPP0ynyJYWU
LbzUiRVQI5TrdZAeM6Sf7zZa6IOeDgN084B7R2EYW1OrVhdERuvkwDOWJZQauNZ4
mL7qPC38Z2CaLoMh96fLrxvk+cCQd0L+EFUeYwdqJQ6Z6KMj0jerp8its4lExTZY
U/pUWPfe5W1D7SnwZKysx/KpruokBLws2s4uR30W+AQXwFXo2b4rARbvEwJpmpWH
IV6VJXrRsJliz8tafCMHlA7C93uurEefQFdorF9zk14gRMDxfWzW0FTV+L7RYcxz
Wl5jrCj25CKjY7Ndm2e7cGkh7Dz5Z2ZfScti6durrHpv7lPorVaCPVIJfsLE7hW4
Xrs3Wq4Xp1joClFmen3ka4L6YBVLvjZ0yIfEi2hnMPwhmFgPr3gWJWIII6Ym7Zls
PVxT0fUzh8QyMButfYd7szPg/J28Alos8yvR8AMMbqSZEe/p1Y3uCNmUcQrNSRVR
gDfYpRQjv0DasSedTvJ3AC1Yz3e3okK42wpIxzp+Uk2OayizGxVESbpY6iQcMnWR
pX0yNQAZNgA3NL8CM6ajlNUEdu3+KJmlQ9danFu2MbUR6xWxtTooAlH8vbf36lqU
pvPOADQBg1pzI+mZfFEH5kzIkVY7WWHFq2lHUollmlRNTSvN8+BunQVdylwbbOD6
44dxnjRRYSGz457S3PuZkySOrTT5mCzWkGfEiX+gr9BbdZbndbGObv9IAhMzmNU/
Fk3BgQwd3/BAxaKzVyKkbVZfDbjgrEwbkm+SOPasRHSnAU2IB+HmHrdbmeFAQDKn
T9tTddti64ro982n3Iey5oFDinWK4gUYlvrXs05BdTTczkmbIP0gd5RwKkdCFZdc
awmnYxUYkHItWTGPYEanL9IpMGQiHNejOAD7ON3Cyx22xi8iUrDP7xEkiQcDks+L
OnWl/LexQ5FpcA7l5UFZKWDa4GIURvQ9v665CSc5JgG4/KhjEBNl7rVujGL/sdXI
2HQ3+Bq+oSlNvTFBB8x2gnNQuAjhz5CjrWhvNb/VRAb4fYmBIUk8LeL+e5AbnobY
wv7akg5pYjAKkbdhy1wdGegdJ9FYqsbb0R+UKJFxHnBCeXCt4u5D7ijFvDyqePxV
IU89Rl2093QWiJm1DZGK0QJYw/ajyqdfTdTVNR0F25ljkT/CnfSgIGkoDi7H5DZn
TKhK9vTJOzJnKdAQ+hCbXA0KWjUvLkmnvpNkMYOHuaD+XT0Kr9JqSs+y5MR/o73E
Eclq7PUGeKUMBWRLk7hJHAoUQ70YkrCjXraVKbMTtA0JBUQZcR12VIaNuP2r1nD8
MmaIbFGpXE4HslNOme4YJ0jDRtrXzf7XraJa94oXPgA5nD1QdYctfMl4q6aeMxHk
UNvINZKHfs/jLUxDhKuP5JmvrJH9bArQumnz6GOBC0BEVFtJbN1xq/6Xzq+wyuMl
3itEBVvslTQOKwqB5g5Yfj3CextU9R6jg11Kbo5Vl69e/rQMzW1T8bVvY+VTo9O+
VgXDg1Vq9Mr8NI+O8Yxuoxl06Zp9EEDVNNQK2aG6Ma9828JKtyM3dHHpATfIRhPj
g9eevjgJzjIrUoBuB5m0YjK0CDgcbAtAn88JI0Ep9z3ZZ6lIY/P2KB1khO/SBQC5
dqGz26RzMxe+NNKKsuPv80gNSsbsAdo62V/WWaq1wtQTZOgI7b7/mJ6DiWxHHAy8
VBGiU2pMlEq82MYXJN4/WVlfG5JcGRoCa/mTQU7BxrWJLpxTvRogsJrDoRgDk/4g
e8zvtuTKrtJJm1oVA009nGKcsPLXocapY3KpwvEc85EZwDlM8x3COz0EKeI+EEYW
7kuy3lS1dwaybVNYF8tA1/pSv7P3kJQJPp/Az38kLTuOJ1XY1vUtX5erzxivjB1j
D9F3Q4VQgAamloCt65/C+iSwzip9DfEZgSbUEcKbM12QekU7XgfOCeaZQSEpYl6U
5iAQp8ft3ZkJVksVsZmj2YKmUojqoOdML5Xvcwpi5Ab2oDetYcTmbbinWB+ajq5v
1+GacWC+9vS8OXP5vOlmlS/2lCBauuSeH4U2HPnYI32lRV3KDI9zmYU65q/jsSoG
9eiw1YGpWvf8MFv9///3DLSRDm2mBEUwJhOtfFrtjCfcXwO0Cq+XrLAPVEznGPb0
kW8+R9ljebFRE3W3vXi8R2abzOS/iyjNFdZTD5OgAGyH5FgK3V+mTlXnkilTt9KB
ZgbKUTZgO47Y2N9TCST1tHsaDXknVC1iPYfFqQmtC+xNSWocdxM/o0WBqOU9AHBL
p3QE/58PMvw5VHO79DYQxxHKcCUkR1ffll+I2PFpu3mDg5Is5lm43n06JEJathKw
L+Pz4CMozYL2xIjTvdw3T0fwpCRPGN6Xlprnv1tcS1Y51INLLDoZUZ7BkwK+A5/F
92bnHnjqzRK5E260cAB0v9Kx+RTSAm75NFfvCPPJM1ReVNdPulcEQ7Ed6VpDDk1w
DjxSbp3wsbp97bRNgXm+blTS55wzBJMQRurt0RuHU2Qsij3+fb8UaCX86LJ1RHCN
ACvuCXgU6Y32MqVwZRo/Ai7NsHtw0w3IMs7BYpli6XnEMqLq1lFptdykejhDwLlz
5nF9Er5vA6LWWerpvwyBPiIuK6lxcnmnpVCcJ568oQUgl3hYvAQU9kWwTuzUqxUB
XXfT1IK5eT9eJy07go96YDPJiYKZYonDEPFGCuDvPOIS21YcNOegQEwJB75Ecmhw
A7xZkG7VujT4E2k4ess1qdbzX+DDZiQ7tv/WHls8XrvlBvJUSpZ7+/47Nq7fUn1R
yGmzAHuUTcARj09wuNcBiF8dP2qJNmEdk1UpV66Y0C4rzWUNOnOqfbs6WOsNqNO1
ESXFqavx6ArikEFbxQG7XuGeGN4x1Cz6w7SS1PkuGZiKOWmTNi0oK3CV04KCv/GJ
r9B8HEongLsir8IJVDq7c2tA4XVuqL3Rwj0zIAh419vC+c8U4/iiiknLcjPMq94p
7naHIttjP2FTFxfuKgREA298qmHuAdUfzGWwgz4WK98VmF8FHOFByHpX6dG/ysNi
/r8kD1FDYBoyevCPNI9/JoY/Uy/gNc2FI+jn/HyubdFRzyGwU8uA31d6Mqs4lTf5
97CZpjMC3STjPWbdaSqH5Suih47OkimseCDimWlx55rY59+bUWpXptBmhzFc+0Et
AMhbq5k8MjBZ+fwdtgCRYVD4O/17qeroCCXnmBSiw0laR5YEFQhgE8pLh1eaQIRq
OYZKi1sO9pP1yYMzdedgurNckGsa8mH2uPA5ev2KGnba6vuqWluq/8HQxKJekDJ/
IzW3GJKzAVv+CSmLju4LqHwgeG/gJaQ0C6VVoYn5cEPDW5WLZkv6czhqHfp004Ce
YvP1KjUVGEmRtoma6535gjJitFBQN7gr2uz3+CLS5JNqxfPMQ6RIMcjwYiw2YIHd
O72ogZY/2vdgkzzp13UHE6J73XZRN2Q27Om+gEYYV+gfnM4IzQh9FZ13QGzQJo1G
KuwFNkmjezQ1AKA1tz/AYGJWcyrF74m28aPGwK7CdFOP21XuoIPlCeLZIfH1Wcwt
iE/ghQs5MH2hOkTgMdIX/+/gMVLbZapFmMAuyFtBn5V3M/xHnCWOVIXl5so4i2qP
SUemiXnXA1fIhJ1KzSXjDKLTRvBH3CsNvkjTHDX0aS2XCU8xYfT2I3RPQN5+Ky0G
VW2po8nXfY+a1K5qTHhUHRLZ3rbETnBqXkZuvof3cRc9lFetaxTliVQl/MGRlag6
jGiC0o0u5tshPnJC1IyJOb3momSa8QbpMt3T2MVQ5zi42ggm/lE+cH7vAN0ZG+Zk
qsM0HWiYbYRhgv23/M2ywCJX4qUhbyk4lIyCn1rRXiQXyaXKwP1MNtiDhewre7iX
sH0dIRUgLBXbKFHDbmozZ1xscL3P2KSpE/eFNX37RgQnkElqiCk1iGQKtkQ/TG4Y
bSV9iSF5LafFTSxciwuOYVGN0/06a1rUppGc1kQ0GrUbPGxULjPxdbqk+v7/XLjW
l+zIkPR2uL+pBOYnRLCSed4xsP1BEPy0hWEaNwWZdz6GH2HSbdr8zxPlbX7MUqEp
MUK7lV3r+mR0syJPPbXzLRzbnJUnr8lEkT1AoYsNPbiwRayhTRGlZhbbsQKYthUr
QNkAfwGtcMUBCEH6iBoN3WE619zpEAlECHZrc4QEqZ2I5aOo3ZtWiWI8CZ0OvyFD
Eb3GGjApi59VSNKpifINEYBxk85PCchYv0EBpxgzwUwAxmq4Lb/km0rA6Rt4GZm0
SnNZ/ebWZFpmgFEObF+H6BZDvrx+7P2wfRYxTpnuoZ7xMJ1/izOw9UKrKl8XlFHX
u8fvVJnPoMrMiq4GHihF1aOlXPDSz/d3QaYXJ1a/xVpz8q3YyzXT6OEObGmvQipJ
7wq28BxDfunJZ9ceyujOR1Co8+Q7meAueSyITHsmv4UrlQIIb4qaZl9ZHjLxgWEo
xoRLQRUnm3mgjYMw3aZv/YgVvyIg+T5VivqOsea5EFiLHiDe0OqcH7LmhqgnLiIM
HVO1D1+frhaEk8I0yJxnWLKA2AuSoAd1/rtiNzEPFXTGPk22jr41ReS5IlRpp+1k
4WY0+MwFtVacf005v3XWwfUFgZgFrUNflSyv2GZkCMKtxkGUWn0HTR2OPoWyr4en
Zy+/MbQTQNjJ5EnQ4Ooc/0WzYvifoz3rVd7RmcKHOgSDPondRp128NUs5mTIstCT
pdHeg07D5Z/oFVGykH7dnIBz6chIPLPcg7ahzn9Vw8y0h9ND7lvPhJ7gPBYg96zA
a18XHS7Z+bU80bbm3KDXGHtv1iBpJWU3AuLZyc9T7pe8CXi8HPYzOvo+qM2Kv4AG
oBDQfKFs/RAY4V8j0US2pRApk1ZBWBOn/4vWE8qrjdncgO1yA5SCE6nUqqySJkuw
Wzm+sCtlEawUHrVBlPkI0Z3gOMLZ6o9AIaIEZLtDGsij+tLfGhJMSsWbnCn80+/l
LbfeSihqzI+UUZgg6T+K8U/f85Dcoi1+U7i+PEuWK4r1IxXVjDeqhFc6O57ytDaA
dbge/p1usqcnmOHT/fUalxnKV4fnw3pBGV9lylW7eOo5UDOaApD1vjVadycDgH2T
DJfA3hJdDYSMus/bWQQrzzxb2rlgSCmsIE72TlGloQ0h95IdNSJVhtYeJZlY/snk
5qxBhu8BsB/bFUsz3rbEKe1jpNvR4JoeCbNLfJJDdx1HCdEl6CMIs4iNgcmqxkwI
o+2JX0oXWgGnGQcTT0dg+EndLDSCqSUgvkIeQY/k/E/VaZVpEHEggILNINte5pCK
0pdAGq6SDmkHyfCMyIC/pmyQskfulJp+JZrocgarX1lgu7i3+xKleoBqudD+trtf
+WqHZQXmqJ8uOZnYPE2cQ7IyIzRHcbpW/ofBlilrH3WtdDATiriyx0VFzcOfd4Ir
ZrjxugHc51Dna3bvPtWCMUHDuK7f18wEokULR1r8XOJSebd5qZC4Ae7qMwAQyiJS
i0iqYfErxuWInzeaSJ34MSW91cJ1MP8ug4MzOMgPIY06RTSXdG7Aw1Xe8o1XxrNp
OH1OK/FfuHsZFotXgHe9cGpJ/PLuJh10gCGYouFB29KbKAJq09WoAEwpBOoLAP8h
OGKt8X8A3ockEro8T+/VzvqFcM4lz3IcuSB9znGuLJQlBtek4BnX9hMMY3fABM8e
qeSIv0z8hmddvXAD1wxx4b5SmE9gvJnOFhqILMdFI5prq+25WGsYzhq7P87pdwo5
YXmSZfSZ0CKM0or2r/DaGmu9KrUPmd1jp1thn1KHV4/5Y9eCvZTtxPjkE3pBMEgl
53a4XYMWvlUnRAeXjH3ciUbaBoA7AB+xnUAZr+EwKSGNB1XrCQVyQaVoMuH9wwJm
M44l2omV/LupDoBj609RPzfBgoFMOIQN2Ca06scght4pXsoQGYBAVrDVxlt7oA1i
FVpdTMKbAV4K6cVr/c0GCgiHD5vXM6745nF5+8krNqsyWr6k9Vh6GOoOv52M8HjX
pGrYFGw1+Y1AWN/W3qAB9fmxzZ5aOwBNMi+jxJ1SqVc2MFi3VeqifRxHFdSGC46e
oe4Z14qzL9Gzh9TqVQStzIT9TWoYaVqO/9FwTQPAnB87zW7CTS45IhpFOfyAhtj6
AVLV4r4dAinB/7Fo/s6ByKP8XcLI936qT42ach1oKRpB9iGToBsx+182ahWEk/Bm
AYUcyPb2pnjU0hQL8qyE1WbkbkPmtvt8fbqR3755dhimhvmeH/SB5rUnLwCxNmO/
EoqRs6sB4Lhd1q3Yl8y9+WHKW539V2gNw3bvJXlNYsOdFk2Z6ef1XKF00/YTfzGr
iODvM4Rtv9Z8hQjJhOhYPVWXeyW0AAgFV8Bgdmnq1iHlJ/CLQz/d5uQWNUPfcDk8
2/yNYT2NgfESPbpQRYuxud7JSgJK+PaoBs8DTzWXWS0ovmaptw8qNZZidP0tnq0D
KTTaWIbjx6ZquJR6bhWOq4mA1NkDd+rcDZUYMLUQmQ1NEvFBLHnJSvAlAbLjJgTZ
AHs9fIx6tm6BRD0vAwx0gaKgeUnXkK3iTPIP0A5XEvcDmUOoB/g7AIIpmXHKzAH3
ggk+hgMPAC/XzIq5mtCxYrdVxZDFJzj+1LW1vanLq668Ha9bHP3XgxcK+jXhiPKC
QylW2dilALwIfwa5IuIcWzzWFidTBtXVrv3dUY8fAE8E36DlpPe6EtJc8AStb0Al
rfeE1/RR+l333JFiKcIGfNb11aLXb72tCKMPYAmey+8RauUvTgJzx9Tz1kjCnwzP
7W6ubParL6puJsWNkbnvcBxJ9P1TV3YdQ5bgvpcG0WtJ6YDYtdlkhF+PUtZyML/b
MUvsAMOoy9VvzG/XbqiE8GkodV5Xk7dGOee7ee6eeTtHkfWH3L52naUQteaZJmjH
xP3+3N758zsvAPWL5CigwdAeNT+qzjbiy5NUQlIBY9B6QrbcHjhoScvSGVjzsaMa
gO1d54+Mf6UbpkVB7mvuwty310QAreg5A+DGpu3NlbjEfxwnALX54I/eSVGKOfgR
XzibhKeHEpK0H2PrrQHBcWYl5xYbt8OQS5ZKvVFEY+NVNV0gcS3Yxiv7uix0cyTC
BHVRLInPtpyNfcmmH9Wdxf3EmYp+c2dpqqK+W3+k+//nSxCsH8xzNcHrYpffTHnW
KxWWEFWKi5g+JVRwU1RDeZeNLVKmdZSbHhSFT2RNXkPKzcoZPceqIWviuRUL9g2Q
K2VoRBpQssuBjVZtBPN5wCL5ak/sEtt30dfRqFfxf8aLt+NwFidqNDW5B7g3dxWu
8mxSR+azrQbsMGtnLeJWSoi95BBspTrkJrmUcShr4dZeISv8FhPsZsPh2HBVMRZd
LibxAyc21ZzEfnFmAuxv65+Wrfuf5vqAm1pkrlXYq+WJsDqOoVQMz0oyt4alczjH
d4EMFnZvx8Ew+0Tp5Z9lxyMT4tC+WNv+DFToc4w/hYrjMo9IzaDotrSztAzy1bmu
3YlutmDmpcDrz4sMuAOmSmjA7FeA4FOz3OjqPRyk3uKxbn+zVb89Igqee6tz6dHe
7camzen38NpJKjE6RPt0e7TTmzKZ1MwznjO+l2as00+oxJWXf8GpKmejYf6phcdS
MdNGwpHkmaa8nr2HtJjBfAtMkhTig7NYXOncJEBXy9qW2MF77jFrsKoDqIcJeYcV
DQemWfg7Nn3nfK1nXJaoB1lPOFhs0PoPfHpE6rqdLJahnLuUt9CNunixE/RkhyrQ
qPZK4/uOmsZ6FGgEy8jihTsFkABwufixKOJ1IIbTE+1NQEIIijhsZ3FtWiRxIOaH
MhpGBtf55oxDCerFvjyQAMyODqltuLNWH8PBGPhjm2zBnzTTNlUm63EDlINLlBTT
G+ve5St+XhEQsd2z7KdX8VjoTrjAVSB0+8J2kMKAnYKx8cZv0LgeCQJvYXR37SkY
3lDKIwP+eBV0OHztl/HFcnHezAkyv9T65Q1YOryDPoXURIt9YqWGKzvQr7/od/Cb
7ZCYWpZ9RnJ/+yWFUUNxFLvpIbvUeMG7lIP5Dx7Oiy5Z7qtm8EQvmzgiVYQgI3e1
j41k/jOjkp4j9Km1EZzK465OspxE/R2LKfoZ4Jk0Mhvi2/1RQyAz39GRkWW3Jgul
wZoIJQHV9q8I5hyg0DRufNMy6aC5o/3xO6t7zKY8IjiMpJHfGV3TCghU9J1ppkZI
XSQ9awyZpKLGyQea/4/kN4oF1I4yb8we9lTKHLT9Z6M616KjerA4/XGh30wuumF0
uPA4mxHDIgeZAV82dDsy+Fxdf80iShkfajvGbB9c1G4WbIJte6c/JxyueMY/UQtD
1lHy0KV6Mh+QHo2J0EWAfi27/ixyPCs04Bij4itC7TwU070fsBZKk2r1iPhvJy+/
CBgI2CXZeWQguUDQTjSSeMds+ftnh+i0mAXXkPJ79NMe5BeyzHM+vWxP1xyAi68Q
uLJcQ3nAqsO87qAqZDtQW0jsqxNS/6OKJIIJEYSZjL0k/OWKm3b4zEsD2OZzicC1
pCleL39HF5LHuRBgypc51jIlG20WK6v8nHPBxhIaP4Dx3K0NY6hi78KFhnABNw+J
ZykqcuUtDGo4mWfzAMaPLIv+kk32UNkuIgJtRqPz1WwnpeVsK4pDXvjf2Ed13VC5
1hEt6Z2PPrPc7bIFU2ThGPnJZjF1NJ3IFdSiwx/880M+BFcgE9Rq5guT0muDN+Vy
KZnrjVTerFgkNim5IQ81b2gNYwWl0FNs+rilWrev4zhrwBOMHjvRqWpCSkLKkCne
tB5qvj87tg4RjOi61IQt9PD/58n6gixEvIdpYA7cJ4UhdJoVwrUUJiI+TM/NBM96
JmY3d2lXf56ZY2QkpRFSKJCyJME1P8183veB9K4qiWHe8b17g854f26U5FziNol4
Okq/DF+mqvPO+MKaKL8PrtjzZgAst2op8WRJnA+Arls7JBe6Y172vcYZAA7+e1YN
/3W8t0K/B2lw/V4zve1PLDAzHPTRWunGCbhLbAF02137lWO6veAt5BsFDJtUVXEj
8HZIkcgr8MYkH6cx9h/DAi4cBTT8Uhh2NzVl+yIa5KDW6E0cA7zzUs2qby691L99
8JQYOU/Ijz3TDslyE0H0tvoXYs6pgtvhgFQZYSagRlynKiHiPAzxqg6eWqbCdUBL
Oh1NJlkHTWJXiOw5lZ1Ec2pfVBb99nme/Ij6MUCjBjFE6zrMzXtPuoiWuywS40QP
OlFqX8NiUYdH9T2CsfWtB+4RuieBQa5+qV89j6s/bPIIcyWo2cXkITmjO9wJv8ox
34tSAvNR7jjlLso9PORELp7hYXJt7Dmb4KhDyZGav7/lQre2AORoe43Tb9fhW1YN
uh3LEZunujW87/t4L6VnejfzIIHpkLCexUuA7V+Sg2BBNMxWVhwqoq5PnQ1+UKvs
o7fXyXB58rBBwjStKGsNQ/FM/sqEXAaAqC6ctGIjJhIeNhipCv3rEIXdOyl5iSv1
cK1ACSNlrAnmzOpnUbJ1CdeUAvvcIrGB0IswDBvpWhEogFes4/UM8a5kVE0on5Ks
zpxzUsVuFJ1gpClnIkay6w8oMUb031vNuesIlbOvd7Fm+l0C5ep1bdNKXPstEfdE
OYCOUhwZjrLxPRkGDarGCmoG60Z9midU3DueLGY7fK/n/j2tdX238VqjTgmKZXZ8
CkhyQefxCT9IyM69VnKhTyokShDbpDIX3xKPVBEn8eJLcdquX/10yIlyhUrsIPIJ
BSF7eTkMMdxElk0uWXME5o+th4GlMmnUj4jO9OTL/rjAm5ZZLux5/nn/NSIRX8z5
K7QbfzYSAh1k4TjVpP/LooVQ45YZ5QlFalm7ZF2HjfQDWupt3zgu+4UPal/I1qBK
eoxrDPOjz9bt1135+ItcQf64RjSupx6EFuKlEpAjk+33i/cylNEhdfHPCkSLYxAJ
O0QfO+mC2oH9dobUpbHoCC2alFjlpA+AgjcJ7cjjoqFi236409ZpEOlLaaRMBX5n
ELJQcCQwyle16WvHfTImj38NI4cN11//8zakM2Rr9+WxJPBoyfewcEKKdu37K7NW
4rFOa4iQlgoU0aZG02POgA2jEo2qPH8QypgTaIZtr05HWKA8REfsYmc7jbHwr1Mg
qpWiCtPWNR+7wQK7XiHSBcoxgv9X6yAqAW3mkUc/5As1WHn8gDpVQQt7CI48zdda
n+bSsiOHQAYSoGHmiwkDl0iHOeGDVxYnOugUwtBHJ39aYbGXCSivmOO2JhcPRmeD
JeLmIS3NpK6RYTHD76EuOQT4hT6+3PYHISf+tRNA4jKvqP3FcII3LieeX1+coPFf
Rmre1U/qlG9Mn8Yaa53frR54DudMNBKsEWlblHbkXqkLSZj0HwL7SzE7nQtJYQVy
5VodED/vVPR14VO3QEneULuAmfWJZNUB+rr+4jOT11BxM79Y9HYcOiBwODCeRxgg
xyZLOuJFU4E0tc3ZhJrJsfqCHqOlwTUehFf1Z9w+pSsQBlGwG/RnnguI8qU4dTjA
BT65mBjPYCFD39vyCqXGEl0gBfqGIeljfhrkpAdaR+lTyKhx/xD4tIGXskbu1Z7R
n71Wxm4qrCLE/V4Vk6qbzjjuZWXthalM/lbZVBnhj6nQTzlxbOKmw4CQRKh+jWaO
ZSs2fFi2yGp8rDtgPdtrO01SJRJxAXlQ2Hrtwlj+nMXfw2RDmYVPUBt3FCVaazCl
S9LuoDPP0xf6CbPd/MeOAs0sxS6FeNCPyRLO1UpB8rpij7gdPttZNFRh9UNxqnLd
EXwAyhzQeXGTJax5eeaKk9png7Tk+uFGYC2/uOZlqsw6OXjy56v8TlYWLER7+uVo
ZPbQmzymk/4Po8TD0pF62UbvECqFqKXt/EIvKrQIQSV2iG5GMFK2cPV6wVD+9s4N
FtHATmswNUSWcKAA40Lt4G9SbesPCnRy2PigS+KxLUG2h3YsO2PWgepR+2Kwokww
msU8VgAo+/1FoLAjQiOCIabNAhKFIW8WJ+JiYU5fQVMZUZti4DgV1SFSrx/RRFKg
IkBHWQ/zGyAp9V2GF7ms3aVYoiM3T53p5rsLmUVF8KZXgh974Zg7EJf9z5klYmCe
FurZb0RNgigklPFCa+AxbvDcETCjnGA0JUusfj1oB7X8pfkEJzIYwUtVOFbTvtEi
z3qmHeASo8D5J2GBL9hD29CvYbvQV/cuD5Q6i1Hl+1aJVLipc2hAgN2S/H3JfNoH
+ECiPSSZQ3tDQHfEhhBILIqfSJbhnS2J9lurlxGmJIFhoiNcJiz3Zk3cCKERUQt4
BNNPq8gosyAG6crMBTqpStCvYUCsCGPw07htdBu0ObL8lsZ/xdVvriDwUwoBDjst
BtisAam8REo6EoF6+suG5yHyUwuRhxBAhBcsyLQRXfS/MmDihdmOUuGhZ+d0fLKR
K5Gi4nqZ6qTFlpAt3Sw11Cf0sSYV24p8z2EkkyRqGwISz1Y5Q3q8ZKGKxhHcvhl/
CPjRBKCzpnpZJvSkHLxiHD+vnm8h4t5XIB6jbCvH/vURqNiQXXmXPAFWF/VfgEIC
i+mqAxAt3mj1Y+yo1m9oBi9+8ef9ywL7L3E2ualnmDKuGazXdaReNadv2mYwi3IN
RuN1V87NX0OdeyyCdxKIwsBGG9APelyxdV/BMEUAihtNH2EfiPDu+q+tmdcBf/w1
wuznH3exHFUGNt1O7Hf1zFUDR5gZPUMe+p3FEMiY4h5xqf9MstiIujJ2n71BZOHh
ELS9dU8yu4//AQD3nM6g33udzqx7s1uhSe0dxBcO3DT8z0mvJcVGnmuvkkoR5XXB
u6kul+98dumDAcb8QXLSKluJadMXXB6eEYbExu8plr/PgXR8m4kHnK1+b2ruOvxh
/Yf8tZiNgZ4rtUmQ5TcQCJx+bm1E8ul8gU32AHP9l13oCods/4kUBZRj1CKl8PW5
DVCYfuqDIAk7k9vHX5azLXPPLoEtpr+gG5LuKU5D7MIBBK0MOKXpKfPj2LLBmXH1
x0DZGEb3iPSgmQ6hsdeAymrUjrs2DYdkMKLRsPvAAfQM03wKqMdjQD3g7YabYZOY
eDGMENc/1hk8pW/rfCnDpjljFWedk8kMaHb2qZQMjRe6GewwapCeIGM0dQgrunJO
W9RVlKdVBFGua5y/hUORNdJln3hxv+EimbnrX0KrzGyJmIZX0TITw60rDiLZhf8p
/EfdTtWqhvWzq2aDMFsA99cEA7XjEcgwWmBVuuRbFBTyOEK82sg2isk7doKi5sOh
Pol5NAXNRKNUXNrGlaUq15p8iC0EXUbutBLyPoE7H34++zkrqCj4EVVpGRTsMGYY
TiNRJNZ8O4J+20n3ForY4Kbi40nbANOgiroX43wlmVbEu6nbufpdVEt1X081/OgA
0nHbJ2JuW1VQuskfJlqCAEHN6LkQYBjaZUgfOVtO1vmk4SRSbIvR1r5JKSgesBZi
aUj4ySzIyCynQk1qJ7gQwW0jDi5m4v501MY5iowJkQz9ovC4Rioro23DAYDPKq4f
VKaB3nS4cvLjIN9M++mkUPR3dvcdZpuRUOpJCIcAIKqa2MqMVLR4pdoNoDHOFvCI
D4nRaa1MolPc49tM0LXHlFa1Z4XUcLQZ3cdyk73d6S9n4q/dG/3U8HsQq7aNCieJ
f2fiI6bOdT/1hqOo7FkSdkVIr8dVsFDrfGqjRSfVZpn6yNJUJrPtdjp1js93O1hO
wqUyfJFoZqSfCXFEWw4kb07BeFbktkMe14iEOqNMUNd8ZivwsfgjJlI/oindiA6J
73Wd3GWXYS4LlIXoUSBJVO3SyOc0jFAVYMb1kqxPrDFz1ctK+cMoB6nZICavJaPI
04eeYI/ILGy48vIBM51YlboSe6Xu/NBaprZuEvo5eAeJELhMRR5D8UsQRpF4803C
TI1ssQj2TwHiP8iGU9Hwye5VCZbSnzrsJG74J7AGbIDc6j0FqMMw1zEjL6a5eahX
hsK/KbOs4oQiUuUmz7ylk/UmjRmC81Dec3Kx8VIqz25o7sVew8xWevI/4wkTKzLR
f6tMlGYIwUjEUQ6KmpSb6XX7td06uiKhfRcDCe+aUcZMpGNrF0v5X2+AmfMRbA35
jWpIbi76FJ/DwYImkKcpE7tEjTwhOCL3sSGJhMJRTmxj02cytjz1Z6YNnDw3F738
EfVpcEWNXF7t2aAWFUvWIXH0ueVtntoSe93KEk/wA2vc7qc+xMc+MgN64c0PmxzE
UrjfjVaKioMC6Wj9GaOEe/URgsg8ZWH8Er8StuxZ80KcOKBt0cG9DaB6m0JNtSU8
yMEiBylDAikGsSDja5CWt0ymaKnWcDkExeUPS+1PUyAeYX++c6QOsDTHv8nAGI3t
y4LS0neS7dPDZrreb3UwrqGm5dXL4WAmTvM3gxQ8aI/d3f08WnolctGkAKVJo4xO
SkEb5svHSQAhc6ndLY+cRrINJudYKwRLB2SgQErxkHdoa0AkFELe32mgCPzI3NM7
vNsSCBbbvlkJfoNMDLw6PI49TIb2UkK9kxEzimWTjM0xyjqEYPbZl/QnZsu+MTX5
J8I64Ezu+crJoyJHthqy0g5YqWQEFdEUKR2cCap3hiIi250xbkpvH4591r2+nI7R
gPfMDbp/BBtLZGZaynFs65XSillfx0KWv08EaRauugvuSC79ugsz16Xw6HsPFe7e
mqymi1kyPqg9iY3+8FIK4X7Jgz4l6EYAsbrXrSLV3iXuRe2yf5Mg+gdCn2xrEbeR
qKhfu0hExPUGLm8+AZCdEpxUNUsIA0FDEQaU7zCnbxrY1JlcVQVpZbROLa79Y7im
yb/BE8HSzKhgYrKOFFB24UUcYLRqyI3g2mdJDvN+GeMHjI6c1NHk8iVpAoWpnnMA
SGMge6rGXjTq0kbDta8yYzq+apRmzoLrYEtDx5uXzMuaVARWREAuoiJHe/qBuJ1X
G4FNfzSgV1azJ7DY3t9JinPhpysey9iG2VswzR/V3tFYeACl5AKVacJ2+6LqwUb4
6aKddD6PHQScNgXsm3PQpz1dU+Anq44MP61DVRljWgqVpHfs3qv1mQwIfi6YWg2b
wZcPHikgn9vz/DlFwknIextvfr1AzduiWDbFY4X7PRgVE2Xvg44nauxRjaqR9FNk
KYdfpnlHIxhb8K13iTW+9pnHGiOSHFxxLsgzmGDO2bQDz8SzpE57l84YoWVkYs4T
gkGin9FOls4fL+LJTfLlYNMQNa1tRsAD1ZD4SFHMmVJad74zZGt2Dv5LUQ/SQHHa
Y8cUSSeHl56tX0yqPmZ39pp9uLOX4YzwSdzIPRwsv4GxSxtMVyTqR4dkg8QWCHl6
yVyqD6XYlVbsrs9/hlzL/5Ru12KnClKHnjYu2/02Jbike/skq015gdxXbVvL4GPM
PqxOkW32Kzh0E1/oqlqLsZR61WkBh+gN6AbfoaEtTV4zpwCkWYEnjhPdcJTOPxrY
WgYd0sTvB+CpXar1IwGEuAFUStVansxZcg5+dxmFAf/BixYAslnS0c3a4tdp1Gkn
mIZATWc/jN1G0iW1nWVL6WAZz3TaWeLg/BkM3KdTn323j61OfkQlt6N9PtYRGHuj
ghg9+WBI27jYv0UVtpa+YU9B+kIAVhXdWEFRLECKEGSnsmhjdc9geqWYXXu6pk5A
r26mv1bo/NTb3oO8juXDfQouS9QdhCUd+JdhIgEQ76bfYhPnytz3n59XjIiImByo
3W71HhXaq01KMMqK6oZD6W3ivjTNTK0PvMzVC6xAi2Ba+m62w2KRczHoiuYGHOjP
qlxfLmETENRbtlYDXV8ASoGXOzbGSCORQDbIkgsEaRWsGiF4snWZWtn4i6zPO+on
8itgSMddok9t12rq04xkBLcWkJ7DTXindKAR11RQMfIvN1tO8IHIxwNiFEeMxjCh
BwInIj70gwWA8K+3ETWVxuiQz75RZuB8HU2XtpIeGqAjaXAJm1S1RBzFPUfbtp5t
xgSXMvanE6hl8sfN6JI83OAoXz3bp72DOy9NrgvfdBeNUQOXngVZUSlN6pmoFxMW
iMZIivCLwHovDNdwGmTGYxs4kyVt/XXlqapPA2UV5SiO7g6uPQOMdy/CEiR4Nqzd
GoHyN4ohi0BoK7e4Slz1itMy4kniCNo6RoDElX4xQVa7SS0bpoaf35TBPk5kNbNL
oUo4zi1p0s+yTVUSLxyUC1Jy0YXBdJ4ixezZvrY0Dv++v2Pqxxnjox/V4GQ5wgD9
hfFG2I+pxHdPb+KIN+qtEpR+TXbQrN2HGnnscpEXpl5mpqHmAatrQIY4tlhzRdyV
gNQynB2EPmXov2JkiGp2WT6kt6F1fRedA2ZNWrvMAJRCDyRCFeAa3y7RSRywtdC4
56XbyR8mdSYvGwKNpYYSgJv3HE3q8bucJUIIS/5Oz0mIO4mEWOXT4fkQ8z7rLfnf
z6RpfCMZSFEb/m+zau5KFC/iIlCh67jHR95u94vMaQeRUiPzkN16KgwNJnE8UGTq
TmrlhnkZCaRZbPB7Fa/GEWEeK3A2UXFoPi7HCRXR30NxMRhGPB0B3mB/FiwYVylZ
4wrsH8/DKAvXHEUlD11p+e1H/ixhBfzADhfC+S79f5RA/OQMM2UlPBGTDyfUwVqd
n/USW6Q6dKtmyynsLFaC7Nuh6UQ3JHq5aYz7CqGjkG2PRc6w1kBci16O4OGsx01w
U3bgi3fg8r0y0Ve1QZmgWiw9K04EA48hD7JOfipdqtZVtjrztJoBGNf6GfL0bZ6J
tlUzDQX3pU01lmwiZmv+QuJwqgX/8qCCD25Y/5DEy11yyyrqz5z5bM7zS4HjvmlI
DsgHnXxEWtY1ymNaVXCSHS3A5IKG2Bfjy3ZwX5Fe1SgKsjwfMMEFs9+uRjRP5WBC
iZcoOCo+JBzkbszKU1hR2KRJ9OZKuvNMTA+QVKT6DsDdjP2nIcTzBWtT1BxZNvol
P3GBguDpPsLUP6V6kuIxfZS5j1fZ+zh5eyFw7Nwldrbvdmagu0OyBpEyKEcFYAaP
Zk3wwpdBlkie7xXwRGcfuPv8Acg54YxS8NwFHlcincr38TdNS4/zbKvvYqIXA8tO
57jEJE+/PoaAEBSH7Dv92ZXcbMD3qXQmnj882UEantCpsY7GP94pT0fCr1AXPdUM
JWwMc2Vyr10u8oKW4uBFhYztwf4bX2+1IjR80f2bwN9U3QmhcgeRHtp2uUmyZv0x
GPpsfQsM7nJ/uOtj9PtChKD1uVe06CM2nWOOHvwMQJtXlv0fvZvM3JmeeFPfDpQz
LLHabGSRTgyXKROP+Z4vakZtwY1ffVbQhlWQfdLu5oViH5EayyJjSfZRkKYiitwo
5A5H3S1sJSOW4/YjZDW2YWrWFcZKIxkIR/FFJYzg92d+jvxPO387o8GHVcmOmeJT
qNbOFjnCSEsB31vAu3mggh/f/TsHQXv73pE29aTbQGb3+s6CyeVnXJ+xpa1K3ZqZ
UXoZJOKr9mOii19JVV7AjyKcef2sn+YJs9mH7Byi76AUoLVFp+GyU3Fu3V6NGLKD
wk3tXxxw79k7vqaDMj9qqQZnbHgTRuNUX8GxBi9sBZKOQu68z6/s2oRWQ0ql54B5
i8WlcJTR3yHkkyP8ZUQ0ARsHfgG2PHtWm08/rt5H1PgpoVYjs5dYEdDzsRsp0fqi
WtmKP7Io6kOlynPLIoKb21vKPRuT4pPETMZ9oYAFjS8QbMFby4EskPfNcnw99qFf
LA/gzPBUZ5T2AfQ8w5xobjyKG76IWNSF/bVc5phD0ETJSfzLuBEvh7hL2Zoa6vaQ
Lu6I1M1ODPjjlXqNZd9HdzGuImRXkLnKRG8gyEOWY+ZwFNnTA0YOisag9TVVF82o
A+T6BIxqasvkxyc6vd+dmaZRKW6lajD3xO1wLp8FpVAq7Cw/tGyy85JiGjcM9LCZ
Y36d3S4a53PrETWJ5Hl1AgRvGYiZ5+MYX0W29Fw2HId31P6w9f4aYYCQXyQYX67s
Zpo/hjeHDhDGiXtoYCQHF2x/UtngBXQOjMvZh4bvMzEQ5MdLscqj4aKrkaI4CZIr
IkUPQqM1HsrbwatDwzG9/qdpfkHsU8J86Mwl5oIcHON2nBtxwJPDQsrUN67zXEgJ
X6n6OABgPDl4yylOkh9HcHY9+XiQ3P60UCI138aYPKChqyKqs35X1tygMboGJS/P
3tPubVsdtLWCuj53ZaQv66USZTYQX76Y10WuPvQkpNCd/aEbezVlBorUQrk1Wrxl
ufas7o0rZ34ofnMbU/TPqTmXH81fGRnel42r7lYA6BvmxGp1kMeFBvzYeIT1IztY
PWYkW2pVvAuI4ZKqPXkuiN/jOCH7gaZfFvd3vLbok1EAL30EgPmqQscg+gs4Ns4g
jR24vIoX6Vp58A7q51yiP0ucAmDdmk7USvQxadDT+i5Cm2om9PRlViSjiZjMY60j
ameEJAzLS5jdxHw5U5pQsn1vkvfu32U3hv+CVvxpeQo3MDosD1jw4OdoaSWo1VVF
YRVoH3ufLTz2QpeK3GmW+xByM3u9AT4I0slgce9PaOh3e7TBHExkmGR4w+CMeWpM
uAC+r3MBoApViJ7MeDbuxfr1cFCmVTjDAOlBJLJw2rLdsmVQytJBo6sKktN9S8Kc
fLL+5u2kTCc3YWH+ZvRJmEPyto1V/pxiFfVrgVdIKXfPjIyvioPSiAMVhme3oB4P
90zktUHkwDLbN2Skn6RpRAv4BfpCoIYJZjctCKRFERrwk08aLD22lyda8YIlo4v6
AO+K1Yp+IAXFRUwwVN3u1fVB/M3aRnvYzq8zV+cCVozIo8WAc1TlT6YYqVPFHBFs
vqFcDoUWyCY28nLkf2chB/+8i1b4AFP+w7quONkzm3uPWxmb0F+NkoQz8INmIYCG
EaplTrsImUz0JX0L6V/am+tOlQIqmWoPdWiDncjKkbAIp4U1PSa+rrXCaETt6IWc
xCpJhbNfoXUhLqYFNqD5+cmttbOVB+yHMNMOoNIMZzTZMWwD6IuOXl1hiVtbFX/r
AKl3gKatz8SCZs2d4ERyuy1dUO7bHzcz12mG1pOZQjbBRYjdhMymYkb9QKz+Xi0q
1aJDslexlqZAa6Xei1hRsWBbLGpdFJidPcd93iD24JQqVQTK9fw76Q6ljT80J8DS
BinovhwFm+fm/Ds5gIDDm43B+G8gRZi4+cWshEyYVFHX+Q9hZ9eMMeIHymA58bZs
nwN6GaItXtkcGaq9HMSlla/kB+UXKLq8oSZUCnIJhOFoR58TLwfCP1Gnb16tFNMh
Xaknzi2FfkCgiF8daLwL9JCqlPf78YfbHVR1u5maeNvkJgf+ZMK5Am2bzwRkwrc4
7d7SPQy+efA737TgdPRzZuC5C+lDy80tK+Gq80bo7B9ok3YZUlanB6jPAlTmqG11
JDiaDwjBePdTYgJ4MnjCAJ49QAfIOeU45/vzVzl7BPcnfKHZ4ptuHi4Bcuqy0j9E
bLE9gXORdErlDt0PiCpNfbexzG8mivOEl7dIuumAaqSKtfXFmR/V0gXZbbCPgxTa
BBzgH1ZiAIAqCcCEyypK/Yrs8UcPgizHGKspKnaVhYuyfxH4YJyWhcXQbbiiKzEM
a8nFDBkvjd2ihPOcv2i1mwJIQse4Lf+XFInhtp89miDm9EUa+dl6VdKdkFjn2NPd
FR8ILNTfpzYEUDHlmN5tbRk96rpuNdgJfAYnR70+QUeyDmicRMWLugGpLzspv+se
KW/ZeWJTZlEIbjERisToi//hJ/FofLBeRYC1M357tr9zhxoV1kOspWy4PGMSVEQH
lwS0JkwwAaZ2uvWrJucS9HDYF+zx8u0mC1kI7VG99ggUWK2/9V4uVI1Kn6yq20aw
WUapHv5YU9ZGm07jwIALOJDcInT1fYCRjZpFlTT5tbZHPplFlmotLozJRgyzZVG3
pvseHaVFmMzFs16/tWzLOUgi4asiB0E5L0k8HNzxvgwGgi6mPb9zhtXHFCjXLxbj
lbmICxHDnNNdxNI3e1vxAakMqYDUtl207ZWZByF2egMPyrsqDfndONTCXPji3ZMU
jE+KzB6uufYmWOgI/dfcT/xFvRlerYPU94zNFdbcK1DnW4MrgugUFtILvjL76/IC
Xt38uGQQ+L7hGEbK3TI7XUxnu4V8iSdiKmV1bt42Fsn2b8OWg5wORfrUm+5YqZ7f
3pbDrZAOm6Zxj0q9LYRyQQYkVcgdkdN+LQm5RW/qvbmDb8SSCci1qDjV93+D7j1p
TrL6q4bUVLfT3NQAknlnFAYeuAzcOF2xTwoOvdyBTJvCAJPXPEZx7mkice2ZcH7P
hXS8EjK+lGrHmVPd7Bxa6cyoOf9oBI/edEwKa9D4y2R5k+ofurpvOQAhPP6yJc0v
lBBF0tC5VcEgk8rzVFk/9RR8bwcoEKjnzOQJdv29xKQORWroXXvZik666LXdHmq7
wuJin2fELiSjthiDymnIuIppCEmtGH2ZbbxLH4ik5CVQ6MM61brNgiubB4nhrZ9D
16TPwoupd9mOMzAuR0/O5UXOb+2KWloc1zU4MlgViCsjyCnfptNWAldhJnZuTXIR
4bvIktlkH2mQolN056bMGev65Gqg+bOO0ZvoKwpQ9yPZLvQLGI8SE0ybO1ESPFgL
t8DQ2D2hQqMimffNz5AGegBuh6Y4p4jzOcn9F924Oa+jxRHmg+IkaTC1Sn/ep5o4
/g1UYRQC3yS+AENQaA/t6ctrFudnn5zPbm0cYo1DUxda64+AXFzSf1ez/NgW2ao9
L86c+mLJqX6Q6gkQY88PHj7JLU2+q3dVSfM0Eh51SsCCnQ9c3dIVVfEelckxHpLq
OuOFUw7Y+u9RXFh2D/Sxj8dAu3xK3XL2SxOKmWZcJQCeqN8OWtMzjBQ4zbVntR3G
mxqT7C3nQNaRSNTt5kNcOS6L1JT70YZcz9O32kSifZIYkpLVA3Pgdv2Cw703RgMK
8/Ebhw1fGN0T6poBUj8y058zV8ae+YTgKbQrJbDtxVLij33YY1RDADK+FEVjy0cb
rnrPr+wWOG5vgCNgOaQr/ZQTFQSyxlTHW7L0P0RW92kinjE4UuganE4cbVcSyHug
sEsuufR/40r0t6WTQdWiW32IGLZZBj0H/6kgVOcIqvevEuzhAClRVno3YpoU51SG
oh0ll1A0yhn3T48VeoMF6TzyzowzJWXHjhPY0bxxWQkdB16ZVJ9yncPVr/BkSzEs
mmcHL9Ait+oW8EVEhoFjRoI25Mp90t6FKTyVIgSbrGnkasLaDCM/oQEqqbuXoysC
lK2vw6StpOGSNqZkI+xbjCIK2U8/jMaUwHM7ifyhHhagxOJaO7zVBjFr9d9R3DPZ
2wkOKcuv2L0yY84wAA3aCeVnl+RZS7tVEBIaE2p/zVqM9hb+MdXlzabFYXIClGXb
LDKoha68UiB+Atwvhq+zq2TpQY/DMmJJYt+kzO7jH+tV1Wlh6eyKA5c2/mJRDe3T
iArOqFdjeKFeUmTMvcSD9bxdVayOz/R0BAQ0PIDoLhYUZq+LuYSqyav4fHeuwvgj
47a2KwCVQ5pHoaiVdnr+daCgSWFCbiy4TjHgTLxEC8VbXB5hx47gjorzxmQa84SL
7dTG1lZHdqki7F9KjRboFmRiMUyNtP9NNWMGeWAfscSSnS0CTImGc1ZtPyZm1NrM
S6WTi9sQ8xiSuStfrim6M3NeAFDSqV1d5lXYlSBYppJCWSBVsBy0vK/blqpqIB3Q
OI6ez4P4i4NvBqUjDbePAmweydAyrRHpskOENYjLCnXNn+/3hlOGT3OhsjlmhCKS
JvD8To/0tD+xMAczEnmEJveNL7+n44aNfUwUFyFTMayifLcbNk3e34G8iOWuUd6q
rs/mq6QSEQdO22aFOYoRbK1343Udug0vMb9MuIFDJ2EnfcWTOzTUrosVkyewo/Ie
f2QlhrG+xkIdB4X9CO0NRPD7V5smIhGXyu88TYEIBtKydhg92JQGHdmcrWEjTYl7
tb/gRQyoZxm7c/jkU5p0BYka50BHJsFoXg1OK4b7n5zo++6IX12+xRvxzACY8hRa
PGlsAm15Js3S2sxRNgGJAGK5CD8etsieWl3+zPUuMrULE9xMGJXI1t0pwYftD/pe
H9H8lwZ/4YSAH7tqsDXegqHWLEyxBPRKWqCUsJRnlWbxlw4LvwABYwCM9y34kLwv
z5PJeudUAU0qAVnjCTcsed4V+DYgzmZGXcngfVcHtEzTjIJrp8JFdjvUfaq+F5P/
/Dho9tnM2ip7kcg/kBuUbKHNctHmDJgPjHL8UF+dDhYtz3ii23J+yL9532IwcO5P
1gPQT/zZB1TGTAXKihU4urCd7pkW1L+WbckGFkkuTivDszCKWO3UC1+WF4hTdDsl
9D9O9MK4jorukt3kEy8xBFPjZGCMk/CXqHx98O/ziajrIumSrIcmlNjrlo1fsl+b
ZZycAcizoGWfQYjQUkhX0a2QPx4TN3nIIRyQXnDcILhsP+HkCT0R+qWg8qgJ4EHT
N1DnS4fIC1bf2FT4hCbVsQ6vZgWt5RfoIdJuVGMHqBOPkbKlyqWbxxb4rUZN9lm2
CqAEgC0E7AyUh8cRUyGPYJfuQJTRn1oXodYpLh7c14+lYg8zgaLjy/GU770CqIMu
R8mZ91m3uQLKTZtwy5CmxzUnVkbDgqdEs7tAkL7Fo+STTkZ+ZR9KMuYvY3NR3cad
CPOtTsAGnV3DEXVpbN+gw28OwmjhAwyYt/kpmA1fGSYJZ/t1LaXr3SdqgsqPlV7t
9XmhOMaxsL/eoQDfUgrAhWRMoLK7QRjJHLycTQ1gcJcD+MHABPPLOQzDQOrZVHdy
XUFoh1yT16uKa5Yx3/QKcqI7/yfTzHol35d08vDWysqAmuEeYIp5JRCDcuCAaQLn
j/Jqgcs9/2TQyJPX3hLd2eSj0PxL6s2G7ZkqGzAh7UzuygWB8jG8avAyJmnTdJU3
brpAbZ89MbeCgEW36DynlFUnjX0sg84QpmV4AepyH7f+VZRAeJCafzMRdpSviK/I
myhR3JxJceT1xbc3XaXR4Ip7e2yD72KrU24MBqwIYPXqOMoCKuXDaVA0FaWfCWIE
Kcf5aUClYZT6zrzdMQhBc/uhFoGsvaJ3V4E2jsOtWw+UH5vY0qU29Ay3wBQg4sna
vZjkgbRGVT1VDJN9E1OcmPmRnYoClOIn4FfK8YK4TDprU9lR2stIl6p2m+45ooEU
CN/yCirzVQlGACdS4ZZU10/iunVeRaaUNM39fFC2J84IbA04t17gVYIANA03aJTI
VtgfAqzTyb3OTALHVprsrGN4OI766mgsYPSzU6fMNJqKTiFYlpCiwKV5YDS2P202
2qkOd0m5lGDgXQ/Ty26drcYcxTWk25PEfC4dJgt/+Hazn6qMzNRwmGCdgtuRKbdP
4CEfK67Fe4an6rxkdrVxafyQnoBsrATD6xDI+jrm9tajtVXas/d76o1Jq6/A0ZJ0
+Y6LZbpv5fnd75XZhYjQyk+IfPDK2CDBNHPgC70fNr+1hBn0s/nnBFrM/a0J58K8
88miGeuLHHJ/a8YpMtBR0a7UpV7aoS9MRyZykOyDpFAB2X3O57eIZWUNQxdL10h1
PNRNVFqsmMTbMoW8KSWn9w08UlRT6lm6uxQIMbL0a0Q+ViAOFZF3VAGmEza3P22f
xSK+h0SHGzaqGbGTodqBw0SG7vG1t8GSOELJ9grCJvIAH08GEroNLKLetbJFS7kH
obhvcXoLIsep0W/rwBKuVWtIGsj/Mm5htUSAcSbl8l0b28QHL2lu30BoRzccehAm
X3qhfieoovb4Oz1czv9Y4ku/zZ4AfRbAj8qOCyN1+sKvK+x7OaO0ycKzWSQXsQkP
Ujtume1qUZRLcKYRNqKdIv148HHhOYbw3Uh2sY9Eka3P7MAvFbGBHxm8QSdgjuvp
XTp2QZ/1euPEGL2GQZxVz+xrBSEZNrMY/c5AxunhcZXOLmnrLQFsJC3K7IBLf+Bo
x/F8+N4bePD2xaVY3lrhLqVnEw7r/unYCQcHO2CGztH5vLeoayIs4LTH5dcRs77S
Fk13L9i7g/UxSz6W+EI/AunvVeYEEb7xnJnD+nmwaSm510akg7s8OFrN7cOQzLb/
AbrGK9zL6u6XU0e2rUGE2SD6JRe8SjZ/clu0Bz6QwGqroAQpZ1egAT3FJTR6JmGN
rTuuij2iE+UN3X7GiaYXxilXTwXc0cVC1g42qvHoDJ6OQVUXpaajfJ873khnYVr8
oPGFuvMnQ72m0hNGwLWFe6cc8brY6c6U4DYey5jd6YniT9arAlcEiEmgZraAnbrj
WG97gvotR0KvWJlcYkOt8en4fUz/7TrSvy5QoC/lfe9DlULRwO+ZgoRPmTExW9WC
I3ZNPMU8DtE8BruALz4npeagH7/W7tg82wxUFPcb/9ZT7Xgn5iXeE6k9a9kTTkyj
yBzJwP/GAsyUind/f00m1BL3+R82TJl/paEXKO87qe0sewvhxldeuoCshG8EsQDx
npU0BBUx44jEg3d39+EMFwZRy0mbzvbJZtnx3pTYFAIADgZQ4hI93oEtXk3ev5WY
FQHOVIoEVLdw1qO+2nHK4e4TLIuienup7kcoko4HmXPgmJBj7eUhK6p5V8TRcLtw
NJsgbgN+mbzL1wcwK4OpZ8wbJ8nMvPcsBSOKbwcvU3okes0nkQVpMtlsONZJj14Y
R8MR9IkywB/FeNQRgi/OtLq7IxQ6UxrjCoca1RfnSDvTcejeleQD+I6bf5U63/JC
3wlhZuDx9rDMGdQc1m7BcEr1FZ/PKeyw84OIuDJZQGPfQAD1gDV+926BSh6AYnTJ
EwjMs8mH/C24roivDj9T/oHPy+4WrxOzj9h2Nk634PeE8G28p4fDSU0XyRZphGLt
uLqYGMZgVIMjWOIDQ2eZUQ/JKXPOz6ZiTPu+xqSufu6fdU82qk5XGzESYemSflFb
k0cDZft1uqcm4TyerFXFXMfLXd5s851oulu52ySCDScyCAeP2TtFv7S6HiiCFkNR
I9pK8zCm6DFqHIo2vq21dxBm9fJKGau4Y7NHiw1Qty22j2kzMmurB5B7vTvEXj06
DoaceFZofMXcOfbh85H1dBfgYhl5S/zI8w+0cDj2mzpcF0u3ZpP4U5k2brx+77ZP
AQZA0BDXoPlq2Ml3a5HfoWtDKtKkkZLkJ0Pf9XNYvUu3VKcxKiNyOornwDPGSXn0
J7TYm6u/ZJncqLaD9WIAtIfm4kSpPa5CQK1AXTBXebDkXYUx8EamV8Bxy9EGkN1Y
MiuWSpJsuV5thmH/kcGKWu1utbRYjSyRIcqPjih+W9HEueFhHRMqYkxhKp3SE7iH
8XXsMQA/Dk2Rcv1xPZd304uw+mDVKpAIjnHv0Kp5V7z607NjUIERi600ei7H94ad
+Hz8OUbzkokE47tu0CFPFDV1e5kGsNydbAc0coR9BmX9XVd6l//rPUKvjB0wCWHi
3QsmtNgH6DwyYdHL2IxD9br2qMXOQoG8O63DjyLXnI34xHaaUucA9/Va+FYJNFHJ
4ykzjFzgrIVciWdmFRXAtrBJ1ElukyZ710gt6fDzDUWKyg+u2f/GtA2ZQltKIGUD
EYVaCXUWUNoYiOsaehzn2bmeaTiIcGHXh3P+yVUJwbNPAmlTvBZM0fx4kYs1fUA7
wc6AVWCBlD1njZdV6n+kuV/BPq4ecJCV+hm9ayR0vNkxvx/0ULqNlu8PUGDWuLwF
YC/WzL9YHx3nIlIZYv2KpxEFFG+WTHJVZs8h+DTc7y/U5YVlqIcCo5MWrGTOduno
JqDIoNsvWlfrT6Or9/riJ1zg3JFBYHqMmFeKwHKm0FUkJWaZ1PnnP78G3MvLKgJ/
+dEvPTKr+NKnDOE8+WPYaaTpNhfEBC5NAGD4SgaXJQXx7A5gXNJPAmYSceZYD7Wq
K20ZivmpR6D6Df7JLjDBXHXF2beZbB4tI7dj4Afr9xLlGOBLdKhADbw9QFx/28u/
IBCxpnyJAtn9R2j2+Bv3lRABghM+JpLSeunRa5eCP/3aVkBsCWW+tykP3YqkO00S
cKRHaQBQ3EUxeU9rECQFSIdiW7etff1e922nJvohujjZJIfai6gi6gavwmti9Gn7
cSvJn9bEv6u6GfXpraddl+aEjomeT6hmGKCSQRNrRqA+skzRB+KHwQV61a5kStli
WWio03GS768LQqvuH+K/EcIMkHseLvapK5rn6se5zWMkuR3fRmRGjbYzxkz3UlHL
7ql1YKKtKx71YsvX3R4MAYlEFaNoyeuRgbOmRh2nTylC9wn9ECMeJlw00yTJR9Bv
sQReZH1BtNTl84fGvK5nJ9B7khh2L/Zs9U7PUU1FPh3HNNjn/2nTqiXErbGmFeIB
5tWIPMnhSG1DoWvM7szfimyJ3YMJDPJE5ZzQBXlJbHtmAvRVoXQDDurmbE/hNKSs
hRAYjOSVkj4erNNpVo8KdvrrVOh25k1umbxchrP9v99Nm3YeK57q2IvCvSGuGk+9
B7klO712/5WNWxtXS8Tr1nQ7vjYCgcPqhB9smrjahRAzqJ4koVJ0rAPEF7U2jF5o
xJ9FyXj59372jkKEjZv4H4MqkBq8lei4U/anX2n17EDqYZV0wuJhbiK6tXcljC13
QzABRlK8VXo6RFTLTHjoygX5C61VfDcjmfbQdliv1STx4W5DP1xD2opWvU0Co2Cr
v8ZFfgY8tMNkPZT38A4+z81Dx2ZhO/IWs7TVZEt5SoCwRO3Vs0ZOrrw1HgoIqi/j
hdE9PPFH7a4MGJdSSEEa/hReJMirEY9MMqjehqNvuvLqoNzvjkw3Eb88ToU2hf/e
R3iI3bsniWmThOvuSftunW2wPn4WtVco7C9CbVsHGynfS0Y1frYkx8Rlj9lqbThq
xrXxzKBzo0J1hTjejIqJmiBbCZDRu0TaX551iEZlHzistbDrRipedtO3PvqmKNth
DcQthqAh6rmhlbpZF7w0P7YtpFJ/8odRcaGHW5rjDkgXhQxKdTMwT+pmR46nDZKF
4m8WSjr8nSeHABWR9pCZCgsr14uVxrvHumROv+LguM5nVwwjvJidyGi6eFSre+7j
pQ9ExpyDo+Ne9DM0DfBL9Js+/iI6skKNWrjs3684wDsLHLNMS9mj00CYybw5s+Pl
KFd2YKoQiH6hlynjJXaixxlXvndxho9TYtxjRrhI4RqLB7fZTtZyk+S0pAU7Mum5
743oG2Sui32SZ96gZk/5dY/VPtyN3Erc4OJ4PIkNuY4faJBFpgxJm3qgUE5xEE88
lpSudWIZ8v/mvVeVPkieCynZONnlEm+EiN4FRF9rAReP+TAE6mhC8C2/V1ufw7Wk
5els+k8ZGQ9GFSN2ruiXUtKVtDqQFLoZCW6kUD/azC4FKXrOoVCen9V3juP0o/+T
c7YciRYLYmmutUVfShF6X4kxYUZ9v4EGEqX2DEGZKsTHBP6Rrk7BTvqk1ErWwpWR
r98W7937U6NQqZl5YAQsNPWTbSo6EX8uPbpZXcAJ8aE9Mzexo1WEFe/7MYIlFTvi
yctaE/M6R4aAwHY0i1BL8YtR0pOIjPaiNtlpjahrHFRANzLpw+OFqa86mpGYlXMa
PaxBi5czNMptNQY8iyGU5mnicK7adh/NHpgHwWfe4Tsn91NUmN4fA9k/Vsr2u1ff
1GLsj7SZ0saqj6eADIwhQtzpntLUZVN2PIdsL2XqRGq5CRNi/LEGuXxtcWYGu+0X
urqMGsWDM2mpvTg6iDpX6PfBeM5eQHXFdePythXkxzNgxJuEs6dsfz0CBRZFjvBv
4fBKvQdOJ1vy3sIE4SG/7Ox6UhgxaEpRM3Mjo0awQXkEsKPi/ABXDBlbKWzFd5bm
pTFb2J17+CbGylt4RNEYdf7oziQut961V8tV/Parql2ieA4Qqb/sj5gFULnYVsIB
2GtLGMXPwmDNI3YfiKQUzGRB68oSTw5TAWSQtyFFb4NOotHEng1MMl7/HckxXl+K
nwCQJFnoWp4oIA9VumpSMvlD9A135/7b3HGLAb8RgMtiNqjTUeBJpt8hTlA/a9St
0r+ffkfxej4m2iO71Ni6RQKSVYkYUcER/j7y6aEqW4DZeIUrQCGlS2PsC1/LZZhF
XtqEM6WrBwPTgPGn04d2awn8wW3e2myT/dRBr36zynhMx4v802gDz52v7z6xiBup
Nx7JRNEXe3CAkv6HA+BM546GO0eUf39f1c9CI+UqLYrpM8ut1MkLqCrjVFiDrpjq
OMmKhp7LsloxqdZeour8nr+24cSLl43MOGNmrM2b5ciNM1J3et3yxkDqn0WOZP2i
gd8fg3o3jyVlcPVTDezzZ5TW0injerxUZHwOYbV+fXBS2H/O76UpEYG8zG/vqmP5
kBzI8h5qcovTVwOVsG2vZvkLQAMUC182J9Ucubgtr25RlQYz6qI45Db5M4ooKeuJ
oZSPLsLvjThWuiviAor5HhgZe1ycU9o3DUxLWSwL91SkuxIqSdWFzoyenAEwMxSx
8WNCuVM9XPbYhtps5XfEYzoxGc6Gd5C7Qq/Ot5fdKqkEzCYXISk59/wap7xi49kz
N3pU/C3V8UnREl1lsv6qVAHvekB0eGmTJXPBcjOZc9M+ZOfQF21e4kvPZxovtWAw
/7AYyU4zQNA+7FJ5NiPfHceU8laUmIBjhMC5BBOczFUjb3VLGFQOL8lC5x6vI9Ha
bPPhLmVhHrTM1KBQ2U4t15tYjqLRiu2bytPBT1piPtIc6lWUfIlkewQ08kJb4/Kb
bBLF1A2K0CE08+8lGdV2zMC8CDkBqrvFFYoj2YT5QL33A4JM1pJqAUjIv/qK41kk
3J0NfFYbjaNDzPBCY99aCtGihuwm5GR5h9sajEGN/gdgp0HkvY5PzljIEZpecqTn
++nSA7vwCYYaXfCHPqndSNF8+LgdqTFxCK9oT6pf5E739fbTsmDVOH5BA0VBNrqJ
pXlsBsyGI/3GBiR4bmAusCsmN8iu5Hi8GgOuWjSB6YHhI8gZIvHy0713SrLwZLwE
Iw2/xp3Tadsavb070Xy2uiCDeZYv8WOXVownkKqJ1f8VI6ZgvRaOCZcIIJdT58vn
rAODxQEXA7Lc3rd4dRM8pkhRYn57nUc6thVXFQqIS9rwqHII4t+t2sW8F4SoUg7I
mh0DOCsatzmo1m+dAtlHcFCqN5538x2MhFXXNLGGlb8b62SKMs0xATcBS3oQGElK
zoodtTMFIsfE0KqOosCPchbgQEx1jlruPSiVe0rv3nJtJNmcHyDE83JdK8dVedd3
n+SSokfNLQFxksiz0ZBbSLLKCTgJ0pJw5dAfQY8pUdfoUcAtM5NBJGnNx0M1VGMa
7CMPohpxt/NS0B0PsC+EOg4Zwu+1uhzOGWbetEsh2ueO6zuFrYbM48tUr8xf06kU
NMqLCmDccxsEKwjzPxd2sRODPtvRHKFdwWGlskAQcbcBOw3+OYjbS4mjX4WkkVMQ
u/eiTsPK6y5w7TzLkdSInyEpXN4Z08n9kgfn1rvxFEdcYggtVS/olg8e0T7iD+pr
Zne783ptYyhm5HyQkkAFNE1izi3uPqCkCqE929QDBnPx46m2jFHwRc5Ed6piugVo
gM6C/59DyowXOjIg/ckPi7KI9n8Ea+3zv0jzfq/Vx8ObScAp59j99bn6azsiOMup
ciVzhOz7rcIoodE6tP3SQN7OyH5HBIjtLpP2ewNrxSwIA5YHnvqquKsCqh8DnarE
Df/G9LDRo7HdVwxnk9JPVhtgx8y9C07jogweKAkIExZXJAYjT868MNk1xqdJZD1N
XYBWNh9Biwd1GstC83V9skjC1jtOeu7wScZ40zw5xsvMTqJooHTZDJOm9G7Wup78
W9VcoLYr9FigZwXFXIOqHh8X8Abvvmfevr7S9P0G3j8Bq2/nseJZcA5ruqcutL0K
uCM1cd9bdFe+y90KTS+5Sjr+u5jjd00cQ/zpTpw7vrZDo9NVcnRMtAL496yLqvkw
u2qjtPn9KZrIuO28ucQAu83nJ0i/sp5oRdiZgK0s9NaLMimMLsdTxJ1sOVi92Hg5
kTYjjmjbjvXsCRpptI2Xn2uXx/HZyXg14HTDFYj/41KnFTToVx+oqPOn4iXA/GWG
76dbsLZz97F3CC9xs29Z0iHT+AgKCWg2txqsdGEEPks4v9hphdapspGJSUOGJZ3Z
wIjVbzpdSljHPK4PuXJvb5GhTVpr4ZIAnPQ6Z7hexOn4HB3EarNHpUP0evX7a7f4
C3hBj0JBqAAL1c4FQb8N34bxJR2LeJJpL6NKBHAWI4kXreV3vbjpAdCL9LG98Qzd
QnxaOpBpaePhjKLrxGJITTwEqlMEq9qZJ8hq4tyIYuEKvA06YP0cEHBPC14fUZkY
J/mERqs+1sq+rrrcKIQb+s0OeHokuorHNfuGvXG322VLlhTD5zZaS7kYSBZTxP8q
oUeEtNL5jnY48rfGG00mG+59JkWPjm1HmBdgPRrMmSRk4Z7VNDh2z2T5QwmMVuc2
7NLL/ZhEQ6qV64PTdmZGCOXsgM0bHDA0xD2g1ko643CTOo1UlPXJ2Ini6xe7Uu9p
cTAG4ilZX12wxJs/AHoLlz4Y3x3USjckt4W7RxfV4DB2Fb9PJvQ6bswBS78UnZH5
m9d1Bhfc3GfCLIMssOLC2WXr51czcZBeaRn0MxLglf4rNkoTqp8X+eWKcG3uuE/O
L/2ueWreOjvWgOEG2ye1xUwL/4VmtUpaS1Jc3/1uHKC+gsP9+g5mXwCoJ1BgLZaC
GmJGKch65NWdluphNWsQizMLza7HDDhdmYdIxl3f/uHOigOuMSmqvS+fWHY/8RjD
QgxRmBNi9fPbnnmoIWibWZNriwHDPCLru61bELDqn+Z5uHa2YiEw3PS3OAsPxXjm
1utkwtauNADhoqsZTgVkGYepXxbFXD2DOuHOKhe8+47Bo6SdSGNNdYqI+l3knrcz
vJjHVXEL6qdO4uMiaviw1rIUdmTtxK+JpiDy3Rlf/2GpzOLypPjEk3ZiK/w7L7GG
ZMu/1Ph8b3fStrjrTEm897KsJH99hna0WNJBD9D8zfhJeo0N2e0sZKxnFnPXUoJm
yw8PiC8yFybL7u3e2prDkoYIu3+AaWo4iZ7VfYBJFTSVvEcAwNpXZ0epJn2UrYTU
2gUQLi0K5KpMhuJIhVdYa6v0KCaqK/h91Ztq9KG+pEFpweRARZ8OQRH3OKDl2s61
1Tk/yKB+zhwEJqkqz30+xFUnGdP6HOXmvvQYNBNO3VaMq/wnSDWTSmxvreh7UkbX
9lkASW5KQfq4+Mo8+GmVowgTniyXPFVl+bs3Yo0015aQJjnYiFMa1slnhDcRIpvt
RGQmGuGkZxXTurvPSf8EhjlQ28y2LGlwBjpBZXiRvmaSg2IpXrel2CGtsMX+V8WV
4VKc+U8jlhy4R8N2ib7EJjkKFBEhlc4+Xee8ND54a8O8UX5ld4va3lhKdH+ksurd
+P3tY8QdgaXNNnqefPMNy0WnnuE4i5RkEm0/gc1LCjZdGIFokdZ8uQixaV07Tfnl
cm0IN2tT0VD7d6fBwmR33ZfZ3cDaOk7ErdH0f6dggUlx31AXAJ2Im/yP4pBG3MbC
cUUPp/9dbKINHwD+hDWQ9eXp1HbDGvfFMyqoi67gdu42/Pb3zxmDAmCxRuBftmeC
yxLAQ14rGEFa5xd+B4xx/O9q7OSNmxtOsL54hL+OKDi7CNLWGe5h0uDXdBV4J147
ODwO0rDPAIVl53ZqQx8kVbg2X6//YMT7EMbbdnSKfV9vViVHwV1Qb29zBdfvcBY9
nRoVSJwIT2HNvHadmMcGVYtUHaueXZvPJ/SHACkdw9MKBjL/9nqaDIQqeWF+OlsY
DQXXol9YUZvfHVbxmaocVDZpbG8iXa9nUvxGoqPbX1VXgiw8oBRcBjreU2MeBLlU
/isu3Gpc74GZoCUTEDX8j6x2agC/Ha2fLAR3JCNjp4yve/1RhL3wbzCLl4Vkg46z
lQFdILPwHvglac6T6iwms0BaFS4liYjcNTfUDM8X58LkB4r5+fqmVTH8xOnh8kOI
H3EsGMV8pbZKpfGW/TdAqWHKYLTJLlJ6hxsetzeFefouOg28xzAouNTFPe3l8+ZN
Gi6TG28hkz6GlLpnn8xyH66yrXGXf2MASOHS7eUhM3V5EGAGjALyTuQk1ETisMv8
gKEBlg+q75aXqPpe4hv282X7zqLf6S9rR8Fkc1Bl4IrIjQaaX2yHohY0b3JQzexA
B02sZ3LlD+7oAtiNCqpZiircl9STy1Z/TbOZCoTCcKSiheJOVvFxgxQZlwW7mnpk
BmIdIlymfgZ0FN9pf7DayXY1GENh3gEh3VLqc8g+vyKGJRCFvDSKrrWy4O05suCp
KEDzvc+fGtYTc9rC9CDy//lcXQnEWAI5ydbWdC+SyD6Dqsv5APQ96zT9kJ1clz7P
l7pc2vn9D6mZdr19hV0Fwtjb4AAQAzgT6wd5f8tT08Grfdac+bg2dlNtfok1kP15
wNIOXRgrmtpPEuj9xsb4JTwCXQ/61IazFKrtb7sbOfhA8TPdoqiDa+ImqZsRYkGM
LFyMVTnjzAzTOELrpuoaGk7hdNCJoNZZLtH/s9JAFlUKgcc3+dlRk9/MBzrMwVtW
amra4Nxlt33nl+vJW0TuQ1vYJiWncej7Qx3O4wOp/odmjQBqi3M4gA8JtHrs4AVo
f2guO6xKQBkBqGJwe/w3eDyj2cMectHABr9cpQ+iVRG4okbCHmotOb5evzcP+VqB
ovzFda6tjAmW8ET8Ejdf9jpDHYTdH29f0LSL8NwkCZu+RF8mbJVf4+k+9gKXLfyj
isUoIc8BfYbfO3yjPGErd1kgks1HjwiN4z/gjA6gyTeFTY0HWXtmgzT0NMyYdDXG
A2tXJasjZHkM8op0Uy6Pxy58mYXA65+P+PjfA8a4HbD/QHMP7+dGLBumKFU3p2jT
B9MQWACmmQneinzW5nmY3eXzJhOSLnIj5OIBJX4Pj9JbrLAc3YwtzjmMbeTLfbnX
kZIgogvshqzkJYFR8/64YgUhuOtCerI1RC8KyYjsuEFYso++ZPZW0eQ5gIhpZi9M
9edoPKR9I+e8iSnhnIrGvcKv30dex9PkzgeFZcxVqdSto9p0dCCYj2TGFQVyvFhJ
sWyHKlgbTKYiyH8pjtgbmCR9vSkjQV0hJRkcsrrqGkqVLLXP08nEruDK6CxK0hk1
bboOhULnSgMEYyTPqgkTrBbuDYzDSlSCDfLvIkx2MhPJaXwvQKNvgftuvGW8jWz/
0HE9rzpPzR2Brp5cUpAAejOvRKBi54GxifQUKKwlKVBoFVjZdKs46UI1Nm1jO2oU
GtrhPrxi5HChLP2De66hhAaNa+SvSHXvMl9lLVIuqS+rITvDhLqUAArzA0OSCwX/
I0l0ORksr5cQsO7/xQATFs3AOkjVg+QPQEWV4Sr5Q2pT5p5fQm4417P/bMpHDpOd
fYtZFGpzKdr5Q3biMX0/5zMYpqDK1N59j/VGB1ELBKPuXHLaTaFghWiAUz6QXLit
4Zh+hvweKPgLGpYsdauwKKH5Fxe0FVCeRstTMfL7VuPyePcELexygr/lN8Qdy5CM
1I98hTjv19vmKRn1cpKmu3lAGJZC9U/144Bf6qAAPah3IQqtD4KiKq4PRPs44eu5
Zd0Pzyi3BtEonWOJVWN+5G38f8mPZeQ0vxDjbesG37/FS3P0FrVuj6I67SGDUOkj
Wg0j7ci4FQGPVBkvDq4C69RXujYjLS2XOaW0yu6C1eStfMyTmlqKSiu+vcs5Mno6
jaE3aZynw+72+MVpQEPWf0VJg3aqJpJiiDSvU+wdN1pjR8jyqb2TI7tPlKGYAmXw
l05n7iRXhwD/hMRDrQoMJU7sKtljWyAmF/2ue/P5b8WVxpxuiQHjfc5wfl6gAEiY
5BjTygw+1LULxeJnxqrOw9LS1eQ03Y9mIwrbeT+o6czG6jb4SxusLXuaZ822U6UM
xZcsMidZ5hpNeajZys5+T4f7Ovf6Q0He5gy+Nf0blfi21KF9BgMdbJv5GeAYvIz9
Lt3nF5z0IXAqWE2H3UlItzGN6gDtAlSdEV/+bJuuhzukyrLFP7PpiqDoi2aFyTBD
LrBna6rsVVrF1icOhSrAJ8pw+Wd233a52vOiRUMb9xFSMp92rg03AxId7Behz+cL
AUBJg+g4pRcBnrRF4aH3PC9Bdp1WahEWpVCF/xiYol6bAV+YSEOKK3P/rEtYkBXM
+gqKfeV7yrZikdadKOeVMruolxJXekNQwh1wMKkGkBzU3XwYixr1/Zhzh76RGnx9
SQop3aPBwMQdqWc5hWZTJd5wbvMGRGKlliLlGSererBt5BjnSAS2o4BDAB6X4+Yp
N3HOowC3pgC1nfDWxwcXRwklrSVS2s/S6bzcPAKLsWjRiTU++AgrEPDdcdFO7JzS
THlkSWELycoAIrtCbR0Q74vHkPFhTtGAQhhJrIPcAwrLbAl8lK6cZKhlExgLPCnY
W7+ouhR3EWNwz8ehcFWb0tEQr4SuTODatFepMj6h3xvDGNZnQSZLROziQh3rihEE
Jbwddjrkb7dhGVR/3WWHqPQyPOAuYTb5Nxteevvys7mPLlGju2oSTKo91ViOXl+o
7um81rvgXlvPwrR3nuDntF+/vwNlsU5CUCNRFRHO/uWUIN4a87ZWl7YxbFBflRc3
gpqmzOf+qK59+Tat5rrCCExDEg9lE1oObz2giKGIey+vqvsTeEJphsdUszPN88xz
WjfDxwf6+vzTFLnrVCWoiDBZfQ+apBTYntcQ9/n6OUlPCbCRhsuD7Rumv3J6mg7A
grpOQhpDMiJfQNl/hrtsWGWZ9yRORs73c7fDS9vQ8/F+jqV5ic5MUt6mlg7bvzMi
DvO83O/+80qhEHCSdzbdcXc9QebsPz0Plivwe4O7fMcfS8nQP0CwJ4sgA2hnq8Zm
+RVGa+21LWj8XWuA5A8dvC5P2si13doYvSrdLDXKa3POCfGX3h0YNOLHOaresJDE
j8naqRkV2o5hpTK27NrCWIL2fioRjXY5avZZVBSW+wFxcWRZtZTwV91faTPNJbdt
A0uJtGTbfow+XriqKGTrmWQaNGThmWmCy5F1Ej0bOHXux4K2zmuAg2vrvZYzv74j
DIjIJRQCP1lNtlNlh8NVzqe9OsVhPPFMyt4LbFgkDa9bCHlEvjSz7HUJnARh1VC9
qTtHGIPr2xPEF10S2ddxcMkeJUeMESh3UVrdRUvQ5DAqLAx+jSoZB0/HJuiWareU
wLjXmoqduwliP4gLl/6IlwHk8sXDQBYHi+6zxpue9diqco34QxcavV/JFBb/By+5
jmf9qiu1RD/hGm3bae4gGSIvHchPQ2uYEHGy/DNpoaw8hXI8xJwZAKS77oV+ID9g
4L4VPGh03RSysuTzWA0FmQ2ydLzrqFsJae6PHsWSSF9Qlzd7VyWin0sOayf308fR
qzJGyihTpNaG4wTQ8TJYOisfitRhNJGKH4eXiN1s3LrZ92ed0aOWoJ6yKkpE9Ye4
d9vUG01egPynjMArjZ9bk3ehWN+e0g23T10VQycxUAjlmJtQB8gQQXG6UPJoCpaE
6yjkLLdLSsrmPFtmglJrs5Ib6kjuhg152+7FMmzy3F4DTokySH7fNHBeJ3qQrFBZ
0A/36tB4kGkg5aaKGxFVCVaUpGVB6LQAD/pEUsiP+wOzTg66GHZIWPY7U7P6bZWM
yGfIOqjjEN1yKZ0KIZAyUZSBeA+4Y74U/iBdTf0ByPL7X3eGfJgDSSmVTxTPmVWd
1Q2Y36lVlcUp2C4d7mC+sV8qzk7HeHQoEA0NnXEElvStUgO8zUjPOzPYlaRXV7QU
bWl63XCZrLm7ET2L5p/Gz/vXsEHGo+WO5zzXqhiDR0a9fPP0K83uceTWvYJI1mIJ
hjX4tF7jlXigpQn/O2pZilMY564nHDlhYnBwyQMQYZyQ/Om8raB4OBwkvDflOAV5
fsOmgwXtZXwCs4CsmuEn23K5L9pyz3IRqMiZa6gMIHZ95vKfXABA2aebq/fp0pdO
a5QWNghy2U6awouiblq8XInllyA+bFvkqRKW7O37wgQE0nfdFpNX6Oxccbk6u7an
EYl4VmP6RNq/OVBkWg145cpf5Lo7eGwfxPc9h6f41+TqldlEPFXUccJkKlB4K6hN
C0xZ8B2zqPKbrxIHi8Gd02CmvpzHZ68PsTujs43fU/JN9OGKHzdCgvzGz8es6DiB
1Zg9YlL7xWW6Oi9dhm2OkkoUimk5rXPJI3Vm0fl1oED9aF/nzYU05TklPUQAGc2Z
z0VpJ9ezhIYevYOxSoU1z+8esVG+AeUoA9Vd0WTIPOjnbRzNGeR85tkfSHVe2hv2
3DzXutwdpb8X14GgU4IXopea4l2yU4+Cu0hYdIDKYsM5Jz6DgUe7SStqCznovjlr
F6kN/iMFcTwYYOm5Zo2pcoPxXAb/0i+GGJ1gTnajg3FrPJ++pZlHQdsvPAlAdgXg
lxhW09SfsSSrVAyc7AB0SuX8Mf/UMDpMRpHEbE/FmLKuAJKfe7GjpGw+8ax6OxPS
sVsDKBRBs/fjcSzq6uWGHd0Jlu5vYcBWouhZNgQYv8zVwaIzY0oQmuALcbcoGsc6
QowTFjuN/oR+k+i0przshAJlOdrLlZNFMomS4ZJbyvr0EzcRMpPbdGY17b4LFU9D
cqVQwvpoKVYP02HCM77G492jmbrc4B+iR4+CVCw68t+TOqOLcle+GixIjsv8x0tK
FcT94sIfIGpYLiRlB0L7SAY0UBjUBQVfPGj1tchb4cRYvVHOuq/3TbpzU/CfHFNo
FSYLcCa1SOADKMgd/pqAr3SdDVVCVnpWkzxh6vuu5xu04bYM1RDGgd5yLktLiI3X
FmQn6rJIRVg5m0t9ewFL6MQVby+njhO2ui993Jq+/pHLsaNttT0UxoQR0tCmdq23
xyi/+YE6+s2FE9Ox7/cp2FdYNAoxGHM76UNxYIZQn8PgX/hwiFW6WPhh9ULPoQS9
btMZEQC36IRYuy/vIxLMXQWNz/hQeFr2ZqTiNoCMmoypPRNJN8Lx7cBazf7bt/GM
bZvMY1eK1s5fR4bUJGYQhcTD9MiWpuBHvkoyqAm/TdTqsiL8IzNI9AdjAEG2S7b4
11j/pk4i+UJG9Xh32pZ4WWSzbtjjsfBhByxXpaTxKmPveuJJ1TsMBON9Bc7Ds/a+
l4zUwwGOLxgUhm+LsrG+BkWUUFNrS3wxH39FCfMQslj54vEnt6l2Rb48YYx271B9
Jmd8fmD4DEEFECJ7+civ5hbL44CucbPw/eBE9fIrh91BORZUzTLOL8VrbJEL1WU8
63+fOo75LwO/yMo77LmXxXv18GZpL6LJ16+EDi8XWAGAfqcolEfunZoyX8OFosvA
32gfE0hJq07BMiNw5dH0nghxHxOpYh5g8EDIgc619941Ik+dTWxJSe/SY1WEyjd0
Z+J7q6h2y+1Z6isUg609lQ3/fEDuzRScT1lr+Zam73rUIY1pMTAL4Gt7IIjdcGuv
+pdnjofDbrAAb21a/DNlJu+4GwUdFQdPh2E+USG1uC1rPTWuzOe8pVyjYi0M8wC+
z4ArOiad759Q5iUdERMknQxALf0ndr5cEUG7moRuZ46EpeyrAHiIGs1n5UzygMr6
wE0bZY06MvMmSYgrN2wM83eoDO+sPnB86a+G4eTDw+Rc5BgiUJhPBrpbWUjAfphb
V6VNu2jPxipx1BszXtXOyF2n11yGzLF42yu4mbdQZS8u8rxX1s/OnXdReknnInL4
a7e1b2mBa6yYHdxEMVsnvu3rb7VH6Vy0sOgG9wu7EZRQlK+TPSvz9qVbD/1U2+Jw
K3AmjGEpsSMBqOlMGLFb4XMyaMQBHhHbgRcffT7Z/RH4JF4X57385fDVHulpfEow
hrtjaxse/lm64ZkbJ9Ol4qsKKLqOxU7lolVsUvDez6+Sdu2tyIGz0r1OrPT1hFbE
TTE7xIxLQh5eCsyzi/8NM/fH+0YM6xuSrVS78zME0lksaOONE0K7XITxZ1VnOZeO
3+D3ZjHGzza6BPwKJQqXtpdmBXExSD8yEreZjwKA5cxDKzORWB2ywkWcIAnf62DX
jeueMdAA94QqsceJ2ailSlGYlMI9cEum2MbTLere/gb7XF/myCHrPO1VMXsZ6zVd
Q8/ou+Zc0Yz52j6QOPwdHMMkbP3aHvnrTR0m95CTUdKqenvWH+IlDF92XtKD9s6s
IvuTuAqNZxmrlM0akR6ttY8tSPQhnMSpyPmnTfqkoFBdf2r2H3hOFJW81hQJ476n
qdnRGi0qx9b2ZnDVLiif+XVwaRw2+LKP5G6RdsZ7CCTZ9f0D4OniqVBh9MuS83sL
23WFYLTWcX7LBaviJBx2WdtB4/sF8/gaBKLB9s1SjpVMfOlFp+8oBeQ5WVbvN2gl
Jn0yghRWbRf/iB4KQ+DjwtZi7X0YwdaOwjmY9sm7t5UGo1+qmJ+dSAF49Aj0i0a2
aiO8wyn53/vraRYvQMNiO3eOg2lE9DVmbXh/Ap0xrbcPvqkm921eunNUTHpW8LD5
UyQhnoHXUAKdQ2TI5F+Yj44eWgjhVD018bRKuNiaWYs8wDKMR2C/Nio1qIAymdAA
OzM2+J5gDFCU2NOs/rB4iZ5PVRShR+KZLISZ7DGSAqgmkg4NT/L5eid3rcLDd9R6
yqwyqxWMVMgS//bqpHNP4Y0Gk3m3hDIo7FL6bkDExgAbG0E6RDCZTEexFq0WiWOU
0f4FqQctyduVMXIcBKcER8qlb5THmiqEylNInLOOUVi6umTDWnJhRsYlaK78WGM2
rzi3YDj6CVTVgbpGnVg5EHhqsj7dRDt+SlI6v7NKfmvd0Dfd7pUgS1KgIgc+pjfK
PgEoea4jslVIXjo//CEQA8ASWfn+eyGSv+G3DTMN2WCD/rXibStG1L5Kjl/ovlls
utgsOvRmaIDwPtRIjv9weKBSEm8STvJOIwAtLDx645DsTquXwB7RgdJnLbI5C6NM
gqB6AFjSkm95RoFslI6f1BKiqgBRLV7Y2vgYi+QbGtcvWo6YDKuAAKfP8pJah05e
xYvUcb0SrzopQIBS4Iw0Je1z/23I9YZ8p976EsmFubxESTv/Dq/nIlFTwVccOo3k
9IQnQc4FTje7HohxrnPb7xiSXrmAxUKv2iE40GcqpLUJm11yu2uAfq6ZbX5immO7
0TyMF794k9jNGViE+NdRZNtpxsJsOmSkSF5MO+Kej1CkENiOw5wqHgG2K6/3uVtB
IetDQCR/akKaWLbbw9kUoAL4EhrzdOxF/tseNMh+6hkQaO451gBBGjZ65oQDnYGY
NhEGw0i/V9aSGeA/eCpQEnOl9yXown9fWd3H/tkToCSJ6SrAhQEORqMcDMoNxcg/
hqJS+yC/Al/W45GLwg2wkFR4CLoSDUJy9ARVjPkldiQvBqToyhq0DRCDghIbC79V
CsD3AkCWWEkkpsxEdbsJ93Fr2gR+4LYwsqmqxXmuoWD+AehSFMDXXngntBz7kwzy
WI0KB6n5DdzT8pUWLDgUKOcDoKZSxfiJXCANiD/Bg5fth0zkLndxVTdtzslIEed0
sqkRl5gvN0kvkOeHt0WvBAOFfP4qDEfbjHejDdB+h/pWXU/fARBJeDkpJKLacWeZ
M9+1CweBJXh0h0y7cdZ0eA4GLkdwJ/a/cWSNerEe8NNkBpQSslTv10tQxhScmYdy
G4OpjwbWjVFalYUTg0blcXT/i+ugyO/VMpU/pln7orrSZ3B8hQ5q0vUQTMHpdYJw
uuM6Bq4+XzVUJcv6c+3mZu/H6/rcnoJyB9nQjHpn9vXqz2u2ikuy9JCeLEqFZBsZ
I5aPVF+GCcZCdxvZv7usyXwhwRCW7+fz3YNgdsyEtKyoqQb7XWed1ZQgvQ8tFf8H
AQ339kAZ556PF87Mkct+OZjctEGMMG/yX9A5spNIRy2luPAAmooscOPxUSwBiFjP
2lzrFT6Ow8n/5e8KbTWWjHQ4GIVhmROx6LXKaowmAWFhAm5Ghpj0R4AxikSxIe/c
GMaYbbIfrXNmq9LEkH/Zlzr6ZErtYfaPEWorcTl0IDGk6UD3K+/vnZ9beBjLu13N
RCnF52/dNV6JQn4VdJlFOtFUapuEUPG/fH5l2H3jI6FRgSWnn/Q/5f90Bwh8agxi
AqKJlRSnM+DVJTrL52CWDNcWviNpVPMCXHsTawo/1xf+7N0UE1A7dfYH8Ws+UIQc
adkN0R3GnW9uKrBTEhrz2HxDzC+F/RS8JrBBdlz4reKPGg2cXSXB1HGG7CnG66VY
nKFEkgj1UP5TbumUss5duf/hTdj6TF+/3AmX2x/n97x2x0yK5AhaGX9JqVogO1OB
3OqLLrT6m44ayd67DNfVVa7Eewjiq8YGjZwmDdxq/ZIkTfQZkz8eOO6wW6rCufIk
EGimkYoP/XlItGLj5/TK59YMFmEzr1K15RX9yJ4ytlhtjyysinwbUJiPhnDFS6ym
I48ffHmdL1udtculixvToO40ufpb9iudOD84/EoUody5tYuhnX/1sOTiYgb419LZ
DiGYYPwN9tFWjWhyqQ4I1MyKFDX+9wUqnVHMPSoZoaHkME8dv109zCbj7kB+r84U
Ti6TTLhWpqm7cXC74/cb7IgKL5GvTyEfWVDsCITub5eM4WDTZ7lsz8j0QgVQmgph
ZI6o4w8+d+BibGGisj5PRHYfOhzr5tx1DKUq/MLtnSc8LZj9RjCpEiV708xOvjbw
WDPTxJ07mOm4hwmA9/QJBMlGarghk8ANDbr2iLt1Zbr6T5kukU9IhR/engB5V1wH
uafI3lcFCun1IMm6qDt9hk574BjQgSFy/hH3AwTlCrcSsZzo64+5FyUInKJWV1gP
zJHLZvu+2eh4O7TmQCJKFs/HmDtkmLq+C7sY3bwqcRagRFrMNmeIWJa+0WztjlvG
H5/sU+TltwMkuUWTFnC17YkS66GPVAJD5/MOyyu8rg5ucktwVACMsYGTC9NOPKy1
Zlfz3XNSlL2F3B/ucBegPKNUB/ItctlKbTpWuY1DXICYXeVgLjWxgOQ1WGnZUGXV
DznnV9aQZJWZQySj9gBgCDJnhFMfGF2uEvVEXTXHbuCB5t/T7TWl/CyiDVv/sPlB
eShym+FdpcrnKB5+JDv0BfJLYtmueyXCUdjq1oOnxzN/mZ0w3AHpDA4CrVmGFeQ0
GpSATRwtnZ1gyEHU5+T7Qt5+btikJTfjWd2Pm3XKRQBxC/hgOa7IEkwWzKk6wOWn
j2aS6Lk6LmoSa3rpP/jkEhJY4ROLufT92zA7Zm8h1OKhHhFgfZzGXLsEDnh9NAxg
AXqwcHqStWUCTaQ62PzSgpxHY2sR5wgFxqB+VOlo1IDZZe+3DPg5GtUFlpy1Fsu1
sHCtd1IB/win7qCTN9TZgNgaN3j454OrCiM+tZe2nR/uBPWbtH7A/ic+nUEKeJvu
yfjZcGDsPPOsHBZGe048oM8rODIjnU6cj06rDBWLhPXT2iP16Bp3vXn3ulIakgOS
YbK7fbJvhnXB0WUreZEr1GyblWC8epb28UUxzW2cYyWdPtFH/T7Avw8tKM9y89rh
xa6Lb84185J4CsfupC1M7FvWs13r7w2Ilz5nRWtESZ8IB9lXvYFsc0l6MiKLlVGq
lqGlGwjv+K1R7ELKVe4sKJOZwxY2HC1YSQmykCUmRX1a7ztHweWsgApS45pS0hKD
bJ/heeb89mDXYbYkE6Dw6GBYRZ8DTJLFi67IGix5HNA2GCSDO3mV4lqSaM8AN4Ii
/O1vBl+ZG72D90gsvVv+tTAwL9poHAoXGA7GWTSyqaFLWlP3BvUiown7FZkD+Ugm
mxHH6dJmzDtgu5aQqLLm2XNYs3mxwwGWor7xpbvNCB6cB7pT8aY3NZLwM5ipWyE3
7r9FhwPUwlY9pCeboUyVS24vDHDHxijryBlWg6hFLtXZZU11iBZenYD2Ym4iTlJM
6IsXFhah8V+f/CF0HgqUZ1+udnc8GGh+Acl3aPVtR0shlCtaPr+TFpzku5TY0/0K
dNgp6Yj0OCQ4WdueC+WP5eJGTPUOhJwSNCpPUH/NA0Un7X/BzGDG8OZW0vSYJGIf
DZJXrXpYC7vSrqHwfHlhcXKMBRgS1A9zPLEs5okHMGRjSb4tkaZELyMgmkAETjWn
HyPQW3TD5JyJqWFZ46xu4TJWzrHCoUInbCEN0/zEGLcjpwRZ3MNs7dpb3w0gfULz
Y0pg2jXYTVuDR3aGM/B5eVHX7C0a3rkoJzAWTdi6vW5T46UZRJdyqpgfou/tQj2e
OIhMNJMMA9LDiwTzBIO/75yVUWPThXYEkAdLyENHgQMreD8VLNNDtsst8cfgsRN+
haRSsrUKNrO3fkrfaa6CYthIYeu1Abo/KItYqaQ3dhwqz7p2FPYbXFunc46UVNfW
q9pDAnqF8+sfIiAO3YClChzi8p09QsSRNGw6jY1aL9ajXPBs7D3/KvDKG55ANNqZ
2A163kH2hi3rMAPt88wJfgqDkr+0L6k0DhY8s/vL8tBiBHsWQDy5JFa0EHWZ6Z7p
F51YvCQCJbaImsOcYEJ77UZser5Vo2kXak53OvG8E06LhG+DBcZ8Q2KXnnG3j+Zm
RLAbWxvC8L9Ccn598lAnSvWxYObubD8NwbxZ/+6JrsZU/5NNfvw7OUjSRwkwLSbe
tp/a+WB2GYHMT0zXv9bpPJQUXkgn9iGbCPMcK5UynS1jJ+FqImCSVsV2kP069Y9B
/f3FqptnC7Ea0csqrWl8LakrO+PYevHR4k47l1c5muc7rbn+MzvZpExVkK3qNmJr
YSbmxo09gTkcD02EOyLJWfDeGcx2k5kTi89aFHIJbOu9f+wRRgymuV/mZPRN4MP3
lvG7OHFo/LLbxAQJS7oUuHBVC8LVumyikCgoTJs+qx29yOdFW+zopOI+NP9Uukbv
GizpcrCerNA+O3jtBA4pDisSKTFFaSjHENzd0G/VVY8xgaw9LJI96ZOd5NCOifpX
pn+QGD+yk4PpoNHLJRLCfVkQNJXvPgdIgmDo8VcWOkmfkB8Po3I2uRE2a42vLosF
z+qG5cX6a35Jg5KKSWxtZ3L2v8AMAAp6KzyzvBQkWtDx2ODzby6Rz+T9oMFyw5PV
Gj5EugBjlXTt6OTEBFCdIelL+m0TzvsDwisPC8B9DzlW2nfpF33pNaAIE3/9Y52C
Ncvr/wWkECiTQWuQTFJhgO0ydgfSsyiIC1U3x/iUlYZVaE/SeWIKhYkgjfYa+vlZ
r0QW88hIArfDbcFytbx/z02vt7AN/3mtB1kF426NxYNXN42zn6/r8ZEV9WJ0eez3
TutAdo0wWnK3iTgqaCLusGham5S//Vagq+oF3hW0OQPc3Hi6uidAHyU5+q7y35eO
vx5laSHt69ghhVc0WOoRHpQgvtptCstXfgNQE/IG2uNAC+8cdD7F00g+Ui8COogU
XqgdR/F9TkIDmptghJLnyaVnFmq5KbWIq/rp/bT+dL/GEL18969lO1qjcTRs22Rk
wt7DexqThjAtZnG9BUWcuBSwqMFp3Cm5QppGoVg39C56jlhSl+8dFIw3bGsKFz4O
BPKRvqWmRH51/q1uXuJLyhpKfk8jaUBzY62wTBqVRcbabqEIPXGKmtuubf/zwpM7
OIVnyRGbb1bl9MBIVTZy1mGvmNyufIHIA/VyewFWu6gXhCymNPk9A2hri728iMqe
8IcTc3ZUzPHyEZBO9QqsHKPL6yuzaMKuhpU9pxpRhdOEYmmixCK8CN1G+0mAv1DI
yIK8D3uakKiSQ6kio3MqNQGJvFF/uRygrmXqRfDBVd3cwT8fb3yHin3hT/bPFtwF
igBNEMyQ5jhYSA5EE7z2vQ4cE9B0ORn/4LzmZ6Wktp9HXq4t+qcUE2sFlWbubKgh
Mo4ijNZ8++g1xR5TkFC3gBHbZ6omR3RXlBRTee+yl/W4EzdzDUOrvefFUgIVXmYO
sOq3Whxf5xFtosUj9rolIlhhKOOgtFsbA50ZnPYtWQ/gDQXdt1gE6oED98pHynqe
RXXeDOT8M5o1g+KJpVJiEdztOd/vIBeS/fWvf4SAfzFtEdi35ex+tStmwlmKUlrN
wKomJBdFf/WQ615ZncanI/sUmQ8qY5+nPmori//cX2SHy2oXokanIscLIHrYA0pw
E+WSXVMP5bQnFmL/l2IJnhT8QxOhMYiRskGmlq+iJuhshZ4XZxUlss0HLoXF/lys
qCzF95x0jhya3l3we99pZW7CJ/uiePXD7X7HC0+UrdtqA3eMcsVSJctrDG6ka7Rv
TishU2d9dkD5B9UPYcjVuqTJrJl8GWuhrq7EUHxaMfgqiJ90QY3d4TzRJef/BDv/
NU9OyxzNwU0uxZf/JdbPd4X2RLHOZfIcmFW3ffzj9opElJkLr9U73pcv8okkWnbP
7S4Ipcm+oIEWeVAm81i/X9O1Dyf5WhPwekjvY5Vdjo3Uc7pR9eiVWmP5uQxiXEev
qYamhtfgKh7Ki/IjnWl6ig+5+sVfaLSAOLmLML+LZDSaP19dw3MjBUNqsmo98yOB
eFe/iwhT7HJBlwB8ALYM8+s/W/hZjM0TzNa5dlCcZXVJj5gcF7ASHFrBq6AfkNSN
yRI1e92GEW2U6c3hGBqNHJfZtnLA9E4jJ1KYPqzwzA5VXNf3UjdEE3m/8N2A7Piq
zEXeLuwhRnlGCFg2QzhBD8txMw+95FVPMCUrqAQjbMdgSGQqcoleAW3QRqQSDzd4
8ACYXnPyVq7QKqxeYVcRC1ZQdledJ7/mmS0aC3D6iqyVdht8E62b4/s//ZxYfEfM
CzQXxpFCJFFrqgLRExCS7KLxqKVDApefQOrdW0u1noDTN5fum2gBruVSHX8HUt/p
myAEeD36tUFISvEe/UHzkn4OIWUNxHxGfyNMo4cmSIH/qXoD2pEyZMzaSjNIKmYc
lDY+HA9XPCO3ZeHponmDxBxmueRbYqLuxidnukxRdtH84kZ7NJk8jSMpIuR28Lsq
vhMQRDaLqz9foGabsxLLtWwgX/olOUggnyxyubG3vZaLOWC2k8KgSWM5ITEnfugY
N390REx5PTidjNdvSsjELC/nDBc1WBDCOlQN8p+2e0SCWzTBBtwI+plGh6UmEz14
PtvxooybLHjWcSHpfhEG9eoyBD6EBCLjTZ1P2QKDg5gvvAo4hD2nKkG9/iEo/wCU
IuFwzLUgNf2Ff26fhlfLCtx2QaFZYg4ewIDRPC+nRiGp7GggJkzPcmTcYJHMy9Ph
3LzDbtUhzwdwlC+cSrCfJMrohBwbj9gz49UpmqNzFjunIdj1Y4xaCk71FnZsY/mk
ibWeXjMI9GHGadq3nwlWbfv2l49FRPYUy5JhUkPsPXB6WzOaDnA+mAaDLx8WaKil
kXLMX3BT1XsN+EgI4SlMLqdmcVJ+Otyca4VcBmEPdaqqo3ObExVlmiHEc1Ax2lE2
SqvD0e50rUelo8g+O/UoPeqcEd/58mzjiPyuaPv9kEKV88hsIghPnrsH5jDKucOT
3FVz0Z3WoTQ81y0Vx+Y4c06eZ+7WlcSo0KxtJ3idH3bQEIK1Mn9fXzDNhc/pTE/w
hYTqZ3DCsnZExzbFyWCECH5oV4IhQX1s6WMSecKlLLN4IhCC68zkzI63wUyDvziy
V8jB7x1oLcPJAbUm7Nfg0RrWPaOAEZmFUrqKk/6yeecPZL5DkfhHj+BhHacNsqIc
ZkKuYppG/9UmDChFZIIdw3VN9aywPlPFcuJ2HZedIKDNGpLj0Ju1isk8md8x5dH5
kB/voD0wP4bJ+q4Xbt/y4shCDb6aUJEVdu3d2MhiQEbyv16SxVZ1b0XuL1pl6dGv
rgnZXkzYOvwFpRiSqkINFblrqrHvKIbKgt79kgjqZiJbfXUWZPsKZS+zPN5U/kt7
WmOU3+B0qNQ7UUDhb46KIWNbxT7s4jhWZMxUZlUBpJt5i/yaEXbXxXw1IuowHAbR
Uotcf4jkhWP2cXPkltiuF5XIGBbIEd9zqP19GATsQQ2oyiIQGvlUBrVaQS6DXJ8H
YE0gK6gBkgXPjqJh0Azo3ZNRTVFumA07yRClhr9sGS2po6jZVnTaaJ0t3yWt4uTF
AnSHdiB+b5zwwmUlDSQ/QUnxn1IIaFgpGO819myHVBGQt3XfwZ5FCTXoaRBtAxhI
i7egaMUfWI0oSXejXoiM9jkGw5ddQd2DJ60It26mZpc2ZhUTXFGBQK3eE1+1slzk
VvzDcPNcD1tHiZ8HD2a7wXbwTd0AHix+xHt8MzUwxOMTtLr35w5wdLgN0DcyH9El
y4R1HKOYjJB0Xn6WpSenbujsl7vW4or/P2fhpgmhxZuXjpCq0/+tQfeqhjlLcp9m
Ko6YjS7jL10axF7WeI1tYEZEzCKm7sjRxEpGMevSXsAI7W1VtpckvJdbHftv2iIR
zK/nLSCaxKFZip6kCjIguBYk6DmVvlx75DeiHT+tKesKgzPQgtQ0fBSM4ry5QyAh
YClK8B7OMvTQKO3tLNu9wCyRPK3XoNHnZng2c6do33n8DAhK++PyoiI5NoLmJaKx
iAEvR7Vz90ZnA24GiakBjnTBZ46JYZFm4mgq699iilxwkwixPjdvr6mZiwXzRgso
D6mF4mCixWiuerBphMRgFEK/HNS/lf4YvBsx5RVK8gF4y2bMc6UhL6AUx5pmJvb8
m1bi/icBtW47hro5xujfhTpN5DQ6t3US+T5VLyBezgJpeotqGP/d2Ll/pUfoszAz
xOZ7WFsCBFwsDlF2LIgsSUnXWWF2bVE36hChum6chJkhSCLqolofNaWg7F3xUvjQ
apKYJVIvfukKPUVvKeyHudAIx+lmXgdZZrG3jgt1PLkviMpsnAFn5Z4lw+AOCjoN
M0m7Uymw0Ow5pg5k0RD2WyxcRKqHLIrqf3b1a0aMO0DdMD+vGMjEpk3JrBEv8ZKp
414AktOhqxh88j8oP+lyaEF/2SVmV1BfMKsiA1E6yCYf9nd7kq9EG9BoNIMYTqBu
Y+yT3sVH01j4ZRNJZxH5xVyVAfh7di29O3WYB7i8LdHuHn3n1d0hRO2BMZZ+ZFCX
ALgxK3hUQTEPpiR3hl/kGX7vG/h9ZDhVCCFTGsWVwYRaqk6Z3U50GfgHrJdXmicU
IGXVGGxwg6Fzct0fsYeps0uCwTDCGKLOgKCkh3V5Up6+rtvQLToT8MODxZNNyRfW
zSYrKNYVUxO7XkkIHvGD/VTiYnwXoTz7OCrYiGRlSjE7RRpxjlSZnlsSPQZ5z8ML
dzQIg6hhHNFsHLr83uHS3a2GP6sgoMk0FEh4p7qq1oYXAOuKmE+XR9YiU3AuiaXp
00WxOvH1eDNXUhdi6UAJpcc5YRC4IieBVpEpfZAItzy/bDdSFnPvWmeepYbqzLmX
bSFmyRLv21EmaR4JCsD3i7T0O6MYjss1Fm8vqStMxMj5H5sDI0XTNHRizK+5VA7K
vHJczGFRICnl/dm7/ifuCTfDLIC/KANfnRDLKPItYkcCNGDxbM+yC0u/EPJwUDHl
U5QkHCTOrhf2M6fX0DMPsiqyKSb3kEHjWKpHmzcx+1sw5U0vHVMfZ7unXcZl4Xcn
kckPU9xxTiMZa1tQzBtrCNR4x0CblnTj5P5rX0LLjV40ngzg5wPxESJy6Dpak4tg
0pvV/rrKDxAd4u2G1wkWi7xpm7m9eDx7/4wuDWgGnBEA0NXaHWR70z2LiPj3MDhj
Y4Q5D+49emD1gSRfydvrujtQOM58EiL6euxz2wPm/xC3iEP/noxjcacsZBZCVZVO
vNwVsJ6kN3WLPU+fqUGRBH2vW+XWbKd6gcko2/4xFt5PA3/PlUKMzZ/9y5n6SBHU
5sYEG/r82r2YGLMyuGbgmWeaHLps2SnVtuoyyrMvm4m6yQ55YbnnIRMTt09zoO7k
/GYxjll24ZN/7XNmtunicPI5mLpq5gHaz8sHx7jJOl9InHfOGMZ+F6Ki6Ylq5ids
SWDnyz6fo5hOqbfAVjHuLQ/LrY3gqCuwf88bxavVNhuEi2Okv573dA66z3sJr7s8
ZTPq7j/b1vwxigaef9MJDeiRgT5z0x6TWRCJRUR7fL9ZqqfMIO59GG5/RpP9ikOc
9zwJZKGgmXTxXc8cC/HlloUrqJp+/3mqdk+UdFMgwhfPgHRv71XLlrzMteUwH54U
LGlB8Vul35v0rK3I8IBKIZ3JFI/aY5LsHh69b5A4GOApItI87fFdS+umFprv3LRP
AxazjGL3L74kug9Tkk15TFrq5zPgXEoo8ONH+efO0qF7fXzsg5GyoLpx86x6OxKg
NmFxyRIhFAw+GnI7a9SljqCZ/vrK4uydeFqIQVKfnNC9ujh3fVjau6QYWQ1kp8ix
UnwvnQR0GnI1lEWV/MRUi/h+7sylRp7DJ3hQ2Fmo4WVLy7dwLUtjI45myIt2ue+s
aQm7e1MrknDUTh1IfwcHia+xlXC9AxHxVHRqKqz/f0ERDPVSZHbyfuJtcxAGT0P3
KV+eOlB9Xk/A+4BuWFoHVg3P7dxaJyWtMCVOrTqJhcyDd3GwHWZXqWLIqa2LxHfC
NR7JkYipEI2BIeNwYZJM0MppDmuXpVxlsxlQneJeFYDqzmpaW/2QVs7NmXoM45XJ
3erOCFGO1WhibXS2R5oNj6mK3KfLyzfsixJ7DH34ufUsbAnhmkHrfMevxZwtkyGk
2XGMiLeZSuhaLZ9uroH2ylbAjUHgosL8Jw8GOlSbdgDXnBtu/nM2nbXD0ElnTdwq
0nhYUARr/xoK7GcHfptmu9B73tW9nu5ecGiXz09exNnUhV3VsJGZKBaymsnVTERV
DcFYg0r93gFn7oE4Yh26p4BsU05t63Bz6T/FySQnw8rn7xMs0ZDncUl4UvRAgHRS
koh1KCVvYyMyEqOUHLjn+n2Q+Qet7VGJzxYX+dM8uwcPTjucb9jYPivvvNDLOWGf
jIQRRTr89s4yO0pT5u6f7749ORgFYIL5K1C4iGnZ2Tdi5UC6oNmhPME3+pY+1Jle
S4r67VtM6VyM5VbgeYrG7BugCIPBZ19zUUdCB01phY0fR874awv4eIQyoXblbFAq
izpu8bMb1ZBjQ0XSe81dVcmA7dFVI6kNO4CiZdfL3DE0VWCWj5j2HcR83x+wJa0J
k9/xSRHDXblsoeZz7TEIs93WAgl6iepT49CAKmNkj9wKxZUavRe3eobvdhmwLqfb
S0Yy0GylZBtXLnWnwk5MjJjlEDTcNchw/2tHiMkYFvHpAzBKjPYNmWnHG7LtamMr
PI6M8WmoIHiBCiN5YQcDk3pQas3oyIw2AIV7Jkifcf2sKd5eRmAC7QGkY85wR2R7
gu8t68xxmyvUK0Y+5xBL0jf9DTHKx2mrKjtNadDJlCkccM8n6uLEbZqNw2lm7//V
dmT4OwrJMmDHlXPi8wTu6mzqfvUBBcfLHV7thvS1d9I6QAY+3MoFPnItRkzfJcYW
8q0ZPgAf4FavekjrzsuoemSaLDhzHnu0CmW8EkRDfMtzp+2/FEcBsnRnk/Aqw9h9
xYcV3PVSDIi4My3y3XGZMmmy+gII2JrjcJIB/dN0tjZqcgkT4B76gBTjUAX4pCPE
pewNkikMBKnEtc6JZ8VNtibKzVKJW5ExU/Bp2Rkdk1M8gdsc+z++MvDjmKHPkciM
rx+pavst/MnkvelNYIQ15l/NjkaSSo9/Xqfredb4KJVTzZUp9HioYLW0RXAB3i2W
esvBm+xcSBA1lb3jSGNc4kmtBPbI5NVkMIHHQ8GvrGsap26fVGGseHD4bGXKQ19g
qAX7oKKGzAv6MiQJULzEK7GxQi40tjuy5NHJOyvPerJTbC83UbfeIddwgPWRpOCR
x23o9FzYynJiAKsLlBy9tyukC2jkVw3kYHF3mZSVoTDmdc9LWCToWlcXoCobi4dQ
6224vt4LhLmd9+gjwP4SSD3juDqsLfv5BkNDUBNVFF1ScAKDg437wFwjJA/skyh1
J/t/x8jx2LXPCpHNqxz95KOpXTy/wNgvbxnxU2M6x6/BUsylYza9jRapqYbNSzAR
tiQErCC30xpS2G1kk7V14LMopErnPwZ6kYl9YcGC8PjWxNC2FFh+e7hUPEPnV9md
nz4C4W+5m8UJmtCCgks/LZNR9F7ck/2GyWxtnFhgN950JVXKGwYYG1QnA8v+7HXQ
wvNiE/tzvlIhge89iMOsPRvLWMvl6/TOcsu47GzSZUUXZZpu3Pqkzms/8Ig25yk3
7I+clEIPMY7TaUhHX7R+5G7OFXUuxFjE0OGPnrFIEArji9fC+KvALU3n6vLl2MAP
VgSebN/5P9A6XX8VRYWI41xlKJ2SVoNZTuKzaBWGLGedcAknEfnsu8Agea9vXSUt
wRWYTSJQ8bKlXvy0G5Ln94B9fgrnwreMwJPPbo8LJoCrG0tBrgMaJy2+BFepOi2O
aJzKH8Qrgcrx0NiH3N+nrVOhJw+iNa+zdzm6XzAF7EIes8T211vybApQlHYMnaGe
hHul+ogg4y6/p2G0OnSCY1i/PoCOUaczyYE68Ji/0DHTYPNv0mkD222kMIeePvUI
1WjoHOWCZh2OyjKGoKrlZ+1AfxbRmZOo10KV7xZsKDDGn9xhAjk+K6uCS94aTSH3
hTG92Tv9t06r9DV8jW1o3QvCZARgGC8SbFgFnGQ/cCAcRDrldMfrpt5gNORDBAJC
BqTI7L0vSVf03SK0YXPD6HCR6eTmZ6ba8obqMR3c+VDFSzsOMK0eMz17/2N3+ePS
LtZccRdDmXBrIQuaQuSGK5sbaXFwsWv7BZWocCUb2luu5zLOabL+e8Sgk9XsXiyp
u64n+Zv2CtcVJ9LAzzFPdTsfhAxK8HJAIQaP/3IGmHFXyEs+tBzTNC4sCdXcUmJ5
j2K23zgtiYdiWDc7OkDaddks0mo9iqvufXsEJFtm2lCJQK5i/cXBDdjKcGPK3P3w
+Qez80WP5VIGkmBPTVfJTc4hxd+OtS2ae6LBPBLfjNdLtNe6WqLo75OTa3WwerRl
wXqTJCsxHA0SGq9LZcQvEcTCUAeCZFw4MGIKqFTLwWeV1XRMPs0eTksp/k5eOhdE
u3O/dv7lyHqa9fPfijN+MHDUxUVyKs6aqj7B9BnQCXJMZqj26VUKwJXZVEA1vfHU
lb3TblqScxfdHe5SlKwoW4/tiZMU1UT8n2SYTKcVw/LKAMFhncyTqdXSc5HPc5il
nYiN5Lmdrtw9ulSg7Na1rqL7q4V1Yv5oKrYwG9C3ZOeuZ8ypSP70fNuOMaUYj+FC
6j39KCVnNyfisSx0x7PY86+olGTEUbH6EoY1vFyMJVRmeWjlsZa5/IzlMQr59FmM
npYGvfIhvCa7ERl7C2dLVi8JLNSEOsiJokB0rwi6bR5d+1kSYyf7oq+yBlYlaRTo
8uHqq0T7uMWDBwGOAV//Tn9C5gshcHggbsUPue6476i3J4Tmhxo8uS6yEFH/DKa/
3FnTsfkoRfVORidRkQQ12GpU4XBh4jN7ImM4T+QwE67iw5Mw3huudZoXpJjPxJ//
kmv8+qN//MFu6dsq4oDESi6rEr5EqkeAv4sfFzNXQRhCD/gYPHFQmzJz7m+fE+ys
lHJaiAs0o3uxsfentSdDZpgrVQm7A/5HpWVoDM9sXDA6dOf3MoKdPbd9GIul6S1N
ZceLHP2ZvYnQjRCMN3vvcDTjbJQbRD+qbtj85ZRODTVksp/YbuADnPRUDBvFaQ0P
1ZvQUDjCS1ImQmgfbu0wJDPA2dWSRwAil8vH4RLSYdT5ZsSbd+NebZ0hLJtYTJsc
KFdW45CzHGSKOONzC3atRtFvBqBEntYGjAYlO1xV9N9oigchkhH/XzoIdhTy5O0X
CKma5TmLYBxuJGg7OvxasAC6dK1O+2cBLkrcz6347MVjeMk9g8m0Z2arX6cQYmkE
1KZOc6KO+FgYJM30esM3NbKyR4uWPOSd0pntaUarj6t+Nw9bh63Gtghcw0JuG/37
n3ZLOJcetXtU1yGpB4ud7dz75J3J6DQr/F1KvjnFwp6wOpf234z4JXHWpB4VX+uj
sDhMcO4tcO55i7taLyls+vM7uYUbaK/s4Ucsv5e0nsmBVTWi1ZE1MGUYkGQ/U5qC
QJOLzgNndg260u+Wr/Djfcebr9TBsrnkxB9S5KBsLOKPSRqQ+HC2WZSmxgaIYAfj
LtxAb15vWQJnY+j9ivY0XUiA7hnMWQRFFRF2wOgPEUJadXaIKVR25CPUWtr38ECV
mBlvRb3cj6vxfQ7Wlbo5nEl3ih09a35tOsoQR+lNikCsK7dhLAOM17WEHllPD44V
GGFdc6/rLf8ZF/PLoknMPtVuVMc9um2uPfPscT2z40YoenAb6V6VYndFksAUlt/V
ocRpnwMscPBd4yRZnvFIkxNNpPUHILtXudy/w0XbzMOui2jz2xYIkAZvrGCJ3Tjw
qq2yHnlChEK5Bhsww4lL86ibec6mTRqVV/6HCZN04vCTeoDi9W816WSp9a9DClBP
0vdQ47gajlEIh7T7HkJ1QoA6yJvhnE/K0/SxqBFrdCAFQv84JZU9VZ0WoJ1UR1mo
ZJ/WsYdfzc0c/A0873NN64Aei8wxZDy6eo/2TpLmbIC7J79F6w68bGsBBul1HZap
FUYyB4p4ITUDucr9/TxoBREzVdjvlcikaN73VjEtDCtJyorK4Mgx4m2OhwFsLShK
TzOa3LoQLBDwMKRoEb61u2kJ2e4G4WU8SMqmiooH99ZkfAoR+vyLinfEfMjkQOLO
i+//jNignNnvkzkXjgVJNXOeAGG7uv5Vs7HbZYR38yZRY61r1cu4BnStWI1zG8zS
bDZHW6b/6ywMhWNsuDuFodzDFrY/jBaVbO3ovPRdUDZ5AjJN+SyspTblTVPKi3F3
5SBRS+lwMYEYArzmo1Zbdddgz3+jn4yEjVYQEcvbhQS9vGObEMor4Miy/yh/174r
XuJvhz9E7Vhs+13kXaJWKZuggDONuafSRevrwrO/sSci+LBO+vZFERrSGy44DKss
KA/798wQxYhT2o8FFE6u1SEGZtOibPPcqr+T61RatY+/WGvxPNMZ+P4rYX0cLimX
oYf8Kx1zhf7c4zS94AVxdrwRALruB7Q8uRq0Vi7k8Xk9CA4Sp6Ci1/txP9vCtuCl
Qdq49whCt3BsM3FqiwUzy1kFSGdYMswznf+3Ecu9rpXyhse8/WZSFfQue9iFgmU3
Rwsu8Z/ZE3omY3Z8TxjFDmxLbjmYm0TwIpZ+fUSVnYCjsW7ljbYOauAUoyK5CbF/
L1LvWG3xCpZtdLCVt1eZPR5G2osF/65hv37suL0Q1CB3Olazi4WxGzT5PFcK3lRN
EoZST10v0WisWg8DNxgq8Akk320PshTEb0fHmg+HqhPprI0wniSVVPPH7JEhsQO2
va56GkIsl6lwz/mSdj8pV3G8k+MdFPJh6xddYinnJn4o+KAx5hAGshc+9TU2h/cs
YecQDE7oSzFap0nr3Iprc5n7rKh3VKbpWigv+4MCqBr+5owCPj9opSWZLde+7QlS
NLApFr1wUUqOmrfXoai/yctNzICUtBavLiEccs/y+97AthVOsUVVMpNuoW7IYPSp
fOMjBZmyhe1mM965vr9fFEp6L/VsZuRXhLN5QmEyUg/8GTQdHtFHcDOph0vGu1ty
RjmvUs2TLJw+gAeWmOkF5e/TNl0lO38Wi+zrGX0zKrzRInW9aSAZZ7Q0IYCuMtZp
7CgqagJQIDy+0Is7pa179Fzg42SqqourZdrPyrxwOd6ZZ80vRImnsHBIe16u0q88
Eq8N+D/Sdm1qokN+j0ALMmlAbwqOg7ngkH4JgyjtYqN9xekYj6ql0iXCOOc4mifv
HV8+mUxMSKeaKin+kfi7L6HyRjBoPc14PGLGuQZd1Kh37lpuyWTsmWKgdmuLmnVv
Pk+e69sqJ3eeA/b755d5133xPG8vXo/Rke8L6+MKYdsKAAiH5emljdErWQ4dJoDe
A0Q83r2gUQjiuf/j09Jvydqj65V/e6grHacLnVgB1MjXlhuXMIvYlFtegcaoG5mY
DG4QSxgyRu1In5doWOC+tdw3xzt04U9XgFj0w/NSwgXIJH3ZSv/EIPwDJdbRkCAf
/LQ+25CTtuRKmA4NaxDJUR4qTha+JcVi8h0xnYHe69A694aQQA6B4FJJGSD9/uAP
5MBqFlEdP3SPYlfmdFZeGMdbLUvv2gGJGJ4lLt24qFldy1x3v0aH7vRniGvTr0DH
nka9r3PqYXJJANwQF+x2De7gIpd3fOCCy+f8IgMpGoWXIsYPHbZhilsNpB1ZoaZG
3oA7x5N0iNSbBZVgR4mm+3wGvKFOZs180gzgpOV0/x8pXiHEnYaC6MLWaoUVLdKI
pAMsI5bbYE9fF2YJPnGmSo9MdrwKMLLxhCW5jqwtTkmd+4+GDbnMWcq14qiAHPc5
fenK+vsSqDC/nsrD/tUHwbUwPoqZj3zXBd/7AlEC11k0kuBMU28BlDZihBAs/pEB
IesHSqxMzJK7tGoHuoLMnQCPycVtwwncQ6v6CTFh1X38MpeK35p3ETo+szgmWiIf
kxfDCF0HrMjcsdjjvlBHEN36YHPyyaMXcHYTgW4XwR9Wz58dLDGi65Jn04tiSMbj
aFQXwOLxpegXw5mI1Iev+NAyroEVoXTlGnfv2DiOxcH7+T5EhEV1yoPLmUVfJ82t
RSsV2143DmQuvgxSuDncoq/m/aF5lG329U0tcP7YaTEQ3hnjQ5sJ7UBgXoEcm+w7
/DGE9wl/o9kUgNs7po8f2fKZw+GToBroFNshb9YiETH8WNOoUIwZqxv0EqkoKMoF
9NgK9LRtjGBrdURxYLieaNRdFfuDW7glcadh5SIWnZziaYr1JiUreZ3R1inRTrsr
GlNQgV64LCfWGAZXjmYnEwOuBAmwHHTgHvumx+dbSA3z1dHLZFghWU9YepUc5iDg
E60oQYvjkYm9bTwvrpQ8LW9Pw1YJPZz68bVP+iBb6m0cvKSA5t6fjdHIrctrvkFy
kWhTcNtNkqaRHA8DUzAZd9iecBXfzcsYJV3KM061HxTL6un8yCCbQOG3vJ4DAmQA
fFIQhJAwXX/qsMTTDFawP2RlysOMTsJPBTpFoFIruiopbDRRIarBls3GF894f18K
wLEmVw32TbbgBWQm/r48/bwccJxQbx2vx/BXakcOnzLRijcv6+Lxp5p43ER/OpQH
xynul24xG1XVldZ/wmZLJws0WIKO4t+qxPRR+kFrTDqmj7/MaseGngVSJv2H0Nxo
oOh3dIbKojK0cholup3oY1jv35amY/90NkhQtgpN8EJiednxS8fLDYjEmxvqZGae
6cCe0Qzpqg1r62jObtBsKD0netLD+c2eDto82+g4yy3VSdkB4RaHw2mby6prNeGY
RPbAzobsxfCbTe4mNQgFaQ8P350gxXfZ3Fdk1d82HtXXRa3LZ8Fwwp3NjHRS/q6v
u5O3pgPe16t2ArXblSsVQQFnI4E9JI/iLE+PxmuFNgStRAJWNmiGma23Gxe4ONsv
ggXzHCEV1usCSc4+RUjeiyPc1Et30UsnecxVv45S9P2b9y8E6/Wx3/fZ8wRIf1Cj
2JuVIdQZFg9Tx1HY3WaE45EVIv/m+zC+8tryfCwgMHAcvDllGM+n22vwbSeTokNs
VnujUNdnRWfAPUuLIuLOsMFrE+nJQRBDsNOEgzL2HnfvQQZeOR3F5wn6hkb5Tvh7
WWlB6YsBxuM21EbF/a/aFc8+kBPwBQwmKBwsQTGHkvXTo5IXAoGanl+LU2NblvvS
L2WWrmOhi6MzsTCXsKkShABNpHZ/MIqRHoKk3siBskTscRJJKT/q1P8Uv+8Mp6ku
be5KpPiiGu/gZhZLdnZvuREABKZC15GJSHgDoyOY6LPBn+H5GCV3+7DA6xfWBygv
pv5okAbjWkrZGbbKIHRn1ypjRebFV6nB6nt/kymdUhWNkF4q8vQFyi21L5LTD0Ua
BjCCR2G4QimR0+iSB/Je1x8GqpsMNofrjPT+hYw9wR3MxP22UMTXhxHqnCOD/OxP
h9A8HN7sZpGizDsy75tUa51ketLvZ+L2L+9Ay2Wi2A+BT5m4MD1GoaCcT22uA2FS
5bLhWOZdYmXpz5HTL/42FB5bKpEq3NhIZRDt2YgNhkbiNIGD64FVG9DgWs5eEKN8
KubgZJS6Cj9UHAIhZiG/K5isqk4JJy4y2XrkV0AmMDOIr/CQAcKe+bWQ8OfJWBy5
JKkPxhJMnY72AZLfqS0jzaziqvSd5+uqTk60R1nMixquevsFsPbhmOSjvmF4KKcx
/+2zcRYcO/LXdetEe07+5hJ6vaFrWxccyjG0eQsMCXhopvQ/4cDJ1CU+V7NTQq39
XMDww/If4NbLKqKOualoT/dNDl2iUWrxTpvPLk7UzsescfBjm/AKE3ci41tD/C7v
3Afb1bNkQIWtyhr3XKEymX/RZXIe58ub35Ap8bsa2oA7rGfvdwqthwlCSdo05xpL
A/HdnxSHdwvbDtvnNEEFZ/aiomPEJ5OFovEO+8khBn88+NIwDB2PzGT6RUYtpC7V
A1nc9G7qwztx54AM3g1pQhPyiwUdW9G6W/EuZLolYKQJuL+vpghM6UjM3u8pzxNz
VSGNu83INrIZJNVRdgdpqz7386m/pI4ql2cVVc4FWWOmZ7cuyfYjUmBQwLHxfQ/3
/h7ty8vJF6BIhj+ZLVkTgG7DUu+ybtO/JeDHrIcxTxWcZtBL+3W31x68lr5yNuAh
QsuvuiaPvDw0DY0ad1vTApGNle6NJVTX09wylOGnDDPsHHUaAzF/3f6SPqe6365d
GNL/7QN0rGGlm37eRSXL700UDzvNGwggAcjsKMfbMkA4kM3u/i/g1OfKAj1hXWVJ
ZzqYS6qjbousncIJPLb4w5DHXG3ebotyazjEc3xR8jQBxgXm80NWY2oF4w+7JeY0
Zl4A6+KprvZp9RmN7GdgaoiB0PvSqo//C0JfyWBmEt2MbHQ0J/EoSZDEG/xodVu2
b7DS4vvFyNzBt6g/QL8l6x366r+tgOnH3LhTr5GS4HdH46+z8NpoS5JPSIdjpG1w
t0+Za59igqMNosPHhVKQRYtNR1gjKDq6KVwVeA6JURKGmq8BKsdpStyTLtqhE4lN
/jdU26Pd/CxIxUsUGS8cihKJHZML6nfvMY3sLIwfyINotAUMvpKt7TX7hJr+H190
dMQu65LvUbK695WBqjeo3fE90KGYVFvbznrhJhHv30m+VlEy14H5Mf8Ufw2dQhuC
LCPAnRg4CtXBWOH+ky64noIaEjp214Zmx3iVxYUzBRDbU1XkO0505osI7K9SkeT/
PCeB7ySL8ZApVxqchVPCOQdIlaYoZu8VXOv042Yv1vtFE0CFrSy6yvXVZN8wYAiZ
cNfaqWbbcUDeaHppqpvKDNzer4tCdDFIIg/MdpS1yw64TPB+7ebBxPai7+19uvdA
KeZLx4v3gnQvnzCsdbQZj3i7w8TtgGqikUhsbIk6p+jEA6ZbPRMeWkhGa8mua6jl
QbWQnkVpC8wGoQnP9fKCasNqez5UZm6j6bFlLNXyC4WjkRmbmIdOeN3KWbHjyBfQ
+MTkuhoH4yms6fmnhX1NUE3y9LJAUrvsiL/75wH3Ge13yKN3j7PtHagYwAJQO0bG
gOSAWxPp8gfMjJbd1TODtfmAfo3fS1qPZguQeJgIPP45OYOLlZlJKC8Kjq1aRRvZ
ys3ijoLLCbp5YAs/mn4rE3a3M38TeiYb2DN6oKS/8Z/CUoHH9TzbhcK5kc/HGDXC
rUvTF6hNJbdrioX3lZmBrGZYZ4nO/5gAWgyrNBx8P6oUExBuK8HrAWatul/RGrxT
j87lKn4kvVvpNK+AZ4Q8gujPktF9SyBjfrl2GJMEyalGU1Sy2TCyCB09iaeAeeXp
HC5MCWGyd0wc6TAibGS8SPpgAwbXR2q9V9K5bZ36Q7EQiDdDbH1/bKnkwOSH+OJu
wjT7TFYGOy8vzH6MVzKLW/+LPHVS5iLHbX9yYPtCajtMSAvMvUhrnDvKj8ZTRhDu
Q3zMlegWV3cL3XalzAGtIG88D3qZ5+apPmhdrd7pTEmQbiuLTFC3db8vJFf0jOUZ
NgNZtn+T/RAfaoGt5YkYePNHEz2gBzclhiUNjx50vA3PfZlsk3Hq47JCvXHdazM2
c2FIMIGR03RnPYeJ9uOyglRigQqYEiKSX4WBVOTYFF+JcbouIv5kJolPGESFIDki
4ekoDyHQ2Etjky/n6HF4LRoThmZgxsGa3VBPMyeJFfV/Lmovl5xvdbnuuqXbCuhE
H88NfEG7KzkEL+AcoUEd1ZQoPVbuV3ChTmN1TnqGe2w/Io5URfrrgCm9KAPX1J2G
RAN27mTy4rCkkJFbECsFIPHT8g8x4TxdMBAMOVpsWSpxRM6eSrB+QIOZz5gWysEB
6im7r8gnT9MtwLuvslyd/8lNr7/BJZSDyBgXM65vFVdnLUxb6ZQkRa/p/r5jPjPQ
SSC5WvvtWLCkp8e6e120XLmLaQEtPHVETKWIgFErAjzk2lcp4wOMucXEUrTL+BZd
h9Tx95cFKMb5++c3sKq/gKCF1fgGE11KUJ5y149CcKAUo69YeR5YwXoN8c9ssurW
7zJL4SZP18c0aESA2Y8zLcsEYu4mKeDGbr60k5F6r/AwX1SfEzfpAFCMJlVVnl1A
CAqKj1LVMWU5g8JVWE3ijbRJ23rpOhhtFxwN9BZPeswhH4V8mrUSf73wNSjSz9vS
5Wrv2jBNU6kFB2ccOv51zsP/GS84Sx6WY3FKF9dGrCluDB3/R7ZSFi+bs+XaoIC1
zQ4s1zuSmjPq0s4veXByDb/F07+J7HfzzmZRReZD2S+dz9j2+7mlL69ugb7R7+aK
4IPXVp9SVhHaHm06WaQ4R6oEt589LsPx938m9mY818bHPxPYtHIpHBuLXOise1gJ
XvVl/VlxMIivhRg+mx6NOQhM4BkfgFAyql2wLIIxTosmkkXet3PIewWg9QY3nbE6
IHvbQTu1l2OfvCIir0dtFtXZmoA0oVsZ+EyfKT1Fjmc2qSHWCarK0CGstfQDTBQo
HOmod/jR88tuBETKLOmMgLWIiGsK6sBwbR4fDzFUJI4wj9YbWZexFBEeg2m5KbeF
E4LPvhZdD1MfAX0Kd0b6cXIoKBgguSsE9AZH0fVnm/UaCfvtDNiWwxouRIjZLSEb
mlGXwBYfRz/kdmytwZBo6yskrwPfJGTOj3gsbhpXWrX5LGBV1Yoe+BruXva21dba
ke4Lq6tx0SozxiYgtbOtABtKdEVZBdxPXq49TPNrTaphR1zWJd4JLDtDwpC8SEd+
c8JVfXSSH58RVcwncfmH1PQwHBD7P372R2+ZeDuMRMq6fnWn5RIkQIiPrBiVMcFa
YPFuEfV6gH+HBH1SThgM+4GUDgS4m/2GlvVmkDGcEvnhkCHXAeBmXpdI3IpNzA/Z
MVBICf5QTc0KcryNyMCIGvUtd/g5AAvZJlagIoPNUN/ADm7SQkB04rH0EOHmiDEd
V0SUnJgbSsp2XZ25snaNj317spQcCndImZk5WwD4Zb6RPcsztdyrT/Yo4I7DMPr7
PuxTMQYJH3lzCsD0mlZRurBjPw18Fe06ySpAbjdSaV26tmEeIFIZWddjaAS6IB5e
jcuZAwWl4+90RKtpYulu2yY9m+3W7DIoW/iHXw3c/HXEttXB6RP2KcaSUJNC2EiA
hyMx6EJrtGPVgxXDCCWxuoXpQ4PQzObIJv4Sd1TiXCix4bE1TQBWslEufviCii0+
YPVpEpReLnQ1d52I73DBpcSBDJ4UR90eBxe1XNraNIGvBOO+vfsRrrcaxcsIqUTM
XX3cQXcTBtD6uqDOLonFIa2hcKGXSWaEVQCAZw1pHf/jMwXvcdgnn/r2T8HLM+9m
iClYUoaQkr3Dg+sxTnCyaCPFjCRY+Py8OxZxN9sd0jemFFt6LZtOMr+NOo67ROaL
Ex66/9Fv3qumcsCi00uU01RzrGM6pvkddOC2Kq/FAoSZu160T+A7FdG/ZMOBlAGN
apkGQWpLu+fznpzWQoKQWTWYQx9k/Z8KVdMhhTelaIcjV8hiHNWm5TGar+o0NPgx
+sCuqWc7O/0lo9IpKTyGsi3ku42YJCRnTN6Hcaz++DqRoYVRr3BDT3vh5yNeEXt+
UyOIP7Y2PCRmHumh1YtR52ns8C2LmFGgj9hKnSwdgz1d8li+/Zkcr8FDU/TbPhKU
XS2g5ZRamO0Et5ZIlZOCXMqDsWHm53iCYhZytW1h3UCJ5iTDpj6GjzQr+pAxRVgb
fCUmO9LPQ2ML3Z2NTV1CRx4nJiFrxmN1svueC3wSF5u9kVxXMxWKInabc5bVj3Ye
RblLn+Elaqru2L6Okm0xlNLbTX7zXlCVCKvvPfI72/fKTUwWX1iGEuLDA+5Ga+N6
5b6qwGXFIgJeg6qmADPapqAnmFw6JwHa8ppbw3J7VoWerrp34zYt/1yu7YoSTgdU
j8YDYvzk+IvqIE12q7cIxSvemc4WywdXTOuhmYx0S0QjNeV0SHgYhCo6MUfVRu+n
/AuIZwltA2MbVEM2FeLPJMUCss+eZ4HRIM4jyhzQqAE2tdJo4ZTEoY7nQAnLdEeB
vr4yiCjTEtCHP2WAbT44G9OxQNO6vIG5sUoslF0oRqGSxz/E8nPY4W5BwC2lejz5
IZUjZfejx6IS644Fe+KMtTqR6eHaWmwnXnhy1w5KoFjRS+Ro4rgivzX1Lv7LmHZN
upzOgAQ1ru0rpiFCe5aEKJY5rustNQkzCujQbQsC0xqytenPIlVGwf5AvkVtchWK
6mMRAcbMO4IsB5JkukXavdFpHt2n2Yy47HyR0uF/qkTtx4Z1qwrpsEu5j8Uk0LuA
An/iIv9tMbW8UqK8v4cnnxvs6jttA4gb+EIyAwkFlkf5VSFy/vWUendWahbJZVEx
A27bjq/9+Xxf8T5u58LZzDOOp/rOqXAi3sjQipqzr0YnR8cokwcEQkfLqaCCvXGt
IP/Nb4+2wuYU5x8fpMj/seRPABtQCIEU6bqZkgLTLD8V/TemJP1R4h1GokYfzOpj
1FrXMQrrEHp2MNYMjc0R1GD5MJESVbilFPdMSjZ7M0lFz2K3PrB/VEa7LKayRhoM
Y1N4TbmnBetX+bSevFvu+Y0XVZXgiwb2Tv/2sq/rgaiVzZTck0cDfHU366ViWn2R
VheB10WUt5+Toi7NGtU+1m64Q6yTzrgV96n1//YfL9Q6OObeuQlSAoEVxJPGK6hK
WBTIcP3QzpUWGyJOZB3+biGUTcoodPe2KZbV6E11QSy+kQTEW5ZNHynH3QjLqNaX
YJtwVXO8vjWtGc/MaXLH6WD+vw7vy6zJVGMOvF3ta/uzsuhFnON4gnMq8KQRdjZL
KstuEPe7QKYJExyx2j8YkiODbWFtPYFqhuby4WEXsnDm6OF/SnQMO9saDG7U1fvO
kR47LmRzSTp5xYZmlpVph4lxEpf5N1H2hV2iW31XoeVlF5vqTh68JnMkUnuUISxi
Qr/CwFRR7PaRJyzGGAMjkqRnEoZWy00HXOxJueFzEL0iWusGjDINR3rYIZIvM4GO
GKcJ3bbGOmihu6/RKxlBqALWd6+jnZqB4QDVA/ZJqH+UQO5+ucGNEJphck/CkFOt
t+ZA3qy0CKoukakay2eerLb5eUmOlti0V2mc6l5SgOZNw59OMdBuY6pYDCFHgiS4
GxuY8dDISAj0J5G9QjMZI8mVF2Ywq+HlA7+x4rF2GHOIvKFFG3opBJq3Ta21VNWU
XO6KtuLv5nfkrdn1ZkNxRKG5yeK2ef+W+HlcdRuxTJuN/1L0wPou3Z5ioX9LlXTl
C7H9zy7uls/Oh2RyUZPvH+MByWHiKIu7UbHnkGKFH1VQJGnBATNiX49Q/s7U13m4
HNJ1QcRCnPEGHhz7Ez7CKKAG4Daq4+vpR+n5XOlXxwhHvnwUDHiF4WLXuKrxLZFu
Y1G8pJkPyiOzz1fRLRSDu4OBiLN8msrzhU8yJT3d3lUl2IsZsjShEyutSsfJD4ae
+6hb/PQ4sd+Ye1wrmFSNZhb1K+YjBwHeCqxZtx0GgzXPup1ScOAtuCWc4y5y+NLB
8azmtoqMopv0Y1osSiDVrGNQCOGvQRR1k02y8ipJDCw3yVLhY3lVAw+lVPe2xcgT
nFaYq2PE5gHo2BbML/yme0NEOKOCMKvvZ4rdkjyUlc85jEx26U0V/6ZsBmqgTgTX
kgynLbr7fwwBt70RwlCBc3dZDAHmR4386E+07IZnFsspECUoovjFRX5JKtBD7WRO
/e74tkgosCwGw1E77/O+GB3lIIQcfDi4zRO81vxEQW/nf1DUUoaYuXEyNMdLVm6V
fTnwrnRDrFgPkIkRfLSc4LuO/+fGoZmX6sTZn+upfspt4mHML02JzGEgFu0L2KYs
PzjWbeBiMj/1blM0IydP17W6yhJ1uAHAYPmr6V8OQyCXjUUu2Z2F2VefOWr7Vocz
0vfkM8hBfNC7hspLZrvPyau31SvAjfy227102UaiECNAPZgZEGu7ak8GPbTpV66N
W3E0/c0dr9gv22ePy0jTfM7iUKbkt5v9OVyv8zgrXPeIH8QmtSu9gwgkb0qUgaJw
gFV1GIz850qouhQE3PviG+4f60GNiQk3oU2XxTrGYZTm4gSrkRjOBAK7GNrk2vdE
hesZIV/B0I6iP1wfLP8S04oduWWmFZijCYgoJFuhxGve4SbNNmIMynDDx1okZmkg
6sptEYhBjh7NG+v2nLafUTvpcFcAkpHnCUdlFC8L2uzwM6GOzlwfbT2aYMMvmJWm
mvrV2++kgLbBn+1akwiYIItymS9ihAK2daV5xzHarsSMpxrTDGsV2YZtXUa+KLiq
Jrfht2t2miGkp+TvetSy3pOX6NGcq4qW5f3NWvtAcQPk0rUYEunbybKPqAiYOsts
p7TjsvOQvZ9gINySqcTFtOlO0iytBtssEkpGrCngC0hLCv1LqgZJ7YhnI6Bng1Dy
hNkjym7xfzFkmgwQkwkRQU1DbxHQf2nrVE3u4GPNy5rGDCxD8UkcKLHnxRcC1nNk
ql3Mb9EttdL5M1FB+M4hvcGby7W42bJn1yWGvhrkXOuaaj5GPNFhP3yurplJNnll
445MGR9Dv25VDyY6gQH43tUnsZlbmBHWpu+WHeRy+yBRJlMijTfdWSTvY+faiiCw
9szd6cr3VfAoP4rvifpIaqL21c+M03FdlkyLcmP/DfFYQn2kJKjS85jHEBYSifmV
C4aXQNEuurbC+p02Ihhp7jbLbbgYmflZ6CuaKy67pYe1hPVjRYGi3SAKP86Myf0l
m4y+9Zesi/fY2vmerWdEweUjGeKkY0n3/QoZem2HZHhnLHe9qOn8xYzZPQeuOGLC
/FSDnZ4xrGLClYdl1zM+4SFcP3auW3XrvfhWTzfk3TI8ZgTV/vYy5PFFvpVCW+We
gvtw6WlyFldRXewk4YqMnGY71B31jlpRH51t+qj4djrfYQYLcW9WXu4R9CF5x9wX
PEbGNOgJT05fG4LV1lmBvABr/CmuWdBKMgZD4ENwbN2gMgb8rCMwzJG8NZjHcyRj
eh/moz0tBzyEpJvd2zK+qaH1VAJdkhgE4IaRHgbo7arcK1EeSoa4MzOJT/KlKQcJ
ndUqP3iX5kh5i9WcymhqKB1QRvHdSs2FyC3gI7H9wwonJTENiGvevMCxvqniNmUp
4xIMCueijJ3k67cR7X2DKlTSpqLrxdWuMKE81gIdtl3RvKtgdbL0bcmnRAdv4sPg
keQJFzfpCHQEukAZMpD2yJ6k3iZxiZ8BRi2Ihi/KV2QMNSN1LUhGcDQWqKsHb5jd
5yTOwJEaifYrNO9/LzXjiqQTTxlVQZNABkO3javU9KYT4rXtfhNQV2XewxWGJ29Q
JgiJKp1gzY2PjE+vAQ9ve+3sHFDqWCtxkwF6vTO6609G9jUVievlOSHTq9KnCxF4
tc+86wsz4X2MBLVsh9YMIvE8+xNa38jMVirSlNXZIGQh0l7qyaYPreHoBnXQ0FRK
asIdxECR1ljJv8R2Q68V50SvFroZmV7Rqq3JOq4w/W01XeTkLHq/1CCljr3hB6kL
Oui+y9rUEUBGYWC1DzlW9Cg04HzjHfEeTYsffV3SWDeqqba3sKl+g1fbH5xKPWyM
YozljHhrUNgBejc2onUnoi/WIoZhfeFAj9h0VgX22LmpNhxX0wcmxV75mCB4245J
3EJsSJVUmBOFb0OvRR+pOP8oVWBa2Op/379iJBEa7SpHNBCeh38gJl7DJXo41nUl
J8P5st/lFTIkiOVXbXFVMLButPF2iZefeiOHvOB7I0Cp2GJZT27orwcvZ2rNx8Bj
1iA6vcm6e7uCAnlIW+J971ShvzPNedFyMq+x+AeLcnZ4egmmBMW/6zlAzbbf4P1Z
QgoE9+5L5irNUuOyOEpPSN5I+bFK+W3xP12dCTqSc5t+U3a05hITqp9zek17KG2J
KhvVUTbVT80PH4g0nvZQcFdm2RvSSdiYNuL5bVNwRwMKLBFWJKZPA/xo/xGk8wl2
XQWKKZzKMHmudDFTRosmo3zzwu/7P0BnqnzHoIaal3nz+8fr59jihYmJVW1dwIsD
7A1MYMbdpTx6R0XGvshBKNd+iJyuPQ2SN6AcBT/sa1mc6e0b4njXwyDf3ehuMSPp
FwZAEvIb/XXBVWKzbCC4aY8i58ZvgblxdKGWd9EWS7iAUwoyNTt8A0L1VMHnNb3/
4VDgkd4BIEgHvRxwEmc7eHQ1LiD8j3LyzZg8jKdqWrh7pwBm/LYqUAx3cFdw1pQP
aEq5mUrsfhigFlonjxgjWnoA7PfW5QLlEJki5aWGEBrlaIUrNS2phOxRxkFsuHp/
r9mIPnAKKPVb5D2ZRB0cUPDRYxtKGjoKjCR6UDzIkMS5QGlyG1Bhz1jSszyvTjV4
FI2R9hnw+aTl43ONUKZwV86dLOSQiho0GvZqJc6eouYzppRPo9mv+zbJQPn2ARpx
QfMjc0uv0k5diPfyKxsESXxXs15c8iw7lITcbPjXBFWK8URfhf1oEcXVBT2OMPyI
vAvT+yQCsv3kVHvvSajtNDywcZs0xNYsamkUwO4nCvFtf5mrTEmFAcv+0dd2aaC0
Oug4UWt7zOVV1/vyhgiCas6PWXNB5UdLHFQowEdaOkbqinHy0waUafmYwdQWf9Da
T3b7urWSsJANbviX0+Iwf/gT3SRJUP+BM7vruJkOOJHLpSdchgiBg/25VU6DkHHc
AU5WcfIVBrW0XsuR3EgvWygq+o6AK0RkNEvGFsxveVYpBM6fRuNKnRPnE2kFIUC+
N+EWAF1MKDn3jRbMA2XsfqkwKgK4nsiHR333NkQqzbNR94RYV2/fV8wrLedaHkRE
xPcM8jseHTjkBhxA6Z+WwFOIrgtV4RAzuib43dG19oEvUaep75VajPdKU2G/u0m+
ZXQfTjKMAk5iCyahRb8/OkAFT9Bp7BzFKsD4JkqhvC08VKBtI9qKoWlTcbdO5q4n
irShOy1sy7fDodPZ0Wvr+buyLEVX7JBohALyTgnIvKoKqBdaKPGuqxB5hF6eOVT5
nfapg9a7QNRwXVje2YjTpoudF+bflr9gpoNuY0LPqQLTVn+fXkGJzdlg/CEjXNtv
A4iNTtziFScYsB9TU4Fyvhvgk3JPHXw9AU2IdpTy24qYi4jyWYjATLsyABZRkBw5
CAqTKiGKC0vto2bW1xx/58RhGD+0g6ORScSQBcI5BLDDf+GaF+1HXD9WpUth6LX5
folZ3/Cj+cP9sP6KuZjRgn/OypuwmBvJSHOPRwadjP0Z7ijw/Mg1mDF2w7U0in7b
nuMSEExOI9Vj8hOCJkZNowBjpkZ6s7sthhcnwEJIIeS8jhIu1TImAzdc3sajGCjP
df+gq1JM+O6eA6F7zNdqO+xYvHQ+6HoMBJ33/y1KJC4j7H/IDoKoooFkXPmWLkHQ
6Ux9tQ7lXPC85TAO03+C2J44jBq0j2wG/aVJEVqkKqik6acnK4ApHvrNYOoA+VE2
7YA5ZCd6UWSl3sqS1rXP7LKCLyBKnZacuk9bqWbCDb2aso6jk1JkyRY56f7Z5r04
pvcxNzYqITPVRa+xUoX5qAJrPFR5ZdcRxq1F1UUSNOfHCTuxpzLdxu7OzkYmbjxU
YXw/bBCfjfwifXPm/1tP2c4bheFK/qnnb9DZAQGqtydYL7LiyOQDW/vEq8KxOczw
Vtd4djNphxz/qXUlIg5N3mgg6Fe2y7z4N4d8ZKupHbE411xUo1/d0Y6w4s7r8OZ1
6FIWhkzarbiUl2HC5wRGWxA9ECqXU/OAu1xoE7CGp44mYc0gz9ZPilCyEKwaBJfe
yiOE84hnYDmeXoEAY+ma+UpCUj6MSk5us1lh+UAqu8AV70sJftMpxVsn67CaaspC
zui7IpHIVOVqQCIZHMoPIIXmyqP9b/rLwafXU356m7J2b0G2qoYQ9De2vxK0VyBW
xs90Ade3O7NuVDPHthS1e471dnYXplhQAFu5mezOTINjmV+ZnfKMooyJkmZ3oB4K
Lg2oYLc4mpJwBXNeNgs6tQufk4Qc3jsoKgCulPhqZj7kgCJ9WXUT8JpZ9/0HSCZV
oCyAx8caTcRuoqcR1umu5fTDAZtBTDDE1fAkWVpWoNM3Yd3M0SAFEWxa532EU3Mv
ipkGjppk0r+p/0DxJji9EUR1SazjxCgwxTWjB7LISCSR8dv0w7UadCbhwDpX9cBS
EhZz6l8PeLkAeitf70O9hzejl8VygFvAy0Umc7bSDb0/f2bZzPeCu/Mrz/nj1WpM
zHhoVAR6AD955an8Ori4M1PnqrgWNBD+vgAg80ZfINSgRC/ETz8RuGzol/zAR086
yaJNrYlV+dVyiAK1pgcPwD0jAex1jI761rCmSSL5lwQjYMvybC8TzjekhV1i4Wcv
a6k3IUO8xRGBYv3kP6lhJ7MnGVuIKAbU/pOmaVaR3vi9k21JSRS6CxSDofHuAmD5
07Q357kH+WdPnSc9FdfbJZrnFKFGAMupkgjJ9kdS3NXcEuIhlWVIByi9QC70OsTN
GaDfKj5HISQRUA2KYk4NKoPM4fk7gsRHo12d7wEDAeI6uWSlRoDJLwMcDA29gAKn
XjwCxphIH14/+9GUl65Rp77Cqpx0Rs8tPo8UrMuX4WDY9y9uXzTplZxmKLraxV8+
abdWnuRMFv4aOoHGsEvi/8A0oHGm0v9H8+OC0pv36MSNaz9LOD63Vj2MbSBETL1I
4L5PW4QG6MQkxyy4MqUnupbtv1LhCjK7/3aHHQyPRYy2pXbE0fHfHsgRIiAopcy0
sZV72NLe1fYJTAqefF3WYgvUV1S3KhZ9EMeubxSQJ2HBneerLqaVlYmQAvCo0ly5
sK/IIdC2pXWSY9vGW3fDZe2TNJ7ZfEz5GsKJwCPSabrfrEzcKZVYjCnmM+k+W+rb
iN2nJn4Dogncm3tFg1VNB0jOh4xz1YvOgVKM1a77Gur9sEThYwV8w8nmuXc6o65B
ka5M61jnnoY3G8Xk9m3i56btGlcAyyR+N1kGJ4hCMtj0lyVyt4fu4rtPPS9iKBzK
Lc/KTs7ov+NZocsImSfJ12VkYnfhklY1gmGaXdSafqgSj3mO+gnng+Bl60qXNwzj
6bqy/PpZ0J2KvJwRULf6U8yRjdw289q3XBfFH0iHqL5zPzl26nq+CQ0ndiKzJcMY
qzNCOyl5hxo41cVP1ZoFrcZo6C6+wTcRpP652E+e39MmC2XHrCOjgBFSMpWR7m6y
wOOIbI3aRkqkNsq9uamJRmAeyG27g+2xsO9iHD1sjeVxoIjI0rCqNUXPIuG+F8Yu
5CFAutLEAt/J1ifg4Lexq9mVnkkKoJM8Rrkoqxr1t2PDQ08nuxQfrz69Dz1Os0M1
nhdq4UC0YyXnFu67GnKxou6v2yE6rLPjbPBzvq98gutGkc28rMULNvfASuBm5Bi7
TBfQuWZUc7IbYJ9t9Y4k64zqqmqu2b973npMMyU/vKswIG1CUdJL4N9cczZlVXak
dO+SpWeVfmDS1NhAde95lrQ2Mzar87uEtGX2aTXItenuAGTi3hgRVaU2KzKkEgIe
yLbQ4fw9FWGaGYPVpTQ+29zRDJvyG9oB4ip25f181OgxuG9BGFL182YKr33MlrNw
wDmKwDOyhzae2gxB7n5keL+YSi9HQh86qVFl/C6JD9Q1eVS12+zZIfdo4QktszLu
TAaLZ23FVNUHZXSVtbtpJ98mspno1WDvUWN7GNfg9vWm5ztaQ9k7v60/Tbh2WELp
tScKwnRnCIKX9dgdCPNgRvUYnvF14oKb45lsILAWI0mFjhq/px8gmNuIfJvAZpXt
U1pfDKyRvHu/P660OFC+tbrvVEo0OmMqF/aCLtK1vgvyLx1S6vftLzGp70U7JdpD
IdB+ofUvV0LYbY8FN8i83zbwvVba9vQE0hWJyy9rpjFaqOizw27tPactTb8VLSlF
5l9rIqw+s1E3n3xjWGsTNAaFoaapa/yHVKx1s6MbZSUpskDPkqXvPbjjDX1ZKBUK
RWWy54eGH3fDuTrB3bcXy2NfBvioT8uBl5tLIdAeuWcFomdycbQ5OMdZ+b+cypuA
aP0gYtamK/N2pgvBVTyq09FKRNLz0JMOivzOKZfMtregvntD2XCLjDK7ZwUMIUFE
5nJCJJz0bHaJbA2EcMODModyLrg2Q7sADZPNxUxna2e4FAcrN5o6kLsSSz9rQ1gU
KVkNExf43LFGhQIxNC6gbdQNSF+mioaZKWIwmq7vi0KdSYetw1fKUUADvGetGi/B
CS6+CDDbfkZFNWLWsrukhK386+CxXkRog7vyl3w7G149J5xvHzN3Dwl7yEOOa37C
RxmoUU+ic35jx7tg+NLylQ5NCSsWtgSpxMdNAf5lvFeQ3xzdgKYvwIj1K32JaQce
JODS3Q95n2ttZ4VhrxgDFIBueTSK5XUDGv7DpK1SKxyDTGV31GwZ+BWYa58I1UM9
LrkA2pgnSXyea5vAKL0PvXMUdPBPKGrgfJmHYk4FNM2RMA7YTo2A8ioqkAHIBNp5
Wdl5yWrGkAgms9WyTJF3gzacvdwApcXLw3PBNFUXsdMKOktVezvB2zQoqy87+eJD
apjapNPXhhV1XUO+3+xbv3JgEPGKytfOq42bTUx4I/UkqbNpbRkEMwu9f60a0iom
d75rYKdcwBy9U8+uTMzDPgXoLNihmloW8j6YHQ2Ba3cwOnbBjaK4ey6lqYpfILOo
6bWo0vWZdFCe6oVbe3OjMiRSZSQbLP3k2f7wDWRAvesZI1AvtF2Lz34JYS+ku8yE
nPTgJCiMaSmkiDBhXKpbBnrzR5PlrTgBzdvWrg9lIMwO317OrGYDG4r6nj2rg5QX
Ahcq/rkB8JEJklHcarZCx2r+oQvdw8Vkf0Nl1Vk8ktWK8G58zlrIV1OdJHhT/8oN
3kHA7YNN8AOnZX8y8is5pmdoDnpKqlsfnw5jkKnmnG9l5BaVxoeZEPT2Q7MHwfIU
uxlbx9oG1nJ8BaW9BP0XfnkN4pmN1k3uQdOzZfM3lwrxyxUvGCM52E/ZN+t4aG6D
6XACEZwCf8uRcfp6NeFZ0UUYd0QMysLYXjUD/7akScpoX+fVX73M9F2hnBeaKMhX
ePlHVJnwtzpRaM/LcMuSNffLxombSFJUOufjciLYN7ITVnGNWlr/X9sdOs22rlhR
rcmczHt+xG0SptYMMC/7gCWMson61+s8KetlVY7RkzXIibx5UvvkLEJI+F+sA5dp
+hUZo6krT8MIMC/GhJQAAHOYzlCkFfdmoN5X/oA249gOgdpVM022iaPbFZxtX7cf
cgdvC2zi1JfUTr/iSH5MyD/SyiHfazLdOcmdOvnKXYFlg6vqoro3eOEOVCXPGIZg
Mh0LxFYg36IV8ZTCicAw1d2W4zPj1fH8weTO1tkIL3Pkc9+UMat30qIIvAgpuqQ1
oF882SdH6wmNNUPE5ROjq8q5/Oi239U/jMMxFIg4ikqwG0z3d2Kcp1cV0DpJPRtV
JwUHjWaaaqazRQtDvGG7WVg+QEwBocb+WaBgpzVHwwZ7EylcQjNa3PFEbCWmdoam
fONrbF8LiQM2NdpnUaMc1ougm3ZmP9q9cdPR+kZ7ELcIkuzz0VBUjXG6csXNc+cO
fP+YCmgaMIraIOLABFn+sUKAAb2Yw0U/HGp+CnS1h9v46GLGrrIGHF5fRQIpJ/Lk
SsE3JIanICOxnylnEUaVsM3GtvPHEVHxsK6TE2e2nFjHs+bn2bMFfaPvbAsKHKv6
Nl7CEM5TpT7xLscjIm4MWi7lTW5NjDDkyQ2IzGTZ47YdvQYAURCJg4hzL6C5KdDg
MJbzHRpElgcmwCn1k11eYOLdl4SKYI1bNp7N17xxE4wnQV+8VnCet7sZfGOgovDX
1LEA8b0euPOw3BFqVqR+5o/TsVbS95NHC6TLgTpuC+5vxgAlZVgVVZAX57SfdOs0
g4OwDt25niG8BI20XlzHLUXLGOcpB82yXJgngMZb4kYtYAOAm+l8dyrg+bYgWOcu
eHBnTp1VotJhZx0GrUIYDQl+epG9+xmFY6w0tTZDu0nyGeninGLo20CIlhu03PyA
4vdEedu307IRQsh2CxMfepzFe+S+jLqCSxnvu5GOTN+s6SL98Gsn7sqH1N2XX/rK
dXndVex7RXJt5fLApE8sbtKCl5MgC75wgGYF5uOBTspCkcOGTwdAMLbLTSsWyzDm
YACsgH9hPOWKM/wyLbIkMxvjesYSNSChizZQeWbAoOU7Sq7lbJmT1aimShbwPX9W
VHxJcTVrO05gUrEvNfyK+06tn5t0MTGzyDV17u5KH+28zZ6Yps3E9myKeaFL5mmh
8osj2QfKKwwlwnqbatCMeuieVo4xWkiRIKPDk0GO4DCy9iaC2A2IGB8ZExm0+F2m
HcS9BfjP9xKxiHDEu10jZejELH+XfeSr6Adr+/uMqMlSSrpKNfzjqC7ppj+ya9GA
AGrRlvAjqACTUeZZGYrK+fRBZAXv+g7nU7mcYLN/mldqXBoj8uiV7khJQRZHr1cG
ZvynvtHy2Gn/s5xHbXS31z2hkAViECciAekhwmWNkyg/+Q0XNM22nLs61cPk0Oue
K1drqSUfE5xo5LJlgFkaf3rqQkGbpQtrwtPjPWWmNSf+autEg8tlVskziQvL+iek
Vdx+t7izg3X3Z117WEbIabzHslddrW9K5fQKaAqmuJt1prOi+cMLatm/6JrNtEa+
8/in2np7m1UaRQ3AO9v/4s+rQfyXOib8BPuBrkr6Dnz1pT0/49SAaEEAs6m406vx
vi/7A69O/r9nlyIax2T7ocPefUnl8iJf+ZJ/K5vv0V4kJ/5AnaghMXDf/vneEu0P
WHU4S3UK4oST7ejmr9q93mJlIoBdHOLVnYBiEn2p80ufOyE8FQRUvGLBRCDkp/Jy
7s0/6IOPel5pe7OFIkwk/4vHvCuk8juaaK02yJu9wsaeN1cGA7WxYajzkHERceVE
ueAkJdNNt6P3brKpYIRPZADKNdemIPKbU0MEBAO7JNCZP2o9PyE3E2ljxFXzG6g3
iZeRk+1o8iHKG7NB5zPF80Tu9cHEvsj+KKGUusPmkbPJXDIEwmSOTZrGNKDsj3dC
793avZnsqfvY3cFMhxtwGuFwijtNJht0e/LT4UZxTbKo+jKO9AIzK7pbMg4GsbDO
/DwY+8ld3tjcJiBjtt0Mz0spJTPaAD5w3PBbTUrf+Smzfh8BLHsPJlu1U8jRHs6O
CAcuiQQZdN6HRWYPc45xmjj5K+4KM1BM6tWs+5uicSXc/kxCErBBW1iW7QGrhYu9
/Yfl+bvm7GGle5KsgwMFAOEba4ACLltLz1UvtzQDEAcraZYXDY4ABDadzQa8pUiY
9ymdMPgkWbCrVEDQqpIRTPGsS3uaHz70hoiceW+nxYX8pNohHo1yRNudsY6kfDNh
ZbSd+vCSxaGifeutlAZmzXMHay5bqqGWVGspii6aWND9WnZmQSZ8Ci3P91kle2eQ
LIOIPuI8o2YvrJIkv/Pf9sUDO+kRbgKMcc9J6UKBPZVfHdKRCj25SO/1GW12VJDt
QMug6h7Mw96ePq7vJ5F0CPAK2865Wj98XbrfqVHHEqOHkRfoqDdtDK0TlETTs5Ih
JGyJwbycYXH1qOLR4+rgcJf3VU75Wpnigv/9zb9UMGM9DHNcahUvhalW6XsKaIj4
fsFqZZBwen6oiGPSRnapDsrv0pVeaM8mE3dCaXBOifRJA3dLGax8GWJqZkmWmFMP
mrXEzImtYC70K6N1V66+ivZMFlHhe9xJl5rf1OVKGTD6RfUivEH3Po4hG/0X8sS5
vNKLHBfdwJsNAWem2/glOJiQ6qDgOFRPx9OkvYGiUEf8aOFU7Dof8UJZJ+yq+I49
Hy/Rk2mF9hjDF2Cy2QaxbEDopvztkC99m9jT9JeDqBztTZwqSw7fQEElAJ/OQ5H0
0GJ/vx5K7cFeTlGRszRpfpaPAciPRQIbl9UAW4/zZjbmKxZ+y/twgrx6lJC+ZcL5
/5fFTLOxEBdnJB9/2HvxHAvpYsR+A4/424ath66O5aJYNNq7PPUH96PK8864H/yj
GFXbNVDcdgBaCcugBYLSxVmxL7kxcyTUF11xsHx1KfyiK66UHvSYm6pwEswaZrjD
xDcGhzB2YRgRy2D6l9ZdvM+Hwzmfj2p1rMS0i2ymLTMBZ5oOlenSex91u2FnXjko
ys8MpqBAahAh5A+kxzHvgZtgWs+LZygAbB0bNWhqyZoAwOnOTpc2ttkVGhh/78mN
N28w1wSDl5rQGDPjW5txZsLck7gbfvnBARPhP3m9g+HgPNWAXJxU7yfrAsfDrdAt
tIRDHuH02xB6qk7/zE3THjH2rnMTnwOQXeCjbjn06oYNV8HfRXEWy0PVlwdaLtq1
kJNKkG3AwTZvQ8K8A1JuXd38HMY/BQnAPn7lhHKeEbml7ojHsXJiDDEUmKHUoVt2
9XfdOycWzq6Up0JWJgvRsk+9iG9XLdD0EzYCcStKW6a6dwcy6/ujR3ojp6CCb0ah
b85rt4IK2fpPfnjOwXrOcq7jJaARYg0xJ8HOBf7+G2ESY99trJNr9H/PfXaO97FG
8nICCzKXEPcDgJrD1mN2nGg3OHImdooHAr//fVBU3Q3yp3B+cBy556YpFunSmwM3
io7/8SaZNiLFvvkWHuk9anqIZ68WdvPD09VtRzN4oVh05tHmz4cSGvmdQ0pN3bCK
WsIt0e4JTkChzQiAoM0S2FVgVor8li6FWqTwKmJuvn4coST6rWjBWf2wfr8WiIgq
MFLcpkSyYzWCd+EEpLGwk1dbVUkFZoOpVzUZFGToU1It6sSNxFOTxLwHgdsrvy/z
ayaO5j+abYJCAW5j3qNj/mYKdxeD90trwHgwU8FAEkRguIEYiG8mrWGea6m8ltz8
qCDKPq+9YctEgRlL3iYXVSTmGUjy1e0l4XjSjm3rIuu6q84Txp9GX1OAUoKFNmRK
oLvmUS89CFrNy0Xq/InSmNbT0X1hi6jzZFGaXIGO5akTUln/qqJ9pXoYjk7FRwwB
z6ZfYEf9N5O65kdA8+JK4Ri/cOcO/LXw3Lv5Qoc2CsUMtk9aRo7yq7Iie+vvb0Cu
WIzODzyeUPjM3oL0+r7KVv6RWet2EoA4KTVL7YLSidsM9/w53Fi492gJ3SPRvwuZ
LtCHW+6DCMQ/iJOhYvDzEcDqDdFUfUsC8Tv4Dg/nGDH+Fhb0YqGkWjxngim96tsw
NeUnC05AS3IwqNgZ7c0X0xIh4I/H4Xv71fX/s+2orHcoRyAtaSVc2zW+XuxM1MJX
HaklWv30hczLCXM3eTwLPJrwKTPuQvX+h2B4naZN6Y0uwgdEKp3271iwtZjyjasV
dfbzrieEmq1eQw84J7FPLm+FHfgYYRfRCu66b1EHq6LDZ4Fj16FkaQNayea1JreG
V2Siq2X+EVd41/NlP/vj47zDCcXF7aqAR4Rodnfsx8aYasdgmiLzBm2qGeKjBoFd
v8XCBUOMDrUNsbnGEbhoaxhdc8vshyqNH/B5UPXT8BUXw6iXFU9TkkZCnA72Pe3u
Cv0idTlLOd6Jxt6/5B1jUiOL/n7wHpvUuF8fVaB45jSN9DsGYKiNHfPRc/0IbAT5
xSasWHm95b2VezFHukrE56ngGS25j7NV8Gnwj/cLfQAkWQyjn+feFMjLmTqm03TS
tD4rXKkfN4w9HtBNz+Fe4rmvk75l/UXc2h8Jscd/62fE8jXDkZHD+H60JnvARr8M
2EcPq/XX5lQA5v0Cp8Sa4S9XCXET1RMhDQj4uCZU8pOQGC5bjgtKhU1GCrYhC4c8
kGdJgQlzkd7DumvPTCtM9ob0Z+euw3+dACC+avjX69lUlof02Z6vPgnJadXEKAjH
k7R/PZ5BDF+c6AOC0Gye9apuM7KR4sJBqO8DlK59tO6OKmKTSKFw42z5l9Zjpf/f
T2RCf2rTxBVpxT649RtevzdG6oh6tQpC8eg6FiO604gm1rkACwNbKyqyziwwkZfg
EeDeHjqMxdcCc5FFyCnw+L7fo8q3QPAnLxsb2MMxNzBi3T/5vMkblw6Avr5oQWDd
qCXnJhXpi1HTOBvOgjV3kGJ9UXOtSeX2JrM9q8mzCylsCJucqzDfYHvieZ4o2aPO
U7P3tdQ9IKD3YZFmfgNMbo8465FXD4Zl8ZOTqVeQzouAdIZp3bkWMJrbxCyPjida
ktVxsSJFb1VkK4nVVsqXfg3EjIVCALoK4C5np4hMPe3tgrPrQkJ49bvVqySYkTWG
5i+XRndcjS+QJ0cN6UyzNnTzloHHVDzVJ9Jg1MpXHWOFooDMe0h4sx40yzHOnIps
99Da/Ny/FMRcU+W5cZMkk9Upkf0J7NDHD3oNvJDG+CnsdjKpjhw/tvTfUoDHWhAM
os+xtK5e6VB1vsTQglTUbYccS/qUom8W3YLb6Iet6j+ZWgQ3tTxdvTnEKV6qb7Z0
VTKfVqO8gtnM+YCHykeQSHUpWZh4YoTzQtrvBBWQ0YapxAtGEfbrs/71HjkjnA+g
9XN4OAMjuDhAIyWbitpLn8jhRCy74yVQQO89HN89MImjNN1g6yq6webYDF5Az8oo
TMxH+Ytv/bEymT3m7wvqY+2YUIlShv/3/YLR9kVaWkhPbn45WZIY4eu23C/lGOqY
YiqGM93Fjb9WLosbMpO1Q3eEIBJ5Lkh5rD20ZPKH+YCaLkdxuwoJFKqtNSPjZ4cf
kgSglw2kF5QnAm5Z1QMyuWqaLV/RbZDM8FQ4FOB2C8m7yIX/UMHGiHZB8PFI4M4r
+bP4qjcR69E86Lac5sVDXwtSjtOGvqHfvUGi2P9YHwE4fHbiVyC72z0t3M7ZHX0I
6OrUBaVGXM9kVOO/QWbqDAAEbJ+7YADcmFGzpUX6gFGrlW+MAN8Zp87FZlqi5gYk
0/6tZxv+G48r/JNvJidpRWsnME015LCXiPxJHPwzRrOm/HENiPnh58bxwXfSzguQ
xVrB20hl2c0fGVt1ryxyx7QJSk+fTv+Qs0UOKGWGEHwaqSBXlcgkA3wcpPdLTsxk
toLwfriyWQzNeOUOprLyPsQAI/uakPi3e2O3j20x0kJds36rXnFza8nPqMJZPGxI
H7wJZ04B4ztWbqjQJKSVH22u80EYrdYZ4SL7SD8drvc51aQcktGdjY88/AfkRqnc
+mbyYk5Bdev1ofRaRyYrGXIClh4HiDbUa3//5VuBOkZ7/3qmEkh3tnsmHQicEpT4
8+NGgncHuj6nM5A1WjLkPMU4/mk9mkWNzMx20/U80IGEOvpKP6Zxpl1I3uB+9Yyw
IkMdWlkhBqkve8dvuIT6crrzG/Uk7lMxpkGZ9xtFvCykZnRE6NziPAmbQlIKunDm
bfBIub9pT8JBQIqSvse9D5F0Mn69FbOUGMN5ZoXm5FkzURmoWXn4/yslM+JetVxh
adpXOId6HHyceyjvsu0r6lo62xGL47p5r5YxDRSoiZN4m0thdRts2AYyAS9/TMG0
7smy32HkQbxy0Mq1+pbCP5uqs8czxvbvcnNEKLmHocVfC+4dQxG3taWREwPhQarJ
JF4r+3cB3dL6wUXH1ILneieoVOicIydvkiks5BZXoTDh0A8l161nMi/eU1vsoMc6
RI0qLTJArgD9UFmp7HAk7/3ZyyMirVMA6wC5q4m3Av1u+B0OvdHreZSTeqKh6UPl
rooYUkici1tjHrfEGR431yTV5UF+Ldo4Wk4B8PB7lBaTXT+Ire9Sa8DK/V0id4gO
uJiF7RyINol8ksZMmnhDo+qjlmrxUYm26AE/2fSAvkOTrxGf1+Rl0zwyHdxDYY+e
Fd8AKIgIsAvrq/ji4Ud1mZTeVzqem/k3igppGkGcExs6+PvDe48qSr4My9P8xUr7
kSi5kM470+q8EEMkX2ymaaY2gH012+1A65+QNhI6hQgSwBG/wtUsmA1suUT6fU9q
yWFc7K6AjgYTogcFjFX1wVdozdMXQdnavm26UUS8/96wj8kq52FLnj/A+ohezSL7
pgs77VlE43Smy2FIxgHcG2/KTnn4nU/q5LLw8NVOc4IIWQGGN4RSr5PkkJGIOQ8T
NDYmDJsUzzusednHl9D9s9I8lyUbGuaKcT7JEjHzxBVGx5pU7IjRhTp2m9VJs28Z
akR4hjtIewcsDts8m+9v0t0/K6mg4QvtRFJjYZLRWYc7I513tMi9yP9sK5VVkAYq
zb3vUcqn8RVu1b+iOM9UBDqnchTSjLzUTM7OLxydKo6S7LVF7cu81Qm9kiOZsFhP
iehEizY59rKJBp436/9dw+HEjlB7f2+zedi7roFYWXoxPR5gErA1oqdRnlJqQKLe
ALjSt801jKltP+USsYpnYylPrr2H0OhPk7bNfamQSak2WfVEyqyWalexALuNcQFT
P2S+wu/Svia9Mr1WLncbscRVem/tErQvBYrBh3eg8eBk9tsciLvOrBE2FI3YF4kA
PxNyNzOOMA/HHcTkj33cYHjx7VWPmUXnFlrIrf3g9vmKM7L98FyL8xJjelcNIeaS
fS9ZcOHMkMKnxDA8hWyktoAOtmk5hOZApoNwi7A7dWMmv69I2tBhZcA0tO3UBFQX
zZwWjImL5963AIB++YENdbRObRaHadkFhYDYsp09PK7Pus8TcIdoLP5+TqXdVrm8
qd52NLo/uCEDBWshGotjplOdqWPuj7VhFmpVwA3OGItRxatrkhmAlC5zul92yu/H
MQ9lQWo68Iopyldzt1ZfXSMGf3wG8zH+GggRqXc5HnPYVWJZlrfuoY9E15i46nf1
xhfzzfYRxW8iqHpfKMRnlwHVg+mV3xrq0tIIakBAPEKQCzxjDtaBcrccEi7Z+bwk
bkRKfhPfbnnhp7MijmUH41/zuF5uRFqLr6U+bfo+Q+luFeS20vtOOSPCo0jCzRvn
4spSeYA6vZIJ9jvxYSPgpozsbSx+QDXpp4XnVfm2Xo+DekoQLq51SfFIzg2+4dNP
pEdz8HteQ5OiHvdWJkSqrmSsQ0psPoWC4e2+a2E8NNdbTnpX5kWzFGI/QKemvd1c
b3lRWkJYXT7Vkchtr81fGsQ7qTJQeZWcTpWDDh/e3G3QMA58ursc7p7Baom416jm
iEUGRxK6U7sg5VhJ8XHBaC9tgy7pIx4a0M0smVldUqvDiKJbDLmIzRPuP7PHatb8
FQxvqhMfsY+EAUhtZ0A/8bZumqcql/33+Xs7eMYH3SfVFogTQzwRuS0OcTx20DXk
NsySnpO5teKAy9PzZkZxjJkypbzSaV06uJ/wWQucvLH2izs/okSdNWwh1nA27qZ3
pLNGoA68JfZa67M4CpElDrUDwkUXCwfr7GknJsGH95jW/ghkluX6nMrtVEk3NSZv
fkMyN36/BFUl1qk9gz8aSDKvcCpH5tBzjRYTVw7L6TU8UUJGX9LUjAm8dxtZ2g2s
qwWgRhWuxxw5rjh8WwyPfI7XXrJ85LF1lzgWXW95WjuryIEt+xE2PPDupJ7oMxMM
oPLDEfsXUrnkKO65MkUe4hRPYZWzdTr+jeQSfBXwmynDifCIg6PrR+NSJIe/G0Y0
z6P/fzz4VMgfQAs9AYAcFtwZyCYmavQdyB5D6q1YJ7dWV3EKE5NAQQps/1BZyE/S
FWzrJ2PEksW2CAFnNzfBYN/OOiZp6w0j9sFc/ez3tPztZMCMPeuX2wXITNXEJxA5
FCSkLf45STGddHBtU3jwzhD47qnDrSx1TsLrv4uRiX5okAmwg26UwsuSw0zH9/k2
x9MJ1muxkRAXOgoiwREEzAUrY17FdgLZP4ZXYruIo0bm3xCaiYLX9Q5blJ8N29rp
VnxIu0GNovyF4uapnffLFXo9R4rQFU6HL7X7RxD8PlzdNBPis37e2043g1Qeyl2j
QYp7ojxdVrhJiuta5SKfpcaZWP8uuGZUit0CX3duHJigxCTeDj6+wVrmpl3P5AbU
pd93JZi+43NcDdpJU5+LzKUUO6QwsoE37MgNcseY11ggXyeUL9z/ORFRZMJ2nyNj
Y2Sge7WrVcWZCY//UEtLif90WocTV0Rx8cwB3o52N/FdPmE8i8GWeJwsEOmDWjzb
vvbIzmFSA8DqJuJUYaSHDYd6mU1iL+8psDRL5YpLqKYwaHCsc7ih8e5pH5mTPSOU
7BtIwHJd+LY81BNnnFyy2QCFQgwJvg4AsvXCvlmgTQcdJby7/pYk+QpCT4qMwjKY
cuQ82/zchoN3Ox7gkfUmxTae0z27YCBrnVkYd2fyag4eTkZYCccyXRF+m+QEeaFT
tSCP1AekBRvLQXqGtqvjX7yfCLWlMmgJkEBkKqdWiZr0tfvXB/8lf9xP19f0OwGu
Ng6IAtdHwDMzGZfNkoqJMQu9ONB11hfW82aIO3PMoDOgkkAXRonnkwAkzHTtE4pq
aHIXpG/nJim4CoQyHT3k/I+e85zHCl6HVs9t9HiOL/EqgKZtgokoybv5abLjzklQ
YDLMEe0MJOZmmNHh8EsYKBhoj4HzX5UUX5A1JXVbgzEnFsJjNvapbPue8tIhcVzZ
veRYvfvuDVE3wk+ng7+eAj34jmcNUbkrYhzx03p3IMuJuJ7hhOzUMw/uiEST932C
0Ka1LSTNtvJpyGVA5rMR3z+JXg0oVn/24M7rTfcjzRtMiOi+eaPQfS18BS2U/nwl
SxDCccLC9aA/LYTq5d7v2JjD3XnCUCcEqeOPtTqwA+c1+U+9ySUjgT9ypLVcmixr
yBOBlUfP6lzT+V3BlunsiNTFCMwS8BxuiLyOTzV6g/AtcnusLmWVu1kpd3n1Iqtg
yu7C4KF73v1BPAHBQJJDSTqhr6x8UGjeoGpD1Wwd9QThBHHErun95BKjwO2YddNr
GBZDdS+FwR01htMdfOz0DTvU9lsQI3EbHLvVsSwbp9FSehScPg8R9DyBUISQ6aeL
bOSQ+rx8qwHinaSvcnqqov29eviFU2s/iJAcHIrgFrOabDvYWx+vEcsnuhFEapop
f8qnscl+kbNA6K/NAC8PTLLXaNzzeuS2OQ6e5p65crIGcAQIj5sEU1YDcmvdaR9q
lwtvHMc2HPxzdef03zbnezFPT/XnVL5gAdMFYX4jB4GooamGj6oG//LyK13TgKjk
JDmwOolMROjzt1xY1ybE95aXIIF3PfgVEbx06i++4ZNE+J3FfdRQKAhFO1ryxZSU
6TOQNNW0PaRB6qBe07/thqaqkz93y7KdI4CcuqxR+zwaNv9fm/Ki1ZMzsd2ZYYsT
ZERRbt3neltGQTifFgKknMyJUG7ZtcM/NiF0V8kKXKiyOHW3wAyQI5zI9X9F6CWb
tasLOsIeSoRmGodyGAusEgaVSV0c3R09fPs9wu37QYf5lvQP1NqI9qPAgIzyDRNo
eZY09Atnv0DSza4c8f8cSjKbiWAjDc+9n0XNs1MR0p3K7p0SkwMgZgcJMugtx7Cj
52v+fufJgZ0oz25HTmfAR+U6RMDL7n/IcFyCzpoKfVqcjFnW0pTeh9/eFgl0h4DL
oXFWlhNQBKsTaEr8EQah7AspEcGVvbFiIQJiwDSNIhUH8mmbVvDZhqQVBg1/ZlfB
8WUJ4jceoyRso1XGqC/qH8B6Wh/pc/F0iYglSQ3WqUTVdgDVzwYkXzHsqyS9JFB7
1uHrwJh4L78yNqMLkyYaJJ1mVXhalmiqZgPVjkJb6G73ADQIlStpD7u1ukVhz9aS
UGDotBdRP7yUYfXkVwFJJkXSeHebezkqVOVxGslUQAYnNgid1Z6GHuQl3oOkn12w
cpaAgNlwq6eSYIv3T/ZPlmcDglhdmz52mJ6xFgCRkXqtNehX0r8/38RXBYOfBuF4
yVVOtKyF4anlT9jUUve2t3a9Rr7O5nhQCv6MdVs63tUxPab1UfHWhTK+dqvOQXFU
SwELEGEQKfUSAodXDu2fy/gB8echmK+PE4PbRD/VFgLrJaqVgnOaO3mU+Kkosrvf
eZiM5/dUtjmx0PHClzAoipLcafPi0JryVDsPAkpGsn8Q0VRa4zDhQKxULQoNMijW
YuBK4xmU+/b9AqevlPFZkHE1HvRRW1OXWzJpCW3uKyoIlrqUvAqfNZa1tYpxEgTM
2u1ZQKMY+RIXPsYn6LhtaiZd4+wVI2JqeOtSDWrm7Z8MTafntmodiHTLNwfZNxs1
To+3aODYOj2BrmVAU1Z/JxDGaTki9yPnespXXSxwRlWCyWW7zJpR2dzMDZTr689Y
+FQOEIV+WhqrFpy2SSXdNOXsZ6aG52W50Qz0l60DoCwqog/rpYr4HVwLgWlC1n99
qDxo1DgKqsuA3S5WW0IMFXwCzjnrIzJNSDLPE+hUMGHspSCH5s0HqrJS0B6B0dMn
WB491OgLJ7kSKrHZ0gPDR0jNOKo28uHxPAbvVM8wrE7cc1aK5gsu5rmLH/prPGqv
NTV+OxUvDd7FN7e96BxbLLakL8tK+ey9grA7D4mA/ge4T6GDeDaoECdqEM89t5Fm
Vg1ypV7BOrfhuZcEMMvFYHFomALYWCBzOvz921hD4k8lABnMZmOHnnILwrPMOpL7
B+o6Tqc4nmrvZf+R7iAhf2CRt2f4SYz9ZWN51MEkqZETNXX+66kTw02c6yMxTI58
2BscfwioHeBYwlzC+P7IML2NNfZUgedtSOwqgOYUejMHxKXerg6BvTk8KThwUfNJ
ywpEvP5Q44UZfAmTHqaPvsJPcOFpwPA23tHCpXj0swW/PBKOJc6sSSUmVqaJQ0eq
lYrPZPxx/krAMSfEYG/jSqWvAZPTHQeqxf3v8PNk7erTKG8u9ZI29b7lJKlcG36X
7bE14tjOMcJTIBpmmO8hoptzwDujrTbENKzy76Ln5qNYXrBZQt7ybK6rMNNgESXG
i4b/xbOOR8wgZhHm/HuiS8FA6IyVedERq6+rt0+/9fVy+FphmofnoO3C4b9+fc1N
5vIZR73wjg7i82sZ9Qu1bB6SnOebPF1n67m1kEz15eOHmLNnWjmOtsi2X9q85h+R
aB2Sxn9wP+CEbFyfrWDDbf4kzG8RhEaIdDV698k+XUd4M2s3L60e1kcqCy+Ve4/m
sKy3+l3VEK3UPqp69InOD8MpI8xPMS9HjFao1BGh5GwzBNv9UG6gWHNHlXGk0vqh
j2FyH8Q7ID2y8HFTTwmAZsQTtikpvTsnjcvTLlpcdX1icVNKhdeeoHTJQTNHXs3A
QAB2gKKBKsp/tRPDJC1AV4a3sd9+u3+sZE6JYAGDKC+BNKY8eQObdM7RDbkXgWLv
jaRcUW7h4MMP1mHMtmhjfY0W86FdhTrvdHZDmFB7J8M7BItSRLhpkj8vM6WA+jYZ
08AZuyCUulJG4Pg/p9vVAItpPOkcDaqqCgqMYIMpFk2iT44TEzpD9bIWVNoc1oFE
+5c/7gOdlxllu+utNfbOiKGCFe3U7Q8xVjcKIqC3iogf5XrhrJKR82yi7hTmJQwg
WSUZyxbilfIat//srFJJrJwRMCcSKwgcAdXHFwfZ7Le5A8qBqEupDQLCIGbffZSI
UcWmOsHeHG8j1h+h7llPLQ6OKH/3lZo9gORTFsa1C0rV6QfizmIS/laNV3FoXW8g
5IS1I44YJDLxbVKCvASlVe4OA2KbZlJuSXN8//ZFVpJbVqYKphzRyygQYHxpZetB
2+HkTWZX2GEiwBuViG7S5rKq3RN9FrxVcH/IJ2XcTrvmw9nVlKGTbodu4/e9EfF7
5opXDJ9IFcny+dXheVHbIMJoQ0qDoHqUqZ5f8BXHOmz/fPOvzZmmKzR3RKECHiWy
/sDuzwDLkyGy/NXJfX/Vb0soPzdHr5wdtvNAADam7tD5+PEeKWzfKu9JBc/UAUfF
9uu1INCxO2UbQTuAg8EIXMCkbdrSPetwFDbgycu9SnKQ9bFyw8uEbapT9g20VE2g
8ruTxg9hY2zfVtZd+8GbYIwDgBzk+NGaJGuGmtgx4tEn2+cjtfSLjqf58YiXAYqj
kQWs8k2h8pRRluznBP45Ay+99QN23y5bMDbT8XxP//fI/CaOxM/YpTJ0VdjQZedV
hilrDcLVIqjF+bOzgaMeewJ3OQ9PwdJm854TxidSutbdNFKIuuADYwCO6JMT79gz
uM2z9qCxshY2MrPslN9t26NCZAwIzHfzKiUXTVJlVHNpvoCYzSk4LhcZSO2kXo0D
Zi6hapyjOHxqEtVsZBbLnbwpbEUohO3TRIeg8lp3nJV70+oY5n+sU24N3/tEw+nQ
vNicynAWMGbKDbobLq2e74rMQBcJxHn/wcHsIKLpEVHIUguAW2vfLK2OuNRE/DUR
MpbEzzzsM7xO8ojzIw6p3AMRH5bVwSNHpdlc/4n7b6BTn6UgUM8WUyueWRxt4apo
JPKFYsN8LeOQjlBGOGd6um7BJJckTotk9aVdnGzubWN5oWtP5iYorUsuQWRkFTEu
JxwKDeV0QyIRmm1nHGrGFfy80L/615XXFmwHAm8njm9BzdiEV98DETSGy1O0K/hC
tn/a8OcUtJE6kRlQUFUx8SDjColyNzS8TME2fXLGqHOLKahkRbtw2TU3JUAvga3R
/S7YxTLvzVhRV7EZ6671Ul7a5FrJINcGGStCLn6cmoHiehQDTfYufujMhQCNvQWG
TVCC8H04nc9+7CZAG/ssPUyl/50TdK9f+oQwo3aQ57pt+ZPX/vrHTowM1oONRtNI
AwzgD9EuplRL/eoODb5wjlWKw0UNMe4x/D09WEcTrweLZVX+vpg7sRUmGRDi480n
OrUsCUjO3a5RxpTjENT8pwTDMSZYS8RcYB5W0mKxYFxA9zBL6BZ2QnnVlclbOZvL
fWWtJ06OglVN3df2q0mW4HhuBnjENc9wdBjnNVFuSk2gxnqg796d7uO8MKX8s2Fe
XssmgR8NL4kWzpfx8k9+Y2YNt7NC2yKls/sV8c4TaRLhXBw2P8mYmgHv/5m1kHpl
9O2X3+511LpNm2SSXKQgWmEKQm+SL+M/iaYFw4c29hhwKqZGZdw142nS1qEgKJAe
cxeIe8DlUWj6xAe9/epwI4Oplt6KzejEVtT/j4l+cinFutmNVFDNrWAaA6xe01Y0
2i+ilPTzunNJl3vJUi4nsFwiH6+Kp2dM7MDOvmL160eXfMHYT4EyhR+sqiMP33+z
U0GJAnemKI76Nbjp4QQzcduTjKf1aMvg124Cmala2BGylPZ3C5ZG/BxKWxn6X18y
PhHN6FiFMYKTFqpGrRohO0TkIxVVxzw4KTQNvqN1aLOrxVSWL5j3JwoqI0vh6FeV
BawSBfWq/heYgQRo+zZyamE3PAZwmNQRny+aYP/2LK6dbN7R8fUN2tfH7iivDYvY
7Pd7vpjwZrYDjlefQBY+ABJL4dw2ihQH1KiLZ1egkihKi5no//bZquJDnBV4dCmc
owjjeyx2UysbYLohTIHVJAyzJqERpQ37UmTxiYOeNM1H0iL5OFpd2R29cgb1U05z
GSV0Z47EM8GNKqLgsHjh/crlrweV8ovHUSvQ2L4yUSQlAow/XFsaH0iOFmLCoqqf
DU9VaJlbt3gQ1Ih3Ak9u2DF0JJ3UU5GNjvWxWjzEnwJm2ObF4pUThxq2NnfRW8Dq
E/YzoGPkJFUKkxd3IAZVg8h9yvS/FeEt+QOdN7Chor4Dig7igGMKxSIgXjqsAwCl
Sp+CDyPx2vrY2catjCYrwwf9LhtcByWdThGxmDcA6DvFTBYUO5b7/woQ2TzCsTeY
lvZ+xensIBXseARf4rTVUZXkEMz8BdKwF5dpZNNFVx0W1pouypaz9B8hFs51Su75
hJixeKFwOmndPNWgbv/Hrx2b2nValxxZa5HN9aQk/kdbkKqOME47kJly7pNBTYNV
sFEZmv+VEnzmscxIjaGggO1KMvweNX7IRn7NrtuD3VZUntmtn0kldTy6HqAnl1N/
uL+y1D8sOsOBIcr75a8Loux5jyANiYRaBE8GChjMFz96fbZ44RgR3x3SGVcWUsXr
dd0nnJ2loH1oHHGkgMl4FPBHId9jagHXWOKKEJA0/3ZtF29T9gZfpIjMtIVxCGuE
/+ZJpzDZLDl2V7Q79DU17CxgQHGY/aOz6eApvMX7ofeBLD7jEQbU8SfBZMTqllux
I9ua5MVY24o1hJk7ORTdvP7Bsub1F3nUYLwK21dsu3VkDGplW19UPT+658DlE1Pg
oL29aBl4MYtDuaEchoTfu5EEUF9qQr2eIqxRyVpMG9tKjbEeirtKIdFSz527wTeb
i9nbtat5afsq+J5GTBA33+NvPyprPONRWPuglJpEJH/vWzUXj8U47VF3R0mNlih2
LuYSR1yhm44acUESYqJilBKUAoPPqmgjh3iHfvzTkaurjcUdRONPbG8ehko11QM6
UekSS3HJRB4WdtIyN4dUrBLEFokhGKwx7VOQd9fDD7z/8rmkeCWazhWTwApMW3rA
yKCTWWJnH0EkptoMwHUosBJwDb9rYyD7DtdeYZaHqQYDpa8/F/4Hlyx5E2Mr8T3k
OdMdAktMYz1+FFXXe1f5rlDJ2iVySKADDzmoi6bJIqyhvvGcZlmtlMkoFFX0M0Sh
IxDwckXD9JSPJNUdroFoyiJ7zOlJGYAUaUzWg/yh27dRWMi9/UwoIoPYjZIO1Qp6
kk+LIqfhmROtb4bCkMU/dwvxJpKxb9FTiq7GIUsOGaAEk1A2Q/aS0ggYfB3TAIep
bnRRqExwHXbZL8+nf9KWK6e2K9BPZrB80X9u/bZinvoZUCsb3Fb0TABPC7h8a11f
raH4fK7t72M/ryW0WGMyEyvR3+8uOyhA4Q6GyZFrkMcjvXfEf7uWuCIS6ntMlWcv
s1IkBp2C80KCj3R8H4EE+ukGKrEep2if94u+ISgmm1FKNHclOuM/CnP047gGRBhH
EHP0vzQKDg2BAN943CoklMHnqwiLLwgNM6PYfdUqcL+HUq5otjaDciyLj9pLWyo0
MIbqtVMCRZ1noAK1MmWzbZR/ZO7lrnCg/DD7ZZYQIw31qKaQ6UUAMbnYtXFeWWng
arGS3NCd2YwdEVkG2FZET4fAVarkkfJx2i5Dg8A4haLSt4fLDMmHwIjXGvvqK6+H
j8kkSbxMGFQVeKct0Ne6boXwNvoNnYkleNXblnyWI1CA7PAsB1eWFpj4XMaHrf9n
2jwCzcZex8TyRam4yoPvhz+PHBcnf0ZJURjqoOvRX75ubzIRt6DY5SPHjMLdSk41
rxOR9Dpql4SqpeXbLpn0LU7/o/VauTiMhpR05XvTQ9yTo5VrGnvKpTgzMaOixIpv
fXj/fLkzA9PSwInO2DykxJc4R1h6rmsQ5bhoWMYusSVQa1+uQtBdKkdVGn8yhfLG
ChcpWoRchwStw/ATAraJs6sMyIEn4REsY/jVwRs0F8IpKml9mP2ama4KybnrWqEU
5/PjLr+AG5LXYqWmFrVac0sbm1/CE9OKMBxKUORpXMmMRxIrkka+Xp6HO3cc02uN
DH9TyTRJu1Zff2y31bEzfPQmvvNcbeJevUggCFhP4FTXQDMOeBI8TUyXJqhSFwa2
xJpuXPYdkVtRGttmnDE7gAoTmvsVZpmR14yOHxFHmzEDURSiW2w9x9VVH3MROBBC
/1YgPJvJOqWMsHDSQpsANj6HO+b+aq4NTqoAqEfu4XpCrH7ztBxKogiL+ZFdTjB+
yZ61QdU0dLwg2gZXtZpxZHKtk9+iaFT51RCOtcX0D5tMbBwYr4PImwNDMySld1Jk
Tdj66QpJdk63LwxTD8tNZ9dAorcx3G+/inSZFpNH8BU0W9q8j/5ExT6OGhxiZiZn
LJqH81pUvdq7qgb7we72gGsEWl2gP9QZREHrJ/5gtlyYkG+3OVqYNlrjKBN87Hw3
z0UX856U+EIyMzC2B5RCBtU2xThrgiHRUEERdY3ka5HSCIqpFZ3QeWQQH27yiEpR
+gAwQaXrzVzyrz3iUO9E0kO6vLGVYuSgORwXGRchi/yE3Hiq6iU5YNOew7mn69cy
BzTGDyDTDe0Of235Mv00jFshP5r0nR/nnQn98Hprj12Bg0niRKhuWbn1IGgaPWfe
DCqtXiT/lR/fZqsRaq7MCe0UhDH+e727om1jK/VgcwvMQT0JIgFWeqjanJQrj4yR
iWwOPOkLKsV1P3IkBnMYNwMeCo9kf71NlEM52+ZGLx0HWOIpX5kTgzUAft2mbG9Q
2jNAB8gycmLHVB+UCymOC7ZiBirrsx6GqHCnhjIEtkO0GTn2EGC25LOoYiBG0dFG
7V8hRd2QYaRyqymnbfEjefAtSC3zHv5gAb0jaNkHOxvW/jEz2aUmr7KEJsui5AVM
yu3D9MoYa4kHDcvnmVFkseYlpqLUXsjLo9u9JkN5DzOcpQ4WiosySJlxw6SOC4GO
Tj3tbP4wJs/KgPNfW+Dd+G4/VLsfzjt0ji7YRLVIcaU3tA/ZjuzwUGPt8E9iPKlv
J0cw2XM8XrolhZma85zhgGHL1yAVnGizJ+iLoC8TGTXyNnJ7AodIxpM9Rn7RY3ap
GPYJ/UVvTBX3Zdp2evp0TjO4MT2kACTMX5BPg4pvQIytMGJceQEhM4aZuWeWMkA4
KHs95qhI+zw9Rv7IulTP7J2XHAmddlzXzuPDSoz5MOHmueLCl5+/6u5siT7HAZeO
zsycSkEisJeT0kKVS15fTRcK24B4x6ly2SHpjU3J3e/9PDtkHHm2JQNMuf6e0ob7
Fv6nxBepu/i2uSv288NECP41r//TQvSE8/PEByR8hLYbmiUscpeeuWBzaxC1NmWE
+PoIUWzWBPxTPTL4YvLuKA0gOGh+brQrBJoxvaaNmi+8n+LVE3bgxA8leFw99DzY
S8CljJyzg/yCs2X5jfkW8NGVGpd7Zm4CR6Z0LdJOweslC83Nzj4jbpgGs1baWPn8
AkNKhQ3wPDWCxuAIT9/UXY/ZCnb5FWNdVYzNCGMTcStElsjR3bGnXiwG1gMoOK0q
xPaxUy1EhzGOT0Sge5mCFly+kCTt6ekmXYOvTrOi1ByvOHC0KAnqOUsjkDyaLtiH
6ydj0oID6g6C313SWieU8Me1/AbjD2lAWVkURU99EdBsyPl/L1lPwfuieFa0hfjb
4YQJfN6gobUSPUS1bECbfSuLbrueVFxRii3FNBIIn5EWaP5tjXYVnxdoXLBZPdW8
6rluvDvu2BVwXVjJgTNbJA170OLNwAKF0CB0SvchhlNPeesXM0zqeO3zV8Q+muY7
wcYk8on/GhCEfyrQeQ5OpvZAni9z7GOXhcSQl+Rh3TcZlSxtCJa7wDnR3If348NT
pXEXxrbpeZ1iM+CxuZJNvrMZUS9N36xf0X0zrmVQH72WuGNf0yErgFRhS8apn3/z
D8e1UBx//X2rY8dtcb6XRl+hq1RNmEv5Qt4h5sa/0JrUcKc+p/6ZOkRUB8+l+L0H
tO+yol2dSjjbDZI/M/1wro0nTooTAtdQCuX0wI1QDGcEwYqaDIssfBHsQrSimDoz
hDmhqlIc8CDiZv251wcBCkxdcYnxUkQpeSl8ZPsETwBLn62oESIctZc2evro5m0w
AojoCB4qIM7cGk6/WISJttqS0P79DwY7wFBH6iCbGB0ltWYGvqiOTGJj7cKJ3L3p
uyJti2KVIsOkow6TpU0YKbluwK2nSOTsikQLjWw0wwlyxCmvtjaZn3cFV2RvK6BF
FftI0Wt5mqLdsVIr8ayfpB5J0FyFeU/BGBZxzSL0dpE+HTFgPczIOkVDtsv4/7rB
xCSCnrEkqdqv097FXQveKET+dQ9ex2MG7np923xzWyKY7mbWlJjYEp2j+Xb/yHpr
wAPJqbfUmbOqmzDBkCDbKjBlUEN2ia0hLUVzm3PC1KH7SKHyzI9PDiPDl5a4/f2S
VaaV1KyTOiDr6e5h16Ya+dmzXD61p53DcOp7qW67VTEQvvOoqQDy0kMMHUmEvuYP
Sc7qW92n8dduFlm/luwa+uTguqaJMkbbNfxbpqGsSZwsn0PDiAyK4j4L6dbbDJ8y
NnIEdooXGy2XKNGBXB3aInvXmLdLS64wjDo5s8Pb7FElYrGIWX4xFRSNUTgkHvwh
gccPwWyG7qcxBpMGJba2Ip0YEqdWrHiaeGElopJQHI+5KWkGEtwWiSLvURj3s/g9
DNcneON30o+/e58ddj/EYfVLa2QCjb4mfdzVKJlMBDuCTp4EICMt5DHU+BGcwOIK
MblCCK7ndFIaau8lJ4vn+UhL1qH+Yy6qLzkmKuM9QyQB/MRljfw/EDshiKSX6Orw
JKrbMldcrV3Dm078XPsI5sP8Xweq+AU9E9CvQaoZY2RK3u17Xmlwvzwpbfkzr1h4
P+COHxi+yScuMMEQepOHxgle/vTnqS5/chqRnug+/Id/E9Uas7SoraA2FpeAvrX7
Q0A/hR7LStnLsMrVfqyqse6OCzeVf8FXDv33Nrd/9uDpTasUDsv4qQ9z7Jmmy1Qf
301eOGIICsja1m+s6WssDafMXu0moZ/ArdF43PMBW+LGMQyXiLlediscP/5Qf5cH
auGiHwt7Yr+eEqZiJgXfDsIj1eXMByR5RIXiEN2+zmGFbyu628ZMztEVSzzKHcO/
4g6NAf4WBJOJ5r9z/f+Z//esfMMWbvVlwNZKIKiJMz0lzyNOqb6d5BkAvzEXhDEW
sBFSWdpQ+H24Lx0OAexuqKVs5t7nuE4kI7O0rEceFmfLjvxcB+/9yzHCvoDCtQzf
8k/ZB/zsy2ipGqYlwmteG5Ku1aVug25UIa22OCzRGIczMvDg+QaJrBKJugrkR74n
slHp0Rf30zPLW1GwN5x0S7zFepqhof9EmxBJCuvHBZGOMOivvy1nYQIq4UtFANB0
YCGra2d20+870GaNxIDRm+zot05aZgMhh1M2MkELpiIabjTlewtMUx6nNFLjE1+C
bIg1XFWM8nfZsbwaw0h4chI4skmCKPIkj6vqUp20OxiX8qG35V28hIyQNdenMmUG
Umqe4LNlCakJNVRkG6+4iHWtQV6GU6CzxNIG+oTNCyLAw7hbGTugRPaz5Igki39d
J15NpAi1ka/otmbk/Zy9AV1ZPSXy/9DMSedY/rSbfJ/6L7SKltzcOErYTvpIcR9l
68/mNN6fgVFgeeHnsfTg+w+jZeI+gCabh4Entl+j2CgbL3rMOI2JoFTBzy5m6pE9
Fwcaa9ip5BkLDXaoJ954sWzdquVcdxUoCFaxNeikr5rVhjyZjQuCFywbeEQaP4Ke
Tr+cMT9Z9ByNiF99GgYnNi3bSybR4c98ltCEtWks1QKVdv6GWRQb7bQ4IUjUHQpO
j8PErurieDcDzIFCAI7Ux8TeSZWa1dRwNV+1CTawUMiqSKC0A/g3NOUFDNhOOoG/
nnX3o8NlnQWDuF252mNxDdLevLHqquvC2pYTEvb4IwQV+jSVu0kLA+T2/+jYXqFn
Ph3uHvGbyEIwk2IUzJRYBsMC6pjCjvBte0N6LEdgHmAGcaoUY68O/NbOHbq8eb1k
PkmYd8wdngZGx7qSO4l68uhcKYk6m6r7Af9pV9f0PqWocC5wHo4PiK1zMmrwNT0J
5P1bPNLWKKS307A/nN2r3oeeDeDZ9r75fCVh0yd2uxR92tIIYhMZKvPDOAtjSq2w
ZCb9x2kBETJsbXO4V1RoDCnZSiQyLOmMF2Zpv6w200ElY2lZ0pMgT03lLgAQ8kwg
epTnFqoH87eig7PoTZuIQgrB1lode05CaTJuHzJz9+Etx8aIn1NJ7BVoJXMuWB1e
+w0LHWM45KlSxv3/FvHTO+ikYuQyG0lgyZgXfAn4CW9b/66mH6W4+vqqI4eX6jCB
WTJP5zwkdUF5LGDSS6GPzHVr1eT+wnK5UJFoV9ptoDMqKKF3WaSuoxG44ye5jss2
bcmfX2kZ5OYrsUXO3bmQUA8UrouqigoKostD/7LQUi9YJCwzvn066lEV3NxhrLpU
CiC5tpq91h6EEedtD7e7K2vhDp/GHqPxW/fMNbu7/91RxdZQhlGGFYSGTz0k29L0
Q57O7tHChhY1ApNTxsmuUUgBBhDTDMF0v3hyfDZNMEqp7gHzpS+/YIRGN0hdbCad
hkpUE7hFgORPcKlMfL9ldaY/aDOS0N6oDnr0jPevIcMUkfy/A63+sOy7injY9dGv
8SeyLx/rUhEVV2PsdZtuheztd50uOKBj5M91vTfq0ai6bWnG33fm/g1rLBhwRnoc
1N0C4MNvDpSbUYanC+36/Ki2JbWrapM9IbSKTNJkotk/RvsE5dmGvP2BNJNcmfWM
Os/LzniXQacs64fcW6GIRakH8p+oUBuIG54JVEgVz2dzjGVa3DpHU/1EY21PZ9eL
zQgXITbApWDIGNxmWDT1P+irN8BS8NlfB3K/LIFsHcB/iHtHlO1/y+6AI0fGo/D5
00eTaV2TVopT7TrFVAHZiYM7mqH4zEbg33KJnbaIzGrFwKfPJ1hogpavoChIkF1Y
vD9bjufLbbjhR/dHLXn9pkRPqzRFfcpejv7cm9qyh3E8gUbG9YKf5kmAAuPb22m4
3JpEuiqerdVe+RlWuuPtt0ggtdHR00NWLBuAucfsekBn5ZHlaR1YuLRgJIIRcqjS
YJfqDmLQ3LI9VPVQ0ITRaNxW2wNUsDAj5+Zjcxo4luXjeIToxZK6Ffe6Uj43ZDYI
3pK1M0qBfFgqNnrIsZKPWN25eBv1yNzYgC4VZLGf7pwoeoXdcRgFrFBgbxIgjNyJ
/j5V4FUk4zyk9cRm2vGglkbe4qwnNadYBNsPWXJv/IUtj5A1pjIOnjmideeWhGew
v3DJId/BXzHi8kwMCKhM3hUPIhSgoj5o9MngaY2iawt3SLiYE7mzNyvYf4+J7kfC
/v1zJMbMFq9X2d7Fv2o59IlAEHRjLHBFkJGJjCUAaAA+QVaDC2374NTudWAsAiBQ
/hAq3zDL2r97HMD8NCOEvAEGsnSlX+kHa7MEY/kjz2q+eBFtuoVkqeOtAZ1t2Ixd
+9lRi27/Kzv4EN/k881XXZlwXvmcijIikWpLXOJ5J9oAP9QdL00oSAgK8r7JaXH8
PEdcE9HhZFQXXZuv/JH/N7sn0+PDRABO+O8wyB5liAdE4BazEArXhRWynOEKg0zL
FxL5ikKcKzmZW6fKqEEdWsXTFjnX0MwVEHqo7uMxbbKRl4BFrnm0k9Cbr3QrLe9D
wshyqxSB6GymOR8yDh29T/fMTWBngevk7jzI3OdlFhaxKRk670NOBh2HPLNPcJcf
PNnPmV/Rz0fIfeXoFB6VCjFpYmIHGW51ob7QKQPuC6rtFAUQ6H8zXCZatDAmMrP9
+IFNrOLuyQj1bJO6Zmh99sOqm0DKAIlthtM7mqwEdLw9aJfshDIbIXBlE+/VUZre
bxRkIphEkTA2dC6l4cps/Paxu1yI3iw6Q+kn2Gvcnj80ZuSEVx9q4fycO2b2QBjV
/9sHZ86u9Sa0+voEZG3XO320/AHBjWApt/mnWT7X+E3SOcCgGiA4Dv6pTZ5kq3yj
DeezVYoEVJXjDpO8WURZA7qVVmvoMPLe+0cJujfww0sSXpGqpEYNCJ4jKsYELHVV
Gi/Lt0maWAC4a2xaXbo3T43utgP67ZHCTMDe35DqqxUyKgJhabbnp/IMyQrC3Iit
QkacQ+20EiDUxHWmd5yuKH6wJnFhyp3QaIsQxnSu3tYRt5ON0OK4g2bcDFM9vzzr
CY9XFUPXNstglfwgWtpNWz7UePXq6Hk6IxLA2ww42CfOi2FFlEnKTOu7Ml27AD8j
THq+yIDG54DV4elNyl62ywHHv+gAka/41gFWFuUkm44FUeuP9Szno5lvh6Da364T
8kfaSwx5b594Ay9yFY0YnC+LmybV339DuIeF4+1fJitm7zmjNzLeOv9uvjXyAEjk
jwRSH9PvQuDLQEhhZ1VKm4vYe3Gp6zoBm8PyaRpRoh+rFoWT9g7WGDQLKylVsD/m
rp6vyAwtGb0f/E5XIVTk8U+5YZa/a0FlBoHKS0FQVCODVk3gnHXqRyuYpuqlTsRx
TmsD62L8bEmKi4roU1JHZOO/tbwDWu1HP+ljQEHfBNrXtavEYXK/AKdNs52UvROb
SErazcs10WWqhbfhC05OEGWqs64Fap0JIMkMuoLUyTH2rjW/Cxmp0MZcEyPnFdo8
vhc6a/rHe0iYx672fEnxN2WyuQ/XDVJl2OHZMYYe2HlJWzR1WUzeED9ROJipVjOf
cBGxyXrH4oVLXb098Wihr7kco+mR0sPeJQOlvHMT0EREJibgWTdd8bfaw6WwHZkk
0pyhXHs3sMWZgxXrk5p6/B4/y4h4sPYpCBDJ6Fs2XCD5akjDaHU/EpfJkGOLHt1Q
Amn8WH/3rzjVKumlx6vEMs9K3RGzyMMr2mBAue65gYRQ0qLSLVYPnGNMRGXS+lk9
bDsAv86Hg4E5Bmv9LjXHY/4r1dqU3MeXDBOH7szHmqhKjvc24XKz6hZ36s0T3eLO
6xGneWJ+SVnUhLA599yF7/1xiYSrVyDvdi8aHIJWodxu93jo35kzVOwpHqsYu8gD
5C2gIQs2k9kyrUIS+66k2fwFNgl4/aIC0N5fvReRAgpS2oOv5Hk3lN6SJrO88eLF
unOiRkmOZ61sXjOL2e2eBJ4B61g+uGCGh9Vp6RVCjirf+cFNonxRVMeKPcjD1FgZ
9DC+sObNxCfKIUIYuefm7UpvNlxGyhL1hgSte1hCysBSGhQ+hHS6RF3+Gf8CvANn
EXnAi6V4mn3+mU6f/O6QFhudtsaFXleKHLtV2etU0GYiwW132FAPKfBgKAgnuzrd
Y4YNa7rql5pI657lJv/7PsqVgq6KehpRklT4QjOtddQqjeX7YJYNZ+MuA1QWZR/8
cKfngsZGdZAuXTAmipToS4y7Wm6NbXSKrYOgbriweVLAWKeO16hfm2TPhTf0/xJx
+plWYn2sPn9fLNZgtu0jL+0Em0WP+wQ4PYI0b+teq+QtPcCyU7+jM1GSG2LCZNgm
sYDLqreEWktUwEM0G7Hmeyk/1Qg2kwz91343TwBB48nlwdDiPfWEAv9T9Uo8UItM
eZQChk2zYRrMPfiy7pPgMoirv6jeqqmFyy488aupgVrTBzttpCJIZm9i73bLwLs1
gMAEUTG5RGKrrTXveBKTYAsTiWAoRY6OkWplL9hXJsYaQmBWNnp+MUOQ1Gok+GyC
upE6TXqD6/Ez51qgIc64ctenxecZLDV24wcgWPaJushl13iDpYtydm5OmrWkQV1i
YG5WqUs7iC6u6UWk1Hmln3qhqmxGvlmVIxaWosbr9RNO2YuBLtAbxMk/YlBIOVsU
9J6S2G9OM/CAHPntNt8jgdJarFKYRp2mBVTnr51VD6UpJiCMfIQy28/Rl1Z/CKbN
8DDl7877IcHjfyQGJCWVaMLA0vaHPB+8b8c6O7DJoPYVfDHhXvikCP4a4FmfCkpw
BuJqY6qKhWc+SSHZXxN6dJKDSdxiTCZyKtL+d8nX8sUXd6CcdKFVb131Dx+1izyv
cP6EI49d61gXN7qCBNUQuj+PrwUtM/n4scqOtk+MkBVHckZvhQV39kbnVPwYcaFi
d5cZU0u53yXokybLHMusYhVmIEjlTHWq0JtIylnD7/NvGcG18vw43Ct8dDj8M3YA
de8NCL7LDGar7UuoEmmblivVdeLAo4T8YgI06kJGyVzDlBXLXVqAHF9OCuxuX3jk
5WBABpDfBeLAGkjfUOzChBXtto6uQdde6Dy4OF2pd8XMgQBw3lMnF5/CPJaGjqOm
pyv2AnjXlGWOOiDVsKdOJXWAIYU+e6HpJ62DxV+TsFeA3ramNnzyhyeO3HNt138C
qO3DMz259uDbql27w0T519UWFBInjgPiOwMVk2PSRFsZmx+OGDxjugbErW3u5cKV
sTKKsShu5virEN1N/tl2tUpwtBCCyfkezx4yOLymZ0CKlkvpcTWWJQ0kVqoqYZ7E
izVVMyu75C93NivY9pc3/AL7/K5mciksB9S/NzQpOkf6vTqScAiarolG/mIj5q4t
t872n/Zqh+4Av3gTxOIrJs3o4BU9gROHbN8fg9vG7A6+LGZkwjivmwBCWOyu88Qv
mXL2k3Ih9b7lkh8oqqeryinaFb87Fl3LNzhkYFnEWMlOQkxmI4HexN62KkA/0DpU
XnpjaLwT1xGJ/Q7wwPvU9FotiF9G81nFTDYrv4cSdPjG8GgvM6ZpTer70q/wX19L
sGx8yOZUcbUIM+eAK0pjWvlw3+zYP8eHvRgIo0TkyYQ5uEsd7tLz0tHURBC6alAo
9ESOGEh24aDMYaN0bx5uQPu5p+WWlR5Rsqiob2fKVxlDI7+y+rPdHMbx3FPMaYzJ
PFMOCHEB8HlavJjPzy/bqyG60IrQn2FBnq+TMMquGlgtDb1S/faSlASM7jC2kO5q
KPbRo0RdQ83OBFMBn1WJOUl6n31mnSFLN4Aydpy4Y2TqNRRjQqDcxTLL2E16SDJw
k7e2r27rY0rjGvlbJ6ghCAmQqZFGCRKfZ33/e4LuTtqwG9mryuGyndnDXMjrKVes
6DCWCACC0u1sQHiIyk7FUSAMG/UQsV0+/84n8lP+Ls+LWHQb9eOqhVwmcCxxytva
p8iHYlW/BrE432rbjrT3nNqbm9vfd0XhGmyR7P9nBRFxp0KPtvYlZDfREYfS6VwP
qeglTw6aMXnR0P43c0YBAHnofTSLFVCMaHFQuyeT8QmvR1cQxW6RED78suWPfcZn
nnwGv3xxQ0gcToMfC0pOe6qNmVpLj+k1X6jRu1HsgOU0bE/N7NhoCXcfmr81EbQw
tB2nLaVZIeiZd1G9vC9GarS+n4B2NUZjI4vTc4XNrrPzDdf5JNR0fBeFMPppQ37r
UoAMaigx6tcPTBuq2/3DsyYkkxopPcQFe1m9xQGN6JUFsCdoluEVyHUvn2G36hgT
QzoqlndD4+CYT3XQTOEoFlOo5bCe1vDk8/afQD+S15gCWQqITziijvE4jX+KKozS
hP/3RspDcOtJxJT1VU78Asn6iKh5sq4GG6oGWdIHXeCYTjpnPoH6KsDbopBKU0DN
keYE2ezY0SOCb5iBMsoS5bmDMqJQSucfjr4yo3+GNQrLAq4sQ56LBH8hpk2nkgkd
t+1Et8nIuVbz3sts5NSEvK+MQ4rz6YCydQNn4/+aa3me4KqTHyaDP1K7mrOeB5sU
KYSSTYDGN+hciIjzDR5XDCfPlEAoF8IuMgH6QfgVoNDwSbqTxg2IMfAWrdIb77I2
vi1smRYMfyNjbaybMuqseJH1n1QI4f+lEhwq3Vl18uqLq2PDSwC9Vu4BtWqN8g6V
GjQOqp8+X3bp6VXLClNlNmiGvwDa9t3pVG3ghD81D9VadO0srxCEhXwXRBuyCIwm
dqOSPs+L7ktJq5HhbkZe344lh8gTp9wCMrBA+0OVnKuytgYIE6nxnh2qDFgVKWDw
ZX3qhvjD1sGs06y5tPFvAR/ilO8FDlwkIdtILHTnhMsY0fiNCmR8qk68QqUWUFw5
C3BOnirh0NLOh2UwDabrtDIvPuMNhv6VURBt7dHcCDiM/u+1prn9u4pH7T266k07
pvkh0vNWPcE1q4LzGE0SmaQuUdwF/5hIecoki5FvqRFBGo5+8SgDy1B+rAiy9dwz
23KMZ1+it2JRk50kkBV66jk/p3p6hnyKCz9HV29KxT+nrPrrA4Pg6VAeV2Cw2/DS
FPNZ+oYsWWurMikyMhoXUn8XXBzYwHHJXEQYApZ555L69zU13pYnwbG/JgLyDNu/
G7KKzINbSsaZ0eYQTLPz4oFTKilzqOu8odqNBxZI7EsYtW2r8h+NUx4CCOgREhWT
uRcuVPpy4D8YkiHV3hvnADVPwvqxDWR21hjJPgM2eKU+9aBiimo7I9uDkt5HVTiR
5zd7G7yzRKJHpX4B8sdHpE9dt9tUOzDere5lzk5UWKYBDIOJHlr37IMIClV45Lz3
PtaApvgdXnfOM/sbAiL1rNxgRvshqTtFgW6bTdbetti24Ccg9RJw6fT6RHx5pKAQ
Bj3n8x7MgVVJzPxLnPqDiy7x6y+iobBIyq2Fh7FzJaGAi4itKLRKw8l24dWPC+1q
z7YN/BXPRUVvD+ji/WNRsRzLEOf+Rz6+ELSpv4TaJdRHsO7hfDT9OvWQ+D0A8z23
Bchkc40rAK3qZfG8/xs93qfY/SjyCoaBOzmB6fln5hy85/K0QZ/8JTsYMclUK/Kc
XJd/bL3WTPXxQR4idRWi2RJwMXDGCosePykcixsBNXmO/BJqupQRhRXtXKDwlY4U
qR46o3YGQ3M3n5oVjTbh4sUw0IBv4jaIX1/A0LYdedjs0GYT8OSU35quvjKwWToc
n744ME6jkSrKO7D9XE5BZeZwQ6kdkH+5JJgqt/88wQayYcEFSTQb3RfEbLsrdkl1
FrZQsGIKRbKB2F0VIydVAvJVmzQG46mJugwKr1Aeljwhnfsg7pt+UaYkFDJ7Wtlo
JHmKQ9cxiTg2zpDQ+xZb7SHr+rsP+4EnmeEipc9lqN9hJ2ym1rxIsOTanb8Drcss
7maUy9BW1wo8TgIVMFnsZLhQJwma4UCOP4AoBmZ9Ey2oAYi6cIA0RDDj7WgjIOGl
TiiSYb7n8aHumIj4HZF60p4LqRBZ//TQEjQLWipxpMT2ejX85JEZ2HwIxdxqBaOQ
sw34foT6jAvDE2P5MGoJFKeoLH7HwJLD88Q+4Pln06pGjLKP0TZbXiwhQTUBcZG9
ulzgG2TNqAmE/K+P8aO9fGY2hbFANedwtTnLC6YXzsxKCeRT/FOEevE4u53Ssvtq
MVqIq9Hjd07vRCbvdrCNUqv0wSQD39SRm+z05xHnPSTc1fLDPaAVSpPtg8UXBUFn
e2qwNvITS2zPnUQJ7iKD/NTFDdTKEDGmDhSenoBc8VOZGcL0UfNUOSnuRPr0JPJI
FNHQFl8uBd47zyvWXc/E2uMeHX4P/q6Dc3WQWEYY1e0bN++VvIrw2eyyewPWspp3
+CmTmy0pt0VacfHygWtfWJivSyfbxBgoS5HTblXfP0AmUyWUFJezgEtqQ/lfhSlE
zcCTQdageURhYlTb+kFvnytKPVa0z6U4S+z9ZT7eNnetv4+8O94HCW1/3R/DjX9+
ei4CYKk8vElz882Q+2bzW186ghD0qWuJ4iI1dptvsdrPfNUdnNEmSn/at6hpBdRE
EZ5MARl/csqG8hxvc/q4k0k52Pq8lImuPs0uifAI1qQ9Hd4qs2y/7jmzcrKvAfAY
GcxjUEJjZvhLnhVfz3jIz7B1B5MEOCUjrVbj7fEh+GkqkPrW1Dl0gS5u+qNd+H6p
QATM8rJXW61O3Zc4cHagXIZ4V9p0QAlwMrKx9up8G7E953rc9LUy4tiJcHzlzRnG
rRJoAMSF6egnGAVWQnc7AH5v29yb3r9YUeTCPw5lmbLoUmV3BwYhu/iBVv0MaTP6
9Tde7vl9tIGbuaOFzUM9kZgBkQS0be424zk0xxtowFYRiFFugPL0ZTGgj9eCyi+V
BhoXQpHOeZbiPX/aTjfmk5PNZDjawEJzd9ZzVRfg6EtMdMW48twVMTz76PdhvbSe
r8PDGdu4fM1o+oRU5sTO/pHoYE2jmWyRHUBP4CscnYyZkLgP255b112cF9tBEQo1
naD0yI5yJBNH5X4c1jxZzLUhRRYe2Lz28uCBU3ksNTz0/YMPh/6Fc9K+KhHTT9Ou
JHCfx4W/GdGp6X01c1rMzZvS8qHSZje/z4uF30s6K9sNaC21/1A9Pt3JnhsRLT9y
U3ReT2mvTm0o98Dq7pqx/RHQ7ay7PqBOjc/2FipOYr5ed6gwthVFA/h2mr5szSSx
9P71/+zFlVSs9X8/4qyOTZUdP5qY45g9KEmDR075a3t6wKq6bxniZs/C7/3oK8gs
ZXrmMKKKArG6IG/Xc/dBkBLa2cL0TaRSrxzJyRmaRYpLVRBddzFVJSL4gxRpGveo
F9p5jIVK6bMHtG/hzL4FyFcAvhwwHVjJMaUdkv5L1ucylJ+DLARwWSTBKI/UEtBg
z86E67uSn+xztaOkWXNk/P/OTsHO82xEBLfHCpMYEeBxbagZybbZCAmi3u79bgDa
INYQ35cDpKLBW1ypDHFjUbLDYls3PWR8a1+Jwfz820xturzmL6KDIA5jaU2/ehOm
sDGelTr6ZED0oBsxl36p5A3gQ0bp6HPcU1/s5KLtdwUigXpO1tHXD+oUL2udvMN7
4UCEUiNA/70Dz4q+BPCmsOE4ggihhxnSqUCKvmgaNwg4dwtDtj50hW5VOlqIlDfL
BpcQUdC+VvYjQYaZzVFIEwYIfAsvQm1OWtcs0MrONfxMstSnqh0A+K/9xNP0WrZF
I8t0KzXhTRFUtmX9+d/3Jwk2F17O9Vhuzub/HEaE80knDcmrfr5PH9N0U1mpP2O6
ygNclj5ugOmLoKIqt1WECW2MyXgeUsM8Ke67gyzRycmIoHiGtZekrHweHthc2sTb
ZSFvSXGNYRBif4VFcfudwAXGjMcgVJVwnUEaoHosvWf/IpaVzQOgy8yFfnLGVg38
OCknfKFgCgAixcC8kOIxCr0BRK+V2vdj8sUI3ThQLJ2fjqVHudr96W0MJSX58i+E
S+tMmT7avbytag+L7d1vuDPp6dA+1Li3MKOCyi02+zYIdgzmQJuAsJg6zkXsPzmk
+gEFhWR2Sk6v9ApBXaO7HO12QLeir+geaeaZGdOfYIlANbfLk5TmFbogHdgX9/Pq
sUgDtADp9saXFmvHKDEg3YBcjoiJzj6XwOHH8N2+5v23EZN8EWFz5ZuhiwQ4XbkW
8DJeLh8/pWsYEJ+7gwYlfANGNuaJOl/WBD/dQ/PNjVU8+YHSB//sA6KNDhVII79m
CC+acxWiStpekrgNRmZ1UWmi4JmWNCHmdRPal/bzSkSpZgE2aiU4/RxCwWLNOyAg
KIniZ76fYjPhQfTXWSYPd/ufrEoIwwqtko9Fsyxzd/lzCkPLKIYvmt84Twn2MZ97
R0NfRonZj2OFfhmjVgzmNwmv5fWpmMoNy7TJbEGvqysyZSUSaZJm4IOti3OPecnF
s5VNUa5kZWyK4V8f1hAaVjQRba3fOH06wh7MxYAx1MUCgVyoTlT6PANEQ6XTe2Mo
w1/uoAcyY0LMmuexVcO3Mc/w6+QCcIWgfQVbF8eYGbbczYfctXYQS45wXnb86Tax
FTcSBxcB+uH3RuHzfOa7hDxUaGJxArjztonuxb9xe6152yDo3HHu+m2onqut54m7
q6oQKw7KK/p1DlQMd3hzczaNbE/hMlf2KEbt5O0F8r/PwSOzXr7b5SUK5Wk+s6G1
L3ySmw6WWEi+oNiON/cvOUckkEgbAiPv+n/wFpF9BgMykAwQs5g0DvBbUhCAa3l4
DfjirwabsNHZz0b7odOQKEcJd03KIMN5VLYLsq+mmmRO9tYUZ+dIW4KxDZsb6khW
4sfQNROUYado1b1Spphu4AaPYPO5mEuYVjWftl5z6zy1HDGuUQsykQmrOGAIpAX8
tCA4V4VKi9fZ2PRrv5KMnc7shOgOcT5rOwlACJAa9lAutlS62QTuZt1PDabWUbHF
F6HhTlhmYAfzge0TugS2ohnMqZ3XnesAYKA/MVFy5K/Z4nIIG6TiqWXNMXsDjcwv
2lF/UeuvTEGUyFQZ0AdCImYI4jDgSqJ40E4Sv1qM+h2P5XNBgNR8beT1qut1FMGz
+/pCKEy/8G2Hiz2zLigkLuI8ZzWsMrOv6DBSI5gas0FodNNiNH9cbByes/K+AGM7
npV43V9r4UsKjU6SsCXWqfTCFdEoUuwHBf8mGqudKm+t06UVoYNc1w+0lYeoKEq6
hVfKS5C25Fh7I4wujWoCXnpcU5EmTcUyO0UsBSVmV3H9C28y6+RyrMWZD893F5c7
llcVNauYBz2zsqocR9/VaPTTFRrorIy6MJOap7j3HAlxas1xBPh0Q1SihJg+RtrT
OxrIvjo805oEumJHePj+2D78YdJo5MeCkp2q2qvFo2TeacV6tyaP/ZcEwibod5ea
NBynespaPg+B6BvMaUdJIlNtzrSksE06W4+7OhTpmf06xeFL4O7/8x8qTBP5jNd9
A7sQOv5A6EZqSo0XiNK3mf0lxmzb5tGBN4vB26cWsGgPH7UIcWZyJSpObn5UB/nK
TjTnvVs235IcvYDI/hs+4syY4nexwVPys6QPx9tLnGEoVWDbZiJvZhb4BJnbBLEb
Eya5R6sgZAn0YMmXcirHPK5tNmDQfyY2e6IeJbe5ii+pBcfSJWUonEm5ylIG980c
LWA1l2G7ok+tMAfsTsRVKM1VtvdEDQAyeE6FdtN5wJpBW1NGYV/CLEuuKjzqziaO
jgPX9CfSAmK1shvtpj9Z78Nebv+pqTOsCDNGKSTaBwSJXKU4Hgisb7nmXwZZhgAb
yoQnIyg2MbYhOW6Nk/XqxPdHwDtvfglOy+NyygjAUOdpLfUktYMD0eyXPjuYRdOr
6zKvMaVN414skJBNBiJ7UhdrqA5A9mvjGsySFploTxVzI0riA3FaHRXWhbFJukyd
8MMLUPmgSxarL4qZoU3nWVlvThXM8dCWDJ3TJgbNQv2ht+T9YH4NO3iHdd7UBYJW
O33OXS0vEal8R/3MyZvRcwjGT44raLYnWYnJdLDDFj2bPYpAcBS519TGFXkF6n2y
vh5GEm+USpwTeXhJA3TmR1ebxUSxj5eh7T8BcVjw1QcEXfVozqGZKROYDRJLZDrA
VTOLKhH3IP7kb0YI6nAmkUbWCknuYg7atPGNghCXfWdeukdTKbk8xCKIkZXvm4aC
+ztKcnEizcQVDuQip+7ylyrgO6V0W/Di+eQIWOlI1patmh/CqcyV/ukQZdNouG8A
p5QUW6vpCgL+AyRYxbKy1Ty9ko7VoS5kaakK/nuf2Xg9KXgj7+vhp8H7rL8keM6l
zUdHUT6vb+6Iaz5UO+Sae/uFCorv+XSfcVvvanFPrcCPgEvQ2sD9pszdAwMSvPRe
PMSaLYIDjpzr0okZoxHox2PRNCFa3xHbvK4bbSx72LPc2J/DQ0JCpwmB2XzUF7vt
ZS8WGX2Y9l+0Ifi67rtgnZuUc4deDR5xpsABzJRErTSe6fgoPI6URq8Xk2q4f6B5
wtGdf/mm6kglswvf7DqhNBeCmdYNIYaSU/r9CbcSgCatBCAODBeEvQgwJrvxB0Ye
iexvbWPOwcexuSX5LreAPX8yN2nE6DSLNhGttY95Yv7kBwDYWfs0RDvNFHK9PnkW
TOWLxWg0Fnx3aKJx9Y3k49F3vLXCHOddwBK88ipECaKqzFfS9VXSBNR1rwFoK893
L3lKOSnqIwE0ZK95hLPWXZdyvSnaeTPYnvmZZjHkVVF9itbdwGOxeyuihhJCTH2t
BQThqa/fkpox6+xJTCU5UlEr1e9gKFXfQM6VEHlawb9Bnfj0kolJ2Kv5OVWNel30
nTjvEiKJS+vJLMunQ73gpfgzTm8WWv2E8/eePFKcjGWlVAijP5vA+q4GFjVBTjgF
Jc2UpHm/7JO6mv0hsNSbdao6LmRx55POqWcQ9FnOctMtPlMPi8iEqJ8zlqnq8bPc
X6hXgpV+X7Ait8ocV/Mm4O5NqLwxFuDv9BNb4B/yRVY8Wuf6Ak8YKQRH47tOarUO
7M6dDseiWMzG64JHCvE87ZuoHqXJ1bixfBTP1DpMl+wFuesjbsiEZ8qroESNbhs9
m3pdv5vc2JviT/1pto8upqpENQSQa0B3qAM024y/digi1ZsYbzM9b1stBpqJXF2E
mgh8YftIY/NWHUbXBJWVah+u2gd7hKgqMZPBveSdldOA2jsztNbL60gyCzBSo9gQ
4g3RI+PUOMwgpsCmuHfXIbje4+grCat3q9iiRnY+X4IkVhyeRxSJieb990Wb3JZp
BwIzAl3GDaIs5jFM8ToPl6ndLCuOX1soFJSzDfHsQ889/r0gOsSiLCriayQ2NDVE
hvTMqP5txxoz9zkfJ4D7KhoCJGOf+MysIEZCdMRBWX4h8bRhRXGjPA7+hWhU5kXR
71J1kIoITcnuuS46gputh7nII+NNBR5KNFpV3Vcd2sIhPjX1VsYEwoDB8ROymTQp
vFa7HAdLgNfGUFv3tOnrQxCsnuVZ8fiucK2saWWdp0zj4zm1ZgKqPvs0Gbx95sTS
2hZDU1UlwWe62kGcnFhEUDWM8T92pkeC8R8DpgXYiUoM43Kkm/SYk5UY06nHscqy
IBr8TOVzlmitPGHEhpPcNkMiPzTqgnaSl7Vy+qNm5km+zVMTi9VcJOyloPjo7XN6
qN1Hquy+q4U1yIF/CX7ZoE0c/x+nz4mfN3meVySkbNv9LDtKqBNJo8ypyTyK449W
RZXYHg7Wn4Oc6QSHQbgCBXLV2aYoJYSPhEaZUxZbN2ptqr8UJaxQlpIpWC/351T9
LeguGWh+RqWgFc9NL4dVDnkVcoFKKDcIgvbYXzeq7taEdkOrE5uIp/BFSvd6FzQL
y4PiTl11DPAv6t91ujNztNyQEi/U1t3ratJUOxGME5aFM5FB8i78Cfi4AbqwjWfy
ASwQSPS9aG4+k1DGYLtM9LTjgK5S9gkUQ99MI1VR0xp8l616LafrXL9at8kZ0D1J
iVhd/Ux9aITw5M0GvECBbBtsGC4iG6xKJ9WAM23C1uCq30khk0bWnQPR1p77fT6a
YZa2SobabQp+xfU33+C9JfRf7GCVYi4xGW5kbWG60pF/FOQJdvCsa2Q0f8TQn+Sg
idlLDVqjp549CRkSn9Sr0oImaHv7pzN7SHDFJdWd7s/jXw8mcArfDHWJUmIrenBs
of/qHjPGP6D6ak/sNceZPZUrVPjZH2C2NvGhgC7iuahaTm+E9eAV3qQfmG9NQ5l1
TW2kvdZoNbnvL17bLwOsXCbGQG9mZtr4bc2WlCyioq4eWIdyMiosKQpyqBWAZnGG
wda+FaeW7nxTHI9OK3W9R5Na2IaQlopaqtgVqae3PbeH3SGVbKFIYZglwRcchpm9
YOZRcDJE1EG1ur5Ew0ejkJIgcFF2t/nm9JWef+eKtg64BansMKZuotYkF/+qX1tf
x7G92VKfDJR1Uko8VI4cizC5vhWxGMZH3LqFT4a+V+O0XIZBG1Zm7FXr7oHRjYYS
ivPIs/osW8a7jsnRpfjrHbAiRCEMZ1UqHviyAGyJDAqzdeXM227xgAQef0tHt3Sb
7K8O7wZKOsSJdqi/4ebdOygD07of1DpzLLhRqYbiqsFrzrGqc8No+/VQljuao4ch
4sx+9BZ1BOKN8vSm6z44Cvck54Dr+i17rs3VSlNjDLDm2Iq4AjBpMBhVCDSwjRWs
1I9xE680jGsswHbscOyX6WAHIBspt++fOSx8NWCvuQz6o11Es9hP1JCbK8ElAqCy
o/02hJfBL9Drlsqh6xOVdjjXo7lN2Ynk88gE17pj9REQs0ccOdeseAIAs9dteS/f
2mZLmkrUV60SrZFbgOLlzIgDgPs8IW4Fnl15HG2USOAwYtnYqVo6pvbBg1O5ftIa
CROk5OriORr3sKl77jVXQdW0XFhuhZWTfRXDXVK3XTa9Rpx9e1D0PtdIus5DbXUV
sVapAUG4JpfdPWuCYq3JZNjZGvTf4fgtqbVDTjoWkzmr7w1SjzMvgx8fcMq5yDvv
h9b1Eakk34qhqYu85u+O4B2whbOqoO8NqYay0NVkG/yZJ1glYR+Ly2+24/ak4UiK
N9Z0OjAoXKlhxiEKespMEKXwVS5FznY4AL0hE5OBKHFsVvJ/A2yG+Yc9+5Blda0o
nhGaRtZclGc8YXIVV7H/G/hhCeCe4M7QAxMIDu3nZ07WjbNiN/q/LguBUK5emIQi
kl7PHEU0ZIBmrbQPp5+cka7FN3Nb896uaERYuOAoc4vMpa7+/Rkl3us/dj3MqBJk
mATLNi6KKTGc5Kck17/JTdBaqgMpXml8YiKYuK2R4zUQyCmT/VkUskuei8Bmt08J
7/P8BfDu2vQgiODZsLElKTdz5/VTYUhd2t3bJgjgkgYBK7eBnHLLdPM2Fd3DNyBz
FZlrLay7Opkb7iqn1ubCEw3iSTm+E+vfvJ+glFSiZ2ypsHlJ5Pmx5Hz8T89601OO
tGenbttCKWuYt1OIBbBBpHSi/dYzPPFvIM8wCUbZh6ye7L8gh3nv7PktBSA5nVTh
avdIvEoHrM07FZq5vCHiKyBsbZ0kwueoA+kn+V0ttq3f+VS5Nr+14XRU/c+WZxpa
IJjU4mBAeLBF0n9zVnK+R3t8EHWNC3RBOR7u40riVziMVNxjhn1fFt0RswcLmn88
O1woNXVHHeQ0qvhwLmRs2jcUIGnRNv0xTsBK07tbTeCfu8saW77QYUaaMJV1MJ48
XhaB7fqspOSSwGCDRyUEIEbpjC5VEAGhJicstTwo9ZoyoO3XtUG5N5LcBVYnPZGv
qSk4wG0q51jnOGIxa5j9dpnhG8hDqnOVLlW/4T/gv7kyHByy0XJ23GS6ypnpwXpe
TckusSVWbkOL3vz/Cj701dQg0mEgnOyZ/pVLIIdBGXDNKhaWrtGMe9w27EviTEwZ
qMpOOFxwXGSdx5+5+TOc8R5gNDd04z5dRu1lL2iRklF3k3lFNy2+HfBAPptXjqnl
wEJuLNMGvmx9m9hiyz/wGUy7NlC68aRn+0IZAwleYZuMmjP0mtIxczVulu2a4TOS
XLfo5+Q+5JQZLdsV8UPAS3BnarN2mCbkhy7ou/addIyVz4gJc91q21rPksFdZKFa
eb/TwCYzaVeTtNsiW8xhdqD9JvLxonFPYwAXyeqee18u/nLsiAuwrhvy5u3ZjeJN
baJf4XM5gR9VZNpAKIg9BJIYvaHh8aPZsnknhnwOATqLOBx1SOV+DaW/wi4DqHUq
jeDNUkjp0nixK8g7fma0h7fdqKeI7yPipMYwfCa6Q74wZ/yYc7XHRiY9UrI5mbPV
jWQ6gK5CZzIT4+PolP+c3OG3GV9LhImwq3skOlIW69DyTeV1MtnGTCBvGuOZAeF8
JR/7GG36e36UfuS+kqLlkAlgknge6+YOtl0X/YNaNKVPhhOnAN7yIcoVuEPT+Lpe
1zL97VjJf3HLx8m06njw+BiWBufOAvyTlSk7FsRUmKTR/l2O8ljB/TQqkSEGVmP7
48pNsV3A1yfCVVL8Yox85opkic1CaRZ4uH6zVMOyrVntxgiZpayeaFCRhqjMtAWk
upbYKmSSIlTPLiQmK4QT/Jfbf1jj+shqAt8tCQAmA2DyJm/XwmW4MvqjTS0Tf3+6
2039okdWB8p/noOB1JsM23GGSFrvVl/3D6DDD9A22IM/YrsHWyDwY0bMrydCHQoF
lEaeb+dzI+5HX63Ll1ypLyibO5AcEz1tg3Nd7SJ4Jyg+ZvPYkzYfZgMENJDl//CO
JIHEM/PJCHVgrDnsICgh4J0ouzQCtrN1KzGNPEl3IRAOzIFBVpprko3Wrbh98+Hi
svkM8+Rx1HCncXFSz4MjR/qeXjkAcD/RqkiwJKPHpVj3FphbgztHeit1m22Vxapo
zQ7xKma/DOJU2z0xrhpSI74BGdLQUvMBlwnKcv64HS1yhsMDaPKPu5Y1/IFc26Ix
MMWqrzoMk1RxL+3s9vqeC1Xpq2cU5ALCjghlY/kYp7hOchR3JoQWG4oXQ29kcWeO
DPggiS1rG0MgObRGTTKRph9Q3rF9BqvMixd07iVIIhtZg51Wqg4505DLW7r9A9JO
UpR1avrkaDRjsgXaH0ElNZZF4RvqgAA0uzOvNo5i4GcCRwNWLeiB7OR/mPC3wgR+
hjIWNdpC4lqBaQm8TKJB+Z6mo08jhYA1mTZz3iXUQ+N1SJ5sc2ZmUw0Lor0dduKN
b452eHv5S7NoXYpDS2B3/FGxsvDSCywlJSC7jWzXzzUOsC1l3fmMfZ/ualRCzBKw
X/qYLDBu6L4PY+VnBuW27F7yd65FOe6jhseKIR1irITwVzsiOOlSyiVxcv9z6kXN
Bp3bpKkw7YumjMs00kv8usyM915tQPCT9/XIhS2jfuuGGY6EyAmNUvIFwP1qmIKu
+KpbDAp1SwPSfoPpAa8WpnfeTGTedtccMVngem6eNmU2C7JYB7OX3ziVtrYZq+p6
CJq7UYLi63Mq0xMDZNYuNzPOxzun0047WQW6U1nldO/RzxYPB+F4n3uPLfWPrqM7
aIOVE7C08kUF1464KIxB394r37dC7rtpTem0KvPIaqV7T2F95PoYvklBVMuaIksv
d2AdpnxzxuGL0lbwTOPgkJzzkZsaQM8qxxl5Fw68mEDi5Y4EnCF+13O3gwEp1kNh
J6Sqff0al5KRmXpC+b7xbnhypnYe/lyj1W5QYfOFNAejMjPHL7VPymQqbsp8RtDp
lRnYf2+Rgqr5Oo/WbOc9WzrG/thDS4/aaYGcKDKBGHQf9tQmpWVx3r0JYJUqSxmu
Qb88E4hDfkAUEw0Oeak29ZcAbKA79MHeJoddQbJ8s9rnWh2Ub5g4wLTqFrC2jDTY
1ZnZ9JDPTXRS/bxUFWiNv1YcptkAr6saniaZd1gXOxbFnadOzcPx/U3aq+tc/0Vo
dbFMmHKemMNDJqcFmLUYiVRV8/FdcA22GzyETaw3a5Xj7GxZqCMov4NbIfWvTye/
rNfVYekxAf8SNrSq7I3rm0bSNn3o694/wfI55OLyJFk0KKeKKD2lD5cyfZGoe/zE
Z6FK7xgy2pWSMX4aunKE/t9qVWErDVRig2v8giDTHlAZ31ftRMDSWyN1YgUjGkWo
dAolIgsJnDB25I2rJ/zzCKNg+wAnaHdU3HL1yUcKD2fuQXV2IuGNMDWqsNtw2//r
vrzh9vViko4F0FRMCHZqaABygyJLTs23avVu9Z98lCc8JnRuNrPCYmo9DLUhB2+m
B1ktg6kIUtHAyO31KGFmMekA71os7irgVbhU1JUEecUlrqASQTNF0XXYDR/wlXXk
3/HGYPbiftHsg4HCNQsg2QOWBIr2w+diFEjFKFCTKVqCmbxcAyWVb/p9eK9zDPld
59AtRcvAPwttSfsZtN8RO9tKpZCz52kkP3XofPNcbvWRLqB37tR/YZPU3/yltOhp
6JSXBEp6TpV/8YnPc8GlV9ZTWtfN/C1GvtSb2aIswoKaWheh46J060VVI8ieyQz6
mVD6gxzaq6IiWXQRvIbg0YykfocpL259aRJPPr21DFA0qPnhxP2u5SMUPPpVrqiL
2tV7+zFU1tsTMB5PGx+gFJvXHg66ug/NTNfruhVqj5qLZWKYcVsSGU2gNNSDUcpt
LNrENzXmxT6h+2FZyiTKa7ufH+B6HPrbenSs7T3yH5PaEaM8XDrHbGmBaSfg1bzL
oZQQpAUdaSR5Mh3qzeiU8XoxYIB50uDn+hecKWKsmQwM9fMGTqjSZZNRcua97Ig9
6gSqFIKwRP6BlPNdAW7/OX6gnrJbj67j7Y7WjT/KL2SaCEr7QBPHtKnAoae7WFEN
GLI8x3SFBIb0AP9O5vfN5V/uslaJKEBiiQrwKWAyYl6D1gecn/meizCW+/CnxXKm
51KZVsiyUaOC00x9tPzSIuMEOUZXW1vSDrIYyHTTbSjwAQ2xm0LrOlbTGqZ6VG6U
ovV1zI2DXl5SmP1RAh63RMFML4oHRERMrXgZ5hHHaD0toHqmmcv52Qx3hHJ6IRMt
kQALUzCGVZfoWbiWdUnZcsSN/bcb5f6Umn4/XHCrbKJu9WF6Kulub49KZQaQHgjp
PnUIJ3idHgcBkjSv1bKJY03ZfTKOFcz5husdSYE7VKqmMAqOcYAbfWLHnScZ8Tqa
YxZ8ecRnKUZJkgGnrIjeU0yh1FXtgzvK+8H44gYEjgyV3V6UWvEBz23MG7vISeha
aAIIoWJiOeAjBg4/f5f9ps7+WUt8k4khPUiEXrjviXw+DCczKwYm9lEVA9/bGPoB
jx8zoeLTVjWLKAEWIrbTUYSvLE+xBHMiuJq7VlPcarVICusSsBY4uZFIQI4c78Md
tu9a/KNwORKaqQ38f/CWbsoLGVxFpFScowSKc/AtxQCVZreJuHoW5F5Mww6n4vSq
y8S88apiJ/W/JjjWF+zc+ahGmBsPL3x1eZICEEHV2VWZoBRMDtz/ItPHmOl5aGVm
n7fPRFYJwG9XurFwPbQ+2giobjGxaHa6vRZLPHxg0Xkji5RSdYa4GaYKLHM3MGri
xrzG5f1znGmxD0lnfLqo2t/W6P+uiW6HXzwRMCZsk+uXqO8wE9LB1RQtI4/joFTO
el6sBK70lS4u8Y6S0WM+TL+xAndiXLlPp8zsxroRq5sIA1Z4qIpebNy5/XI4Ha9W
U350hzBuXIDKDNg/yQM6P4VRd+W5R/ofT1ueMHRQk7G8E9mRIfLOxS+S4jtAvBsk
o8Zye6W4D35fi2rcCh6UGzU5rkK4pd9ZOM8cqEuE1D2eldJ0W4c9r6otx/TxPYrP
YhLBgZ+UY2ijzfD4Z9TMimKBPQH+aprU/Zr0hpcaOMI3pZEyM2PE4BuAlIPF6Ouw
wKkTEn/dZHO/kaO7dluLKmWJzrNO4VOYk61WyHed2QDxhYKlolNqAQlvgT0m2f+O
RWBOoSg/de9FnTg+hhETA0fjpV5owWm0EGVMzRbAiluUa2TGXma1n4KKXHpUursF
fT055Y40gheDPc2POlCaNS8Nt+c9ggR2JVTISuaOtAh5BRYvRmP/Y/H+gM6/EcnR
NeRvMbMbeH2sFT3+SGcQ04tb5VRGsYT0N3mRhPb3y/yOg2vfKVbHbyxnX0Rk5nBG
9+UlXiYiPIMll0bHAprjTICaxNjQfYAMOUJNW5Op5lhYJ+q6ojZIHerM66FCjDV1
4bt51bNDorokuUImiSYJ7N729+4PYYpIZT3uGik0mrfmm4EOyXPZAy3MzjCwfAEa
hXF+P5npdqX4oX0+NST+2ER2fKl09uKDBjTbC2lgQGrJIdSRlYPzcZNKyHLBk6X/
88syWWeDehhPrBA6rPvOY8uOqrQv7dBTjPvb3CC3p/RN5/xIkBD/JUAAg6Uw4Nya
LWJh942Y2NUkXV706KAQaexsUCHFd74lAEtFj4/GvO2Q2FGljR+eSlaZ07SNtQLU
JR1Q47YVTnojmcSOqX2EEBnyj2b0WmLhmTqGjlkovzgFiSNtjBoIsb3w22WPG2Fz
kXAnStTFmVkh95p3aJj+NP10tx8C1KpR1TqPK/meJkKQPomBhZL+9h6GMaRS9mhE
7eumebEbjbiRPY8oKkfsjkZpuHtkpDNrg3wGQmONupxJqTovm9afQbDAETaSxI4u
V7edBbo13+TkYgvTJEtBRfuks0TWafzHY63UKE+PQBg9i4o8iaLe67Py7rHaqGst
x2MkQuwnibLA1Vwxt4ZS8Q1iwSpBwgA0weZ9OaNyw6tIvm6y2O8+ZBv+p97h2fuG
jKEKl0324UbiXcjthiOg6Dxpr+ttLIn3xmCHG6SBBvnhgOFAeIwJxXXFEWwqKgQY
7xImJGHeNTqevOp6q6Z1ki36EsSnnGFudsXnmXxkdVx9t36NwDo9ptH/gQm6AmHR
sizlEhphf5iFpi6M8vBgmhA8VzRkJ0JAX5HslmHgnNjJ8HydK9ornrD3wJ+xjoQe
OQJsE/+h2rsUeXkblWRnYjzPNiVxeplqaG6dtKX0B2Fsb3AZZEMUPnzRiMiG6NbG
oiJVfUjsdN4PIt8+W11Bv7r0MfuPvdMYbGiCv02AhK8g8PrX0jYf7mCfa56/DIkk
aBWLn/EbvBNsyKotGEDBAze+IJBnb54PFwtLkQYHDSeZCmu5BAmgwdvb2f7bOCSM
ZXjzwSKTZ/9ajDQCTWVsXgsnFypL2qnNQObn3H6jfXem+N8m9XGxb0+uwsCWmJsd
NmqR/ItWU5VVgQuH3K/+WHGnI/4tDtFyXStKC2T2adyf82qMzMreK9qmxwuwqwkF
IhLsW3wYgC/RgKX74DPvH6YFT4IGhZbWRg/r6EO1lOVdFcP5aA0+qjkw3auRvMLb
7plwofkeV2o7U7utSxbwo+HA8vyf8NvpKjhi5veKN3RJ/+e1jUaiyCNRuxVXntOy
A7BUkdDcU06tS+4jwBgHW+cxVMwStMlYrF1LQX+PPDhxLmhAGncOqOfQos03SUDc
q4Z43fblz/x3LGRwpJQm/0bK6r6dCdZe9TmhdrzD09/JCtl033VsuuCnlcXfkB65
tPr+5qX1dlwdIsDcqQDmRw+z9F5O0sz5bZMwozeTIxwV6elF4DdP/Wv/pEHY2Uxa
NFzEgiZgY7lfUuF8cFk0u1Gt0uLqmzOmG6i1iH/xmK1LyRXx1c158EamBkq2qtfm
7MLt89Z1I20HnOzfU3hfjuMg0qW8Jl/MFV7yf9cTtyZaBACId1Hf6OliFi/xBJjj
tx6z+DW80FM29YsfR29/WDdMajy4UaH1TkW5padqbWvoRNNC1Tp3XeMU9mKIjq1S
W159QMaU7T5NMcUpRAl919Fka03OEtS5RvuA04tCbZ8m9qLAo/2C8zNGZ5OBGO+r
fetEyZJQRU+JmV2HyEeFPb5xVLmKba+EnZLalBGVwdlTv/5+0a+prw53Tm9p2nld
bI4Vp2B9Gwt2sB8jpDIAwMOgTqFFVha64NhJIqDAWezsTIiANXUEEI6MmkaAet9a
d5dYav2MnuAgUAwYF2T5MNJeagYbny3gO0t2vASDdxnmiBKmgv6qXM1jJV9IHNUs
14Qewt0ZF8JEnNsC0E4YqjoH7PGvf9MG5vfAKDBNW/xAF1YMSA58Vf8UpA/NuWgB
ECBk/VMpRKbFKlpdgq57ddeIKu3UTHgKWye+cPM0JkdpB2GssBBBRJPxc5CO1pgY
Bt0sj+f566kOxU3D7V4aglw0C48XVCxxz+X2mM6d5ksQ40OgdQO8ivAHXVx//1px
HntfZ/ks8AueoE/oc2PqEW34HbJemiBh0xq7Zy6rp/T5yNJulOcuGuZNcCgYhPHD
VUeoF7aenbbaV6Sna/G0LYRQaDXq1e+bQUVbDsUgsdPPc7jlIFfYpdCMEfPdtICS
TxguOJoCntNQ9Xyjx9v3ATJjEc/ryuDykWRwBj6QCV0CF2YJExst+qfMM4/YLobY
RKNKTKBjbMr6Nyi/B/mRGb3bQrfLSlzXI76Nd+L240Y8GJcdbb5+ul2d1ZYeBRIL
8FvQ5MxlOd9qcFDeFcSlttwQNiZjtQoHRE76dTYpTAARpk3rKEd6Ga9D9a557Jxg
+GRbBdkh7DWVbjHg53mA9RP3ahnIDJ9zi6xGeIBNDb8YGL6w4GiiheK+AB9aGp00
WW99a0D2rFC9U4SAQRrZABreklGlr9Wx5yhAi6D2BnbZWavswXn632bnd3NWGni4
pH99g37sO6Sj12Y29U1f8UqDXhiQm/eTL6Uk8BGjbKjgvPZBzmZtmUjuCJrlMcob
DFIyLwO+0R9IxF5ztXkWkbU89j5s3kC4V+mkaXPkHrXJZfKH5PgyPOUF2rEYm1ti
7u7lACQA4LH9O5CHmp9gNZC2GTwCBD6WjPiHYjCENtWTDbRCGI49HVXlrWmZhV27
THYKJ3hFv5O03NN6JF0JEx/FdwBiSvgXEkBSAHESRTbb8hS/GDhR89oxCU5XjCb8
9cFN/ZVNIs03DqmCTO5ytY7PUtDETYe7XcBDkzvHGXcKfB1gWZ6lP7SXoEs50V4I
55xN2TBgUxF9AXgWE242KM3WGPb4fZOTqXtrOV5paKAdn70VqW0srROfwqjUrV98
eve0cWjvOCVYnezsyo7X0n6O6SUi5+1rqcX9+lOs9RI4OV4I44FkHsSmh0+ud40S
zaoc6X2IJJUIyo5nwJ+M2wDLYLSfWwXtMbUscnVapItY76Uu2B6EMFFZ99Vsbjxr
M1XtPu/5Cam0pPRuopAg/jYqB71rSEg+m9VXDuZ2KOTmlqt7ycmAJJx0fnN4wpaE
l1SDF9E3rq6DzWuClSF2sRqCYph34vFYRu1Vo157H7HDu+0Phiu/Gt+T7pGP8jH7
yHZd2++jh6a+fOiwtsvcMFHgWvmNgdEQNNV4TsdDhfU8rjUTU/GnGoyMyPRhTG44
SAcIedCifk1oyF/B35OOZyLdopy/xROejrD6ZXsuci0x+I7AJOnXTvvUDP1DnGpi
hVJJs/wiwvXOMO77G4kFahT29gWGqT7y/gknId0BhNL34H6b8KgefAAzWdti7bUB
mS+7l/0mnoWDMMi5uFZUsGbWyGwrWdPeJL8inAttmacKlQ4kju2oRU1KJvkkk8vQ
DOgWH6RyIz01xE5+qp0AY4PB4bLHN0LXtCixAwVcKvxdgFfYiOFOimMtCiwgF7hF
n7ynGGMkGYfHYrAvUIlMcb/MQR/IMmf5s2xMnHhCvgoXHvf7rVCK+z+u2C3KkGv1
rzVHYewcNSmooKUiW2g3WRBmHsFHwJdvjWBa4Qpn6m0idx15HKtff83qXG0WrBgA
yjjf2cH6fnl/E6utvDsS2zYJt8BpdBd4Sj0roEgV1xhUb8UB2LYYiKc5WHfHuDLi
+YD4DwENGVxwDBxsbmOWZaGOHsFu7d9Su6wXt6v1q2i0bhxnXUUNjHx730SGAlt0
wiL+/CYxzJe27e42l5RP08iNQyLat/c5iXyYF1Bdi6bGpDDyZ4YBrrhZUP50OL21
C6PJ6mKnoZX/xKF42DvtTc9pjLNcAgF3nnXv696vW20yBSWDYiitSiohJwrsLsVj
yAgN/hGVJUyUwHnENcpSDsmVsts5ZTb7etE6nVqsY66VWxn/fvDRLjiqFtpdedpH
RjCC9t6pha/QnyMExh2UB30c/vXNDg0dnrGtx0Q3aCj+Qo3LADePkWMkqfAUMRf5
mwUs4MG9JK7cEkDCA+UyJTdubnYyHMpbQ6LpQDJR7Hx/TUL8FsCg1/G3izIzCfOr
3CV7BGOBHYK4BMbTNJp/EWIhe9hVfSgBwPEVruFwcug+5XGN46vRUoenzmVaur+K
EpiAfTp4RfZHVb0i+3oDC6BVraRZyhQMyhLoXgmz9y6wTotYMdLQWbXt2J5vlMHZ
gpgpj6k5SWbC0kJ7dVKqTR3oMSPwGrCu8FJVXWihgJ7loaHOanozKW3Yb2LjohwS
8Y/wt16zHVhGBrAAmnKzOoeVM77GJYhnpeW9GtTxJ0lUVemW/UA5qjig7pByi+3o
hOcDdluIHta7AVt3fnaoWQCbvXqjeoSBqbvlJS5qtWOE1j91TzqwXt1/vncVtSCW
Jz66BkldxMzd7WnWQGWPPFdwK/+1C41ewB6qdofeqSaKsORbKI348o2N5Gro2fmg
TY4cBJNUZ0a7/iBqVw7qPvGXFMCn65aTYo1P6flei32perdgaQnK6IWSEwJy8wVE
0Bbwa/aNjrhWyN5skEJw+80r4jFL31KyWlDjTG+l0yxzG8Ce3sPm9Dimr3AlLlxk
94TnUsLesHZx3pLyeYZYsBCk3YFvftABoXZPaGfv4HWbz46M8HycbQsGCjwL6hMS
2uW9inpodXzzfWxz7xRH2YlUw2d0bl+w7Yx9j3MwLX160GsuhMvfEtII4bDUaByd
rkzHdf9zg26kKAVWu1pbiFn2x7EHeJLrKgciSwBvHg1tlsexG4WpDLjaEmcZsvYL
tJEcKdts2/JMz5ZLB1lqgka5BlBz3rxSx+Jc/oj4OLmR6aW5dtjEwp6rmsrKzxTV
d1XSDRPBcGanc8mVsbq7uBSTXtnH9h2ughKtl87SNoErgOE5eFIUo6aYfoqMlKmA
91gwwmZ362/pHs0SWCwSWwFryrG61b7WfezurWtVvXbkccOWMM7dOAnTIbcF1/Zj
GZIQx4l/K2W6tNHG32u+4CF3Uz0iwjTY0b+whwktLOoItkKA7nJZ8I1s6LmziB8W
WORgKgdHaQEyIOGOGQjzt8DdM6xdOTKRtYWm9ZTScmSX9IiAaWI9VwQwP14JNJvQ
nEtxnY6xImC4fM6CnbGx/qP/pPkjmhGjc3d4T2J/VRKXwknx7A+/3zpRTsbkF4x4
YWM5Zn3GQdO+NyyQ/zocycpAFZkeDAO0xJl8+zdUPjB/alSxwigtPnimCAIKESEH
p/EO/Bru/zJ1BPUEfzK5h44SimQX0YrgpfDw10C6qQ1L8G4BPZ7I97hmd7K/nk42
3/otwFO3j7Jbsqb4mU6O87LIrHBX8arJOMSK81UmjdqWgjsliH3kA14C6BuUsPsK
RzmY9otnVG2nmB5QKXSEAhM68mg3pUNZq6cPbphzOkP7n028qBUvJFpHJplR4Tbj
FI3lsqP/cfbG/DN4ww3x9DwnjI0rtkXv2KkM21trHhZUHK3A272WpsU9SOSahYHX
ym/+mbybgzgVvUHXtp1aZyJanbgLFKJLsuWYk5pcgxzGocjaBgz8Q3NOgL26EUBQ
tWBU4cVZmlw9Llo1BW1+q7w1Wj2ASD5HOLodGUHAYRqZ3DMZvBbrXEvCMVc1ePmz
/l+3ifD5Nch8UZhR1NmcQvBtC+aerR2Iste+zkdcxmNUKYErKCIcZ8GjQAzTzxnV
kAw/AgWfXi0jtkHsG8EA8Cei3uluB0roT70az0zKstq/tbzl7WZd4KeUhlRekGh6
g1PDAMHAMzo5Hmhghj+IfIGpqKWO+FDGnE/gHpKUrNDrgADeRjJrrTBVOUIIzo/T
gj1Pm6srCdFwUMOd8nDUTzDOoO7EMF0iUtfVDyaAX8/GCVWtTSD/t0CDBf8TpkHG
7ZBY96ttVRHJ7gYOSWwtyRqXLVeNF4Hj81aGbJdaJouqFHPWJvGAbsbk8RroAhHN
5Doquq3pSR5Hb9U2NL0R1uP5n1Gow46J25tol1zsrMfrC7XQY1arelfkYHtdXurd
bA2zbS1WUhnQFD++8FXYd7OpUfPSNyZOOoyYqdkKfi7TPiO06yp6pSoGAQ+td7Nc
xl+Cu+69deM7wtcuED9xsjWYCA9fYVYE9eLPjm9ijLpo+UKef88/1w0B6cmSh6Yz
UdwZSGx6mpK95PtHcS3fKHCuwen6DIeNcVjxLMugQ6BGelKOL8uN6t8q33sR4JBs
7GDBPDodbZGjcDU1/OxPAOZayTTyP41g9p0C/RIo44lhEoHKMmybJ6sEuT6yX0Mj
EdOjmgJo/kTTJbfWIRS4AzRiQDN8hIbv58PSjLVStzRztiyhDQRlB3qCHI6VnZM0
gAsVlCnBy3fWvgth/JeyDsk3YQf1mNKhj2Lwl+R3U5SxBoAl70Saou5AbJyCI2wO
dV6uXQS7e9FyCGRpKhO9cHp67UH244nVgwfD8IjUU9FxjBHmz2OKPRVHhd6SMQ4p
0Fj/8NEi/Dz1x7wtSwGvn6PPfjw1/vtzKv7EDndXR6yphKSnYeG2PKYBia1J96rA
oZsF/o4f6x5+FlcE5mJPjs5HxJo4LAlyvmGtgdPo67HKEJupby4sU70UbCzKGuy8
VFKwrhu9UQNUmaiKg1AukUc+6fM0LdNsSOjCnrP3ZampkBfivHbiqo+EGva3Hffm
Gwcs2XdZa4DhpUk0r5pDi5pcpLGw4c5zl5YCL7pYXPxlU8vaEa+bjcOQzURat2rT
CgL3pv5TUB4EZsQ2uIoAFkqTbCg8z9YIYzBuQzJkVeCPAr2WjxBAJdAKJ54gwrTJ
dtxLhYujTIHKwtbwQkit51S3WUIfUBDPs+dZ9G6WmuaL1lsmEN3u1JqRoTEOb98R
3p/MMe2Y6Nwat/LUF4A7S+iV2FSJivZf6pduZBXtGptv54D8CyFf2CcqFGYbYVfI
EDjgmH9OvkMxdtIvTB6XZhdu/V3JAYcWwhErYk7DFJickQclSW3dH9XF9QCb6dh7
CyGqcnEPBtty/Rairi+sqgWTYNu9a75vxr8DIOftE0cXcxKCXyFirFX62fVh7VqB
ZtNtxQAFMtL+/wFBeHcvn44bV9ViWsa/gnngThumz4JNKFghN46wxiNSh9vnjFuo
bgzUbrL62ZocFcu5mrHJ29iwuVf5WmV+OAXy5kuyuKEh9i49F6AmEt4gG2u4lF43
ue52yE6RdF25SpKGuEq12xUW/1taiZvT4tgP0o02IxSrOSq8H0Fjm1rV+7se/hEW
1R7rA7CAX2Cd+V9KfKk9rcvDHwcCuqNw3OlEjmT2suHSXcT3OgJ2rUBX2ohDVQE9
0uPNCdVRH7I110E5DyscnWpUV2f/4yUzXfZ8aaG/mbtAg3epwimHsZJk/TZdUQCG
q0JtyD8dHM5NU4xUNjvvuQQM+WWxmHeOPRtN0H3LXAcG70FNHQxCMyoh7+slGmtV
spSj9kZJ73xB0wwq04pznoww63L0T+OSKO5fqJRUasgvQQE3I9ssDeRxlN1v6SYy
YQBSxI2ecz71jC+jnpd+W2cNrD4bZPh10UbSiNFdvrMlFzVqNqo0jVjQVaF/JVUi
sQsPeL/i7krv10B2AKTKORjYAAizx8bj9RoKYzIif3NtXXAh+e0dtCTTutNaP3qj
AFfVH1OWcOO9J955NBtxPWhjqKErSqUKB/g60SEAVtMX2crI/UfQbzUD8QawnWt6
9I4EOvmj7c46AMi72L6R6hkigUYftHJ9tVm53S14SgkZN80UqAF/P1NSLLZJO5Ti
Kth1At4HqwL7Yz2YH+BTZh9blOeTz++9YuaXtB0qzr8huTZ5sVKxV0Tm3kHgz1Lp
6vksF6v7ppkJ2gVXnV6K+2fZLyFlMwxAcnkfhieMZ4A0VHr9BrsMu+UdHedqyiWv
sQmsgNb/DiKFTMTaRE0n9tai6YOUXc4sNPD05K+nXraG27nl7BfnH4WWttWSWLpP
I9QEvciKNTaQ2+1NSKkSVSFlaAgrxlgXb10EKlMZXiVlwch79OeBs3udtImPNuWj
BMPsROAZW1DftdlGoU+kGvKhdIo/etR7d+AEUEoigxrsvedr8V/2GnRs3UmMA5GY
wiOqrjQfSVaAZpPBZG7H8Q+trD/AmxhvCMYmo2Wi5b0arRnzywF8sMTnq7B+NYoM
hfgYLYGAOxIpNSyx5ApNCAlmZsIiLHO5dsDkVHr02AkbJqTI6+MlUpYVf9Ftg33x
R7T/CYU8Izk3DsD4PROF1Yb5hjjFSkEEGCU0tQ12aDAqGtu9ndGjNTHeWnxh+537
kgUrb5EQK1wxwydfVm4MQEXjztJnh4YbVRVDMLJyDEvSp805k3vRZkv/y8l0HmNA
tORujZTJj9jt3MMHbxi0PQllKdrqa6dthA7Ggxx8MLsgHpPSfvxj4GI3F6DFUnwo
FrMYsvV/o2vOTsYt+TKJnry4i9k++3beNWfP3Dtqj7ZQmUxLLCBmTPIDdJ6oM55A
/JJKo0csV4jzvSYOvlO+M8ZbkmsgwYww80Q8K3wTx7/Es0gsOofRdzpB+tZJtcwU
DXTuqPnLAkbWI4nqddJ+xnUDFREmfnt+fdgdNOt2Q1hFK7YhSH9LbtVKSZeo1aLi
82fy+GJ4/FhzOtZnWcQc4bhdVLU8mXKq/kg12qA9NxvnisUB+drXEfzZAaj309AC
Itoptu3njmvgMVC10h4Q43XX0klxHvf289+mToN85xopXJAyrRD4hQA8Q8Bs0t+3
M55pK19ovsE6mn++ML2El5lwBMS9WfSpF5NU1jLKjUROJFW3wrOeZMLAgpd6AS70
VsZUgU/8ChEJQOLEJOqgergFGfxDDM9qUylJcL5fEUGzSO6HO9n71APujDJ4vdha
mj8Xr9i+ChCafuSmzE9+MHb30LtPrQlpaFkZobBjlVtXmX79xpqJl+SBHWDS2vMT
CdwRUrQQ/AUwmJ8KE9zAjuKD0ZOZSp0DqDA291mrbGNmGQO7TtFhcx3EqphjkwoH
0M9XMK/jkcJFgS+yHakviRoyl9XlVnptqgh11pPenNTIsdGA6bYfdCLPeIFljwC6
SZSdswfvlI2IlFns/ZZZ06Z5CsIEqZ06eH2cDe5+v5ZwS2U3lU5pc4DOGwkvosCY
aNnEtnzRZ9KcPdIowqyx8r8BWG7diF699VI9GgRwDJM4XKlJa4LJb2pOKt6g429T
6QelchzoFN0k3QlZqPec8aB26ODUj5YG2+tyPUrhgH5hP476DErY3zcnOSNuCrfr
6DIdhofrzP0cM5OC6HYgq4jb5dhI5kP/Lw48DrYOmyUQT3jqc6lQPR3/e0m2YoTa
7z8UNcndK1oBF/OwB2QmWN/zUX07lsC7jqGwTAmCuX/I6Aa9sUH4E6sLQ9EsQV68
1ry52LYcMBpM32MAVfmckh5sqjCAdtVvwfPgau6JvEIrDJZ5rMVpmtbVF6fzYRVG
A47G+lZ8enxVUTlH5YfW+vXp4xbPhZQTqdHwpwqJtETdvD/msnvgnt7UkYvoNGls
4NggbwX9p7OAFS7AahEiorxFibiP/4nNk+d8MucvZFwO4H9KfduSd7n2xRXZu627
JMUzBtYL7OlTDBUdUMhpvsKbeTp3DCD086uw40CmwKdPlGJTSp57gZu6iZkoxREt
Auo+FTl++FNbrY+E4K+YgINWrZg+WICKoMgYxtF1BdgptVnVzwkZRHsXdGEc5ljF
pwHkkYOj2szyYDOPxghgOysTGQYZhSI0bweWKeDlDHJ38l5jKDfFelsh7ilflJHY
xtD1zoUocj5WgVjjA/F134EYprasVCECOpskOtzotFdYiaOrEozHkq/prv+8i7qh
lsQW9/AYWJV0UtSY3f/ENMqDD6MXKis6zmjUqNoXXLj2NqQohr+f1jWKp8ipxlLr
cm/+3zW+xcK1VuFks4fW/yyk/zDnirIgjY0qm2REFByki6D/TS2qMaY9V6r+fIGy
knwGE9NkOpVqOxEqOrXYFgORqSRc9evbtXYveGSY5Ud1JVzkc77ScDaJzR8zyufv
adOdTENXhvE1/52Df8o3p+9XUWfG+jzVeBtdN1VqxbZIdfrHla+NoGbKJZ3NOKsb
WDGGcLo9raZaJw8XS507E885hvcNBiWJi58v67pxrGtAlUymwL1EuN38Qq2LPJPP
wGmDYWbd7dPT4LpD+YqCuhnGiicnvYRtwjTzrubHDBJqCCh7vD5VL+LM62jSpsgu
0Gs8JyQPSxssflbh9jDY3Xv1HC0quqelqkvwiDDyldjgVwW7aK48S/5L+UvLoNaY
IGtEYo4XnXQSYST8CLqiomrCm4aAK0BQqxsWGzb8AWu/oRE5BXv/FFpZwbHjICJa
0E4NvRPhfE/XB2HlTcq8gU6XfY8ZMtbFmZp+m+uHwXaC9S6r4UydhAPR+1Ko4Af8
HKOL9dXzJt4nnPanWQOIKmFFTpSIDQYxT+BDpYji+pM4Pc2Vgcb8Agu8OgfmJkhj
7k7dVInNJsqFPnSdz6WS73sa0sNUoADVjksxj6d/U8FVqGMNmv5AGIr55D2TpZ+w
Y8DBXouCSayw3KtAfLTsMOL9szhIT8nxa1AV9apdlsziZQkYU3yMlg6m9NcACI2Z
krQkid2//aPzimIHJjRy7AIvtbZABgYjJP3sCS/f35CbQxvTk2fidjlHQsHrbqA5
BTtOfEkdzELbiSjTb3URv3Ytx1GS5nal7SZxOfLmzukAL0NmfGTGPqaxsIsb/89u
93invzGCtY/tyU2SYTQfo1nM8UhDPeH5A4s2VHz6UlI/Sv9ImZN89lc/QUC15BNi
KfzJz4MhskRNwz+ZXYUCc9vn4vYkOGQtqxAD4mWCjqljSSwfw8nH88hrhBfnmhsJ
iMjN7dhMuEkVV0O+GczNVmW/MY7MGy6CB3uZt5ktJRTR+J2s5oz1gGQZOdc3GFpw
UnP9nBCad1d35aQffFmGXNcD4Hlnhk9+jG1ckBM4LMz+XC4mUQRikwoyb/f1K7/G
pZIHcd+xnMXyd0sGnABlrO3jofJHcyku4YRrzd8BTlaASmjPXttu3fiF+eKWML/d
gorgDU4dw4jhrs9EaEkuuzg7XnmVb85Erc8VeIEXmP5ca0Msv3WsGv7tLtqMHrnf
VBaaJ+EQHJDTP8NzwC+3RNsX58LHnOqcjhoNEypl/wTI5qseGlYxa0nCiVmjlKWT
j9Zr8r03cJs37I3KdUKDtlo7vRU4J9isl+r0ZcwVES1oAiINdwelGbVUy5hmo2kl
wsOHwhlvz3n81foDGblPVZ9WCm8q6BgYCltxkvb/qn/SLvB5hvUebE78kYJedJ1Y
hiq5Qpekd5hR5lxul5xN1URxg7NuCOz5Cd1CuXOmUy1IG3SL+lHnw07PqGKEdcjk
mMWY/wqKi97fC7NoXcHX6eW4JeD+It0Sgu+4G/Nfm37khMtyb2psNAUOsWpY0sDG
tMm58fIQP6R5la8qy9BcTRINBLd/uojEYiBObS3+1ow1XGlS9UmjfCLfqAzE6btI
1MISciQ2XPJD5MhoqotufnM3yTL/w9x0f91FqTyeS10fXHJBHuSf8eHv952+s1KL
7Y/YXvRkhYv9xqi2v5YMME+F2QZ0a6UyMJf5b/IETnSo2XWynxRXEDrhXiXO8UIO
VPT7SHL5OMe5LD7Uy7FLsvmhp3J/loLX+Wy3e0YMQ4jatjMb5+H/Hb7ZY2i/TfUH
dzvXoh7Mm94+0hhK+blwU8LCMe94Y/R5QJnG3dVbtBEvaNbLAuU9ecoKjawiqc+G
wYwt/Qam238Q1ZEuZ4XeeywIzIUuF/Jtmq71cZwms/YjxtXEpFcBFBD02NnQ/f2l
hTO0/78IjaBWHLrq6Sj6rgiJMTIxLqq14vsKhq899SwOTeNvwCeaMt6bBWbCWSYe
ZLZl3koLjdKYth9jIAOkot8LJ07k/2RitcpaUkTCuJIrcqTv268cYgxPRUARYKFd
I9r0giJn9cvszQetaJ5gQ0gR6RLW/DFquLmaAybAAeGohBEtffftU2A9OkD0hcok
Tu5fszACbl35/+NlE4G5qPOFe5CCRNjEZVDaBlFygY4uVQ0BG+T2kQfw/m7D/RcR
TP3pu2NsUWK5KFLa0HJ5kiCNRQUchk6e893yFR9wdiO8IjSyjepB6fb543L40Mla
xin7YdabeAPQFmcIVkn13ciCn6eCAaGEEiOEhQ/4Zd2SvaBpefUlE13WaMiSz9nA
ZowbnIH7CWhSJZ9UBMxpwTb8uca5Jq7qzTBXv+FGlWUPgaHE2i5gtpu6MfOZrKoy
3QwltRXYXH8EwEjhmLozpZCuFjOClHSYu8NDu+YHqYxRRhW+pYZVDAhoVRud1GXL
qJCw6ch52wDeKv4yQ1GQfkFqcqHjzTnENyDFimvRzOww4mAhKs8wS3YF7VNhbSf9
kYsWvH6ac+BApN5v/iv8+BzI+EgzUjcJd9JhNioCYUuoId8Ahi3RhHlC70dkRn1N
s62VMVAOGLHFe03rk3dEEjtsBSozGM7AmMdVDFflfLz1+qrErigIQ3TXGr/2oz7R
Mk49ldSDv1BoikWhw7oHLv9ZmSM+5fJsjfCF1+r0w9nstrwmQhAvcMdEnaP/xNwm
ntHMJIxBgTVQMu5IKxHgmyhftEsizjS5a22FXeolgDJKM3uBV+hRGHcXMuzPivSi
d2gRKH+O7l1sAT99iToL6lkwpk4hVz34m8hHZ6oc3mR//IZStQA4auRpxtt/EQAg
HQYhvIjiLSJ+75hn1VasVQsaDnbXwsvd7RV5eqjVChIQZ/5fw3eLZmweL2TCVSCW
BfOe1ItfsEYcyFa6ych/5JyrGVgQ3ZpHyFlE05nrBBnAx/MQl79j+C4XG30z5bsd
TULt8ythewQqb1PAqmh6kyV+tX3hCY6TMFsnyE/Li6wB6KKpXFNODGvW1/NjPiPE
N/OW36vKLF5XtbG2S4q94p1rMPQDaFP6a1yIQwYA+f8gzPRXp2pLaOczXKc/y1oX
nJpC2xHgDNGiSs7Ou3GVbwjGbeFUMYpIIHmYcMnXooSamOMm38BV7rgEnW2flbla
2MQKlonKB/VY0tzEJnOKF75R2fEgb2WsgVBNF+a75q3wKYIGJCyU92ByCtJ+YlLM
u0VbrxsJQc8XNppswGAPA1SXZiVpmx+jeziZzQiG0PoFxtidQ2sLM1nVcSjhKOwo
HOyWJUDO3VGXknOiZ1sWpa9VcxIQQl0emEDAIGUXWRZukrd/VuhtsKR/ttbDxQ9J
yRN8oTAYwy3PFVqyzWvQhClLzbzpDZ07/TcG2jNUDuuoSHNfCJzk0Bez5BJOpzw/
Pfg8YNZ8d2BEKhFr94awx3ITzjJbwXKkog3IqZHannAsqOHROwkyzSViQaTDesKn
QI5YnechJun8eCyYIBCFnJAvBtib1DGGvq0vzEGOGfdkML5EASmwmkL+nozYIUK8
PeucdsTUzFx0xvqJ4NqNtQ6jJe74kHFjj3Gc+bZ531x/0SKK8UG5GTo4wZ31vJfe
eCs+XI5VST/ey9hAPmkOhDsQ0X3pu1QOiSejm/44gQJJ1jB2Y6cHjw9VxV98QSmZ
3W5lqDj5BSE9AM3Jh8zZE9SPbejhlKrslAb88uld+iYFQJMEYMqpSodyWsnliiR2
urFgAahzGYeSOlpjYD/IK9pGjPpgKzELF7lqKD0q2lHgHVZOkW2hXIOrGY7OsXA1
rB2iUpQlM00ICV5gAvRn9ob7HtqtqP5+4s1OlVQjzNGuyFV3nIj+dd2Ef6XW54w5
ALWyGAiP5Zi8vowPqo57K6378jHGQj0uIQIgd8adePIQGO15C7qEvEZaBBZ1IvG8
/JgNx7GY9xaNXNDbTctmp+VrnWu1v+b3S84AAF685PYb23gZOwTy+K1dXSLuWf5c
WT7woWMK7PPvw8PdviIH41iLikDN/7bMdzGuVjOl6VRMDsF19+PjCbykIuYgVn0P
jgDpniNwvOSDwE9vsD8RlUVIOuPr4R+mZP37ilD9WfdH0W2ieSA2MTKwPVWUSL6u
SydTKJytdDL//RAxNWFudcDmxA646wUWmPCjQXos2Ho+0j6AXTGSNkW/MlAizsQd
gJ83ukVJfTrLcd+zdSswRI12vDpeIhlupsZtViJvCgHNJzIcN/Lu/6wjeEDw32X0
3ixlXBx6P9MqD8dB0gKE3kvP0pWu6eZqVXJixGyBMEkXrA1JkvQQzFFdS9j6uH00
M4x/PYrsDRqVy9cI64/LNM4c75SINgphiSoICgkoCuCj/Wityx4cAxOBZ41YuXQQ
iWVVCSxvMsZJNj01o8kOKhY/SSk5u+Pj71reP2RE7hTNMoeUAYUuNJX9Y79pEp6h
tbz/jnE9aL3OLUSkoNLgzuWokuN3wGw97enlSA3xNvm4/P/oe9lgB/+EEpItjmWJ
Ny8PEVF0ILU2vNSzA6VV0hdWZnlQVdg7z9iS45lxgIQC8PTsW+cLWYOMpsHEXskN
00RcWLZS6bJTmxbCa/POzOa0sVjs4ReF+05CUMt5w+5YU2Vi5DFOVTHvNhYEJnWy
qqy95Ke4C6Y/pDcMspX4TK3Dp57Yk3JejeIqvZWXYTqlTF/N/acuCWBdWNNiPjEW
1MlxFm2NCYKBcmyoSJ3fwA3252K2iHybMVV2LcK1858YcBSoFqqGIaBJ6N3fn0fp
v+Y8IhRkdeFP5EJy+CAhRNc7Rd2cIg1gE4asFP+aZKKYFJgoavecnLgM/YXEOpSP
5pkZxoFpECvAfnwGmpDBRlk/HMRg1nqeRcWvjc2MAnFMn56MiuSe7fGm5avRqP23
SD3Rsxa6c6Fezvgql/oVwL7ahBk1DmoVDh77prIZaCMOKilpvgpL7x26sFqz9Y7i
f74fctIfZ9OFPM1g7X/z0/N480ADqzu2aLwYnFqUVhP+FdjPczWyRrKPERjSFaTk
Hjkr5dcEKT2UbFTJNwVQZFu6sFWDxOyvNMu5rcwhq0a85RenakyTNxdVPl8vwt29
o4fNuyvTvkd4SfXeVW72Jqnu1ly+eILthHsub/RkpP7FKlAslwZT4u3rxPSMERic
LK2bYNvyJPWyRkvoC47h8Alu7Kfo8+rn1CxEyqRmssT2Ia9UTK3nRmyPGPC3YE/F
Y8+vkoo5eAbYQzo9qVgCrnjveErMKq1rhabSrXdZeXkqW9LiVUdFvI470OXfug2A
A1ZglUSxSXTg8e6rjBs1JQzGC2px4PW9Q5U/YF6ZsdPYF8zGXnsFzEu+adf2938+
tqAR9IyFvV0CFpYL4OCdeIdKsOcQvd60h9yZQAGQljf1GQ7404gCrHw/uo2jl6zK
rMVYmUwA1g1bsyvBF5gAhDOSdhjxULddPBF7vG4W/yMAOByjnQMgfOmngoDB1/1N
BisqXQeS22Yj6uEDVfEWSM4e7j3FgqHXaXp3XO7V+9KOgeyv9cwnwZQ69ULwydr7
yLOuBlTyPpJko6MNuisnBvCzHqolbWCkcxXgHsVrjQ/e6Si5dvHHQHyoOwN+sjJh
toWryZf7AAbhHCImXdgOz/ye7ioTwHIMTZM1r3Wyl6BsfZ+xueqyFF9jnlHc9NfM
3YdDZ5ncsBbim09CCx0YGsTnYQYA37MPllFItkjSa6qVmk9Aecta3S/F+sbcTpHL
hd1ARkNdbZ8/3gHaDBGT7iPwjIjnrLAJ6EF36CMDe9FZCWJBRYda39+2azcyalEU
9MkWYKevERRyngAJxxQF715knKQwrl9W7AHnpEgBqrWEmdcn1vdrRNRLYZo29HCs
AsThk4jW2jU5yUZAK5fW8NjmVYeXT+PLEJZgiAnrCmFhnqzqVSHXLw0Fy433UjcL
ALKiQ2nWW5m6S7hvDdHFoqgk36C7V49qlYIBwLV6NpOmu1Vbr0L5/pwYyaulvo2Z
FpZCqWcZGMVRFTg+LOD/j+irajeTKEYKE8f/DUN64lZVJAETb2qws6zT9jOMjHCi
W6PQTWhAe3iOPHXH9GhpSJ4VxzeJHmCQ2WlTkb7yGG3UFO1XEV9CNIP+/WIlBmH2
458TKlQEQ/5ktmNk2Lab4XJ9hrrJCNgCHaCMBv6FCDcwUTNKROgSpVnXu9tbRmvd
N64irKIspuUuyL/0Mv+KMrLWRS2T4qO6+J57Zgx2fTwpEvmP2GRz4vT8m6HSs4yq
UH1vFMCWnBxqOsYvUy8g59IL7f8u2QwJKR+pLoLoKEVToAV3AZTS4v81WYT9tuSB
TnyWQVljyw4oTiVgEIoYMlRpbqCNuF7upWgLj3n4cM+lQvwSM0dhtiaNDJHft9re
Rv+BCX7GaNnbpfNQAxHrD/W4cnULxEwPn28J0KJkRR6SOrf9qv+H8IyT78gkxnp2
bZy0R5Pf5nwPN3It5NMZ69H+LuOXDOGTGwT+rI7EVEgzcHnNbaXzOJA6f8+BfMM0
qTW6E8RiwK2eCoNLGl4wrEOJe1ciM3QroOC3YE6sYXsNNK4ZSq+/3f5HqA8bal91
ACEdjieKwUVsc+F8CjZAESMyMgi4R4kazo17kTPz2JV1AVMtzmpaZIJZlRna0Wop
Bi9iIAAGUCq/nHCqR1DhW2/fbV/pGIIfF5WsILytTg+jkgl0iDpKoTUEOkYnCi9H
W1/UhTocnpP5WTklLNNxX+mPaZErVd70MOVU4mvIRe/S6App3ozqzUFB7U6jhGLr
1s9SHgwqSAO9mD1EqXZ0ZaZSMWmvCc4il/LFs2FAtiFQ9ZjdZM3Q80yO7u/7NPJj
5E441xdycm0qgSubo7q5+eWE24kTsKqjG1yApYxnXGzbBxKVIuiW0PqxFTHqZURd
FBixvXEp1LEvi1PlqgASlFlAaQvAGr9J6NW8rQHbFySj+6ggLKxiM4nPHTEMPaub
zL0Tx+VPNV4RixmAKVfD5F5+s6vDiHeyvIHuHG0eK6ynUC3YqpxamQXIXkIhuyE5
fU+W/e8t9vi8DplIkcVNQajmI0se7k6kUHNrDGq/E2N6aAJmm+cwFa6KK5GhadwX
iGCCMy9fBbrTk7S4M8To3qLqjF2Tn5rMQbtwGPbc+mUHMfIpjrLtm6qAeC6TWIA9
onPOCziKYwMwDtsBMPg36mJMigRSTv7EC7iThaKFk2cqV7nZDRpeYAlEJ+6aPsho
f/ztUX1Yq0RefUYb14Iar72nEoXVZ2TFFnf/hfMnw4RxYX0VN5lxiGKAaW7RAPBK
k4L8BmrTpk85HB3JuHqoTYj2b2GSOKLsnhvl1DKCTKSiTvvRcjCAfFHVWNKfY7oO
KxU4ad71uRHJCfL+ak/8phAgpqJQuvD40HUsXyAzDX3rGuDz0vfCA7SPUf2BVknR
1X3P7ZLLk59B+ReIih7dwKbTvw+CRmT+bxZbm7UxjL2vvecFgNSqq48ehT737dBG
9eSIjQKhuKK7orW1vo6iyVhvTWndkREomZP0R/OD3nF0c2Bc+NTJdKvjqLX4EhvU
mtZAo804jGgb6xw2dVL4kMcIbcxfjTFS/ExYfujHBQQp2A4jHZ2M8mNbNkCNL4f3
Osj6eo7WUgJ/45AStOcOe/XLdiVMdp+IS7mc1cP8iJ6XbM+jrJLZkvCeeKzI8KKD
ZIW/tUwuV915bBE/UY+I6wtVzh5kNrE8nbzNowDBOTI2THK5AxFLaENtGbx+zw+B
vFrW6tF6Sqevag2muW9DlelLyJvycMMFlddkctINEli7CYhbo0bbEBKSQoMK0KFb
Wqk4qTmh8Tzlqs8HfCRIn7CDIlzGJ9VbzEju6gYf7t7vSxpcZCG+J6hSQvqpQl+n
N6p16tygPAd+XxU3ILj9CdzBW7YXn3ihcB1LpY1+SDfIMHesQCkKq0U3PMen+zOl
AlIg/P3tJeNbFXYXBOvAYG+0SblaAF3K3uMwu3uY2b7C375mOhIMolMk67cvez/4
PEXFALjBFsAhjgSHAh8efZ59e8oljBAjUFMFZE9XACRw0V8zCQ96IEnqguO90y5B
DhV5Xxwa8F7tEVJ1mk8xmToLi+T+cxVd5XDNKNz8G7HLHPmBGNnLk3+FLslpKC5B
m6IR296Sf3a7BHSJMLJIAe+PFkmt2H+nMwObtFpu4j4vgepO7pT0XsAg03fGW3jE
HInZTDAOlle5Zo/P5Xo+vbHuJ27/qMaNvZRxlmCfou5oabXCqG8ZcumLv8SMw4Gb
RGa1jCY5LN5oci+yS/qQ9y+t3f0t6BigTSZUBXSXwYtJau9QYR6HxWckUkZs3WO5
LbCqgxGYXqanw4a0dKCml3d14a1a0roui+C1xhOmxxQq6B2lJDvJp953euLpn640
rBF0LuDF4tH+695ZKFthajsLBHzKZoCibECVFfEpirs1GhoBAyEGP8fTHhpFt2uf
ro8/Af/SQrqOyLrtC0wbjEXViYmBLtdF3pfHSkV0AbRFYtP8AzTNqoldiEN8Jd3H
qE7n5Fyy9GdDJnL7RgQSKNxxVdZw9vlTlJwzFAljL4pF1tOgOp38MsonS/VfHnAI
hIVCx6Y7utH/m09vymoDaOqr/4GDqfQFM/dN6wbbhVwwkexRAh785MugBpJ2/pGb
B4wYNRKh42WXqh4CidcN4j2UCDcaQ2JeGAjt/bRyw7kpzL3GPZ9DXz7hJq/bnGvD
SdZrMi23TvIy4QkSBcScCx3H68uzrw7+9xil2IgGp7CgMM6wAvDjgVNxRqGktsHG
qORUIyqQdO6yXuaeeXyT/f4hheQGPH+6UKhgeFTuBjyUSZLcX+1TuCR6Sfog8Ham
5h7ydyYEZg2WnDcQj6GYrva/VYywaDDQpNwfB4SJD8F/OLR1AHKTgJiZV1fYJLrL
p+KB0Aw50Yi07tpGQqHfstLB/vllg3CNnQdjL1yTqgd/WFcVEcYM6/0H3b7mXsz6
fUCtLrvGmOYO9rN8eu9RrFQLlfVzoCMCscQ0Cfc605jedsnk9SJtXKLuAB+eky3m
4Ay+Roxy9oRoNrqvPoTu1NwUzVnYCeDQqH6KIqglQvicPNUWHMIhN3INMHe8G4vd
b0gOXMdrsE8UNvpF96ydHTTEdhRtDj0WMXlRzhlo5A7taqy/1zqUt2Z5rWrLDjgb
mDGSs8zd8A8lqTZqUu9mbt2f/Q9tT8oeVm8PHRngK7NWiS5xzlhWKmPXIQhMyv7s
5XFdHIFyNnJ6VMy6FPGpFLnJ/ZpQIvFkeZH7Z2Ut19axSfyTheFhrWk4eNryBMJG
7V02YklGOKEXO6V140++YabGy8jEUQhIAp9ATvKnVl/80/lgMgtkP5hoaee9FsYp
JvLKncevi2i3tOnoF3TGNCGOBrSEZCGurdJOdLZRYWUQ6ZgrdPRS6bdXJOh2S53l
o2Kv3Fdga/fBahPZbRsnDvXyBd3fRey0nHYB8m+EAKDWkMofslPZEebFf48r1GHz
zkIS3TYzFX36XI/Wb2EMOZzMM/uLzclvSCJHzCVCvEobSBudC9HrA1kmwjF78Umh
IdCcVBf6auNQKepHUQVG6HNNTI3VsUltdE9fEW7afx03XhDLNee0kCQOXj6sdA5N
1vWm742+97IC7BQl3U17AsJ+yo+tRAThhbPw7qMpWzz5plc4sKSeMsGwM+daCnfS
gw6TXRSHLMT8TRBaiZCf/8ngjjSGC+ohKKJSL4bwbdckZFvkPQuQSQL08cnW8rHh
6yYImVM3M1vQNoBzxkK/osuITWLZDh8AvmEYrxiMc//vciDnEYDGrzL7TIWLE9ND
Twrr/MOUIiFYEU7ygDNTjPz3PXTrZ+fymFEh6yqtjPf6FftVEYi8l0i754Twr1/E
U4Sw4tG7bRE5WbRUniwcwYLNKz8YAEUAnGKcdPO7vtBdhbCB50nXKHwRD4QIbgWr
6xj6uB6b/pqFkfF8X5bQHF/ngW6j84BR7XN9H4wLeAglV4WQ/8MxgWgT4X53YnDR
GhicmV36CzF3lncbFhs0rkhU2psZGnyAdExH4m4TqqoX1vNKoHDBwHR+xmiMQv/I
pRhaGO8a6ctfnpB5QNTl/NPwm6tUdfOXFYdZDdCv2u2b+JAVgREtLldATAxR7YCj
6Feok4Xk8cqSkFiUK7C3QHbm2tdN9CZdaQ/kHFojpMmwDY/WCc7pljxl6sG7VGPk
/frYjxKXVEQRk72xCOG1deUG70nDJVJVPiCFjCa7y7HBPcskR5Z9kSQK3DQ53bVf
TJfgED6AzQtv/muWTBZ0IVjlEmDsKmuuPCH0CLfhVuCdgwzbPgmOEd5LgpvDb/yF
cbKHeYnxYkM7OY6dET4ZI1zxzPpS5UQNp6Eb9KuQ1oghSnsHEgS3lkkZ/GcIQjlq
8zQQhJQ0UiLY5eHNNfPvzBbBRZFOVE5psEGNR3n+v0GVLBi6ip9ehr7rU8DNy8Op
Q3VT3nlQuEbN6uStLvP9BoEsbdrAjyONu+NoDpnk0pSRF/aUXc1QIma1kd5uqhSQ
TRsProqy70JJYQBPQZXEojAefXlUskUrJTHmSzorwrgt9LgXvof7yKHn5z1a0QSQ
MIjGQZEeMUXfvVse9cv3r+ECfIEdV4KMu9ItA1Q0hiKduA0itWTpUgTOd4qNa3GF
CEwsYJ5BX9xKnEf/s5RpcMyW6UAr7QGpRFHvgtTfXOEFIuCQF+qUXkbBRDQcw5r0
dWTFZ4/zh8OPq3ELtTC1QGUpFbW6ww60yVx9SJ3hq2fKJQ95GEJtkXFC3j3uIbx+
TSrUT0306Vwm+WizeDdSIz1JbaUQJHeeuQirBctxVn2ngWQO7+1PllpBnKPu49zY
ZBD5cOTzrYTKq+Te1BC7QJ/CDe8CCceR0fYBQUzIz1gNEfH4AJsSsuX9L8MGgMqg
myESoJ215rUo6tEQsQPpN4tHyI3cv4cZOKz3wNrN2vSP5CDtzQkqEmVrQIl+ul5r
kpOc6qra3o9tLn19SOJbsYdrngKWe0diQRp1xq+qUxRVNor6TTIqlaARb3Gn9n1a
Z20fYQv/1qSAqcc4Q9sshshUwbmb8y3wP8gd5L+PoiLzruiD/R7H932wMRkT7MxC
vul1dg5UbsO9frz/F5YHAvE+pEXJyEDHPhnOVu7Ri/CWKQFHo2j2MrbuGHJQxOp6
pIMsvwymgLb7MRqLZYFsmOQ9B3WXtxoDt8jwKRtZs4/sUhqiqZ8Zb0l3CsAIVkRP
uzTaGmc2vwANSv1jAtyjZSA6PWgZoJ7BaGOxVy+S+kLgEdy7s5Nb7QVxDdZBxvOA
4kXvPIS6WGIcbAvJzsUudNXkfGIa5fzrQv44qM4v1up13NDYYI+e/aj9TJjQJuIq
d4AFHBVgtUHRDFND7QZ45tLXILAOhH3GMYvaluCDBWQ091IKrTZqqflrYFBa63bH
eE+mS/Y4EN/UQiQg5o3kHQD8htRCj3LlZsbsMHaXznCB6fcpH80oEukKs8U2rPXs
Kvui7KgnjP/YOzcuNciE4dLcw80/b+Ee85YxkNHAJ1JdgIuz0UU1QBeZNlix3CN0
9iAWjhq85dUTxapKpExsetVzLrl/kQeG6Gmvn/fuFeFsKFOoFs92/leatN2f4zCo
im4K+YJjijpUPWHyeGJPbY6pM7/fDOdlgd2EB48cr6klyR8tpjbP9p8bcy9itLcK
4zaWAiOIcZGAMQQKxtoxb5SITwjYU0Adny6qyUbCMDarQaETB5bVBjigV2PvWd9Q
Md7fDy4ADzVHUlblTh/u+rBnDoWO+whJ4LiS1A0AJC1UtL8sIxLomTKgVkugIcg/
zt2nXfoTNQFYLVDPEUNVN8iBvyqIvklyNMjgBjtKL1ImefLYeDIC0DL3akBAOg4N
DbYSZsAxmPKZSXXmsb4dyVfda6nCC2HODF7R1qQ0DxrW4bhSqk7myATC5C5VLJsn
Zk/oeFLCz45e4LabMoFCN8hEbP/kQMAD2QiA2m7HjzBdusl+ZoVLfFzjK2Q+bfuy
w6seZGLdxL9ViCIgnBhItRs3IH/YvsyGP9xNoZwMCRrItbQRMKEVJffJOL2Ex1jk
8gEFrK2xwOrrYhHJzIg+BIMuI0WkfMmzZgoLclTiCQ8kAOEKATGwIe/ogHC3SzZQ
N9KQ1lm4CtW1D9AAZ5eE0/qZJpyUV9y9eBOMjz8d4bKQs7in+cMhBNiI/h06WqF2
mNr6eKx2w/vFV6wVGcSXYB8aII537N77kedLpYFIzD2mjfaXT04yZGc4k7pWvS2A
S584K3Og/RWT5VyGH06uIUj85ubFKV98KWYilkm4AuBB+sRMjaZmCU3MFwVCeS4W
AqwxWV7EZea1j8jZ1RXtqvVmkz2BQ5KBm9utQDq7gN9raddwZIXTd5c8MGdwUZze
1gsZpPG05X40AtWQgOwtupjcb+z8mIAXF8a6c9OdzBmEUELDuP3CDoyAQkgiipIs
II3ZEquiHTIOr8ywZ3XfHtIYNOMN4weNsqunht/JLlsmcRX1hu40a+27wTK2g1K5
WMhwIdECKSV9z9D6LQZv+vqxI/rNUuGbHEMnOGvPtTAeQcuHE9WXn0H4oet8Qb8t
2yqhVPE9wcHLasoXVuBYWIEE6LwNkURLirOsZeDvLDXcnYrs+8YT/QLSX1l3728w
bKdfilWuB/z+28Fctef6rD2RV0YJo6yu9VrqvC6MeYvSAEhi9P0p9hCPM8QeNGPo
h0qE4Z66HD+zduZVX61XBnnKU5HmYWWPebL3q2cT6ShyhNqP1hqWhvV9a6qX3Pp3
uZBDCu0xTl4D/O81Si4tbfxUckDam9OSLPCXSqXtHd+tJ3sB6Q4PJCpASIBoD+di
ZgQctfPdU3dmPDj37FeW4N41ggoSyEAsU0ZtTk250xFC+GllSKLlSeEUX0xBjJQ3
vhjeLRcvp39mGGFGwTRZKJjpsOR0yL8MKHFtpDsfJAvF0xfrGRIU4gozDg+rTRdk
K0GjSlK1cM1w4bt/L+HxV77B3XxziwCM2a0tNugvqKlS+ab1+KfFmQaC5imVhWhx
qNMTglKzmnUXNp5vupW9zqW9j8yv29GG/J0drzd0GOM5Ipb/NiegJ13lfp/jIlQr
S+jUAEY25HpmJG4I48telBM+ABAP2YEhrf+BXate7JDvR3h4yR3JTbYlODCnJfLZ
OeVCV0UrOkYNA38HIyaQIeA9MEyRidGwa900LvC6MXcek7z47/eFk1XvjMEy572p
wb0V7a81xBVhn9L+EuuEfI1Tbbuzcd6mKDz/W3ezSXgk2ar6UEDcaKnQNjlTBop5
rIMwnFKPTgF5RId8TjHs4v1CJdOeN1d/MJ3zeXRq4mI5tXQ/jK+3ibNzkyvzQYiY
SPGe65OfLbTF/IJxHexQ9UxskQtlBM6sMEakIrMLmBrULCpxOWZNj/jwYC4z8zoF
qxoZUrMSyP8INLYrazmHszYVUh9cz0kNF4WW+UC4wIlNGVH/Zj0lgV26tt9I3E6S
VE7jlBsPr0P1iuFugj66g37Aovqz5+8B0EOVmv9zA/ZTKe3vuysoyaVuaquomEvs
M22/QI/j5eTqTYnPCQAIuJE/lfUtGiNCAmENEJ8k4ZJxPBfcbSjRip/7aj3z91zP
+8f8MLLvDhFCNhVbtPpvJYE6s5Ar+Uic91nz04f8ZZkLfirBregzDXPF5wsv7SGB
KbCdWtoztkVvJ/zR24hhbkLDJ8Ub5SF1FfweRwlDVdavQcTq4GppiWTx8NBERB+o
bPhYbII0H8FiPO6Dbl8pi6DtT/QWmc6otvJdcLNbR6CC4BBQeNlF9Vdm22+xsg2K
9FEMfA4DaDy/Y/+ut423w3VkM9HwLXgnDEXc/gsSk9F/6xr1vJ/SE8qwSGVF042k
Y6RT8EJjN1RHrGw7WrVYouASHuc6B4CfqZ8wp4D4MPa38B6LPZQb1/w7tQhqKn5H
XdKIpsoKh9NmCfYHvdQVrMRqdCAekBh27qsVQxBm+0n6lF/tI1P7lHDZ/T2uesob
rkSK15ditK1x8jW0geFNdxaTnRKSrVMarn+3bqdue5W+SL9iN+dAvmKfTcqwZS+h
j848etAcMVfapembh3qwTNefREgSLeI2mgN9mJTayLKElsv+gGfaeW7WcCqouSlV
LDq42qNC5ILoSBrQWtgtysikj6bcwviRgAu30BtJnpBHIF9UPo/zOPOMw4JyBwbv
P+KudrZoatT2UE6CjDBBQCiX4NXf6pSCZ6tgFFMwSUckHYQIKYss0YiaRkjwr3xk
6dpYUMaVIDWT4H342TVF1miCyVeLSd8LUUCHzmQ58VWdg+rs2AXUqR3h8Wyy+CAr
3H8iXJWfQ6jBjNIGvxSPIMiSmLgqsw2B/oxMRVW6ou60PrfgFOx6VbwXx/3VqqtN
04RsYI+ZpqgdSd3LYPEeuiOVK0xeNJdPDAufN8DG9ZRWNWeorKM6zhwT6+yR9nWX
xdU/6/Q1ieZPoyG/FYfNh6M54wHbgx7tkSM35wDSaYC+M8asysEA7d89sn9JZvbO
k/VX77LjKAm4j57+N3SISGailymAz5cb026V6UY1pkKiwi0SrePg6a1zsKSmBkva
AM2Vkgn2dMEhSXW0Wl34kjfGLNAyiBc4gvlW71bJiuf7s3erC6tsUuITpTdEZxHu
yDfnj0emrhnB9rOqUzo7PS5nKMhgpsa5FQzpSqNJC5XRc/FBi46Gmjotr9aqTqLE
j3c+8uQ5vTCVXwSzdJ8vFwGGAZnvUbI892Up2JfgMgzZwEEUmQsZfbl+0NDPsqvi
8cg/atoxl0N+oD2WGc3RWoG9x46KOcIcU9WRunkEea223b+R29TWaEWteDTe03Kh
gItADRpSolBhIKO7sHxweacfg9mmDCTqSW+VWlmIljkD2DPUaB+a1RsCOYbTIbhU
TBRWECA/UiNEI9On4Q0F/LnO8+itoZaZTy9/vuj3OtZAY5VI1jAg/Z8wpFtmlriE
HJv7VS+TreyekPhwHgE5C7uc0p/s+e0YZ9YKlClkiULMRosvq6z7iG2fEa9sYLJf
Nhcv+f2Zu/kvCj5Be/vo+APihSFfeVP7cQxqMh7fcjBJYdf0R9bFXAHM3Oa+LrfW
o6xChSRTu3IIulEY8hmdUci8bn1BcJN4lIoM5EH4jiM5iTB43LzqfoewPGzqwoW3
mYkJtBXosL/aRssDCnVq+HGAxW3h3+dke3JMVyVeD1kn4TUW+lI1EMu1/oHQhVxA
YxfIrg87W1svCGpst+4sc55Ee7lGBoZuuGg052RIbMdj4oHJNtlxLXZAFjSMqudg
3mjNd7D/xTebPHS6/uhyATaCU9rsz6K2cVqj3yQ8VRXLgiBzRTaixP5SPDjindxw
S2QiybrUKm2C/BOWd3VBccql3am9bnluNKEpaggtbAgLQM8mThwF8iNdD4NCm21Z
YJFfzotHeaA4CE/FDFq1XMhBukEhbu27ZLnTJV1AH5vTpgezJgOEpm6qZItcKfyc
LanQFYS23D5wv28v1Rpha67PojlNo4B4iEAZnkd6j8llD+O3dlFJEcg6G53hP9Ly
JE4m82bvHm0ds+K7dbvM0+FvZAM7PXW/hVDwaBFX44XNDHyNVCRDDiMp7taCHbzW
UkapA30lpPFgMCfJGcGdvuNjV4fyBEJOxnknbiwebvKxousZfMmHvNLxiC/jT62S
LVGt/z60iUAwTMg53hZ3hFg+gNSbJuROQBJ8gehYyV0x8REsSBdNJhWj5rD2El8W
2GWNzMZ2SFjR4btUF3F/NGrQonNuOJ1dIyapXgpAESHoRjty0fBpBT1us41aMiYa
LUSYq/FoO03GFr5iYPV/VULWejNqwyfsBL/Bp90fnxdtkYxlajlqbvW1u17Ik4PG
cWp4ne/1PcXmGuaukFxTdSNHWrYxWJ5EhAU3fXc6KccZGhp1RU4BaSIJU7ZDmqQr
qYHoUYkBR1PrfbUTRyBtauHwCKfJCn286eVhI5TcLOj675UqZgA+9UK/KQLbZ4Bn
qguYj0QXz07hMXTgjSEfZ3ojaN3pnUeULnJusqAWL1dCl4ZK5HTeGGOxDE/V5vNY
22sK1QEq3caEVnjbx1WecvE9nWryv/RUmy4llqwHLjbjzReloQ/o79TQkuuJOBYa
9OWR3uIcsCLRRRCnb1xOaizsc0HZb/AqzKHGbtlgZlawMbsP2mj8yTZq68YThFkC
Oip0J41N7JKKIt4PuuKvxCEwv5fkXrPIUNZ9E6ccvqMrcTJvZCVlVfTc55YlOnoV
4mm18sqpFfpPIAFLoV74Txk7C28FSGIz56j9hsJlzZPk3Ghr1leUpW/EeMKnLOP/
q+MARWORj2inJO9BcF9NTfcUezxjBDZsqs7szSNQiW3sC+fC6SA9KwFVktMo1BYW
4HyQ2SUxYXXtqV/6EMNoPyrMjkP/DmOg5uRbJse2hOn2/Uy8SBUTyUmHrlBtf2Rp
AkVMwIgM9js+HTuNciRby/nsy/ajbIOblbIWoSE9QsShZ0PGiyVfrW+W8j08c9Ew
Qi61Tqt31l7TJ4cidHFDwlLI0eB7CZOvNJZ+9aIANTB7DiIawk89ZEvqHpW6FxDU
FKksU5ZsMdNEAx37Lnpi33whwuYtzP9OKb/FlR9Ss/O/Dy7wMxILH+xNW5RQpiqM
a9bZ5fNqQJ91nW95AbGAfQoiOi4kmRuPdQwvOa9P6DoIQRawzODWC8m3scD98q7A
+x3eAFpTNAwnDFj8bT8CxfJ6p/2rNLpJpn0esoSTa+IjtfcZ9QL6oiIf/5UV4rDF
JvCC41NaS0jyuey6MsloxJoT7ZXdg/6bY27mebTEOcWdkqnewWBzMbAsvix9nQ9X
rPA7KktSw7hB8Uh6lSDxOWfbHmyEWlr9DsEn9MD/M1J7zDgZKwcbtf563av8T1tu
cYoM/FHKrgNdDXQ2LX7oCj8zf7P+Cq9owGZR0z5unewnOYlG/MJINNoRzWvLzfEQ
9FtQpMxeaJOBHGjqVJV0BZ6vvtJSqO+fGMK0EFyATq4xEkfIVtegWFgaK+RNhdyO
jv68v9aWdF9u31EL0Uqa/ENrIUdYD8EmZPaDkAdEh2LHux+JVkVCU4oBKQywoc1w
8xv9+8szjZYH/uuSx+c357F1bVjlRnLOAG7lkzwjPaI5s5SvTguwomRFtl5uMRKC
DrlnGBFhRFMCD1IpVNrGNweAizI0FPtjpdOd2dmw2nH7/vcZjbRFM74m3To5y1vC
aHW3Ac7jTUaYyPYJrUng/qHUWGv1WgtEpoarrkKt2s07xOx7qCrlguKIJfE6j8BV
pTQxNFSbRHGVqfT03TL0qqYPBseCvJ9mN+1/l3gy3/2+rwDbs2Ct7H2BGhzal5+y
huZLOtlhzHM+W8TUzpj8imvt0CxhDpqDD2B9gfhqxl/r0CcbckrmmBNq7l44vULa
V8mRiqibTRWMVEl+uEosoIMA1oFkuxz8WB5fIhuinQg8ugXknh+VGv9cmO68+0Xh
TyhkSNZooQdbg4Cw+USo+AnflfyB5/UG0L9B4h5CC40lwtmdRmbYQjCKVonWPBkx
1cwm25mfK6LgtqUapF+KOBQK0VDOs+CdGSmdvXfGMdYeOTcybKa+aqA5mkgABe8B
1swPouXUKffpwVZIUmOPZljgjndqsgOyEKWMK30pmSEFCJBfCJv+yZCwEuHCyEWS
ABo9kgLiKADkRpJ69dB/32TqOcp5x7hKssxoEhZM4swmU5zYl8TBH3JlOfA2FfFa
OS9+gcqz+zn8V9a5RDfZAfdae3eUYh0eryvqq0hWCYT7YYGM1LyrgINFyT7oLzL/
lvN1Y1PtwwvXaij3ZgdxelEvVqVREIpVhv9gWnPBkrYZfZxSMtqAJ2bMf21BreHf
+AezLm4zm1zTiELoe3lxsF19ZtU90Lr40s948q4wv+vtjCcOvDXE+1XapKFhEmLg
84BVotjB9WSyQqbHpyozAogWsY+IckJ466Q5JXfPwzcrUICssRRhnlDv368KLtf8
+jDyM6oKlNEX8U+sUwNY9fLpTIeaSc5FZGlD8Sjh3TcddU9QPXgL+g4S6P79WRc4
yeiXPmWM8rQm8NdaYvxhcbvu/jr7MmfxLL03g704zcgm58r6xT8mPdDpCi0U4Qau
763XERFHVQmjvfTUB3K3anxxE6kAKASWo755eMguX5mP4JRW6vtvAQ6SdBYl/xij
NcA9lu3DFc8yzQ8eVQNqXqy5ICk0yoNevjCdKLNybzXhEoAO2zjAEi9lij2m3Q20
TcMHnhlIoYJuXadu2O0x9t2O0R8AgRZsVhYlgReQzespuWa24TmfUHPXnPnzHrOR
02IDHw643+QtcsB97zsX7Ad9gKN+XOV8ER5QbLHAXoiACltFiWcFGM/8Vpw91jjU
04GAyhFJiskeEudsz8LIqMlcLtS92Mltq9IACbPRWmXqmJ40/S4g8HrQa6TN9HPW
1Ir5J+d5lhU1z2gTJVFV3vc/Mt8OrExNFth7RHmS+zcf9fukNRpFXGiWaoQ6oRD9
aAUT0q87pisSXEhOz/+4ZY+gE6X+wRtpPBNnZigFR+S3fwkTSyjF7J7PX92fcrw0
Sun7aXg9v76xzLmh1HAGyt9wecKnohSOcdkboVsUz+vTd4rFBgfjiI3XZMYsYKi6
ArPsdwuG+HxvbQh9gtkWsNTO6MLBeQvjMayEpB2984ZV0FYxXwS/478C6bv6RE/D
N99zWA7q56KB6gscfFlZ4CfS0NyA9Ppmervf/c/ajraxPZIc9KiocSGXAQ4uiqkJ
hSilqlIJcUnDTehwwwIwTCuDA5qEEzPO49onuDveKMzmqvUktnVFkt5uAc+1BvKo
WHSuX1/vX0iALTHqbOZjuQGmmSehYBCW959ZP+eifGEfoP56oM8Yfo2nFiC7yYcf
7Zj6wsLbuvDoYCV7i7eDlPTKQM5aUcNeXYYRnOZ7+MY0DeDWu8vEMqdqxdilxepZ
r64lxh4a2bT706L8EeQHxn+0ag7TyZQuAYeNAwLzR+JORE1NFcT4GDK50O5lBXxm
Tou8NhZbtWbaMYrAa2j0gPoBs4rE0jzySzz55MNqZg2ffYd2ebgIKHVh6+HucVge
pm1v9QYHxX7au8n/MO9A8DvZteWTik5KPA6fyHVsIjiafqf0hhyaNS5kb9P1JWjs
qNf3VU9CNGSmYoRHW/vrae5DWQL1Tl7k2JD666XxsRxXsu7GjK/rXMhAUZ2AxYaM
4EnbI6FsqrsoplwgceDsk2+1/fp+9HSGw3UjhEAI/XNJ9blWVkKDJ+pUsffCEnrc
OIquDTa6q7RadpCjtHWPdozfTdQkjdqUxlkoDCtaG8Kxc/8gVY9RwTr9QFBpEIYa
HsKq88bkdJmp6/x0GffZCNX2RguF06vgGq55rCSy/IPPh0uxsShgC0kgquv/fo4I
CXL5XmJBTNQsCokppGHsILD1WZSFdLgbmzr5WPBeXq7k2FYwepIMNXmvF1y73lAQ
dXNpxOHgA+cmSK6oZlxBaSzGa+5ebFBI279RKBhjuPUcO8KK7zJLMUO+AGiouFak
4UGAuughAMX7jxqOAz+p6QHdU7H9z3wH19wGrz0Sksn+V/B3RjxF8khNLqiwViir
wjoMTcMTr09EIkPJKK1k53utkvFbqlTw+L5VwqodWY7t7R4zALca9PV74dkTtw1s
OK8xp6a5nygfLwcKOHq1t5RIAbKDe53pXIZ/qp98UWBUQxv0mnL5oFVv996qn8fu
59NWUgZpq+I96Yd30toGWVk34cR4N8VMD3JxHzjQTohhP7Cdcd8oSVAiz4IfsxSE
uLJ+RdlX/zSj5JC9lifDh8dIRQjz0zOS9XcGupG5KfJDFn95ftEWDNkZeLZnN5hi
F4dVTkFwzdMHm/b09C1+wpKGWSIxbVVp9uSMwtfZEwsC3ysG0gX4Ik+c1tBoUEWU
zvqbuR6eErdhXAx1jzcKSz5GYOF4FBAVoxBxtoCFvriGKhvcN9h9kcMFhFiq+ld7
CGFGedCVlAqrikgqVTohRHhjxeV9SERKnIMyB5luhUJLOdgch+Kkfv1wPwAhSCKr
rFpUeaSXp+u0HL5g0VSmBBL/TQL2izwUV2Utbb2qYU70kwW2Z90I1XTtt4AFb0r3
u0QVRfHgY8P4B/7Lz60/QfbHT19r5fflipFw+2zOYoeDVapvQKMLijovE7Y0xG3c
KnXrilmUNkEizwb1aI3MybCUPUg10YVCA6VjI+M1pjQko1w33PhKzfRNo93GJBia
f5MQ7Y/9WeMvfir2bbJBI0hcInGCjBunicTZxjZfCztTC9gboCyQDETUPv0yG/py
6ReoRg82MKGzzA7GUNh5cL4rxzESQUSTEoI4ndsfrM/zV786HNl25AQA4RrUKmfL
+xIurpu9kvXuj9aZIbG0yKGIZQQLXbHG4l4U6gol9Ph5HCNNTmZqkNpNsFkzmQF9
03q5dCU463nAc0VoPTLHqmV+nENF3xIjOLjLosEkhqj3jv0+xOzPHO30XpyUamvM
EY4Ca9aNiU7lQVzXgwlvTDAR7ixF613VBdzto26ufGL4S0L9BS8+PvG0AOsXho/8
ipHNsg4/NgL2ugMpQ18nYKjBf5A9jcHbWtHWLqHAFUPINyxnYXxvcnTwBHnmUk56
JMNYxiOBFQCY7wRqvUQ5aOTOCrqRRsvMUMh+xdZqKKfPbVqPar5Mnne3RRQDBjqw
2sSQRpVM397hd9GztdWSgVk7l7NmVxlVBagZ+4TY75Zhrkj4Arok7YRzWmKCfQfV
yZEcdLpEsC3vbmR2/NYnVSIZQfPCSmBcRCP/uULIo2lLkBkWldUHpDDFKfVyLZWi
gfQevRvfjREmXpZEUtJGIVnhADVeSUhka2ziI/TcEBVoB1aw3jH1X/7itm6iYr1U
JxCH6qxbPnBxEeSC6INBjHQwpRQ6bt8zuKr/UacTt1Pu/yaG/H9CMaQphFS+QZVA
ya5KdUR4PZ+UsHS5ImXZo3nsuLGLZOkmG9KVFmd6cdcPwagq6Pc/bw7Q+mjv5men
JRcsDAzjvUnI1LP5gdDz6OS2TRVxX1r/PojBxXdUHmqSaWpBRZHOf603/gqMpJDl
dhxcVCuuAmOjAbV77pO+qJVbDb9ppdAtjd81yT02GANaii0Z0DNDkhIjknbGgiyB
4XSuIaG1IjQhJFBPSO9WOqxMiZTuSDUGi6kOUeu25CU1IIkzZXfbbFl4vFOr8qgf
XW/vqGA4Ir7KAz22bqMEYt1PRSB3IvuH2kI9R16XREUbtATKoR9uc3+IKiJM9ybQ
C8qsl+KzuyApv+mk39pCA692U98oUfGpsAfUdW8PKBzTUe9FUqX0KTZlhvnTpemw
cgoGG6L0SslN45RqrCcxcvkjQKmOEvsHZtmqxzCZwS9c1+Q6QRQfWMRRtdZ1P5Bt
iOWO66TewtmEo6XX0HcEhztOeC1Pu+aZZL5GiC3eXeVvXGf/OEuPfQ9aba9m6trR
PYpqG3wMYEKRLQChg2n7bFh/DUfX7DrJ9+W8cmlE9MPVwKQBGegVa3i9BMoMOGL6
J+TqAZTGKXh+t3vLyLREWZEBmtQqr7xI9J1Lwix7KwiqBwzqBX02TjIDs9gbAcaS
66xI8ffMxjX8iG1uPtSgbpLUu5dneBn9tITsKtItlsm385uFbOnk1YCcRUUx7bVa
UgzX7+ov/9Bj95X8pHg/DMx0Bv9cyf2ft9S3VmIvj4hkpg1CbBuRdDC59Q2irBBE
l53Y1KQdcQcBKdIs7fLSHiePT84HVlCXA7PPmwaD6+nz/WLhpOuNaou4jURFloDS
2UBbP4PlEtlivmDAPAEfJbEMA7SGq4iOhsEfcRLlWOmKbbpQhCJr8PwWPKWASLMP
f9V1L2/Heo/11ugq8iNd31fgv8aJzcLnlFvlUaiC4pp2hDvQJ2G3fsa1Ie+EIZ/6
xmnnKfpMrH/Fhhn56J14AFKSivKbpltWp447fwDgdwiPb1+7fTJLzh25AXnvstk6
hgQOhfS6ZO+LOnM+9bqXXUTqkDpfUja2olzdhpiilyRI8rN3O7kMKkv2EbGRhPKO
ZvPulqWUWnv4TmNfBMizChNlY39YwOaSLkClbjgv+wbbrpGRZfx1Bhb5c7s0DkVB
NEUWrgmR4fBne745DC+VERyLnO6CXOdJcXi5BCI/I9vqBlovPD23Phq1c6Q37z3o
8G6jx+JxJ7QCzma/EmoD8xrvsfnxDYhqkv6iAhiMtpM1+Y8C6fYgH5KGSYtuKvtl
ZI46PgmiCATamLDRYSL+EgC0qQrVwnHXz9sXeNQARWUBK2RxfJNqnCGZS+qVc0mX
BG4OlfPraU999N4lyaCUSR0RU7A+ecQ3/kYv5TAEbuuR/AeY/n+3IrB87o6JyYGe
ZMqsMKAZOfVl8Nmp9mPURK2DznO0U5NzBe05lAWpEP8k4Eg28n0E3D7UNpRtp0Ec
by7BmJNyvX+PGUO+w8KuPl/oJ267ZP4BKm5rbQ88v0G6ejgra68G7ZYVVj8+TgKz
VUU3DJZuv76D3s0JBeknp7GXZ51ll408BSLELeuYRn3guJbLcTs/TSoTZ5kcbThy
PcYy5rZw4MQCOM3auHiV+x/AA1W0/0VVTzsYTJbSTHCXLTyL2xo29oz8YSHKkZ1T
ZHCQxBzH3b3cd053gYSEagem/68DttNMUmiTPRL5JJE0HeB9+kxF+KUaaVLd1FYa
LJO+betijPt+/2iGrI51Sz9nFey+Vh5ux+560Tf2uPTPJX6qpaBqfirJsLi4Wa56
xs0xEuRPKHNY8wUcj9Sybb3Ggxo/Ke2vk5PaDItvm4EvqfU/8QZCjTBpSm8l4gAJ
1TjZuEGvn7qFahkOnADAY1OfEt5RXxlN+OXVkqQUPeXyym/zgo7uh9YqxwaEdRWi
I77SdX7iMSxTtlzd7cNEvYRY9TBG3iMR8R7ZCcKluQYSZOw3qb5T1wWtfokYW8MP
U9/p2a37cP74ziRAhzKmzo6GD3OSyBVaLyBKBJ4g2BWiAOFDbkCeVWNfe5Bj5ZZT
ffeOVMkdXNhlL/mlWDHFrxSo/82UglwuOCXiuf4VHnTKw8RfYo4Hb1Gl+gdIfCTm
pFA4ClkpmKkcK8XvdK3QXIWt2DvS+OLV7bsLcGSDTlY3Pc3eJYBSVArAChQJtVQu
XnzwXMdK8iKAt+RDTVxcwghTBRibYV2rqgjAtiuCTxhC/VUGE8wAIzVANmlkH1qJ
9lfhQb+f+ZsIJBEsy7cF3gFauXdFrz4S+pznw8jP4mqxi3+ET43WkdlzxBkyARlL
C4H+kpB3s/V16/BG8tNbvkUAFTw2WSmqjfZzSUOfMUHeSpR/dlrjpEFPnhdqt6bD
1v15j+9m8TR8FTd0tWgYwXCDs6EP51mJwTOG7k0tFnaqnMSjauqc+DL7t9gMQ6qV
6ika/2/bxpzgk516deRVEqeEOoeNbx11BXboj2whrFVyGdE6xk56Wq5Dcx8Ut78m
NPlaRC3COPwx2/XNLqy4qrZSzB201IOsKejF7z1vPTEQj3bGaE27F1/WrSmaiuVt
6INymQLzzy/lzlfVZQ89qmafSqsF5LJele+1bxOwms5RnpXsOAWX9TcSseqC8RNf
KuM/YWt71x6bx6qxBZ7WJRCihcyvRzIzKL0/P3nOmOp73V2Ro81+S2uAhLv0/lUT
RQSNJE3hcN7oxMUAkf1CxQOppyQvaEjlml+vwpnCESzr9vAlDAgK28bcpWVz06Ht
p1pcZm2kHfOfhlYGJOZUmo/ri7SMF2LtpA8sGfZbxMlUg4+9QiX9JkFi/LoMVZ8R
B/zsdzz/FAfQFO4xtHZBGiwhHLGVOmvL/joCuBn/TOm11pJbFXR2lkDwrq3YOOd0
uW9a3+jOf4fSReyCEAN308YPul2xc8oJHDIJJUQ+CIpxTN4gDtQChPeACvLndTxP
spsYqFinQDmDr6go+9WyhJNgfH+okCjTm5ttdETti8e9QdK+tgl/2jTvglPMQ6uC
IXjNIc+fs878pSz4GbHYmnP8PdR5nQ/ricCtIb4n2NtyLpHgPvcEwSTAWOxSUUmc
f9xN0R/5r6430MxhDpt2n/zaNnovy+VX61G2cNrUIrjuZy8pMnPEUc6QzTWqBAFV
iGf7xR4MlHW3KMxz4iPtrzNSRDCcANyCAXpuG2pedjNDTztJcnCtSlFNuUwp/sih
VXwoWcEphIQVm70/JMy947tL1ikUOFtaLfwHLLURv3i9QJCimzyhlSbIiVFFnxDy
X9flGoYMqOqx1IfoEWsvkV5CV5lL14JbG5kgkGhZVZ8u5L26iNSHcFjKsM5XggXt
pYesIu6AdA6b31pOgDhDqmvBdYHsuf81zyApu4+EpFX5RHhRCfmwFTgngJmydxSf
TiL5YCZMCjXTxhNDA7HfZENcmwcHHmxIqZ42gGPYv8pvZz85UVKgX9/pK+nItmbD
BpUH1qzOCj/EaC8L5ENRxw24xvY60447X3hqb611kGaHl1rktsCwyFxZf/731KtL
MJiPJIy8lhPPuirg+3J1Lpy5HZ18TH7kf9GTcjLcSqccOFUdC/D4igYM4r2DwXc8
kENf7wx691dKXjuDfKK8yGb6LOGKVBezvj8YyFrEsLCWpM93ewZdcackxC3qXojV
gumFVwtxrTVUDODVhyRMZlYlQn4rT2op7oWp0m/MYJt1WjkUVPnowvgfqADSKpV0
U9Ut9wuhn9k6r4uBiGcu40Dq1sEkpraDSRc9Rsq5MKPnLNd/ZUza4Vr0nSHAJb2S
45k+SGS/9QGB+d0/P2Sb21vgLlvNjSLlgvkG5qmufH/BviBU72xFSKQayCs0pGlE
73z6LSgbDvIckni0WUf7/y/h0RxcXBAdNmUa+r+PHdnKRZ31yeIThru4xANEw9Nm
OkLnIZoocFcgAelCj1pau605sPXeCPKcHx1s/iZKaekXKTc0AvCpVh4xDL4wFaJc
jTBHV1FND5vPU7cvEx0XTeSJh8OLH4+mfwvZUkwo87uLUXzRstRpe6ap93DvD9ZG
HCPb54dnLKk85FjIwNgWWiMxDDrSz4FePOwRZE9Gpqvct90PqmqaKI5Mc8FfLeIG
3OEYN1dnUwZ12MSo73RFsF7v6zrHJOzO9Yh5mPUQx37VUb+wvpiNW+noC8aos+sw
O3h0mAKLzwepdu0nmibJpy7E0UOFU9f/jdeDtbF0v99uk/HYZAkwnWoSX340Rv06
mCiaFx2Z2RdsG90lVHoPfr3DBFVZzrtSbR7V8qfHRiT+XNlXQ2keylqhnv3AkMFO
6HovlQrs3yDpT3l+ShrXtJ6Nb4JIqy5eY22++HXTbqnkfFhBZKddy5IJH3vwI5CT
hn9LbW1VTT1bIvZcy+ljK26p/US2GrHeRceQ6gaL7aEjfvZT/wgbRVlaYMyZWso2
Mxn5r4uCg/pCVdYqQ9CizNhzTOxMksyoTX0dIJ3J0xrX24++vYDuNKbyZFVOn7ZI
35MDEzcK9Ip3bNH8cT7W7LY0/b1CMfdlDjXoDB5CgnWe9Q7sjT42GmsWHgO76zp4
M59PmnofMVtiU2ekRvZkNU9jBRLtjB+twM3aVnrgZq3rUet4y6K9Twe28hqDFrRT
E+7Iy9pDLThvdqJuIXEpC8P3SUO8Jf9/fTMYH2DsyC2CavDMVYI2ExX9zPDnn1Jx
FpbzKXXiSvdNeQhgnkkH7v87Zdx4xiY9P86YE7gyZB7WjX3oGPg4NK/Ozxy3DvCq
nC9EtMnXUUnbPVvL7K7t+pDYJVn9CIG9kHMgcCCPLl1aLBDUEMfL65sQJFZTog7j
oNn+9CPOR9zxj2+p0O+cGP3PW1J+FiOOdC4SQbPcIo7dMwS+pFfwFVBklD7u88bx
3ugxYEwY2GehFRWTnMv+12zpMxFAzOXWmnhK0a0tIfuGVfiLxiXwTawYV/1mtBh+
tncIzQcGaS51nxwpi+4c8sWom41uYRLnQ9q95Jlb4DBCnVT7j5YcPpZswwjqi8Qu
bwX4kqRYcaHpo8/EpAjJ9haYUI/pUHZe7d6KAr9XEkoyHqgtZ42kVKiSOSk4HB4k
NeFnfADVwd2+flNDOI2cd8AeKqtDJM51ThvI9SHnyKDUv+tr8Ky93jjSOtTtnEG3
G/AH0Ktz0LA+YQEJg5gIeQ3nUT1ajIBfmFzV66bLuwEZKgSTYWJJTO8JANhsKFN1
iW6gk8IorRJRqVe/svqUbNRdWbNYzeBbUsknP1RFqqRLs6iHN+3VRPLDt7EYrfG0
XD39ApY95/dPRArRGrC229t/O6gbAQraUSPAyWVB5wdk/ZKu50Q1dxj/3260xthK
ugs9Z1x6x7aAbaBRaehKkQDdpcQGMX2Z0F6wN/+I6D9Sqw8CmbVLbvlziZ8J/C5a
684PK2nJ7JzV5UvmQfobdac7IcmMbGBJtEhXFjchFqIraxIpffhEThKy2UmlUy5N
PvSQxcTG/CJvg/+/tj/AAqAUwDOOBpiDyBj7weTeJjjriw/akWmV9+k6dRJ5udwh
9P9XqJCUmWLTaX7nJspbYtCNBz2v+jPW528Rf5Xvojy/vLX8tyKNyvxLSnsacfYK
3DMBcJLb4B/KE36ImXa5BDYrTfs7xO44ZQ55FQZt2EiIkqzz+csfUQhTiiEhMcrf
XJYfGhmWB+WSn5Yeumismt7402UjTpuTXlXPPND6QFnaC+++g/RDuBTIVYSi1fvZ
VVxrWZDBHfDjVLAzJH4YKu9wsSXehfuIhkKxTj6FLE3bkTfq6M/JCkBH8Aji0Jqr
U+dI4j27jirxcN++ZzmtUw/5g26aBa90padacmXJh0MCrOkBqW3S3Zj2cXzFYc6V
EM93hNrQO9rGKPzSQ47xhtCE9X8vrrpQ0RI48P0CoradRg997UDHr0JCRG3E69RW
iNNii0GkKiV9g4UizibYgo4As66zi8Z5pZShqRxftLuqN/wA0ehDKDFKu+mZdKiy
XfAWUqBsODkZ523qCNxstKWiLNssYxhNHhSGnvnRm6aHtgDqh5qi64NhiD26kFar
Jdyqv89bMH8HRb0hE20NEYjnT8W+MaaVm9MiPfYXFXrONS9jRyiYsl9DeO/YK8VM
w0VKGopZQb94nKw+BMGf13YR77lcvOXa83BpfVTXV7/kwZ1MUo8ZCbp/bu5w/niO
blot7MhWJviAhXyc8uHCyyT9kVSgR30+3b0VND5pxX3sXiMvclOBai0in2a2w5Zb
8q8HhVsHsidJDj/pVC3wrSGq+EgqVEhg2eF34eAvJUbpKtXhlpa1eiH0Nf7fBJ0L
FteYG7Ap0trHEJZDxWdk7ym3Cqkpn+fY1jRdsFvYXvm7jLnhdz3qPUNHL+p9WIF5
xpMPn4LPnKgw5Oy2yKcHc3xy8NkTw2yBun4cRCye4sYjll+F0bw7uNC1Su+CbXD7
BXzFwEcTew7YXZ66sdtpJC5hj+5Npi4LxifrdYgrxois+xb9bgFzdbCmDsxfdSNa
KY+aqjB4fAvBFMVSfWcr0idSx9WkjM0oE2fj3m/W/cNFU2yQhK/NiPc56G9JVvq4
D2qz8jpt5Hw46swTGbaab4U9UvM4oEQLmHy5x9DqfAwPt25s4SpCvMQ7nRNWh5F7
wf5eimSqDVd/FncN5QCfZXvbYtEZ2NrVGH69CLXLPW6vkL0YhLCCr61eM70klk24
eBPF+F639tbPncPxd7crXdOnt3rtQi/WyoaYbvwEWNFlcceoG19xUbAe/JLr5+5L
De5Qv2RT22KqbZ0aCihQy5CuQqwmV9afz2Wn5LbLUrujR/28CNSl8xb5zFE/4+V/
Xc4wh9+XNxPaDoM1rbeZsCaF6XodfcAQpbICdjIU/qxs2SQZydQQ6KGBCYna0QqY
uaCoHPuy6sXTt8pBnjSKqbPnM2dCyueQcLuVSjdkfLYZS/JwN3ZqmzufDjS68NyE
b9cCaeQJVptH3QokfOiVxuUBKEXBWL9WP8Dm3viSjc14zl3MF2/QUxmeJrziR/Yv
6MGYHcMVf5XJz6ZaGKfIlQSn4IrglXMuWvLx1Luwz312WlY/DPY13yDVmyFJkN6l
eR4y4bxIMTBBR1fat/oMPN3teQS5GvLP9E6YkOqkEC7aD0/zQXrm/Pnz0hQTveyr
0SAJActssMkiCAF1xOXbngSnQpxCWckWcZnVeYI3RRXFC757pL9ZQT/zLEfdtR4B
vk0OfUdd1dbiQqyevoehx2zqxRlJ5i2QyItl8baWJ75HX3Y2uf1whFA2GmtuEUvn
hbCZNTUILOgdcjTZSn+rXYhvLiZAl9NCnw3uHTXAla5a2Hg4j/aMdp3G/WndvYDj
N/+haen0N3keDyJ+izh8tS6z6GRMTD/fGL6jiJqKcZjdcK5N/J8jqaflyMC3HUDh
CzH5wFRRDH14tv3RTKpOgb+z49cAWF75iE7SLtOF6EtC4OXxasJOU4QfTqJAVDQt
HSbHFvrdxA+va/twZyT5qcUL0gaHuTvVAWZm4CZEbxXU8lSZF31IktYhr1OgA1D8
d6yA5ezNmIv6gnGvS208X/QNjjb/G25SMY++dhGDG3SmxDfXAjdn5GiGtHWXc8iZ
TTbYHvCCLQtvmvktj1s23G7QBP8YND/SZHZ2sYzXBCIMyaKAVub47Fe87ttYJntn
r7KTYSarJHUNWE8TJkVL8sKxMJLL9v7XMmVME07Pzc7YoUhIxjpGjj4ycNLINHhS
JuXRsNv3TI2l01/j5wp/MMJVeqkrsYaahdf4aL1hPacVusb/zddmVQ+xkcu4fWY6
dE1exVNijWlT3vZDwqT/cRVdRsOhn/vpt18/Dh2wQ42fnvLLqHDtcATnHbOO1JVE
Pdx0egS/UFsNeaQ12DyteC7T2UdnKnswhnfMXBKgjuNfCkvcaMUxugx5Powdpr3x
UDe/qhiqCernTc2NYqedkYg/5jwjAfw/u34O9dYFbO+YnaP/BLwWWMSwSv1uYlnA
TuyqB2K++taoMzZruHXJnvKU151N1hkoT1GYokMAGvZrgJ8lR28mvkNOZQXFfahH
6x9Yd3a+oKGWO9dvTyFaciffUKoBOYevEnld37O2nRMicE9yVWcpr8z6LrAQ/7lC
HYp9lVGN7AAK1dHydOkkLMgvk3Ic360Ez6XsA1Cad/LOOqqj6rXN1beYmqm6jmns
glhHAtCbrKEWdvgpA0x3YrawU8Ybvl/thqxf5upWq+l1Jk92SpLensvAFjxSwBjc
Jmu8tJnNOKR+H+joVlMaPGHWfRWPoDqeJwkopuaarSpcTUOhcBqc2k35vjzkXAXH
rflF2LT7oXJ68d/5mmp0XzoKnKWm1udiwRvKTzSSCoQ1hfksZzHiHcRBJrwc4Nrp
6gfMm1IqXElf7+QmGzbw1ARf8GAA7Wit/1nAea/dFBPSsJy+BzR+olGTRDa9aPAM
cJwHZ/+/Yi77EFkZN7Z4HVs8GksyJ2NeY7xyoQcOm70hMx8/x5RhAqKWJS9uipIG
6yiVCzZqvkjcfvzdp7fJwRVi/kAdv6mhz0cTFdNWTaiHNfge9bN0yvuB3PcqODIB
tboBz8qzLQ8oKdbQ9wjYjMqsKTjeN46gFe45pDVj+DXUNa27GCDgX4v7sbUNQOTb
vlpKOOvvEilkwLBviDxPLblpKwg0E+D1ZBFTrL9+6/jJyZ4TJ8tPYOyOMUOpfQdJ
DbnPKOfepDwCkrqg6UxewZJ92LBA21/3T+MvA6WR8m6P6LrxRgjSq2oi+807nwrO
dRYEfQKbta0Bj+qc6Hhqc7kt8OJu9vlwWAJQDk2BZ1mQ+Y0emlkS/8xw9eWfxazr
ysD6mGnqNFS9n97jQqiPx+PNhFEe/qCU9yB3G4dkZ9JN9rS1Kqs8cNvIkwglj7dF
ki91G7iwH+0UXfoakUINlpVjFZZ0zXsQM+RfvISuCOlWNDDtvHH5/1kWSqc2H6r/
wCMg1rvQN9Cim1DWLTqPPleuhMKb4vEY1mibs2KscQdEumkUSFYGW9EiwvYcH7K6
2meaBz6X3tcH9eGS3Lp0XNOiyL9fsN6AyDhrNjo1hvapatg+icf8Y7OUmenpVkpT
irQFmej15cVdzmobQ0rgCIutT7bbw9SiyiiQPLYuH7Ankk2ZgQMYICFD/8wAQNng
up0kjGhdIsLIqpd/8hAbFEI8WuNk7CCar76Zd23eoxoz70tyXH6Uk25/TRXyT6fT
RgZMt+eulBlz4RrNLmXVNPuGOEKxUGT8kc7XKAQ5Z9ow9x7AbQkoV1QS75rbKqQc
4vfRfmib8e4Z3crObPJI3Gl2hIwM2i5292fz1jRJsqkXlB2XV4eV2Vm14K7CkQj8
rHlhcf7UDZm9+qVz9ECxwAoqnMVspB+bhvEaTq4X2MSMfoftC68phlZFIh6JIIjQ
clin5n+iVT4q4qMtry6ih55EyuZh83mMw0vqAZfUUHF6EdN30Un5fwIW1qdFe1Rl
tQ1rtJJcHFRPTQAutKFCL41fll+VoMMIMUoEDwWmopjg6uUQPUWNRjcUQFBYQ7s9
bpkuQNzgcuDYnVbwH76oQxcRKphKFbyYbjuSai07M8+RLqWYUj4sXPT4yz1QOl+n
4I+czMhXmF3H+UjAq8q66/URMjbwmfGiX4CQlqRUg20cTPHHaAb6LyKfOffm2ipX
ezfruWHEWQQ9L4BpR3GTTCxTMCmuJ0mI+2RxPEOaDTxwGoO+48BGvFu07en61kIh
n1PBimdqs58B5S86WSzAJLr15TZqQvFgrshRA669hfQdfeFFJew4j5SvOpFliEXO
UtNIHK8i59UCx9ecbNQPILkJPZujg9Ib/k0FBI7w/86NRu/TE69zsBW3mYCsfWjJ
IIJS6h9BmE9CivtqKu6gVIvk1Y1EAYltzUuc7QVfYE8HQaNgKCHsks2sNCqXZtih
SN79jjYIMEjGVjsZjLSVY9PCXv2H0hclZgPdNIy0YHdA/xr0ESvIPLyDGsaJfmOW
0thPMP22G/I0JyxuuPNPLLQqPc/sKDmgHtQpG+1j6/bpj3HVNxqCjiiq3h5rBXd/
pLr32fipOb2cLJEYxHRl/auAY1xWuetGACBc/wySF+3hbP6esBUoQVdc09lKAaX0
zGkgZ8YVgGUwnuHcsGp3eOohzfBsBJYkUwHbE3TvWVlTzPuDdc7KQM2oihirLrj7
Kdojo4urdxRORvjIBlLRdvt5rTLdtCuOwUPtjC5s3BiD/Fcy2qXviU0z6y9RR+kP
/uBZKxDxIfsLHJLBqC/a0GpugU+cEjvfpfyvmbp3jDzdSwOP0ngDfAB4RTUYEKYI
NUSlFxGLIc194zbRj6UFU8KnuUTZyoNqFnZbst6WAc+kHK84eh+5OywKKWbXozpU
41TcvtjCR0fEgYX+OMMdebLrPGVuNXBzkVJ/rDkyqvrNztFYWOPLJ8Gn947nGXI+
A+bPC2u32+a4mZI/e03It+U9fu5C3I6rUI4iwCuFSOmfHSkF6fYAfvQai/Sq9gDS
3+nsGF14rnMAeC310X1gwrnmcuM//PFnfbMxvnHearSzzg8J3BECBPVIebDGD5ST
XdAhBS//zNcLT45gjCk4pBvvVTd/8pzuv8d3NbxMHCshaO2y3d128dUplYseKjy0
/Dn9i1nO6lmA4I2Lbf/TxB0KFvVTqEzOM80inXRlGY/EnyGM97todeENmdMgM9aD
uhxgsgf2ORUSRYL1vvLUgjHHVOv2jz+QMLl3W21sG8FplGr8bQW3RagLsBLeQtFb
N1EiH/v2vRa2h8E6mu85OMJP79lgEi66AS/cMz6Kp/Qrb0nh51Zn/GWSudKr8dJq
O7FTMMNl1z6UXRUMkk/xULQtoG1ST6KCQuhVoOZGZemlY4+n4XOu0xmAshUbbBS1
Le1NvJhF23/EMDSVd2D7fTaDHcl+nSiVrH9tyecBlzJ3GN/fD8e4FRi2R3QekYvx
dWFKhzc+1rfhZ8wxTpSJCmXU1vVZ/pDR1mKvOJtXRrJ0KyjXKUidPY8oZqRt/glV
gesOAd6uIqkO9uzSnvYU4UnzE3x0c5yeo7gz5daszi2qWu23gUaHw+MneujOEaos
DqgSh2qEZvNE2Fn7UtvqjOP64Ipos9wQDRLBE9zr5lHMaEEM4/8f7IyodjiQ//2c
/3sbCBqiaTlhSvEEsMd2g6n24UuNhQtDsH+uVKCfyzjy7B6/bpoVAbb2Wpvygoe2
bz4q7lMyNIde51omThwOtTRH15FjnWKMaZCnmEY/jaNDAfIqP44b5S2Cwjp7QQ3Q
o/cdmykaCmTcxiQFFsLXt1BjIl0VxsiEM+CbSyVqndRevDBNx3dmjHzxbyNU+BwF
t8S6wQTlieLJSnQZB/hfbj89R8MrNksoI7XW0suSkBUFOwvxD6bR0yfjskiAhdsU
Jr57v5bl92vZ/dKDviDG7Kr1daOLuUYbN/QlbCmMTiG3I1EVPtJ/DuTTD9vWKYP/
MP2OnTivZKzrvFJpTKGd+NilAKTo5SDS8yYaAewgCaMkVinJQB+50v0P8rILOVIv
iQ6DTvyGddsgsAOR+h2ne/42YdSHSBGeY7+HSenbk1uOragCcahcUkwPv3Dlz9Bp
wip7k1VUv/GHNWiS1KlyuJqVzob2UnhL0nKCEUK/ZMpDyuBbkmNp/MqRbcLzZ4Py
f7ODFz13XV1UvClad9sNzMtDtWQZUIW9fDEuvq+k/Pz0nkEwo9WePXA7lG9rLKXQ
M7bDxr8xO+GWHFQpN4YE1Q77stY4i6HFvXDq6VROa3mBTU/PQSE3Vl6jdAJSWeAK
FQfTZDK1yHSrsT9xFPovOCuxFsPcpH6+dfpkW7AbdlcpM7J+ud3k2iEXt/jWSZZE
I2dCWChh0JbATdieLP331FM4NyQZlPkw7QOYKPZ2Ia7mbWy3SVQnVV6w+fYihJFW
7q/R42qDReYljCIz5XA7cP83GJghx/Fyvu1s0TOvjuI0M7idQXDTy32b1CXaLaey
cw/o4VEupfwL14B+RHZE4+x7QMKGHz3ST6hheNV9CPk6bF4hJhkTlzHHjRGwK0th
+dWz5nvym1qqObLtcss0YVZc5XjYjyFQamnwAdmkI+jgzQwMuneAnk2TJAWPiXUk
iV2UmmhGucPcPmw3jvbID1ktadaaHkZmNuX+vV2PJfGQ+YL8jwTH4CiUseAz9Jto
NVbszTAtejHbfJzfpjFZ7f3+kT8UUxtCdcvejFQEi9AXVIT3DKMYqcV7mrqYoxum
B7s8On8M6ENlGvSrP/PNgxI+4I108Od6MJzeXq2tT8dJ5DguZ2PYrAjhX8yilhU8
81QU5rCGysx1QDanYZqnoCSDFtm1ooQeY5ziLbLXE1QHx5cM0bOUWTZnzpaU9PVo
rxca7jnKWHtb6diqfgE3jD06lR2P1fyFmW8B2jl1BdWQieM5tG7SDDHfXGcJCX3E
uoI5VTvWhoP2BbXbFyYWkNpPf+Cx/BpeJJDvqGMGh8io7nN3JDr4t+p2DWAVYdgo
A5ng6BdUao1SATSURLMQ5T4oyJx8OCx4bojLdl7vn9vUciSO1A+3dA/esQhOoh3w
sHMTO+UYxxKjAjnY3NdFW09sx4zyiyY+DKD9aGbsKIP3yuY3s7e8V6mnUT0rJQch
Do5CZfOy9esKTFTBeYB+h8jAwuq84kR+VPL48Z7f6RDABGa50Xr75IfxR1jRNvy+
dEDqPm59RsTXIuMT5OsqBlIwSGqF4M0VptUNTinqGbAv0wM/+Sy3qpAZiIWHbS9H
GsafcSugVdzbxJlI36Qcrzb0CLJod1lMfQI/FPyzX+ajc75ZAdZNRXXvGv9jJSit
zDEv91PltDiRHkhaUZpVbiv/LBCaPAR2DL2RyxDqXVPJBDKM4leaCHgFgVHDQh7n
tieNa/L4QLUl7/eY+CUOnLid0jGzo3OhASa2MmRTlnHmw4tqKDsJz0bc3faKlU5S
hiig9oeXYWkcWzkucaMUYE49VwZHZOE9HUPc5BXsuCutVFp7mISneQIbiCgy86Sk
HNd8HyIhP3PX7xdZ9uEg7llZ+jDQ9tqUWq5iWJeEwTn+mnZKnbfXK2QL0vW/DYZ6
0Gx6KO3Q+D8frPxV79Ja3lUHidSWqaLohN4HgEmTx5emG91pfpUTHsdpKaranQ76
a+kGyLsOcQaYYKMH0EpPWzsYAcWMJ7HF86fTEw4X9fEH+KygFZXkhx5y59AFu6bP
vhmHniGVkPE9Yu4ZkjCmk2yB+rtSvqbynu6MRBTK17O9OZGNPpmV/6z72sdXYJSs
KdBAhuFHs3kx+Z1SNIy9jBIDQNNHBEiZWyr3pLA8ItzfepngWH7JRSPVAHs5TrEh
3+902Vv9nUpHAYf9zzT9Qcv0s4rlU4DY8XYPRIaET6+5wL4TPGl3/wLZY7TSP9uU
8vAcBdh+3DZZpSdmCzeRPPCKXFS/p6QXMGjKrcAbiBdQMO29V8QV+wmLVSLhWp1f
idkvkALw3j5t8KvgDqNmuKxA/zbf4zBZ2ER60KevYsvgmogesPLsWP4garSI4jBt
VNuHSyrUmjO6Niwaqy3eEQ00NN5nWfDTg2qOQ2YbF9TPuOUTH8KyVh7rGvQoAkr5
g3x3bAlP36j4cyszbKoKOOMnxroFiaqzmV2DvhQPT/0g6VQ95S7+xRKWEdAb4jBt
5j8cuvcUJhw0a+aTod56fwQ/j/tuf+gY+9dNZcDVzo8Jv6kdD1JhUMMdmIp9vp/j
SoqofNNcm+IaNgutLU2LaLRqbS62Dr728FYvCpPOHLABOOtnvncqtNdI/tNZNznn
KQgYXboBCcFmkOTgUMcC7Qv+wHW3mAycWdzQlKprpNPF+hRl2dSk4XdkEhDQShgh
14Vm4GLtHaevx5ui/f1dcoP8Gv+hP/8d3/ph4Dygvn+pbcNOIRUHH3QNLkkpVWr8
fCKq5s00qZzXkbqWaIUi9mrX2x5873HQ08ev6m4pxSq/Q2/DdnpCDnui60jRJOys
hQ4iQrJ7Apvjh2UaSyH5jnMKp7O96E3TrKTbA2wAI5QgJPHdXHALV3CncJAVH7mr
o3C0LL5VtyVkSqadaAYTXmlvCqE/CCaDv8bBmcnyEJLDNOUCcZHT7sClV+JFscUt
cErvyyXHWuMXtHN0xyjvhyKswYm2rTjyWnCnP9xVY9J7MA96OOu6YMx/AAit3AVi
CR83M8FBAFJf2cGd2gldje4HIu2oknKl+XcAwH0zjwK6y6RlvPPPcidZk7cIVUYv
0E+me/Hr9XhL7DZ69cb1kUFiC5yqa99R7zr+IJKtEgHx4jJxo2iikE5cHvTfUlQ4
pNMQGZamaoVX4mSUZbJsrHTfim2y3a3A3rOQaj7WGHaMh/D4V8asMoAOydMsHKln
7BtAVvXRuWbZ8Pkd+cZFEpsrnLqcZGFyVA8BGsyeB3oDmZBCZgbgM1x2HwTNZnGA
yS3en9K+oxx87F5SgmQP6oxayh+N4/Dhm83RNnxPBI+XAbllw9U/mALk1X3yYRvH
AIXTM9l0eRiQamaURWF3CnqVfzqmaqoPIemLDTl74InDTJQdazTgZfvsRuByTIvn
NZcrsur3+TKR2sSAfQd3FhbTgYwQv3gn5IHrUFVAzOydzS550E7jJMftrBa8bHzy
L/Ir7tK5RCZs4zOU+VctvjImTXqezzoupHJcnW3Y8iBWd2AN7VCItPZzeBwXcLYg
Rrg9nM2H8tzWdppW7aBei/+m3LlG0Ved3XeqqXjkrC2jTAMIPS8lbyp10p1/sPgM
sIrTUpEWX/xBGFd1XUGxO5clV3HUXEgsNGm7eJNVhLxvXsbw2Ur0bILX27rl/TUh
j/Pj0+IRPFhEEFOGpLdYayqbepfUBSBhAi2LcOBgWrDxm7tWPNnzJPADDkjqt5ii
C1L2Mz68Eqk5xqkle2VrSs/px3/49NrnzMX4waKAgCElqrhXCMSm1A796Q/q3ZMm
ANDXsCYyC5IHbAnZ0nZVkSiF7Ifp3psUaCAg1zrcde6hZHixCUr6NIa19+dPA1x6
nTY/YpRoBvsV44TD49YizfOLhJbdT5cFBaPcmX9JYkEeZOgmJOElunKFhwwBqsug
jDYwhelH7O2WPekCLHIxlG+uUmRkHbOjsaXIdUrHLeob593g2SDH7TEBLcH8nO/g
YPHaJwG70/yBoDc0qbEiOfCZvv8JOLFIExFsk84V4J18FcJKhjw6pi9qXr67wAjf
uF2i/mkV4VrsGFhxIe0cVYIgrOKoh0d2+js1Zm91WGkq8vUwtxyTmnAGBcHOZJUx
Qq5JKPyIyn2yHrLF/ro7yWP+9DaUYBaaRTNU/VoOeFubaCKjh+ghIrtVFxFbln+C
5H4yikoDHOtTsyKi95i77ZsRMsXWz3PJGzE4/E8czMhHaprOjVQhP3wZVnPxdknC
dx0Fif7Bnxul1sZvcptw/4LaNTkevDd/hhYhnGsTD0ytOQdT5VYMM5CW0OqHLjI/
v2oka2oJ/3qKvgvXHjCEDGF23m/w+r3xeMwteo99amEkxO0hgdZ14ycID1WtXwTz
FBLrdozsFMPID2m9z3/Cj8WBEt0N5+jg2gwga8ncz7dvxnPhPlnN67M0Zn1Z92E1
jwkWtV7kE+DKvQjs0Ojm9SZF8Etz+out1528BCA6KAgUCefbyge8iOskD6MmDmH0
tEDANr/6xIYdIlCam6LlJPNJYPjHyJVXl7oHJL8x3yf4nkD/v31A+hv/+ryfZmCv
ZJ4NfPju3A67UID0wtNlL7HSFH/KywFSX0mfwWjCwtSKNF356hRxAVrAzx5r2Olf
7KHZKdmTBdwCrtDbXm7d2nvUC0msHC90MK9RnHZ8aBfVtL4lUzZ3awZ92TUH3N3a
Wjg12Gr1tMxYwE9rG0gGAyBW8vxa9DUuTfqstmhMqFxcew2Izqm5ImeZQ7ivGXjw
rLTRjcS+ZmSFnYkwlo6TbxMGmy03JffMubEXilPdQofFuUHf+xnzTYiup5oMyyk6
tZ6ujNL/ePtiK7m9aAoyfLq9eTYTWCCq219My/R47rW97pSViN4yeAZdJOBreEeI
d6qUiWPpfBdq9ATbhU3YRZQXs4XQRc1aFZ0fiw668S5YXDFQHhu/2SE43KaWCdDc
/XNhF63+Cv8DL/sMnL3IWXRcdhG/9rxKv764Fx5SpPu+tKwEAY+9bNr2cTRY45xA
5Af5YaBDeoxbFai8hxZDp+YrD437KEcK5zlhLdUBwhge8aJroNBu7tGf2bFNPd6K
G7atVa6Y0buZbDO1b+0Iv55bn/NM49+QEDMJggHewatM/M7K+2jig7qjrNwFrdkh
N8TgOHp0o3Wu3cT6Xt2m5+fRfrPYEACfTK99VNLHR+Fa9V6ZkrOITTEyxQSJbCRc
OU56iahwoChQbzwNyJ03AK8pDoP8MxSH4g7ghbzUw69zdI7FB/Fwt+hYhdZGqMM6
hMWXD6ru+eDB88Obym075d/V7BHmqslg5PSINmyzlLmOM+lZ3nXULSw2DJ+Oadbx
POgvkWOizTFmVbnh2TOR57Skua2ld//4h1VV2ARh5DitvBlOGwjuJePtUI6Nd8Vu
3D6SjPeE/l8rSu2qJzwzliji+iURi1ok3zf0jUr4pOocRofLipFYfS8ldZcZgdIC
h/Kpz/Uh9zNZHlgitHbs/o7K4XxN65BapS49JcF9BkLmSOyglaJcU7SEkD8NsViB
Q17O3w3ScljkMIcTKu8D35UC7lc0rTWOm5fPcIXBo48yUQE14AMIj4KLKyvIjEM8
660rXX5nKSxBeBLdpCqAuy2kfzIdNJrexhSL3l8QXVoVHsRvnvznLKpphRrqLyet
s9C0b4MsnPc7JP+k5htb3wVvtjWUuLq4AJr+Ma/romGte9YcZ6yGQDKqtQfn7xYY
Gwhev5g/wymXc0leyIEl/AWWitcIydpl/gOiYY6tE4vRZU1WvunGGp9wNvi80/7q
IotRMagOImQIAkqAKzIicotXnjIpzDfdWYUoc4M8aADd+JGogNaW6x136VGtLuSl
Otg2KM2JklDrRQiop8s2rtLiWsrl8YB4eRuNrV4bGoRWHBCv95HlDzp/KZyjKdsR
eJBr46rgYQzMc4gQdm++d3EVp3QFtRbn6RLqKsb6TubSs1qXGDN8mHZ1o3VBc5P6
g5TCRBxhOS8sTCCgeD6ZR9kNS1JRibt1QsneY0RrKd88+5KKAdJhwmnOPOchMTyZ
ZPwkb5H0BeZpi1Se7DJSmRWdClEhsvAHI3btpXRtTF+iaYcM7vlucZqzJkG0UL3O
+M8F6fZrD4n6edtYkY5TQTCI0o1bgg+lA8s6VDEa/LLOjK6/mHvnlMKkJMW3Y7r3
iN9vHYLsUrUz5kUULSheO105jSmHe4Jgab0P2C/IqTxj6/eYKxcilb/hUT2/1KkW
FSPU8/+3V9qrtFX4Cfz4y4dTT5de6Rk5PBr3Gqu5aPSv6ByvTBcu2fkWgyPuTOFU
vr29LKTtF6DQ4NqQi1NQvyADgsXD7Ka3dMjQfCeX7bQSQ8LVs/eTu6cxBJPkU1Ej
lhouiz6IK44yCcq77Qe6iaTgKCbbPn+vlq9U/XAA2NSBPdVMK2qToosqq//GN8yJ
2LAfTSl5EpYvvXSkfMmpB5ap7Qp+4VDsPeVGFe5mxoDdF9VlXMLHbn14JXX3SfME
Zzhh/CBU6AJxmz18EXvjL1KCcmGqYcuhG0l34Wtjbih+RDyzhApnYy41RrIiUGkg
g1afajsbLZI/dloFquurft8lIpCGcmEbmKzdDZAeRgYLoMdwTe4hN888W6AzQH0Q
oD4n4x/4mUZqECTJTkRuIMIiN4O0jSwIZ4nrCMhOTpuFOuRuronXTYAnV+NIAAgH
NZxkToy0hVnENjyiS9XnXaRB7uGTHjMwC02bcC+j/u2fmxn88M5rYyN5JcV0zxvK
KEGK4lG0XBcpeUVPyp/NCBScqzT51HRbYcFZ/yTKcvr5820Lcll2yaxtlt2aQByM
iPkQ6oJqkZFh/cGeEHILnbfBn2LH787uSgoJ96A0yIQ2x7bcHkErkMya2GcUYwlK
nFujyTUr+p8T16N/nv0t0NEQedGQjcy68vdzorfxaQ31zufY17x4NZl0y4Fruvsh
u1Yemb7ZYAIeJPsu9vTwIDsTRkeFUSV11jeEZs3LEkFH6nB2fG9il2VGNLycdZ6g
j2ehEXnRHRbFwYrE+3EXVGbUy/jm/x8+ztkZN6X/D0LMc4fJmOpkZ9peUdVhPxhy
rWYVRxVzCNZBE5NRfiCx6xxG1CgJcftlRzFV83BZ2kmSNvUV6Wgd22SRiBo5ICSA
lDoVAUlp/iQKaf+SvO0GaFFpNYHPDLeZdzj/vsb+zMofBpb6lY+ECjAVOg1TYAiB
kBrBDf0iCoWvUvs0M0rDS4UgOwqikWJ05RelaSx7yyIapVZDA3/M5CakSEzLYrgU
lsPtWFoZTF8OzLl9THnd4hxYCrxxKyglijDttAqBOQmRrEQl53SbajlPN9MCXDlj
ufXhcEa6/S3tC4YfSfDfHncC5aXfe5EGTpGpTapc8YHNnb852rvI9CIZA5B3q0xa
PTxqqpDJTC4PfaY0UM/rSNpMB13tMlY3Lj/EwtPsVqttXfklvYstCt0N/2zpvoQU
QYP9E9ArUJLOv2svNO7cUMgKfQwuA5NRwbH7YFuv5vLA94mbIJkhTNRaXtJH5Eet
KKN94rNxBBimS7i7LpJYTW6657JiRNPowzayO/baOEtULLtZmMLdt+i/ec1+34FW
gqIjqVu7Duv662tsTUbLlHzl0AonOlOZQ3zHHnEC8LJaqGupE8mGnwNFHYsilPK1
p4XdzoUse/tDp/cCrmtpwEsHbkzT+fa0CVkVtS+u4EPWrLWhQ/o5B99jM8xnfZpa
BxcuShnXTore8H66EvhR/a+lXbxqRVvytmyucNrh5tS2j/CdRd8iPZVDhH+5BvRA
Tcsr0ET2k2yfZhOKdyiiwOHbTKgbGuOXGqRamTCaKVOEMc1iDhn9E6p3oS9vIQFF
P8GRaBwZCBZQpRomWY5g+XVaTna9PNr+SxupEoFgmnnLquANLjeoByMl/mvUVPu1
uFdDBPztZSa6J7o3L92vSrSK7yBpRDldvhg5uO0PiHZz2Yo6y/YOi3v5p1/zlrft
uwgI2qfkzSiVs+R3RXhp+mCDD7KqwPmLurco+s/Rf4TrrDkNX1wFgamvvDK686hX
J0mtZAmJH2LiNZY+2ACj7GiIDXblz08Y4LXxV9IejNduuUiH/pmtv9IP4er2QBXt
06775IrfIWvAjgv/C3IRiMMqiIvIHWUnyLHN1059vjWQmF+E+06T5M9sta6zztG+
Nl6uYPfT/2+EroGI8tfjO3IVVrZgfzTZXMFh916F7PtqmRDF/3H9CQ1VVSGxtCbY
fDx9WcMfdCCb0sKrNSDPA3ymhVL2oArsRXwkPxmpLAo2Ka5OpWSR9tzNhjuJQtH+
O0X4sGS3gG5ZCUcKAARFhtWExioueXgk/E45t3/E4KM9W81TxqGmCfgoTxJIHorn
voGwWfXWMQ0nf+NbBUkbqRyYMHbmNr3+Ay5qUENM/PK2/LSwdT6OgV+5vj0p82gh
jhwtD0p90BOJS+J1fblYAGF2lHPH1ijTX4KXM4a4ezRyJzoopRNAR5BgGV+8sOwc
+Yr8+qLWTZn3VhdYMhbFc5T57dEGfL9gP4i3gW9rery2RHFvUcm57sr3IoKEoVEe
RTl6tFCJ/l7Pu2N+DemZeRcjRne+YMwoanNaJNTAZmKTLxy5l+lfmkezsdR7qaPP
+hgw2tCIK9F+JZc4SQ/S6PTJVQ4pIH6/B83VYI6HSanGYn38u7hE9pemsh/iiLuO
/L8g2DviiqZn0w3p95fpLoUDozM4E4xN4EoE2Ijg584InNTVXIT+lwsJuaCRgy+v
Rw2z2k1SlZGEVSj20bTAWS+B5fYiaAB68UNdT2mrd2DH0NHUcF31R1Wte1eTsx0x
QxRW03zT2EfIEj5U5y0lwRfHp3dggP1bJIeKq7To0ZarkqW0AlzC9kHtuiDrJDTT
H+73BsHM8d1sCYSkVoaeD54lcuMxO8q9QSg18Q4h/A3h02EXAPTi+GX4pMhUiBRS
8iqg1ZiEx4xXZU3qM3QLf260kZ8CSSOAetBDq0Vb9AlUjQ4xJJIF81GfrhL63rRN
fcr1m+UUBjdUAU64gEY8IdY1pfUAJ++BUe5aig2ZICNxMOR9vqaP2/jp/8pDyZkV
4wzX2oXE6uCqAlFf9FXNJLCAKQfJaDN6Ye8wPh0UmUa8uaQc61s1WSw2PyKwpa+C
AOI1B0VQ9o0zyfAxJIshwiwNDfq2dMjsXGauqiHGMX37pW2m0KTcRvsyOjgeI8Ou
BZxGDyOLW50i1SPRN8rtYK5kBgEM/qrNR0kxO0HAlACOSnxUlsWnUwdX+GeTWowR
+Z3L3c25XCI+z9aXm98tGhzYBTpG840Q6Y6H7C/fWFI/5PtX9P7NRL4GVIFXjuqM
0ktnywTJpGM0U+EtDHcEVOo3XTJI1LUwl4BZ3SgqfS/6qUlFYI7QeZjdb5xeVIbs
eluNf4X7XdILIgmFTVDSBZXQhNHDVFnoHkO9GiPy5XMibwXft9nr9/4NxNniTiPW
GQUKLTlw6xdGAWZBVxIzt0kpMQ1/QjI7aNxuQ7JYlEvuNAhMsJ1IOhs2wHiY1Dwd
8NRGCyvezpDC8CtxsXGg+ePrLR+vYqsuNGAdhFLv01XBOLj94d349RFBOfelPm95
Xl5oXLIJeDRB7j6x5YOf4HepGSaEJmR93Z10oSb4HsVYmLRQDiiDlBU6Vo6c2rQ0
Ks4q5liTKWyJOTHObo1Fcn1ogTd4vQedcREAG/8rENQhN0lQsO6qVi2TbKS9ZJ9P
oHu7x/aCMNShVK7eMsVL3udXuq5WKXAbvKwpoBnZrlkaOVCFWFIsKVbOqhRnmVqK
h+LkJX9ecoUhoXUzKT4JFBx2b/4ScFN7QvBMGJV8nPeY2aoUCVKLuM2PyUXe6WR4
ZcYiDxvtuPhhUEPLnrkLRChY3nWCZZhf0pTGG6l55bhY4sOymKIX2Poul+vrNYYe
LFrI6m7D2L0Up3owlWDUpT/WID7RlAHabRUuAry2w7kMjdotMoEhFhH9vFPuDVLB
cjB7O1YHUi6jwRw/EXUWvJqJrTgWiZnWrQVlVEZZcFkPk4k+YouL3p6Rjrx9aybZ
5c8/IcGmeXQbd0sxCWXHKg+tNmwHWb8P2YG8HLb7LQYDE+wUtZS5enegmi/I7t6G
es9Wwc/BEqRrwXbulZt3A0uNrLDElTO5fCXjycGbecttGOzk/F5nzdn/h3KbGALg
0cs6j5y/zWPdBqf0+jXXPWlhpAAYLH5/eQTUT7ip6UIwrom2mdnwVDK1hgKPOcVr
HnG99nNtl7qVcG4lqKRmb2dpypeXCVrFkkxq7klgcwSMTbqDJoYv1sWv9fOVsz0H
X3E+fOWNeQM8TIKKphnAy17pXBelgUzAj5YbqO3yHO3P+7fdsqjN2qzzOS4baPty
w+BNtST1xo3WE0o1UiU7lv8S2nD4JfBIlAFBEFqdSk0xHWY25REYIqteIlJ6/Ckm
STxq9HBIh0PH1voMSSKjLu2FaQXTve6eKhmraGwX6n9WJDknJdcKhNqLntJ/1Nhh
KXldzul563O06IoKFVZ/huTBq/OZNnoDQ7Ppwb6EVz5l1fSUdn9PIh0af6PW/BHz
gBSPoA6bcMdaHCM73pORxNkmg+zgW3t5tKfl3BTC7jfWv903tCw1Z5tOmVQBhH+e
0yuynoP9YuVP2WZiFm0aAJMCQVQMLCG9Nnj94W2mn3/S/3vWaYWOqJ6RRnzHsmGi
fyShQVJcqP9ljDRONWjQc2nmCT6OoD3B4kPga08fDD/+wEg3ZcUiantCnyh1iDXF
4E0eYcc3QvmYgMlQVly8bM0DTqPxvuNHfu24QhHn1pI79veilcu6NfSZlLRHM6Ed
YmLu9Xmkj0dQK4XbwEyAEEmvNbEoFQUXGGsXRL01jDl1YYksWUIvMPeeCs1kbMB4
km50cQzPNTZIeM6WBSpTapVtQCqX3kFcTaL25AGqiDERQYFAHkR1ZZPQ8ZAqaEu1
3eZPGBIoCXnIEo57qIws/N7G7c12uLFEJJzKdJlIYH4b7qhgH6aNp2FJu5ZxVZcg
pZparS9yqkuv3t3gb7dGuQLGATWzXAT4yahGJQmWdGMGdAar2e+I3MzSqGtgRAqr
EtLWq5w+MHKShLw1SkYyOVbozMz++5Gow8uj0hL6x8rRkKDv6UQCMieUElJ+vhqI
GziVdMt+sSIlaq2Y9tBdQ7kuJKOfEVOxcE7aYxPWUxOTqsI6Bfsfmmeyc4RiDVhm
M5DwKucmMIqzQJQCrlM/DBc0ahGl/56Q/zvjcY/ykpt5dLK1824dG7A5WQYvXU6Q
UfXl063qm8orBMC5LZiZwLCR56QAbLhiJLBrNkTgQcyfZECAqNGoQWabG3dJFr8a
Ao/Jrni05bEpoduvrl09OYlucjEHRz6FmSWAyPGJGG/2EsZBRp1UD/fVCyub/d8z
uFGY0HML/ShhJi0VrcvSYDGeDX3uiT6geLoLBrE88yhUuNfXPQzLa280M5TGneng
HmmBiqsczHspsMM3uitwFRjnQmTmGfeFKG9/9zWo98V8uk+qQLpvCdaIKD6cp59K
BVkdSV6UxeldULy5eskal8XFULkdztobO8w1d/65wmfWVKKnfsb5fD8vZmAESyPp
YLrf7r3LSO6Bbq9b99q6nQX63SpUdcd7JiojovO/cleNHAv/fOPK1LEHx+9jawuX
24zBx8JhuGlwlaba2FPXOBnL5staSxL1RuIJEvU/WiGNQvKaokZrEw5d5Aj9pBUQ
hcKubywGDvWgDeNiZAzafXxXRL/hXBFBwOI4a27LrNFGwid3x1JgqTQuwdviEUj5
RzIQAQ0vsXYcW/nG90FUIgCqYXedvgLvieGGM/k3lacbYG4zHr6UHyrxsCLkJR5V
zuAGkbZfDqWIBjjQfoIWSg+LPH3oFl9zblWuvMb7oCD9D5Yk3Lu1/219E/BabrD/
IEO6RH+SsPy8xyZmP5AktQf8wZC1WK2awnvx5uuKi+STWjdfE71yzBTQR8eDHo4q
mq7Iqp/b8s+aR5Yz/kzx2q2b72CH2yorLRbefOFG49UAtjrnBxwLmNVBo2KFd9RY
PD917HEujUujYQK7ZHTvQJspWSxyrnDvAax5UjngCw4NgV/XOghT+CUwO2XFJ4uy
6eOs/ToDjQyif4AfUMOiNEoooKZdDt2bwWKJ22Z8UP/YVV9UoNOH3UbidoVAQvcL
/GFkhI/8hdhrF9+HUZVE+XNYAUQBqLbZt1cu/iit99y3LKx1/1KxAk9v4J/Y78VY
4FdTL3cLiHot2K1gBMQHlbPNOTzPcg2loFX3bC2J4GsqICYWFBoRZxgDv1+bbIec
KMw/r8w84gqNdPqBWRoZkKkvRC7Kp2SB9yw4TiqJZ+XeCBhZd2oZWbi1EDcJ7Bdd
T/A1BDgHakVMnsL1did7ltkkgqkTRS6192gw2qbkdbgPZjOM4C8o8JWtbsNVAkXN
ui5RasR+Ij6M7WEvNQA97wiMozTIsUXfbnYnE7h1ANIr7eqxIX9OtR7bcTixyJw9
hrqghvX3xdmvNIeZSwc0AzHcQLHJwL23HfAQJ7IVlulYWuwT3ixrN5RRxOVBAlV/
0e9xYLb7hzKbOqxvVIACmHXk90KghiDXaPKejp6deN1nIKVmeQEWwHyNlyPUF6GX
5s2duW2OCezQ1Q0TriWIoPkxMx7XiZB1qmOS10Mx0ErD8L5i+x6jhjl8mVMrb5zO
qBUoWvG4KNzwQrrusn1jBFukNYOA+rTmIAPxVZb/UUU76JY700QFxAhYwUz4zgXS
DTlYR4duXezMIcHwlUcXatHHooheae+ViHpFOaYxjRF88c/IofOP5/1H5ig2LVHs
hMSmac6NDLg56WpgEpeb2weP+gtPtoT22c/kfmndxQgN4YVqFGh65FlR+RgQPiMo
2YSgkg1AH+ZoIjdcInVH2bPxl07GZL0EnsiW0jADlLpv8LizGBUL0wyw39Cmq/TX
QUyMlf7/En5/rNZZZyhYb07DrER3Mu55fMgLvg2zjdX2Oa578VolRnuwS+a0VgiS
N4YTTkfGC/FEf+f0oDLtY3aRcVio83Ihekyo+SFHsnu3jMGD1KkYExs7pvdnDFte
KYNKloXruddlw88vpTpuXlFdmqG7kVCO3hE5jC0LMlk2Hi3eCTLemfFRxb/ab1jB
lhvzeqK3M79GI8aaic5/Nng3LvoEqufmeVcKrbP+NKvgfc1XhArVnoKmEvN9NdmK
4mo6tq0T+wvMQuEMtOuFqme+ZeLwXxhTNG5CEVbPT6kAywhszQqoeBToj86AJ7Ks
x9fai7a15K56zJkcGo7R6RVGZ4QDf+JdZZ9XkjY1lRhNWLBqYcrBI3i2jbBwetFq
DQ0KwQk9yThlvLLTX03oLF/gTRahyEJGjmg5P62bfLrxQQkbQuprlS1LQiB6ijHV
WTuRgMC/Ss1pD/TavUHWnAWimoAZl+Yf+G5qYnZVXlrQnFuXH0ZrtTNFrfRrKLWr
qUFf9P18HY/n+wb7J0z3li3vuafsL/i4p1Sap3FcUV7+Oh1Y6/aQB16l+N/F4Tpa
CyDlfy7g5ZPNTZqIY07wRkc4IJDm4dQVNNQeZO2tGAx/OJQ1sEU+QU+cNUdXSCLC
VauIze+A3kNIKVXbnV4R2jwRs5mU/P5x8SHz5/zaAEBTzkiEpD8QZ1OXMlr0uxJb
AlbsdLYf1uxwRbdJVX4GWwioyy+ba5+7pY/Yx4KREuRNKLkw0UKF52E8moanTBId
4TGJ87oaaKfxPjKnGniVJ6kOVYnV71yJdUUCCU40X8XmtV+g818ds9c1trAKSXTd
a53u4GwVPdlIYHFi8u6Tg+B7/9sTJBCawOL0TFsOAG5UjKqDxhWdX++P1f5h/6M0
iYkMen1wobMWdyTu+F+YxMqKpJSieWOp5zUYgKqbVJ1VZPteAK72v2D1eDWFRVk0
P4D64qjkiYC5GzmmdeJT/KZY4ozLprX4QkYCF+k5ObKvpvYe8OT/3fHgVoww0kKd
jgWwIS2oecZ/0SDHy79GhVmf8fpIJt3bVSWZ/lPThmIdzMwujXJnbjXibD3wLrHw
gi0DBWy+7QH7WQX0BY9+TKlI8HwLEi1wkj6Cg7dkv9stHzN9RrAg0y3XIv1jN9Py
6s96q81r6PJS17tgyuO3KkLlVa3wXeTz5fgfegqxd1knmZD/Ml/PBwtFeVCg9KxE
3PO2aKt4whoMVhqvocYIbf2Kh1WBCTBRdH/hOD1B1DWM3bJ40T7pS6IoIAzuw5Zg
kQiVCuu+VeTnHRwtNe+QpkX5mx3kikRMX9cUI6TR0dk35CPg0zT6aB9ipE91qfnx
SRyuyTf2oDybxaq4L6AR7FrPAn9aL8vVj+iI9oqt49OfFE6GxwcCtoqfQc9mmYIl
R6HOFaNIJHh7VrKQ+Z1LUjZatk17Dr5SJq5Fz3L9q6+bO4/+IAbUCkZ/i7wVVexn
FmNibGvWTvc3MUZIllUvxYK7J/z3vHppbwkBQw1FzijcbQp+xOAtHqEOO8rnjneY
ectyWiwuQXlB9G+7UnXj2AdKj4HrlvQcFXn0pso/kSwN/VJulRorQst1a6sqTY/C
j4jW2Hzt+9IjYK5kQxsZ2iLI/IeBuqEWy6e38nZVLu+nzp61S1AB+HyIpQ/KapmH
84/+lzsusUG/fbD/zZnG/gWBLlwYk3yA032XPukpeaINOan6GZSVCjQAYzDSa6bX
BqsNmPzqjjXfMSVEAmT+V4zSboAgjq7UqUNI70lw6Qs6Bu82IsIpI5ATVdP6brY5
d8xGARrgJO4s3sieJN03jZIWSs07S8oPgUo1cgTBHQV9x5bH52WHY4bC8oamdlc3
Sb1zJ/um/CV8w2BW2+K/wCznV9coOYTBHltyz82MNhOuTMRI4LhBMMpNQRV6oFmA
h8rOQwKL4KB4+LonYCrnm6X0R2sX/uosk3bYFyghd2vjLQ1hgf3yR541h3pmBSVE
EP7KVZVgw6J+ypT9x4oxga2X83YxJVJwv8XJlvrwSJB8afwVy84oao7pb7WlpKPw
hPePPvW3D/aT+KAXxjVOctqjsSiY/gU7XZg8jXGKw01IVIHNuwFYQzVTTJdcOGRl
l3lYSGO68FBhemzUy/rPvsmOXVEAdeS512t+9GM/luaT7ZzKK4jnPYcQZwSphd7C
+UbiJZ89OD0EBUxlOEtwWwzNM/CoMSwTLNIwC9ftN/EYCSgw8JyUa/4DM64fCvnK
KM5S4HdPSPLThHY98AvdCf1HmkoOcNdpomlBMRaf0VP0STIV5UYbY+PGf2Z55H8E
+en3xflSJmt19GIYWGykUtgIvFWRo1ifxyaGfz2v6OZ+oL9Vt9ntogUo15PHiZuL
LVbCZ+BiUNTmKN73qZSTsw1iJtdiPA3eWbfiXix+RQBdswcVM8l+hyFG+w+lv8R4
yK5JNABrdwmxv1oRPYZjKg2G6JveIk1cZVttm59/KOvksTRiHqc+tv2kOE+P9NAG
/fNwFfQqpGP0o9SRaumlKqu6ToS2wNdjMXMk86OibBQ7TfNbTY2kEindv9hMpDil
X9r0a4Bkr7yN3nrTiICIa/yd1DCGXkG4/8aCcXcmjylaidwORwsm65dPuLP6bMvE
WnpI2E19Ri0scIKbARnBxYJ34g9VB0jzRkpxh12lHGQobACNYjoFAve+1svSs6wz
jc7NOY2yrtAowRxruPv0ZIX+cyoQEcDSZM9GgAIV225KLiFJMPUVGfn1hdPxX5+l
5OUdJkAeR8Fqon7nYis2mIepiAMAfrQFQbxSGAnQkevnZHxeRDE0zBzXAo/EAiIp
CvcLPbIxofWbYzONKCAM0U3C04YOfCQcI7rkbKc4qb6A/CViDlvvOCyLfligKroj
aK+4ucKSZuwtfNdNiZ2eYKWtMDMkUpjBuUM+n4UHKn9DZPQ+g7DQRvH9uuFVeOhy
aCc2Fhs0HbL52UIFMUTQuxomfZ3CwUMkBwjbvaVaYa0HyBhIPNS9Iv6gsvvzUIXQ
E6oIq+3SGIbUuf10kiq8/+dF+EV7JSHv23dXtsM8hLvLEmGgs9U+qlDnnL73M0OG
dZS+MF9SlvXwKoe8ssd43ztKNvMuGCklkZLnDNSX6CXheeSPRM9/J8FXFfzraAL2
NrcIbEK99mL72qB2AUpPRQaFcPyAWwEyfU+ekBFs9zTtXP1JSInScXrdnExrmFDZ
rw548gJFJRdhaN/6FzRIUFWtv/xryrIiSKQP+Bw1hYpISzgwZ5H57d/T4f6Rdwsr
qZdr9klR9uCF7j2b8et+36RQNSG8iH7s/VE0hTgr7iKsPeE9k07RGj1cyBwWla5U
FxLpL+SLuAaGC5uDkc560jGYE9dYKOF/xqtd5AarUte0j+2KfpLYvCaVTqgDAbUZ
VflweHCm6hKg1dACwp205rm6ObUuu/eqBuxyoy2VwpSv3eS5cmkousdzk1/r0BEl
RdP68LRhb2kwOcjm1M5Qa7OVwHv+2s1I9LnhaORO21B1TrYD2zt1yU+0/JUrXLZC
XnADwBx2iu1E1+kEpIr91SOJSyxh2HynpsYqYKSNWiaP8AqgiSngzVBm8txC7yUO
A78+zr66UCsoFwKv9CNRa00VtFWbvVyHQ2ew4HqhiR6/jrAc70HtieJZ0giSvfQ1
WrCZ2BiUi42O3MdMdb0zoH50B1J/XrksW4smhn6JedYQkBe9mTYuSmNHi+kItJp4
/jqStkVvtpMSnSlPGr/P+qOL6j0Ea+X/Urv2JZSGfbWYc37P8SDJuE9mfkcH1tY8
fYEip43/Tk/am0v1am8G0gg0WbysTHSIbZdS7Ii9Fy+tpUtfKifTLXy6Gc7BA2Rk
7VDXjCKQhfn4/2rTCemtjUDxY9HCYRyQz6w78aIYbIwmICwLeVz+ZvUsrAbmUsyF
8lPfFNp/eCIANQdfS81K2q+KutyGwiCVmpfiglJDl3ThTS9JegDNVELJA9Hi49Cg
m13whUK3DzLuxNRPmyK1ysBlmnmF3sdLp6OnZAcY04YrvoACvuXoGjJEjZb9pc3i
o0DbsHA9pu099D5aaurHXr9t5kNZSFwApuCLHc6zujoExSgxJAb82BdnZpH4tqy3
Nwy0TcwW5TzNQ6APvUGdxcsJc+txFVp4xI3nAAVFz4MOGSmxHELV3clpWjS9EuoC
snCCSVLPyicuZ4rKM0+osSRGMByFTMuKlEca9oQgX7ZZG2Pzv/Q/pFMa3B4P0/aJ
FoTSmKPgjhdgctyMImAsY9xZ75v7I+b+Pb2lHCBGcOExI5f6FqttrOrnr6JITrrF
4istQggg2Qlu4d9LOJWxk6thGzgD13Is9VIaYQbP9l0eVsf5OrUDioWvTYF0S3QM
Js0HuIt2NPrsqf8GKHk4VEe9DFOYxvO48ydaJv5jflDotKqbYPkyBzzj/VromEdB
2bfIfjZ/ZOhWJs3MewVCNz7e4ir4198VZyuheM3NEUZNxTz0MSwdinPQ56A4OFBz
VOX0bNFTO/4YYloH+36c28k5lqtf7Ev8NghUZ58qCJaDtWvQcYQlFSR3YcdHTDFM
9ZUPHGN8+yy8SRHhZKe6fU0fc5U2bY/OmkVxkYWDAfT91etbkIS9tMdId+R6+0jo
B6Mn0tm98HSR9gbU4xwZNs/esdI6VkQ/rZ2zDujHJFTUAFwPqtM/r6vcTamGM21e
VXLnIXLYwnBWfzpmH6z31Ksqkf+k53JUEn8vMbTAzGifoUozlc1M6kODjTQZWuU5
nf9fwO+7npJbiHMAxKZtHDOlLL8sWH2OojANusAH5X390L+9idTm7UGmBygqMtdj
rQ9cFqOLxFS5Qujc5P3AzULOLweBYVRBcykY5gvl9cW4ppfOwBbDxyCYPlxeNw9B
woz210Lgt05X/A8N+9GjjeFE7Y4am+SzRhFjFAm4KBC29DtbOwouXAHv6IUxT5jx
qaHQvbbBOsM17Gztyko6iUoVJTx7wYnlew0TYlNBKkQBLV+CPzLeJiJ2TQjGmeOl
cDyY/MjMH6m5y7Pvh1/JfncfQgjozxwmDr26nBiEtWkdIfQDqESSWVmKMlRa/5tw
ow4lBSGXbtIngsrTLI6FdIpUn0ZtWprDrin8YHmcWBPV40KMlsN4XTUeVmtShFl0
Y2r9O5VW0pHL6g/GWxSwOp9qG9yWd6V8iY0er+NY8MTE8KSWYlxwIHjlcMvaflwf
rHvn+yXmHAgWpBppjEAKO/eRk67+H0y1v9yy2fEqRNcHXxGkr4C8bR8RiFNo7HZ4
fj62gqcMpBa5iU4RzTnAydwJmHAEBHKhdHemBF33NP/cFXccXr5xJfJxrirK5OV+
5/H3f9erL7RRvDn7rGtQk5iZBJQGIIYCyUv5ZhxcqhfsofE7GsQExA+O7ft23w95
WAF+TH7G5cRWIYn6HsvnkZ6rjlJtCjH79Nl5gFm+AguTM0+b6w9+vpVuwJKgINh9
0TqCu2xMAtzi8RKcsQulrWlY5FFLeGupYBGvJ+CSdzxNk6yam+2cLhSOJ42nj3zS
PxF3wV8bnqHRtcKqQiEdoSUYS0pGDAjNkSGf7tmuNnleOsBw1BeCnjtdisGwweGm
Xx62Ih852AOJiHukiPoYUaHZdnn6QPcmPNQDuzgQ1jIZTfdx9vDzy8yTajNEeI5C
Wq83QjQGcJcbazWPOLO0yUoXEISEqHso4TRnr/60rVV2lQ35FFn7fyriXhqapIUu
/R+TG7UEU8JUIsyYvNl40hITlUvJJ7SfRuUHJoLh7gob8FWoBeJ+cb+qJDu0KAoR
ZFtx1cvXOe7u2ffxFWucSxdId6W1NsjHWLPcbkqiRIjpcim1xNAmTq0mcDTpAnXj
wwE7dzrj8IZ7dcQA14us0E6JiiHl1AQATNRplmaaHmmSBciz2Zudc72LC8AKQsno
1fOnBw8+hstcoP0mvZR95Ht/freizF4n4BR/kL22/UCJOlItv4xG9swFk4hGtWxn
qM8+RS7MOT00M6umXPuU+ugJzPgYiKo2IdQ1gy5hVngi5n3IJ9YwwpoIng5bDfLn
yGCjZ2AoM7p3mT7I9F1UEDbrshNYIinZKbOelOShD73TryV06g7qWdxdeBfdauFt
hyW5emC7dfZekD8Ic3JGys459ryRyYTGvvIu8o3XVx1JyrfPoMU5EO1S+ZK1LoJr
KCD1P64S0z0VrgvDXYhwbiSDBtm8EsXV5Hn+GTUcGc7/F9DFF4WcZz0FRN9k61FN
5RmdDllXeSB4HRt5BQ3NxwuH8LESk7zR0psAH18nDQfU9xYFVlaJ6Gp6evdH0yM3
grpr3pkhIprvMclYeICcCHTznhpeBU6XdxgdJrqXqFgw3eGZ9TFmvu6XDp1+HrHE
nMNKwj115o/YTT0Keo2bBWKzkxszRKFPOAY6+b6l57d9R0cqd4pUwPexJwDSYHIn
b25YHupHNYf6qQDBZCz3lD9/p3VqJbdWiCSju0wGL9bL/HBvZHlxGrkKDnmbXKGF
HKKw8GIpd8GniNfvXVOtOKwsCRC3McfZ3fsfMcdgS6cVbeFUgsB2x7pp2hyzt8fq
+BiSsEKOBmZgS6tu0XftcGy3sKyVs4Lj82oGfwfvfZUCjTAauUtXT06jGGYH0Mtu
Fp+jV2HsV+krDXBBLB13g8K6q+RX+7mzjRFLQ0Q6FMT23/6zIqeoIaNU4+OO2h6b
nrX+xsthVcQ2gDgCsVPXUh6iFwcjq4QSSOHa8YpEDKRfUPqQagUWlfvyz7ZppHeq
w2i51x7s8aSAeTpIpRkrlDV/vL65ekiBa0906HI6UQn5epP1RaqTpccfFpo1DNXV
3d0MvdlIUMKZAXfYFWt8YNeSF5lWcK2kyFylIMDnQ/B8bo4DbvPVMRtMM1BF7kD4
6RHv6V9wzSawfelVhgUhRjT1pBSMW0DYIv2KcE8JUiPQdl3572AJD7nsNWeLeSeR
2U7tGkLfZI+hQijJJXp5zKVoNz5Lq9BUdXS9AZj+tz3RFA7sQ6uc9YV5gRXQdQXM
z0KpWoZrjn1DBNZUI1rr6xABtmLcTS0xlyBmdoI56TD9nRBnm8p3nQXRkl0KJEBe
sMutodRVh+2XhiGdFdhD8mFcMo87G3Fx9BWuPLiZzmCzl4XItV9YFVqh1vlf5vic
S5pDqFdSGonVfMENwLDq4iZX4JH39Xr+6fVodwtz2ztuIfibPuDTsVuHwNwfEtG/
e/QYaCnPQGkYShUelFoaQPjj08Z/E6DHZZyR/Nkzxy0adqlNi8MfdaMmQ12F0W7+
eZDv3v/Y5asbRuEZb6nmtnvk4eREe1WxjIIRr5+BsrALX/wGSAW2l+VIjqzCkP0D
s4TWjGhym++nMT0gmgnzkDZTjkv+2JTTWJxXlnfcoVwM6hUNpFauDvIG6TQSxwSd
DV08YNlzAWf3gxcxIbLLI1eQbmHyTLAIz1cGXVHMZdHd3GGBk6iXRpT1UQw2Mtfl
7Q3A6+gd6MmpQ6lARwy9lYnaGMAjldPJHrBSU9oOgISqGBzDZuUbsZmtg1gpDKEt
cT27DEJLdt/+RKhjjDkEIt0ZAb4AyFnUG6B1d2oYC0L7UWnsH7Ka8FJQa4tneMCe
BiIUhL3T8gwA0E3NBNwK9Ri8SQMra+OIiIgx2i66PkDrl6nNeYug9yKThuyJjIIB
4wcqEiR77b59L6oR3c20dSuJsixlYTalhYMz0mZyyOdc6E2+Sx3DJblzuR5sghXO
UaSBaflQviTYYVSZDeS3LrUexeu5fPaKwIL5Wjeu50vKH/vVainbdlYJcvyhV6Co
Oz7gW2qRCb5ZIckoTv91BEFFPtV/IRrHFJQKysxRfS7P3vfiBTljSB2hmeMyHcc0
ACK51c2thW4Q4M3ZD4CJOI3NL8slnGTHKAPhR5ELEFXc4+y2UW0Dmr5R9Zq+fW7Z
aXbqwk/cTzk9Lv3eLdOYuuZz+UyqNM8HOBXuXr+n1L1M7Y+BaI6EfcW2V4N2cgTU
F4/VUGT4up+0emPaBO3Bnod7pqpZeOHWTyO7JXcGzKtoPOR/WvUQpBxOdePlC8YI
PWSxW34alicfnJC4RvmxrYKuYz5pSOdn1N45R/S/4uBbuc1APM4J/V18wKLhlDZD
Jy92iJ+AtAoSJaPG5Ak+OuwRong4y/n1X3y/+yLMkrB5waj2wElXSm4LQ+Ada+9z
g1/nWY4IKYcNvFYF6elrMwiPHT811rCfeBVwA2lJDLHmtz8+SRWSUtTJgb4CNpsv
ZSpQB+IGUj0dwdsISvqOR8VwnDWYhBogHUIK6ZjuhoUurUWRY0Xvj1t+FzLOIzoa
tdFr+qrGk388bsBPxAgZ2hDxWHbzABHm5kSITKL9t3o/W/fMHJlE2OMSUMekUiAY
rQJYCeJYMxljkX6YiJar11qrNsE1TCcs+OGeD1ov2MHrywsrKhbO+uUvY45kZ+Zv
+aD54xNIz1h6aqyGnleQkSomdyf1cd6xlbSwrXe3ciR1ROMk/Ft/WlopXEZCROtb
T26E7IeK6XFXv6NdKzlq3MPK4LzEAEEME+N5+ySOqikFRCv58k88t2RhrY44E9Is
S2M0iH2vu7Yo+HS/Cz15Go2q9rLyd2dXKLWZ+51+eAsr/yRMrPjJXW8P1MQQZg1f
belZN8PCoTghpXMOLwwiODP1edAb8kHRGbSkn38QEtOjz3Ev5Ny/L4b/O6d1mGeP
CElPCWb7IVMZ6pLa1wKLyFCkVrZeptsMS2YVXdLlz4mPR1pvKdZfkKutC21gMZQN
IRH1ZJOkUp7N9pEzYZwFE+3SblBV8TQ47uwvDMcDxkBIi+nno/WE7iPdzafVEjOQ
gAI+gAa6jucV7f8VhZFF5NNpPl4HmNknD+xtvSA6Fd+ctIgPzmBkCskCbs5zgiyh
YCuUVfhBNye0B4Hpbyg7cqznhGG4dSl13xvsUkn4JRd9oSV+GfcgHV/d001vM7Fa
XfLgvHGBkZNfN+68QpqcmGQMjOke6FxGFYmFshlmpTgFKbK2t84c4RR81eYA/3M1
0Jd4H6zpnOX2cMZHBN4vBtXnoRkR7vSZPnQ0HZAb3zmymnv3apwntP018CI4A21u
Dmnr7r+hqg2wkrJR2KpJy9/xV5Thza675TBuuGubBEEbgb3VIXkNDEL9Bvtp9v3Q
YvDNKRLJI4X8YacwqDT8r4052NdItLaPaFoydnzDeMNzNOFDq37x+j+PBkR9dqjw
daVEf9XVr2j2a9txWuqv0TXmmPTEVlzSMoJe3TFAosqdPw4RVu30J10jcJFHqHK6
SO6+bON9fmIZxMG8wwYfHcUre4wwt+6e2Abw0PFKX2C+Me1beWnJMtY7+04KIU2A
pU9FChv1gRZ2PamSs6tY4qzHBCB46BfQQeKF8sc17WSQkpNDI8SFBLAKRNAq1++n
z/dOhLzF73Irb5gsQYK60ps/3rvl8CPvGESWLRiiRqq/MUmpL9rD/UtD+mQT9sPm
+xZpYWN3UqAxODsTiDUMP49SuRFGTbBSuvjZKAE0v0ehonv0DTE8jU69J8t0mYsH
2KoyOU2A21tGXqn9USlpzdYpdDKeUSOpgZfhPnprix18cZTqBQo9uxKPzBXANlb5
zspZ6e76t9oerH2/rjvGRgHFNn/w6QviCVLZT8op2XagG8nkXf+TrXiJDoi5oiCy
TgR21aWrfUEYdWJVqaPPYTe1D5Htt3xidcMjT09xL+XvZ0k2z4q9XEl3TJF4KoFr
2/QJjMQyZsWbIJR74YGqNMak2hfRafqSBnL3KLxdnI5a/CHcpGiXVXLYgrCyjjpu
aAbS5b7hT6ucsrNHHKRuCpVP+bpzj+W6D3fIkSa4Gg91vUJNiQxUxPVVtb5dB/73
QGkzy/Ncz7pI0IAYeW1SvBFtm8Db0rwxqyjP2zo1FKrFsDU1lOmbUMRidc4WAjoU
GHWN7qsNzmF6SBD3AVLDy8Phr9EkFRJE87JiKJJYFZpwf/1qTJ2UsOqikbKDAVmb
TJH1ya30j2eVLQDHeU/JSqnkige/p+ycuUGkqEtP6RfcC+ZK+69vSrKVh3tiq65i
bPNQPb0UgrEtVfOhnDS84pC1fsPjT/cOedzYOeYVcasp6wqcd8UZugFWswoH7i0Y
8bt++2rAQhaAswz9STe5VQTTfcQevRvNu9Tleou+ltNgXbZIUJVUkXAYTDmicClD
WTPsbVaSJHC9c1gWMynP2XAGtvSi+COOdc3c+QhSG/OfbWStyvybsCFNbVTjMynp
hptU1oq/TJnluzfUPyQ+p7Jo3fcPPSSa/IU82HvjV6Cd1sIBWLfx/AcqCuslQgHF
g958t9l6BkiCHOmmcuGjlBiSYZZ5CKJmP5LH/gQSPt63YxC2RxaayPSqMajCN5NA
kcYCjfV9ncrOjmg2UB6MrmxNUcIt0Ih9bepbTG4xYQyd2OY+Mmf1HqQXq/8qKkMN
pX/jkmjimKFFINXsB7/FUTP7rpjIhwoilageP3o5YHmhRLLyZ0L3/omStrxtaoAw
pShppMnIvKYAvDHZIh0fc4UT1uwtlUYuWvoXhCuSf+pJn09QF+eGXfX1Y3f/ca3N
0LtEsPcGsO/vAaVQdzIGj3eqgd+AiVEBfNvbJj7K7RfLJSoEgvPPeGhAk6UOf3ug
AVtfeCPPcS10NAMr8AqW3Imit/VCbG9SB4hvvkivOrDhOs+uhVkdG45kvJw1P5+V
nqP6vDOdyhPMmFl1Dsywiq8jgbrDOfXdsdpyc9nNtGqUuttCWQhVbt5/2x9XUv8s
CH6D9rq29cdz89MBdHMUWGMMxrrXh1DoylmwUSK49GLVUadS39bQMDc/kH3TD7Vv
3FxkRvAWcDfSxy8fqDGi6cp7BfNiZz1HyzfEyhDg8+JGt3VjdqqsuKC+Olua512k
ealJYypWyMjT5RxvaSVCKT12kf7DGgfdWznunyWBpbWSo0s/gBPCjTb4YA3Eq1BF
V5rTC5RDa35nVVZEF1qgNynd3t3L8U9fX26OBnk4/uk/oct78keXo7UUw8136jZq
M673u3DOOxJb82cIMx4hxz6PM+7EhuVVMwwThYFMeE7CKOrJCXAcicO25K+mVfbS
1cfnmvXgDPwQLD0FUHsd6i+KWtSkCPtKHP5Bmbq4V72o55aggNBoS89QEEAuQ8Nh
Yj+EtWsnlIvvf4L4oIuirZPNLS5AsyL9y7Aor/ULfPlvhp4Ri8rhQnK+uZQIXThp
eZb8SImWwZcUm5taAxzyP3SnBRPYk+UkFe2BYN9IpPZTE75m3mgxqwDuhjK/c0lo
Xs0BLhuqevNAcrrZdG+nk67s+yohTJ6mnPsezOOSQDcsVS7aq3a4CneeEqmtZz2Y
LExa842UxhqfZuUyyLmuluYMH5C6MgXs14Zfe5nyra1uoQZMNHC6kB9XGNLHkhA6
0Sq8oXFu7ctrZj3s5MjYR3fOtirE6XSdb2dXd5pOpvq3Z9POwXax5GYNT8eFNfTV
iW7q6nk/3e4oGAafXQ7N52fvuv96AV+vK5M9jnDqBLY9VuXHsREMDzOvwOBsbxyI
WepZUUV7+Ro2e3i5C3GBvLKLBcOvEtEQj7EL3Wy9gYdeJhWPC1cB8aCfaDVjH2in
R1XqW86nM+nw0NhkQShfUxXMEK+oawnnrawN3/9fOqn0a6qoXaWhFDpZFGtL1Klv
lmzl030bcfN9g/n7akigaE50MSFB2xk4UUOZhRt+ANVeqmumsBKTgyCGujL/bRQQ
+d2KPFQtUHyRVL7le9w4w3cZkIx7FAI1w1DGraBAOyWYbrQim9D1MbZ/NHJa47l2
YglfPuFbqoWty+CRDce/j14A6qHuanXc+bSwZcm2R2uOeEqfRHtegurzWKZIY0ZY
l9suWjWp/Mq7tT7b0rPYLh6WmSmoRzXARCmkSpzYpJOWvQ7zqUkmrmp2sFroedY2
AcCJSu9IL93Jv6KGUE7JKi+jMFH5FJKZGgDmZnMU5b0NZgXorZRFE/bNGqAyGwiz
sB1jvsG1Z+kLgH211iO00ikwUsnoFp3loMf1xQAywrNhszx2Ve9tol7CPzrU8x2r
J+hLklD2/uHyqYbRFN2Tgw5f97WE9+rGJfXB3ddToUhwTqWjcKpjkLX51TRP0eDV
YEClAKPZ/d+pI/q6fHT3YWsuU3HTnyKMRAI+YPk4zx1qFcYv+PxK/r89gl7KtdR8
+tcGeSa/EMguMVpR/0QTNymxTOgCUaWhPr5/Ot/stfj/MgYS3f/7SKHHSCJ94fq/
xGIoRmsaAgY/JKh1QrfKjhnwqRMFLXKRyQqFcNeLfgJv69V2K8972skNx7u+I9qS
G8ttl8UYtMtb/+FVb26MJ/FLMlO2d2G3z0m+WyVv0IVZrCKjd/LzHz4yzpLXl1H5
1cFsN7X2zBF2S72XLkLpNAMKb1jneLmiovHAFSr0572q/Srs1xg3HXaf7lk51I85
5XEz4/fDpu5fjVC+j10NyyQcvu+Trylv3s6BqNXenNgDacIpiu4Ccc9LOWF4Fvln
b3aLgdaO9IvJZ2Ay2TODtWVWe870nH/Mwle38sFM47k2eFoFJaPl9Egf1jSxzMNg
/n6asdsg8R6oLfEvttNnFhMLUYDmEIuHISnQ81gi1Yvu8E1KxwoxPfAsFnKg9Xv+
D12/E+tU5G6KNc+1wvotpw7KRPEzU8f5quvnKrFuUUVU/eD0M0lE6J1UA93RySqn
3m7yLAWfBaNoGbbPuF8tSpsiZFrqUEZT03Qc0ubkWsGgKAkkiB/JPMnf69rt4Xt4
QanJ3rol6hpeMhDCKL7Is40pk2HT9OKjBzYDYKF0EOXIp1vad6LULD8hiFsdpg12
JQZXsmf0hm8sJFhmcLPdXpqFMED/VC4BblI78sVY/0Fx8cC8ae+Uf3ZfQJUYE8GL
JIIzR7w9PVge0Jc2q7gvx2Ixh+U9zuHZuxyYbU4AdWzBIn41ebpDpIOeFveTYQ4y
seRB3b+mYAMry9ViH/UXTR/j2/eFraUSo8X1AQ4uaCqQlIkm0y+wrPJwcG3LE+Wh
yP/wpCTlNv7E/SME8u8E8M8Gu6HTSoK+aCWNXiSje7FKjgJffLCmngMzDMZjv7NZ
MEGhrempS63IZo9+u5I3wkDa4Qa4+gJLwNO4DbNhMos5GZHCU5SaSPH2S7PXFpEg
k2slJrD/M9LqeM//JksyN9E4pi3F0uRixSdsYEAc+apW7VgdafbOK/oNIboO1qoH
BPQo4etnhJRF4k2TI9yiywbplO8O5beHZHZlbDKk9X1ASF2J5N6/ces7V5kzIZy9
/NDqZ3eV5BJ4DuFti5GAnEA5YC6WkOPvqxWjRu4MlPQyFFmrJ0i8DjF4KyK/2SzP
zPj8wycJNlR4ScrH00Ac35p0NVIFIYh5LwUbQm0qpGDizd5KmxdIlChd8rDRkowh
xg0E7mZscB5HnU4HMNBY/m/K8pclpHNrQnKwIBS/Fjz0GfJBS3DkabW9IW8xxQfJ
gJyVmA0db1qtFXrfkIzf14NhbKKbpyWp9jze8ly2fadPhKEKaNtocNf/wemJZGbE
/P4X4aflS8KpDgz74vTt3oZfw7oRR7JkcQSHNqosq/bBDFucxceMyw7LWZcFwj0j
rsLEaIwtDbgoTuK6fYPCz/lQ8QkMNwU+MEMqhi+5rcnXhk2wYwX3kxrHjtWFoIsA
BLATbKHIpAVm1ENXzdB8u/vScjM/OPjFc6OJSpnH6M7btYTEvz2GKX6z5VddxzeQ
CzDNeVWGTqGYrP+ho2IUobqMqr6AMlGAEqYgXsWDciB+7RnjnGIFzMQfhtLbYKi0
cdQIAbJha05bBd3f1tluThiPJxKLTE5f6V9KWLlIvqFcq6i6HH8Z8U+3YrtpDu2m
Sjcku+anCNB/FAQyApBamcuK6DMeaEwaeQLHRwD5QvVKwF1I3rWWJA+dlG0PECOG
w63G0ql4/yn8wmYMjC15XCOL7Q9qS/AOzjMzMPNTuIetuQdlu8tJtxao9r2Rxjq5
8cGagnpo8BH8rT0VIQNxVbI6t3t758b617rnizDgPO8S5vphCztpx2yFw4cw5D6P
cTigIsIURQPDkkWhAdKH3rlDvypft6VnGjn5aFywAN29d0uxAAStrWs1T41x2Z4U
7x4qVWUYTrb09tvvt8wtMyUlM7l6eAfkDu2Z5wUjKi4phMLp8elBwjSx+zknnujI
CKifTOzjz/q4+TxlslpmWciLVxSqsZ3wvdpWT1rcwzyc63B4KlBxnb4lYyfWPOa9
l/ZZ/W6EfW+YD8jrr52Q8T+y1y4IIy1PzCVRVTbl9a/WmBNnSoFDcWKhQLGatzQn
24ZAbZM152cabvg5qr3nt37zqgOIZgxrOCXjM842+bIeyYbh+sETCLIWJvLSbJlE
EF5c1tc7y9y84DCHx5oN3RE5i5ViUR6MnAHTuH5pcsHa2v02HwmeKvSg28MgtMT5
1iMghyAHKZtRIHq6Q3fKHLIA3HfOnfpe5aJa/qdQmr1Nt6M5hNL9lcYN7AZvAWUc
1Wq2Y/n0PUgBDUoW/n7eDQoFMDPF2ADm7O79YCmX8s4eA5if8B/QdRAMDTUXBnjv
pcoKS/099CKDq1cvrFft3tI1aVnRJFwQqoEikmne4QdOngHpAAc9bvUtjXFMrmCV
5z6zO2kSk/jXl+HmjLyRzBZqMNZZpyWNeTt30C71oHxL7GFT7EPszI98QEHTKVbl
z9p1/27nfoF9eBRG61Q20YO6PsdaG6VHInujrcTfn3sTsetPh/PH+2dGnW3mGVj7
q9Lur78XXZ9GeXTCnM4jTjFT1oqEzmYPdnpA9qmJ/TF/mS1q4DF/KkpM0Ml/sO79
fpQpqcA4GS5LMstW+JhgxPt43NKcpeAfZZo6fS+fp7d2aJhcHIg1j57MTIGnWirE
9S+lPlyFxD5zCUcYgEoII+T8TdumBRsy4valcGA7ftD+JMrppn+URH3gKbQwi39b
n18f4/Q6sPyX99ofFObYJZcMtDT4Vb37703xuK23/2Vn/7DL3QBvBilvMDmeSpj6
ukqsu9ScLy3v7A5M2Wocgr3Vyq3yFhuK5ZdbvmM25Y2h0SdZE/yit+qEeo4nwfuB
qlDcJ2q4rE395b1R/NFHwjKcoDU+/OJ1Cil2oIcVjIiicR/basOQSRgh7YK3o01B
/Vl2VNkAt93v5EUQS8F3pEtKYIEgrhM1YIQupfHAZGDXYWV/KGj4Tyc8RLoff63j
j2EsifWoRTOBEtqj3aks0kr+RAjtMpXo3J80cIzUfv2dWxKiXQyKNPuyKhamx2uH
ABhhdZb21jcs5NgKP7ncDSkQVsZNAo+nzORJysgrdDb0MKoJ3VgFztz4oaB1CYM2
DN+/LvtSg9GGFE6yO2zRVhoXgeaBPHgeydoTsxDEXsGoU4eF0kBvRQyrGQ0pew+O
wjyzHzAyzKKDuO+x+eoTGlKbJWQG8y9OazNqLOK7zfdxbr7Jk5RVBENqhlfVpkyf
GFNcnYaM1Y7Am3p8nlYtluVYm/bSlV/EU5JUvKtBuZsITJYuJLens1Hyan5uwTMI
oy+CYrmCabjnI+Uhm5Eof387uOmB/GMtSt/L+TK2xUAphzvzLkOaLubX8c02u8aa
DaGAdA2QANTqVvObcjjUICUbQjMjYfjaHE7iv4rXIYISndh1cuU3oosQuvReercQ
Bp+jRVl9lgrvOkA/yx2qBFLqt4+25E+NJjrUetUh8zlmenzldTXkk+DjMf1qIn7W
HkUPS6dJLZ3I1XmWDB3VimCdqQazPwo6eVoKdBpHPUusPJntXhdiV+3OxeUF5L4c
WqR+MYdB+Zn3hEmWzLmU0gQGD+aZ41WVSKjYwcifT7rE+4zhn7m09/gwiRtOzQna
+eOB+jmeYq33bRUKuEbwm+sb+IA231txB5EpJdm0N9yfz80SaE/JQUGtwLPANeBq
q44C1m21UlfIrDIK//n0u6U9GOLTtmEzCUk7+JvsjzXTsRN37Db7amZIL8QOvH8a
CwPJnUnN/Tsu2vXLqJKa16DJKOAMcUl3JZ4h/WYGzldFuce7PzTuHXd6IXYlxBun
kR90+ge50u8h1s6vn9e8l1CVpbXYebL0yFzdD6/Ss0wgMf/KFndunWcWWw1NSz1i
n8xc5OR7XoPevZr8upIQZuFZfd69cefwqJXEmt0ajgLEx7Cd4G9Q1OsRcuVGeuNR
/HDst4O5+xtEgJOzbMDpAOn114l4jhZR0/iPmMnNoGVbQlELuzAHfLTbjnnOOiIa
L83NsB7ZKmvPTZp8kooljgYianjgh8QHNW1/PUoGIRxjA0pFf/YENj1lW6FEzj+V
v3XUbWjthkziopT16k0qlUsdWyBnciecTu6gwH2ouvLakN1eaBzRH5Z2EAAzdTAU
AtH/8taPH6bKWy6LibAajO9nGEU1VcimOYyKmv2ZtbTsofP38/yWOrTacromFhkC
pwHKMp3QZEI5CQyTijGefxTwv74R2IPPRn3bLM42byHVdCDcYI2gmbmpl405Gm7i
Zlt2u4HuKbKpgni/qRGNPop8kl44LBWDvuCKBZmWVb33OGSLPk9vGpusLpJAsSsE
XL98AKbQMIVqLbXLednoAcCyJvs4NjMnhjoEbbClnXetc/vKvKeuE/p18lZfUyjm
NFfyIg65Po7FlSORmTxadFxuBKNqwsR9u8OjcsMvbuZ1+Lq2Up5LaPgu2lx0f1I1
R1KGUfHl06rFJ2rAXh+Du5MYtopXavCZDwggZxWWnQMKcD54L5zoWZ0IQiCjksGM
18xAIgR1FYLcyNJ1Yh8S/MYDeGDtvED0tkCG3sIXJaxQoSASP6M40DhIS4Yp1rtr
jhRXLAcRZeiRz7Ty2yFX9tysJoo8iNu1aEX8MEvdP/w20ru3GHxEx6/Li1b1/vTJ
stXqMlWGJQXUIBMjrh+0u6/Qcrl03gDOW1B8b6QvyEiJHXjrx0h1QikAXIo1vUU9
/iREvRLKmgzQchS78tqZXC2QnVDiBcq3rE93YA0MGObiSXfFncNI0UEi29SrRmQK
9APc6SC9mvgy1rO17LfKHm1yFhdO1FWxcQjAybFkIpMJxMhFAmy4dIzT44nOvt/q
qMOF13e4cm4lLONn0dP5Qpo6bNIfjHCZ4A9rCRHvZynSwJxFMWqZC52Y3f0ZHi/T
Cfo0k3CSY/C24KwayC37so5ItdhGbxMVKUaV/yahKQ20250aqeUAsmMJMwnalVUW
YXB9QFg+zsZh4McXRC1OCi8qTd+G9CInhiQheNLYD/O2CMDjr0tCdlzbRHuFZiYV
Y2y37Cj/rdjrChhYVWM0sGYdBex4gaB0I+z0M0fvWlbQiwVTup+6Qf5poPiJZy2V
2Xf5QIDcOdMmp9rAuiDwAesodbjWUd4gVg8Diltz5F4nsqYaw3xNpdH8y4BKZHLE
Ia2QQS9FSavYeiynREkOC6t3S8+WDtfDR0iG1bqmkunbLCm9xJ+gkYbzGhi0/exh
5OvgBY9sjo94AG2UShrqqw4duE2NGaXr3fItLQjz+poMkydUDloP4SQNSsAvWl+Z
dbW8cCQTw6vVus+PfDXUbLumhiq9HsEh5VhjGDNi54FdKK6qfohWNN7xk5oZBj4i
QEpZYWWsz3NB57QVOVK+/EFAeBPE+/iINGU0qREb2/meplTLYuSQSW2AETgzjquj
KpMuz9wRZ90f4W+4pEIpLKBMHWnLP0wG3ooy8pOkCLspgU8UQ5+uWLUfp33+cp4d
Pi3C2T12uAQTORHWcPf3hitYNRcggdx7wEKgRm1Ie0pW2yqi2XpbFeLTvaw1h3tW
gFQu69VBJ+E1llCGDiBRK5GtgvqxFKWcb2FN+JXJpL8jArfnWSLoKjszaCU1PDXX
+zrRckMVOC4hqRVSpxxp1B3nFZZpnN36OJ8kx1rQnPD3VEGj2rACGGlbqnrKEr1D
PPBDKDyzqjZdUCd+eIDRh0RoQJZiwkLbAmvwIinxqXj75GrmiBlEo75ELQhRQ+6+
o1b85/+DhScpYHQMh1ssAbhE6rQQ2WNSzcdv+L/UBrW2wt4Ythiu0RAl04Uek/wz
AeQ3htCdpEjh6XgeYQRLkS2s5ec47MVXyLgHsatbp/rDDObFJIyymN27Rupcq+kQ
VabXQb9TggK2ZDto49JPt1axi4QmgR5ZC0AzYYXRB9s8Idm4+F4rVfR24tnnczZZ
wC3cddDRuTRY51yUP0BhjzGMTAyniXosMqnGcunPSr93wZZ8aAJlEVh8qcQIPtEj
hpoi0fcD7ac8AuaN8DYNhIYB35dLNSmHLRWR2YiXFZCJHXNaLasAJ3cm03R9hxL2
LCAV5zNsh2oFGN45EGdqKX/rnfrKLK/VLh8m0OVR/9Zkn20bZLRHaOvJgNY7pm1N
RqZAb9qzkkpEJ+xpQ79zmky+lLYyx56go1t+CRCJo3xGvmX95ikRKJsCRrmPJsQn
tlGQNSRwmkhY5yGQtsO6zRmJYOytEeILrl50FeUjjRJR8dWbg4WWefGHmYBaK1zP
eckozexMAJQRFcf3xyZ0qQFuCWi/w5/RC5VI5uqkIomV4Y6Hbxeg5Bj++3JPsRm4
FKcUlusb9QRaZQT9LR/snHfmjeeeSamno7x2ljVR6PJ/gBNOuyvsOjuUaHBdhLVk
1/jVbsQ6ZDGbiXqJEEdbpAJAxrqmlbu2j5cDU/NJ19ieRzphDytEPaaL8Sn16Gsh
1uiO0oIRSz0RC5Q+VdVzR0tIaerXD/VH9idDEBn5hBIJbWFP9c9Dj+HtlmI9BEmR
snKKINFTAiJz10/ukOw5Ueq+uGdMnTSI4fQacmmmLmrBGvgf3lCtmd7WpVhBxM5y
E8IMGadKBqnEWjillAZmOtiR2YG4cJ0lQ6sBNW9xbZfvHMPEAPk0izpgSZt8Jshl
iZPDf38A3Cb0Gs++62DwqcZqcu3SO+BTFf924F70rNZWuhdcAhOpevtpi5BSG+k2
P005/5rDcFExWUqFFSOHa/KT/O8090GpE7tCO4UEJMbrgDRY6cve+ZT0NkzEmRRe
/OXu3HDyXVNHMJPK8WD78F74c/kGWGIyMmhLB4tFn6/vSmEKgeS6Up9aIi07nLb2
dMMsu54DCQTYdVpeO1JIcRuQ4lROdfcjSa5Fofix0AdnBSI7um2kLJZCFo2gjxhB
wsQ97mBlcM5JHlzfLjxGCkylvVDwjHLGuEkeK8Ltea9TQK8lrKxIQEmT5gk06W7H
NwInaOcONWgYCUujTssjxyGbc8B61iAgEx2VOaNko1d/OTVCQ2vy4kusEiTlbGBm
oyk8XllSZB8uhtC94ZDWI4YbCghFzKx4XOc9eswaRsb6FEsCOxqngAA3t6sVzfnz
8doqzXmqKv7z2leudstfUKtcCD6wmrBPT1TvTHuRGsCdbACFxDAWe0gUXGhpAf+/
zKGgjHFqoTHhQQAsK6zPHqQ8dL3WTRRRvrTWUFdSm6Mego7kaC0xx8JieZCuxU/w
4SjOiNOj0U0RVNBWIKbLD2r4f4QqusV59M2MT5upOkN6Q807d94IWDtV6yG7WrpO
fE+R5wudwd8g9VzrAl4C10vzDaNHsSJ9qL2ftLWZOrWUZrZ6aQB0gTknSU7AiWGg
0Pu0U9WLq+OknnbYMFD39lukW7erJHLY9LJ1RkHmND5HjmW8M8llSTW5GHjhz083
Sv4iIHIgMy3f+RCQwIqx1BiOW8TNWGWz0362q7OdX/g+zkSeQDuB2MacxNDgDgU2
EzrPmooxzUepzhypG0YAmRRdBhTnSdgNMbF4WMTCiLKzw7iRyjoUUIbw6uQRpBma
W/tL5lSkm1ZE45zc6mH/o+vvK7SWIHeyXJmarRH0FzzLPPhBpCkbIUzABtEhQhCD
+T9EU+/XrLvwVQPxSRXNTbZwX83cuHM1N3UVbL8JPPXrvzN1l+iSfQytUsrbd/sf
PwvpS2JJrJw6YzwHy0gDgkRMxfS6DiDYY2jY8AI21UeV/v7T/73SVDiLpIYGaXIW
yUwEUD/VvASHhGekIxApBcc3+F5xrkrE7Ala+UTaPD4ygxTKgF3Dea4gbfrUsjR/
ANeanBQkgriDHvlFm8vQD6IgxheCyIeB6QA3AVCShtVB4Gz0RQUcJYnTjdTBOGMD
ho1OBh/IH/iIdIIDB/Bd7oBFDOOZO5sd6HFmjKYKaQWxYVUxSAt0paNbqgPJX2Cm
DJb+eqoR7ic+oyu/qKvvh6TadLYoSCyCp6jewnI8xnu1jMojjxnjsFxwV4CJqK/s
vXUSno7P4yNv+I5VvZKZ8h1RWIzTJOEKR6urqdx6wy6T1QNWnu5PR3SHQnj5Qfsm
+al7pJmxWWBrRpHAOiALtCkdIL0/QkVI6jj7ZLp8HNYoXvfXYvn4kbVvK3Gp+dMn
eN4qPsJ/ZKKBfxGvjtGUcAdbHgaooPVoVp0GLDfwAxin5ZCOYRTNNjcWXVBfLD6R
0fJI4lwRiGve4jUgv+x/ndOBClQkjyVz1tglZnMQfFNukUgRVPrmuSK6WtXRZhHu
QmGiA/1HBHjuOYeTXewJWcU7aNor0fudbUfYdoNeeANT+sYqUjbzPfhfxpNsTkNN
bgPQxhdkxoGkG5CNHsXHNXPRESlRRilEAilvHnP0wqji1V/4DlNwQQZmTXiwsexU
AKewjZlkn+fmEEZ70oDo3R+ikB9SnwE7zEawSHfHQgG0nGAqVYME/XmRaVhaOoSz
9PXALt18aRZ8U7vlFjKq3Ls9pBbfWJb9gXKQRqoyzM+4hH/Ixa027q77oGMut65B
4qA8VCJ9qNfCT0mAO/ZKoeDqpesiB0UofBgo3iezS/BIiEEJZIizmzokpUsF5Mu4
zujitSLpCDYXwjF+LJEx2CAvEgmL4fma5+tTk+hr12fEcfDyJL0d6angenA81nSm
whXW/8elPJJUxG6SwBkkD4RRA4Kkyki+oRXP3Kca5CGxjY0QwfPlqBsr/VKb+pxB
OEq6aWs5DXrcUNHSZE7jxJlfm0miogp9H9gQFO+FUODY/NaMBeGa7H6b46YCyeqg
+N8DlevphcurwwVvYCfXaJedr38eDX+6ZSrCZorZH/3ahX1Au6gviGVpjlctIQ1G
XTduOTHJIlPY2XJlhWZY2v+3bMgP8FgobJ5V31yH0yOrPHFxv/07/UFhLbsiCaog
1UBqfoNpeUs18ZiACDJtNCooEwXjHgGCpNnrxXZn4bLD94AC4c9JQisF5941CDqa
iKaxH9HiVjWlD1WQtBg1GaFRISZfWAdglWco2tu6nqcm3TMYfSLzJ9hcLqSiwBEB
Jb+2xb5Ra4xu+tmOHo8VyoSYgUFn7b5Aiz9yuqWlEos/8BpLfXdIDhfS+DBnH0LL
kWX40T5AzqsxWlthRtREQk/iUTAPUDOh7mQ37r6N+fae2tamzmzVONOqChed0QHu
aFzXP/P3lWC7lnCo0s453Z+BTslbLBdHYWGRDWPFNCzlfne/MtEh4rtj9E9qj7Fr
WAFxQKuSsS/TCYxx3tqb7tAyHi4fdPMb50U8U0ApT9NCT7NiPQ8IhV34FS4RPSi0
xyMcM46rHqCsAtYsVtDX1nYeT8n1M9Zd//GHA8b5Y//fJBS60VO7a5x8TfrG9bDP
1X+LIV/rX8RMBNI3ymop5mU63RH+NP5hCYZii1Vw97dA2FINBsFvph4Q8oTJvdRl
QACC8wxqew5ixDW44IHUJT9OKzX216RMtUChFE8G/0A6iWsvoo15UeB7sUYPIwED
KBV/yzlrhfUkCJQsVuxvaTMqPpOi99xAmzxuEqPmKOEuq3F5+qCeeVXATxGeMIbM
m3Oukh+DIVOsmWn/Of9HWrBi7j4QbwC0dAud3NYf3OeqhdZW/Ih+GssWIdJ8Kamn
EO8ek6+VfltfumgecZn2V3ebdvVqt1vEZaFcpMBFkvzE3xjMpwoVhZ3774XU2RnV
/17S5tiI1AXXxi5huxhc60nnTAv6YdcK3K7XlU6trLEkex1Nz5FB+Gkd+DIoaxgI
Ydu9j7MEkWNktfdN2tsBAgwry72iKNQuCOOD0WPC0T9MCNrYIm/RlVBgj9BmPZ7s
QPMTXP6sDjJG8bnkvDFOBwmiff+D+hozkPUiW9wqsCR/sUmYq4u6dJkWIBdskR63
/OK0w41zR5usJU24VbuWWSc7o98pJUp6SHBBTQPmFIMgQcLd3uoLJix11NpUoA6V
BbQfdkgRE9gmTSL7235h0OMw6MV9KySJPSv+pr1eFV6YuiiC4TAB4X+JlQrVXdOM
AaFdnskrOhxZGZCcCFdfkB/s9/GvGJtn5ejJNHoPzdNLp1V4wiKH55Xe3teGnZd9
xx1FyucX3lwMpkbINqfVjEQhMcZRV2qH6H8+mDN2h7DJV8nnjsTAZbMmp+2sQQG+
FunQfCYvlQDiVWUV/lzMpYFYG1xDKnEwexjeFAP7zCYbQ15hs0cGyTBB+0RuF8oj
immBdHs5iIB/NU99L04LIlMqxK+A9og4IJYM7YEGK5LlmRgjeyn04H+/SEg8UbI5
7LOVhpHV8X7R9ZP1gw6MR9Grd3JbaFG/dwiKz51nT8bQoDB4Q7nKMW50WgEeSLjZ
3vNeCwakDoPRWJ2yDPwmiPlrrikLjS3+Z+jUe94oXK70FmPd7N/iVX6a1OznoHV4
z6SS7RX4d1iuoPuRDn88ZHkTlKyXrbvh/uKa0PSwAniDzDCKs2hGrTtvEsoyreNS
M4edILKKgJBABaa7rY/DIyAoJCMnxOKFUiWLDmjAsLoBLVdVYGoSUw8Dwhyi+Q3U
m6x8e1eV+gNP3XMbnx6lbps4fGlQEr+TN2SpcnFMI9+bQ0u+sjGeY0henYHVpgFu
AOhxrIx9GbnLNpDYEDAig6paxSsAL7HTyKI6ZDqJZh1RRCvlcT0z0zITE/uQdyDM
f3nRCY0Q3/2P0On469rbYUT1Q3EVXJcjFEE8MHee54Tb7V5TflLrA/K/KAGDlQZ2
iVuQtsl/Kdl6lsqPLIe3zC3rJGDOYssCQoARXSB5vwpKLsgBKMNguGLOhkKzs+LI
lA8IOCaZ/yC79b5aMpNl/wHm/fVAUXNrsf8vGF7xDxbguVhf2w3BOnztvAAfGFHM
OiyP7CyMqrORJ+aD/6MKQfB1JUwLyf3U9nQvh/gH4TwN85Stdiqgk15OzjGhiSSZ
HO0hZ2Kc9RyMKU5zbn8NsqVNk/zB0fuciOtka4ygp/JUU376VEoSnR1m/nJBFO/E
QeIeyFcukTf0DvxU/uDbgcoCOeXZctIvQsYh58imWL2i+tYDeonk6eg4qSCNP4kz
QVkwITR4yDo9QdtItvRzAaJgO7zO8/hyNj8RNVIsZwT8EamEej2Yl4ogdLNf8AOr
P+xcBDFeUUSR7UXRDKaswNvQd75JwU7PVzjrUJnyfsCoeC3JfCBTvopyQMOSnZqT
EkAjSdSruU1xluudF7HUbGbtTIsWvdPZLRllqbRKceqhQK72fl9AtoWLmSefg9HA
Fhg8CvoQTQ375rQA7bS197ZxfqD34EHXInAn0f8d77VX05Kpz7GPQhpcQBApUHbZ
NhAUsQq4u3herSLcQchoF8vAslR4Wjp+N34+Yi0IsG2db7Zc1+KdCgRSRWVSgGSn
hFmh8rQWUkUxUnsQ6A3/qr4lIE35uONZw3h8eWQ8gj4HIWSlBrxZW3vJDpe6GI7a
kpA3oJk2hcldKwAA/ownPbM76GePRyZZqVkpQgIMgKryKeJyTYIvZbiZhfMUiOlk
tC+4e6VagEg2Gumgr2ovgoN9lv1+czRNiWg7c1se2E31g5q5NaErTxHNncctQ7Lv
bltJFz2fDwc0qPcIr/oTOaM76WtA13JD4bXLL0E0oZAE48I97TKiVr7LqAB/FsEJ
Hime+5nT0uXbn6s2uQYUZctYOwElSj0iw2gksbDLpqcOB9I+luFTajAYOCFmt3Ry
pPFJAONHZrLHBZ8JWobseosiv6MQ4vsVazRt/1djlspi32oJEWmJaiYVbbLRJ4Is
JiXYB+Q+wsJ57DKe7wfixftCRvIfx6bsmuVUtFH2leVbIV8uo5O48XNweyr5Fduo
XKmW3dQt4XUwNd9fH6TGNkXM71EKADV/4wy7u415nFmu5i1J2Q+uimUckABvZztm
gtUoanrH+DxdP2mSuoBl54KGxaxu+Rq/b1/YkOFO6CYZjjeFN0rxjgIt75cXghGr
Qvo74P6T0bj2yW7pCWzTidga9npEPJggCtdSra/wOtgk3LVtS97EeNDf6t7/98U6
q+9LLuvv/bsMPD0GVSN9pzG8zC2jZ3/72wb6NJ0NltcTKhTt5hctlDXEnMQkd74t
pXsvoZRlSDm2EwrKLFGwUvNrIFZl4YUlzMFbQXPz6tBHdtyoRjbka1njNjEzCtlW
XJ6yhrTCIkEudEpCrR1n4shGKxw41+ihkFsr5EAVCBIwIiIACifyWJggBLl2j6zu
yWvWfcVSEhftaniIZualWbew/CpT2iECwoIq92zyGvLH2NT3iiSFFV98/vKUCTcs
ZgZZfdja+SIq4FSmJU73I1TjLdJ+bclVO3PB66SUL3WNZ+Pb0X2YZIpNWiAtGbP0
ux7ZAnTvgYHY8fJec3XTndJt+I5HSbVulF9npHkQhqadhNuguoSDBIBVn3gQdSaj
1ANVhMj9idqhRxu8Bjp7M8uJ6v08RPxUEVDxKzOzRVxZeFTIujAnDDj6cQhc9Xdx
SZQBOoGFN3x+HST4omRa6ydQVcRKgJkgFtTUQTw4vsypHVVQ+TeqACz7NU5xzlwT
tZ4Hu+XEWafl/r5ynHj/2BypGWAhDxCn+WydFdh8qT5N1XvDXA94ZNI/CmOKDTjy
NmkUObZ6xLE9TxpWbOemAU+EsuJHTLyvmvEZs3KnHaMFynz46rFYwMDyjlyO2cm0
e6IN8kXy2TrW7OlNa3fNQy9b9bd9BKQn94TLUNjx4sT97DAJevIkRoY4qKwP4C+f
P6plCrLx7Imsw0ia+GuPsOkpdwGyWa3bTIb/c9IHKejHdB9JS0VYVkA+C405zjW/
ITDxgtNGbpRjzmcv4r4CHjN8ZOxtv7Bz4S8JhujyzADTEgtjIcYm/MBNdsqLVnv0
mxk9J55HGLuUkiVfHZPlVVAsEPYtV70r1l7iQes8kF4D0MttoSVfayeTiPKbiIL3
QREFrzhNZvOjFoR9SaY8+qePymMPYhulw/eXWiDePpZmccXYPynX2NlEvW0RHi1C
yi4pYASU2zuCBDgoedldFkkD8xuixOMwI22y/jnWsDJV9zrqJGrL/F0TfMX25kTO
Sec1XJQdcfh9f6TVDsZCy9mGATgeQFrDkeldU2uwW468q7f7Tho/P3Z/jtXviCNn
kieAOF/y4kbysZCiTUCyDe1GRUAu9PdRs2+CH9Z7LfOZTbTH0BhpCFBTy52FbzPH
I83nigWTog+7jo6Atw5qX2DpDWuhCdyoxL5XaFIwY42mXaueXtcR0UPhYyvYCw6O
O/apwsTQqxlfIe6T8DUz8xkkrYptFZJSnNQjp+6dXRdQoULEuBqFDWPorkxBQ054
DR7Dve55IXLpsdwuEV74J5v6pddKJbXc3oUoXWwrJ/WFqac5aVY+hN19KQ3E+20s
mFAM5BuGbVWwruY+CDtP1BY+8yJPwc7glhu7a52Ka3UHJlRi3xn752dyqk5vFrmF
zp3ty15xfWDjHINaafl0zqjww+ZGcfbHJl+bYVy2tPk0NIH9xKePCreIFD8tEC02
d5RhGn67YMyxbGCXngUoqJN6L7nX4TYa8OND16PS6i7OEzCI5D8BEc2CtpqT7ITy
8nWyFKEHky8KqvKiBraIIQCm11xxEnJPOmf5g4UpmYyxNn5UQQ/UiLl5JUwh60Hf
wOUH8T3l7OV49wws9uO/VGiDESwqiCfL01vZrMqMoc5J2ITIN+pdKQkGcNqBbIjC
pX8TAuF+sNiJNDMDWcbpCKSvbNxXlJisDvCNYTVDwgXNxkONWJEkpskhpTSzu+aB
bp9OrujEdpdjTnBV2LPeMxSqlsV36LJ1dFYEm0jrVahDu1NfsRwk1IN2vx4ZC4iQ
Q9hhqkzFaYfLnOna45/YfIZ6zf7+EmoK/BxU7kCX8iTRGBl7vpLyy/B6U7wEPzlQ
2xD68+9ydGX9yUXQUn5baYSt9DFues36ARx9gFZGBUMscrXMQdCjSmQtV5cLpNQ3
cuDdZsUZcmf/vKsMa4N4n8XnN72mFum+4JSYaRt0IQ0qGQcMmAAw8e/pB+1adF1b
+/p/JFY0i6tZdDHg1N65X72cpvDN/BOuoWmPIkORFKcrC9NKj0nzD5NnXpIO55lU
DstMjNVswCDrV8jYVwYg3Qg86TUhXIEZDt2weyQHcFFv06xUGOaGhZDJWAAVB4K7
Eo27rrW9VVbafSXp/D75ZnJYcz8/4f66n58atxKjzLf2sXchEhLTyojaNzrLsagF
BAfUGmMGC/7SOtt8+WEZ+IxemfsOlUJkVz6nDZNixZ8YaqMoo4WhvfkU5vIU7qRB
RFkwV/qX2nzWbfuZb0eMxwSO1rOZKItyIQVVfV5qwpt6iJZXClKKjvgT0OP7Inap
RAx2eHZ2OY4gM56MgZ3cSLZFxOxVZmFA2daBb+HOUeCAd5zKnzZ3DUE5gAVp8kLK
NS0/z8uXQhqFL+eMyuQCz/XD4jVx2Ke9hyqaVTld0QALGEu2uHm3FEyvCZGru+Xg
eQqRqZr1Kytd8ULoEeH01sG+HCA8gq2yNR0EBFnL1/uD/Elw/1juUYrHpZT2XMUq
KiZE82Z43aUi12gokt7fcunCFzUluDxcFK/l6Gl3qcjQExnNz6ppeK8fVrTI2oBy
+WbNfVQcoPOaOx53UqEQdQ6U3rNL4ilE9kq28liMG2XGJX7AdVnKdpqAmsCXpn/G
WXEHJajrKiWqdo25QTIpOi0+jOTwh5HcMvXl1l9W+/H036BMcsvj17s9JaQUsF7u
t7EcAFBltVXhJemE1s40TGhHuF+okId8+l0Hamipm8Wzvof1OMJZhT+y8gB7/1hw
qjIrMUTmg0cGl9XGRoszw3PlsUQkDt3Q20nCoPyODtz9IB13zq2jRgUDt0OsgoyM
rdHxkhgRVyaCjOsPAeY0VjN7f47jdADtxBRI8R0ZdAyHr0s+FrNZ8R56SqoZONpx
SWL+VhAyLvbIOF46j958zq9SUcgJDzNx5xKM7grphxgl9q244DcxAPNJFPFofYf9
UGpQl/bTRFoA1KywuR96C5MNbCYaEIv68dn7xHnfjosDRvjJqge00A0iMLXMoQaJ
X4jeyphLgPa2cukoyyqVEbSINyrnlXjGr4/w2+u5+SOZ8WueA/H+I+tBBRKdzNi8
C1efVSoJKbwfiMzDZq/lYB9ScUMRTbP1g2wjWE6/wreaXtQEwtBfSmQ/OesFVsYK
j2SGTTQaxuU8FAdi+MiqqDZ2Nao5Ts5JiE+Z9ANj78O0D6YK83VD+CFvvuTVpMeE
3SHrHtyD3yPGc3MEFOIdGq5wc/9APLInFKYkQDOjZ1r7z7ZLiMvkDuhkUQncKEQP
rBq+/rskYDnznOcAJwb41MAA2JKfnzaRnjdvRnlDPc9ZANur7fOauDFsWN52gYav
18ahBFUhTBiKvHExPd4gXZ+gGc5M/GbYQA1yqwWCwaWWilGzxf5vQozM+00kVxXN
PC1Z9u76IFLLw7Mxsos4Ou5tBdEN739qdzePEu/74Oy6GoJ7b7K3JHM/vqPJGEs4
LdG41UGA4mYLPDVIbTzmkk8+cpPtF0FzC31lFkno4VvQhuw+F2w1NXLuqqa0hOwF
OTCyjrKUcBNJgI9waPSgl3nUajBhmHRdJ0w5z9nA/5cZPFViGD3oE4WFFS5Nvfnq
Vx5Z3OQ/W80AMMRbFMhXA2XaiJ+pBUQoSxE/lOlrf5P6650RgnPdmvB2fjhH+KCL
DQcjZ173NtA9D9d4yxTceniFt5PWQOb7RC11te7QJisoZZ5bIrfBjlYFcWT3Brde
4UgRYwuTMdD0IqIE7PpgSg2nQ5wSP2FzWTF24gy5ZidZpzSXdmdzLeN+GerZvZ6w
oxMc8ZB4YvuvMtmUi63fxgeMneW8iVe8tahUldYzbHRov94cUqSN7hlSmMUc5dlR
Di2ckVUmUKqtcd5/Mvqfxm3JUCmjcf2arv0NjzNGfsLaT1qRjK/koRTgD8psPuNG
Fw/Tf8Z6GgXz9BYXGTwwwHQaEktkPKVVa0Ez5TuKIe8Cxw/NkwgfyXy/viO2/O5/
eYCTqz5v1smLKBuJ/zj3BbK1AXtUb1YVrnmLzvyeWU2h8l3zMnSohYSC6+yYa38r
ZFtg8XiCIrqOkR472wXbut/aHZ/SGxGUkSK2SHTJCsLB2SUDYYMHGK2PWhGjoDXo
e01SXoaU7YVsHsr2URgPF1Ej5l9X6fPwlCM9Bf5im3+vghDe/YIqgSFfOmo6Z++s
9VMFslVczCZs9YTnv0TtV20aDx6IXY32JGNMm93LlQDl767syQMvCCHwh3HOyr31
jrIOsnW+ooTwZRMNrn3GHFihysiTGEjceZmK5P9hSiNhKFjXLkjN/JlVEgjDfjFd
BeJbFUt6dtxe0vBMChwTAXKv55dnykx1SqE8XbWKZzM+kIAWEaVuK+dYcCWWKkC0
2PNFdtSQlYbfghOFkbH9XQqrL8BEzQ3s6e7uzTQI6bgXaL1t0HVJVxyX0BA8w73b
J3hM49GIIf1B19uHCNt0PWUFZr01v+TmvSLwi8vdqURFugyrt0WZXNKcyvOY9GEO
V4VD3dCPKugD9VlG3HTHxAF0QWQmmFETm2mpL0w6NPYzOF7j0OPq3ONLTp5S77iO
X/pstLG41ynrEhIfdUoEqhXtpMbN6KmWUTnZe93t9sFBxYRkN+UMOE1Y7+RCDpby
ME7yG8D/LAa4sv7kGJntgP9NY/1qen/YqYJm64bGgO67WmKz+VeTUYwR1lwdUCQS
8A4oFgmoavZtUPfRGKpyyQ0IhedjxOMdCFJg+Y1gSr7Sr80fhNmbRdVL0Ce7RfLO
u8aflOxby4Pzo9xXTAOvBDmD6d4rEyudb/isTken5twB1lq1FnaaaJjaqe9zufwf
jI63NVozwfE/UUB1+FFaZxioOSpgbbNfKCG6k/lNWBWvegZMnhRbQjxWaDvX1TV+
IN3yNOMOWt3srxVUmuzXzkaaYN+CoY63ZPpWBXbmLuKP9FwaRY4x9BJ82/RyUo4i
veJvxxhCf3Bsx8QXnewVZwfZNf/2QO+R67izNE4hSO3Mp5VTLndAj+3qL/KSrrne
akbOqZn2Ytpz0h/VzlzOIyOO5cHIbSCyTy4NqrNun8xvaeXkG/+zdRpJxWO2Vpk3
k3UUyKcKTbebjZjSHYPaAzsxIuPxXiEHKeuVAxV47f4mszwhI2UcoWE2jCWs0ZXw
l1hmLT8j7TN+QbcbRRoLHk8oAMhTwKvrWy6jDF+6rRYMz8MjhATMrVjoniDvqMB2
OQZb4a8GFJCYQrzu74Gd+9iK1WeiHXHBNrrCM8a/LZsHE4wSsLTcrgFYjUb5zIUZ
Mj6YAfuRAOl6qbVlxsB2ivJ4e0qA9U10+kLeryc1q7fXgznBR9NF24brMojwcQzN
j/yS4LUB7MJIquOzd01xAbDWMoVZ2SvlEYkLeWdEenpMrDcjK4//UQn5m6gy40fB
R4WzxUba5PyslMm3hxJOxK8jAhzIPwaA5CwHPcLEMg7XmOP5lxL/4fmIikgk/LfQ
vb6Ebm1ALI2ayKIffDDYVrPmCXU4ayu6EvQ48uBoLLtc8mjqVug3/tsihpST/sCF
p2W1sH6EmezkBHlXhuG74kyu3OvaOLwWTxUV1DGB0qS4IgxPBgejEvrJ5M2dgx4O
6jWORpTw5JAW1bkvR+rflB2ZAlSUA4aQ6ZZlpvDmlrgnblmCjwvcel6OuestmTSo
iBYPJvXA8MPdWy/AD9vGU4HqbJBrVoBkTw7Bsj+206K5t7NtydynNnqG84jGY7HT
At6XqVsCmosdZCVwkfMM5cV8aM0Z5Z8/bd3LDheFx6S+KFed1+/yKcIg6BSFKOob
4KUZ4+x66CvHAgwC5buh2XCPGyTsnsFAYnEZ/ZNGaTKsuIS5GgvPuKtCWgn7fHHi
JV622ZcO/dIBnABMllBqQcY4NpICG7kamWe0v6bGjzvyiFLkdq1OY93F7RIYOGPt
7zM2J1LAO7EnL1H3pJIn0Vs7+sGgmedvDZ+idvlWUmVYTfz4e0U8MzXkQfYBXaBa
hyn9UOfK2otpWZ1NT/9Ew7Q4fSn+i2ZnGKt37+/2+SLW5fgH78CpacmPhpvyYd7t
96OBBmBG3MyuN+L0wWgQpBgPrXRlWC6sNcM0UBQP/xwoDofClsEbTT2GSVr/VcOY
1wEM8xXj0kOGsMr7JIozYqtMwW6VLXUvZMVdkhPKFKkOY2TbEAC82IPW+KdxqGaV
Y+G3cecQIUzXCyBO1g2X+Jj50Z644OPpPS/n+Z0JABOviScZ/rLjbmZqzG9YfBny
JDOnNpvjSVaLCj48ca2k8lQdtIz/DE/YdIjRVSfEnZqzFpkft086GzYIlSSNRdgz
zbCestVAQMTPOIVngo7aKKClrbPBfuIYgHhfVORC1JQsjjMb4VQpKLGQ+pZDrb3A
EpV1VgTBzGppooKqwLpI7jW6lQQUVzzBmTYqCgqmWNu0gWkmnFmAC3J1RAuT8xBV
Xa/QqmyridLWolAycnSnPcnLjuAh1V2rQQqISMbK/DDq9Zek4VS21wHkTurV+i3z
7UzRj+wLOkMMvBMpBxUEFffrMxGdPtW3xj7yiylBE17Av+a2+IlBejRruaE77a11
3b3bNIynTAkRMoFMnvjsy3vZEFLxK5ZOQkzuoKpdtdDoDx7gZizdtqm/n37ZtBkf
PijHrwmTdR9FZp8y39JWrkg7StOSUKvE8M1NQosnSPTdNM5uL7tCBQR0wKrF5SuP
H22//jCxK3cnGeXlEgRSU1riBUnL1WxCgqBRjmaGCigYhVo1LYMGY6xyqp/4XIPg
qVgx/5u6dZKrv11qMEyqlkPB9l+z6AJzDA3C8YnVIPV4uee2BKut8FRotCM4Vm3B
wIeaeZcslZJ7ZH0KzAFOWKxyTpnOv1tYgwe7N7uP9Ugouv2SRkza3gkd+hdzV7/H
/ODelli3toygcreZKl9XYr1IF635+gIulQ/6qEEDu2R/3rID06anxZOr6Zm5kqeB
+iAF1nI173E+RPrghdP/zck3Zt7t779I3RAqt6waibtJ4ulYxgyPpTjUSYa5DcZc
oba5usmjoDPYliiYWHYBDHc70ZN/q68SjhWSFPecB5zXm9STZ6JAOI2+5W/Kg1ab
x87yYp4QBS0bGST9WoFpuH6gI+INBaWqrw/GfV3Y4isCqm8WXvKjic8bxTSWVuA4
BOpYvEaA9uBnvVZuwU6Bi5nFXFFO/RYIoRJlj09v1vzG0EeOM2EvNawrUqXHJpB6
80Ftrf3lcgl3/N/3kNBSfYmArdPsM0VqgC8Lh5mgA484HcWbQ+ePtnAuQ3Q84Gzk
fKiRKqFve8YNyhBr6pChSnwUNgpnRI6b0K0SE4e/WJ/yjUitzW2PqBNSygl0FaRA
bYjS03QT/Ne/scyyCHlLzClFrPglqbLGoaDm5sfNGw2rJrFOVhFsYlgIk9smbeSL
v/e4fsssWXPoKCmZqB4hyPZdJ/R82I28QG2sdVGMEcBEjvfy2ae7eHpN/ILpmE7D
DzVAM9evkeCYEDlws6cu8fZ+dzBCS3CGilNaA85df6N1f6SCAohX6XsD7QoZpf8Z
VKKjB+r8ulcWM11lsjVIu64GPXtrtKKA+pSeVgqZ79dfOe3TU2GVfo4VtuGJF4K+
kwrqSRJcc/G0o0A/iS9d/eeDVuvkPDPVQITvqZAswxLdCsVtjI0HSuUF9fW+Jtl/
ZKbdsh8PqIcz0TRbjf3I7DVyuvA7OnLLPBM8KdhxiQVlpviZqCDswmJgWAijhT9r
g723qdtWLQeJmbm83+ZH55CPElYAZo02jh8QlIs14nITi4Gm7GODMMI1jF2qhxLq
R4WQHu7bFc3nPfYasoJYJbmBD7w+TH1r46pMJjEL73v83IEqCHSOYjcRIfZoPlIU
C6NMgKcBXalJ/A0sENZj5i8GGqCchMGiitB6UlpB/WMPysNKeLBeZY5eMGos+P2x
/wgRANRE9rFSn2BfWP4lBlRY9mMMbcBuFtQDjgBChB/l/w0oqLExcPqV1RlewAgp
1aIL3E7B6F7rF5pjSjUfP8hLds7XzoeAcl8Unmi33ZzDrI2dPXi1KDsKQ3q9jxPn
hM2AYCVy6Hv6YNPaTPPL707C75Fv3F83NJQ72vd712KpDAKXP0JQxRfLAr0gj7aw
JfDBwGDy1H06rxGg1Zef6Wq9SJTDeek7xNXAYTGNjPIFoxg7YpamChvCJ+pYprNx
M8PLcwmCGBNvIYAeOaBvhiYxNxT5VpbCGwRoONunTGTqSS/Q/adKgt4Czw9iUn0Q
Tu6eR8h8rPCbvxqX+f/+mJhgZUEPcWy3pP0FTj5N2WGXy7yH9BJvgH0RSCKCMOhG
0Fy1KfWPhv3s6S8DOnDurV1t3dnKrVAgX+5y8L1Yno2oUAIedz/4uX1x6o4+1qTX
jFPg32rI+YM6uWayq3Ei9/NXUhOg7rWi4CRDZVszk3059j6RHI1VhRU5h/OdE4bG
xU1rx6W+XCukKGou+Duxz75Ux0yalgGl1uVeX1adCcwIhQbzCM6MgxBoBpgwASlp
X4LkVqgWkjF4njuBc+EfPBz88LQ1qZBIaa7aNWW0NSZlkyq4jph1tCQbu2L5Wfm2
IALXswzTk7T6TToQNjQ46YAuM7ud0xpgaGcNf7bsnaAhta6t21QP0V3WPK/fpnxQ
snZBUPx7HLaKedT/55dZeenOIIGwOJdDzGSW974ytlGQUbPzv0OTEUh1YMQUwkb/
V3klLiv8MrcGCwV6+2WGjPpmPiqDEi5FC/gJVTIxUcFr3CX7s5+UH5mFnoW4mUOu
FvBprELVexZqIp4H5Gmnf8jdeisZ5w4T1D86m/IAZK05IVvY4qpD3L0AZGpKtONE
/ugwYEuK7EcsR6QPAPqfHk7i5tMHsnn2H90M7xHVb6egEZ/wmuMKFPni6dlXcoBq
c5t14u8dfR5tFf79ZjAkrcLjdjOs+IFFt0UCdqJ90AWcdDku9RmvQvkBJ9nDrVSb
RTnUmom676NYGNXStqHPwyoQojCftlIJ50jdWy7lI9FMSFodv4mhOEOqZbBkJiHs
1tuhuqXeVtDVM0de77mYAcoy/gMSljQ9N3N2zLnnUPK9ZBfhMBa3uKTdagKWNMoe
NaFwTeRnNDG+JqlPM4z/N+KshJrgIdf3JNpgJ6oK4uyg/LIVAwGJihAS7dii1nXO
X6BW8+SeI/46NdL34tkNxl+5J5qAlVqvCiDIVElw69KVLcY0Q8LHRWmq+InU8zUA
g/bicivJgw3EkuikFFP0Kw07KuuiYjp482skSWvdL35/1xWCPkx3nBVnJwyPmXX4
v6r/TwBckl9hnB09IfOAW7HbBDlu7+qoc/HYTsc2OU/OD5cZpFht3cNhUiNSprqL
RGmQ/2NXO0Lsm6VOuHpnzz6aF/RBY8f6X++9Ebikmw8b8zqNKx4emTcf7NXSw5zM
zCkHOKugGucKkDXtTScvoLRHZY2SsOPfwLnPDRFhG5QxiK4rfrgNUK+XjHF0dCoB
AmMiY2S1FioPiJ0ZIE+0fxAQFfxa5I+PSzWM2woml8Wq6RFWLDIUol9uIM3NdDwC
uJqPB3ctTvsVKQp9z2Rl0rubukVsN4/0UugMTLk9ztlF15uAP1j/gZgnFwJABumA
d3sCV0d9IYyepFHsO/ABvTe8bybmDENFeHDJYeVO6kPQZoSGfwb6LUkdM/e2FB+T
PNfCsB/cuYDbFPQ2G9ewZ9bx8EmO0qDI3ZlHIyG12C+CY43R6rjUOD1eMl+Q2s0h
h+pHs6JEc0+3qCVt3AxUekDl64wMdRD1iIpnyU1vGPdkzYpb5XpcCICMafpUiZD8
kRIgjRzjtT38l8xZActdHd694dzazM3sFGzWP5OJ0wfzujKGRzIKzyOvBniSINZU
oaZwoN8OCcnYq1R1QoKw2Y3O9lQy5Vc1Oj/rgAFypRES96NQbocAFgLH63SKBO3g
llaCxM8wYbw9SVaxGVOyNZWARn/wpDP3YbAcJQ30bh21RMd5Hd2JCtP7AW566yAG
sQayxvpOa18FizWVuY2s/++08FOm/ztfWxaciu/4mDzUN0FhWyrDuaeNMO0oML5w
WYzm9/j4ha1MyPCe35zNAo2cXWy9uIr1Uzcr+bI6P7TCLmRupBrb+Uaxf6qY0wee
Xk9RC7L4hNQ1RAj1ejVaQhlE88hDY3plcIgB9d+2trqiQGum+7y3rJQeo1d6XFf+
a6NbLAV+9JfJsU+rzt+TneBU9h6cSc9asr/3E2zI7jHoQcNKGeowGBDK4N9WMijt
efqlwzUDskRDJR4Q6EkaT7c0jO9V+DD2hHZCe3oHG8asEVMOBTypsJnOeoiqoRDX
aEiesqocjJtQyzbnv64PUJaSw2/zSFNtQhaoVXcHRnHqUL7bk/+lab+a0zi1WVOO
ZpBMKXWXXBnzZfaNO6ZE0KPgk6iZWheRYE7Rq+40bqkw0HjwM/ayDflR4fxet6Fg
0H2P2FoqjSIbt5Req5Nj69pw44UQ9wWCQ37UTchelf0zWdOicq5uOucuCsa0M8XI
a895hFEpP0l596+AxuN+Uj6cWUDcozp7EcMZEaA1JmT7+Rtv1QotFp/85mtM4RIU
El4RezrcZDYsDVwQx5KGiUqJq2vuT8vbVtodMozqnEaPaqeDjwUbL/Ufiy+iyXfX
x2sP/pUu1p8qeesbWaEjD2lMEiv4/9qZWA46QzUWd9X4c2iGZlwDqSr0iSK9acZ6
EeyF9aH7hyuHSQmvJki/qX2zS1uYdLdYrEC6r6wFpruTBq0fqxQoQUZHIgry1H+b
ZWIjTl/9Vs7idCuuyp5Xk628T9D6X/8sBJT9KWz2SuKH4b2FuxtFFZH02o4dbKdZ
4b2GRUbMyMyJNWGmE2KwP/U283HvyHtAbUt52x0zAUMiq1sy8EF+kO4DEtmKTUsZ
G26onhwWRy0D2oUSRTRUEnEdDwNK5j/iM3B6icQeDSESgaO7/PgKxk6/ofrpllqy
pCj3mnKYwH0WMhFmI0v7KH+IZBP0xHavpL9ZEEwzeK6pPOoWwDPg92nZDJw0U0i2
a3hOWIGpTF1vqbdsQAKC65bDOdjFsPzQfiSS3ZrOyHzrbspIJ7gYYqF9mo6T6tnY
rQhtseeuYXeP/FY056Vzhm+b+pzQKUqL+fmvH4zOeaDDKwwMA5QcFFdWZuR7dERa
/OYtZhMRpdBSxlGx15mB0fTgVb3ZOG71YwjIAw08acz3lIHF6dmRQOzMEO8FkEAi
3ARJ3Q6JYRwfNCosPWBMfZmGEnh7nZB7EXlJCNQ2aLJLbrMkNpmQgyEAPYSY54ea
RismaOQVXGmVFSnl+kwrMHY1z0D5kaO5DiXOM+ZJjqWrIpfF0sx0bAbmsWsSvFUB
/PggHlrNVIIxxF/Ziub2MEjDUfSehho2QvyFNlk1jAEEuf3dK0vCRMadfNwlyHGR
/RwYQIuPNMthuC1ORa0NKgMyoCFo39lbnkvqFkBGJyxDCoYCpH+2UkJRxdqjmQCi
5W4/carL7IcMjOF+NJ7IZUgbZFLJKWYTARNGbuY7+jPPHXgLpR2iQ6vUja0bxLsS
DVO2pGcfIxcIUOme+Gj9zBKzdM+7YwEHQ51r0wgZQmc1J1VbPofFPA6ileSJ/Ukg
THkjU+0n/vAORospgLduaZvkjWPFAHiQJrKbHNrxvOqLpLtuYItVE3ZWgGEZE901
FrBhMviCLwWtkN56sCXN93bylBmoWjJlJpr5IK6kHMPBOINu1icpDWGoPLmKU1jS
0nRMcikuKTlNDkSXefb3CLmAdP5ku09br+WhBUM0DElNEeaV8z/n6A6ZXp73i1CS
uebNukt57eVBjxxavlS8dyB3u3nF+hUDC6Dg5w8YTMK8h1fXxIO9kxQ2IpvqeeHr
6RUajjdVQCpcdH5MsrFRbzDyFT7VyL8rmJtVycdFrOFEsTxW6iS0lSneMKF/Gfkj
JTYOn7xHQXbWt/1U1lJiSuU7j0uTAlM/h9s8CiPu+m/3E7oEPvtXoNAzdLdoxrKX
EjIRnEsRf5fu+HDOdVk7lE3sWWJvW22fv+CLySMLQtO/9KQd44LM6zNo0iXFTFdT
cqN2suDcUjpPSgndiSD28l2P2MONFclSXsPPhVSxkQnoxDmMFg4py645YD0N8Yze
upREsP/5qVoYuBw/q1fTgU7iqOH2+4Whvv12tDLKshIW/zzMfqEecxxATZGaUGQo
qkGIw+mjHScJkFZlssV5j+CrH8EQh2Qp1eEnbV67VBe7iSkWuqXKDKO5YGl7HGbQ
pi+zpqAfeyGO1S3MXOvjzkwVx3DHLfqvi/jWjZNHcFPMgQhHsqxEWiGm71IvIIWY
6tBq9XiKufsflgcpf0lesKDdwbjYwoGOi5YDQi7gbjZdAhGqNagjHEUV27XbkQU/
hgZZCMK/eb0HRoyjTJdIScwLw6ss7y1LYVumGyAq3UNWr2ovQUJmyflH5SjZsS9w
1DHsmMmftAYi2S/hFa8sLX7mM+0iVTwpdts5VAdihabRTqPxAAdccDVi7vqpD8lj
W+WngylUv1LFKh7fuJ1uVrs7TmC5mrkA6ZlRQzzzFCDEs/qrxY9ihSzPbamfsiKZ
rk2Jrf5LXUDbGZbE4QA7vLnP7BZMMB01oHlT4rdtf0Bs6/n/PlBNZXGGGvq/YAWn
Lmsl5PKxiVmWJlfyl4dve8Aab5Y0ygEZ2+rVI6vdB3VJUPwEVkS98Ydhj2kkH2Hi
RNIVbLEPl8T6SEmIwhiyc3p4rgoSa8WCwE4N95soFp0xtA4gbgx79EGpacOaVNAs
X34McKxcMetvjkldoJJhgKeW8Zdweskuo/OGDuI/0xVwIspO5zJVszOswWzMyJMR
HZkZSjz2RSUZgqR7tcvFCt7MJLCrlGSrXRqNIDPQPswNwWYJgNtWofRuFQuGBQ/s
AvHmckI1Ycsu7Euq281e1wRsB7fM5zHqnVHb6MiXpp+MnFodhI+oiTJm/Slk+/dy
efIsGDkhQiFXGKBsI8506vbwzqqs/2bDyiVZ/cYF7eDQ+vN5C5SD9iRq3TOzHrZ1
xrobSt6jJCgjEhtmiLYVKicYX1Cv5GGZ16r/8fOJjcKz/9BxyLy5YTc9Cgzo0aqI
zam4UrKQh9PWNuJgLHPP6v0VTWZjJNhX0ZUj0cunhNulS0v8jnIeL2Wt6q/lpEBM
mmZazyvGZi6t26PNOi8BExI5Zh/hmBypE/xw5ieKqaUmmUGe39EuZoqQa7CNm/fq
DawrFg0VyjRo/74Lm1J/gsRpIuKePgzx2FNU15kyUykUoAW/rkw/07shQnc+B8OS
0vnMnvA3pwwZ867i+3D/2pQSTCsI44LcNQjjZMm56FqKDnJJv+AjJ24RqflNL7fa
yN47bBZkxyFiFGAWQpG2jT6KznA7Mzp5PqQX4nCd7qqLkYVUpbUkpyKLVoIO8Uhp
+UiGlgYI0HFZMXLGgWvBjz9skyNlJ+YHHEPuosDdBIDGL3JVVtvh27IN8Xf8Wsow
hCZI67EhabVzKVYhlLY3TnunbK6jxyHLJC36BjDPgHpL39PVJfzRzC5SFqwMJmra
X5eWJuhRZ6g8lXXIJ+Z5w4z5psYYQumQjrhJOVTJKy4Z9IvctcXk/fGqOGrHayfx
s00W+hozhjK0Ez1qxoS5qZilRm5HjfdQMnWvTvHPFTjlUp4orNA2c6R8JVeQMKOO
ObNLgzCHYnOxclpX674zqaUcLXLm+wF25uybVZXSFsnTfb3wFG4Mrhfo/7URw20x
eK1ppRShIt7Y36hxjAuq6+YZbe9Pn87gvkxMRxHtoc8UDmU8fK5Y7M6G2DHtSHXn
GkpGeadji+NnVp6oejfmhX++2eWmh1O54bqZfPR5DNKUp9TfeZLeABHdsZoGRgPF
jlvb+6865AzrV1hC8BLQ9fGXkflhHDzFksWjYk8Oes6Nw593Ky57yjTx7rUSIcXh
uwhcHussrEHePHNBE2fRM9Ip6dqt+7upvnmVT93tt6Tacirme2hR5cOO+BPt9JwH
A4rlnINtQvRTle2COOK8Ljo5OkZR6n7gd4frfzWjeCsgyIG7s3gmyQpqameG3MU+
eHJuXOCZMejkjxmR1xpHnk3cVsoMGkvAJ208gpV2/4MaLeI6xTFaQMt6mVyEIUhT
R3J7InYGqyzdnnRZH5kWv9I64tgFxCKld/D0caerMoM39Im9pXXusyGEx8UWEzyR
ioQNZHNerbdewxDORGVzHxASKVYwp30QAfu6pH9CRw017Fu5zsh9BZqXuiGRxVTZ
Nj60js1IXw1esZgj7vJDqfD4kya8C2Ge/XrCe1Ka1vrqfksnJTj/i5BtFOLRaPtM
irsEP6IfHKd5nDGnVOY0dkzXVq2BHlrtGi3JpQwY1kp5o/5XcZbrHFl+LdTMXVu6
QE/v4gZSbuADh7HIr1Wvo/uRKYWgzKqzgEZAYQV2PgLhwdotg95OhqwDf8H1qPth
g7VXWxtjtr//GhCJKzFKmU+f7/4Ay24moou6/7pSpNfhcr+j1HBe4t3bRfapqfwB
V3+yLDsj7x7X18J/JnV4r41rtRgEHoVy10mKS2lDiJteKGkMbdEAtdyhc6Ta1UX7
yHOrjZqMvRy6owSufLSqGE8F4JICvFkAltdkj072Q27e18JphNqNsWO5vAdP2SRJ
t07/ri/JrPd96rljM+oCN/q/rdTxtZZuE6LZZI1keq9GqyZ9R+Lsy9DTtFX/M/vF
gEh3fRqA2Bq27Sb34EqlaUCIr4U317t045X8uqC0UJWrIFYQx5Qgz3MErd0s8kuD
uWnOalF0zLuDc8sv1/juHKrJWVgQCb/YZv6x1c37P8XZezTc0CZkNURjh7G4GbQ1
De4BZSUeHGZOkD3u+M3VZIva3F1NSGAx6hvIXhBHab2iz7yHYxoiwy1zpS3ESTQ0
l7pMsRGVY/Nay5oGOP7e+E3QLhUnOJIPCLE1Y04pQQJBKxwZoD6+T6VHME+6fo2X
JAD0wokvJIZimKOH6CDRntThDR+1hGhWuKKVWMf6n5vJ4fwruVuQrHAn5lexVXF1
dBZDcEbo5cBYrjrGWVT94mR5zpKX9E8KgcouGil2EZiKtSsjN5VPctz+YWIWJXSF
2Te2Yp8+cyr4W5fJGFLcYlHu+CrJMVv56a6TKKUMI4ZZMzc5vnk2HFXO7fWqeBtD
3ExFHDzJqmpn2HGe4gV9z63xmtg6Z9kLnWLNc4mMW48cBn3H82TWLFfv+5EQPDUu
Pvb43anUokx36aohPs4fjhn3Zc8l0Ve93afydXf/0jjorL53y48GD+uQkLs2yQGF
gT0tVPwoWHRoDomWsMbfxEWzeLfWoX9qAfqPIx2QHLP7FSQsGdymzIZ7uklZ8qT8
8zkcYBsCQIMeoJR3j977YR5asJn0q0N8Qo60dA9bcHw5/yJalO55QYJhUwBY08Xc
swnWz7BA9lev3uE6krum4ANAU4k1Ml6ouIuzQDA4Txovj2b+NsqX31DdwN45fXIV
qVd6Owly03W9uAqihTtzTx0+zMpjFzgYq3NAW5XWwFr1uzVO4lMj+wXcDpnBOl6L
cCIYMIr+nBMn9dUv2X5OnUsIXYrf7g37FmYJDfExEOK1BkKHKqPgRjbCne8s5q7A
yTnrgPO8OqI24a1ejX0mQZjphGE77csO1O17fAs39VYDZwUfsnHTzTN4BBq5XwJU
h1APXNOMqRbEM9W8E7Sn6Y5HBviszcb/43FyvKn28Ty0w5fSoX9XkV7q6We2S3Uo
hfNAsBX5nVjj4kFnV+yXX5hO6A3P90540yovPo8FquAduzRJOnXh4EPNKum5k2al
5DSdX1lwtoPVBVTgJjUt+uCA0dPXxHcD61CO8lJfyQoH3OvbGVwXUHFcQPvD9gfl
do6ay3SgYCtzwsEDS3EMrs/CXoDnrpKjtclClXFautMFn5ZELqeiEPpLHwkFknZ+
LgJUClYIXSyxWJb2HCMnm7ADQsB/4LtDMDlNG8vkhK3D792lZuP2Yx0EAbWWk0KY
wAEoxft8nkkH22vMcVpok5i6GZgap2jdZVbJzCm492ItLkm43DQ0b7oFx0CYwaQ9
XkoYB+S2FjlS/FIAxbsbkyiT2J0RrfRpdqWC64E3j2MBqTAWcRNhlk+BoDArFbYm
b1XBF/BjSnmX3zn/4LEu7/gTiX5IBIquxYk5ru2zGfBZZe/5ESPcVH7jc0Uvrz0m
nP4MnA4CoEkMGPgLKc6YH6iRQ1CsVfL6sVpoG02nN+C4R4zoyV9M3/K546YXvCn1
lWeDG/pXaiUQ+bBnNfc72ujScokBRg1gnHdn2ebPEVm+T0axf3s0eorY8qYrt5+7
2xrOOtJhUu5zy1yz/PTxlVtKaGeQ13h8WGTLZJFb/ylC7OaN0bJ97UPoqrFhZdPk
2beSsWT3zgYKYn5tQ68hDvZbmbCd1shFKU9kM48HwGcuEG0B3Z/wsEkhTzR5Q5nU
Le03YsK2pK48CnVMLS5m3iT9L8RLF46c8O0aKT7a6et+L1GQeYSdwOuSJK9hAJRy
rx5+UxPmOeUSvRfUxo2SVrXMtRMA9nRCre2vn2wd2bBZdzm8lALCofKsVW4SWqv1
SHeqrrECRbXNjEyr694y4zxQanFlGRRC00dL5rgTuOOlirJuxVurl2XTnRP2OJlP
FEF8kEOMtTA226gtT4UGWuVzf+QS4GCcHcxcLm2hM5MwYxlzpjmKhJqcl7dj91gO
4aDcWmKtAROzsUuK8cIfG5QA2g2+H0KOB20jjTJKn+5k3cPsY5aNBr/kZDEybVLh
miihaXmN2yUWrk1vd+13ybs68qtsPBwZB7z5df4/XtX0hrkPMr7FyaPr9NhOPOTV
4nl2tIa0u6uUM9veW1kC3g02g4inWeXdxx2o5KNjx+cxRmZhl9EvG6D1AkxnytOC
Bbu+JnL7NHash7c2TMzA8skj9Nh4FOoZT/AvnJyssCYqa1/qAP3fhnKbScxL/VAm
Ch6l/LIE36xlH2Sdh1M01Ez4w0W2ZKiLkcugG6kwxi4ka4wUkimSj7VQjFH32fOI
aCSNTv+6CFpqejwfaVlYUooIMsmZsp0fsFf0XB0SsEh8vg0nmE7WiRrApBC5ceaS
4fNQE30hiV5ll4bkIMvqNv2c0woIzVJ+3cS3jscnPA6IjQ0BvQpNxWVLMqB0Kbsw
hl+Y6BgAaBXy0syFH2GqIerJ6nHZZOUf9inNFQNmps/CsOzBZrcXjgf+faTxkHoZ
q/D90kafQN6VM/EXB3rbOuXIWDeDMn5RFpAnYH5mESfTiH/vID3a5Uasgg4ineER
8BVC/K04wMoZbpp6NQvjrjYeEEnFP7VZ7iA+WkQ9YPDrqXJ2DupYg9OYKQyAZh+j
l5ht/ISjZRoujode/56699NAYx9+iNbrXVAuTY+2IOjWHsyZUfK0P4+gQM9vhXwa
4JHFu/JtJoDa2A0BqFPXRrlIAT7Vz0YZIr2OQKx/sP1H1fUKm2LEMrZWh1PpngJi
ebBWiwaXEqXUl0YA53I85xJlOepZJmLh3xRIvC3zai28z+SLRAiiJic+unIrf0np
vz12lOBMqlocdOafMSuI1rIhjMCfwybSkVdOW3PNrXpbSj6t6mvGxUnCinv+S8t6
4EXH6DqN6dOMwpEHVw5h7zdO/q1MZFQu57k2PfgTIXF19cJ8Pi+ckWxQ5q4FQfiC
/KcxnxmDZixVjbREl+NkCJG900b5gb1dllVeVZIFIn5pDwzKzxdDyQZUJxmdjPh/
zvGnOndKHu6s0BZqCENkCCqrAJoT9vHe7HEMEvDlda/+cKB0pYWHLPiFSullu38H
cEyxDEivucxV1Lf+Z8XyliXICfOl1x8QkDGYdsehvgVGmbfROnz5juWk8muTe7tr
ep/rTGcBRRJRCqaoI/lc0lFQ2y1fjhbclfq/WSqfTiOM5bJi2NUW4FlY5TxFWu+1
otzSPd5eGlyDqLwlA2+l/ykIVckgZ/eS1J2T+5ZxCng3CUvSTVWUneIPLuA2Vk69
5bR8yzNMShJPrXgELemtcn2R25LWtNyDb/rzDbtGmg8psGCjvlhb1BDymG1mjse8
jSFut/zPLZMzeXfQp+9YLcrjxGz5MOiSzibX3YHRbQYIHtfyz5/utNQarvT1MIOZ
qAZ9lPn4x50nSEBFR/f9tuDoEg01VzI8yFKhiTOMoIOaaNLa7MZ/lTp/fBYdd1Ds
9QGvGmU2RXhlwnALRpL+4tIQN0CgPtIQ6SCoqcku+0cIgawk2ceR5WbAvuY6DRJZ
hN5z1bI4+TZqzw83Osl9v8qcISgXoW1pLdcN54DUssAA30st2wKxrRNalbFfP3sw
MZeVySCZNfkU8MjPGv+xHrK4mKzHMeb09SC4sqC+kOcO9rQj2rA28U/+TGtfdQV6
ZDK3sbP5f3if4EQC4CRRwloMVTY26/c3XukCf3WnGgHZ4+DNOYBJKWnL0E/ZrK85
MiDf5eQEWzojDbwFw90Tz4XhfCNRAled5EVD6/R8YnkfBAbiD0j5XzZhCsGmoo7J
SeZAKMYxokjQgyszWYjoYDhp8Kra1wlNXLBwZPuePgJLChtSNxlndDRsUw+/2fj2
CBkTAOfvwkX/IAt4nItAd6IEZ0EAsbd56/Afz+RQ7dRE3PfeX7qL7fS+gnHwQW5n
Ff+ebHJlAEPDbuCwS2Ih3p2V2DQExmLqt9prFvVH4w+/+AlOkq8MVJ7FIvB9ENtk
kh0xWEgdSxPrcAuMAxSZmMdIcTmCljh8vooljOD9u4B7BFYl2tR8OqGC4MnvwgGb
aQfCRDHtfEs1doKY/31vXhIaILzatVLRBcuVAgOp80Wi1h1arROKLwWpDoq7JZIS
GrmRG2MNGkuRATAy4EzEUX4kKyiWaI/KAQtzzRFjR5Rhwd3EHKIveRRaTdIwNdEK
n5FpGrsmSRTnHokLi+QvAGxc9/BgUzuYWioQct3/eFrOBjnvZuDCOuBObQQ1OAAn
nyE1Yjg7xhbanne1wwPMQI25Tl5T0K2lV1VaqXM6VwK4q1XHcN1m7O3Js6jKI710
raMDyOjy9SuAmwGp4kYTBFhq94o2meaNQNoKxMMnBzPktJ08FddsEQ2rEcYvUP14
lM3i2NSVg9+toOzZ76VQaAkRd9WNytZlbKUyTCiV6n8Pa5ahMR/DqDJNT/OGWsoj
g2uQBvkY/IaeYrs9VummMbRSBKPuhXBY8cMUxlhxAXLf7DfxdqhYxrf9BMWLnPtp
1gZ5q4TiReA5HFQYkvCazkwnt0GlHNrhq7EBTCF9KgQ16428FVtbJLMf3/2Y6ybc
kaVJKFhRaRSTpUGLPhg5dab/ZPL0FXHjKqtQXxASDcnO/DVNnklu3S47RVE8V4ue
BzcE4v+J7UE82PsLP1MqEsz+ZyzVaWgNPylgOHbqRK2+rNOwdN9pLJXgj1/ZjjTR
EOwkCuF/AbWJvwGEg5pR81JbxqEfWWs+9kypKe0tOF70CeYkoN9q7TBkgsHADj7h
egL1iHIODnxADzxo726mbEqFMfpSn5t18FJTOmAwA/nuGDzo3+8N1Gv6z+r8vrg9
Qpi8b0F192ZWtIL/0rR/t1l7+pdyEgjru31LkbUMcWQVV1h5QwwvMwvuhGwaa40B
klXB3qqQtJYuKLPE5LpLdfLTVQqD7vJbbSOzFeujMR5TP/CWX/pL6M9FFPFaC8RN
oG76Wb1y6o3A8aVbUYi6yJeYMDWizgGEVHyXd3knZEdnF7xVHs9TQgKxCRTPvhrP
651sB/NrtVL4eMNdzNFi7jnlNFeSOa/GB0gdTW3xkKs0jdy+iS299vlUewBIRsmb
0XRlnrg3e9A01y+R6Cpc+4TIEogL/TDwmb2j05N7P9Zal50uqTAJL5PxweWbLKO8
/W9kSPm95zL+sKIOwScDhyMDV2B6UHrxzpn6vOCxBXcNkGzJszegBUfV+ctNtLzi
v15c8yp96hFX/AYH6xDjCPsITQorl2IpL2piOn+cS8NHvxRr0THZYcDPitIDdFun
Lr9L8LKxKxa4PNEITzB8Bg4DbojQzhYtN01g+2JaUGNZjx3HH2yMmuF2S8rZHm41
6iCRoZrGlcs8M3nw4k7vj+pqx9Z12uhXuwwX7sS5A3axOazmFgYo1+IPIGMueV6P
ILg5gIN6h65m+RBhon8RwrNhYcydx5ikvW/TCc+21Q9nTX7mB2vBqS8dZiMkgPW/
Ptm00YmMxcKTtMdncqfa0Ipil/Vpt06tgMI2Z1PRadEfNFwOPqizhJxUdBXyk7rc
YpPeoWdr+7Z4xfsRY1g8ZJ7XYGsweDmzN3eKzuHxqoeR3Td/D2e5SzY7yErc3nzE
MgpKhaan89xcH75UovNshJGiGVjKFpQivGsit2hMsMHgjdZ+jO3UTFMKFFlcqdYh
Sbs17/BUt7OeOzeth+i6abaqRv02Dq59EziNBlHDiB7I19Rtf8YeCQjzZ641ipvD
9O5SM8upHQr8M96vDlyR2aRgWg5b/Su2OEFDIsV22vjD5PN7HJCeYVg6OeQrEv6w
8RaN3T2KTnjjH2rlptZaada2gIQClmok7MN4PQuLbSawrrRT6ywriZFL+DtqEjKm
D1n2s0OFQkIrFXV5CqeL0rx2xf4a1dqAgjXT3Pw7A6EflGqHvtWIqaDOzUGDTxRt
H8CWwB2ApYQ5lFJ5M4txymJH+fmDcXLykeIrBzNS0hx40DLTqZbYXhU6mzGYRuRC
+PjGIGy66P9PpYj272DD4pMgI1Sz4ra+YoRzglK3TtU40RDexWNqd8adkM7r8xzZ
fxeiHMGI6aSY1/pLrZ5s5FtdxttZNtZulq08wVcvFegHcCDbkx7eAJUEhCY8iEg3
FRFTscl+ifzKm/VoigrB9fYJ/pZyc3NlBFiq2a2nPcU+rLIKYDN5rKbH68JLqc1f
1qeiBVpabGt3XMXl79wXZ1Nyn5gE0xhJCso/C899F5oj9xP+cHU46F+SY2v9m8Mt
KCrqk3n4ac5v8QiK2AQ0ReqmQjDwuP6mqwoTvyvmlr8g7q5999jfVnzSywde7kqN
ROX4M64aaLkuOkcCHW6yzmLhB4lEB2dclRLwTx96t9dPmOiDHP66LykasMWBQ625
HQiBcDFNiZMOXBxHyHT1Ghpm/yvwh/G+efWIyDxCw2WIYxvc+wXYwqKxZyKBUAID
kvLGvbstjJ8YiirAdbsrPQOZ1szq8QNoNpysTAy2c4kqAPr8wH8Sbb2xiYtcBkpO
MvQ3ALihyb9Q5JmnIPNrfsvcpwFtv2Io+IUTYFMF+4hrCS1NfEz1Ekz57/l3rpfU
1oo94TjQd28njkWXDJGzSK1gFUFxGk/7L5OYJt82eE+3LM6IxQa7ybqYmXOBHzSN
h9rl84paNvBNMjbYAzVqlNLMNttSUE8lZ8T7c+52on+qefATfq+e7BVoMfIGqaCO
1zQMBxdqQCrZo6zjBUwsw2YJIaTWK4v1qoRtr8DrxbqmVSrtDQ7QLBInf+sb3ArQ
gOf8WMNJVWNCDTWVi//lvoJ+hj5ONDHvJUIcr6rfdQvCorGEK9N69yPvCpaU8VH7
1wVYWrfkjA5QRq/QQvhrUlOwcIRvcv976HvLZOQnnCUcNv0JlpSj5V61DEQCWKfu
Wf41kHsFKKXpFt4RKogXen/whLsM93TEMOt7rCHcxcWgG5b2UZVcTV+yvHhGkoOE
2W34ydYehA+UYmH2z4qy1DPGWM5NzbFUD027Ixh/yq0M/IzXcNXjE4SM8g1TyZAL
1C8IOi9G8n0E9ij5YW0py2J6ouKsE3zBS/Vzkl9ZutH0CswtAEPeQB4uswyxeBA5
oRgUCzxWPwU3+8Cg6sodgt4xMttpqEPHDQSxW+O/tla9eHixnWSuT7cti+G3u2OC
nq35ug5OjPlMKdUjzAkxydh25hWQcezpr0eJ9fKAujKoCwfG9+49uscetqNHJsNV
Vqszac2DQHvjBCyWfElifwFCE2sk/4bk2IhnKuSBCeXIfmrvpkJf7xPv0TPv/OxG
hAmqVjJiXU3Kw3i4p2H+HoQujwWo2jMMsLvnUVOXgrknjraZ9+SFM2or9pI3D1lf
FbAhuzjjUcZuYoPfRFTWYImfjJ36uzay0+RBp/arLe2H24+zRwrCyNrMSVIqt5PQ
A2fFDhzfkjGB7PuLwF9QEy7WOKi8u5oc3dFGeU+08pgbjkbq7XA5OLt/RB53FDFK
GjRQ9l4VYqD2he+qBtLxrHOiftDqqo2elEEmstSVi0+RgBMzqpBHQ8nV4xMOSU8y
4T6Y4zKQXB3TWMJ4tnCrpdo6qV8GNMwMl1eQRM50WzxjQzHSj5ioor4+Egh2AEAC
aEdrfMecqFCZXFovY1qJ+4WGyqayhuHkfpIQMfoKs/Az1KKkPxGsG42/oje+4jwQ
InxtftfLHdpsFQ8glB3cLThlKlGwknaMRJSI/IPSKaCbVWkq3wloGarWDNO8w+3D
s/MdjvvLhLN3C0P6sZBuzD5ptM6WX6j8h8B1CV+uMY5bk4AiLYsEOlpFFPLZpGhI
+yer/0dlJq3Uo1Ljaqecr3iwGRoe8NvQJefFB1laEBuZQpIyT9urjn2JrRvA/K68
yOabdAx2mgiJ1Y9uYIhR3soqdkihoCJWQIKKYLixYPBdwD832Y9WYkgO5hoOhtne
lTCjYPNZYjljAECMHyLr4/Erge2WtVtR8ZFPRn+uz4u6qAtuqI8flM9RQT1jKobg
OZr4sVgLMaFDQnsM0v7OUG05cQkxymzWhtYLS9em/MaHyof3t5A6la+lE6FzzVu+
solRd8+Q1s/TehsVckHznVALHqomyBMT5zTYXyoeulg/hqAJZTX6cm9Bmm7XR24y
Vl0p9mi4e/ERxOsxwEHAcFEmx5xIMeV7bJ1R81Iq8Duzih0Nm7s2U3YHnyViN5cV
rCFeLO+YNOfFBdjLXAMRQ/y92ShGJ4+es2USaoxJNBFZuVzdeAogNgt4J/L2Ii4g
u59iHrM25bQ+vTrEknJ3r6I7f7RfsrstBerW99lVaW6V1ZKlElBa5r9kMHNIOi9o
Zl5CySS/DAQJUDN/5jEDdo7/aaZDRnN7nBxWB4kVn+TbadlaQ3djXTIMExslZZuh
/HXGoEY9autPAeEewSXhPpdpe7E+ghuSjr2fxzvvsciL38HoLp0BWNsfwNzMCnPc
oL6hL4q5kMlHLLnDVCXZgk8PLJBdXuDm6vZf0JqEKp8+sUcmn5RRWiv0kYvF0B3Q
53I8janRWqg+GN6bkX8l+bjsV2cKaAKXiMkwNWw2G8rpMGlrMKCxbSwgbfosRMgg
78CZXCzvnCuGNDu6mDgXDS5p+MrrGVDEPSiD/NKIXfQgR9fMDpUUhRzgqYC2bbcB
8sNz9YDcUQTbpetzbytoejG9RljO/5+Yu1+Fzwn9A2E7AwaTsbPPMHnMr0aGe3+2
fpd3dpKuGRDc22qB1C856xjUamj1Zmmmn2IOPoAXx1gH5UxJ69YVLd1oQOU7vr7P
H8DWPiW+cC+RMbmRlGHNpvPO5t3RRVQEe0j0HG/GqhaEnnTj5rA87E7UCDft5KFi
DJMu1e2nOCpnXfibwQLJCMW4nodoq9zYeMpGa7p47KL0byZac8yHABSRQkU+QCcs
CPEMp6EnIINQtX6WCR7nKyE18LsDeCWdr/Z3TMP8lhz3lr3XNO0SHtZw83pNV+tP
psF4I010/dXXcJtVTLllb3m+vfL8tzUesknYa0hDjifuZ6VWd0KdkOb7aigbLZY1
p84fz8kpOsnh5WTMXb0ispEjiLKFoy8nDkzhJOl88q53zkeDJtq1zyWV3WlOOvEM
OnXz27A/+Jb8p2+YTwl+rnF8IDcq/JrSQCRVOMzrN+kkZSMsr8CqsdN4+r8k0fsh
zT4ep9KMl2qrL+Jybp7300Cy1b3XZkpQVx/0VJuqmboaUamAe3mEw6785+ATstam
DPK+wk2oOBsZ/ST5/mTXIqEQMZDFCjkJs8pTt+x8Ah4rt8loUlLhgffMferMqZPl
Hh9dPRRcm4EoQqO21Q9uxYoulMkahXPOae4DozdsjoET4yhA91CniXeDrw654yq6
eGkFg4Yqv91p+W7jpUyj9bD+67UpouuCQAuejSKt36xjsjgsyjYuxP3pCwHr7RIM
feFRilymEyzmXcXm5oitzEeKfCDwbJuC+iujyjFJFhhTQxWtbZ5XkZaVanum3Pby
hXCiOtJjcktpjLshyLye3b1IndWVT/C66bBSBxL3e05AvSoU32ValbIRrNhmSwKS
JqaqXJleOMK1tUG9JgQjvDNR5lLX6i2Dw2oAXbB4eK5BTMC1JmAHxUxQZgdYM9h1
4nwD7gmJjCkdJBp4lCJgR3FwrKI4wO2gQ5xHjF4CsJD8XnxEeHJ5PD/jAJp8p9dK
KTN36Ifzdq+Vp5HOLVNZcE8xF1PcfBiFIcu/o9rIHA06T1wM+JlRh9bPjfW5+lFx
IxsD9NEQBxcRHtmtVHl17uMhajHsm9RwgJmtOJhy7lx+REjIsFdc+iYO490da5L1
ryuboz3vT+/RMGsITeMEBP5ISOCLK6wBjROQlWteTlszeVKKF3JGv8qdcRXUHRbW
uBtqMmBXgTuiZXnHkiVV6SSa6G5LVxOJB1pA4xzNNxbp09Guk48YFfHKn3O3RbV1
lKtncdrFBhfZPVXisiAlt/Az/dFcuQ+LE8K/YVOZfHTW60POMJdgDJ97IxF6GPVB
F/1gnPKfm7CHK8JPUMW01Yyw3tAIqOW4BMx+cl2C62tEY8f9aueJGJauhnjNyFyV
AKTxVKwazuyawjcPC9z9nmFrpNNydx3Lp/6XHM5KU591/ELmT07CjWk5jBSi/nsw
KUZrQCflcCW4K/hRSCvyfBENyV3wlDKRhCUP9WWd5QfBVKXAc6BrQJK0gJK2tQI0
ev5+F/dFS59RBHiZmoLDqtZ7fA+SbbP57+Qjl9kwTfyhoaro0bLID5Z0wUYm4Gy+
A7MrwgPPF276lfeQybzYT/UrTlTxp1JyMuwIL5d1uBhABJcawm33i+4I6vH+9stS
PaCB3GU1gnbUpnQ2xlemZbZ9Y9iXNwam8Xqhf/PDIik88AqnKzQKz0kWeVtiWtT+
igF/YRNnt21+PcUb/GRBmXCVBR35OF7J8kS8L9Gd0NWrXTTpuHe8BrgQeWmHSuHo
Xacv4ykMm7L3Cb2wb+yXfnVkVKqf4/M/7VHJ+i6q55Kms1W6M9mtNbdJPzta0xOO
oZgwsnRlVFlB6zOKGJRXs62+UWv/m9U97M2i5i5/hHd+zt1Ov1mPlaRzbc0qujyf
MxeeUCUiRdYsIc59ViOdifYMcA83HpT2z/bPiOo3TEXiAd3bygWn+pjSuCFYeEyA
IaXAPLTDp/WrKR849lx+E7lZlvn+rI8O5/XM1q5MxDC2VSOPYUXBxMFLpyED/9vT
oS9xHSqefISMtIXO6ryS4UKAH5ct0eqYxBSNLUgZbVCcmssFNfhxHVNbtGadpI0U
krcODCU6zcfdC2JJ/Vz7Gcw1s1dP3V1oZJRFvpq72okGM493kSKtGirR3G5pvogR
uAbjgn+9Yazt4E0ITasCFDeXMJCMPm+jpPqY/evuGHmEIjLotQFrsypYGjfPM3ME
pHyli4TQdPz8483E3h8eysHKWLhxMkJBcgM2bzPABITt3Cv86aRiTyugA3QajgYe
Lgbtkq13aHe0PsxqpsxhSLq8B/RvRPpkL2xSB91CwLXA4jhR8BuOXu0t17chWD3c
/d6Fl3LtxC+ctHUIk+xzR6/PrGO4qrqiuekgNB9BHyl2qlVTfO7hdG7LztNO/kxm
v0mLun194Qyxzzw8ZwFZU7YvNkF8SuqHayb/vPqcwXMhkXqY+tGkCvF4Xmb3fwmH
ePBtH9iRdK8qDMz8Q153Mgygsjp7e2zEOc8ILqXAoR0X+YZpN7efG+Olz1am9kyN
DqLiwO2C4f2dn+fEZDHfjvZFc1yL35IhE1OAGc4LRPuRSlavh8exAETeyq6GRJFt
Kt5BM4jfjeINr6KtQiQqgk4QmpOrAqFyAkz/exdwPDsfY/wqPXnkvgjthbeYuM7d
7Suut+izuM+fyvZoMVGAbQDPlr4Hkt87bWTiUqTogTyHWS8GnMhYUgU1bMzMP6tY
U9E3z3jPcT1tS1YiFrSLZZOQT+odr91LyzMghSN64j1lBkAW7Ul9n3kXQs86xH35
vqXfiiLwe3L//6MXSIoX+Vqr1nG5fqUQDOJ4mirmH2ywjjFSDO5I/ttDwYSBbv9O
08jWSfVEdEUUWrsIUkXs4KT/MWyrZIlN76VPliCWh8nUu5S48fl4a7O9hsnTmC/N
xyt6Fc62airHnNSTCKARhZgTGuI9oDBQZk1hsLJ7C9vGMODy96DZ6pS2wF7USFt6
czEsctTk6w3zCnwrz6DhZlsi1szJap72m+1lUCHJG8iB83GFqQkPLeVnok+KDtb0
BDqViEbY9+Nul4VEqr+GZoOfIPbv8fH59qLaQqGsvitLKrV5eWpGufZkm/ukEB5v
BFp1Y8Ka5j4vFhCsnZ4c8iFykU6pICCWH1ahKxCCLPoKbkZ6kusoFNbWbfv1mhsV
YnOlFeluDW+T4JR9Kee3jzY45n+4MMKTiM/svp2Rvdj60tnWh2KE2rBU5xBAxUBY
Vr6xLLd3qtU6TrhGNN+y1wP0ESFJcdXTEH6FhKkmeB3ooyz8EumioArZdEKTm73C
YczhXyX6J4TwLOktCRWgRtQR+9+1Kiio3f6okylPA/vAIWga/LCDikM7+C+slJbE
haRyFxVsAShnrRROeXBoYLLSfBRHLUs04Mq7EStPbsDHzqTtdCQZKsLYaJV9lk6k
pCQ8pAT555TzZpKyPeIZKmARk2ykYaC3RZ4/MSxgGoZlvpxqCKcKiJxarTtVTOdL
8iqB5Nph85FqIH04fQfPWFdXPIt1hW4O1GZ2y8CqGgwZ7WMVDAd580VamC9OzwwY
SGCCP/rcrgTPIs7H01cTiYY7y45Yx+38kNv3fIw3/ofFCOsWYheNdnyinj4XYjT/
eMFT5Pml0rBeYrDIbHeVyVzPx0tQkCQyLVPYkKDN1j9HdvwZkO8yYBtfLBtfyQnv
l+rQ6bJcbZ6fI/Fkig1UrnTiT2NuMFTwiWTS/I5Lh4Voc85zWemIbuxTvlhNGPV8
BODpAMFdQL7Cs1XKowmGa3rVfjnCitc3cuu0hhwiMhGpuQ+MfCXX0U4RYv7K0CH+
7vqdKDEbcd+AMYLjfPDclcQn82E6YM1y/t0MXSb/XRZNqtkJ4eSz9NcJFjc4u03Z
FniPokSmvu76cRoIPyGWyYlqOJ4jfmN8wTTAlpAUKMBqeGpMgTwJFYhHzsiuGCBl
jWJ/Z80VJ4TuuQxYt4TKl42+cO/sGbZRb+j34RIQRMNuYquWi0t0BqkiLzfg8Arw
Ap+Bf3KpRbSX2fGAfYPfnf6A4oeyDh3nVZfWIALOJ2YHPker7cwA8ZCHhpBJce3I
WhferCFZ4kdnzqnaTTgZ+c7sFkZWvaJznjJY0jfUpbXvvpXW+fxXi6Wor/6Rzs9u
1vW+aGR63jB7XkosiV1LP7a4zCpdVjOEqcmHGECMHIPrqF784b8WuuNNsgNf9Bdm
3IhiM3urWxCJ8mLt+DNfv1davd1fuBIbLGdKVE4cQ+LGltMioJ7L0FuL4pGA8/Bz
f8sgRz1iLtt/xkcPq/cPQeqlW6UMkgqOsCm5P69sfo0LczDRyx8jXNbmOKF1gzQY
gzj0bInaX49JEPN1/msV3/46i0yOP9psywlNY4/iHZmHLrZ7qd6ubvLME6MaBc45
XFW9QUzBGGMpn8A6cwHMZDYvwBzJLWCg3emFE/A3lfw7IYI1olaNNaYljAPSISC6
LawE7EW35y4HMqbPwZ+bpv3uWTRE6JROY7vZnlV4YHCG6g6rPYtJ2VBauuhEQTGY
BRNyV0gB7AX7iMd+xV9lJ18uHB65yfIZYwDQ/UJ1t9eHclpnffNEjQps/7nrVbZl
TOk8V+M4Yii6TwCgvHuRLZnshE/vvKq3l9D6OOzPDrgyBhQUUcFEEBTJzWZylsx5
zofzluin/urVtzIwYIPz00glVv8YV4gNiKEmkmThMC6aMAm8Btg42wfMhi5+KWEo
z2ClU4qV+LGh9wR7rJUvOAveErxFzgXtDPJxzkNiMTs4Mif/Pt/z/Fb1rXC1WAv0
tOxqTCzbzxvbpiIQAcXKp4Nx7tFakDuwUn8x85+fydQyu7bfN2rXpGkqe4gsTqjI
LwboDIW8CmvgfFR31SYQeYcEnkoSjz49lQ/ivXAhM+XQobkTca7YKLOFuDctgGc0
VlpGMH+wHxi4y+pANuV+9mJy/4Zt+SZherF1mNXLLIPmgDnfzmufZqOgFyhVbEPh
xPF4H/tPFMtINlCmqnMJEUCVleY3drHdD9lwzePwIP2CDKxReB7ocePrO5N7tGdy
bwy4WhClUI1u9PyhzkLUYmdGAINYxxV/fXrfogicoHdk0yTYDg2jrALTRREqIUqS
rGbTKJEpmrYQ0coOqcxw1cxTN4NZoZHX78tt2JzbyNnUmrS6gNTYvamhLmBZoigI
+cyx4citaS6xC+rmsaGlFv/86SX4bPt/YISOxwYVv9yPVfoWr0MGSx1gGdDAXdTz
BtXdJMerLhYIyXdY+LprhfCsCyoFCAfDeieWSqRXKTqUqz6O0WikjeJ3IU8Ybd+e
MGveWgw9NJeMP7Lxci6XBDPUwwAjhYU+81bNNYi6n+BuKYkW47cs9w0ivf2WVop2
/6rQ5xoiHgU8huSGklbfs1w4OKQo9WgrnAL1wY6UjMJe4SnLBLa0BRiNzp9Kz7iw
Sv5KQDqTt0ljaJboazfd4aTduTcV52puguVyexVbAtvW/t0mS+RfujVmlfBMDsNd
aKFxVoWqZKJMZ9rm1aPDVPUkwnZG2GX5vfBzD2EN7IQLog3lZyA6lI9352cDS56t
cVdCuQcyUv1YFNmY+KRoq7KcuprbABII5vERMRSTy9WJ3ghITF6ficzBkBzCdwKV
ITLwHkhcBWzhKlE0SVwlMIZaUxCgfL91mRBI4jB9BwUejm1yGFlD3EQtyF9rRNSH
0TvtHQvrhEho85tFWXupXbszD0D4JY7ZrRcUNhYpBDuwMFUZKUSDxKhVrpwsaUt1
Pu5t4MwwldNV+QE1Qb43RYhOVin2FWAGGkmorhkddFh3LdNUFRj31xa93qtEg3mi
dYra6YFT3HNhfui9OeiVKI2GwyJzf6PZtYcMVjmKAvCBw3SqRbZl41W8Ha1Y1LCA
rNaEYrdaTILdKsvmqaucFun1/IwmF8NuibhMIFLdGITHZ+dBqlxWxpaq0hyMCZmc
DRAjDyKb4nlIbs1FUCvql3YnY6ip2ksWklu2VYsP3CpuFxOODT1LTxgumjflxN/p
Sz2i+OnMNWGDbJ9HhQ6y1erR/VlwTBUMtrV2+ocA4vkwpR8F+ahKuB7rZEAxVbwt
z1ySwt+nMjLDW7dzNNJoIRae98bcv2wMEIMF6keYjzQkObePKCle8j+4huwg7iWG
UgSfXTvtTkPbRKtJCNioHnVcKXmj40E4ELqbc7ACdyTIMbhqKti0hhA5Al3T8Tes
J3M3IWM9JdkL6EsCYrFwnvupEBvW/HL4qFb19kkFC/EUuC7FmsuTvWu+73iDI0i7
F/jSN70poX5BEmh28RTNJ1dMNmKYwwpeyqQLWoTyLvAaiA+5PnjNQL6qrXepqgQu
s+QwC8Ien8myPSW2H8b20CwV56eUgxNcIawns1PFvOkwIRB1UrOTDBw+wx3zO12p
ecjpxhKnKHMMLqyfZxylAyu7brnkqc5kTdaWSGIZxsKhROaocd9g8mf8Y1rpTx3M
34IqeoDt4TugprcDq8usvfNcaKWwURUPRXlNNU7xn4xokpKeJS85DDQd24WCCKzg
fFYWnHgW0g+dxZUDtUdii2O1I6nVnc+6cVvyWdr5EA+xSzNbcL+9+cbFXb/nI+Sj
5LWX8YqE2NcMMwfl82h/Bx59yW/O18YAXD+KxIsVg29EW8vwkIK2WVkcy+8CCKqA
R0D2Tw9jLpSbkxIlWp8ly6FOpyIkdVZdqFNqybHYLT5KObG/N+/nRI/vj61gDBD3
ZyVHLFrEwmW7ndcXgTk7Y4VwWPmJ6MqcrYYpD52TjXN4kq+3ifvkFVfrKh5GfJWe
DaKu+9Q9pwgBusA+bx0lYPF55TmAGRRRzVA4CQ0FEEawpdPnL7z31Cj0bfqwKEKH
pR2aGjX3JPR5W45NKKgrVTjc6ceDYSoXruQM/MeXfSiuJjlwFFiLkjHMU3mtomIJ
P3l83Gu0PWroYKRDZV4j4yMLy7ainqcD8jAfLlUDv5gH8xRHx0jdGchph+kU2wfv
vsJvPRQJAr+WgWvFrW3TIIELg9wQD8wyuhjwrIMdUOY2RwQAJPjLac4X8HsOwsc2
/d/7tsMYWtJkbcXozXxzDhhSUN0LaMEP7oMLQiuBZKe4Bzpc5YN5syfgsUNOM/M0
T8YQXjWSkRUS1IOg8ugCfAdStdAsek+2oWn0G6hdnV1gV2ld3SDh3oFONszlx0AX
LM347s/euLV3huUia+BZG1Tq1uO7XS1NSYM0cHBPvAgA4UIPnKYn+UUqcu8iMTtV
OfHrspikE3lTyE52UdzeFRihqD/cokAHZXmb+AWk3s+BBVK1oJ4NwRIs7Kleou9m
INSnoYUXOSptxQZ0t8DnDDtpO4FTkOmnemBPW47ni4f6EJ2Qni+Fh/K7f7G74Vnc
KW6Bsavdx5l3/nB1OeezP0FpwsuZLs1mirSc+mIkYofPlVBDV1WNl2VVf3DTVVky
4j2T4tyaXXlPlh0fDwPHMrp0ZgimOAHK1FenIjRIYTngVEdayZb4T++P17kJrXfB
t/w6VqMuOsL5z7PLcIFWYME8zL+z8d3qLsrwc3iBj4ngxMfakEm6tT55U1Hu+sui
AWhYFulWfznnPQkNpXBZLwV3YFAF39uwFue7Bt9wgoGbqTARDS347f1JtrU0V4N+
tRkcoozCt2K8ZV6K9wLJyK35K+ur3SIThvd7G2+vaHxoW9kqzBw6Ks4QfDkUzDqs
QKv76ESR0OJVphMsNS+X5AYZAk9Wn+h+TUoFtskbGNrX1SaAAeVg2MHMpUhP3huT
ZV8PyaqJbsSd0/uEGcj8e1OkLZDdlQf7yK6aMtScLors2G/i700wct3H0GYWQkH9
9TqULaehe7LKVPGzDvf2JPW0A9IMLJZz/UD1RI4rue6UlUxNfLjUrBTMsutH6ybJ
zrJ7GpvOu9AWfdc9i0MQMydgRZWsW9lietZ6nOZLogUJ5KhrN9OPHY3A6AJccQtE
syVhv8q+foDn4HwdLvHFEIN29fTVywryajNuyBIpHY/yzsczsQ+AtkoweFs3HpHS
TuqtB9e3O6n1WsD8xbz2GtPEVPpIm+kow+usvFuQwxaTeLZftYdqBiIM/Fkxa8SO
Q4fIKtnReaYMddRmA0vxk+FDUXNacxLAO0nvjSlmjOFGRBQAwytf56X6OfYCb41N
FvJGOe5BHgj9aZKr2s/6494LR+2JQHB8HBlOH+TtAUXjw6rkyN4zWIXHpv3/6FHT
z5lXTNRh1FNWJp4zu1YKC/h6WKQS5VZavNH0bHo23W8RGme6FRa8l5jpdFIFqUP5
V5e8n1K8aNRw1OevCkJQu7nNBq5/7w0PffHCUIvaPRDaH5u2Zu9N6OKu6MKyzomt
fhJil/yJtSj6+bC3RHd2hfL43PxDIhlG2Z2M9pNu+OzEVMxSjmkV/fGTFzpiOdeb
SEq+ArSfJLH/zNUuLDXtJGFiKtV2D924FbfrLcU/FYZQJUVcgQdLA4Ykbv90MddI
h04b5riMFhy86JNKCkKganlyHy7JbXYH56EnslDZtRlZZsZrnrhoKyts8Ue3m6gr
p35ktyf51DUJ3VEqxTfQGzfHOuzFDdhZLnfx2tt609T8ot8+ARnnSN8Ss3wmxEiW
KxlFxs8BshzogT6Hj3tM5pmQBZWCu6l2OQveZCrDDRlYZxkjzX83/wWVc0p5Kza8
ywavpyNx0mo1VjKKFB7Ac+hQVN9WzzTrCzcX7sLea2u1tU7udT40itBqxEBxqv70
3zmGjmD88FBNbn63+QCrQ9JwzPA6Engzm6Hp9nKf0xh7Ex0dBWjUaakL7Ee8j3N6
5nWGENp5EdbIW6TGs5j6Om0ev9lKKiLItHQWBQMCboV4ctPQ/rtu3ijg4flQObMn
QRQ39b6CmwbNoD97a9tBuYHNqCAbmX9wwjTte8a2vgb4Peix97a10pVkpyMN/uua
yrKrhf9lNLCqpgZD4JeAMbnfsK3P3hEBNiCKA2QaKxRY3mUA9NlNgUl7nNkkQT9X
wqrIxjcAjIGV0T2T9ESgjQzNCZdyW8ouV3kUVsv+HLnyOHLq/ax+pc/pCJG22i/J
uztKsC+ZnYGhzvVz8pn4Zd0h55sE9gL6LCcvjcaXIXvzj9dzX1vFmT1J/fJ/GmtE
CHpkUID0gQ8wv9kJewFUx1WHPZiVl6gqCpVTA5RhARSEoqOR8m59FeepFJObMYBy
aR+mIWRH5SjvqpNMecnftCbsq3OvUbgFPSB+t1DZ2i4NQgZdAHyBC5bdhb9G3qIL
4YARGiC9WuDv2JW0XM63eaqIVvzoPTDFpdEgZ0e372VZS7SkTifNYY3qCZwP+6DE
FkbI1YfPSCpInJSepnL41spXFzrqHxZR5zbn2IIfeJ05JPdI34SGhD9O/QN9dxZo
9NIDLIN82KDcyav+MbpTG0FnvWmj+L4TPHCpy6b/xdvEmby9e+P+xZ4AERaMljwl
hg8xkqT0z5onkobW6XH3YI1mHY7Uft/oRj8cGned4APTJ/4XAjB+vT7YR0J4vtAg
K71JBpLebCRIATtFPxSHdYu1BD6uB+EJq3cEFLY1J7fO+ZyP/HaR9SEKyRUfAPMj
onkauf+/5om8f50OTsCwppBzaXc4tFodxArsBBIWFk1+MJVkRHLjzWQ5WaC5VZZO
2eSe2yamtB6Jl8T2cwRUY1eb1rG8ktGpL7XbjF2/f2y4OSa21YG6jM8G5TF7VG70
zLgCBaKkiaTtNF2sE5dbvdcIGAYlkVGNusMxnb5ifK/BETxLIaoADZcKn3VE1V3T
JrYTx0cq6uj7/2VxxZwSqPB82sNBKRXLoHdbs+0G7MWz/EBycrZoikYTAXmn+/jt
4/sDN/FuJ9gjdfVHxHxZXZKyJt9ZSy/R/LKcMLyIoizoXbSuJcIoMgLXbVf6WM2I
tBrfdB4dTxKj7IkDlgwE9qpmD7i9N9B3EBw075It0508B1MNyK0+vqmQBUrETUtU
hxhIEzYXv+JKgfKcmFWHXEiFD0AS3qTv6FlQonqnl9I3/PofJBGSYgt3aO5LG5yB
x/0FDASxHaMUqnY8bS0wrz0a5No/QVcPflftLXiDrhFc8JXi2fACSxA4OhWk+4u6
dlHCVD3R4oUBtJ1y7nHTRfCVs+R5vtKArcvmvclEok80bbQKH7w7HeyXp4DNP8Tb
js/nPc2OuV6gKYqhCzEd0Au++l4BHjpmuuqZQLXfjOB6VbYHB0VNbIbUvS3EVjsT
Fpq8JvrRg2dsKYktuB6QUJf38XnkUPf2Z6+P5+bMFSgLcsOdz9FYC0jOVP6xXbOD
IhZLA3ZcphyA1h08XZN9zX/BvHC2PMc0gxU+1Z7xXmaifA5uupH8eHw2Gf5kaNzK
5390zHtjUDEcY/pHN0FlYrFuYZzoZSM/ep/g5bLy1C9Qp26EOEhgbvemlnnB2JU8
IC5bw2Uok6b54jiwU6xx5rRxDU3uCJBKordfK3kWqyVdniPFsbBD4Adbrr+KQ6IY
rwBiL1aDG0x5BF/9RNXdGnNOlZJXlTnFWpPy8T7Lx69JKs8AzYR5a2Z697MVzY2Z
h1Jwq6waz6UMtA0yB51RcuPox6cetiq9FQ+pOFl9TzX93EaRLitfw0kIPlqQH+Vh
izZQquQN9Emnm7UD6Z0GqiMpm692qbRMcEvefdBCDBmIV3uwAp48XlBexLb/mzfN
BD3W8iPbzqJww/+C2oit7lNRyyMo00SX538GYvY9quna/Y2EYD5mCYxnxtckBeSg
43vXKIccN5a2ko3Sv3sgJMrIlE6VKo+y5y24CwQsUMcFZAT8cnWFEHWyeXik9vB/
kB00DnPSvZ91uhC9Hs598E2PE2x/6HqnURkJ4qL0/OQINTXE60bNhD8GbAmtxydT
vN4P5pHSQFwzqE+e+FtsibX10AGF54EGiObpv36yF4o7CyXLYZNVgsSGL4Vnbkif
vlr77/SMqzmM46ELvZA5NudAx9hGXPKco9G3cw8cys3z2wA8GvTgRedyyk9qi8uJ
xG7fvlf6AxMX02sfN/82xvrP8+uMqYsjmNJc98uCfEA2+1GfvgPfrWURbW5N3PpC
gk9uf2kWn+atyVwvTNJbGMd/1XKuvuJaM836lHpIJpM1VuWC8ZWpZ0BKlpDtJ95R
VkdtdA4Po25U76GIg6sxZzHFOZZ3Sch/d8d/q8hYB1qfWbzn4cKdGgnbmAASnQQi
TKgm4+JQSGLNfGeNE0qgKxGSLi4OJfe0vqVHg+7L45CkzcqKWRhpdvlP5W1c1loR
LiiAZg81XDxcJlxkHME15cWKT8yUgjReuEt1RLnz0LlT8tgypJiXZ7A1tE21qX2I
So0C/M4xIkocr3/rSZd+1At/ntHa/DBHuK8yfEDtNFHPo7EpAMF48sGexBpO6/gJ
+VOf2VPZZyxhSP9DNs1oDvqmW+N1Q0HfHWduCav4fNlIIPhVk4vvvdjy6HfRQVz7
TsfK5WlWhFgYSjoQRorbRQhJpWDSE4PjMAzgezEGS7totZADTe4xJnZz5T90d+hP
WRSEiY9RVnONR877pR0jGuyEGDv2QLYRI7pM6Vb+lq6cWrFF1RiRBAoxjgHC7x0R
5CTPHXtGzsn8ouwuht1YAJMbfuCjY6UMpsOWVGBKR229+sabh4yyyfS2FO1op1/+
gb9bre211ebKWBTpphMZ2RrbuhrzrFjQ86O9vd/WSE+/+tQhhaFOv3gfAR1Nq4mJ
7hRP/BNu0GvlHdN/aitmR0Ck8fo+4/8Ego5WEAawRRBpQ9y/gmBd1YIcnlZpJqS/
/px621HMM55QvFeUS9cQUocgByOhgjmjyzgxQwnMso/6nDj6zY84sxhrgHM2r/db
T5ifFgcv/GjGpnzfggHrIVQd/TtBYumGp9evgzR/PwN+Kp8Lu2eokXOPCnOZ7LXO
7nrAW6C0DNUgiPeNsVGwBBJC7g9ge2UGmXtooYmHfAh/GqY/kY3RC5XwRJf/SDS2
cekZM6mXF9M8s3Im1JSK0754URfoHEo1sCxXrg24eJ+4Him+CF2GjfV55oQ4UKvB
Gr9PL2bofaoIrVPs8ZP9KC8o1e4F4h1Xnhg9bVCnP+bPwvhoDz1O8nG1sahEiFeF
ZL3A1tmpy3XDAdf1Vtm68lol2mijSj+xr5f6vR5ozJIR7kgimg3htAVGaWfy9Y+Q
qdZ6gviqit/KJIN0xS6nuiyzaLKkpNl6TAX+dvoXvszxN2kiNIo2Xs/l4JJmdcoD
dVt+poTlsKTo1TRMixsV7bPI3mzjJAqDQ7akfCsx2ILJLDDhGZ+eoYILqXOGoLMV
uFop9BPjn6vIPecmfyN3cEWXRmisxhL4qRbhgdSkEioEMSgz15eJz+yXAGXixc5E
2HVA8i5gURPlYWy9OwJR3iSwY9LRKPc5ID1H9zGiI+R0ExhU23O2n37TRk747V7b
To7Xjfv0r+FVwyXVSjs+blxGbZYg04Nb9wNGUIdu//oR/6ZPlC24UCH1tFrRUsCi
vp4KhFMqCQyu7B0lH+TV3Q93wVdUKTDgJYwDq+cUV0SCSpAXsMJut3IbRhtqfgEZ
9mvKcvi+lIR5RbmJZLpPkln2jViWK22kFE4IIfr26GwnCjgmi+VUaoO8n8tofcPT
RMjHU9geTN2GpEe9vsBL8sHsczR40uncnHjmBwvN7TNMNLhzz0xUF3uct7bfUHEe
WJgFryyA0m7blipMUqzpjemKcatRa4Le922r/4t5vcbXuqeklMVM5ZnQyS6bp9f1
+s3dVrwgbNqr/TWIJJAWBeiQ6HF5XzFc+2sRAE87jdVumT4Aq8Ebh7n/zM3agtSp
uVWCO+q1jMWzrbfiUZDhyvufxSMxdvEPjKoh3MqFggzFx7/79Dwe6A6y2EDIxIjw
GGOhI4nJNpL7wTZK8R2OcqFbxEJhvcUCXprehXSu0em36d9wBbbCbunm8fXbFmhW
5kgQINByOJSe2BXps1mTYKPNAIJAAnAZ1T/jrhhsUN0ZXFSYUAu/oZktX0VKmOSN
vQmAr3O2K8WXaYuPixS4VJX9LU3KgAERSIIifywMqPHNZnmTiey++XOgI4k05a1q
a8JC/Qp+fCvBC4q3k11QBL2uTR09qTaJqQZp5G6EtNyP4WNy8rSrzpMWSdIxnV++
c3Sxj7LW9CyKocgm3M/+jnJtkplX97VyviyXN5/IwddX++DNLIeUoIYwDkJkx/iO
R+KGC275wUbOsdPM4k9U4D1/+COgMyGMk4KARHJ193x8bNjixMv1PkKf9TTUX8Nk
sKO+r63A2Zvp2OpvJM9k30uw2siWA1HovGIYFHQH+SUkTPiZtoI05yiO8QgP4yoo
cs7JumUGoDctbp27BfvaeDUuClhaGRAH2PmWt9nZBIUTQdEDbz0kqzNaZ5DKdO3V
y+XMx3L0RdQX3HHLmCnYXzjXA7Xf0XhiKtyezyEb4uft9vKzlaRVGZujtEifl9sh
l8NQb4AsrNTW58BlBo957EVys+wppblOssZzc47G8TgDJGkGYO2hDdEwYCJMdoPV
fFfTFEavAdis3xvx4HeiKWjxwHb2UeZlww+3jaW9Jry3+x8KGwwUjfJ1S6qo88fM
6VcAUfvN9Rb1gQ2Otdbd5dbcKdXTnsq7ayoKTgGu7Jm0wyUFdk7kDDbYCw/wfNEK
GpDz1bwAZ5hBPUdFEJtBwg8fZt6aGz6ImYvFbXF9A3HhQacpaWZQYrM3OAJdNoAD
Y+EwmxTKkRjFua+DS+fMP8RWmj7t3gSB/8NBwWW3ANsy4l9M0sGYYFlbqvFNUbbF
lXCsVzp2EOorM9+P5cIIJUPsET4jhZVCDtoIwRK3BRylW1xup1HsS2/wDykELyTG
ZGQk9QodFPsgsxV/7tWRlxtHQOxnWtYRVysqQ5JFOUUkGkgzaKwc9jwd6gVqJ+pc
E0c2PF4nCpK6Qkw3tjB7bAw3Q05TQs9pXWkuQ3q0KxCPxPlTg7ss9EIpeQRVnUH3
Yb63xNdI6/Zu0h3JMNteW9xqezggVdRQdwommu3RmaXTofP/9fFqKbu8uuGSfTVs
ZujbJBLj4EU7UoTMvuJQlDANLncaYtovo7nEOf46ZCnixlOfyXJAwGENcss62Px8
6wptBKeVmp91lowbZ69e9gmYCs1Fm+HuuNgilcbIVBWkNS+D5cL+rCPwKWs95c3z
9dPBnRZ7tPZti2BSUOI/k9TN7cDKSvKMtMd/V/UA8IxvgvU1Zh2Ql3kdftonFr+g
5SO1+6U4uv3+Q+UMf/ykYTxBn8X244X4saJ/LiiwIyR51XoB64VVL3Zvtoe66R3O
FPJoU0PVTz1/jrE1hanobjNQu+UqEI9VZCoUYJRCIqib5D81OKtXpFPmlk1A42SG
e/QYtkfZBP3Gr3c71SIMcs3S58/UAxwKnGwteSUPrxxQ0orIzUD9Ra/1jjpBAz4R
rd+C6GJfefEp3i5VyzQIi4h6plh+eBJ47PnFu7RnEluKu+GCeTIMa9bqfAKDUhLy
W/B8QQLtRpIq6IA5uZTFGk/2VINQD3Tf0WtS/J+JlhCp5pmVBHPx8eiYCBUffkxU
dG+HRM2+dVAgSjhNqdrmuxp06J5silsM2PZqT6YEI8A+R7YB6bwu4zwyedNOfOKV
ZuvpgeL03fPP4/rkg/dvojdx3SRMDr36CVatoLayrotVwknejXv7IDFUIRK4/xbW
558AclCbcYp6tcWNB58k7vZ9QR7YL562MTIalszf4n/eN4X9Fu7aovj5FJtMtmW2
+bLqvPZnBnPeeEc60JX25G9+w9+Wgqp3ru2xTm2RdIswZTXJ0Wo+7nhL+BueFXBY
BmvoBVRGot1sDGrPYOSSpbDVog6Y9+YuJVi9MAawtAZNMtJfmqpZB+XSROkD46Cw
P465DKvrDy7gOSqDT5qeIdi/62b/U9jupEACEiOMUaWOCCKwD5sq2I8dfeNruspx
e8cCcb4eAH7mRcJJGjLAihY6Aj0tYBEW/a17aRNmMPIjOd+EkHhqXRWKW/ZkbXdO
MVwNPKnVMxSPYlaD7ELOmcgdljGVNrqEWLvWxNaCj0SQ/Mm4bgy0gvbEPZTXiXKs
HcKoxT8auL2q7QzJwZ/J0SQNc061mBMM+mPTh4ST11LgCPXlNyNPkOC911cdMf9M
4ZaWnZU1CT7QL9PCwP5Zs6P777TS55yx1JzzotLAl3Pos3/66eYyXLZiS4fGsX32
2OjU6V3gY4eAhdjdmlB/S/TYHXUD4LRIXf34pPIJOEl5FoL+5OP/DRN86Hv0CJ/8
oAoSxEIr77kYqwvYNi+09wxEs8p3SxbZ7Z7+NxnbgzA/g+VCrtd2hj7+Wija8qUK
FCcJP7BuBcXXzuwMQ2v66fxTIY6+FNaDhJXfBZifnRO0XWTIsPfjMdHmBNOS6S38
hxKY2IIw7vWKJIsg+NNO14XQcUkDxJhBmdB+VHC1pAL+2AcVXPqw50hjPOomxO5f
Q8KT3XWgWRpBOJLYPKOdckVgdh9XY1lLWsPlC6Vj6w7O3nkhDOHXvffdw09GmuHq
xnDSoOTaUxTQqt6vcvxLij5UrKRXgt0IlnYoQXUYJfLub+Ai8mbghpVD/7bsQ/cJ
pcDlX8o48dFR5/Zfc59DjJHt19SdTqPhWM12sA2h5E2HsCrGXXGCxx4QO5AWquhb
xfVCII/P6AiY5EISXaB8ASnk6Sux4didKNgtQfq08imLwyirTr/+Otx2m43X9lWR
hBQWF4VpaMBLbLNkpWmWEs4oVhrNZVxfdHFSzd/zINfEU/y2Hsu55pIi49GwsbzP
ntiMErUXS7FmA/GAiRD3GMRBSGsgUbG2VZ6uNFev3laeqvQwLWCiyxFCKfEzlfo+
BQgkR5wneTOKMg8JeZ4MSNBWs3ors50LQ1jxqD/GCJeHixmNrBREH+4R6AvIr79R
B+hCKvHs21mflmsgZ+/91/4EGIabo4rAh/JrH5YvQ/+4W6mELcMiypTHOmqQAmxU
Os7/8X1VomU9yp+TBZUPO6qt/7dpDsgt35kn06o16YMrBbe27idr7v0JaXLsCRnh
XR10E91X8ZXDjL+ZKB8Lp1Mcs8C5DidDt+vxQNmbLt8crVfsGxTDcpIJMayc68gw
oz4A0vTvyclf/VHons3/3vJ2yNMcApeUlw0SKB93raOO+YkWC3Tte8MCL9BSvC1z
lawq0d31XxaHVlFQBByZEsF80Z5aB9XW71OaRaXm2lbMBPwqouBuRn+BV788Lnoc
nYYHIYSeXDy+VEvgnK0YdaWU0Pbw7bJCwN7q+hbWPC3BKE9Mzs3rHr9MEBHHJFC6
viXSnA+DklV6R9tO1WgR5Bd8s3avdFe+t3vLiHJ2MwLneFG0j4jcMiVbFM4kIKXe
RqTXI7oxUJFqNvsvB+evYNgycEpiw2uLaPUEu9ffYfZeXdWi/5Q/XcZdRjZ9gdtE
UhFv7spHdrjawKwsROWpaswf7b5U2dt+zx9hQ7wjlPiyC8hWabP9EoXsHlyE77Cy
DU02Kv+KIs0y9TFzoD5C5EO3BI8l2J/QlOJBxmfnolgid4ih9FIOQ9FBlOJqEzzX
5GXVEtBeiQW6IWiPZt+z+/1Z+K5ILi/kCS40e34OUIl2PcsuTx5eTuCthn+V2zQd
/ajdSAwC81vytKRSO82ANsrdBmMU9u4XwnwgQPmfLFlIbskxEoHYYx4ahzVFO7IY
vyKiGVTSprExaEKGcFVj0CMe/Ud8LGSUGNGFjdGRuNzu3kMPsZr/Uk/GbOwDrWcx
9t1T31DL2BIiQneQYVfxTvKEKCk35qsBXmOZC12yoq1EAJewXKshu9Um/mNPjHof
UwWGkOVDzuvL7D6Bupd2rlCAkELl4o9SB77n4FRWfud5mihOfJR/KriINUT34SwU
Pn/AnlP449+RKqftz8nvW7PBE3hxatiz8mkOIY7A9dT8Zx3Ek0QQ6i9CHvOENXE7
uQFje38CdLc3frRGyYrzn1nvNivZEaLgEJm7tx9+qo3CuUghiedqlQFn9wkEUFbE
jxTsh4e0UqD4D8occuYk+4KV0krP3jo888E06ZklSSbeGqCXcJAA346UNzrGu2gc
bkUItwf/F+N27NJQbeZleGWw8V7sIxuKHeImsOSrB1Uy/d22LDPNuFVBliY3jf2H
UAsPWEas3IY4mrhH/rz4zKumiJsd4hNte/47Sbsr6BoyV2yP9KXc0es0AlCPQeH/
2fUH9JWX87+kkxYvIGsG11S9zCUJCKPn/ibBSzXUIBWy1tl54bEQGaOjOiZvrZyS
NPQJ4LVgd/g5hcU1lFC4yRE2D+l5rg2D2vun3R7nfxck7affW0MOnL/ezmtmMyFT
IbMQV0+qJv2enn4VOavJQpnsc7R3I9G1ZOrv/5ITM1wKG6NZVQPwuQJrK6CDjepg
VOFTcqxQKvfN2byKFyjmKzj2xxSgz/vDYPJ7VZSl4s3FX9Ql9CFHztDPg6y24PnZ
7wTEzVSu5OpEAoLo0iQcvELOeGQJg4wSTc8kwj9dZuwi4uR3z9lx9936edV+iLb2
Ytb1YQKA4Py4qc0H7S9b98u7haXTvSRQDAV0AOosZonS9ATXbgBpaBogciPrLxVI
LdV2vkvj36h3d2VYbccRWGAIvIWTURq//HnBdLlDqzEFTgWo4ATa6HnwHbkQOuvz
wqbMiaX/85wjyC7PfwoZ9HohzBQJWOEnj4h0Pke/4XvTdNkU2ecmVd+qjvlbYdpm
aPjV/XxlIUFE0ABbhZcb0sYb41SC740Mu46nzjNFmwdf/a/HLMkrxpBBlLym2s7N
Fh0waBxDAE6Zx3uhGyDLBpAiC36srM9l1eG5kfBAAFil326Al1bKeSUA7K56uX3a
2z0LAJhE9HMdGoWYUU3KLVnhkWolzqVg3w/QUrEkUeqSC04GodTGoUVoB7hDiA+l
02YS0rjmdBjFyrNT6yY+AIepg4ClyBbiVXhk6ZQn+4O8S/5PObSHh9mluiEMibQ0
Nb9AkwG1ruLPR9oYULW+9yOBPEw1z0L3s3E4JzF2W4eerC74YwSMJBLHmpGJ37ik
N5xSpMZOwxVV3CLEieCiOOcHsN0eEIcRM0KlCjNIYL+dGtjf9LA+3PWCGJeOEx0W
hJi2fHaTXAmNooV6UPcDBBV0NJ6mgMx+xpzj6LRzgGUdcw/2K1RIiFbyFNC/twW2
EypTlqrKUAbiz95IbUpalhPIOnnCDMYx5Xdruq5Yp7Wo0CkJQywCz2wtnTA6q21p
CxgjNgXDwfNfFTZ+naiGKgRmOZVQ4Q4SBaSStQ8jIgQfERgz7aCYh0he29tGgoBu
pacLwWaBQxtatv/rmlErjqKd/fMs4c8+01fCXaFXNBMmWkUJlBWj1m+l3q/B6F6T
P4nh5cXZ+tugVe0zjt4A/H9MyxZBgMBtNg51Jo04XPfoilejHXtPjrQFVoF0FqVF
q8pTR+K51dZt6xKsJhDIGwWYILXc+Z9aLd/p7EpiG0z7WDh1wESQDFPjH/66Rldd
Dz8SsQ94uPOhWP2cObFzph5lL/Pbhoc1mnW0/dxNjdaVXO6HjsZwl6t6gHD5Pzvv
wQHUUSmm6DLIae6J1hxNFPGlfFq6cbXmXnQvphWzNF2ZAC1OtLK87O/mi3em60Eg
/93fkaAAFAvo+/fhEqOe08F7GyBIYcLdBjb0I1z/JoieNweYj3mV7oUSOePxDY4S
T0Yvtyb6jpC9wp5T8gWpPIEHhvv0rbB63aDUY6scThiu7FWRvcxyv3P3068022qG
k9gBZXxaw49N4uQA8tx6hb7OX6HVrITy4fKHPDQX3iPuEjUR2GPYTKIbpYxlznK8
qoAAVSMfPw1uBgykVbEeNh5VFmvY3s+ldKH74I5DjXnTZSOb3eKS0zq6q5CaZcUC
b+3U+9WeAIOe/d7FD4spEuA5W6WxAgayKA88m1PFpnOwYNOayn0GCIthvTvDlUO2
WhuZ4QXqT/GaFw+iWZeGRiUKR+6LIT+VsZJBW1wqqh+wbGOlXMfp1oFCE4Emhb1/
XDenI5bOGiDJq0V044IdFzMUxjHrCRX8Dp3cm8temUOOsl/Dy4QZqjK8R7qD7WER
oBrVuzUJb1oiaMZp+woJlmMpp7FMSLzl4XGFz5nJPMEuLBMYg2mmeyqZ/Li0g1QA
1Li32cuZyxtE69k6ZHFw6SsQj9NWfvnaTIWChtRpXA8ldM+3oMBibIvPlQtAHzWt
KQDJICtn7dWCMeB/7ueEa9FQBcm90GeDfCsIFLZyNNUsI1Ev/HuozMdL5Lr0aXFk
U4fcVVow+MLxbNP/dj0PKOlf6K/1oOD9atVpaj3jR3L12TBuobLJUSxStpQQxqdd
dq8au+CXzJ6I/lHwDxMbUfXLWwHsfX7JflDBLqybz7mEikr1nAwxdHEo60jIIE+1
1Uk3ZjBb5FILzWXmvjIhC6jvpCdLWEQ8qeddEJGeXC33D67jfA2PLuvJWqoIVmY6
QLS2qYaV+n0Z3oV25Obhfa0zpRuFctPCrAwu6bKSJKsp4/CUItC3C84IPecIz8ln
avveNLwYKtA3t/nTtDJxJl1bG1eeSTl9QpA8D3J1m6vdjjQgdbn4hvBPeBfEqJ4m
3ZnEf2EPN/p3zjM7nTwYO9YJL8yXsfz+P3sGk+sPPs8q3a+FJj7xJH6OT155Uv7l
uVUlKPYWgClJ4bDxpEwvdhrk/6ExX/KDg6hCgCmJlZlARJqCOwLzkUkZcFJ+jjae
MP1Mn7QvqoNcOGBuK6CI9YWUYnuAC72bwnuBLL3N7/GutcyselgFH+/nD+uDT3uN
si46U+tJ9zuMpUOPpyAtEqb4E0ADRZBtAy+VkGnWC300x04jZjDJaW7P+/lPweUS
LXtFsWP27kNir5K0tgIcOhUjJ8OnzS1DHe799mWcsWWhDF3vQ/yMInIe68p1L7fC
XXInYGtdfM/LUbmx6viAptd4v+bT1yDwnRwyJ2RV4ivoXMUL3bvh+VagY/T89ju8
yLQc5xJPeiQiTz6bAJCdFZ7ETAl+bIqwvpdkzPhguQzrp4uKzQHu195KmG6Zhh1U
0P6fHpr+ePDfPzplPAmcp44ABryo+aG32mnjjT/jRmmpzvHnEnGrbQ9h4yJimmKw
lM/T9WXI46XLhSi3PAmpJlzgdZz9VofhhTEv+ijkjQ8oiZkWHeSbXlcsCj8u8ITo
8DynVt6nfQg9wLPhzILvDAURqYlKpx6JY0EDgepayySQokBTpZlQ3IRfaFydYoYn
1Ibe5G1jDjx/ym3LEmjhSn5nrzvVG5tphC+TlG9Nf2jnwYR7f+ZONKaA3eAW3M9w
mosags6Iyzpg+5kgmGpuiGtn+WjPuyn2Jsr+w5EfZHdezml7i6Etf18j3z0XXNJx
o+GqVx/QeXEz0T2psnf8Bm8Z47L7JkIzevK11D+crrfrL7hED+1dNylG2mBbcCzN
ywI4zAhGcqT7PQv+aI8VSdmlSjApKYZSkShG8xy4cqRyxPf/8OnjXhfVQLYt6kHz
7AKKns6WQBzgv86fUp9odduk8ImbA+6CtlJARJWpMjede9CP9Wfk8C3yjZZ2daIH
sIKFML36AWOxUWunSJWaDJ7/9cRjvq7WY1aiFBnTdl2QvDLXB3n7EUjalLzR4j6U
e5aJ1jTvCFC1HXaB5jQQXHqfMbGmwaMS7gUrz6i2885qR8Lhf/pXglqgUb8GY0FV
q9H9BLeaYmq6DSnFo+wX9rkcUP/x0/ZDayWYDFUftysScFC6Bth+zuzbVOzt6UpA
T8FF9EfLt+l6tb8I5OoO7yC+FlpsK8eCJF/NKAAYyg3uRxMynNZyRBRnzSJhpMFV
GsDYruLd/iORGod9q4Z4DISEjmOkH5tOxd1R2bWMB3spQyfCEPj3Mb2cSr9CVxoQ
yKZTZJpJcfVuCKI/dwYY79qoWE05c5wqtML3gasqoC4BP6CIzAgB/K8E5fwrzwQW
CSYOBfGznfyHv0WN+TuN22VYiTKDd345ioZ5kqmCRDrUDKhmnh5V874fIc+RstPV
/tGz+zKIDsm1Se1yr0tzSeI+MGBGWx7vtXV5ufrqSVCQEwH4OeaWCKo7R8mtPiBf
uncJ3AiLcSKabzc4r3Pjy0K8Em7QSwFTJYMX1Uv20JMiMJJYFNcmW0NTqV+n/Fq3
WLe2KOX+LUEbLVpr/+1gbVhPim4cRjGbzLkvad/S86wouyjprqf75mn1qUYXAYW7
bml96FBbxiXxL5i0aKJJbrC4GNX+89t2/okGzzkS4Zpv19eGRuPG6Iu1H9rqXArM
Kk2O3bzyeyVkHEHnN/dOLpezE0byQSO4TRLdzgYvS+lfzGtLFwCSbnwlHH339pCD
eozYpSbDYHC/0/l7QFXLIinavRykJ3gtdkh6fw62rJ5XQfZ9PX2OBmKrjjOljHgF
34yIyFVoh5jQqHnZE0EHo5nhyDJs5yO1Z+cwXNJtiP3O8rEOr1SQLw2bSGBKT8Uj
UwZazEuZT8Rc+fV1XYLzFNG9pJ3qLJLvXBv1F1kZ0K9mdcwbI71/1wGnL5TuIyB0
6bJ0zXGw9lw6yDw5HGV8JTcLza90B/dAYJTVUHb7lsYAyFJykKJuHZDPgdHC9BvI
yWc//vRMKuWGoiT5VQfredrXu+EDeVBWzEqIGIItykP5afdDVaA8qW9pA4BHzy3y
1okSLM3zV3HM3dVQafwUrFAND5vCiJR7a3Zljt+rETT21CYz5+sCYneQlnn8pTJA
6jCAk+Xsw53/6uCP0Sx1noVX1VrXELMHnw15TgrBiSSF1VLoDIbXbxkq26ljyW6i
tyF2xXktL2amTNqXrRR2Ip24XEm41v7EqtnPeJqO6MCxiYr6O/JuvohBB5DexHxx
x5VoVsHBHAUbpYAQh64pxigUTip1sKAztkmvfthlQIndURdxLu+JFi352Hk/7V05
n7BGMO+BfkWiWQKsTl5mSZoAH+PqbS0JV+QZX3+KkjrNpqykXfiVNgKp947niPw6
A5haIBSo+Sl+J3VtWpPqXLMBJSioAl75l1uLlnILGDHN+EnqM9DK7Ky6tfpSnjFh
B1j4EwXoAwDxjN0q9+u0bsxpwvsXAd87kz8ShPy2zan/N5nJmG9aL+n/1YKdYqEd
0iS7RvZ/6YFG6Zhzk/moP5Fp9EsJ9AagkeKSPQTb99lJg17JtuCllZiqVuzVECgd
B3K95KxWELiLbc4uJgIwxYTGjUh7/cdR4LjLXZQJ7gQVYxvBvRizzzC1Kp02oH7+
9GdZ4mn7EXMKY86pxtzK60YUy7o7Yi81pmUc6/UASpzr/b4rHPwRNVMokQcqE0lC
Mz+uNJbbfHdcQQEuNhVoKM5kQR5/LYNgm/PlRl1VQsoHeMmLCm1niIM+8Qq9mqCU
cnEyA3l8y0okaCsFvmmpzoj8fwgmmGOS6csQ78JMD1aU7DX9K+VXNSNdoOXHYUOg
aQLlbFHW86ajc7dzheoXPjrt2dl+wN85NtcrftYmeBZFnnsn4vzkAaG+6AOgvjQs
kXIu59OTvrfDOKnQV+5MNvvYNthlTsCNkw7LSQNmyVF7GpqLg4GJVErlwwhWkmyv
VASExToBn+wuMDKnoxQEQHjYvt5pZj1qJm/D6FbuOy71oziItBNcCelKF6saNmnc
15YR7J7Jv4akk2tAZ8BMdDtuVVjA19k+2Co8hQd/RFdZnogkrLbN+rJ+qV/F8qv7
O6KpSRpIDJ0y7N+E/VISeNWnok3Yf26ShfEeh0LYz4JJ+r0VHbTrO6cktJEcRKDd
n8RHwFG2kQ0A+M/ifxVBh5BwgIhJ3sHHURsIPtvC4IuFIih8UWe2pVxf85aySCfP
+dtRh9I8IkQ8Wbv/EYEzb6fbk4Ddp6ura4FevHfM7qYUqXjDhh1qruhQEYCumX/4
eHY1bbYcNGn54nr0BBVKhEEYLyMTXtZyNLms/DU6G8C488K7cH5EeT/yyMFAOUFL
BrNPUpP8rkitXjyrgpI1JYX2/D2L5pbnRR8Xux5avqaKKOLOEsi6Agse3k/JZjDr
xYwZsOHYS1teFMI2Y0YBRpPY5NBYIJmHXr8aDGkUV7vxekBjzL7nBMiJ/SO+YyUa
qzwLubxXwVLCLQRPQkkKUBHa+0v+tVbhGffW8LEG1CA52nZP03ZglFkc3DPrHavA
p/E/v3Pi6gPveTDzY5+ELQYAedCxaAzAH8Ut7qmdJlI9tT+6OHixMWQG2T2ttMli
DaHvvsIu9lCMhWObfF1CsJDa2GUz5fM+OYXZUuilHdipgUbhS3fcex6fSgi4TsnL
c0EpDxFR+H/TAlNUctyDdpgvn+lYCb4/Kh/F1mVAgwh2eVjQdou1Krmv8UwmxdIf
kfn08pMhrEuvOW+Vvr8K+rwN0PyK+imPb77IlIW/LAaHDkgtBGexgnhQBp/OsDyE
2tTCr82r7RwJaLm6t7U0cClFwbjUA/qeXJUE+QNTQob0486rw/d20JWZaDibNAqs
2vz2/BmwSDdqLHOSkudCY7zifUcML/TOv/Xk23Wb6PdgHROTw2nES5OCM/XPIfga
vBtTIIyGaYQhdHRJiPrB++sBI6jEe1ddHx277MxKUB2d5slmAuQLNO28ieVVJ+nQ
numKP9VEP7bAOIGZ+M5kXaRFlduEiYXgcmDnLfN3gBfKbXHJIoWc62adjKJ1aa7H
++8HjxVPEHSiWqL+5Oqoye0rKHuzCdq3/6hD0ADYXfYNRRQ5eileJzWQmvoiZYLm
+oymddvTJ8Eg2LxXEjh9EFx6A6vCJPD7Ktp6xATcyz2rk9OBTeT4cqZQfQhnU3uB
KoOkkM3eJtzVD1jDQurF/b9UQjp7kDWLWXsf17ladTXzHO+Umfn3QHHZmPHlrfn0
5/f2wORmKdv2c1oIhqEZ87W/nTL7VrKZoXw5MJxdVXImCh23S9hlz8E8uagKebhd
2GpVCjmeIsW/KH27lQ7J58xiSPUMJQLGwfau+3/ZiCgki5L+oYv1fSJtg5/y0DIO
RO4Y5M0xTVPBWaxoOqlEIHxr6jyw0zgalWMEe1+Aeg5mvwDZLWBdNjpC4gwAxomb
7UgnovbZPEyNUe/p3RvaMLwxgRr4nU805UtsWL7bOO/WEBJw9wa1l9fYRwVFopgA
W9aZ/i+5zT0li6glvQH6ZcepFKBuJCJdf2lvrmLwcJ22M13j2NnrnVTgmlketStV
cfTnS2FJ5CD401v2WaEF0SFbhz+MPwMrBi0ecVN2WsIKvuCoGgiXcuApwQqeDvXx
Cvwv51a63iLx6VCx4R0AFYTsvbBhJkMQaizY2bQG8B50aULiYOkMPGr7Z0d5VGv3
zGubooRo9e3GFzHXFmNC7pKt7F6x0yj91ymEZdiBWl0+1dnVSdHimkZLNhe7FsjZ
YaLwxGFPvYuq6UMgt26nlkggDq6ypZzmauzNhENbLXkNovBuuURlZV/S3TCZ8QtE
e9KFASVvs89M2B5l8I/e+leZ1YXaWyEtKZIoUNhcSedPcH9M0s/TYuOk6lLFqasJ
YOTVlGqdvM/fE3s4u/Q/Bdp3ak5Oy+88m3dU4aj6jzyLagkPISAabi8iRlx/bjkg
3vYJwjehesUhsRxlbF7UFy2l2EI4VsNmG+9iBhHnvYzZDhKuT7uLd3UYcYImiIui
QWR1t+9e+h7jGagvWwQ8QD5MLGtccDlD2EmcZXFY/UUcV4hxxDkkA0zxTDTXr/3c
79OeZJZsalv4RPn0GRodJfJg50W0rB2/UZWYPqZBt93r8fPYxuddzA2sp3GwzueO
Uqbo4N6b0zdzSy/Z1+k9Arz7J6Ib12axl4RpGtcAwPv0pOuPowfRr4GdSF+kO7Pn
0x06mq+EQjNfO2VW+OxF6Ff716iBYiGLbWfgXyGUIe3Smn2Kct8LcDG7RObsMnN6
nPIxebu/nkMDtfPcyKwa5l5HE5E6TdT9Ghf6R0D9acnI5VMioysx/n6I6P+/uh2p
LJpSX1o4DBsiHnYlvo8t4VQYtxhJEvvj6jQiMsLlmpvgQquunWUQzzeURXrIg/Ct
pLaHExEzJ0xQ54gQ3PrhDVzuw/HAUiEop4wV9cfCJuWskThTpi9+2V/u+fw1Lf18
XtCpSvhLhsr5MvzRnHjSc1RRf5vvxDcW9VhjyzbnI5BHEbkMbhFBkLWPbAmWEuFP
TeixYGcb42DYPAf0YJV9aK/ooA4qLxQCU+VQGXap7xJ7GeH4rTpKIYzpwYRe04Bv
Z63nz+Eg08HBnNgZqZhCL739pDRE7pMputaruvQbSdOf5elNu1LCIs/zB4AF6Y2E
0M/y6FlFZqLKH6v0Pf6vf/s/rp8nlAp+XkO7YaTaAz+8KASn4NFEQ6fYow1AkX7r
lDf9Afo/fneEQvKkOd4vp2l6pdHBsg6uIyqNWFRYxHpVofL9jtFxPI8om3TEYplv
2HysKlTdYS/GpwlsBMZnIJYxI0TVlMmCV+SUm8lK6SQA4oNtNOJBxldH53lqSzgs
C5LhYkKTmsH1IguA86dozj2ZlWa2KwvHuO0hWuFlrAbC2/ItZphwOG8KELD4rM/R
Z6XUZcuaOH57lU1Ep5D/KeRR8WLkXOlE1C8GNAnYGW3QpqoF5CosVLWBTjVshKM9
xKBXXo/k2Dt16RagKoV/YcbvabcoMS183Q/VQ0YVudKzJhLHq9tXbo/K33pLFNj5
q7ih66O3FDBw5Y2ph5sjOmy9Pvh4141XPlAJi7asdZaI7MH0C4nhsWBtdi7oK829
LaVZ/QdNvZ0UaYbbqdnUndRErCYAWQACa/JBlO+I4+ZNMI0x7yMU7UuNh7gdwv8v
5j0NeUioo24xpgr7RMXw8+Ln0l2dAUDsnsh0PpYP27WOZK1KEJaa3hCQmBMZEb2H
4BJqMyGVwCiOV1ZEsuixkQzqQJ10VrfidGbsWYA5Ox6aP8LCcLPIcHyQmc8IFR70
qIw05IUD9jIKcKqCNjuuVJv8O3+rQW/SA9jgyNMvKQAUlrlzG3uL20zF79oUIxj7
Guhz9x/KymDc1Tp8EwZ3Ucp9F48Dm7BhB55MJSo2XSFQMq4ue3OABUhz6KZsxv28
CtsypUwHidEhhCvDZS2r2ycbHEc0JibtpSHU/CgBz59T8itkIetcUFLVOvYF2+57
dOhTZmXK0Lq/gLklMsh9jGyWqeUjXpA61dUknlhsUfsB3JkLsYDazN4G0GWp/H0h
v3moW3Ysxp9mV0VUNBS8dLNdnex6FV74xTp5XO81+lk+ie04kDmUCYE2it7rItJ3
DZ7LyJo84OxsTvQuBd+s/lVKFYCj3Bf04uGDmL7dPXEA4UQGakrdGpGrgeGbbphR
mtU2Jfp/zE3+sKB7wAWVNlCH7pemXkfqzFD++zrpvLVFfz4RQ9xXqh+I8u0EBijE
FomypLHNtBisQO9iQOqsI7Tb0M3Ej1kOZAKAteOGxTnzalV2IZlA0DkkUCiTD789
H0AqyJ9YCAIHOuN6oqeltNSw5ImuTcDI33f2sDAdrdLfCmvNZcg2UJjNNTNV8a/t
PE7MsCTuEwqyy75Dmo4k25ilqsz5u7NRxP+3GYwcYmqf8RHDBApu9A4CFWLkfBZ6
eUto0gcRT6nVb0AH1Be2Gqso3nt2NZiGlQXPXf1wbvhUKgHGVsDXx1AUaVGZXdP3
2U1uRdbbz2Q9786I1TeoJ+s2QIUYUQB4GoPgz2Rcq0Ob6pYx94eCWbzLZ4k8u1UL
O0n7zX+7VOdF8G2QRrRTlOtrDmn92JexYWlsQ0GxdLjXaTZ0bHktc81XhxWhEo80
9Xi+JJZg5eZNpiChgSTap3Ha7q4oxErwwO2XApD5t4l1Min/vQGu2F2LrErp3J2r
PY6A5tnIlRLzbctJB2OoONCecpuMZY3/7fbaQq/TMf7zPFbKQwbI7V4tnlFjtJPJ
fCYglyWkNevxDogQVdfq04WLfCBPCCS/ZsoBY+JwM3Fu2bd1uiJMl++blj02r/Vm
2i4wJytAuQ89PrfR9VgO7AUNyf3OujgsWYIJ+64p5UuZ3zyo/d+7laZh1neZmITM
vvvcplIRRGcHf8ApQGwewfYbfgj2y+6qtEGNkECdaCCuB6q4hnahE+rVaTvDl+DN
bW01KVm42LETsUhXqEpttCAYLtk5XbQRn2peOuVwTCywi7/5/iIjAJuGEB82qokr
EfYYP1ZLXM4smF6NXQX3SSdPG4l9jhpb56+0A6OjPjut+mF6b5zoYCYpb9nBA5Nm
ekt+kMUG8pNULxGKSg3ZwLhWrfROMvuTglvkcapv7W5EXT7JJQRYH4/GhRYVCPTa
KNMTj8RFwFKcTp9Xxc0KIDiCBnEKDAxTBOw27o8asA7TdeKJc5XT0mNSkRKA3Ola
3+t8KG7e+iTm32NoelO7Ia/YIxG+KdEMpawG7yV39b5DNs8CTa3PUe4olndNHsBv
gxTfZJle7cOflsM/oZ0N/vALzrkmbva+DMHLfuIh3YuRKznSvckd5bRnq1yryoOI
m+7xBCRzqwe9bOc7I0+y2LpZ3q3ENr7RG9h5r09Uaj6/jJqqF4lp7Hm078TBnN/R
z1QlAyW1GU4RjKXNSaBzfYRj4Da4Xy7Mb5Vt8LJRUu4Mx3b3E6qrz5yg3+6uQXR/
ey4zJ2I99phTjKCuHMgHOXSdDpKA2r0nd/7Y7SkwbMnzUeAl47267WZgIIqyay0n
TynoEjjm9uydZvY0yJmmBW9Am6rI7oXUEcy2mPVHrXNQ7MBnexhVtvmUQEknPS2i
tYbDE43o4DCbog2/mHiSbwATLr7//x8vU+DXrahUneTPijil+YfZhgAAtUR1XEpp
/fuvG54ewxXh3+7Qo0RNbGWhuXEPGKEIDDZhiPse7gla6tVebxKOKw5JgWnaQTiw
TKBzZ4lWFsvAjqNwGv2wIFHeNtJ+zVjHXS+wPhdmepNAQoSYoALMSQ2XN8gMjnxS
a4qdN/rbcgtbM5ei2px41VY79Xri0ymxUVyi1Fl7WdjfCViBFwtHCD5TuwZUJX8N
cJFJanLygZY035PY1LQBXvnB6cV9Fs5Sdg5tqUTdZN3F/7ZAmiK4u3PbLsJbLU/d
0stJFqcbi82JqMgW3k4MStLDTVM66GBPD3qURbs+eQL23nfIO/Ho9eGR3pNM5t5Y
kzowzDX7+BTPsvZ/iY40eH0LyladuvTKV41Rq+UqELpp4pu9EYwTXcAw7AY6vXMH
Dl1gxgYfhyXhtcP9TTz2a9Nofvm5aesosFh13VYIrejlfgtc9NTIbGV20VpuuG+Q
H+NjInUW/EXYLfNi2pK0ZgOQWinmsrWEbbAMpvVQjjqT344RUVj/uwdivFFaMZFI
gBEulhmU7BMoJ4wYMtLPTMNM2uxT/k+xhSlK8JnSWSm+nloT20af8GLqCwiVr+KM
I3RrTaRDhT2bmhjKjWKMa768Jcp/pFmFBghjtlu7z6hWzOJDEyRasOnenkyhas9b
lwcCK88NKLYw5Hp0ZVe7P7eTGGdkHrdQbjs3vFW479pki2D9DwNPi1Jit2qtawzx
6vJYC2lEC7ZwhHy5tEo6BaW0KcWn83HOMnfxW2GPraww5p1Z0+hKgiFw9u4JvVvH
pk7as8L4NfxUxiRYoSSyDhhhOwPaOPWar7/UyL/5CssPW0Uq3x1gtbQfqS9OqteF
wNPCrgGtXhvwzaST28qr803kqqtXa80AxnDGXF2HmTF5NnKSxejus00oAeCL6UbC
YAKrJ0y7efxQWF0i5gu3d9mmE9tk5E4N4nCTkxxiw4NMFqR6l74p060m43581joG
x5NBMydHOFBmwqU/aeSznojYxduRx1SzPs/nyPrk1ZF6BmL0v3N83EJiefqPLkuZ
2WBn1Q/6/JflXcG3XzlqcdNHyYHaZ+Os7nK9kIzkUdLWgQc2oghHPxxdtbEem901
gpWSeXt/1W7QVq39R80C3nxclTN0MqyFItwz8ZGkS+YOARI+KLm7Bd0gmt8Utf3n
/s9cicbdKjqZkbfVwAo/1ZB6EW/FLmGZscw/ejiTW0pIJs43R6tBtjjo5IXLsgvt
gyknH+k0cJWB77GQq+f2OLMZof5tzWROvQiSQCJUAp6cGtvLR50tYvSwZpOwZrTh
mTItJ222fpskFQNqAf7ayVFMvGrzk6gtLWHsoCYjCHK4ECHkMBSZN4HYmR8nrqp8
SBQaGXq7fl5kzDvR4Juk8Y5MkjCMYwxMegcqQBukr1xJM4sJIGX25WOScI4+5m5Y
NLFkrnKWGk2FSKspnS4938R3Z982eo+P/Cc+6wHveGEo9gz7WwogMgOudQgkLq5c
+esyQpPDXLxLTkYPHFjL8qexQdEJfe33GJDJc0OUksmfLuNuGNN2YiBtGD2NvSGN
XbnUwG4VrSVA9kqx5y1vDN+4YutEkuM2nLpoAXYdJ6i+8TLrtJPLPNWIbVMsHIoE
kjWOCkdKZzKf2BTB+axO+dCF6EKu7KhsIigze65eVLgiv3qlMg+7Z9DOcU70NrWr
DQ4PbvGA+Ixwv8+g0kdP/R3ylbs4hEmv/QXDOSo8TsZGiihWlSOib+gTbATNPKWC
REETXAGMs3/IanlixQkhLmKYBgKb8F8jirfv5+bUmg8rpl9IirOiJSF5HeFOkuVi
BvwigAZO6B2TRAr/jlqLDcX3iyzNz12fK713Lgp9HgyDZD+Rje/w6dZ0kJKfzExB
hWe60sdYbjR6+lUCpfZlz6VIikapXzvHYT29jTnJIiKtl05E91BuulsIUWkX6V8w
GRAnzgwyWjxtZ3HXZYW/PvI6cYyQLJLTG0TCAcyx6RMFwDpNEF2in+GI625YC0nS
dkI3g67bVmKCOzNaWj2PsyDHePKDWp70hxtCq47f74NKzhrdVfu5Ie2vXAosJdwK
ejpHRGU1GTZNkHl+CPTteAf2dx0RHbPInfWKXXSNOj3Lv0h4Pa5+OXiApha86cNK
rVTsvKUXuatmhT+iAHlbw1DirqLgW0pBORVtJ2dKaZZodgisAgggbnkkE4s7kIEq
CuSdGfuN0UTzerllEt4exMb8r9y+iSnHPfBF3Io4+aJqfevN/+Z5p4Ss7SVJsoFB
Z9zMLagSThI0fPZtu4Wm1icvXYzvZNoqEAFfrbGV6hsUdjMpONl8uwGD9t/JP2jw
AszVFNpjyjSVu2PnWQAFfbue59olur/QDND4pMtyx5MTChnfQT9OoS0OziB6nz9L
1haTpg+iCBqDC9uyIzZe5ZAG1V46tWWaPYNCIrjuiIsJP2+/nj97tDn8agBIkOjs
0oXUUlgZ8njoQANpB+OkALkNd5ieTCgQqtviAp4sRG5RR3OwOeMC1kSdJ+EeYFop
lXC7zjp2jHJ7/qMMNFlBhbP6GZzrzAxxcalr6rd+r8wU2UXK7ud+rhT3ZC3GZIRH
VUnLHhga7FjfmKlhzrMQg6o36fi7bwOp3K+tg7SlFyFuJ2fBCQYZW5txcu0stSvf
nL27p6m1fsJYd4/POIruQw0vFMA76N4hNOuJNEvqafe4cIvZTOcEX9HvgkvIZ56y
aXdOki6znhMWZyMtaVneLeJYZo0k2Q3rhNldkzp0D6zBhLn++kAEdfHg9IaijUm4
EUN2Aus1g38YTY3foQhBobhbLWqBq+nfdiGKZHgxE5WBNgDjxGQy0azFeLop2fbV
zHHNZwqHztRYzJIkjiJaVq7Y+cb/KCD6ZZVb1R3H5sGR4Ldkc5Ux9bGdjGrvKbKk
yUa8ax/EC88VIM4d3lLd1nnV2168Gz4NRzI/SXitQDqXYcB21+TdiHR3qpPM+xP7
RO5woy65WVN3wq0hZl/q99/i1XzY44xlmXvcToAhIZYLqcrwGksDAxFg44QisP/r
co6NUhgw6gekmStH5w1KhHTn7hwJyLtzHnZwgNT7rcrXw60tmB/D8IyoQdnG7rNV
ZBDgFeflTQ598Db+OZPiSqCV6R1OviB7fOxPj2AhyOo/40kE4LAzFjs9TFOrM+vN
OI5AfvMO896kFV25s4AS+ELRW7etPvhmWgfhPCovpGnjWKBw56LUU7ZJU0HROb2E
M6qT12/r9+t+/AOP0qXUs91KePH99YG53JmAO3vqENne+xjIc5tKLYSejJulMf2W
ukS/Cjf31Tv0PjSaquCG0vyanm7v5WWXgAeEiSzFdn0pVjBB6SbZDnAXUOLOqHX7
8K6dnpB68hOCRpoL1znxIhiCOIXDBuLBGOm08AU1Tp/Z02h3oMmmrZKIYW8eJW66
IDfYzOb9LVKw4Ofk8eXx+Ia/NwC39qArlvpLiW95fWCXtpsqpkDWr9vTZRhKeKcX
A5LT2Ty7zCtii5Hi8xHZ/iy4MNcedgzebyJDnPgBTnoCjOAZNDIGXhR65iKfvv23
sLZVOijFinVNJ/4YJtka5SLLIxU2Lhb+DnlrbcuDzOlFcRbJ2AcfvzfJdvwB+L2M
+40vtxMrmSSUrqk5rYZJQYAzmJsmcwnaUXj8JNNrOULKGzDkLfynoKpQQmvbhBKq
c+aFr0YmxDsg2QcGOU9Q4xkc+Nk+0sCwntywzCuFUX6G73Xn6LZ0gG6VvuNfe02J
Eide6dZfsgtntzdjny951U2tETa60dG8+tLm+zlC6Waz0DYEjQMblx6q8Whyb2hd
0wyaEpfoHjK0K97OA3XEr23MaFdFXBYAE+JYnOnpEq8dRj5EEVS2MWdLMzThpmie
n0SbFT8T435pgeCrVMTdkTilAe7t4FKpzVuIS40gdZu7H1DukfDLm0+sfw2e/p7d
fcdBSQyyzp8mXCG7wZVPT/+1H6b8f73KcgxPD5XDT4oUPCMvRH9pjfzx+rHjlTNP
+sCzIFmGCUqpSAEyJLyU2aDMrz+3Dx0tgeEqlHGlfgdZltcp7Km8YF2YQNjgB7b9
/IfPfID3VKP3S7SP7KRd7aaTjSHWZlPoiu1wBbpypO8nErJUzPTfTwOt66kvRf9N
7ZnvJbKjXntlFgfzR7uhfoon09WZh18WrsRWOVAlOZwGXWKTy1dJ3ql6T8+jXMTM
5uaq55TDniiBhO6rqQ4FUxc+Zmt/ip7SwiCuKcuAGItZyRNaCu0YK69izXhaq1td
+zYH2/ohy2tMCWqPb2wU2dUDwGgvrDCLNDeR7OOqLOzTfD7bEpiW793ahZUVPtRC
YoaRHyEaqDxOWey8f47i/4JdPuJSJq8gmk4vPFY0X0Aabs256ORzZWQry0qmqtCZ
vXSZe2x5huoHoX/JNmMKj6skKoGb+4MLYVK/ZHRaK3xzr6zYczUCScw0JKylQ+ce
haR37ibI5gaH9bqpfzGPFRm+yfR9PmUDNlAhJ2fDM7wz12ts6RR34vZhuR2OvBjs
HPBomBYzkMkAaVl+ZQzwbAdn50rUe16b7jIzgTe9Tgd1KOOvOQTveBLA/zhZvdwQ
XpFBdVvI3cXipFXvKyqZsSB3E7xjQKTknVUnlX+4h5HS8jsgIVMwpdX4xl/p7fLi
uK1xsh/Qu7m/+git97OuPcZ44BUywcOT1uCP3/2Hkc/NxS5ffsdFfOkQJk67gHuH
UNJ+UgMABl8flcXuMxrL1l4Erpzh2+LMXLJPQ+HeG1EbuNgesuFya1wPuhwoxuMV
vxmfHr+WaepJM8ZBXk8MZDLhUcfmy3XQH2C6H9t+POQ7Igfblbc7ZqDSXt0FJrct
7EIwBtdxtPdzE0kqwuM+10/MnC7vGW5LaeHkD0qIW55/rzWd2nQIhqX+Umvwh4Ja
CSt1SpkXPV2fBc5gz2/D+uA+RqEXaQxhVqdxPBwha9wdpnyu2Qrek3+VgTocGOHC
CYtI4rcxlRsIwORrVDall1t+im1gpJoixQVXlqXSoUALLNH6JOdd4qF10ilL+ivf
vv4ki/0gpjhj88FQaQ3KGcWrTAxUnR0u6/9YdZI1Z3t8dXzgsLpBSaffVRxFYfoc
+usB+RQaIvxqUaC3qZbqp40mZ7cxIYhHaCIW7VYzZYObFUGJEhMfWeHSKt158JsO
Jwp8KGOhq7oxWgwexj3m+Hvrw0ldIAI6GRucrb5F5gB2d4U9A+JTQkammEvQae0w
JMfJ3MzgCgxKeLMTYe5BawD1UhJKdKX53lj+U8zN9dzgGhBaUA6DsnzGXqs0aHYK
aLWtppliu6rGrVBdwINTfVNlrS+I3tLmb5MdLLdxeH1mDHLvpkMQTjfR7mjeAm5V
UuWEOHkN7NyF+MEhDddKi4A9A5HN/3R54wn4aULJmYlFkrhLR4KCSkm6VvztHH2J
xthcEHSP5dzYtsQRPZ61z48V5pKUBgvfRR06Loq/gk0rbJcRvXGMYio5Oze+bFCW
ZzK2b9Y+OexBo2vrJvIVDg0XJ53pjFLeXwIKE9ctwTJHArrbPock3NJTFgNzbQID
lco2sWyazx9E13C9ghGc9rtrJ+sWo+QYGGS2XSljfOnxRAMIvUm4+ENwa9r+xj2E
iQ2HMneNKztJ01bivJ/NxDi0mKOcg3nTxbEBS7GpwsXUQR3vpA5T6XqnZh1hucWj
sYE3QZhSqiM0CAir2GYwc87uY0I97U8xbh4GkfJVnlT3s0Y5d65EzVdLcgpQtskx
hBbCwivQjwOrwQd674ipkhB9HfD2KWiKq74cxD8j+1IqH6kdc1b3QOKLGaK5Wt9P
Lhcw0HEaEFn4jLgTyO2nfyhaXb5AlrN/A/VeZ6Ir8x4pr8O1kC/F9MgSPtaVJzr3
dIRGFpUhPsPBdZkkGlsh7iIFryEG+M5eBXhzF+9Dx9HFUkia5hB8Okf9f5FkVZrI
bTJkohPkzGdjKzSClo+ZR+UbkSCT3aAIO7v9fnZAtVXs3S3RahItI9xilysWmID6
BH43Cx/cChg3nwyHgSi60iARoMYgxI4Ry95jW+ep9K67TRK2tL7UGvkAUMt47Am6
bOf0maQ71dTLc5wUsbtpjhyJm++KQ4akfMVYQLx+s0RMqr1eu8IMJHG968GrSqUr
cQEFApclMGenNJsNYnoaOJqJfgxSPtJhqiw5COgv/qgcKajRDat9Dl0B594xj/FX
0eVRjLIkmWpoaAunO6jvCIMmVR8Lauqky+CneGML/Lns/DIM4aJplD9hzsOmhIkD
NNx79YBJ2DTdaKHTuu15bjdEiREVuhzJ0qtbJD67XcNF/W53+Si/QnGICs3K7wJ2
hKVIcqAvTXF9n8esVqouPcsiQp8he2W2JHdvbZGRXOoZMryZzqffYPax4ZSccPYm
Yl8hgEdvobsxiUvVI+zcDvSCmMpbPkDyKCZJhxu9XbTX2OKC95Qvl2a4tWqgwZSG
qBP3Fd9aYgjrhaP6Q1TJhVkqEqTXb7WD65Ai+bbXb73rpQ9o5ThgZPO9ClfH+MAJ
PtB8tFInD4OvugCXi+jWFNaYgq4Xt2Z1Q16ymupZQVEaSsc/6ZmMG/X1wzAPWmbV
ISNK/KMPbpu5lIuPaUdH3EczuLF/w0frU/D4Ix0zRt4md8HjLsOCW66tljnWxTvD
wEDcGWN2L3BUxGS40Xk6kTjaWnN3iArVmzRBt2X/yKZi933nDwnx6legu7r//Y0G
q1evvzzByfIkxG98qMqzY0lbsYRvpG97oUu9nW++0dYvEJk1J5EEGJcKGdFliCMv
Sfp9Sjjz8QaYJGTLnuotKqSsWRnOogOeGFLnbo3GCYY+LSGm/fpN92uYJafo2xcL
0eobMnDB/lNfZcViZTvz9rbiyBzvtiJWYXDuxPO2l0NWZat7eQWcg7fISV+khzET
LYxQVkba3yhUaKOmF1VO2wBlFO089D5iFjxPtWAAsQOM6b5b59YvxRLbd4t0moTZ
I/MIE951SM5RcQHrmc7GEoGbAtl3DyZigcMQEsVVNTHlcr27aN82rot0jLzzcBUl
LUlw5fISkQEQtS+ULL+7kMRXZONu5qseJyflM8squLMF8m7rBwrCejedm7dHGTrT
zwmJLB8jlEW6/y2A6YYj1xzOupYDej7Y1rGzDrjzvU8a9BO1FhP/uwPY1AYqoDuV
aj8h+CIu6f3OXKkaPYCPnhSdMjv7+VsIVLAypmvbIi0gHFxREn7fseWlVA+clyKZ
YaiW6slLV656HCi6G9dQ8b4FIHHLDSUZuAmRfLXrgHw9yN98OWI04CgYjCjNmlxF
FZTYaEblZYo+nF0eZdZbeRY3t0bk2lWLvPSVJpmaX6LMkfde2/QDHWE3lAdDAIgC
mjlJ2ZGwhBcyyzq0wwIh+uh6VjwZLqtJ4vDIAVd2I/hW8eIerR8TZAT2tz98Eu2p
/O0MEXQZgLdYZefFUurALGWsU58qPZ9UDUY5CA8cL3XqDoxbmuJRceRgFSzt/dcL
LeYAGIC4fZdyD/rRgOVrx03hGZQojt3isE0eTOEh9bALy2V3oSQ9/BdBUmUV/kqH
zmurKSepIYwY2252fpF/1nDeMZRbX6d+6Tb91bf7zFb1mnNQsO0PzsxMTsRjNI5B
5UwUIkU0H9pmZyADXqLA5P/1e104mbbWFuZHYtRnSYQ6HoEzY5kJtsNm+lu7Wj08
5JamHlIpA3MLZ2g9Qzny/qgSVLLTRQ4FrJy3QXJUcjwVRP3/QJ3rzzbpDU6Fyz/F
pGOtZWpAKb9gGuXRDKsMNt7pPnDKIstdFcPmisegTmcT9DFBnGDcEDaW+/XQf+gp
pBz252CMwoMoETIxXz2nGGxVa1XPa5LaZER1fDNoXK6YrPULD7/w5clQ/t+3tedj
Ef1owlxZxcFT6rm4zhI2iRBdx+uZwrJj5G5B++/RzNVumm8ooW2u4KBsrxSHJPQR
Lkj1GM+dXN/oi6wK0B2NeHruizeFPBuQWXG55FIed9rmTcIawRZrgbDMRPYqyk2w
SFkt8Rz811HBfZSONy9rrhrWjxdPyJ/r68xVV8VvavClKz/V1dfb7l0cxxaqJkBz
sV/3sag11UOgKRAQbGLqBQaWerI1SR/pltVQb1W8RMyTMEydGQdw5YP0EW0O9EOn
f4Hi8+L/o+wGsbY8L11HMt9LHQPR3MnbLiYBm/ifr4D8G8lTTDIDiIOBP2I+4UlX
/x9LAWi5A/J3F/9/GIj0HpkWLTOmyHKOYWZvLpA2dN77qFS+zPNFt9W93I42ouEx
BLtyCSsYonAnoEPXa1CRRyYM1TNIB0y5xuaPcj9jBg5cs3DGAuEfxvWz+rOGeIF+
7Fq/QzBoyqkJ7Awh3qWjyery0chHKv0hxrCkn9mVeMbCei0y0goatR3CdgNgjc29
WiTCWg0KVHR985mvszG0SCrzriEt0IQHG0aXV+Qv6yrvLdsWIzirxhnO3FZVVZkB
65TTyiHZwlcpb+m8TUFqSESRny54fTAmhg47q411+urOAjN3Yvbmf6z3LakDCxf6
O3pvQ4O0wRFccbUtqIdUuiNFHb3QHKRfBo7GtGYMP+3cCkCK3O1tj6WyIDAXgfNk
gKmocL3GBn4JU1EreySh4wFbrrH0FMu9U1yqdDwTk3EuXs98NkHuFDf5GQ5vdKql
HJ/Hl/srj4FVSQzlA4BTLKLOoIcHtT122fYyq2jTZ1CCFq+UNDEWsQq1ihNWBgDr
hjoZPsuFOvI48i5KWTwD7grUfhFlYmswjsstfCMp1HDyhbwZbc3uPD0n0f3AR6s0
WbrMawo7Md8nUVMKM/SFDlj5PcJDS5+MCEDXVd0B7taZHBX+HKkU15mi6+zklxQV
VVwvLgk7jNKF+sX4sYzhd0ULWLohrwGp1AHNbZ3hJA64zh55Byvr4+gIPA0p3PGz
walT5fQUuRCqxHOPWCMUaRkVIBO7oHk9DAGExQ7q6pxw7+xeWunTYjJ4qHEfyCtR
Dnhjai1h5ZFVh6/9QD3DjjxYQugZKWcq8SD3rK8qvHX5d68PlDAtyMWo92qailg6
z65ss4eTpRcx9ndP7EHo1dtH9g853hppYT/JNqBHhyJLoTdpE48Lo5lbpluU0jYn
A0lClf7NNoy9pgD77m16j/wtGcPrlgNUFV5DcmUrJwBZ9Z+yWYvv/ZrxqGC0y9lC
TkT4c1jMJtOMrFeRpW6XM237C/o4sEZCpOTlardwCngNAjBH9bCUcfb6OcsvHNqM
Fa5NUc9Pr2MUL9rTqjolHnH/q9Mz6QLOzWJHAXt8pEA8xTmsKtnUoc38h9SQ11ZF
9kAMKGlt/XKY6jqh+RzgKd7ZVhTuhqEQ+cY1qVvuPldwxAvfRggqqJDncNAiPEI1
I4h4pY7oTwDbNmb9QGmIUbO2KkUvdg4jpI1+eQKj4u9QIRZT0xsuDspG/32Iy2av
pQTrpSvl3J1yvBSOY3ZYr8gfIj6vHVAywLi+cb6pp8lw37JeyoR5BNEV3Gr8vydt
mBQVLYJy13SzxSNsiPsuJqZsxqrPGcpMkyOrJ1KCrpzMwPKFYW05M0x1joi/dtvl
7ciseyuSC3ERvoixCXBB9HmV+MftbV51tOAG+TX6LpGR4c0ZDqGqM3X4TFTmq9yD
rOqw3EtHMsSdi+o+YYLnjSvMZJ10ftbW8XW0P3sby31edo8clzYQzATBIOPmJona
FNLCeTd1DjgCLNYf0UwlBZylKuQZNVc4FFngqXQTP1HQf+2QKY/2u1MIGyyZDjlJ
E+0Va86DxiGzHqB3z+SXC0e2E8HJ7BZDriVcOLaN1UtNJw8O7nKnXQNLfzQhnO9U
CuaW52Yd+aaXRaaJ/XzXeDeOp3vljQPErFYXjsUlccedobqP4LIeZYDIRp5R3j7f
DVa4bOO54dSSW4JUGlTWzrrMOwLk/01Ot7mo0L15GP2XD1CHgt/xAW9FouuwWb2Y
XI5PY4Tnd8rG7ca1NrCOLUl3zI4gynYpu0sjlvye6T38sbFRZDs5zZEcasPeFZpY
W6mjOpBnaqKlT0qSuuYQ7s0uhw3LAA/lQbSzCC7wKujbrzLndySvcC8e6LF5WboT
YsneYRdr0kpxc52CKkkfrawpTLv7vBoD6MWueaZEqqqIssYcLdXs61tTwV+H3wXE
KfENJuhF6LDRk3BS3lihTTd1q6shMA5H+0IZILwGtciy5WHUW6uO+sRpOlVGjJa7
TPDb07cyvrbJly6GAgDnnHR0fP71tqaFgGkoZcNQ8jBRZIkktJwJnmim391Bzy2R
KDps2nuXoKYELsLQ2EhWOiIK0p1fLGfDhssSdRwOm9fdw43s+nwHwj/fYvicRUOp
HqZZgcgSjZxvgXaR4SdGgcN8KPeoTjlb7kt8tr5Ubzu5sP1YU0ss2CbfDP48BupO
1IwQMIZCuPEw1uXU5ETainMMUCsHmYRs6p42zT1JFvaKh9c/h7P/9tqiKFHJgtW1
99yFu1GuEbanbrmkrAfDGIWB402DUMfzTjW1WwX0aViGQywZuQa3e7vtLNHft3gU
YFyuu/3uIWzYtElDkBjVRjNokLZMQbB7wA1YWlbR8AAlfw4fBcaSwfngUaGhk6o7
s5MBLeYZV6LX+IsSuVAmqVGBgr46dO/MoHvZjjnCqxiCaaUSHhMehYxH4YZZF13B
D3wqstVLhM2OBhtuwxQosOXnJ4higIjowurTvGsT94pF/KG8u1P6W0sxxpfemmeZ
jyyqfxDJkRW8ye1LIMnRivMD7aos0lSQSTYF5Upbt35+FwveztRMLiPEPGCvC3Fb
cJ+pdRBrEtCZTsRz95FR/uDyKW9TZPhfgMmsrR/8T2wv1a6mSJXBNzIwsL5fqwyG
rXHWq37i5PoYmPKtDLwAzN/mh3M6TpU/Sl7rKTqtSu41YEUFBc5+wWsSG2xal2Qb
5J68wZ8oHV8cxyOxlKYl7qD1Mwlw9RfjWLdmejRY2oHsy6TTUoxHuQTi5XvEsg70
Gd/DJtVVjl1Td08N7h7G2bKbl5LHYL19dQRga9sSy7WTwwMCpyPWYdap8BoxiKzJ
12g9RL5MkaP1/KCO+X+3oXrLReTlqciT0KODt0bMzeHzTapO0IJ1EpiBwKHCXNz+
ugRRg9nVNRTTb6RLJVR6t/cpTIbxMq++AVGHOafs13guy8O0oVc5I8JvzniDoHZR
R+oJpuo79IzO8YGhkxoP5UM23M5t041ULKyajB+x/eHTActa62ThjL6u3YM3BJu1
f6jMle5oE6f9Qs5kIWeakCq4G7tiUWGgYGa4IdSKheB+ua1nnJV9+ZYjogpRuB1M
EoAgbTuBImOe2h1oBnoWeWTGPUy7ihnahw3LF52fJYeHy42SPSqGk9h93Q+PiNkX
pjCdRw66Xr/raUrQG+jFpyPEgeR7Dm3IJx0xbGpidSyP9s8Yp6abPPcqWj6QGTZn
+gY0sSd1wls7xbCovZjr0Nla9kqsRj4jyHkzrbGm1d/6h+gXY9vuveH7DTxOzolQ
+LoHkTre2ZC1/A0wgUuD1gzCeBP9vbFMBW5GHfgNlkWY/DC6QHuN01jXpEUUBgPw
GJympgpIqeMOAsasSli8uRDI/XjEsgGChzGn7Y3+BUUZc2qptlV1p4Oe9IO4q4OV
7QraDbLJ80zPkmzN2luGAp5xMz/do2/0ETg1lvsT/ZJpIGzZdmm2BipaoRtvK1Zh
L/FJzdAKoroz5Oszi+5o/XapsHVwlS5lw+uqPlua7uLYoUej0a8xs8gpdaMK/qDu
N0LTwtwucV+pQNYTyNjqrI3GpqNyBo5C1urNJYcKK1VhrA77olgiobqv0AHCUug2
bFQTKgaLGZCUyiKuklKMY80m/w8DPe6zZXoZivvxiEKQV1Sk84Or8k80LPFVKezx
bZrTj+Bmre49RDqWIlOIVHw3uyKIAXyA+a6zCF7QJvm/djuSDwbx5mlE96SUlu0M
PltURHlr9UimibZ8KVpQU77aIJ+VbayYFs1ulqj089ms25lzjg+ED6lQ4OGBj8Ya
1ScAg5gnkeWJPBywVhl5dduOwrPHoPMsVE0ijKDx6jDR0dBh0WXr4RAi2jHuuOTJ
przRdo0wFJYvX9SDW9RDctJf/vbJBWOdQb/ujAbfdz1tv6kCunRoNXPYYTrWJPew
TVMIioU2UFez2prvqCGy/H2K1zo8ab6mvelByH9wI+szwfFGrxZfrMVPLCswIDUF
1R27IwO+zXb1vnQ4fJ7pw6mdPsqlyHuaAE1erHpl9RZlTKeMmYn2+AnBXZZA3gLN
8IdIGbESICLPWP9eNPSrvGSGdoOgONCXOHTBRO9k9m0wUm0cQLTWZLNJJUCz7Leg
ZkKW9M0LrfdrcqtilWN4lCgTaGD4xv39CUj2ZSsI05wnQjVkB2Lq/X1nBrrcCQET
T8afszcqM3GjsHn3Eh4AyuWPuDY5S1jCQGC3/XmjC8VCMSsrBxr5YiuCLRY7Z9b7
d5nHhhSh3BEmwTSSLd+w98yfq916t4NJXAsjiClhB5cl170J/TfwVjzsMRxbuBoS
EqLbGUxGgyh/xPfWviLh9LRVxZXPGSQPdaFiyKWsWvaD6lpO1e0X5qticYqBnI1S
5eCwN2rk7DVrN7r3DNdzQqRAwoKZHEZLDVwldf0lahnu+qgnCaYC4kU/HfOw4DgU
XtRJ3e0OMC67tkJ5Hy51STxDrgxXyrBRCjdgHZR71G1FRXGOe53aXzY+yzKI9SyM
j6+evbSTheGgkgNyJRSoHS1PdQ/Tq5VrNFlm63z/G6bjCNp6Pz7itTbLpv+0TJpv
JFcJQdRE7qtFVbPCpIAOmh0Nsbn18V9wqIdVwvV4+32aXEZcy2NwUYvKMT99qZPY
RdCIEU5Ylo6klSWgAN8xghZ8lFrIDuHqyZhNEG4KTf+0YraPfZAICIYcCammjZHk
6Ox/Jtn2NXSKKWqI5oz+GUacP4VT+bBpdo+PA47PZaFnc7SANezmrXh7RGPrvPCA
1rHGnDALyZvfJ6G9v7mVhaFM1uE5vY9uoC6k4Ub81pwO5n3BzILGcJ2btr56lvBo
Nngf0BhvEXTSuqdtWLUupGT4V+tLAcVhksmEsn1dBz4tKtgWHDPiWkpv6DITOzGi
OgZQjgJ7w1FBu34c4KilCRYUVRFE8iCc0Qze3pVO1F4iut3aO7tWWr7/MhZBoZ4g
/Kpbrmznbl1TTYPt5uxErM1LZthGP62rEmjy6/bF1OOXqcEp1TX80ycN4KR648jf
h1gbRN4NeLUyhUKvEkO8Fs6OMNFhdDWcdfEcPP+GEwjiMeRdh7cQ6v7dzmO/+LXb
LcMPZll+SLwSB77zeQ127kaEHCyuNM7IeX+FMWokGM5hsYQUSxsV0SG5dkA3weSr
bf+bvoYL0up6pWsPC+HaycHI5b0ztn5xVQrUFlofeY1wvs/LjTiQPKhfj0jsxraK
xVsnprZtng6OFMYVXEyyCGVBYhMYYaVMVUMfaK9L+2elpkUHgp20av1xSRVvZXaO
aJ8EpReEfTIAp7O9QZD9TsIf8M/GxH1Tef4EN+fUvpF8npy+B7JWZTikQql8RMJx
5zW1OyEfoP5DCMV9NQi11eryeQT7cgACLGXibCzkn5VvRUoCzLFJCzmQESLfUTey
pj8NIZvWAUik8AhDW8jY1cDZ+Q22nR0oyMpNX0hpIGNWhNERPjCacs8zcHc9XwMo
oBv0vbbGpAH+bdDoTkYBdathuBE8MUR70HXHNzX15HomxIZ1+KoGYFbrpj7BCF5j
QLChXU537CIvVk3SLPK91QaxIUsJ1sJ8KAyK4ouEl9tvtv3eLqm2F7bg0byquiXE
qa4svTquXqC68FUQrIp//TDrsTdnqSKmIgClu6nVJtIZbVzxs+jyXg7WtpUD3OvP
mga91iaLBkUJqw/JD8PvfLnf2i8K0oY/wib39TH2WbNAHYP8ZTBMV99T5dYSv8vf
yFAdsx8BFvef8UWoV9msBn6Oknm9jmDSmh4j8G/GhjYqklFxzDdpFCi6XlqQxlro
HkpVnho7buldK4q7VXZXZmksdB8IyOR5r9+vdN4QIs+Zt6n6EicI5Ty2t+NB98T+
2+meYG8TZpT98POLpG/iEs0t1EKwX3Q04nAWV0g2i7FVXZ31mliNoIxTMF87igGo
O6PMnmWoRAZdhtNWXJ/gMAgDZ7PWj/xTP4HBxIqefWdytQcOB9Igz4V/UTYlEwhi
v2pLULqsJnkVVDE8HRfHx7pYQqcYJoV1ynP+hzLPgivJY0Ho0kxhmTT15V/WxuZG
UqQ0Bl67e71aJk6UlQj/yuqea7cfmursQvkEpjEFDiPikvxzMgoh09jVf7dgS+CP
u6HK7gTBZet4sUThUg9gexQOZp11s3IQcmm4DQ43z5jc91qSwRhmXKt+nSPv34QX
Fv6WBfwfT6/Obtkki6VXyn6nNQEXoEOGjxip11c3QLniTNC2ieGfQc9w4TwJvRCA
c8AyGUSBgX656JGhOzxvZr7h6xO21SYNHphl6D0v6AfVsxB8yw/WZcqAX7TV8aoG
c3NRWTxi6imMdO4Q0jrxg6toovkWZsqHER3X3pTXh/yDjF1Y6sYvplIzZa6r96qE
PyAqTCCqVa27y0kjh1dlM4Mq1cgMBMpn2911TbUKz0pKxfmvO6FgZWnu9qHQTwuB
Nwtqwc90IHwpZwKzdHEBmZ+3vMib7txFW2mIHXslk0/tUNTUNMO9bEvTMKwoNIe6
k8HMoTpAUHBFw5m7WAsfFZXtaCINeK3iLm74ChWZg9oxYxW7g1gh1zq7ryHl2jiA
hc/7OuF0uNXgBJOToYaxMQOyyT4dcR9icUS/IcL8HhmXxtN0yut4M76RqvoovqtE
vtJlLlJ/vYRJXfjG76XdAf0CWlIdgh/n3ONBbK0+VikBgZ7LTp4LXcGrSjgdH+Ni
w5kr4erhzxwSJgAXz8oLDQbxYgkVVQx09wiRCY7GSD/cMC7PCESlDrIqZ0Gae9Fr
EDVmM3FLl6Qyo40A/SOLm6GidSVGFRgjUol8xUQW/Hee5Y4UY/NwLdX5F0fH8GVJ
SY8nh2SKyzXNuKuCs1mM70fclDwU2kni/bVnkpkI5c+6kT2lMEjdVspp0mQAadJw
7pKVcc2bc6YhWq6eJl+NHKccgrkkIu6tFT1QhS6KKj+TqWHusWms2DRQjsrGalaA
bmopm5D58DDmEjtDRqjZ4s032amVZovhsZEDAdr6dKEzyv8rrnwty+6IeDER5R7i
kMsMyuE3lDfWTSRl+kyzt81AT4dVQWTmpLZCBY3vs2vTpq8Hbqt3c8h0skNMOubN
l7ZW/+psrBRaTPPeY5y1kvDN4vq/5iYFUkBhnyWsXSSHDa8hgrxxVP5KS29uoSZf
txIxka1uBzOeUZ/CqN7ZEdIVxHw+0v+9yHLP4MrEKDnoCkcdDUTaXxjpPlxTMmtf
xCa40Aae/V1lDwiGIgFw8D4d5AthSS2zmMUTPOp3Avx1PmOrSYoCFJztymoSiRak
OWo6P9IZBBQx1E8hjiwsbZMUhv/V+IM2jMgcv5YG6nYYKwatt7gqXU2wXT6qdk7F
JfI0SLt7ieRg/ZAwcr0ZK259MTk+f0q+UbUvdcrK99CyjIUfjuvTzEJNmwTcrWIX
CPbG4lOo7fCasi9xCxpxQxfHUG82SHnpUY+OeEV/R34BLG/caLKtiBVt0I5D7mVv
Z0U978hsmC8a8292iQ+i9nbiCuce2F9pJgE5ZQ+zJwQQ019WxGqCK0520FSXT59b
apHDrcij7O1LXb0S0QNY9oY/1GlTkXvtIlqr0eJEDXsrSSnbojhowLvzFj9BUntl
O4dOdZgMCxdl6EgkOaOa/0VDLmVP142fUDwSU6WgSzXbr+iABr0vo2hZuTOX/UD2
0Fpnjd9n5RdcakMOToyTarrTI5vX1R13j9UpthAqn+GvYRCA48AY0YyU9VkvaM/V
Db53KgAioRI70SUD0yszq9BuuuPCRaEIakmteH8Dfx1PuvFxp2o7x4ZeV+obnVoH
2480cgjTpoy61mJxPdZXkmbYgRlN69kZo6pGOx5Z1H7hhhRmV+KjbDiZMAxlsN3P
Pws1e3BdK7hJiocM+Z9yPg2Px5zJwYGt4VqgAVTliaoDzcvOsaeiBfVyKyv9Z3ol
5jaGu5/fSB5EqgX9TlfPMb5JDvP6keaIk1AhSa4ObjpN5mNU+w3VqB+crF08qEUO
o3zwfneZeVaJv3y8wbfAQU2leFIENCVg4SM78rFOCcDd2KiOBolXfuIaxlHIFXVI
iD7I/4R3ww/34XWKO+rRJzsPDA4wGC03kb8VBMPzTC4JQAaRGOSk3BLGOeVH3F3F
Iq14v1f2ZUEjF7PgmLRyTIBi18rRy9YVl6j+5/6NrPQthH5imCmPJS1OHtzGgfUl
ovSDckOk6uv7CAOaau5xFn8f9C1Hvgw16tv9t9Uj2HyQgCJmmbCBKfzPGzdr5xt3
cT+zBaiBUCtJLwrUqbWIsKeB/8IRB1iOVxELoqwsWldsr9idMR8WzEF6YxAMdbCp
ICoIgytycoe+Vmke1eWwznsuzEiCuaIjekQF37GLcXKLimmteAsWO1xF7sukwU+l
rKuq67d1PTGqrMAsgJtcGq8G/AaLD7Fl+c3ixi9Lf8yl9ZA+MzUZ8Y2xkehtOhJE
5bcfkYnkHL1gaqSdBWTKAQbJkJlpwO87ifug6KN2b/AF26IW+AEwpmEbxmNrM2Wc
zK2/5lbOzBZmYP1PEQJI4q+U5duGt4z9LN5p7EN4VcQKh//8QX3q+SjrCeIjF0Jv
OHg1WYQ9ctopEVq8bwgt4fOv7WNasEDONzmUeID+xp6TNP6I45iRQ6QCTV2WcUHd
QzoVJltjyzxkiT4wjFzy0ifBi0uE/rAyhWV2W7epaJ4ClYFMeuKv8pzP/ELm7zw7
0HpTe7OU7GLHHTDdyACMVs1zIX//Z6NI2PENSO0/hHvtRKc5yoAoZDrUXZPf3Tm2
Af4LoBBnYAkA//0M40o+39qzar/pST2tG04S9IZmccn7ZowG+CxCuNY7JbzLvcv4
/GMEI23IkK//lbQ2vIer0lkmqPc0o7auYfcjcAlC2WDmsY4p/fqYqhGgWwOCkV+i
apH7ktXPylzsKAgOkZutfLScWTZ+ZHS5yeDa/uCX/tZbiSH4LNv8/6jZ68qDbKBr
ZHbx5J56Xqiw1A7kTog5p6V+g9r/wS7hevq45cXfnB7hwxVdSJUOcpUKrVPy5YUn
wG3KPA5N4PqBVeoBB8TS0y4N8nwvkOzR1aJR7CISsZ1Bf5BCoZfgiD9SrdqyVkaK
uDbJ9ZEKEdDZndJQc0uRW4vxd4c5mMXH9DEf4nTIGovLUljVHxS1myvWHROde6X1
aFB1U3MUi99c5b0znK0gdvUza01uxhYSM3wUO2I4uwzqz3iMYcR4JsNx2hZUCxdo
y2uXlRDDCoDNYE9jEWu/ak7bn++dye3Nsdnptng5JEUBdz/VyZZuEwQctf1vzGyq
raNimjamRxtZjhSo/BtWkUnlTFmHjmW1uG1vtEhZpyYooeVbZFFHa2pK19fc6Knf
NIthhNBOsL0YThHk69DBlTAUl/99s1RSuWOrSimMyWlDzkSMFrYWVZOROD4gmeDh
LiY0E+cKHw0nYJxgDQBigPjtTOlIW74Whi0eynbxrhxMeZ71XEzIShtWr2E2+xJy
AcqsaBt3xXe7nUW511mbIiykW+A+564hFBImQo7Y9iL6RxcxkQILOci13Ptq2PaM
LoCuEl3uC1Dx4k3WPrgFkwrOd+UlR0DpyPKG+MblRYqDR7ayKaBczMgg1godqgYc
dHoVN+2FK8jNFl8I5SIHV+a3pXjWFFmgvjFy5GduENjJMz356N2rrBpOyRJA0zXf
HUHWk0eY3rP5ir6ZY35ahDbHiqo/oZ0/1peEnb1z25pPljzp7XGIrzbe6eJp2u9d
FGPgSU6pY/bJcCu55fe2wXUhI/CuslFGWbk8txq0NyLlAbep9BdVAuEZAsiZiKlQ
GqED1fKINMlPvZyERGUKBVaTehMJ4BgEzizw2cr/T/sHcFWdpKJR5Ljn2H6MnzUt
k28SFOd3po32XEeu5ZxhdtTry9d5Tk3ZuAZCZEMtExBg0s3kkjWLo8Lh3bKzC+1C
0gDW1FUOOlwcgpAg2cJDlvLbtj5wSfw70zIHHRgPJ0i7eXFXJcNsQctxDXGi6HVv
bFv5pkqfQbJpBBDTHz7eRinZ3+bRDWzgi/uSFVf8mLDIUd3+Ehe4fo6yzmI6jza6
B0lQ6YZNideTlgdP2csyIuUJTjAkaWo0dfIUAv2HvX3jevVMxxYOiILWJoB6SIGZ
HLUZJFRJJvzJ3wInu2k9PDq4fd4Z+a+iw+0xGwvf3Tdp+Mv/soAysKR6Qkj3l0q7
P4HBJ7N2xPhCcmgpFftsHWXZ3UjbgAYPW+aek3nWyTM8eMtCdkQ6R1OdSVrwXTYn
JCG4i3Fwq9NR47wYxEgzVcslU8grn5VjW9NwpvUkHM6hkxqaoTbZlSEAgDyX6HUw
Ae+T+bWL6C4yUSrgrLm7ukidOGgx6vj4ukUMpfJFcIhBTMPDByfuT24VTzuBvSGG
FWP4KiAcextU/oh5OJPASpt2R0ukHuCZY+0hoJzRqgii3gCAzU24uWZVMnQUFnQD
87wfjmhixXblLR3b2jNr8AVCO7V6k3PYotM5RYyZ7San0NQPy2T4QjO/F4m47pmc
KN9WKKimn4TasaTV+geEXt7kKJNhwZnu8aZrctxmyGk/D+WgT1te8gHeU9LxgV/K
EwwCB8Av6GTULTdKs6tFNdc9ph18mC0OLSb6DvCrGjFoWi7ptg+lpTe6bKH0ujdJ
fftYwNZip50jMQAmyklu5urbUX/0qypF6M8HrE+HiCWnrByry2rpwzY0/JCaSEDw
0IZHWlQfu0+qiydtCU5383wCDz4P3P3MgC5nMrNolPEg39iQeXDRcEiMoYQsZFzL
WwJXUNn6fybK/W/AtziPRWd4cxjQjTj4ZKylePYvldTZxtIK2E1fZECmn2+jdbQQ
cV+d8GAMD9/OZx93LF4phRWecM7ahYzE2P3A5y8Yj7DlcIg9ni/Dnw8whx86HwG2
IGJ9YQv5jnsS330B7DVwXjd2+lCyVkCJM5fjA+kiCsBf3nPoD6xM609Wtoen13KM
PVHa6UmQZi+eg8YlRuerjR2u0g5YImO1hT4gk7jfr2/9UgvU4+b5DM/pzlACKUkD
Xqn2Rbt0t3UaW+DZyw6pvbaTCQ1t58BTaoUxtoSGmtmldGYeqs9awMjdF6WK+CnY
m5ZcCaUo2PzvWPDHZBUC5QF6M2NRPKYa4Ez+vWpETIf+5WHbPjkinjQ4KZBHpRWC
BbmsgmMwr13jrle2fDzY+3rKzjzeO8H5DxVugqR4RDbh8+0CK7LidSV4KJo0FtrB
J00VJDmg6UwkeGgaemF7KtflVGoU6Rc64LyuCYErnpFclLwhqymkhHJMdFMRaS67
0XbC/BJ+/vKb45XhSN5U8WZog+JhelXPJzib3RzI16qDwctSfWwMqcYEibWFssXm
JJbzWQcAvT6DxfNIzK2XkAn1sv3s6QRtWZa61BG+Yw3mFYMsZsQecm9FyW673IT8
GZUWWOlwFJ/xPdzoMOorqlcRevewL4Enau/aTJoUdsGsibLs8AaNHj0/k3AqVuKv
ZC2GH/TzedAgvtAYV3aOzS7kSmAsfUQJJHGJUy69Jma0uEzRDpm+v2dRkrZx/XeQ
tAKGcsnYHTlOsmprAWkr5TcHoYKs7dTI42IYuxWhtP7hfSq+Xn5b3CdLOQdfTmyP
Kf+hufBGnFfH3P0jB4HmBuPd+N7D53K8R2dP3VgKiCh31ApBcfFzjOzs3bt30O3R
dTU+R2XpBodDxhYsRGe6vZmTwZ18MDxmCXbYb9v5SYE3FzN9jYCFfVXwLTlRojUR
51EWHryMHLqes3VsySOMissQE/gC0MiL9Kbb7nEbl32RZ2fNs7TJA4NLVjKFvN2v
zW/T47Oz4ZJ+tdUEMAT0ZrPLCPumj+BRbn3Qiedj0ooC2YkcMLtWpI/gkL34242G
VhrFTidqzXY41E9WNvdbo0yI17whyCXT6sJGiP64Yzk6f8BFF4o16lLBIke+/oOn
dM/CJ5FL0p6OVUffz4I7FKxfOYEUWJ5G4DcgmyBHvia863kWI4x3cwVdxHepLW6c
XxyaaBgEytwZ2RnirLHR8x7Xh3lcrh1WEUwKyRSjuBvRLoHOeRxNGUczUqJZsagP
cSs8TxIjwFU8uUGHmiyBFqQj8dIC/UmcLH7s/4JPI+wo1lAKAFO1wPHVbRR0nIwP
I/R8fotIk0sstPoUdF6f09yuBYvBLgXZ69xw9nrnlIu2ygvlEy6KW3sfhdFJ4K/5
E69l8U1l/WDqAKAbX3W6IqlgE0rdTF3g1ZiA4/w2Xn85ukiDlWKgjVdonH8mAxJR
zYqWPAMjRMiwwbsoFP1YMKjI19by6RRukUvQ4gVPTLr2ExLzI8C8bGSfgo6N1SQ8
bAHNHghjDC3ByLaMWjAOmS93GUc+ovR222OSmZK/RrLNgeQnTE++rZmfCR9/zfZM
qbfZrFctTv+Jg6hYIVGTgC7z3+4iJANoK+jjeOuDac9jHZYTz57ek+2x0Z2eysoJ
KBqcTmWAn6kX776bbyyCVp7/09VNfp6IqCsH+5vW9m974OzsSdX5xOHxmjzPydl+
iH4wiTmBZ1lmOSvzw1SAREF0Dzhg5e07aE7QpHORBxvBydnknC564x4RBnfVhfTP
EnRsFcCrtvU+MdboeZCDuuvgpHSrNHWQMakZXvV+plILMX5T+j/vsbfq8ciYmi3/
2V+Wl1/3x/mpeWGjZD5usM2zj6C3DiRXijnp9eVq9dWmC/TqEVLczb+EzOD/4vCc
kadIn2os67pIW4ctnSfcku8RwWiXPJCHHbqntsT1AhL/1OwOA7//r/tzk+9ErTWO
t3SkiwyJPH2K8kmtrksZandLMZVlnA8cEzqZbN5FyxoqQnKanoRPfIjolv4txYv2
dPFhCwH3LYpTJh26xncIdzG0GK+NyxwxDMGIwC1/fCMsW8vOuYIBN58vFcjJ1Oo+
DhgJrKLWiRLO6XKxYI1+k4HqxHpKbG/0HeIwYSGG2vJ9ZWh5MzyQ4fXcd/817Pu+
SOW0WMW+phtZZNGNqOcIUSDhTdM6cILAOvlvT8U5ZONLK5PeF8SLL6SPogCxutuz
GxgjbCiV9rh5NK3Hb4EWzI2Xm80J5VSjIDveIrlJowD4im6T5lUD7qo2wfmoz16M
kpsxgKqtPBI3owjV4TV6DEcdE8AUTasR3ZGsBNFvSw92hh04idakgQ7m1Xh5f8r/
zAtVAW0akyvu+Y7/tVa14C5xLEG/de3NEijOp1j07gV4zGGYpA4daDzVCr1n2/7r
6xcoM3G8ZJivWzRlDAY7ZuwACj8ka3Jg5Nme7pNtUrpO8Nryx91KmhytbsZJd6W2
JmSB63N2O170yvYK04CYYVna2imAUjVY9WTo7bTEz/cVVfyZ/SvUvJiWkvkZ1tDe
MKOHvl3WC+1OmAt5yyijJdZCeHE8Qn/hABy9wqFOfGljkd56FOMhbum7ogryZaUJ
obyTLm9w0g0VhBo53hS8zpLloMpu6BvRFA6MuLzYLGppvhP/k46z+eGAXpDyAvNy
ixCKfa1IALLC1cD2eWUQbZrvHx8NMxbG0yR/pkBp8pHA4IwVyeFFBbyJZmPdk+Ag
GZI0gWktviYSEfgp6tgj7FvcZIWMc5aOydEmPTr3IqeSVg9vpBnX0qfs+0HuHyRQ
yph17yAkDXZajx0x0zmrwiSDNgelH0FJYnv3JOH4uBXAR0doDFwf9Mk2SbY9gP27
hxXKWPboakCwlTT0SoA5Kic+iMC+/xUod13YatAkwX4DxViJzqZPBF4PHWc6N42C
YEv2uupvm4UhOdRGz7VEMrNDLoGmU98HTT8Cz5D7H9ej/SIdSZ1zm5u99Bw+J+F6
PJxl13Ic8wEa9N8TVNFm8k+15P5xc0p/Wg7Nbu12CEeQvBB4wVNwUEOAxSGqqVyX
4WQMVwG/YCww8VloMR+Sw4psaoYh0j0saaCrKKBe/j0x64HxK3C8NcEg3WC1Q8KA
u4qf8zdCTT+qnoWHuizRY0+M+WIQOJ2WZnWrMpv6eQ7eYU0Lx/cP+0lLgsHofXFZ
WGVzrs99gH/JwcCTLBh4cwazFrRXDcWn5HOgLZsBQejceylBTtLTyJtWU36O89i2
yRCePp1F9EPmBfwNxrmkFP7nri9AXqMVLhPwlRUCLrrldE+RmfiO+YgR7/37RQgc
iubNoVJvFVndhAwOwtXXw70n9gjDPttT/kWAMHd8CsmqNtN1UVMKJHxp/GOry6xe
QYhiiHUZQZ2mO6sZEQ2HLYw+qX1osySAd4rAlZqh20KmFM7N7oyfrC3EJpk/dS6f
0rO3U18CvSai+SBRv7lfPpW3Zr2jvVXxT0A1eWUXzH6SFSJ2MR9hAqkyw3TyCbyS
RGkiWO23LfmejaczSEJhkOV5ANikYmFrUdhV977EcoDhWXOw6lwzFmKmtStSndnp
DxnQ1cQHmQLBdeMwxaxjV9o4a6AupaTIwjT7wErc4I9p/9FXTje/rjxzQoL1BIhL
2KFp/NJ1yE3n5DajUKmMYlB3ZYmFOhhFLKY3O80hlBijdlpxpDTaWfHxBVym3i1H
pLwxm4GDtVGjfktVTJuYvMzf3wvP9Y3vpVhOSnKZp0d5qtr2oiMTT8XGD0RUWn3Q
pQVuzhXp9HZ234eNpCsEOiGjobNQiBEJIPKvJ0uTZ8UR+TL9Xyo3dvDBNndGxTz+
7DFnuiGiA50pgKuXvKxTEt2WJBLwbeDZf1L5bW0jVM1UnPr4U2oNEQTB7WHTvQKe
rFWDLkhVhuDhkuTAK01kMWSqZoAwiUZMkypxQPEgk1LLSS/d9981RTegCf5IIRzL
E/eLzXKWeo1VezOVbHrpzTzmgKSjvBkmSyOA6F/5KRtlB2o98tlaoa3pEZ9pUZ/V
NAHYRf2oKa0YmBHYIAojNVBZxyDHadD5sXzoxwf5czs41MoJFc+4D+B33umy7an2
qvLLpx3+3CwBA285xMz/dgNmwYNI3s1Pqz6rOkUSfXKApmLr/TufqvD6HDGIo43h
LpjbvCE85dfZ1pXDcK3GMiFYsEzE4FUXQUS8jUksebSonwmBS3iOHjnH4oLnLq6N
Q9l30pHZJD2qfDEMuMf+Yxw6cUckJ+jKQg4Iiar0XlV3s83EwoyNC1ah5zXsnV5X
QFORJVEKGs9aYHsxCX3L4CAQld+wtAiyKXYvndUBjdWrps9MQDo+ObYD3Rm9q77I
IaClptRloyIXbye+fNu430fJvdB48XIJngUCkXOqLtHir5uPAgeH3JPv2aYvw5CE
mCzG/YonVGrwRCF+q6shc7y0yHfyimBK8Sung3sQoGl8VgblKzJHzQA5enkL/YJM
cn/oxqqE0MlxZjAcTE7yypKU7w7zoMb6hbLBjq90rTqZ4gHYlBeJ0xQ3BqWBQcXC
bpqU5tQxam1N3EVZzvJtxsq0fX4/ZYggxhl5ohh8A3lAM6IFQxK5fnEqRqNgV7lQ
1zdyu/bITY6e/0e8eLCXbqrib0KF06ZUqgj4iMciMEwyAPTVyHWXRAB6FUIj1qLA
tX5WoL0bybXloZr7YFuSLYgIilH1PJaS4aVbrsk1Ni8WiffkFhhiHP53TIzgd29v
QIlPFaoAKOjcZ/GZhxd1Cyftf9Fvv6AbA00L/T3hL6wpSoC249PIj23hHePtAL+a
PtNIAKVf/6ggTysKH/DYpiQ1zANgP2SXrO4b93TSUflJxfAa8drUXXX+rKLZNCW4
z4MijwnzWtyKYSWnhvm0QGV5lmIPVH2ltxcWvd5fCnDnY2UpRHKQoPwc+bWY8Z+B
tqqPkvLB3yF5NGSOs5vdYGPo8CJwLCLsekXjxaMcUMpdpHZEUilnvI1SIGU/KPMM
dCWNT15HNDwieuDVVGyTVtOm+jNjp3atGNSMqONR4ebOP0dDjpNaui7tKAd78JXT
yy2f6S88FotIN8CGAsF1bne1HxeyzYsxb1CuaPx3HThZRwwmYqmOTnpRTiaUQvrn
EWGAemkIQQ79rg6DNV24TXg5Nz0Gc56IYVIqmKY70t+RFMqvYXDRnTahoJygAUJn
W+TWv7lGz63kaa3Xjo+d5gFwtV0tcaOEaeHN/OdPV6jlOzCrBpSc/BSBwrpeUI+U
mgehA0RNytkDPBvJe60tnNpYQ1TH86WATyTZ9ZM8SD/IWV5sSYH7UezB7Aam0b00
MMujyRNvpDctJ3uzuhhwGjA45CgfgdLBGB9NpyWwRbqBpFHL1BbmXpJtStfg/fi8
D7RpuWb8A4RQ4bAJLmaWd/CXQZa6nXlzyK1jsQqRhcN+LiKjJsYQsECgEqpHBmbj
GPi0bDitnJM3+36qnG9Sg9TMEPoJEYJSjbR5ws1MED+TES9UNojiJ9ICkeWurdUL
mxUrP4SMav7a1xyq8IXOmxBH/r4wpbBr9D1WZSP4GkB40VYSN4H6VhlAEQ4sUzKR
edPL/0JxLNkswP7ZMfG4ECD8VzJbWsplHsP2ZfBH0eexYmbHaIQWOsxng0R6RSXs
rBNFl+LnXHr3WVwaaqgozGd7nOQKJ5CxpTfAm8t6tKbECK49L2Vju2F24Qztcv/q
Vd27yabDlR/HQDJjk74QcrwYbvpqwVE115SASsIld3W5yXpccd1vuxm0Ibd0H3IS
/GC0Rjy9wJflOTC4vrHauK0M4z0dbXBR/NINLdUKtTZTXOHzuBjsBIk9vYXNZOfZ
agoUJWu3s1aWBc4sEZMRlq9T9YvWiMWrLtPoix10CiwzV/FOjb77RvSK3ZAWL2BP
bNSe01uL9Y4l9QJ8yzIQdJHLitZQZ01u2SBp+qKwnRDRNRH0cn0FzSfxabBZqX83
F6MIVSf7dSCtTxJ2gT9OhM7nxO4rbWG7vaj41MrNQCj7+ItTLbD/AyNczutOxO0Z
epuN716Tf+ZsqRsQVEnOc5iet2k591lKtl4t7jjrFOOZOjbCwwKs5+EuLEf8weLs
A7jWHAhrts60AM9oBiS1UHBVC7683WLwW44UinD4HTLAp8V4r46cCV7zfaQMa3Jr
Pql9ZEfwuspTvDJipw3ELsYdQ7VBdadRdsjKN4i/Ip1NOClOLtVLApUEiM+D769d
FsQm6HIyen/KAcfExCUMmgj+PzOCGHMWGSULkD7bxEXSUBGu3MoMvmBkNYk+Jw0H
Xgdle+4fBD2N5DX95hpaTr0XJCLE5dcOjvj4PdLamI2VJVIXp7f1PK33ipqOqboD
7MXi6W85P3pHlgTyTVdhWI1E7ts2pPULod16KEFn3pwfu9xrspCAb1sh1zJHKjaQ
TTagdoGPfKL4LVOyuwwenZj54TcqtVAx7XHamsxjXoRPVbBwOhM1Y68dVFKFv+uI
pWPOVSS4dvJqk6wcYOHqPNVhwni9SM6OG23D/O+BaNgnNEje3Eo5Flg0031onbfx
Wo4efb0qgAePkcE5xLsysWiqsnHSY5/WUmRfmLMzhOCy79DR6MXBFSITWI+GX1oW
snCMoiWxX5pJINeyMhBFchpFCyRU9LK/ZO2I+KJz2VoFIHocFJ9wLMcp9oO5Wbv9
uNmQXEEtf0Gy7XdS+IOEQh5d7LYRNd9jrn/QuEqFMq4MoQJBSv0jrWj6sssAvO3V
6hoFJtA3iHkfh2YqVkxg6dbKHDsYq+1wEJoPHb5zMFOwrRNz0YsSxf2ciktkHzTZ
9d1i7AnSNyCzV2e4JcvVOUTV1FwtUSOZG6ZUGiH7kSdCM3wQL2v+626i5NViZXzX
z6j/bOEHaD2qB/C9MACIQvRNvBl/CbOnHStm3Oy5l5q+k6BLs7p8JDd996PpdlkJ
o4yrSYBJs2w8Q4aPpjOBxLBjZFX5g0A9RLPEOEwet4fEeDe04dhcAq4UNzzpj7aH
0t8FNb1MPHisXw5m83evPmSqnkyTklHe4uAeMRVIM8YZ1kIzFx1CJtxvW0iVn6i2
2B9Iv3amUMwuVWKGulgdwAoeyujbmXYGQDZG+T3eynCbzhYkZuFDCks+GcU7mog7
hvcQPPRI6zR7Yi8B7yO8jILZmfPdFyNQQyYLA8McDC14lRfEy801xekEU3hG/FuC
2JMMDC9C7wVn7RvT0MnDxMCjLpVqq65Lyi8onolLqF4qW1nM8k3xo20ZjYkjBIq0
MG+buWnRdG0dKUrKjqfguMTTXIr2Saf83wd31E9ivjl+JKAPXbAt3tpoVcCKjy1E
syWeaceB6IyRxR50Oi+Jyd9O76y+57Z1UscfvOIb3/uA2UES/eWrUkojA1+BYM4c
caa5CSX8Gqkgu3IHd+XWACANaZQvzBobZt9VIA29t0UzfxGWgc3TUsM8IimlsVRS
t19gcZemKU3N66Ao/gyUISGhYydTbVOymshwej8EPOouNCBe2lr/B/FKv6W3BSo4
HC31MWZ1TLVe/p07vVJgmRbt+QJGWsgKK2Uc9jue43D1r8FXvz/YtQ/AYhXCJTU2
AZbpS1SeRRisk4qt8rNazmD8xk+t1HyZq1+ddntVr4tx6kNX7muPV5ZqBNnh13Dd
wHCXgtMpE0VmzIqF1kN4TFab2PaJ4VagJaUQziGgzC1hxWZ5LG7GJzJVpIj4ZYsA
VJSvW1bgr2cIzYtimivQuk6U5yP5BAxBbwdQvL1+MNgtc9BlOPvx/l/jX1CyC8em
Q9mLyeRaWnYNiI1Z6kmLAUgVwsVUMvPxwcgLK6W6OC2L8xLfo6u87iXr1JRfwumh
ha3RmKNV3ZEPGdCa+SuSFKZB0451ZqHa8AZ8+jPstboes7m5YEgj7XDl2c9iCXK3
4PffqAtQa8k2UMCf4nKWM3+dzgNCdDx7J1cDa8Ktn3j/ziNzzdsJUk9cpWkO+uTB
8puFp+nx1F9hFzutfmI8pNkRa+5WqIjzmlbQJYRCju0Tc0pJlMv1Oxhi23H9Cjo3
+mcoT6nHdaZyoCG/xWTXFezGHWoDE4nSmrR7QhPxCzQFbFQwDnJC2D4slXy5Oz3l
IAkIZrJ4iPiNVgyLUueVG7C0uukQVskao5LyfzPiW6hjBxOQFuNVbqdW5wkKePpk
pIaldHu/2rBxyP/dU43Ih6qz3aBUMpNVfHkWRyCAhyBT3UrCeGO21AUYMJDxHO7u
Vt22Xc0nJjv/LaMna1SqEOz2hypSRSBB7tc+oJEZkzsJdyJzhNrTiWqTUsoxLEe/
G3vdNEowcOqpcTujPE+pqqRnUQEw+ysL4oDF+wXQswweiKmNhY2sZEynlyWN3pwj
HncrqLt52zP4Gjqit+LEEP86bN0h0w3O2BBtkjR+Edz2xwM3CM2/sfILOuZWuzN8
PvFrRMhYuFb5eOTntp1xRppCkHPnZDdZHRBRyLRVgCRK1Gb2PfbGcEuOBqkLKHe0
36j55IC4LpjqnxKV6g23Pcv8Y2QcMYt4en5E5OqmPdZdzWORpZmPlYea6d+m0yPa
LUSUeV7saE9XlaYC1DeKuJoqIvFAafAX2mW5f09OtaTKGFnwCfukRRgXmpA6TA/d
6CtWwZ9O3eSQyagoYmqSqB7uWdcGTfrR8kIvz/4SrVrrnQN3WqJ9vCWZ5PUaxuN4
08BOBHTGDnUaXexFBqEmSP8IuZeKa6bWpC05kgGdbG7uMShqzQjeTIai3PohPJZs
DRddES42Bm8j/93r5KPCeyh3tSd6RlegLqKCmcYdIn6ZmvgrasyLCE6l5rOCrq0j
WhvsWQn6sv+llaJK/vxSXguU6iNi2gJX3EKyBrDOKowcoCkKlzf04U38A5GM4Ven
GpmrsPPODgtuts0pM8soGgEsVBi1yX5kx9vSc+4lpYMwNe/nCwn0S8rbz328KjIu
jebqkmK9TuHb47OI6+0zYzo5Mh8HRms1Lfr8csHT8ZQq0Pd9DttG8IN8Wy1uc1dD
HzGvfwAAPsR9lz5n7lDr0+kFlPHbX6XOGPIO6WPB2ev6mBhTx3ZjzNkHYhgQcVZR
vBkk8QBfBulvweFR9Ya6FU8TRd7/hw2zUCTpDCAet2pz9S3yY1p7RxiPEmaGv8VU
aFHulVXMTxv9BsUMuS6NAuLjXnF/9OQ+eP0oBfi88ajndHeYWR0adfaPkZKPaoxd
kg3QJF10BgG11OyUNRGCq75+FfNpz/sw2qfNYysX0xbbyP5C2XzCHnjPfL8PdDRG
4ZRGdDvVEzHipfU8jjGUGRERdSzB/WaxFvcboZLJQ80ZFb2nTjRp/xp4ZhX8/jYp
gZHpNBPIP9+ydIUQJh0Tgb8zJyD8/dB5hecGnuCLy+9zTY+/nUmsBmoQvqmEn7tG
Yk0LDpCSXyU6Q/fdVsTOEW1Kcqm2AeqSrQncObTsHth7CmGcbEBJFCg80Zda7DM2
sfLQMQnDWKauZapaMXY32NUZ0o5zhGT6gcV4fMvvW9UWgjZadCwfCzgO6yQjWsLU
6FGSK93XP+WRkjX3Lqn0rBrUq9JI6lNJtRGlNCb1xIQ36FyeTKotJl3eKfqcwNBS
p4PEryQYWz+Amh+FdjgPkLhtqDg3xTGVkh0HtKmEHBsRrfywtVAstGsoIvKHVyAC
qrVGe105MbfvLy6Gvv5nVttGpmBfwRFN1jRPSKSPJ0ZvvG71PNFukbHs+OaCROSx
oMQZ0crTcFuLE9o1MQdUAxqkp/FC7vJqSj/WBYdsjvzptC/SpOlOtJcgDGtLZY8Y
oKS/ek3mjveAFmPZUXGWHiIA6qZ1zSvZm15/pRFDkkqD4UzSBmVmkzDGW2iGnAZO
9F3kpod8oUVplzU+Il/e+nt3/d75418cdlC0zSK0qRK2m2RJdNJg+ae8Lmm1pqjS
qUR5s/C8urF3gd172oXRi6adsXqDJiUDJCtI9RTAIUVwAFri23Xkdht7+h8Zy3yW
ZV2R18Ph3BmugVvWw7sfuWUWWYGQ6zQLqXdEDPY+mQxUd9wkhhrXpBEed8F2DvDa
ftDmugVdyqfRQ/bSPEUxNNrGSo4m4C4ghzQCIIMLqbcubRFc0o/S/WlSVlLojox4
dWC2maGSCFFljnhhbh99RkXevEz1fT3RI9b7MdpinW/h6fQ/xtmSWoZ6LFl8SAKQ
AEhF8zWKiI7krmuBIK3mqaK909MEpSf7btuu2lVIWUqyvKDC1wcnqTDZ/gAjHJXO
cRStrS/+SEIcUkFObQmKKRlApwHaEk/+cH9JvXh/QkZ7S3zShmi/4sIRRSzrIfOV
SWkxXIJ8ur3QNkTQv/eAatZ1sm21Lbi4G332Gneh+P5DfxGBbdPPX3qbg7BJ7pTA
guSD9wt4SH4dz36Q0C+KCwOi8tvHT6DE6LkrlywWy/xIwna4Cy+bOXkUxYbKgrxj
CPBFsXAqP4IdvJold27YTj5SIxosqbjsP7mrtMBTW2prI55vIF11M8gn7IQra7NU
xD6SosCI40l+BPuaNRdrVnxWGA7/aQiTT8T+mIZdmE85i/lmPHpZY25mTBrhhFUX
Zq1Ru3xCX61ebd4a6IogbVwRW5K/jntAbBj4DbTAhh2wu54WUZOH+JjnuLJXULN5
1IuswyNUI3uv3rPLqAOYLfaB8SH+Aim8RIQ0l/Q+864L0XUbi0KckU5m619a5dwb
SCH0So+NCYzBu/mw+yVA+rEtuYFVPGbGROwncd7oBp+SDAuaA+ospUA0zaceaN+Y
Y7KuFT1czz4RlZcG6ZkwHNipqIqCNKmfWJ9ilrBTR8j+qSbWbu/TwpaP7VJz2w8k
EgLLcjmAK7ZZMrHK0p7/97P9TTH4MHzvENyy3YmKwpj7nz4SxVfEu/CLBGNFr3Xx
cdJ+e31LkXy/BNlTAw5M22mHzpn7Q8cMZC16wRlkhjU7bTrlTdjwDF0+rdsTn+7h
cjDWvX5vc0gwo5kTellQqe4kXCabiy0Q4eHzzaAyjr9xI/WhFgZdoN/K5aTTA/mT
mvGyvPeOUL+EtMYii8jMQJJxLaLseL9ZTAE2fO/+gc3U6oNicfOYDAKBu3WFc6Ot
rhYR+VFyd/C2Z4SwbprSdjRyKYnWugwFuxh4MuRV2J31Sdf7+7LYkBrmYXOQZNlW
/pZ9KR8y+zPM0J6XYWjneB+DTtuXl/u8d+Lw5wDWuMUmFi6LcCkGgeDjQSjIy5dt
HabmJwh+pwFTV/M671heVVgLUmDGte/6H/LIvbxCBeI6OXnLt5fJJixuYDS26L+U
oLwjEpejiENERu1iVp1G2LuUDrSBsHUyh+bjCsJ2Dc7gqN/vHzEsIF1+YFwvwE+G
Ipz/LbePXMb8vNs4Q15MAb+3JjrmBTC2R730hiDbhyVzsVIkAZhbGyOl4m+oHZZX
H4JZpAt4VyUbW92BYVaiNtLXUDjCiwkiQEWy2W4xe6vACy1P1bhUOwL8eylGQQN5
z/VrSb5MPlwnoE+5RCPCyv2pdlcPsvogw2FIpLwT8T/4Q2997iAT7tv94+7YUTng
gq5247GccEWpPx7bFrDuNKGjvTRMnyWzhOIMb/qS4dRBfti7P+5nil/0skv8BdZU
tj7qB8XccirXcgq/DtnNJrSN/tbo0qc2kCBfvVbuXTFoKfEIDmKIUifTYy22ddrm
6+TYsf/iRQfI5cvzW3Gdpl64wbmN38/JV5nprP2Q9Oo7pQJt6sKUogZ+3jZGmtkg
KNR+setuSB4DR5/zBPe6GCcwlbSvKnMmpB93U1tyX7dNlCyTrocsxfScL8GwvZST
ivRHYmfwfWFnxeocyYHSnTLB4dy0GtBXiXEgEo7idrd/vq3BPR0gWgRpgEG7XOCl
J8oD98im4hOB9YrV+4+XzZWPa0YdM3+PkIywFSD9CL0zk51irov/HB94d8+GgkIG
Y6uE9WQR3+xfNEeswPLsi71cA6kmovgDGmaA95Add7G0EgSTmgphQMmn4ptrqEGH
k/kTx7XVbKvrEbEZjfiKEh4rnrdchWTnzdfVjsSd8XwdgsZl6nSg33oCWsqV7WqN
Ne3G84EkPX2Q7xNJEnnyN5IVafOq7Cvnqw+3aHx5l/A+B6WR2lmMqwQgF89Txz15
i9HfFyEsfvhD1UicdGZOVZybTmGb/srAFj0Xr86yQmr3Y1oGYbyujg3qwP4kL7GH
a/cs8BfUmynIOleJQF6IkhN9e9DAQwWQVw3QSD0t3o8INU/scdjMQR/HmRN13rfQ
N7n912f0KODjN1hOiWFuPIn1ydW6VAd7lySHxsFE0o9d5/FX4zGn6xeF/pYxs7Nk
4Ma874BE/n8QM/XjI0pPX+va/RvLWfLUJU5zV8sAYQYEzM9gYb1MZq4JwtcxL8YC
rxXGypvgy0dVIIuML3WeDkhWtGHOJmDpdthx0WKIHxzHjXq3Fd0YhiwI1If21Fw5
4E2WqOwcQCLkwZe8jw903oBBEuOT7bZwObehTqO2mD+cQf4/i6YXZ1S/XJ0Lgro/
R6NmtjN38xARzCi1WcSMccnHRfeeAfnIwwT6RGcpXWk06RRu51ZfYJXkgGGN5wu3
0o9NlHzRw3qN8Tv64jiSFIQp/JZF1pnc8Whk7N9zH6718WXV0EoSiHueqms2KCAX
IwKZZ8Wgv2wFNmimxUwc8vPRJt+l85wT437RzoJs/qYwN5iEP6QhOqetBrN+QfAO
QRfIieRj3fOEX3qka3XDtJx94PA/I/M0IaRw+DUWTkFwBJxA/SbzBBU27NhjNH/S
xDfZdacLDmWQ7cQIBa/65sN7m8C36Pkvya3MWJTa+qm6Sg91qNNcGTGJSEAFrhB4
vNvuW61E7x0LIcYz5bqworMz3Ub+BegPd7ZgICk9eQhjRVvU127XvyaCDyQT4zx3
cwYKRhjz8wbM6Q7YyVSYEROrsoHUJasPEKdyO72gApc6dx1xYhG9V47qB7YopApP
QJEJ1wCSyXQa46Srulq8fOW52ExG3DnWLaDk3/ycB3vIzQ+Zs/YucMzyezsxSnfj
vN6KWAh9jncnMi1Btgm+KNDakF16FJiUxtuYIBpnS4KRqZCXoekFba+c1QkwPeFd
5Gz149TXf7kOrPjme7jrWp9pRzAfqpPsAyZ0MEH1+6agB7FEoabriH6LYwZN+4OL
9c/NPXlT+RG4orKhqczL8xqOej9OqZ+dKCOhl5XPAFf4uWM5WV5q+8Omr4griRi5
xsEJZ5Y1ZT0yC0cwDdXtoK9hyP47k+UXxy2pmjrXaRElzuiwL78R6EfX+GTtnDU4
/As2RiFRANxcz8lOOy1/rxZS8/qH9S38KP69hU0lAIT1IPQrmtieYBgXY3s1pmiD
bsg8r5/FFmdVfVX3PSTdPBVlqVGwNVcgMmr+k3tgufcGkQe+qukUCMKHdKbY5kSa
snbuNVrJIYZc3zWqjky7vZx1HQLVYWldzQEgHkLow0phEIB6nkKxoHT+lcv5kFUP
oMvRUI193DV1HZoqKKJWgWo9IW8TpyQjVYqi6omWyAkUR8Uv4vZDockPkE2Ree1D
Uxx4B4ANbLxemVxUzfvRSxZoBxvWV+tyyyUuAfXu92rnh3BlTjSvhhvs82ZKB6Z/
wwc4lLplMpZaSzoXTy//M1V+mSrDwa3JwAOu4eV5Bfu1H/gGPtYUL62c6gKdJPdY
X4k8zWlPHINVqkuIqouxiQYEr7Cr00L9j2Ktv1ziY990xmaOnuI6A7IFTy4BN0xJ
L2FXXmPIqtslSnX8Qc6D4xobkui7Ok0ZZhUMglCgHJ3LLDRtckQj9gT8Ei/nPiSr
nc84AgrGUmY6MyqkTMu6z27ygg2riQK0Mn6DKVEn0zj/oQ6HK46CjJA5ayIo1mYI
jh/mMwDbJvAWCUL6jBG5wiaWj6sDNatuwiBu/2wh+A6z9kKeOoPyko9eN1NmUCQO
dPSdCvCS4yNpmnByHLGgmSxrpLq7XBxpV6s8wl4O7wyqO8R7ledEGWdBYTEjw64Z
6gJ7RpNLG38/zzv/R9ehqpt4Rlyqi/am13dgK9O2GIU22VvgGmY4QyvBL1xT9i4N
0/HRIsWNkpEW6vy8fW8hOrAmLfnV6mLzVF6bwlkY2M6rTb993xBqqwvdDmOdsluq
k6AmJeex/DEAj4VmIM68UJgLlLKGvCHtNoC2JD8jpZrjl4XVq63C+gZHt0zWen2Q
DOTleVw/i1R0SHHSiFbMIJi6AIt4RW3KpIhUQhfoHyvCZ3EMaW9BK2pB1ClJtKhz
5DZu4lH1jiIJzTo+cYjm2JIJ/2pIMUi1DRLPfbX8n2naDtnXfu8wO388A5gSYh3r
u0r+rEXckxmDovv9y9pv/49rvwRfXxPU+63IbMVo4f0FZtjBP4O4CuQqjx1Z+AxE
Bh45wna9Za+yj+qKu38zD92K2vhexuqe3qI000WB93q7t+NeR7rWp92N9FWCOwaE
SZHO67o3mV0lWtnyJqNthCN1qQsUicp+7N7faspArBSnq7X1W0vhdluy2aBgrAqW
ygd4Q23GIvoVg/G8PgFi3jEEwFOatwPyALorUqczQZ7ph+I1+dLaZo6hmgtC1SCv
HGfxncTE1WcrAEF3M3BbkfB6yerjESyRn6QJz7wrcxjUBlCbTDUcb5OwkVjdHqwW
IZVizpKBZNv0X1RlB95HG7UTU1minlghF4z+bDgliSnf9h6ccIs8/XDNR2Ft2SRK
l23cN9Ghr4fe6xOoctJjVlFc8KXaDMVrXVbV0eaxwjJkKbvi89OXincClRyiChF7
EhZFqofP0y6tXv4+pR14fqu0Lof52vc/ngUoS3vC8RF3E7AtiABwJqlrGFhrM1d0
n4u99mEgkjdr4IkXU1UTdhlN5DyzYY+PzB0e0xigU5VDzEE9MbeeZdGBcEoY/cJT
eGohCReeFzJxKO8kjA/6RnQE7z/99ZNkAfNDfqFvN3H535+AvdbVlcoi5V862hec
LV5jJ97/t/ccXgwf1szluv82fezWzVrrcAhMd9uhUhHkYAvrPs5qCQ1hT3lbXKWO
pHIOt/YuYqwW/RKi02Gs3GlHXmHsfLessVEq6LwGlnTlDpgxzBf2Tz/+JU20xKn/
Z3tMogYSXxU7d0e6lwiBEgnaLaA+dbmyPCwbKhYDCpsfne/YVOuf7q4vdExKb0Cn
sWXJdjttINfn6ZyhChS0zP2AE5zif24dO7yRgsbVmVIYX3rSZwyvCiX/vob91/10
I2gaacBlA32gHJAT2sFTdbjtx2ua3HdTXkDtzuO7Pv36GHLtFMxO8sxV1r88Epwb
banCf7H39iDxk+iF07idjbj2uuWMM3lO2iU499+vjmVXNhYtBUwyPwumM1XPoE3Q
dxfks93D6ibitkJC0wgtqhH/kY38B+KbnlVgN5aXG6p8XB3AzjV85dIfV+bBJasG
GBFHWYG/u9angZahC1swcHSwjQoJC3BpTjdE1ZlPLN8/IgzKJr01eqijChGEmwcf
j1pvZonSNIIXebNFZQ6ngCi/4HFnQVbfRKHjKrhi+kc7imFSdYzgbKQMP8y7aX6M
aschVn5J6ofv5zcMeNTnjmD+QexRTFWwTobZlhzWcLt30SnzLeQgnphjfgOUI8yi
m7pU8fL4RwcuHIW6hq8c/B+trdMnXTeNyDqb7ctjWI7K8P1OnNyFSJoldlrfPEie
Ptw2HXCjFE21oB+RayxwZodkSdk/eovuIn4ttlnt76oOWn1xahyCAwu9srIEowX6
I1Xvrc8fCk6cV/K2pIvBI06UT7P7TcYy2s8/KUAIdY/RPFlPsDNSKo7uUTl0eRkk
w5ldD4sCZRykKWQ/TbeXLLLLTMfbO3ec317fWSXejRI1d5MxBBfhd9M+btBy08F6
nTRCkt/gKT/6dm8j7DSpzJZ7G/b+r7bSXJBg+WiRsEzFOhU0jjw72x190HHuEwak
2IUBAGXXWFOilGqZ7cpIfUnSty6M1HrjYDlLgExCh7AbfFoeA2I4CkqRPZghcR/E
hyquDttGfSlztcb5R2fyPoNpmMQ6n1w2Z3/1PZTS4Ikhw823P555Mw1t5QLRrXJ/
/gQnw/EsHSZKJB/eS93AvncOhDbqoe6eyv0Dra/CMTSlamlDM8dTc9zBvbTi/Arp
5QipnTEBy07K9Fi3Hik1qEIAjQqV4GQtluVTx7IjOIxuu0pwcNykkw0dpO6PD8Jj
UG3XT0GfV4fesXVbRAVXveiV6yHQA5+2s/Laz2lmZG/KmL5rtlRoQCT6N2PeIpiT
2nuvaV/xgi1fseu5EANqKnlKA9IpqBbkBqP1zN+Juo8mi0Kll8IQJsJqNczMB8qO
2iBUd9y1z2Ir3UgJuvM455n8isi2YQ+as04Brq9RZ7anymHhf1+t8GSfSziVJ9Fr
7SSieT5qEwr/1/Th48fqYoDzPc7ohwD7AWRupk4cga7nfIiVpoBX7YkfIBJl9WZ9
7La+j/N7cqKbQVhyPPymu6sdOBpFC4jT5KNQrT3T/2B33MJztAs6cezlX0QG687z
cerrH3ex9/yd63b13KGsg1KTwXAmUVEsrrLoq5FZdWOpmp9rkmt8TbnfTNxZvt0R
tKfJ7wntBsHxgv5N6ClxC//yNgcsj7N27GeuinFCpfQ+FMNL00uVaLtNg/bwi96E
6d4UIencE+0RGbdw71AhC9JlPWrVtRK6kf5f9+4OQeyaDU4to+Eodaaq85PyK+S3
oSjVQk6IwGEYwS1mFXSsATdkPrc5KFDiXaai99NdD/dfL8IhxPrQ9evFoUvwpsVO
LrVkX7yjwqAiUoa+wtUjGK2YjUq/N0dJLCfc0rBbs2zMqARwEk0NsF4fnpeixnwa
C9fr022kAaP+5P0w6j5KY7XpKBigW1yMa5p18awyCICu0j+BGgy7RKijrKVLKkkj
XEW+9tKS5CyW8Ma/HeCKEmK3egFoYugEYP1YtL1G+GvWA1LDpaDA4N6JOh2zGG67
KFbVv0jhrseo1zB4Xkx8dVjBHFViJf/O+B3j+oo7M8lCO/jW8FQGZzRt9qp+TpRR
sy2E5acPK5OrNmksSLaF7X+YA/t+gElcRX9fepc7ZOz6kEtUOM/1Q2HFB9wMdFbl
HQmIdTotJpv0v4Rpggz/dLXUKjBrWs3VUrdt+Pe55gHyEayNcObJllQSlGbyYVF1
XJ6euL4Sz3vSHS9dmAKV2aeeBOLAEPkGZa2scnScCy1bj+aFgszoqLmNfWc8caIa
iAKd0XwYoz6wDjIwhAm8WsigxBdqMNEgz75jUlmX3Y4gXJjtKZBP2Du8Y/cfZfxc
x4S8AF6eNqh9P8f+UmGfG6lR3mZ8kYqazbZFx4GahrpM+wh11H5+sH5iMWv8dG2H
sCBSngAoPCzYKAdRlW8pDYQl+aH0BsVxFEEOg6OkIa7Gs1SnqodnJtur/d26+YDE
oNfVC5GsUCV8UCve2Lj62cBgPvvwxB9Ry4BvZtPp962l8g9QXoCaxZjVO2IAxp1Q
iHXUWg7PbREFZVH3PVrXQ1f8JILV5IVH/ASFtwNf7MTwkYVAE6Z12qG1VyVxFTCE
Nx0ZhdGjwRcDssPQE8/+at6E/KfFJ1yR/T1gEVSndN9Jt6mcJgfUjFm5h1oDhGcD
g/4vuNYzT8oi/nM0yzT4rgH4qBFqjlQrw9J/w1BlxD4WZlUXn1BybNmuZxRpNSTK
Z/jNBC3mCQJxkhKUTF8TKj4SzEiJ06WQ69arfjRUK88oXBBS9ySCOlWxc0gR3Gr/
Vn57z0p4VeIiTHzAU1TUIALFTYQe4jxuXuzaVKxgOYngr47EZUlVwmW8JVEwL1GL
GT8geP4pc+8c5CTYR9KpEUecuwFjr2XuqhO1dxCbwHM0WmF/W/bKSxdCtxjEN6Pc
0Oybu+5s/hEYsktO8S7ztan820OrgePHqK5jqDrdhBZP1T7CBRfaAYDG/76agmzO
/+YGkxW2QGm/aiJZUavIyVrqMoRuUI5jJ2eL+CJLDm2guUt2M49PTpq5+qzxIBQk
KEcVVLynNRY2GkZkTEw5MBiHDMEoMsleKvCNFlfUJDaKpLc9ZOgyy+DdMWBhvS4Z
dFjzz/XHMcsvbtRZ4CGahcGPTm412eDcX+rKTIlEe5BYlspHQaKI3jWrhmWr4vLS
P3TXxgWzO+4/axMo6cTJN8qE4LZ+ZdDQVyM3JSsawr31mWD8p8SF9Z5jKWYr82Wh
ehpKf53eENX/cH1DRIqTSev3Pv7SNWk9Rm8iB4A+xUlp6Iu2K+gwnjjWCTdUclz+
LFt5v1ucmjwv7l02yWDIaS6ep6lNzEqdwkPhRNI+1MiAotVdBmw+fQwSAMbI2oSS
vwkX8IaeDrnSAX+rCLl2l7USEFJwdTpXdNuFhj2pBBhV1NBMTVVNabA/l6HoWAkr
sxDvhna2NGzgG7OjpNWCyyemAxbMEtvtOtoGVbyI42S+CSxQ8xApT080qN6Tbj14
1KbAOrRLF5ZZnV5+yCmbkrVOd0qnswT+IuAi04xuH9MPeDM3e0Q8H4wvrg6SsNnt
l34wnCI7BPW1WF2d4+q3ZmpBBzL6xjDPZgRVAeYcOkROXkDqjAstm1JRTWAdvzcr
N3hBIFIsEi+wYIvfaSIMz3RGUt36RWYHd5dKtlY8d4uzvxGAm3z2w4QDibAr/5la
kbgXc0gzOKmeFo+dGjVtPx9W5tbWZ1K9qcvA7gobNxGHSnTJg5RtdZFA5gJTxPmB
BsBycwRjZ3MhEvhnrFoL8Qf0TprEOf5i1G/GFYvuuZTdNF0pIaxCJ804rWPdfPuY
nV1ia3sVF05XjBb1cOVgBekukgIpdJBluZZ7cTzdh67+WPL69kkLkSYgn18pmjZv
fIbDnhZ+OeqRmLA0tJ0EQgvnzZSHzDLCjyZNDNXWzijKu4yH8KYfJEYbsKz5fUaH
NpjiA+BnSi7xodzRJEfck0KagSysdugw/5PYN6Q9K0WfXg6bt4o3MYiLOHh9fH+c
I1Iw8HC+nHbMQYVeQ+ujJ5/t7AVA/3bhn09x5CKDZHn5e6RNL6uxbwWeQbOqBtMG
Y95mAOBUaAgU2aJCWD+WuPiHWdXsH+P7vVIxT4Oix/P0Q+2iM20LVrFHuk4ztY8b
GVUa818PB3TY0PQmwGFVBpKUNV0q2NIVYSpikA1Fklbxwj8R6axgPjd4fCkdzYEr
/3ByLTMEwrBZSBu7LydAbWTzwDqDoTyO4NIo90d7zaAlruDYc4bk+Loi2RuvZlDz
1daSjQ2q/HBrnDJDdgPYQz+ayP1oowUqYFsrQ2pvsl0WJHGE09id4LJufVzJ9NED
iwLoYf6psm6MIGiFJhxMuG6jkjmHCRRo1T9RC+vy6iBUdoLWHGPYa+68PFeANPYm
Mes+YZ5Wbwc+tC5E+RmkCxji4KfRhKVO/rXg33upMGMEq9EEIVEKj+6omXqkfaCt
9b4v4r9ZVbVtVnfxf2TCD2I6GY7//7uILOtyTfGECrLNasirMmtNV51N7OQOp0R2
UZaOC9/6jEjdgynaXUMNxpKxKfCfd0cx3uaiPN6jqmoV1bPl/Jfg0iJfDYNfpzIe
E938zsdEbvz4BbyZO8d/l3qit7FuuAYi8CfiNzbokGS0ZO6ycFuWpwDyeMO7aOme
P61hhyYlsfEYj0szSMzegCPpytynAnqNX3AuSvy4yr4OeBMw3sGMD+hzf0fZHUtX
gENJH3Xwq3TSZ3yy+hXNMMD2izBrhXUvYdnyc8e2zi7p1T1t/8d/Fe00i/SZTbI7
kInV++wjxFoEWpeQEcBZQP5pK9Rh9g3mem+05QDomJLHdmj+6W+xpmAMPo+1WBG1
xeTVWR3R6lKZW5z4h8dkhqjgrXpDmreM9fllWJTp0ZmUNiCgme5Cu/mRGCtZaVnO
elJti8Do55DvrLJv5GWoR35xq0+ggolBTSXk5SBjJcBN0wyEcaMrlEaPVBaAbZfP
/8Jn9CT2x3R9AGXicXDoDb3IZisUyL5nbFElMKpUWVnYEIC/82eiM/Nk8tTlvmOZ
8/vJHp1seAOcr2xM2DKCrOc+s7SnwOgsorbJjJ8o+ikf3FMQPuFHXKdNEEp9ngtM
GiRi7/zvJpLIX/waeXq6Bb8urwym2ISW98Sg8ktDLgMulXfDeolf/jkBDUankNt7
6jqFOf4xLmfMylr+NG57TP3xWos+oXQ9pBmDF/eukMr4qtvW2Wi0tC/9+knUFsKo
YRROTtZMjPyEL9swF36QY8uZXoI7pE6KayJE2c5czM9eT6oLS2fMs/UygzZJXvo9
AL/o7mZqDTWWiReuXf6noCwNGqKmKprValsOpI9FgOGsyUIQlxnkfHE1KOpJTPR8
HU9A2LjcvLdtcw4zey3jtQ5ro3sGknUNqBjJ7F4c5IcorDmp3GnBtJx8A6e9/euv
VdRSeXZqs36lk7kjZh1sAk+o1prsYJ+1ZhBGn8QMU8+KirNIHFMArXDwhU7d6aVf
cA+lGT7/elagYJgA8m/VHimlKG03e/6h0bSn9+78TC+6dJJEV2LInAVLOWyhG7ua
rdmx0mYvuZQ6s0ALxLzaKL91FJUQoHPGjLd45i7EnzOs5qbnDkjEGkh2zafTOqpe
hBQMHh7VXpHlqa7PTZS26hvDoc8pvGxPrPlgtUdgLEXnwBrz50jM55kuVQDY11Kw
OumlALiskPwckM8Uy/mEk94OEvsTuMKQ1PXw+ObZkWrlwIeOwaMJlAUve+8RzbtG
l4dTh+lErQR5Lde/+QoVb89xWPVRsuDzPjNH9a130IOnipyuxFK4LfXXrpag4Y0s
9xH0VYPu+EPZK8P1l6H9Y2+EQ7O1lB5BmzHU/h5JmBsI7hQNmBl4HojH58tsYtlC
4o5xv2Imv8mMasqoo3vSaXJ53Dto5M4ueJM74N5AJ4v23M2e+hyJ3Pav56Kqgpjx
bjSom8YjWqdSKG2BtYyLSRlND5RuZNcBtDovvJ/NzlsPZTVmR69l/tr6GK8p3KH2
BCdVN6I/11lBfNpY5tHZi2r5jltPC2fDtMvUj7YEsftSK+2sxmIXeS43lA7lQ3p2
HpaIZMW1oCwHB0GJFi8fQpKG3ibCbZX0iGDWIC0/rf1bgZlU0vM+KosOJYDpoa/j
rpMcv1dclsQzvjBbS8Je6pvA8gGIENrdhk+C9ERzuJEcYLjVJMOwOcqKwMZA4VQ2
Gpttlxy3Qhxy2n/2aOHJz03u9OAKkwDND+Cbex5YqZZ+/vCtIfvm/G03FI8kl3Lu
+c8tHGway6I9tyZ/HIzRz+1yiEG/KjUfi3UZiqUZP/1WxnaRrh4g9Dz5Hj9EcA5D
hSJIORaUqJDtpSGkUsnwlQvkdASbTQP0RRXxyh4h6wEsBV0BwJJMdZ0pn5Obgk/e
1uszmm3z8O4BUO//yRJUvo6X3r2+RHZ5PBEVNjKJNE48GKuQZ7OvY32NTXhcTz9Y
f5qPPLJyfhO1bAgQkN1zROVUSM//ARmDQpOqUli8P9xL6D+6x2kNUUC10UmmDV8y
Lp12tboNxzfenhnuILkBf6zrghdlu5CpJFsVfM4X9z76uUnIRon/fAmXSAvUI5Aw
OaWekf+tF0Iy+Jjm3gbhNn0QmW0uZFyYlZ+PbTWvw6IlENrpA2sR+R1X3RwyzeAE
m2hFihLd20GDqJQwDsV18fcNHpjdvvhncEDoLhRyKFeLXZ4cDZXBTscQbJHgQ/FJ
3NoB0DBiy+iNs40RG5J0UYA/d7MlRki4TxUxCsMDJQKHW/ymLmbTCS/O7D1I504d
+0UQ9cwt8gqCMswamOO8/khxKnH8/BhQfxNirdx0NAoZvgkMvPJB2LPyYWeP5EM8
xFWljuGWRRC1K9mAeyXXDkP2Gqz4BhR4kFZKF0eZIy15fPa6fQYVS3lrOnOoEsSx
ipcBeJmKlMmkaEka7Zosskeqs//UEQDtX8bCcMdeswtbyTQncUrNPHxNV4qMugJJ
cP0v7QEzXKlKiOJWvgkL/Sg7UBjxNv+ld55cDfT8OtEmfet+Oz7+EEcRUhdrG5HF
8g3gxEwbilUaM/g/XLlWYNtOvGXvKGDDOkCA2Sm7DS3hh4KzzNruxAA9tE9+qU+f
0hT/P2sSxlBO8xiyr2sZPaEZG0D7SGCr1yZVA7xgU2w8GaaU//yqlpZORIBvTEpR
MbibmA95qJwKCfGV4IMKQP22230gsDiMggjHMhwEB8z4KqKgO6AORFqoqK7qOXv3
CLoFetECoEiNvqUqcE1Rh95czHrT7uy7oktZW57A0w/CyvY8RvwKkM6c0ofyLgck
QdbwukxQCS8R6AgIn8gt1jF2txUO0TUxhds4Lmfo1c5SnCY7Y969hKtsdkQ3o+bA
eqe7VV1PzT+eSN4XJXx1tJT5sLC4lOc0WIye9vsXwVzfKJyNl9M8Z9/McQTGOpus
egJapZOK7LyGUu8q2RVEL+8wZ8XXuAmwPPzFbZODUczHDAC9LAgVUod77m4RsTQ6
cUNl8f7CXXtf+byYnGka198N4wO44SXZgCClLRtiK1WlouqrlEWhAMawWuFVe1wv
CApctQ+7WWBpd3CgdROxeA7oAaW3voK2Z+uFGQVMWHh4zzwZn5q4W2RQpKIYEFxR
cEQlmjfWuXalLVfAD5UiEiH3h/bCyejQFbVygpcWiu6++RTAHo1/QKxyW4/ACFw7
GehBRBTbOlO2AlBvuLRJu1pQq9ygfubKv4HDJt1S8rwJFtNbQ0PM3IqAnD5O2vHL
LNd4Rr8dhbEdJVPDeGoktHt6CR3OLRtjbwS8i+deKilBBvPrzebDNCikXZyYeIEy
Czv6y/oIJHJjRzsgfnxXdaOeDnTtsVJTX9ZrE6QPnq/yMqLTYtShR/SyeESCdaFF
h6/YS98yV8d9GPUMAfxdR+nDE913PLwsZT83dlaB4n3jJOl1OEQy01B4gPqqFNuW
wSSrdKSE3xJQi6olGhDC3U3CU+PogeC4R8I7G3M6HDB0TtlFLwpVu4B526LNjyb2
uJl7Z3sWoLbPGEvyr2mLMhx328gxchbMNVQ7T9BAAlaRUUr1nuGm4sGNmHbg/eEW
eQ6A8vag88Lhyd5lV+EzsvtY302hseMMk63hDo3vJ3dMtVJEPdV7FV96jqLoyCa4
4rj17E3h3xlREIt/Y27QgvCF9p6mUwFY9F1lhk+awuClz6JjXBW8PgIsJdkTg3aG
DJ/8aeetleUlr1LhrWZjD3mjsFA70RW+S30RAIoJR1XHZuNleyj7fgZZ9ulkTz5P
rRl1da5OjbF3Q/9SBWJtoJLPbIqE25OxvNgkHvAlRsbBo90nWYd1QOBElK2m+4/c
6xVXgZF3qAnOe3O2ad7YXUvNC/WBnEovm7CJlGLBn2wlBAgyLgLg8ERst1AoWEMu
ifIVexzEF/NzufkJ4D/XP9C2q0BwdgSj9U+Wfx0+wpPtULhP45VtnTWZU6Hk+gA2
uFsACmtS6W0dXrHkNLUpiBcMFUG/ZoYWj1EOG2HuAvvNzR523FH3GD///yIqj8ng
7FJGw9k7rFJC3a+6qv3Z960JRhuUiq5UaXpB6aJ4V6xHx1mgQkZ1hlKRKC4T9K8H
8pxzGnqemu3IsR1zdlKI3BFLH9wAr79ugmA9h3M0bfog+nIaQmazfWp0GljCxeuk
59yCTd6Y//x4ObBVnOiKXvWNCdAH7YOkBeCybbQlx3tVcRKltw9hsNg5xW8v9Rwz
eitQb/7+LmLKLAIB7qDAj/+FQMBSDF0+/pAcEbuGOa5/+n9IHetpQamWdFxdsNkr
xE7L6u7r+EIhRa0XHfPk42C3LXndB9aie1TUfYWllRuJ6zl5s9wxqRW3IGUKvRD9
Wxe2b03wcNH2fyrWHQ5vAaaxIxO3iKBztEUg7L1ytVvRantTbWG9epjiBGOHxLRQ
8bVPwUAstrcgXXDhXsw5hXVJbxG/TYLYX4Yhoe4enkr+oCXd4WpDtzDLlxmzTVhs
w1YyZFwkU52PgXaej6afZDbgMcmMk5kgtObZqkh5fhIH+NETB8wUPqnHpIbpEx7e
yB4XTHp+GQwKVqFmtTmrSU5uRVQrX6UuE2BjKZjSuol3qK/UJGRZC1u3mDigjRmT
JaJeA8ML2jwXSXiqWeFg7TuDTqnEC213YBCf0KHNkS2fUpILVBmmGfI8dycLoXnh
urM1faCE9sWjPPTmDaaaX6pjEXT3Mwq215j18AQX1x5SCu+/dt+ta9G9WbjpyTYk
OIYE2qNqPeY2JLH5sNkTUskYX6R7AujGKofSZWy8tT9iHREGGlKqV7ReZ29nsw3D
YzDplim4lpZu4sEBmoxa8rrrBxArXK3v9FFWt6X66wpp+e6kkSsUgSTu7KaDLF2N
tnpPXLsqhthENyIaAB1LfLj9PkGikJLaWY0AEhcRYdofQmR8j4ekBcGdxZ2v7fIP
4+wBsGtxfuZXP4N7goCP6IrTAAGbJXR7ScDZgZExJjcY0Qe5srJPjcYKE6XafYf1
EdKYqksrpaA5BiSTlzOJspwZYmWfiH0QfwT1zVzgDkAjr+mYGv1BRGkpgxkpcXYn
dGV+xckI2ic9tQ5ff7/DDYiBbWEKgwwS0s3em59CQVoO4bYzLV0y1NGOoFWfIB05
rnS+BEQeGc503eRly/rnP0bu+1pjN2YW1yO2I3IZR/CumbcttE7D67hrXpv7rPnh
ixtq5Ra3Q2WDL7EHB34YQGEIjFpnoW3AYBktQRLcNFARCfLvw0cz7sdNn8UdD5Fl
wLkmbRe6iNyfUM3rBnq33fHf7Yd20ithL728oMw2OMJbxCx7hCaVfLPUGiI75lpH
TJZgndInUNRYmRcLNaiYyc4BYCTOwnNA1Jcu1wu+GgEplWDPb8lww3XHT9a+ZeOp
wre2+9yeCnDtu/oBbFJ7uZhaje0h7Rq9EMsvioImHBdGHrNEflrgtUdT7dDBeyOl
Kmkk4iUIHJL4p+0dTB/v2W1/LadW5ypiVN11UYsXru3PPfmVAAFrD1zXNvM5TceV
E0n/lvrWJOs36pG3YHR2drw+BjgQZ2juvdQyz3QpdO9GstTr+ACsddf7TQZu1RIx
GigLcrQycIgHBQRqbugAYWCvxgGMvSMBbKSFwX6KILsTJs36Z019q+/ankImMSuY
vmCY9zEZqVvxkVr2AN2AeQwhliZ/vqjmQ8D0nahX5ozy5/rLZ6bwtcTQs2liCojV
B58qbzzdn3sO6P6PfOt1nJgBxR5R79E4o9Ieaeo+kjRxe/YyNc+INMUhzrrN3n7z
h0NWsbGXTBm98ua6PGsYTp7gFelS5/PUsG6tne3DqbRfHkQ+74ZO6v6HzVbnyVP8
19GAseJbEWyNPdML9i6wkyWcpaYuQMT4FXkgS6KbPqpav+qICWgwQVuifBf5nCJ2
GQq4KMSOE/ynLX/lW47FY+oLcuADRWX+ZW4XyppT1Qd95SLXSx0LUMyZpdecqWPb
cs8DELXDxfBDGQED3YSSuJ7seL73TVONpb1IoHfxkw58hiro6OKt0/rlmd0xWLpY
PJc3OJbTijB0qKCy4+edsrs6qZmOSj2tvW3Krs7Nkgg3gIjYwRvMuJnpHCwOeoj6
NREfXg61Rab5U+2MVxaCFA5uFSZfIxzUTyxbRu5gMqM6R7M47u/Szi2XkWqss7oJ
tI6Ez0FOkpLtbA9Sm66D2jRRPQb7MbX1FH1dZ0cV25ngpR3tClJaERy8K5gNvP+e
i9HM7q2LG9b96bTMtTZ9DQM9JeSj3ayQT1htmrlpkLsyads66ohZvpbDoV0J0wc/
nNxxj3sqLsPKp7oR12tP3HcWOagk14kMHw+G2+CtLbGKe6vkQVaEKHGns8r1Vbw1
h8BShMjAS3/YrYJOye/joqo1OqEAciKiOoUtVt39F1PSHWxMwoH/dqMAR8ftdoSt
Gi5GuF62/5gZRtc9dZ9ELuMpULGoPt5LfOL+e2hbmLj5TVpX3QlFu1y5JNQnew2A
Y1VXuDZe6VnOv5u7CEoC1ubOlVDUzozmP17qFiY8C7ut3BjpY6E5HkrSpSjGuseC
z/BPn5LqQb9zClsMXK8+WLCBAqFBzgsbm6c26x/h02nADyqph+rh99lkbz5x4dR7
1uEYvYjZPUNUTN8gLPFdeNizTzLOF30tG0DyQcQx29SzM9Z2O5+HSqS2ZY4+lV5/
RL63GzIClm6e1n5WRgm2moBg9MneYvegT1azsWwvvpsl9vrN2FhyzbPADw3if5Ab
FgGGZDaOdPOcxlcYm8sFqHZ3Urdr7Wlad7y8rK82By2PbjggoJSRcmx3OpCyqxNi
0OEzicHWVH5ASBVPFaMSOB9fAyrKbI9wt10VC9Ztt7GT+jENzjPotDJz2j1ziz/W
gGpzJ5a0rTmB8jS90nSppAuDjdmoJLjS90SwUIkHw63iCHATLT32sA3/IgJpZaqG
ETVMzf8ZymBvpbut2GWwYLctHQ7jgKeoSX0vNytlat7iAuEdO/0iAbJGHVRs9MTE
Ldn4yqashaf+JZG/rtNvD223mFj89xaN5dcNOHu9zgMUP5Pk8XBB8ancrOb7INGy
1zLqdrYbh7Y/WIXXRh4mFDBa401F5NIV9OwwyRWx+bDz5+eom5JukHf2gTs0aNNz
yqdQ+FANzVriH1NmX4xf3BqXxYDL6sM6raDz9s1uJ4AYIHfDzSayDFJ6v4CjshYI
vWlz6LBZcXQ012xHK8xTW30gbLUAo3OyKtk9u4tcrpYY6EJi8C3hrsVEgilPK8a7
gs8fC0M4SnxwpfWH4+vuZV6Uu7exxknDISX67uiFKcfyPpVHziTesIsnaHoIj0f6
Znh9SH/c+Kj28jLC1ZdSSZWxG5Y1p0zSYhJEPZS+keUsdtDPXHhmKxEQaZqZaSNC
smxFM/dtQovfG1IAcwTQUSViN1kkCEoR9Kke9+I2VVM48iw1swLgoD0W4qgOVww1
sqNhzfS3Xp7QyFzJ0+P+eSHo4AWqFyk+khPEDA9huGSeDCBC5ECY3crVs1dWJKLW
ONWdHgH43tHy1q6r2yQBngmefcro1mkmvpN4ngppB5zSwN3tialJQW8ocNEQlGAE
9YsjyuUbVh4p69vGTe06K0PZaZlzxUb8cl4jiWx2iCkojxXGnkBacNUWKnYInJ1Z
YvjWjOAsn6xnaMSKV4FIYJoExLKKzinUMzeVA+xdwu9PKymgJcqrf6Wf2/8xVDNU
xP3SMZU2/GLmwzW+sLmDcb7kIs8c9UuxZIUFou5dQv2hpphSBxUy11gtGNBheDY7
bqCPqdVMjEyioH53LDvsPdcCBc237XXsGSq9OwWoQTIHg7EMuTis2wDNQey9tjlQ
rRxgk48DY35cD36yGOB7j+uue4ulAaahTG4JhlSNOKRnIIkZ+m0sPcHVkJKn3wVv
HtmS1fo1rCENSPQKcE4dWu9KRFBaZxfNH6WIOH+J61JVa6nXEiNnKQ2pQzjjy3N5
5eyONTUdojVBE8v8xxRvFB+edjCfdwQP7jbPzyEyLCbOorCitsRJj0n9PdiVApV8
gU+Nc3dhcolUUtoQI4o9Q4WJunhWh+fb2yK9GQ2i6uCiWR6zWvgj93mCSnbR6XDA
+3OlVTXsg62WyGvxxaFUB7iHIe8TTwntjOusU2TknOGwDQpTEUfA+uA+UhzQA4UN
Cvi0wbCahd9x0k1al83WAom/yXQancAvXLw6cMt1edyEqcmbIA3bwrpqezhuHwDb
O0d4XStY8OTkQ6czefWmaO6euMGUvaOsRzn0HGdveN7OATtQ6JzAuRHyNNxpLcE+
zIKsuAaBPElBS58f5QCvchjK3wTSeElFCVasPe8eJ7E/dwRJ1Z2y/1bvJ2f9tBN5
xib/yK/upxZqNUVb9ZrFja6G7vmX+iu955qG89tbBC2NfE47vYkN0KDkENlBU/3I
HmQ6kxDCDmpT2CBJZiTBCvWjHFzxNkHuqjoPidw+/Sc0/OXX606vmctPKu8MPT0h
W7UTWZgMjWKz0IfZI1P55PyvRIXh7ls3QLyJeRHg1LXtLdVQcyWNFQO9/Dlq9kjt
bXfRAaIBGBZhPI89CuesjkaYC64aa2YtZGvmweqJRQdv9H1rYnivzWdNgi95TArw
vOUk5934xH3QsxLfSNoJbjaUWSJEJynpUPWgVyUJlyPlY5Bf0U9DTmFREThY85lt
ipKWFeDN1K/JAJjpAvSPqLmjU7Zr4/wNHM5dktJ1SybPlzsiguBGyqi9zeNRz3uI
IgNPrqmiFGQSlUeeiqVcW1am6RU2aZ1jtEfUp63AyO5gZEscvRQy9ShLw9DFisTh
ez2fUORvNVv/2ZFop6w6Zt3Uj0YxwUIRnSHwEWMHzsI/JDN6FpviJQZwhp+2zOxb
Nv8gSns65cJqK2wzJGqVaYdir9gQLlKWvcmLo/hHjkF1Fzt6oCG7XhlXchHwsi9D
lavXLCmDJdOI8bTgVjTs8aAn0oOsshCmCD2xE7sVDa8flXgF/ZtoGN9zDVxYez2s
TIXEsZ0upghoMNeCUi20XFI+3tYs7vJhqCpxH086blGFP7s9YVXoWq5QKzAgcJaE
SVLlEwWW5RrqSyq7DNBKtNeiKl0xbnwV9kQF1H1Q6fORp+MqOo/w9Mw9C2nP2BwD
uNVw2FgT7fHvZYv1JXZq99cthMIbr7z9TWFa+ltL1ZD1QAo8ZtA54Dv7GF+uBf5L
ue5B0GnOXU5Glb0yawSg7ioMxgH9nerUrI+rmm+naNExMGqSiJorcUnh7CYb2kOV
PVCAA+1IyjZvfWUKXC8tm0Q8+TaL054gNddacTNM7mhDqhmrtJE9pQnN01Jyn/i9
MO1NzVYhcPcfZNmyEw/jR4rOccMiSQUN+nF+kbgir5qEcufX+5ZcIgvTVdphixXt
PDILauuCqx6oeIwb/iI6eYhl2OHV7Du6YnHIE6vgVL3QcjN6f4x9NfhcEjxldUiF
Q5UxRUkKgybdY7EBRTxprUpEOpgdvSEoUozljxM0W/pukMpr4DQ7Xg6mMeFId8vh
rYlJFPE/7b5JSUIaai1DuDA9G2OXxsI+2OB6b/C+XG/ptHJP37liwHB469yQOXIX
EZBxjG2l/TYQDqb/7gGhapPGzDFh7VhS1fkXe0Y/E9/wP02Y0O0tn6MGT2JLJOET
qURBAj+WsimeUGTbTlhZKaRpTmtDABPJzHPT38bcY1cj2PehpFHdLeTU0eEhtWsg
BQNc1Wx4k1psRvHwpc2W397L3gATK9o7lNTiOpVTivI+NAiqycsYSyiTvnvA6Ho9
NjUhIQwTlhELJ8IV5DS9EM4vfjv8lzv562n+/wsYeOd1uYhD4/LH1e8LA+9KNtww
SmvsBdPzZa3vQ2/50c6PLoqDsOn8kQ/63bEkrcf92fGC6ucKhL/3x6PcMQkzxr8K
fZHSdjXOtRMTkr65GCPYKHiBhbgP+t9jpgGcCFLf4SDSorQsli27XrC+wrxiRm97
iF2sgI+AVzvhFP1ozFY5FmAAG25YW6hOiMm3toynmhiNEQj7D4ap1wfWOztoqiHH
r3io4M+M63VThdaqcNszqIWk3YMxc+ZLOJvDUPreyG40/831vauMtS2cb8NNqe5h
4iLy8mfLpjhTBybVfTF8lhVgjcK7WkwJ4eH+jSCMq/cUwa9Tungi8nf+AOkzlacF
U9xNMv9sriBmIkcJTuSvV86ou6EvhltWFVQAgi/pftFP8uTKSsX4aBhKPxYgaxJ0
PDIknpTBWo5Yy/Yi1podtrrl2aCxXWq38FXGbcTOZg5CPHld6fMw1xAwx4pTrI4k
YYycOIEz4iUvcSugqFlaT0q4R3skif/IaoxGVwFUXpqU9R+VegSnPj5jj0tBYiZM
+dFo89tMDQrlg1ycwthBBxGyRHEp2hXj7n9klRzBXXXlhO2aTXR59JkYvECPWUTw
/ZQ1RWflHQrzIzNFHnkBaxEpebpOEU7JwrlOteNua/NA31LosBVx46aRp8JfRXEz
sERV4otgLP1piZOuDwZhgh3Cm4qMx+YDrAm1lvGeUhpiRU2bVJvwQkjsFnA3JLS6
wj7LebJixgnAWY6ihh713fMrLrx+PMiEu50nAtnfafJuO8AVTtwk31JYmO6VyFtA
QzWwvoYEjdLrsp0YKCXxEBO2ycwM7EkCZfGgjnbb5Q69JRVhYsV+Rg00VRZQVE2n
1l9lXUsscmcbimapBeHB54yQr8wAFJzvrXJ0xCKcb7lJ+KrYs0oVD3zPumH7TmGN
FbO/q/0/p5pIm/aLi2aAi6Qx7IpbScuFWXMrXzw98aETf8lAQ4yY1nuf3IpBOqCz
78nDOX9TZP4dObDQQebhBw8CKxoVolGtJiZXOziWTJfwg1+gSKcjKN/E9G1hR9m+
2jUFrU0QUJJaDSEt0lnxahEXLhenP2WA/uwpPCbMd9JUlbvAO7GYJme60Wwr4vdk
xEhvARGg3uQDzIpYoWpTB9JkWOJ8xZBpUOZUx++MRWOSgzIx2Q5VJAR678peHXt6
hGSaV8qvZqpFVi5gLUz/E1CtqhgOWJ0C+kyUkstH++PkBDur1+fl8pJUyvsbYARU
Q50Zg11WrQIJj1Yb5aWm1DjcKtNA4GCC3JOIb9xGXAuqzCEPq6UqcmzzkOBH2X0K
osgH84NC/zpm/s9QxnO55027tt5S8sxpSOR2nLBJ3qa8lh6o3reWOOpDeOPCMEWH
kCEL64ZOJr2pyo10nQOBBjXfxfYgrMXp/yt/1IfcS7bMnE4NKAzJM6lDQtdHYyaq
srVVH/5dnYYW2+RWJZs8b6CSaZxFQ05Fw5l7UKBwk1RcRauXQIEhWS2oD2sV5EOP
zsVUHmX02Z8h2doD9v+16WH+ebD/fA08v4TtRjd1zlWcRM/GpePsDRZS4oLz6zfJ
0AYnBkbPcPxV7xxI+kahDJz2WiLcyNsowQ8mfqnlyy0wHUyGqcs1qmE3rHLXIpT4
zGr2Mihb7Z42n2ym3KrfpVNTsEc2ypzRAVQz60TYInlr359A0zzA0N+mhVu6JTGf
2beWouwVkv3YYBdJK6tC8CsEd4TExurlm7qiUIWDWXRP4U6xQh2TUekYhPfWRadG
3AcTgatuc/FZ40OwlTZVRSu/4GDDxl9BuNiIG+6fdRjLPQk77+BvdLR6zTFSpWe8
eJtbKQShmzvXNDbdvpsZQXpv3MsVke6Hfa4kCBY3S5+O1jB8Y9EAaeLyO8cr0xOt
vESEqHSvyVyuihteigDoZ3JPjc15K8KT7WYl991GFGwjJ+t75hIQGq1I4lU52IHm
/sv399SkGM7iBRAMNxB0ZcQZpFuP81OLnxH6DwaLDC4VGeWD49oOHK03xo9Bj8ZU
UM7jHHDbFtwaykcAodq56YFyBDfau2GD+kpasW1cxgl2jOCOAr2ynmuKTqvR6R3d
nPrGX8HvcELWiA+QSdpymYYI7ktrghtd+QUr878BgNq6UktYznHsaVvPIsIM+PlK
Jdclsd+P3HtRua6//pvylCqXO4mr79K5q7YG+af1ag7WB5gLdqtIHVLv1L16EgJ7
HbAYzBQlvgfJiCcTyuJoLi/HLnN+JHk6TsA+lbKZ6vwQEcemivNydyfBWq2mILsh
wIaeIsPgu5Y4I3Vig/jArHGUSgIHWqpeIR2w/MJ78R5HnqMON0olEIaNljdUPgVw
i0My3P+Ugh+yjUBg9pQt3HZNgL3LS1hALkuVLx0nA0U0wdeokqz1pZVvoe047fLh
rpMbPC7JkH4Y0R6LmMgMPpveO6kCyZ5rDdmZjvc6jNGQPx4s3jZ9WFrrmfwKryxN
e6EHqFOq3svsggut8SoCgFZee++dNK5WrwMYsClpdHjJmSkokPLupUfqcBNgSuAI
yNRUXQPijP0t+QRmX7kZlSRuCodMX/4shdA94XXj7hJn9P7TqqcHcqs4Tr/uKu+P
ceidAGlI9lTTX1w83nlVbjowVuQC+t2gbWxbsmISf2nawN5448KvnHpZDcSFldoT
U+2j0DK/aofoq4uUFdOxzg0SCEMBRtQQagUw4I1pIo6lkk1ofzPVenp+Fm4RMv8A
t6p7hp2Jg+AgAAZZGXxVL330ERIxLnRPoo23+EuMmCowFf/kT8lkxb4LbYF27e0c
luJx7jbTz5UsS3G/cmGc3CVHpNW631EvqOa3gtaB+PfGqVa8c0+iSSkT85IsH75C
ZKWaMPmQwz5MMc+J6l4+NMt5rXDDUN3EtDl6opZm42tlIf+P9fE87w+/DoSDpANK
Z3Art0ESGrPSajfd/1o/adJ9s4KDPYjJ/GtDgSetLDfPRIv6nIRul0FxFLXY0CGT
LfPq1vFIRxAaiAOoZVEZQxgcmh458nKgIzjSa5w3CZ7s74NDe5EwZkTuvDc8tOmb
lw3atlY6+3quuKcxOPB9nQuftnIbq9Ma4Y4cw/i3foXHwIRhkSVZZiRIAx47XnUe
cHYhlDaz68eAxriqt8gKfJNrxxl9l9isAzGykOOgGbOW/2wnqOUIBW2rnPJcd5TF
aQWWSmFp5JwN/GAaRNgmibMBXBm/KCmzH4XpfHAabb99w1Z1WW6C6BH/baW/VoeB
1KafjT7yvY+ooJ3hyHjaM08tNJkHxrJIUK9hbY4BYvv5i8I084b3SWML+a5t4Uc8
sz7XWicCpNaC34bOPVZ92pf0GmloiMvWw2CPDQfbIMtq36bAbTpvIPGHuJnaFOBa
NcoKCoAoyid8ABhuDRPP6pIz+6XAywxPBpjK0v0N7p1q5GvqLYgtvD2j0d86OuI3
187aiehG0YyppthegfgV2cVGxDeE0PPvCGXuaT/LKu3BCWAOPp08G709v3gPzFKf
UOgKFch6eG9YBWbvR1q7jSN0x+mpGSZMzVu3Txlk6+lN4tlcqaZSq/PAPrwEMrQ5
kLvBDi0cl6XjmRP0RiPurpyQ1RziiOTO/yzQdTv9xUlZEoTbs41PvfvH971kZmm4
IyBh7qhV0wx1Yl6gsfQWPsDq4F5eEkr7KN/aG2k+0pYrAxzYIJtU2JHhOsY1gEyP
/vkrQvcxrYtKinIQ3SUMrmq+3Nl/uMeJy6mTgOZYdtg/+WnjFBGv15kxOK6GvMsR
6YoyKOJVEFbD8EFgDAL4AQ5C1V2fqj27otpdG2eMqEibjdDNthcYgJeFSBEs/wbr
LgMGqjt8vH16q86Wk6osfuymvixO5ph3vdbe1kVL8M/EhuHfgUiBIpv2EfOpmY3X
ob78zIIGDTVt0/KI3Il1S5VGJ06haeGuYlqWegYnuwkafo1vzn4JRHYnVKm5DTw+
3NJmYQUMMoE0KijIGJ8ldn8YEXwxz/Aycr8YFZAZHVYCgPFB06xxyvhGRbpSIehC
pZa+J0KWlrUzoQ/N9O9xts8C4NlxGkhSY7hcq8CBPbBKq23Ma9Wep4CUDfu0+FMn
ufAD1bLU9RZTucR/JHDqOM909TUFRcQn9tpnSN83D0gFqRd9RdTRz8QwQqAyES/R
GiKDMt4v58Zfwr3Mv1ViapLCX+069Tg7aY81wETQVpiSD6d08kcuHXWJvuUbzpYm
WUqCywaDcsqGRIaVhMDiK11b7wR0H7RkEhH41hCtrvBp3KTUEZ7r0jvJoQmLxrsM
nw0swzhZg1mrLI82db2aNVtKhLdZ0XPMiKdNOSS95NAh/ysiBvgYjUyj+f3s4Dud
lCYrQnMP28puXVqPrbv+v1qhC13ulyXtYnL8guhhorUjdiBuIsq4AZaZ3qqS2GEd
DlXCGarS89CljS7e/BblxtoClimadjM0dDCQt7sd18qxtpqKLW+73Po9HygvnPAq
BPc8okuM6HY9f7oXBjL9U9gxWMlAzFEOqbHNhEP/Maj5n0n++AHklrhcrb4YpTUG
xiyWmEFtGm17Z9ybQt3fnDsvv2j0dkYztJsss5JAS7VcgDyNvlidePomCMkn6Hb1
SG2gQZmIkxV6qncRevl9ghV/C7rtYtVF0YKeN6VG7+cLZAo5qJ6wZxYSihZV2IAh
pGCQnnLFG13HZk/BomT81xN7G9yrzgp04MMMPTVxww/wqC+jdy2mNkMv1/YPKH2R
tk6epra4XD30pEnobxl5VZhjHAeu9PBi91zDTWFA8xwbAtxR/ShMlIkauS30WItI
XiQj8vn60QbfPWrQ3UHjqKpIZQ5+aIoC9eRqwZ/V4UBDE9JU8ZIyRd3NlYFlbTqo
aku11t4JrjO4eCvJ7ENJKcdy7cAbyvUoiRdwNa4So9JbJoOQ7pcxb8UunezPE/ay
OiP+Cu/o5+JhKyX0ur8quPxTgXswnavHeYVH03EYUtZDo+HyyMtMLUM9CyiluCgd
rIkvPy43hPoXjcu/klB3CQSJVxZOLcAewmuu9JBG2pCN0KRbE42t/2Lwedf1E2SG
kSI6jCnqKahG1l3oCRg1c3PmzzmKgBkjT2rXsJmh0QUfX0aVo3OfR0sfkyofEMFz
qy7e6oXyPXnyPlSR4SlOgpntYeGFnwwEoU9jOZ37eliWH2w3bJ5X9xMb/L7LmYVV
QIEQbgQmUqB2Ooy1PpPDOpy2c3M1ZYbdfScbWLtrAuNFCPNw8inyRi+FxFtYsZ66
HBlO+By+H6gRYlWzLKffdxBA3xzMzMmvAnFho2zeib3c5miAdLeYmMGxBtaM0apV
k1wGQyzBk/RuMUPgo/HCCPRIwtKcgqrKc8WH6NQjlLE7PmyCHRXuQQlQoOMzChYz
xh+TseC2htBSF9WCA9e8+7ByUG561JJ6J6kCf3t7ABPEyAH1rc0C5b9rHHZGKdAr
HO7kdQoYt6LsHCChIq5ACdJX+VxmsUE1SkAV3RiVLzlO0qyzw8HjgZ7yb3SS4BPM
vz7KOhPD3RzSpVicG3FRT6KWNVbZtJwcAfMDI7nPBsNLNzuWjgUcjYfcnto8ClTP
/PhEO2PKYTNLIv8oFBQ+4FAsjUSK448LZgRLFX6oC1ZA7pjUMnZhypa+nI4A2EaY
naLwxqm4zLES45LJkGCiBpoBb7Xkgji6tjBPd9qWq6USJR0VqvpsGGJC37+KNFKn
oehfX5+Tel1odeNeD3BtAqJ38zYJuqNFDgkoJiKpmRLPGFHAbC/ysmnv7wL7OuFB
Rztt6B8QnXb9mKMHY2e9RgbnH32tq4WbjQLyICE6N13IbFDoZlR0b3UiUzwcs3KR
oEUSB5RuEJrlplDXRE2BC3/w+7Qk2iur7QaLRsjjYKrv/+rloNAXenpSObkbwAgt
cTNevUCZTtsSRqGjS5qhYZcmI1MbRd8xOT1HoyMtJF3HXfY8ZZfn04gyXx/bDiKt
PjORBENnpGzYwZzxAa/DxXn9WMKmPDlLt5xD0y+7vY3H3gxw4b2J+5xezKHNU5Wn
Blc8NKDEeyZu+vyg0woWkDrF+rXjWctBFa0DFyKaMuyFA/1lG0c5fRIuK7fkuaCC
8/byZjO3UFzGbolG0qYLPNIKPXkTNwYsGepMGZj+c4/P5jKB9TSgLjHRklMs/+HZ
m6tCbKUuqkCRRhQixYa78yGmQEb54WoVUvPvuBx0XAQM9v54aCQ3FCmkrnn0fcCU
kC6Vssw9+zF1CXHNf1vGMJoLdnVpqfH0SwUsnrGDsqG0h0ptyv2kEhoJzt77ByaN
xXIw21J802PhrOddEN/Cizn3qTWvM4arf4Gh0dm0XY/kvPs5hf0J2kV/HgdeDajt
DGiK1PoSqmOyfPgKjVHkysCROX+uq5tAZgXR4jHdUeRXSpstIZavgCtgTTgzm1cJ
E0LMH1dbtyI5ia6ywjagbzEqsm9pcZSAG9v76wT1cWbm11fDLdNfyX/qdQUW3oOn
o2v8FdP1Sn4hzH62uxI9ejrY+IB5oK97jx3YR1Akarfsrq6PrM1TacXpmUN6o6al
JSPC2QIoKyELEyucfmUYJ+IDb6yG9rCckU3esGX8mt4iZ9qyIiVAEGeCGxcF2BmB
F9DmhLe917ogdNloyzL2BIc2A0wVRcn0l7Y5XlwiEhMEob+jex5oQ+HMkrMzmqq5
F9xDh6XjqlVFqdeVG8kiVIXfC15HFgN67QAQgni52Xw1BfyLba3pmHSpqpEC6CCg
ea116H6Mgg6ESV2+XNNrliK9XGvprjMo/vGaW6TTPeaXbsHgHD/GINv/jzJaloZm
ZMwTkOFd3IDvJDWCjDOdIIdEAt9Rl6H5cKM+NxTq05yR9xuDHa+E0BHH7RV+18Kx
NvmyKlesnzlyHIrsvo/31jXyWkMWGrWCHkwF0wQW1Xql5RmbkgJ9os8R4/K0VJiV
xMMKbn9NDmkFNSVWyEQknOqBNBcyDWXyTtXMzwFhR2CTV56Ev7DNLs0Xj7oTa4kb
Jjx+Vqvi2Ytn0WdIGejzQAMBtFyEP/S1I6K0bKz4b5lNaAapHEbtLdbqd9sCyvXv
LHuo4j4mSJ6N2HgsZRmdwBxOqU41InjgRLze6w44DQwFanK5A3dR/hgY7yCwWHtK
tDv2vHxWIfjrlMZuGvkPpLO66tL2KhhQ0CGrPmjGeJmx2xV9TcBrblV9jNJXelFb
l2sywqaPZy4/OLziWiW+n2Lzc7AVkHsDeZpYxVOa2KWSfMf7o/upw0RBFUT+ZR/c
dhR/VT+J9XnfeR8dAjEaelaVDpoMvJylesoKRCa5NST8hA7Qb7wlwgrRLe7Ce4qt
8by6UhK8nnRzdDUS6F3IR2yAXqBeThWUzhXgmjTcL4GBnbnKlZqVBaYtaETalfhk
+mza7CchbUnqPZB5Klxel6KVWDlH0U3/hyJWjeWH6TS+yMgnbgG3Pqr+d88qqBG8
+5gxEYhHmpqdcJ5cfdviZt4ngk1t5jA7tQKFXT+1RtDSldZXwAfAGBOEgyh3spQs
xQ7mBGp1Vmf0LLTw8C+YcBiXitD5s7O0FmFUYzyftEvnZTkg4qKzWAMbGRx3VuVj
H15CGL1y+7xxY975qsg+O1Tc3IBvRM8kZry/8FzK/LuSKrkam/FzBW6elvDCTC42
9o2/r4QZfHMLZyioXNWkU3+rSlWzA5bbaGq0C52KtHA5M3IdEwS5DhmXN2A3zeIW
F2d/4E7oqEbqTs3smt3jqLIclUqjr6DGbyY5FEfUWaUO4QLRYtBeWNCnOHFZXZX/
9C0OOD+mqjA2QDG7uAE9zGHGw4DRKZAPjS6nCPNQh59LrmMBQsI7aFUzCJPvYmho
3qTZkopYsOS/C9Uok5F7ekJaflsSwKQxsSG5OIb+kDDpKSYnuFaQFNuJGQokbKfn
F8VkOfgFNu9bI2Njvl5WbnqyknZ1vjr+xR6+cks7h8sqYn12to7+xAUrLv1xN2yr
mMgKttGNulEMeUe84jniBZQCN5gFrRQRgLu6TXUYCmsuUr9+WaTK2V8sVg2RpZT3
ejD8+NL8xgH1Rbpo7KJNYMymJRBtbfVJxtcfQbzEZ0eQpbKpapM5PvrBEmlxd4KX
l+pV7plGaHE394AWaHeme9HW/YYWSVXJsrIfo56Z/GAKA8LiId13YNcGDiiuk1m8
yG00+jAKtqYxQ3nZrPoLiGPqmBU8M7UC3MtNHbi0w1Ay5uzTxcKgwjztAYR17qc7
kzS4uvwsDiKAP6t/TmSTlfawZcuAbBanXJrjfeOkfuUNj1R0pbGpmHlXW5TbxFzt
A6wBqMUvuHQbqHh07HxPPzc8zEowkgYGYmrPK5F8vpd52oSp8QNACuq7QEGJ3RTF
Ne5d6m5kyzSNXHFrH1swqcbvxvbEaMXhyIXzlhK7xgjdhnnxlxJ0tj5N25MPAuY7
Glad6dh8EDwbA0iCSBhNvjnDcJ71NoZUSCvGOkZaEyIqhZM+q15B/d/68dqZwrSL
eGQK68BiSP9f5+WrTDfwWrc5hpSByIHl535IoYeu+5UTu328HLscm4RTDSAbEFHf
WjQNgp0D1s9Mt5LlLIVwvhTLbIuzx4INGSdAoX/AVaXUjs3OQSGmmB7OaFbaC2VX
wjsNUYdt/dhmHzc/rQhkKOTxThXTeoE7/4iLz57I5HFv90/eD/rV/hNdj16ebpUR
CC6o3rtgL4tIWQX1b4Tn5RS4pMfbVYX6CIE/k8HBw3VqUeoAkcJFgS18i0BG6x7q
xjBsZfNZZwQ0/2skuOguXtcLqWPf5egkYUpWl/slLFiYFyedaLcDhVKde4UgRzUo
f/X1OiQdJW1gEL3yfNFa5h6iJDvmKDq9a+VkqSMNHqMxrLzjK1D+WlxS+xqJqXKY
tRkYn0sKl5Z+JrPmasKCEcyzlibF7I8jIjSVxqCdn4EnpJNxAf/NuTV/a9LAaVZs
My0h0ZZSJEpirjNX+e5tG4cclnA8TYQdPk8fOQlchg9MvrLoSH0efIoo3gdOPBz0
xkXYl662m595WqWYAMtgCxd0YRQ+6126sO4TiwOEswGMrqowq99xPt2MUe1Uqf1D
8wmgnj4FygQ5MRDNLOg9KlJTh3W/aLSc056/hTm8+azR6e3pHUn66yLDVZb6m+lo
Kj4AvYISVE5mwxWM0EeYHJCcshDK1dtvbBhdvsLyEEgRCGPULmFEg3t3ABWnwWpQ
svsXCZRdmnRCt1uphuqc7IaZQPmBlsliX/F9lvZK5XKn+Y/aRBiQ5chlg2uEQA8p
9YOiW6UcsZXiX24/DGtdVDufRoq5P9MR4F4C5ImXtV2tEgAbTN7TZVg04EfkZ7Fr
q/rE93OTaO9wZ03y8GoUnC/xyS2ypwrRUlWaf+NW0s6dB08bXLVOAkzzyHkNnS2a
Uu0/rssgzi/Y+7p3rM14iWvOPlUMCCm/DoZvhBkrCALaB+prEfKQd4YMTWyM6nkr
kpNDIFGJvwKyRpgHITs1qa8v+cQUfRgLZ5d0rlrfRYaP2OwqgP+oQqvKc7wZAOpD
oDZKGt5bO0aA3fD883SvUZ5ZQBMPZ983eyFufln0uuWYljIcuqH/WMB6WMRGtqSg
MPy+P2CT7Ju6PbqTMrN1nzFGMAO1EtbwBPf0/teNf9RyGnpoRso9K5SP+84keTgk
AgucNdcwlAUxaotiAh+l0jHOSdIMG9Adb3f+VlczoWkTURUkhsAIUnyeixH5rY6+
gKmonuT823tsWgdLCk4OCeoKQbCbpZKn3uPnj01G136gB/rVhJU0mGA387hWgmlc
b51JnkmxExOVkWR6SQujCZO5j5wTuk8zrh6r/jAuMHlRX264u9A3ltKrMCxJYaL7
z3r6zn8Hc0buDNjOvTmay8JgOkbMyNAHpWL0rk99r1JWknyVAEjyhz0LTllCBg8g
fVMHVnvqG8qij7jeeJr1dF8znfxmp/01iwKIvQmpKoLvBVncmxbfMWFWsB+9nQ19
QePaUJm3n8hrPricsABTxjVdR/pTXIbQMUFuakNqHA9BHzfN4wmXGJ0dfQMBQok2
0oBHl3en0t83yyhrJaYczJDHjaYKXMfEHMXBGMCtMKA4iO8dOEHy1ZuQDquAyV5c
BiUfjWDaaZKJNK/DfD/LFcvit0hKrZ0JHrTgK2xdoAyr6jQU3qpyx8htTS89/V1f
C/yjkUKARGqYkLF+45InVhE9UVWUu5pNEhZZsi+fPCxCUnCn97kmEpjS0L17T87E
Zn12Q8Av8J0YlBWY8tuFNHjZauEhdi3OhCUiV/20AkOqBTXDi+O6dOtMhdzNh6NI
AfUywhGYCKUQ9SGeuiE2fXLxh3eCsjr+3xm3jcP9ApikDmghRC0uip982vc5mEGr
dzwmG2G3bjZgdfcb8p2apfer83AZP77EEVKphMDqHnYcL/4NJCg84gwZTx7fggKK
ji9BazTsYvqeUilZve9N5z7Kigw+54mJWnlAnVqbNyJNkRzQB7PDv7DiKbf/gGZo
XsnWCsWuOcd7uBPc5YlV0HdGKly16+59EC8JZstGtNMt+waSYA+5Y7L3M/EtnsWU
TS6TDsw5zDtPClLrGuiYmFr7TNOyI0HDQmQ4WeVRUv3x4TIpWyUOwlfDaNIJgoMC
A9NO4MOeWHjQAyTFkQ8TZCO4+yEtdTwEIpCTE7bhMHbR95HcOCaYRgCvD03I0cKp
q05S+O8gIrcHmyTorgMACHPYGjN7ZTLFtzCpirST2mPAn+AaP4HhChIal2ia/oXy
vIbwEmEduYYauDWnxJBimQ4pHdgQXhf3ssWni1/xJWxGSsc1HErbUcxrhweddCEm
wjM0gojaFXPUr0KAaD4cI0YHfMl2hboFWQHHGBQvi9aCKSTYxupdz8fUi2D++kR+
Dv6YfUasonQK6To/bPtLTJ9BVsQvl/Vp0uUGLvm/7KfN30OAy//EWFaOadXQUgNo
RWiZcKtuMNeYCF5eRNFj0tWUh+nSl1DNcrSJ6Shcz9snE/go2/XHkzKCuFHW/aVd
CY/JQE9nHHJNJsSY8UsiDmA2GCTWmHMxvGK4F7CRF3AjZfLen0PBU8aBqi3pYTdU
iEhujeCu0Ao28WwcJOIAXho8XThk2WdyHJ/aNqW6DjprN1uGcoU7L0hzprBGf6Hd
ZnVRXx2/ayhB2OkyeMVbF4IYi8ndAHctgssSD0lCpoMvVPWZ7EBt033iYUP5Vk+0
ujscCJviP+VoW1OYo82jz/PuFX68Kn5PD1zzM1pxiesAS+kDnXr9Cr8dXiNPTsWr
Hxql6ttuRqt7f38Mcqm3Qo+k85mL4FZt6Ne71qzjkdVByB8CKF25ANI4ASsFiHQl
8Ci5Lf9n3b1zNtsfLw/U1wZ9hAyPFFjR7uHvUm8ptKUPX3svGTMzjCg2Zm2gU8ec
9qqiBMayDNuDMZUIgjN1dNTt3z+g3ZBKCcFGvxEhOXLuxjiqX8psHEH5MlGuDrZd
37z/ApzQJ7/EC5PpXjBXO5rnoIiPUL+8BC/Bm5Ba5GMDckttC5P1HEBNGL12c7IA
jMmrT7Cr4VhErmC7q0iu4NaJeNIN1BmB4cNEmbZ8F4486AKeS6A8hrgojboveQbk
EW2+CPgpHk5m3RZMHIIXP4LpfLY1bz0xpdsVrjuMEUa3xXllEWz/sIjQaJZGIHSz
2UotFrudQozcX5OYHICOPGK5aD83CsY30y9PPkb/WxITmTfAqiy8wZYhZzD3GrPD
u9dDWnDxsTVgVdtlF3dvNMY6a4u3kS+kY8rdtY0IdlaenR5kkl156S2Ej7m/DtGm
C/ZL1ul7GlIuElxv4ABFC+mWBvZAyQnc+cSt+LbyAM/ZOSKgqh/G/0+kXqx/RHT5
SvUM5+wgQeF+Po2Zh2+0c132ur/OjzCLZoxJpXSA5eN5LhP6l88b7i19ZuSQqRnz
HAyZKk2vCJBTpi2czOkp1fQycLx/kFJsru0B43+NQzRFUfiv9gbD0HgZ8NyJcYR6
hIrY5cUNcGJrGiTkZ6pcXZFoqhbr2uiJtCSUYRZWM+uqZIBJ1K90juu28Q6kJNmw
lGjuSzVu3/RSI7WWs0+27WIbiz9ydw4N/vDatj3pyMfV4rP4ReGPKV365Fu7pynW
t7o+hJH+jod3bH5uYIeVgFFJrUdEvfy3S9WXKyE7kuRtVzcEeaahyFU6wZiymwHm
OcrKiPhWunLa1m8mV7PAr1K6wlfExZh+ODliyim9Wk3wX7VadMy/6r8hzDybA9C/
NcF4I5AsRf3gFyUbaIG67/AUHc2lYPWRl4Svx8gTgRZAhm6RqADQqajJ4vtNyh+2
lVZ6tVfqX1PUTngKxx5m7Mcv5CL9vSSflBJ5h4C3si+kAJse3uEmFBnioF+QZKpP
cEw+TBtSOjxzlxI2u1VeBzja85qP0ZrwQFU9GngpwVE/UNE07nXs0GVqWCR2AyB+
V8aclhppsIq2AM7ZKI1uZEwQKATfop+u0yyAK6ePptJKKFHndVH1mw7h+vIJ2bke
Z5nKBAgiS6pz6xRp1j3L95aOr+E+u99NIXzgSnK4W1MOx2thUUEr1GNn/hCUVemM
3wjW9CYze7S1OzmrXcQ4Y9zls7PYuBgmomlIIcWx47i5V2XzNdfWtEIB8aZ6t5Je
a/CZHsMK7U1SINWwy7Fr0iyaxkmomlCOMOIKmoQ3Jb1ytooMNtgUHxfeOvKrH5h4
04nt5ha/BAxFOTf7oU91x8/BMIsps9D0I5AiXf7s3mGzfwihdNkN8eQ1BN+1pzYg
1IMm3jGqa0l364ZUiMl51zTnp7WbJVqMrYCLwzDatOHm1uf4Vrmh6vlHNohoZhtA
rFyw0UN9CyfC3mpY+nVAhSWQ7FeSCD6mevoU+yJTiBd6Ofzm09R5GdlTiXLgUBek
Re0CpydenOx++ECdpvC8scZQTvicZnqjMNHJXxQ1U1GVKjhIpATWc+ZLK5j02q8w
7wNIDEIDYCcZy3WUa0eaX2QLV89D1nwJtUOrGVpohej+5ZbNKC9gPVS/UkZh2m69
kuvnTRq0FJ3r0wEn+gvYANDzlsivqYCAtegXSU+6eXrxqBmAUtcPLIBCpqbR8gCD
zjEirOJwagID3sAPq39pS/4RUh6wbQK7LfU3nUCdG9nn8ecTt78qAIOz3qqSsdkW
n3PfAxvePD+1uzk4FXelMmVb2RhAgSDH5tX572PABHHFE1LehNOLcXDhXSuzKNWK
itGYeKrKPBQ6dfHyQ4DyBOypCQsyJ5bJHW1SlddVPP5NoTqpn5GPqQpeCv6XVTQt
/5PzlmxHe4XcuKglhBMZRkiU6HNaad7suC5RFB/b59lx7QKczOBGJR1ML1vUaaHf
TqschzyMLF1SGNEPjDEDAoLHWNpWqLVG97Ntij9CpGlt2vd03/2jtQ82qIWfRZIk
4/AkUwIrbKw3ySOa7+AXgh29BWRp+FKZ9Mtk7wKo/KT0tk2VzDqY9ZHTeUU2s2QB
/jmxp6VBzhwZH85sHoeguFORVHzBfaZE+hc4gA8NsK405vqs87047LeYsIB1DEOC
yUGgdT48l5Bsi2OG4XiAQqL4xv6ik6tFyiH+53oDNbmtEhv4Kix29fiE3pPdAeLh
mH5FQKpy8huh6zrSgbIbDnCtJQdzP7i8U/0XiqkWbRZUhwZU8YQzoGNQhB++geje
TDUj+YN82SXbcLwjDGvjRexmUq9e9OaelfB5DtHDkeWsI+LgH6V1np/oOO7mHfoT
+SyNehV4lPOBXLA6899AyGWvgxaohBCy5fnODNKhKvNoc5muGmL6TX+0XhICHCwk
fOnVnqhLrHvO3gv2M1c/jcvwRQcFg2xRxgq1ykWNRkyHezL1e5atDIDm5H/UJb+m
fqm4p585wiUdCXWqN0xNAdjIOKVuyhIcsM4WrMS09662MhHIqzaGGwPIDk0h+XBx
Blb8XvhASqJPPpSY2mIufJSpkOrtZx+nDEDPO0CRuIkB6cS0LdG5eNR0bCPBL0Oj
qGwhiMLSXxcuq1l/E1oktJFU8D3g16v5bgkL5JIOvf+aA4py61rEIItCK07zweGe
ZXv7KOwuRlMmmAvnSmc3X9gXrsmzqURwTmLp4GDQp4WqGjL6+9dgbKhLj/JKCMGX
qhlVC99MRv8HYEZexgr0/zyqrQd+4uYK1tor41f3f6vgf9uwYBtk3I6VBJwX6yT5
sum2eP7Ag54yUfo5ztKX5S3z+Pqq1jynnLbJgXzrEJCqJ6yFpDCQXTT+Mr+vhQPD
ZCu06bC+lWdhrLbp2ZWKeBt+t36l1Tu8SSJkwJsMXZJLlAzs6a2Y2ABu4GU/2nhV
DGL/U9e7wXf0i1D21MmT2FYRT6/6CPN51S7LsTH2XWhqzyRKlICouuexXqnytWJq
cA+BbBVE4waaPKp13W0fhg6/LDLNlBWH96h9YSebeeH7sVPJ7mm8IfCLny8jsD+H
XRiEslYvSPW8IE+RMgGOOm/o1oT4idUphL6HAzv6DAlaWjQJTmyWadpZBXLRxBwd
6jwbXtMi0GH+5V3pTj7rO0k4duXpH0PaeNaXHoyuv+I4QhqwX2Tk8OEOAjWWTMeI
KcqcD4GLRWAuycy1MfKK9YETBmM7e8Ts5l99jk+/+UV1LN5ZLOZRXHrDLBru4Az2
We2LqPbxcSv28zGQqv93csxVcsfIMxtSBTBvWIWNh1s0eTmMwH2AIk9AF2dEs+EI
09meLxKAztVkf501Ebl9UY/O+dtoa4BpqiW1EejdUZsbylrf/emGjGRDQIxHNiwF
QX6L4PNhjGhd3N2Dl0Q0NZ5aKY6qGxyzredE+aOWrGH5H3BErnjrtZg+sdMMc1aw
hQ6APDzxbEpZMxNAModF2O07QdDz/dyY9KUUaaceXcF5gTXhDyKA7UWheEOqfPtW
euFvQfrrnZ1DNkQZ7YbFG9aAhP8Vh5a+/kofobkNW311F8CpT4oVcnioNWCUHzql
Ta9X4id4GJK2h9WK47daMvgDdLZzk3uDk+dpo5LbZHSSwNqSMrSRTlTvP3sOY0+q
jWSQQlf/+OGZfhdReN1t8lI+I5yVI94H7BMmSRQz3e6LDzptCoHWIUldzmfStk1V
ByEuSi337Qbo7b2OZZLyWdF744p3mc3WXuvZsnvqJsNaJhKiYBFaMM97kTEy7jPs
a+i5ARukLUWswQAM4qidiQyL1hYk/biyHhoc1YDAzaj6I4V02O80Qtap22ENV2br
pYFl3XOhltygLCI0xq8PVD2v8Qo7JsIRzGhjR2EG0kTlSzHTAqAoUPjrJSkwiEby
Hu35YWZs6k5UZouCPzB/TNAnhUYhKj0BoA4DGKoOkrN1khMgdZY6xYKB5IclMDKd
pZG4VU25OicYc2TsS3a5dEIuVnrZQfkaXbSV336L2ifi3k39o7P0jX5HfZpINuFF
6e68IC9qkBwL+OTKykpzcN79riTH8LeAKKN0lRZ2Zb1KeARSnx91YsL8+hcH1941
rIRbsgKVzvL1vrV1euVKSoOH2lDHLkMwCGTFR/fX/g+l1u7YS6Vms39F/Ch1yXVD
fR9FtBLdKZBVBXKiurhvK5e6r5BgSMQmAbn+2afg8kDr6tgdbcWJyDNP6iONcFZL
ABaWXByvm8S+JPB88GrLSRGiX/I+lmYz7HoEIWXowMsKysc10Is/X7n1vRu9x7ck
BC6HVNTT0pVTT8MGxVnjmWEnMrXh9DfSyW6+V0RuoPAck/iEuN+yiC5VAizdJF2X
EnNjO3bOklmAOkiaEzBS4pV3OIt1VsCSU4WUq3DCNqaVRq3BXDNFNsmo589sXegM
X4Eri9tWocnnTn7qg2dqasTTwSH/O5/dN7hnfHh2uMsuv2kttXAV2LJGgv3xbC99
iT06pel25rFpO6g16+KWwp9G/odxCf7pCU6rM4pRqjeEZ9QnyKH+UGcxfWQS36gm
2bNXBQv3Lj/kZFx39YcErttgWpnF42F41GHI/McTLs0/gPGtFZZTFk6L2Ns6IRSv
gho7hfglzSMxStf/fbd+P/9a4fIetT6XxTnkIX4LfxP/2jBGnyB+HRZt9b85MS0I
8T+Rqy0cMvkuH+khsppXLRq4vAibukZHPCL+AFiKYjsHCxPVrJtdN6X1TZo0LmaE
EoyfNhTsixRePIiaCmgX4TaKAV5AQF0+HWMi4EQbAjlzUDe8t7o1oJTBa6jIOTJN
V+ak/O06ZUNuDdJePoMkb1Otz17zD9oeOuE6e5oe6PK5WV0CfvjP1ItYQRHMQiYc
IjzWBEujv8OfbTcg72SP+nJSkh0oNzZCmhMo4e9zoEmGcfudHKNk67gSgmUZqITK
ZXYdD8i4mu5JfDCpD6xbIC0RYOYimBp4/4klJJEiuMIajLCOE+WLqd4GhX6ZbM2+
bQXktOIp2+r9ft5+zdj+lOja6bV51P6HVxbg9K0x5B549FiXTcu6x9hcpQFyf3AP
WzA62QXk3gxO7jQn7aKKq+iQsKs9fYmbDN3SZFcxn5CELyFNICo9LnP3T8NqIG4T
uihAvjkWUpLfXx92wEk06N8XpaQv0aaxrS5zNGcqzw+ytK1xFvQZQeOMhHS+m2kk
Yc6BNzaRW1/0JiZvmCUEFbeSISMrmS+ZAEaV14J/hUHfzWQMHIdoHSBYQOBmV56J
GS6ikxZwrOnEqn+KgTAoKCI1YVf/iVTuTC44p7EI0Rl+8tRt6b7CxW/IishU105E
sBJbtFaTU/SAI+3MqLRoXlhw6k/2WJlH92Q2c/lRx4YwrJWgQthzQJHhvcli3ek+
BGR26CCeMgMvZm5dfx4EbT+TPPiyfG6UA8WMoYMLBuj+n+eKqkVQCH907GFoPOuQ
buOegv6ZbFVNSibdMvOV7thBIDB81bB4bhU37Plr9yC9o72Q3yzzLX0RqkGyMoqS
KFrEIi/iDi9m7+s12r31D0S9Xd0bVxSjGnQ0f77WLDETMgrO9jvEcvrCK6x1/okn
6Gq8TllyJZ9EbOf46amnxvEp1KidXCcTaiLfeDSJszqpZHF4BuIgpimHq2W6pY8z
p4Z6/DTx1VYJxM8GJ2TdEOU/Q4GfkTED4yGU+PhnzZbpxhHWTMoT4qbDB5XxDDdJ
ujnzMtTfzGkj6ZNj5ryF4RMOoNLT8IyzoVSf/1bpI9+kqJn73G2afRjEalK8iVit
4Nq7SPbH9eZtd59sYRGQXcP9OwS+qPmndIt+mY/aRpfefls5zMgIMGHx/ysfUi8f
rjvaxQNy3sBAzAfscE80g3XXqGTaMJYGsi8vqMYFtjaZy/Qk4oud6Iimdoz1ORpM
ZN7GJLDPTOBplVnLGct2VnaW3G+KQb8/hlwBZQNm+SqcZb2RCts6xezo4QzOYt5+
5MFLYxdla559sd68wDvpvmMDAnjfvifFRqpjZqB4nR/U4iEWosIrWn9Pc4kybgPV
YTR5dOIVPV21SRfAgBrioUCP12oDvkIJYPHH2Jo2CV/+1yI01gWLxSqHa1Wk0oJI
BPYIYVur5Rrll8uTHCjmEaOMz7Z7xUqsf4Fj2BdDCahSVssqg6ecxggUHFMKObgO
j3k24HEnyYfTb+ReO46BYhJhwBMwdqz9YnIxY/mufWouXDlFFXclyV7Ng2nzkaXz
2mu9UqWO83SWU8PVOHgAoX3LQnEHil0XUGcSevJqkSt+70seia6xR9hQ081orPQJ
HlmgBA4FKKF2YFOSu86SSSsgiz45WyXk5e/zUeC/vgBVcadzYvmh2bDqa2wKge5X
C6GHsZIBmWj49JRmqHlWI/+qwNkkCQhNW0N/psq3xdlHt6KB7p2P8nUbkAqem0If
uaeufltSZMt080fonud4wRmU+Mil9JhLJ0h7BSDlskgJvOPxhim0Y8W99ZCgOgAA
mUj00sF3EfrFIs0fjPnRYwczTdu4K6VOPnvod8AfqOewOVV+mdWpEVGHBOoaMUb3
g6m6R///eCefWVXd/xkG4JCI9xtZ5j9C4f/JuF7U7bXX10sCtzeYGPo+dcgaAUY2
XeXoT0AO2F6qfvV+EyuqArRVAkmnP8lZKozGLjURY/fkltBqrIxzHUt3qSzV5Rsg
uav3K9fPpU8FJKoc6hbBRS/cUZta3EVOIZyva4Vx74rQBoFi+2JGM+joIfxZhsZx
1249LwmCqkDVNjqRATZSG0OLDVsWeq2Pg7Jid1X4i9WIpy58AHk9+eDRB8K2dGcC
MIX5mSFUc7tuPgVoxBylrvTqP3ujWRrJCeoJRw+u5Jh6Qv37VSZDQ0kLrqkc19Ox
xyxZIibLHDw94KnKcc+nTFct3tTMLrE/TEEjjiFaMauNHcSBIWW4pNlJoUhl7JEv
/KTqKn6TqLMXrNWCvySpd5f9sz9/xy9l2afohE/jLFFnWupsOcwqnC5voX4jxRq1
j3XwYmUlwesQm6jYVQmDsMKtl1F5Uwyvl2l97nZhMifn4HFGj90/s+4vQ6UhJ/q0
x3udwntAzyWzOpAoQ9+jjqZEYIArpn+QY8fifUDIHPIsTgev6amf1JhM3Hw7XqyQ
lbsS+ywmtAsN15rXBAIC4N5AGnxYWvWA2HjQIcl/EY22HMTE6CBe+BulN5gDaxGO
XiALmQz32L78tfavIwHdOerEMw88yZdwIyJ+rU3mKpCGiqo9MfMov5bcLhgG6P5d
qUeon8nRDcjWzW0LClzYONN9x41wAp/B2adQ6VMXc2eZHrTYjH0DsELrITZEa11b
euIelzI0Z6lApSmBfWTBHSMMwa+6F0+El1xn3PcLOl5yxfVloZcSAYrFh0MvVO4F
niBcb9BjhAt8XqF55wZVk+GzJ86vv7AThn+737Sr6bpdfvSdCeDkAG5AbGEGPFSV
UUXXjLjPoqR1aCyPup82VMT6UplyC7xCMvobFVW/YeZFM5EKJg9D3FAKxkZ72+p/
Pc3dHb5fkRI8dtbP/kSf4JKs/ZyY4pCGcb5/OfXEUYeSrFay+CFu+plH4bbyxVtr
GcTeu0JgWJeyOLtb+D02pPoyJyrdh7ibA0lGRiaVU8B71OZjtoqwfhP9GIqo4Odz
rIlSHo9lghwU66dR9QP5nfTIFDqAOV+2054F5RN7e5tYFM6jRAsTPjzUd0b7l2Rx
L80dZpjcBN1MJczlzPsGv45HXPRg/Fu4mm2f0YbcJqnyDo3TBJmqMnQdZTeeF0DF
fGTmSh04dXvhtv0zMYNYaHjrVyNNQHSNsWmTi1B6vJOH8wBFAxj81Rkhu++z9PQD
SQl0PS+AioZjvJ+Kc50osi9AtWRXywhdCcbwgJ8S7jZELOp/n9xZ7AkejN5Qrwr+
ECm8ZvAXeTlYK0XZpz5qGfbfjW8xykb1n40zbRReesaBXgwakOKAsy+fxQD+BbRn
P/0PqyLnsH7dV+iI/kgluepLAip39nO4kJRUPsVsJgQE+nPnGXO+R6bUkiZ1IRFb
CM0LCTPmVocvTcNS2/X8HkuVa73QVBkmFjDJvbqlxm0c/LYlkVDUARVxlVO3qwaH
BU18+nd4nK5X7lphf71aAf5Rkq8z5ryya3v5dHsieygML/03UrfF9/iu7odjdynj
6J/HzXl6Tg625UqLP/iwEFgcCKSPT6hYXhdTF8+xcPoBf3jI8KrgoGFRldFsYxBO
w3LQqXl9PKuy9qfvJfF0/4JYTKqY/p1gPfGl1fWV2gIIvhPEakrYtTKKhzISpQbA
EzJBDpPxW5G3cBf1WhgLcgfsknt+9PNdDDtPaEJy/x8Kr2TXwHPUTRNjqCtynEvZ
VRp62yH89pEGJ0rt38kcn3vjGYYj0lMxYDj+DQhuz3Pw3/0ku7TJdTGBlWuZmZIz
0087DGpQJeyTAZZwdoe4OkHRk3z6tnbXDTUTLtkYBlklWJbpK2//MhX0mylS550W
oD/NWb3jfzPW0rEI7z8sC3plkSO4msIJ0iGQ/uUvqQfUWIaa3Fq7PNLcBOO/1TR7
bbZoydPwmxrhDzJRECo0GaTsQOFUsIdu7aCEulLmR9A23Fsowfsb0+YSJkuxhF1m
iVwbQDpb/TqYJdWL+Gys8VQ7OTEyafsWFowaBhOGafyn5gnogshliiGIgKh9Yq9g
o9hlAXdv2WD+TBHm1IqUWLCzTIqbpO5s0vYLLoKrzGe+4HK3gaLT4Jw7A4QIE8PL
9wEC7YVc04d86WLhVICNj8qnKGd98wGItukdcs02mzaC4Gp676vuUL6tbRf8A2dG
xRmKD8d5w5rwenFOFJuq5BeE8YlsdmllMzxlKEUdEfrHKamjNJ0OxtI4DDk7gIjT
4ZUuk0sM5x3yNOemOuDVa1v/bc8aLE6ru/CpXPSpKNOtVao5rOS+qn3FyxzHpHOR
pzAQSYpbSlpl4N56yVxtnUrv5zb9MCQuoCY48mnt9NAp+opI2qoLSyVZgAriF6CC
iLzlNLnoKg8ujxmIky0uHb5CqD90G6aj75Jqug8y7zmSRrlTDAmQdC2S4e3NSh0+
onRfvFVT7QyXm+qDFOCWoYB6tVFBaox36K72z7DAzjLP5dVjAhm40C2kjBY2lX4X
DICZqiJbu98rsvk+fsHv2iSy5hN2oo5kQRxGiO5AKUNCBnnApy9PhclbUXEyjOwq
H05hms6rT6tFrfUr8jLrZh+OgUippCZY7NAeLeyC+R36zep5Ewi3Ew57+G8LNsgt
ZH+G+KTMbLCOXcbeVwAoWgeHCK7VVQOJvXKonaZ9YXcSn6dsBXY7e2kyklAyXHR7
RqFpWZKH6PGraJw+E1ZPTOa8MEw8GKdeTb+wvnazoKCTLopMv1xpszV2R3W9Ybsi
cVj2/dEjjOpeDavjA40HjU3A6PUYeeQirldYzD+pDgdVgd/AU4D0oCXaGMZc3A9L
svBK9bu4lvBBqY4swr0XpjEZqjjxij8vAHKWPPRh9hcwuilnnlF2cvKjU5q/NohH
b/+O9mQaqW8Kcee2zNtXCCt5MKjB65POzxZOVrBZ9uzeK7CEKfpI+e+WR7V5ukqG
EbNSzIHjEuqq+4dUvuYh1JQRPQ5Vkeb8pv1tCBF0qBZ+Jds3rMkrAQnRQjjTPoKa
LICTHMz1F+Wej9UBG+9+5GLH3fFo5LUvs7moT5R+HfTEJwwvXYneiPEhTtNlfg+m
0Yp5E4VYe9BkzUQaEL/Ew1JrjFSbIR696iD/B2TdePcMZnYuM6dhalE2hDmI1ujZ
Lszfc+rMFWo8wcgUyi0mNR4RHT+eYAdoTvbMJ38pKyuHtdhfS+OKahyNbOkXOo29
9K5QTVGwINzL9PmaUXw+fwTiAgZDtvXH/PtdUKBO8A0qGU3T1NZYBTKUpRVNQay2
EzHS/otMOyHTrRHmqnCLsolwNJ7IBhv1Im/NiqBVmikbUOztJS5IN9J3WTJgG/JT
3vdmVy0+uaLjO++7H1eXZytK2ml9YHdxcRT7Kky0AaMW6E6NCdCtgtTxmd9hNIRC
YzgPjZCA7lrfF0ftAxCRJklBWc7t0kPphp7OUisJt+h+ANH7/uOl1oZPNIUeR6o8
PtLyeD9BNwZr0m8DVJjjKntVg1wz9arFTVx11Bf7zHjJu8uOyMaKNwR7TfPF7EAG
Yph6l+46rH5ytkUeVfrYL6ucLFdFVyRGcMPj1gApSsnWdq2SkheuMYEvAriZaGRt
QDGFHQ3Gm3+hTsNbyMBu08rZO4bsYSuSdFG2Hk52obWGK56wmV0VOVJZKNGMKtZB
tn8Chr2NpytA8nJ22NZKLcfIEpiXNzgc6sUAq0DcQgWtozr/FsAmHTu8XjjYsXlE
FbVQyVk8atioQ58b46TCzttVX2pXywDOtL+ggFwhzEcf8hWMRe6IjaYJyVZxrE+P
DXEQXZRFcSXn7gQ1J6NwxeaLoYKCF5sPU68FQX9c4pH19DxzxbFXQUJd5pT5Qdun
+rYSuu3PI6Q4CZGV7C/v1cQ3KMsQKCtbq0X76A8t8CtrlzJccOEvBFUfw48A8sLB
H0Bl9q44M/lOKhqfQSn2ZlsiqoHxCgKpV8aLQzzDTuWIAAFASgeGCcA+KwIfoisu
7I9CqAzG1SniEwYN0JcNdRASbt/eDJmsAuyMAbtufJcTaI+DBPG/PRE81NHlliyp
AFBy3rQfSYL11LooCw4sz7bb0UTIoJxJLCpczdtFWBwkhU83vcxsU59V0o0XMr1D
Oc5RCtfQoNVTnjsDEjqdo123jVWcV26SUyfdbqCuaQW+S25/biDEZOfo7WhSKU/S
CRyP5Mrwa9Xdm6NJYs8euXsoOmz/8Sgast7gtnHof4xR0KqUA9Bw+HtjoKW8KhEM
xYzVXSHTZPA+K6kBIRArV6RgW7QueK1Oe616ofnCcICwLmGxNU6j2YoKYKtPGh5u
/tcPIZpSt+zvv/YPNqgRDjNHvJ5OSBFfChUoe+TaNSnULZ8exkpFdctv89m41SCS
m38LocHcJfzGhRR6DHLTjSw9OPgYorPp62noTsFXoS4sC59ai/HPlWVHGUI0JUG0
H0Mjdb+CuyZ8PVFgmU4k3O3x2vQ3voBpMrQPQz7KQNdPQlFKxgb9oEeZnpc1VPK0
7s2Q9lzoow58ZTsrhG9JYM/bMfvxzRDAPM+K3UAH6upPU5IGD0ag4u6ggWSiWegq
Lc6CymrmAFWBdFhbj/1bDU3OJRpuL2+c6M97m/Z8VmPC9bjgjCDNg9UCxLLRPvBQ
/AuOk5H9zElz3YfkmHsnibrDluBfk4etJ6vID/lkixUlAy4GoIcWkWlDRjNyAXvP
Ftm1mW75nUQYTH8TezpW2NwgomtT5gXycgWR4LmVA6VgzeYKsK92QYgLzYEO5xAz
KG+Em8DOmSUNiOwJzkmMDsDFXsfOQJcZ6eKFy7VbvMBjI1/osH9D5uR8wZI/kMrY
dsR0Bw601w9Ci/PzswCNwxfcyupK2xBXEwyocIRdCeZfdsOlUfsvGVT9Y3zRDvcb
9aXF3Qtis8I7h3ioHFw6hywVxFPwqBaFMKYuMUIwnYr8Sv6+9rz4UwPYjiqNI29b
ApBbF+NYNlKtIkouYr8so3oYaQoMnB6aB+JB1Qfj3ZyUK63O9txS1q8PcjBFBjIj
0SXQdvJJL4UjHLv1+p63dl5EU4XjuBUbFIme1/y6y8gOktCrJX0srThJTDYUjPji
+bP6ZYP4eERDmnkzPlqKprFwo+nk67F3XDSQ5LF/uYzmGEGAF8ckPPjZc8sMU2hD
J4b8rpr9GU8TNnzpSXpV3ztsmfX9KvZXhNFacaImeT1sc4oyq5vMTk5D+VVnjJQa
fj5VSs9McquRSDDLHWX71ZfCE83lExeO3AItcJbtKEBvJlhw4LLkmHZsssY2yxoE
e9atcjL90LihEwIU4AjcELJ486gFdEXXu4FrHSadTNzOzK+GT9SfFZFw7XAR42Ol
0YuOlpx8wiKOnKmAeTYaT0jriOIIuFe3jEGXom8MGaP7oPsUJ0oajDseUr+mmYJN
glcI/nYMeDT72jcRUa3gVFW94eBAIqG8LBoFDjhIeSH030Mx8lOgHcq4Ax4Sl3PQ
mKBJ8MB42jcDSWAPLYngF7kJnQpIy7YZGWp8EzLWSwusy+kQot0EfmHNL7plQeiP
f7RqIZ721xAkgBG4uG0yOBs5FWSOaqpDhuIQapY/hha507MtWo9Anqqd0mbHff05
mTOe7aUbGYnVgRuYjbqPKqW/sND80Gc6DeVofwAvez4T3lTSg8RFF3dUxgcwynoj
2QUXF2l0Lgm3T4Ns4hzRD4MHNizpSi/Av5FyjSGdfE/DKjiTeFy6OoDufnb3LpI6
lfWSVuoksm6vLpPgc+iZt7zsfWaQdJk4Ieysl5jfKTJL9JFe1ac53sUEVkoYiRLl
7f/50HUrN5XJsyQxBK4RnT8nX2fxGu7S6P75p3tKK4v0z9tZrA9y7Yfbf0jcUDGD
jOI5IR3svTVAZqmyyacCUHn67ohOQhJDUrbnoCyEVLrn9oXdWq4+PJxrY7WuchXj
LNEW2s2pG+6b6ccJklG4LHKK+2/XD88pIRop0XDgTyFCKyCIBSDuZCsRF3Vn1Xya
/H9zvr+6EOhVHNVM2g/R+YOCxMUUrqgAm4gxpg93DnfmjHiseAoQ7pycyvmCxens
t6vDOJYkoahgVl1NHTtksX24PFd8OB8qNw5Cn6yNbPSJFi7L2qyyEBisXlxZyZi7
3OW9pyRDTfR+VKlEv+1hndxQ6C39mRQUwclVjXV8nXE0j5UzpM916XWKDe6MaOuc
BR+9KyIUgQDayXGXJpOcAIEa7oS78yeaNEZe4HP5QGCWscYQpdTQwa2giQ2eQbDP
kShwcYK/q7WZHWfoUT9V1jNFSlza1E+SYAce2Tyj11jV9H/jNo+Tl1fanr3v8mg5
bjZRX11w6DGoyHwOxDCcvNYMLaIBRfrZzmYMo5GZcZ2Z+jeySxLTtV9qSCUvD+bH
nPEsIaC1sr3xx90laNmIzpwrHx8k2qPrtXR2ZJ500QE5Mu12a4gntbyQH+ECu4CM
S9TsWsKcDN2ml1sp/K6mNGpLxOmnUWJw0x3JjdunwWGnd+txWC4fvg0/r6P0k33k
yEVAuskQM4cyCq/qfztfqAgm3j4RCdOJaOoaBqEml7Ou3lcmjWq80S+XHi73PpuV
jxeUjJ+txKirU7wicdgnvc+AMAAZ4xDpMTClTowfKDbWEbUcoAYmX4vx9czZGQYi
49X8tnWFPbRuvkT34siOCoK3Ibj7inJQ49Oc7utv4xgejqMLbnmwnV9qREPPHEUR
BmMmD6JTOJEi3d5DerteQ+PgKzfSq/Uwbd2SZ8/kaIpwBD8Jf3Hu2wqIFWODMzdJ
XlIX9k3zH04sJGJxGK0fTvvqYxrIRw+vV828y6RTwgsHuFePtoj6wSms8/uDPiyM
yfgYgNbFi4EHHA8VDmWZlyr4dpy8j0SGeCspHgAgfmOQpO+PdAEofxAp1onTTJle
DEbyv8HIVVwP8b1HUwh2Gty3RJ/gFYDZ9EdsHQ2OsnUESbF5xUYZkEwtdymi7LJK
g4VWppJzSqayc+rNRFF50DweBLEYdWG3HZkNdMOVIQyzooJSLRlf9hZUaDxh+E2M
qy039ZUlx/2SRaXpzB7cfo9swK6tdoUyHVJqhBvT6YHWxLjYGV9b7fgd4qM493JD
cWB52GQeMNUZkAcC1DmiJ5EUN1NogP459JrQufizmUaiuhvnquuMnubIQ0IRiNoQ
/Fk5HZSUFXs2VYs/gpfqjdv6L+ToEd5M+S5R3wN8jdnTxXRP+k+1kKbrEMm+8p//
O6guopf6zqMrAE0DjqDCOTTpEU3eofZVh34KGy0cG2RzWsSfOEVyqf9LSokPrEko
HG4aLczDjavmEdmcAnuTrbUe2X8UYLahxNuPJ4kfzatAcT3g3w2l650xj3m7t2qS
MEXYLwnRX8lD5zH/o5DXafN2KTM02MbZ32SybuHpPH5Y0Mh5QaUidOovQ6QO7CWo
OPuDP3t05jGF17pzAeUwOkVKtIxpZKDRwF0+BM/w4M9uKmZdP9+Q5xrt1xBimpww
6LtcrG62k6bozz4aGidR92lPTNU3R6vK+3zzi7WQ7sL861sQAvt1A00tru3Qpl2l
6C/PSCvIAzMOBinb9Tz9/NbNcZRzMjLRDzoaXrC6nXOo2biXXF3zpLVerioLCueS
OtVGo11Z+pAr6i8pFfJhHdyLsGnfQ2G1yWf962AOHlF6x2c5AMHyQixnE4hirvKk
JRpeI5wKVecbJFsinlLdyfymGOcJCDVyaOYj0VOkprjr/vK1ZijPZGRHnREODCaH
K/1p/jJAA4pJ7zv445pz7/InwVDXT7zUERR9Za0m5T4L3hc5KZZVRYBjgqXQnlxT
Q/Wd04ifTGv3xpBmnwRpM0CJfw5Ei+LtNYREKspjUMjjp/Ci1WDxNucP0g9h6cWU
uUVxgv/pjV8hUqzGL86QNAfjqq5HVOMJ6yHilp/nwh/neGL0/ldHc6o2Dqdqqm/R
W1d0i+ucVTQMi6H03exszpowdPJSW9sPMC5dXXhthBAfgh0yuC5AL1oo8uzaR3BA
fGiOOdE8k4Ze8Pe5ejrElEeAcA44h+RZWsSFHPES7Ud7qwl+v/p6aFu6TnhNGZzK
bf4h4GMtIleYoo03QZRNoKU/2MZgibdnxbGG6SleM/AOx6YSEdEt/kbtThBEN4N6
T0++WnTLB8G97uQI3LY3BFwjC2B67so6+FRwHcAj1mfBq+RnMp6Mhty7oSdmbNyD
8ISKV4sa3TnIwHHhRMVBcqCfKsS2B4oYTqlWM8+f8eDxPaI5eVpg+PFj/mo1XXrS
hRhMJXROPsSq/61JDVE789EOyos7Wt6uQzsGun45SeiEkzdUEWifgKPPCY/QWnv7
2hvd56zV8xrVqt2DDMhCW5aB95imWzUFo/7nxbxnk2o/whiimjij/VDc34Lo6ZTl
7FkE/A1rKhwWN5RSBWIBIJZo5ripZn2uEHIaRXKJpzi1dFkeCAoCWzkAjdATy+Ls
Ks74DZUQgxcPOWNHZ1bk+DW+WM5dzXfFbsjuJYQTQ/NrfO1e4+3A7SRCpkIKK2co
MAKbZKS2uJBenyiq87Fusz2GQVoC4ASmuK/REZEkB1tqwJekIh31y0RSCf0ciItf
1qxSNhDjmnrVEUaKhFRZlae+b2YN78jXx5fJdsUxNcgzWmep1lhcY/QY99fq029B
wTItW0WX4hurHMep/Xx35BhwnR/ytBNMInutwasHrWYyDk2nCUsdOWFpbaMDQvVV
8yS/utRjFx7amUEyQ1vJU6cOtFqDoiT7e0ELwzomN9/EPmOLPUrpPGczhKi4KPC3
S23fyzEDt1NtW6Y4Jd+x5bzvvtY0OsLrnvr9BzUgVUuUnoH5Eb38Qi1kb7TIFRw5
qRcLDxAVxPrEg2m7RLxwRL66YjJRnKkD4WOPLhFo600nO5afow8JJtfMyHqx3YuR
Bc17oPFy5itu5K741LWuLF0+D5e8Bi8cSOzY2IMBhR4eP9R1tWM2LWckgZHpK0+b
eqEv4qVECKJnY2vUEpjpkA6S4BYiH6a4TRcf9an7JX+jWTtlEEp1DBtec6yEER5f
xEiFDvWKk5vAOQQ8UcYbKlKGjcazsfRd/jb5PlGwytbIOahUrnnZv2jtWDXwId0Z
WSssvtldYoLs/kPCfl2vcWt0Mk90CzwAja/MJJQsnjw+Lp64RyDGbqhFBKcib5Nt
d2cbvqZn/WhaPuGaBD81tutHtxnoBXO2rHSpfnRHQXolKWbyhDR+BCbSutjFZqmZ
wPo2W3I9wH7CLhCkxtf/vxSITnkhfrJFUfEMENjywvVvKCRNTEcjWWGRpFHWZTEP
QKwHD9jXxTcT49ocUTa+XCua/RMdXlpQrIE4jdzJEcufngyu1kmjZI5bEeYca4tV
O5T1h+KXEz//x8dlp5wGdowrEdhxnx0ApO1Mxal1j787PdKmaXvWE5GO+gG2ybKW
U4Iw30lwUU7VoDrsKhqLPBMGXqDkY3/6me7jyUA1UZSZS28E4qoBMZ1fTkrQusXl
P0myx5HTo7WcJN/+/h0PBW5VgYXiw70Fp9GI/48v80z/yc6BgbuLL02sToiTbmda
OhiPZLwGbBH8zt7cM1/M9kqbeNOooAAEIeQbVDD3xJKPkpTXxfy7pVslrUh7Ykcm
xeoYTjFYlrBwmUl1wGfF0+tbsA0rhLxwu5nZqmDSdzW/SeM/qOU69DAvQPywHRVf
MEyoKQZt4jwSQhSTsJlaVbifBdU1TQemOqrYBT2jp2Fl/rPtnLW02/eGcHedRGu2
EZQDhN+FQKejTQDjDLIqKl6Fugcp/vgDUOHiW4GjJ3xvxbq2LBN9hmS+l1R82v74
CbQI0mBcbYkS79S0ioPm9jfu1OBBFFSPbn7OCj/KfETGVokK7+uvduq68yRFrast
MJUVWvfJCBYL3nZrHGi6idszbu0PsN3HQblR32RfwPvJVZDqzFtVDeDPWKWwlNpw
ShDzP1BxYL1ofvSfrg2SwwBbIuQbnQ+nQiIvZ0RuaPZeLmDvEYPoQThebsZNrbLc
j36sCr2Zm67ebAopl2APx6FA3ghKWRpKfMqf75odDtmOlMOhe875sdKpocAgir5Z
vFECw4eZJQhALTwcYmrYghVHU6EqfEEAKbK3pIBmvps1fCHg9UXnKirY7N9y6Vkj
M9mBeAHsPsj4hVega/wUaTGgk7mRGd1Tcw8flYj7W5RnqfWW/Q4cLYBGqJvf2zQO
ErwslJy4FSCbYt31SRXVpnh3I8nWIJtjteSd+hFjF9cdtEymvcE8Ns5JY/AkkCR2
lHPtV/0VkPVozQzFGZlheQ4Rd5jx5skydUnXwYC2gwucazB6j0+tufIC53Ekh6m3
YQ7zfPTdVyiSbbrzqWW4Gmn3iamyrDXGY6+EOYyDlowTFh4MnI8gSUDncjvgcQBb
MVS82GrdiSCGGZQHvmtuZ2kPdZre9a61FvDGhDhtZ8kbUgGL9LDxoVyl2rhqqQoV
aU8I9d2oFQlmBqeWBwjOM0hZaRCbEwAmGiMiv8VZadkPScVBg6AHaw+otj/CDBrA
GyIqzS44piI0HMHZxQKwWSe8uJZw5Qu/xKfEjuTAR/ucx6piSXGtDvtK+11UnFLs
LzGM+rp6azfKJvcuEvyU2s09/rxzKdORiw+K81uplm1zERaaolmc845a77ezZUxC
RAYN3HmyM6SmI4LF4LtSM1RrynH2u9Ma+jiev2lQNIokRMh1D9oNwRbWOjxCe2mQ
DSDHutLycJ+S2bvtqcM+/EaK4Bucvilua0twyftguyyTGCqetrWZ0Oy9pb2a7bUZ
/9rvWGCnlJuPDYetdqtX3CFgCex8HVtPP1cTFuDRSHVIoM7TSncv/6OjPqsp/30s
GZz+VVjyREAVSoi6TODRasr96OjN8Qo3V1mtP9j/Wju3bLtw6h3KE/ErUoDU5qHl
4KmOUjIM/aPgrH0yHrTgGrkGSs2d2Ocns9VtKAQglY788KSECJQorl87vLm8t+Gm
ZsFSi/jd0h4DBYKg9Ld+VDDV5X4iyvnZ02i8+AX/7JDFYxuSnzGA7CCR1G77KmoV
0dPkqQHDq5lbi2CTVOmXL1VJgDpvf0Rlt4U0IFQmqJmjwqRd/WinA3ZGGSZliyew
hHDdri8ZOmmn3/+d78kh6WAl0RIDo6LVlCSbs4gJy1wPKCP9KB1YEZ2QPLw5ebwY
0mdFW71/xaVtpqS4yo+qZnD1TYEunv9OM4OZaVK5Hq0PZAeG3DPNf5X/KH4HeDk5
1AMkQA9UngQ8hYiYfPZMfWNySdiPLidN4+e+AkXOLI9rN7m4b1BXQFFhWsnauGZo
KXNVTZ49emIb+u7RTYDQ62hCAcy9LaulYMGUN8n0+E9lGKK+kw8Kaahz10wsycdA
z6pUChu2tJ7hDz2zpUvCGhljbFhgGs7Nz/eV5157lkmdLivHW13LMiPdiVG03lEs
wKfX2p/TzNSaWhmfK31MtrBWpB1lkZqzOlKyo0BgAtBVMPD8clm/RtWMjxe4e539
9z/6J0Oqdi27oz2Cjnm9OvZ3fO/j4WmSsO6NXmVnAPP77xClT7+pIlzx3Q3lRIQ9
kcdbzif1i+qGDOQWJ3Z+cy2eKhk7pBObEcmHWp37cwsNKIjN9pSjc3j9AMMxSBhv
8tm6D5RABwut5oW+Vxo7tQcKVT0aoUKEI/cfAh0QfeS7SkQFbKw9V7HD6uFBMeh5
zDP0ETnc2+bTwmP1LMy7NUNwu7HUC6F+KxtfJYnGRqTb6GBQ7buKmc7PX1M8g+Sj
0yI6i8Qq8kk98GGe3TRkSMl+qs38FB38yYeM8B2uRjeuPj8FV8fK0oxe39Sqm8Zv
9HpW0yvH/dqUnJOdMTXWW3iwWOPuCsT4v/dPQHh/LLXXjIfNazJMl4XpJQgZJj5t
rL9e77YstbmTJuXkKSlXz8ymvjnZE+hs06MrtKn1f1x8HCvZ9Epph+B+bc/P8IdO
c/H8TRSw0igKRCQyym2WccHyZLwLR6Il4VmUlN/1QWJPyZXUnxFNoG2R2sVhR4pr
s+DlWVgvmdLgy4QXCkOriIDLbVBvBGvS5Gb3pCl53ZZVddSl58TnEmhdbDJ0tGp8
WGKnmIK2oEJ/d849TcfNrPIvqL4czsHmsJ1izEhy7vCou9hVw0aZLwjsnQ+pXpix
0X+J21vcVPaffWm/tC/u68YCy1xfeH6/UI6nymUDyQ7EDXnPINoQnQnCl7Dd+TSd
zGo6HJ75A6ksYmBVT6dbU+eZFNDFJEeaJ6JalsCp4VZRSz+hp3bbKheLd2zjw0YY
BvIMXI4M0IXLeKe3maTvrkkeU+4F2wnDoiETidOOFWz/xK2KsbRfHhlGEzCz9lql
spXlC2V+Zf73/9UKkNmOlwQhkSesapK7FaB/UO8j4wG18wn391GuSlgbJHghxg+f
03uQoM/jq7bNi2/iL3o4qAxZmJyPPO4BWXg6ypMq/qlcDwocoGWGB5CixAxUZlzF
MZC6D8EKkE1FR1jB3MfcXyTzU6ueraD+CZQekY4t6zFAc4mA79HXHx1xx198bvvG
b6xoxRryBvPyTBLDf9bf+KtryVD57VUYBJppVd/u1jHSIMvO8tRcF+1KQmCcxdhY
UOY8DqPyPZkU11etDSrqXbFw3+5UcrPxR+V1VKAYKZLHc7v7XMWfsWChOkwyi5tz
mIxOCKgkWcnYLcIdoxyoKOjhZd12qorXiZysd+Tp0IW7Ip9GLTny6PR1zdPb4qID
TWTykClgxd1HSqSJGReULlAN30L9+A8X+B+tDzCGUosaPkRAp8SJWtH457sRIPar
MZ7XeC6XuSHRGkVKARoinRcncWsFaZ5Z875A892onh6s4YITtGC9kPwym0XBBw+1
Z9LPnwWP4JGThcYQiVPsvOq5zEh4r79N74fQi90uPfXRB+DK5J0Ng6CnZ05zaSFr
Qf8oe39nIsXgXPJr3AarqxI6IAV+LaT46dM6e9LQ+M+L6ek+bfy2GNloV3HFiCQx
mA445SfAQEMNExQ4Wp5GKgOgnQJjtzB/fnm00vgbde5R5igWsPRYvrayV+OOMwtk
RheikBaF4XQGeAam0MtNk/5C0t8tXsYBuiKa2uEYH0kTsP7E+xZar+Fc0l7t2CYj
8saqbW8nlgoi1AlQroqAiZstG9d1yyvYs8hBANkD1ONV6bPxTFuLRE3R+SsbWSfN
e+mMNfMppKxldI9Nyt4unBq5KIm79ERHy/OFreAcZR4ehvaTFNDmEnlT9UPTHRF5
qc+B5xTyY3MOiPR9IJatdCRl0bmO7ANh/pGaIKSK4D9tfOD+Q1gAqa1teFJPNbfT
Sqx6TdowqBtFJqSgo4/u3z6mdDN1YcE6fFbetLTJDbjpsejRjs226CVuBeum7bSZ
qziPyTxQTfjLK5U5SF1+4O1GBlba716O+eUyy/y84EmGKTzTXO9NArVG4S8SjRiK
y4OKV2CLB9TsWprVgLDUjlJtS8pc166MBIzKYET8yLeBKcMan3r/JahLnAdEs4HF
6siqxsoZcAJcPKm1jF38Q7z/9r4S0tWetbbPxuVQouQoM0dil4jzbpjvpPnVj+cS
3w6zFgNVSNSgHkc1aFl/72T1xwuU0+rQNpQQP0xJ6yzuwYr4KTyIL68BQUA3sPLB
tsXI/0XvK4u0ZP9LY6edsal6gHr4/pbDCjPFi3wQA0/l7HpisACQ6nHOPaSAX3I2
RJ3ba4Ui6r/RYFFOTYpEgZdXOMrRKNZ/C4G/CZov/n5JnUpC7Moa01WrzBZu66JX
7fy0peLPu7q2O7xDNAJUsl/+eDcnP4PDl4k4JRwQSpHOI1tOWXPhKD6k/U61kRrY
5T/FhDyjdAEhyHZky/Bj/dCSiOUinwX3g64AF3ddyCGdTzGZC/d29E9XW81XPIYU
ViBJx7HgDEwLBhPFPQCXkFXQ4oPcrjKkNUGCbTP5hApSEAviOPQLOBq5qC8QJI7Y
QcZX9NcrMnX3AjCCLzSbpkozDaUCi0BHazUVrUjvnI2IeHsz1/uL69JqYChLXLb9
/fooIyWHIgt6/B9tRgsoa9/EvniC7xF3zcFRABwOAuHcP6hStrBW0peGdRiGkRN9
ySu0w90NrpwORcZX++I02U6b5UQVcCnILHJ2ZXC110lsW+57+UVfTIMgHplO8QCV
Na95Uvtw4cGAwxyN7epqIN64rkdwuf2u32S+j0/uNDyP+6EGlIW+cTGVZA1HNY9n
Ii+l16Us97OoBqM2u+J4Y5dvBqHgPmGqTajp///j0p4wYcWSERPMfm8olrJuvnTV
XMgcERXelXh3V7QbsCsGly4qoPodu2uU3dLHrWbxDTc0ED60iStkdNQI7a4Gycd/
fBKAK8NpJDsay1X+4ZYafSeeiBKpNUogc+Q6i4LAatCONK3EPuavFkp0iaOibr21
d4Tgiw8R77W5MjnHFA8uqRdbH7SncXJeQKPtENKykdJoElMmXk7eJ7aZONnNl7dM
AL2Q1owWmDku6x5VDFKE6/hcp7qAmGazeZ+ORkIfasi0HlvGGOigdZacUfliDdmg
Rkg536WWjXaNAK2ettrYVoid0tWrDVHk2HhDuRUu08WGuBGj2eLnkOD7qETh8DI4
J+w4FV/WN0CibTBbIxJIRGtBXh+KL2yTTcRXez/OBVpoRIHG+WG31OxKGvnvqKPz
D06mX7M8TmjQ2cJnbRFjBbiBSdEGRcCMEg8FJ1+MqGYkyohtY81DJ2koPZtVKogZ
hFSPnmRYO5ZXgaU0RLokjCZkM5f8upC/WCaNWSPrmmNqtqtL9mFI69obHfAl4Bta
PsqI9Dud9aD8q6JZ3fiaAFLIyaqr0pkA3ZIQn6VB1RrIHsorctgkX17Dk750NsgC
NC1ynzi36XBJDq9x2mxzGtFwtD2KXtR+9eNN2dKnwKubfxPJfzYQr78vxbJrXeEP
kKB/cUbWdqqUdYT7ybULHTuEVh9AW2u3eljwrN34BSJeFx/OcfruvXY3zBaTRKkc
8uChUAQJfWKA419i8sI2zMnxNimdNdpOzuaqx3Z73yVKmFOaGiSlITTiEZzGcZtY
chHrO8oiE3dIbveh94xRjGl+wEqYkXzyceQYeugwZRzVcvn70aeNi7qWLq6W5CK9
H5yItdKCEHPuWxf1uElL6wvGdpkqsMT2lohi4yZBukovb4gpFv4tNYVyM887ay4l
XmIwYGjbLKEAuHmKaBOpN0U2qD39IpN/eLlaadJf5n7ibdNmwBRHnw2rRXr+fUh6
6hceocoPE+lzGyPGSIz/S6KsYQeDY7Dc/a6/yS3mNyJUH+42RmP7w47ykpOo3fbA
3f4CM+OFcJCQMGx7W/e+h/S3nTGhIENoojR513pXqxEtlv7QrI6RGh6mZXDtklHg
cBgIAtPC4bpEzfH9wWY6KK3OAeWoSNUvBGoEgKb04ndZC4qPdzeL6dk6vJl+shuY
v6NVR+G4+1f9hzBRVCX0pyhAWfuCGOgyB36Yd3mge26BPAX8t4P1wyAFeawDrEMU
B8Crr3aM2rzivXUFpTnHDpuzuEQzbAX7RpxqKR46WOLQXX4Leqb4+DTju6eWotTn
e+I8jyNzZB//atcypQDqPmrQwvDutK2Lsit5NBKyqquK+dthb5t16v2bMxF3ln1n
/OiBJ8b0ovZ4oO7tjwWCiVv5Lyii9Afld39AfyFRiehy+uy///pKhZhTer+DqOiP
DV1vy13BK9KIvV3GUK04pqYp84yFbXLa7bLN7N6TdMpXyBXkw0z3UewIu7mVJcd+
p/GmGcGLo7uep70B9Yd4pKMjHP1mNvWXmh9RlxdqxrZ+lDaNdbnbgM+IQQYikga1
0wPRARdQOpDw8yON3udWvkx+0fuK7uuS07D8Jc85lnfn1e+/W6fzGt0P3Weyin8x
RaMdHR10Vzh0Zg0SWEj1p0XcWqLanKyOH1DDYTbhax/OgwOVihkx+qukc48Z4uxp
Tskla14G4JbODUNPnuMYTfBNgcLpDJRfFd67Ckbox9AXb/prC49IBuZYfL5JyEwr
got9+Z3ZAibfAR5i0hmaeCvUJs7y8NrglZF/V/0pTslVQPKToveB/tny5HwTFTZS
cQiEVTKnV61lJcSUFF2rU5ZhUhIvtAI2ygIT+J9IcRbILBH7KPNpEjSezwppXNdR
c2PGs+3LQO6SFNYq3KyrKHybJmv5060m9jmo4a/giKWQ7yykrV2t1Pccl9b37sJr
tr4vi/qrB8jW8fH4Oc0a8ot7wU9bNQKMpRQVdu+yuMY8CYf7xck2V4bLDaJmdQlE
lfOXBqXUH8ECUrcGGGUb15XZ/o5AJWzLziMP/mM/2Ly35zooDjIEpjXJYzl9ePmo
XmL9xms4IO6JjIiHjfZbbg1VXXlC0RVA1yTjPYIoYDPwEd6QC3uOgLSCtC5uevCg
ATyBfZgLfJYNxTsIOn8NjEY9Vuhs0jVeJxfbYREZwVojD+hKFATrWOR36DvOO1ba
FKN5YkxAF6IsQ9eW7GTjX+Jh+7UsYu5nf80JW1Vmrj0wMKrSiRhr3sjzZ76KTikz
HmrYB1G3Pja0b+RiMsEiPeXg2cEmECMbPHT33eBjI4jirBihInFra0ZAe6s0nzy5
riuk++t4LzrnAO404qsCGVomeamtrPNmeklEKgiG3bhx+MI59Y5iab/wf1fGcgQj
cKOqUu37VxeVmc1CjbslXmPe0sTJopZ/G0lJKnl3f29CoKF4Gnsm07PsuonTT3T5
++6eEOHPoc+LODjkev8/QtSPfqE2OPOFC/5yniU89Ew0PTLZmGJhht+WSyQaWKW1
rTQJyOgrYkZhBbjz/lAKvQmyKXxjgiVuv/go8tN0/BICUZnH9rbajNGEbUgABjNV
FlN9JxLDkHPV2/gHatV1jdEwQPj+KbLKDGCpSXD7XCtPzVjVw4Z0sWbqQ/0m7Oi8
BmXCYTBTXqZsu4A4Dzrf0VQFTdqexm9MG4zkWFezRvng/YfcAmN9/KnaNbvvzg0O
iLxqcxVZg8LRcUkpqHX9u6mzs6uhAJaBMmZu9cfM1cJdl0tGf6u+tMWMrKUfy3h4
X12MxR2Xrns5cYKYTuJbYR7Emcem2RzSW2epU4F5GLpk3ObzaPgx9myUiwBiUx8f
u26uEqQnfh80vMQbrA+1CpRd/V/I96XKEC3njcO1IjT7504wE4mrTGuqYqhiVCIk
ftynFtM5ChSwHQKMYqq+FRZKq8XT6WqqvbTsKZOhSYarQQId4oI6KmQesuNsELxN
lhuRxBMaXTtQt2XBoQlr5jXFk35xujIJC+2Ek907XhUIn+jjuWTACLx4CfGaJdPD
wusrbDO6ljlPc1dP/W9xS/a+fd+BPqlXQ5XTUtSne4AVNsrHnxTrltqjGwYP2Rlb
F/OvAWPHUPcn81krGXK7CT3MBJsS1BGQZNXY08NSy7zlsY9E671U7Chv69GniM9F
ygp0Hcwb1NNbqjCoHT3Y6/FlqKkLXlF1cW8tgIOcod7RHiZTKPqtqhCcH2+i60Xs
ejk5vvsMBhG40uDAUUO147A72hVuu8lRcx+CiK8IhOBc0dqBCaudo50hhNJKfdFg
T8LajosAhBvLV14rBMy2uaXBYmK+UKFfe+UZZQYuEByq92eYjMpSYyXPx18pV7iT
aDBLg+ciQOEd+Ucye7s4iIqwmoEMLf95GI7JWpN8X3oemMzx3wkOVxW2qR18BcEL
72bbaJ3v5HGsjvfW0XUapkN1pdBJCeP8Xd75JbVzLTk8l3SpE4FwQrNm0duZQlQ/
R50hEa6x0nx7FiYhDRv90MkZZC02DCz0j0vKLENGNn1AeV8HCZxg6rRjoKZzl559
1ATj3NiRyew5KEJhrUIWrzBR98zA9v6l3gcxIda/f4daTY/f7hh4vjAHind7TmM7
oeLvPfF0qbDcfKTIHcmwA+uQ9oM4gCVqzPBrawB0/7/kKMRRayrOPiKdRAPT4tBW
KhEmkX4pEXoBtqY/PZC/fOUdA4AhVX030Idfx1gs1Ob8nM3V+eiY8AGdLVPgvIPS
80wgQuuuV/11q+ArVtCddErOkscBKuecNtjUXgkYdGC2CYjx9R5iG1EZwNEJsUYY
NzkUQxhw+ZFnKBORPOFBSVDfR3+k3EilPs3cVz4bbQ4/2b3nPz8q1LLiZg1fPN0o
WIFLKd9vskIcM/t3ULh2oMlljjgcuR9qVdP+10NX2ahU/PVgKOt6xdv/gPYSE7AQ
QdWWtd3+S0K/UKReGhnqrGnLa6BvSi382UYbJseCeqOp3otTJGMI22veUvGq/TkB
CDJf8FhIuDPPLhdqgKerfyBswJDLjnyOJjj5HK5PqsQWQ6vlZL7IG29CvIE23PbS
9HfQFbeG9j4LVwbOqVenFKF5bYY01J8bvYUbyH+UyiDsV9Y4dRa1GFfNV6KTY1d9
wE3llGHxmoVu9ktKzT0O5xqPyiSODQBpvfbw0AG2833VGqa3xb880Fv131lk48vF
bUMPw2nXZPJgsFfk+izFVIQVxXN1SVvIB3ieQ8srzOSyK5eJzBWQzgUtV4q95B9v
EElYZw9kRUxMZuClRUUg++OG2PoVFMi6/Ubv3VHGJk8kJUOWf6dat+MRt3WzbmiK
SwbIOGq4TN0TRKo8rv0JOH6S6uRlrG9hhH2FX0S4G092y/RQ7DZqkAerBLD/Qk97
EtKnhXd/UK6IPIWkl1MfTswMHPFuS+xhKL3whb1ESPLDK1/VppMfzSZQAHKK/QnV
N2MlQdSvFamIA0HK3brR8db5iiZI7SqFF/bEqdL0lAOF+WcQSLR/f5HlsX3lJ9Pa
jUN6gD26ZXyJcE0//4ICAIk4p1YzZltji5ABOeFSgsobHlCdHomneRJ5Czun9/S3
GJx5OArmpqhigIt0HLXazcfiyu1gzeMV5opcnbKuAAafXJ4C0WmtHoMhTYBGYnxz
ITSsh0BH0lNnnoHGpLyCRuoC/GPz6Z3iVhFRcNvcxbaNJ9vIUFnN1egD5G5MeOUh
3vIiEWLthfV6qbJeWCOVgvBcDHZAAROinDFFaaK/4z5tDtLP/iuWaj+0RqjQhK10
erwiMxQA7IK5Jnlk1SO+Ay65oDg3CXGvMEI4aiC8FAsBgSsLGXTGE44rz3fL7UBw
5mlF25CTa/pCIHzxxxQ9VN6bS3EX1IUWO400irZtmxTtZK5OXjDfEdMfzb0rOK+B
S71RI3KPA7ACAQa0ehMbwoQOQu9vvHy2Lnsul59SDmKZGtWrmnlWcrEPkmydlWvL
Djv2nUOVSSDIAnIIKdBxqPy6W9T/3XdCX7cwvuHxF6QTeXf1z6upQtjED4fASj9T
ogbOQxxEZ8MXR+rY4ai6676JaTmxpAA2VfZDbnlyO1BxOcDApK6dioanQ6p+Zltf
MT/25k8BI4C8D5mTOAxEt75+WYU8REkFbNlr4eXEYfd+HZlLKZVxiyeB841HaxXY
SmHGeewsW12L5oG8AHaGqftmZETnW9LF8loE2Yvaq90qn1eb8Hq1qAiwryGGz8/a
pXXUh4m4yF99UqFP/Ue6RSQPDP1R3/VdBfGTQEftMq3mSCHlEUgD9eDFgwy28nSp
65y7r7IYUdFhr0GvFfWxRBUZzjD6cI31sEf6ZTCOcXoqme0X+QHMlZNvxJAypPEe
h5lPlJQcVW6k1VyvQc+oEQUFFQ558FI+rDioRUjzHy9EmERjy9GtmeYwBo6s+QoE
+9OeRMDF6BFoD6S19FoObPrMkRtCKQwesvWdyDufV47PSTH8ryjIRpNLsyOqKV3n
wHS5PdiLSOQh0R46V8YOrGCd+DoEbQfNE/O+CXk/8/JLe9Hi9q5yJlwwvM+eU4L6
kd3M5GDQkc8+7IPDK2sjuM+Z8iUJzBbVUur7zf1NiVLhC2h6jzSHgRsl/4Zjncde
i92Obd+6vrlGjMOB85xFYay7zOjzbkG5aemT6bKuhitrkFIghhVfYcMeEI5zwcOU
ujct0Dp6x3sRu2w4rdPEqD+567+o31SCtXgLjl2bzo9vOn3Poza9d2txXJWPQw7j
CFgeYtzOy86X4u9jxVV8JHg4XvMQtKIJcX5yI9x5iT/4H/8bMizbMDWLTU2iuGx+
DoqWxenPCWyYp84HFOK3CXM7BeF+xeIvj5aAM0K+1qwcCZ3uHICVsSAV0LJ1DsdJ
6ZSR7undvOygEq3KBEkMFUAdqAYOVxGTD6ysWwYBYH+E/eBj6G0hIkwy+UHyas2U
UfnL3GrzuJC4YLTohr+ApzYc9LFkOit/c4JhS52rbbC+eXTmJzwcnNVonmYJhdnT
fZQofeYDWUoU6NImo+PNFD9kchKX3UvJyC7OYHl3wbN54Gh8GT9FCVY74+AKTYbu
6/K7sCdGm97zu2F6J3sDN94cNZlY0ODhoo124DxgNVGt10APSu0agGIgsfaJ1t/U
qCs+E8TuBpPY8y5eeJ8hGpXDxcnaPN7OXn/lJFpuczas7tYfMJiUWGuNwuMPXebn
1MpvW3txlAcqhh5rYzaAZY8goRLqhRwSdc3dYZvENZhzduc/pGpHmdWUfRognnYh
jdqjUpGb4pQ8DIQpqUt1asmZDqZV6aFs7xlNe4n5QGiOqvqCcj6lKjX7Cx9IqIMh
VfbrTVhZRIfhI5+9QnMLm4O/wBTM/CG7lVMSTsOnYLiU6jdQB1TLoxdRvxo1fItU
uelk0aBI1z/K+3QRZZkc1fWgJlIXfY1PfYcgdNZB14gb3OBdyoteQjTs9eJPgLmA
svo8K8GFbdHNcdiH+njBC87pjCXxIe6XYaZKYe+QA4u9PkJ0ARfOnH4wSYK+kd08
r+UhGBcbHkQxPWUvDTFFzpO88k+htMXUeX5YOM2xpb7zNg4IS5u6DQ9I4L5Pa5NO
gQ2WgRCfqj5vFrysq8KDcDcD18plXMjtMOZL7m2vp9qq+pd+0tHxpupvC/OtSyes
5+vikiDuWmdO4NTUZakzgVkabczNlceBtzwSnU1ifl2HJ1DYc1o7uXuj40QjgOiv
zVVrJb1vGKFRxsc5i1dIGbx7+EZ6sz2F0sQw7Z4jMCgZs1UZr+/cnTJHm5yVWIgV
PsyXbZ66Nb+y5GWe++WJ7q9LWorE8isknyLxMn+aahuiI/rjQ3/rWOrcYGtl4ucq
HwX3dSN7WWGuwuOz6sV1QyFtfFA2ZJZX1S2z8dYevsg9uqJ4GcpOD8wN1SZUF7HD
hEGnIYHF4SCMG61djQgf/DbxDv/CUhHUT4af+pFFZR9mFFCkFbtJbqGHH3HDOU90
ebh8OrR7797wLguhn7pxk7aPLBkPqw+XT1vulxd9HND8/iQBfwORLjVbjVD93EEa
ytby9afulR8CpbhOWz8ql9OMJAYjtHENRaq6oe+C2oq8F2ahI9ykX7Af8+H0lS9Y
pCqMg02LYo7vg0QewQ2GBB7339Iq7v/6V3MktgpJUQ9jLpna8ewcwMqO85nwzohy
QGrvxJG2vke+wRenNT3ywVuEpHRZe2pkyF00L4R3FhKTtbjx3HYYr1RFwW4rQDtM
6lo2ox47hYEqIIIRPlBX/0JdRLUCB1YTkBhcYKtX0wdsTYrYZ8gbjmXf57B2JPvE
IRNZR/d6IQjyzrM6/KT6A0X2PnjQ5yZK81WX5+xstyjfSjlw4I11GFU5kMajPF1E
Be6Ra945/CymF7MgEOMVW+XxCashmY6xgXWnif9DCpc5nGEXl2zEWw2EdztxgcHJ
5IOJW2gAD8m/3M372q3iZsTOuW4p6Q+R/Srt1iQVx5OcPePsOxhec3FIVnF2YnFI
HfK0C847c0BNy1nhPjIvs6OPcoKOu4l7DUaXQ2879ZYJQytf0NEniij66qvnF/+f
/2tc4cAZjWvQexy+GocXe1QxB6SgEYRjleJ2eBM6rLNQs3ERlkvpQEkwVHW76jB9
EqlqsIFmnGZncURdyP65PP2coLlXZtDzdQPxuIfpA52qELH8e3+9Oza9t1IT6gsh
DCp4wQnt+043I5QGwW7bzAqZLedC1XTQQGgOJ2XC2Uv7Pqqpa2jnpvymfzixX7n5
jUY5NjWSjkoTZB8CvIDPuKCyPiTMoQaYgJW0qdGMPHSPqF4Vtt43RlbfkxKlQOkb
/qITXpxBjRnztfXpRoWnj5TVNxtE5NO5vX56Ke3Pl7sPx6unxR3Rxd1+i3Ujko/Q
tibZhvsfiJ+dzpxg6kONWBoSwBKiPKU9hLAUsInQQKHtQOIagIxG6+v6ikEM27pz
XOlDwbPpe1N0nKps6jiWEM9ItIfbYlY9MAu/bnJXmGkxUgue2oekmi7tp6EgvihK
DC5yz+ZbZlBFoKicCJnOp0+TRIlfoVI9aDDZCMjKsXlUOegbpb2L3FcHl6ScgRFI
AWEzpeWxiOyeI46ViRsdp5yfsDx/p9jZsGASEBg4VgFj22U05SYZesFCTKZbQLS+
fE+Ueb/6dvxXyIZQudn72kcaTYBM5pjfHPLW6J5ryTBWqybAyf2LmCW1pUeK+VK+
Fs4VakuznjEXC9jKu8OmZJ2DD380242L5B9Jhz32onPFR8oq4gJCgwAqLlIAVgnC
EvhDQl1q6aM8SEdCDoExURSvO7HlENNQmgdh8Wz/Rpt8DGC9EQnuRbci7jUjAY+C
BlS9+oIqcjb+OozhMJFCNiGVQ5Cbb5VPdVmBU3DcgipEaEvgtfkrmtb0oRxM2Z/y
yVuzhtJjeRN68GkLkxz4SQLivAtME/LpPtP19+osv1GZ2sYN2gWcxF9es3+M+con
ndWLhz8q6TD0b6uecFhP5EmdqlUh1BJMSDQ0L30scuVf42/GcuWTAUZokzaq2rJL
GBX1y7pKBV6h0UYQYfB/Vw9x+UrtA6lTG+OWlmqISUJXhVo3XZbYeOw4tIa+FGs2
hlGTgeaZfDy8YxHC1fVfXrV9DR1hl/YOPZzVA6NgPTFV/HSIvnEBUKbLMXQvwUVq
bmBHrzLLvOtKTHavquWCHMtTe+c1m9BMzJcVv0ihDENWzDFDVBZTqi8wMEUk5cww
6aRjQovmSK2YclDpCioYwWk9WTSzNRsLSzAtC9X0o+iTm13cPb/DYFbcCnKuAIF9
nh9mEZPLycXqk15HcT7unZ2P0HzoZFAZi6tOLHDLFTYKAyGBBJX1/P611dVYjmAu
RC3aVSFs8RXlt9EpdrKAXEkxdI294EBa0XW6XjSnHE+CJYmoAU3l/0UozbxCWyc9
5lGtd4svXM/2J+1qegaV6edDXsd2xx8LN35ZB59tuNfaqIzzJum5tVF08uPC0nti
PLIc0PfgeMe1CHlv3MAfwYIHfkKF3UWZF3HpVPCLKMevrveUjCx1QaEP7p8Do+YM
SqoZ7cloy0DKBcywwHKdWvCxejUrWQ6Xp+gunAnLOXxyxGWA11WD7hUUpTtgNLZj
l6ob0LdN/D0/h6ctdSiT2WxghVq0MiSERpHsrTwnYMl0yIEAYLNOGgPcx61NS012
Pex2ANHEUe7y2fHxUbMmDQVypMAUd1SF+AcSD246vvpJ5DyGhU88lakJPBmRwvqR
1gEcDNXoPUzaI+X0nh7vxuQdOJLp+SxlZ5XZk91k3A26ACLbfTZs/f97rVHF2mVM
q7O8p+UwHkK40Cj4ibxb8lMcLWT7+Z4y1N1CccOGKgmTh3OUKRSfmJWqVzMBM/a/
U7W6yswigzMDKZR5LVL96jsYjhB8sM1UZpIen0DiHVbXeXUtkO4V+rE0ieQqdKw1
/QTwqDN9/GQiY9Oh+t5dJAaYhlGMSUHdI/5DAqcshwGJHiElbnqGvUiasgedg/ec
V+XR5Gpg2BKfoxxaz1L7TgBDw9SVqcXO0+OgM+kE807ePGVBI4I3z8mby6ppfVLo
4p2GoErseXalsplaKcDFjKlREW5AiIsV3+jKqCTUMdgqKShhMsCVfTrglPqm9AhY
QhIzBh6RTMKCZoCWAqsOEOUj8FWkETWlbin2YD6kwqeDep5WTBOiljv6tE6lQLFy
FhyzITCvdS0TR0v6ALmgmJJbp/3w79P1gib39Su0FLI5FmiTMW7R2QRRtyx9Wluv
VHYr6ZXTphdvbxHKbRbgCuk0+vnHjZBxIxZ+gHUFyIIJylgk160bn4Od91NgjS5G
qXH7eNJ+VNUqTENEq5K6ewPNpdGVymmc4+v/0w9xBdLqMHtcGh2RiNGmJvDjbowZ
304TAZgHVQvRd8p/lUQbVElcuLqqL3NW6rdkOGxVxHr+wQbKh+qb2854SiAE7hQP
5L/fGuYfdS8IBNownRQVPL7kbQDhqgMyzcNHitRiq0MT6gWkC8E014GYT0WTNPlT
XytNTDQBD7xASJZnNJRoHDFj2A0E+6OmkGtjbLBC3xiCLCvKS8aBXDq5MqPXXV44
TSv4IYppqait7tJVlcFtW3c6zFlpSxvh06EAKINJliRbSgJMy9LWvz8lXPMbG4f+
AaRq54wl4w49cMVqYv/V1FnLme88LXPBJzXZ5g6A3Df/jMowqolc6FZy9eqNsMVc
152oY0Ye8FHqwMm8aZRsYSM13y0j5nyctO/5VQ1UThmoGdK7qzrGlrlzArno6MqG
TOrCFDg0jQ+12cNp1BYTynXH0q3SZWVdlGJm6mrjTWYFeYvvFV28Gmergc9DndRS
FKR4LYvGrKRGiIQhTLyjF1NvSuDfDzNnpgVeQUITJvIx3vmEDU1IsD5BWI2OZMm1
ZDiTSRlXj6UwCc97XJ3NOrDH27O+gQz2gC7sc27pqpzr/CL1MTOV7HeCOJ4uW5e6
Y1d/jU8V5hzL56hnA+GMDxLNzNffjEXPjd0F+u52ev4ChtEkPbGUWA2dhj41PqPa
+MB6MJEa+u5nsnXwkKmzwv1DPPHrInVbTLvdmpxNJBNgVxCeNhHK4vwtOhQ9DChW
dSjN1OjhjH/fynj4CvnZ4O6cN+w2UX22j3js0LUOTECJwcQd6NGH7vlR424ZxE0W
zLsqYSucejwqOg7auJzJ4Au5i/Tk6nY3Tu9f2CLsEzYBWP1PdG+XwWnlS1ekBv+9
LTQovp/CPi1e1XdR1oyUtE13GVvVd6wo3W5jqIzuqbeWmEBMaLccK1ak1it33Nof
ZwLN65Sxx3rHu7kjZrq4xUis5u5opJn++apmvwan5L788870ZX+VlDNtRRhot6XD
UEZigpttvwFHR5dUdn89Tuy6qBZtaTN5goIiwsOibPA+zG1ThtEfp97G/a3ZOGsg
GQlN+6JuKcfSFbSl8Tg6CNGWRx0ko/sPDKcriIIKq7V/D4Jt5grCmeQc64h83LBw
j9OzJ/ox8hyAlO9G+ttJ4uHhXBFjbPJ32uzotB+y8bpyRQ1Brx9SsI/xSkIw+ED3
1gjQBHVw9IdWTq8vuYWVA7YnMMisn/s/qmtHXD0o7e16ZRN5Tgnw53nnHd2oD/IZ
N0S+NWHcrNK0Y6Frb17Fsbfkly7w3aSct0/6AtR8kDzmzma39cd6VGMnLF6s401m
NHDEbi4tKxGmd10nRsw8DBwdojAbAcYkRCNsWGyTXmazcdXOBqjtQicQ7R+sVE4Y
+L+qxNQgor7ovAHuGvA/TT2ZtT8d0gUDfDu6/OspHZiqzaas2tjZl5u2aj1lpmYj
Kpp1JRPcHULnH4auPndAh+wgquJdiEoonnHiT3aYpsOx+dF2Me7o953UQq+oplVl
KgM08dVnLjT/acwWhp7B6mTIbteNgMf2mD01A02YBsyqOzO8WhrqaC3YmFWDXszK
Ggspsx0/buTRsUyfie5xoMDRI6NPKs/mWY6YfqAy1TF5xJ0dzaqTv86ZfanD6ZoL
gXeQ4s9IDyn4IqYUVjOvFv4UavYZd8/Im3u117o3DJQqPq2Y88BzvOEjhsIoxoar
UI920iep8NmNOFA/lQe1adzUY7jnQS97RXOnn6IXjutEpbZCpc4M0H9Jx5/vOlFn
2Q0DerKXL0ofZSS+i6eDjZPDnMZSXtvPbJHeLoafAUS0ek8SudR5WCAL8cU9d02n
qT2Sr0nLxYznuS0Qy/mHHVhsxlBpsM7SvmonMBLibHnU3KnT4H73mcMdD3XGHlFh
U9Pr1YV3U5pqcvbmZuEPqqu01uBVMNtRXxZFLTHzo3sprfI5RIfosy4FYR1ki2X7
ESZ3H/OycCG/illkegzorzs9LAssIvmptAxwRLnnb93FpGf0A0F4FCCsoY4YAdcT
O6qKIZb5w9+jVkc1n4PHrbynKMEnexQF/IDgRCb4GBFFI63Oum1ULJMCvn3EuldM
OprRb+5viCkN65qcyf5yr4cCZPWDaEMA6c6kL+p7qmmMDtPQ43ZyPcigfJIGN9E9
B1FHb+2GLPkLWj2VaDqrBqH5LPYiuZgBgfFRd/oJ2SBtNuY3zh6ms0RkFoyZ42B+
unajVnm3Ifqz//GEy30Lt4O/RHxWzcEoo0q3CvRxdYRN8Yp5zNspH9AfZQGS5waV
C522pJgBHhUUNQ4VK5JoJsuiZTuz6J4Iqjx9rfllXTfvFcy5OPbVvoO52w0WkjI/
Oe/rhtDCqTbESIwBmCFFGT8oLX7M6r7wzvgvixlKN3+Wnu0LkKuXxk5Tgv1n5YbK
J0hV5OnLafcYfEFv0YDVtTQ9oKYMXv8992SOPKCjH/VFuCCe5lHcXVlbXy9NlZqz
NTA8ICTanXHu0/a3BSriLtXuTUP3y1D2i1QCBbt8NfPhYAz9z8w0ZSWHSfg+cXBG
3Hg4zbDjquDirjzQ0/VjIprDA8XNDG0NXY0gxlbMr15lOlvzEn8UM4adMDbZNE8C
LlZ2UWXukVFUi37Li4tJCyplh3Fwy3bbXt/5PHDnuZJACJmoAu3WKS9tI2pxyL64
ck84Ehfhn44JngABsJX05DTknipourPJtfLZQogEd3v+iwpQAAK3vEkny6jF3sPy
KddT0hwGlhQkanS40jzJE1mnhTDmZG+2kcC/t1ri60UWbwW/N5Ml1asvnxccvdw6
86uAPKxdFATlIdjzegp/NyAjhqf0Ivteqg9st+MXz8bryMeB7d/eUjljmdmQ6I4j
J+/yIsmL26RgWi//w0vqKEFhwJRzXkb7uzRSrWBRyB9Y/s9cdbA+Ogu8zD8vY3iG
v+1A1JlrujS6O+gv6WF/R09dm89UBkGUlrJMFk5kDtaQACnIzvIN1ThCeFmkWuea
1S+G1eJ1gG+bQKA64UD/PuI2dLAF60i5ceBr3ZPodT5irLA80AWpWRpDwuDj8zZQ
0HaWw0hjx1YAGcF1UKDZcyjr8gd3ayrEd5p6GPA/AVqyx9IJAl3lAC9qM+jqLc1I
RxFYgOdXmCW6p3Veo/3b0NY2Dw3XknjiI/4FO6zWswRquEf6LDDCv3umo7IZlrx0
nivhdgTepBqbq++8GgOZiPPsQa0e5nL6IRe0R0Z6H/ZN+o0QwTt7NenTERxhPXkF
dHkPqel2od2aSFtxvJ6lRhX8GcnLgI6lMTf499DPQZy1m1aYQHEL65zNNEiwIkc+
2t8y+E3pcfMCcD4iFt8lfcKAz1ojTPp2K+6mMLThd/oNgaFGj9dof6189DukAMP9
cO673Pb2h7IDbL7qneQLziUcGahw7Jt4LFeRt9vSc41e9zX5170oYkkkwV7B6lJ+
mb6nGrm56e6kB3G2i2B0gdPNSM5quDVJdWTOezzsJcFioH1tK4YmHAFTah18qlGP
fZT7b9o2ywhjL1vqEM8FNmi6nPRHtse4NElBBmXaPjK9S/WAzhmeiCnwQ78/MZWb
78oO6F+kpsz2hU78bM5xYksomU62aZznmJXZ6N+2H4ShBrtVpnq6X3uaWHXLDidQ
WXCg1TGsS0phCwZoMCRNRcJspD3fjlMibx7gj9YRt9SHJy5hwLuB4auVk/C8o1/E
aS+XbzqIa8AsxyWN0K7FCg0e45ptfLE0FuQQt+KwV+XZXdSSmdFpTRYYUDjO4TMZ
rDZRgKpMMookxuCUHYtdAQWCYDwFuakjvQTg2cqqhx4vmC9DM0YBC+sR7873mIMg
RzWWRAjQNiLtA+YB+4Og2fHL9/qUaNREoWJaSDoLejDZz3q7EzRO540wMzfbWs/a
ihiEiEMkzaMJNkKo22yfGOKZ1CG4l3V2hnXtjGxZC0te8gptvSbYGU3y4/HMjH0I
PRR4y9Co1NA9k7PtEGVoKEQmTqWe2wK+ijUV5WbGYrUsIpXvfpsDWifnQdWFQGQv
0EaUsCMNnWloi9kOcHkWqeRbsQ7ia78ayBJ43FIxOguCLOK61BLIDL/Mr+9WehtJ
t1aBgiN0hBwRqxctmpSBmTn+E57WpNatVArahx8TNYNChW4M0Ais1UJXb2DgkIWp
5SZ6QuEMlkHnKBzrFnprDJCg4YeOI/qZCePLOqitTRMJrY8p8Piw2bZK4kIGnO2E
K4WwjjxcSy9lEKM2kT1XjBpHUtmZuiZXOwP879CIT3ulGrZg8XW1EZLsw2RLZel3
f//BN0rlE6b74KgRG8nXeJxtOoap6fxEgYAI4gEMMViq5L4ZbkqP5mk2BDLTYYaq
tOrMNl3CH5KUyn0XBtgWzYsUKnnBh/SoFC3cXa3SZgJWHYMP0/bmgIU6Gft7V86f
51GM2nBUWsPrYDp7imRq/MDsy11Bi+D9UNu3jhSUgsVKuruaJ0rQWH7FdEQdd99+
7veEy/ytf+5DN18s1QWFrj12epI+3sH0Ct8jxmB2GWtG5OL3eDagELlSSU/MYfWu
7G5zaEofr9p87yAeu2NIKF9/0xbizQ62FGU+ndRHpEwwqjt2kxXmAyWLWxJGZkpe
wgwIoB+AqQetrO+dP6OMgZoP9XV5XslGLZtA9+oDShIvJ+hGzeGbQobi4rC1bq9/
vHcqD6O3z1vWizqqr4Rt1uaT9/28psngry+S4xobKJSbJqnaLqeCALOOr5tJIfP+
K/isk2PSf+MffSEhIbS/T+5Ty8WCYpsAUh9Os4bkx9pCKuQm5r/bo2JOZ1DfWdbc
0/fPs5z+ZdFfdf1DNTJHMIUgIZ6V17Beri0bHvZhohBkHAypa2ryjTznDnB7lz5+
wZzgfA1vB9OVaXBk9ajwvpjGAKMulwv+LNdbkGjXwOfPmy4TB17RW2InNdQWSD3n
MscEDGfzVzgL4JInbt7Yno/xAVL+1umW71s0FUtKrrPoZ/59YA9zonuRPWq23gFk
3Z5YNOkKB/JkzwNrDUexryBhZyLfGU+WTFd6DI24Va7pc2S44T1Ywf/fb0pcVmNP
Fi0UCFEXpNyiCtiIgTH9USbBu+HqhW67hwvoNfoLncS3ckJyyjNAwAFNk6hafegF
Hojt9AtrnQAGkhTih55byoiymYc2SaPw6txYqY8Nno0F6MFsaSCQgTjaOAVnWa5k
1/1na5m8VklOK+Mqz5KZ4abtVEAPjd18SNucyt4Fc8WKTKk2tSuILTeBH2A8lVWr
q/msP74v/JGsiue3hdpRr5vMbZLoQnHk334plNKugJuaWtd5FHUqX02aveWaE7Z7
+LAhl6ZuL5Q0EiEof6dJnUSUgruhLmBLmriUoGGiiLCK9RMn17QR4hJel8R5JZfY
IgeL4+XGNXx/wboIqq5rPXXelI7assv9LXt62pMTWtjnSHtr5LsHLwR5DMzvWkoQ
TiYqzaJZqsscKmy0gkrkXcxSohEYSfGDXMkfWI2KB3IoBukxQe95MJSjc2XrKJ19
QkKWJODSdQvua7vXh29VH6kQh/IryE0zRIAuYLzwHotkZvbwHyxe4dxhVdz9N6pI
cmlSmKTN63bqY7IpMBxrDubBxXv2a8QZuZg+RZAcpJgbZvlmDzehRniKhc7lsEDK
Ud4cwPHFc8+3BXhAbjUA7aOExZ+UjF8GS33KFoYrBEFjE7BI2IiVC1X+rK6dMdOx
GLGyXwsvmSJAnRHZPDUYpeWjs3fG9xD6//pmr4+0SCo5eFY8K2j7pRwz7wdZOddm
P7o8bVDgWKBf3fedFhxDpPw/lS2KbnoU3dz9K1Kc5lpKN1cvXn+ySA3gUxDFVrq9
IHdk58+cLS7RvIyKr6KOIfi8ZEfFRwVMNmwm8Wp2hj3JxmBwLuHGyTCwwJxjSq/V
+HStSCFv7iDqMVeAGzTXq6AfrZ+IBha8KXqPBJAZRcSqyXdiSEmvYMS84KxL5lN3
dLGZ0yAB5xIhuR17f/Cz4lJCV3ON6j6Iy6Vr+hcWMvsCPCDT/bvymhYkzmF2dMTH
hRWHc+KIq62pl90GVlRvRmju+QzRkds8RbF962j226aGTuNrZjGaJsKWdpLafybm
0hsj2BEvcZ/OKmCSNca2k108Nf9M8+nKArT1dM50aTjTftgicMYHexHhfrqDCVKx
jnAqtVeWVfVR5mjhw7c8RFBLnH1vRFSiEHteVez1lXZiQk4FLJUn5TqFelS3W8LM
LqEMicdj+17mclN0INLxOXc+86UvReFrwgm96tDZPf3k5BWnS5zqW6ffMsFAvfa/
bG1NlIsmCpOdk+EzVaKVyXrxlt45wfN3a9Rw1f5wa0aZnGSUlpmYAKV07nKkLr0X
z0ioZQ5uz4Xm1Gg6g1vlD8IKML4Ak+CCDHFBZmFqUbpRv7zZZ4EawmbT1SmvOhdh
pDurLrh0MQ0S1IQvekiEm7pBoVup4twMEjp/QySSwUT6ZB7ql/97SMIvgoR6F7RT
FOpwJgwBZ2LTaeRTJS9NfPTV4JoysmQKUqdwP6IgH8pndWCUXuWiamfiMZfBsWLV
5Fb5l3BlPKkBjxxko/u9rRzuRinC8qlpAM22Zhm5l1t01vTKYj1ZUVDDts5OQJjB
lst1WcFnn9FHgH6Xayg4n3Y1aJBNZXwA+WY9Fbwxle5atJFhifRdG6nkTlIhdhSi
OpPAiCl+NIZrNt2WRSJ7glR6xbTJlN5UKhHOG1vLkhNoZyyg9Ybxx15v9XCSxRak
aL15K52f+TTl9I9jA0sMz/bEGdWWc0BPcan1qVscOGp4FeaIPFy78Jphq5Wt3eyR
2vKBuD5aEW5+F50sCUFgjiUBDL5uwq+74VNj5qmfWcbeUhKFrDKlJnKStxGjOSQc
bGNSx/O3rFPHYU3eGMGIIjjlqRDhaqwgTFA1dZS5pgc7JF1xR75BOmVfjkaPOPbn
IIa+MP7jeAO6O52PHb5mlrwqldGIxiapXC63TD1SnnmU/xMdBDuRb2rIohIN4D5V
BJRzz5DPrk645IUkqAoFoV1/nHwKOZeefuiNwUaBZAnXUd+rEfnbdUEBTDT4SE4p
3fO8Hh5U8QP/U4EZXJ/4wESQjqveOx40dEQ7plo9TTDR3oXvKZ05jtOwGf17rjbc
RDjYESUcYlQ3mdJu/kQaYEwpFS+VRgplxnWkVw0TKA/NvFMvLMQSze9S3qIxDOex
gdcTQKvude/9pXYw8Jf3qRja6PpVr5wuMuKO9k5CIO1K4c62xReUWlvycDkDj1C0
C8/H4jL7Css99qkFa18wpTd8jbeITiRsboOIKOpc3zegZ6hsbAiXw2E7W17rIkUc
fXgpVYVUtzJjoqaL/p453mXUxqiKxKNV7moNFPD6tDcR5FcFccMRMe6B+w2fNGKJ
jH7GzQ9xs0m3tat81YvZzacDcAQC7cxBWheEe9Zr0FAgCTvHZtiSZa3IH1dZmwmq
/I59KGmcA7m7KLreYqsCn/49/zln+n3B+WzzeA87W+EYNfZIdKFrkc0Tyka5SVPz
0ALrSg8FtHL8xIRuNLjbkd9snLYkvPXbKJtklfWrSBRfmM6qBF9I33QLa/Uz2Afn
iS1Cg5ScV/LQigLCnqOamFEP32LNIn5wQdwKetKn80lBAiPit0lGuQ1ImBzHY++P
+wU9aWwK2Nw3vZNp7i/sb99StHPSoSAbG5Jq2nvsxTBemZa3fhO6X7dBt1mQf1Io
tvNR9wJac6Ym0K0X2ZmTVUh8l2nBtL99zAim3ctL3Y4hSgPix5rnPGe7cS+XOUEG
mj3ymMgw1GKy/v0E8b1SKlbyrvrIn+D7GxBshP1xhrFo5uwGh9ASJ+xUuSlvjz6t
516IFXsjEEfR4SOFN4/6JojSdqbOK/1/AGBLrJyHUihNJGznvdTZRJRCr6gWVAqK
v7cJ8+r0xGgUIx3zBfX+/+KKMGbwDmuqBd0z61d/rSqYbEV+yzikrvCL7Xi9A4nS
t/5G6riSEfNzhaUd0w8AzVhLW16eur69KNojFr/Tit6gssePxbTzhirtmsjedaA5
x6oewYflFVrXenEN6vVuCL8JnOGRfFjb4TDLvppRcuxXWAht0aQ7MQsjpLx/GPDV
QEYvRA6AV5hStkQaeZ428axnf7uZRXua/Ni/hUVdsWvmAKDxV84kfXnt2r0eIBnJ
EwAH8L3dSy3bYLFunKdWZi3g5CjfrXq0/kMJoG8XllTM2DIPbwY70co2qsnwBsrq
zDPVqPRu/3tMFyfsn03RiDLR6oeXE2sM1VWtCGQWiBI+IhVFBK5ffuJ2N6+gt1dC
4RtDsWd7vyI/nMr97p0LVlSjEmJ0CDL825+Lalvdmjp9sKT4ps5tiOFjCS5ABdIO
tZ7slghqkO9RVSQaIsKnIyUutsYMXxU9OQVP2pFWMpnGp3hdMcnuLQY5aiAabPU7
PzMjPhhD0AUC5WwCoht3ZiytKGjb0Hkx7qu8lBaGg1/6Do8M3Z/YRsooyvE6/YRR
RCpCy48SnRYE78x8jm9+8bKtIzMemBkfWJoG7G30bW8DfOYq6t7xPyMYFKga5DrW
YS/YgMnjueoFsXS1kJLJGEYQx37qfYNjhycfHBKgNFLRBscQG0RswUHISMGthcwe
r33ZZuOZlfyxDdRJm9xdkGbTkX0tbEz5k9sM1wGJnxhSVVRuWNbJVOg4AcRJEr48
y8/2HSTOjktvNCUiTWm20SBdPF3y57vFCDQWB2NUgJ6MxjoHq0omPBQ2WCkBpI/T
kPe2tUhi+wim+/zgA1W3z3IBHAi8lTeKqH0WITPZU4Wjv35FZRpjKWwytGAjeRPY
A8v2DtfMW0UQgYsqefdbZIqX0MtJxlgC6CtCLXP1fz8UT6XgqaFAlwxyu5id7WnQ
aE8IE6QEMFkTuaWcWC7UeUptloBaAmNns9ft7WLwwNhkSDh7OdBWHbeEOanMv5e/
Mpvn/gPOuxaixY5wwfpxJgSkLVU/LhO5RdiA5wFmICPi1dZaDZdTrr0j5weaMvRb
zX9aWuQEZvR9cU2e6o58Ex7jxdl5ssiq/VTwVL/fsMrhvIc10AZOB3GU3UpVtD6p
coNstpNZF1cmvkq41nrSCCla5tKw0rEDZJMdhDhs3fo6D+3hOnkRALSQPWlbqlfW
d0PiwYapAnO1lNpAR4FILTfDabzDlnSoxiDTX7fSpvP8gtIS0Sr+mZA05JMJKVbB
d9mGZnicmIrSVaMecz+VW/gDjOtrHehQii/uCrs3TuXgohn5xX9mbtnBbzyGUs1r
C0a5ZJpwvPSv41E3iX3qD5UExAvGVmGVr6Wg6cdOYoyZnc7pncHnoCu3OFtEEmeH
xCJbizb+rOS/oQv7sXdqkKro2TeKcVHPMe/ugNypFxBsS8R4CPHZ4NwCr5JrrGIi
W66vT4U7U4eAwPR8Ir0KpTptd/FiPxk65Wp14BW5G/wNadPkUs2dIjLlrXHlM3fn
/8saMIp6CYTtrmbKZO5NHUoD2f8E32SdgfTopNzFD5PtuCD+E5RwYitT1rGpfBvS
gPLf5ivzZACy7wsf3PFE4gRFEvRFAwSm3j1HhWr97J61ajqNXDFwlImV/YncqN06
DYupHkBAbPDV/+NyfHp74FjqOhNv4SYYZGjUhhKb4XPghLEEBq0BJ/p7ge+bClPD
RGc9bSvKQWA7rtaGvohhM/VwE1VOK65gl2YyK1eA8C/wqt74pC1I9xxsCas6hXmc
5p2fkSGbeCT5QbhSV+gk415Px29ve35hGINFAaTgqYEgjkSqJf3JBUWZIApyyncS
43Rx9nyqceToja3HQB+XHalMcnkW9S1pCGFzKPN4uONKEOdZdjhfrgPH8PNH4loy
cOYaW52hdAuJIgNS95ZrQsp698rF7pY/i3e/M565jzBYySrm8oh3uTusHlt4AAeo
8hqbXmzMdiG+JKMFcIqCycOkcav9sZ5c8epxxYTimHpmI8y3Z0O8XawqjTDCgIJI
IOFCAP0hDHOaBjZPZEMiuBHX5XiliEyQFSsJ+yP8jij1SfSG2vEQl0byBYq66AHN
zoGP/EU4hRScoeIEECVKS7UFOF0J4p+Tf6ycMphxTFy2iMJoXabS8N8Z1rhC1SBU
6+bj33IzkiKCQJTqEES3oNfLkU88rWyIhRp9lChAVq88WixKUqAz2WwdE3lgWjRb
gS/liGOVig5w6xwPGIckNqBLlgaFFBHiIjrMTIyBGBRmti9xg4JrcygZCSGZtIkW
TI5G6WumEM13TaY3TjR6NY0Gg2YVoSGlyPHSHHZIpq/scBEm7s91URqlFlrevFA0
tt327A58vmMBQANCaG9Y2vM3zekDJiIsRSynWU/qb/0g5F8DSoUOFr5Ou9i2McQ9
1UpzODps9z16jI0rsdBYIaowTH1DdRkJMZ/d+4qQSm4Ftoq7AMfIv6v6bmqJvDy9
9h6JLfVj11OXC/me6du31o5RGXP3hnyaXbRGdVJJ3qpFpSlSKq8iyDFHvzo6+QEO
cmKBCT1QMrx/rv+h39fQrxK3CXudRI06qM23licGGSNW40PbWsNaaGFXL6ABz0Z0
SmTqu2eo0aAmyf3KFR25CLMzcUJyguh5uiz3/LSPwL/q9dBuCBK5BWRWPdvpSJi0
SuQTR9uHHGLeFflm3Ue7nGAoh9jFTZzi2GqB9Yh8NPFjFY4xC4h5Nj/7+riSIGAV
v3SBojkOxymsZK/s6B8rmhXjxWGOuowO+iAklCo2KXe/WO2rha29AFBJliN6LmRt
SA7AooQUu3E35DO3qik6jhj+SunLRAc3SGTYV3cMfNxfCBFLrA6HRAnz7JMzd7I2
c2GGTEdc1u2jELpDX3aVItrRbDhrnIPgQu4dWH0TSKSj937oSkJCsUbhHi0nLGUs
sI5SYUM4ns5VCI1VXDvBpSJyf4HdovSBqYq3yvbnLh/EZVugAzKyDtAu3dqckbCt
UZvlBQSnxr6EVq8qEAakp4c28lt2FcpgU4G2v/Tb9TY+HZ5Zgins5efRb2veRIwL
oFzqSPqia4wGwz++JVVz/iwXB/pSN8LYWsGBaGiHdaYEdzeifj7sNmW1TUfJ4v1D
cnT01ITCRdM2/TGPEyiR6aXvvuu6j49ReHh/KgfKoeUCuJYXWFuUXd1RsePVK4h2
U+vboIKedjCcxZYrAXh8ZCyVjpRvlcu3AuOokdHtTJddzpUF9Y4IY/3sQ4BA8tAe
UtRXmshWTtXWvAWlZKiXlvy2Sk3cRa5QtzeQHLm9f3a0N6dBzLXnZURrzvHMVcEv
OYUAh3zKARrs/zl+/q1ltay89k9poLmlcofaHoOAn3GIV5CJ1Imm3virY+Nl2c8L
2MNWFbAweZ81PaNokSf4FZsR28vM2KawdHspDga3/b7WUxzmqtNkz9hihXBWmWvt
dxe63r0GeRweU2f6ERnGeuFI0P/3w6JX1RCwc1AFp16PjL2GylS3GUlki5579oTu
Gc7Ov+yIUxUzIQjR76amJFo6dztA1YPzV1CDBzjqnDbrQMUPWqDwPIJPTbDuwNrc
R85GSLKR1F76OlFyKmPyjwv/Zjcse+5gd1dDswJFPHqSyFnSB7Gl4665riD62u9e
mgN7RkxBhnJ8twLCsRPpUQCEIfoFhhq27vmTd/CLuXnzgcdVwbNWIgUIyAsaDpKD
KGz8UGjcVGXQs6eENjYJtEPBVwM29vZrLl8d4sJI6rtHlC3vGi49wWoANCnwiaZ3
YHADld40p8AqzbKEeW4TvZWjFZQd2DPl9vyJ3YsPcLxhRz8DxK03iLcC+mAwop3g
FVfj1v0FEKJd2us7C3Fu8rsmpDyQ9mGyHLEQ/FApEay0t2299k7hHDA5RUF8dWXj
xa7Oyfcyd6Bf2Un5DO76gGaCZZ4wB2dAYUfb+1D48UdQW3+gKXPSxf5eI2PBFilo
W0Ea7DgHFr/iUMzqXaDet5MtaLv7iEnf6Q1GApWEhKnTL6FFNF0h2n3uKb4Ct7IS
Px0NfqPAOMObbuGB5HK3WHE5xN8fhCSFPhWKJOJvyA59/TK9bYvg3m6frMktn8rc
oVdzHC8RvdBO3BCsvpKTASWFzU1PiTrpueAgjjBy+VGzDJ4pf4zd/SWjXXP2JyHI
PgC/2ageXiPNhqaGfVzykJqEq9aP4zF3uzd3OgHaC/bZdtFFmBMiVxo3Ndbm2npH
62asud/weIZ+S36x68HQ1eusy5bTqofDPjhDGTz0vrHjlSnEOMVtrewCSeLBtFTG
k2yYmhfKXzeiKSMvbPpoDj7SbyWtt8PV7H3OzpMtfycA19nYv7KkqOD0rIbIRl3+
AkxGCuVUv6w/5yLWORpkVaztThF9x3Be7CoTVaSu7g3QoF1lUqrqZIbtmGXvzdJ9
FAC+0YoG1xD3eu/mgnlLuEBPsHm+iXiGtFUOVxYdcsvYUuTFrtMstDLQwXBp9Gj+
qfScjr4wvNwytXSGDd4WfdmbCXMY3sGzSXIHb7zXTX8TB37o6BaAl7um3zEVpzQM
GDGf81T63cPRcamc+B6zVk+RhggSzlxwmjGVEa21+5N9Vr/DFfl+2Q1TU2jq8z98
L5bIV7+kHtUfe4x520N9eqvHa9PdXHtFi05tXerrDUmpHALI/yAPu9ZUqtTQh1Vm
+ifpoJcHm87Aybny/PFsYrvcIMNlvf6NZlSxrx50KGjT0mBKRkBrpEc+KG4SXa8z
zBCxf8B9e3xyDlt9FKDbRfjpFTl/wtLVjDUYojCKfH5cPsHbtNi84cHnW4oAPEtE
xbfDfzW8I4JiC5J3nDyaKCTdb3smHzX583KZzHJH5dpz1xLzxpyYRKbguez7RddC
qQLAbQATviVOoVnmwoqc392L6CvPplZE/WBb5VUfidX+Gv8cdTspIaDZAyf69P0z
LY+IdgYhsz4294/OkwxBuxxlVsNFGo4rKATxjyDLxUWZsQvYOLamrTrQW0kqfXJJ
lNUViBf+cg3qe0PPxTGR4sle3JB9hN2AE6dC9V/hnmIZUB3fBB41GIkyT2eMyKnF
DVdLu4s/N77Sla5v8z7QwFWYFFqnMHm+xyAPuNmjSzFRTDnDO/s5N2qEuMQQIJ4g
TmGSkFvKKIb9nwSQYvHIKqfat257RhwW5FM6+SLI123sj26IOKdrA9buKn5STRrp
AZ/7couS5tVPR/SOQ//SXud25Laxd1rdtxiVcoGg+wOH1NFzutwnMONHEzlmm7/D
h1MOCTG5REDKBYUvWR3hoRgYSD7wF5TBDE4X9Ja8U5tqfJxNnl+epM5vOpvtZz6b
0dr5etizcDi9WEAlZwyaH4nnxmsASENyDuwJkD364cOMxLwOdNk412vZkXpFc6r5
bjvN1RqOR4M9yTzf9VHHXMjc6JiDACZCUxx9mgzyKCov0M0ACfCChPeoVVor+QBX
DvZAjfxh7+sRCVOqfV/MeyF3mIgCF2N3ZMXqwLQRAkZm3MyIwFOPTVb2l3neCbQk
SI0y5Nb+mSgKHPlvZy13Ky1ALgt1/wmdWIoxAd55qVZAXuaIUtjs7nvbZI2ks9sO
ACvFTVYBqWVMzE+IwoiZgFpGOFtmFfTDNg/zy2D88fQdiAcTBBwJztoVbZpANitl
rNoqzH1imFv4NN0JZ0i6ugVgfEBZlQEs6kh4WYi/r7vTQVcdQTYC/EAMc7hGaxoT
E+L2OPEJ0qW52Y6EN/bME1iRmVaH5pxnQHvaI+lLJavMpGGTdrhAqYd/XkDKHP68
SclEMrCwghwzIvtooeDECDWNwH+2ZBpns27xwR1vW5r8+FzGM5LT9cjGQCFk0jh0
Zi72iy5tM18+szYlKZ8kvsdrBb+HV9TkWcxg7r2wSdKH++wbb7fTSYoFXwg8eAY1
MIGsvqT07nlHJy+MGgqIzImIYO5UV7f31/S7/aB5hv4YmQvO7uXI/ocwDfMSXCtc
IXfQAgyPnwn27pqWBG0xPrPWDpYmuuLgFre7B39d9p55TNdogfDRZpDuHQ2gjVLY
pRh/W2E0nYYVGh9wG+veU1iMnRm3fSYrsHYAM4yzO1z4LVIY+6Zg/bF32X/0ncJN
/wtqyIkzlRsdf+STxkLyyEmSG9JSiC466lr0mCPrF7ohjZq77laPdSW7jbfK0mUQ
PBizQKf4PFaVEWGNpoGGqm9OsZlj4QuQ/wiHmoTgbYgUU877uwbsJcpPnpk1wg2R
G8ktXFgtSvhypNJr7yd/1J+xxsGbTVJpqRZim0y9qCq3bf1W6VkSSvD2hVh8QTda
yQMs6CSreNzCbL6LWbagOY18TDg5tCvQQm04Ogq1WC8Se71rRHYw+ZTYCoNI5GGt
ZVey+LGEvthx/h6XlWHwSn1kVw+7S0m5OMw94RD5h8OnPB9alm5+7TjN8AIg+69h
RVAZmZ+e04EGeX96YobKxduNUKtLOjGdjAXwE2IlkwBuQn6eNTlbYaLXx9IY0wpn
KSN+B2rRiDbait4gwhIoRbLcZT89DImTe/fKyyKRu+PosUxTtIBqxw7iNaTMVBFu
RAjebkpWa1jCrIrA+RlqtIzjVEbuaMKAzb8AOk4PcZ6ZRh+e08NqCU418qVhbaA3
AN5Ip/pm/gTtSp7M/FsC7tkragzGrxjB+xDEykRLD+h1R0wL77nwiBq9+HjaENWS
WRchSJO9PFbu8pSgorzJoeeAqqWcYCXD0EZvDf+BPks2SMAdrtO5IwXaTd45VWWM
+mVGEbem+Opixi7//JkhjSkN4xdETgeLgZYJFqRmxxmAEge1cDHO0iRXvlnVoVkD
Gn9sDQI+CEMIc9lTmJ742zgGdgar0xE+rzXcPEfxh/I1aRNl2ZxGNTynBTtHNSCf
q0oX2Q6jmbcJp6FRWiskwPELBSihg0Enuz45kODcj3VFOL9dYc2HgpZO1hAED5ry
vlJNC3iFjc2DsoccXIWM87pvpU08dvPICehrcbanLxRkoY3q7quCLVX208Lweip1
bYgyQUsxiBIDvbTVcnAy/t+qbQgr/73UASgLDva0p7yopRE88PzBS+wtaHLmrpbc
5l77WTGwMTPQ//r/Zhn0TwbVqWQTUBy7Spja9zpxOFNe0ojLbYYFt/ZBfxuwOeHS
QAPOALY2ICBGxkv764HFmTYxbRYT6jj7YWACQxA8LjiV8q/QZkArP2FVjAz9RkY8
6zsYdAxDnluJFBEJqOAqavXCV+3BvAdGfzFHgvmhf3bBL2upwbgzilri6XXbc2Fv
Y7Vog7DwsIIChTU/998ymKQDMe5J0Lm0ZoHKIzm/O8vsXwmRxkj6ErlLQHqoy2pd
qWvz7wi5pMP0kNwKAb1F6CFIWUKbAbr41mRtJCaC2e48yl2nnWTp/PEuwjgARPSE
OH+U09WDWSv4q+F63UveEm8eKNrLabL4D4c0bjZariphP2fXyW134eANTlISKMTs
RIxcr/k7nji5rxmZNgReywgKRy9G+AFGAIXhHyXzmpGz+WuQRrOLyYLnzyffV3v2
YKe55Nz23vF7+t5euwTksILeMdirP676t6SyK2tKLhmcu1/lZE7FaP7F3vFwsrAk
Du7nIvyZA0IoijsWBevfz3T91tlzfpf0s2olCUoOxY0c1QzE/+SgpmpDSRc33VJi
361X/W/9L3Ce1JCKNocc8/JGKg6JDv14oDmvjEFKTF6awqYNvXbeTk2TjPsoOA8i
AueIyy7vC5+tVjrV8jBd+Aro2XxrHsi2duokyJ85fF7TrhOekof3rwlS27ViZeoq
UiI0GzFFyRgQoUeAVIjBrpGPNtAd7XD4shbIjuBjNxurRdJM57L8o87t57sNDQVV
V/NA+3UlzOSLZXAHemJE2iWcOdKSoQrnOy+moU42iog2/WlsJ6zsG42XnlbKdWpr
A4KzqWOY1rmFMwv9KcddEv2JyHaBToaIM0ryNSpOY5Y7A+SqQKQh4l+2Yph4uBZ0
gHzwPBJ1xLkT4RSpSL8Ii0fBOjr5IYC2d3yznnmHA4WO2jDAkGClHzVHlXrs37Jw
9dem1XiSgLOG/f3hB8TMx7cGdGTYVKCvxJCqG8o2rHilIYxAZLcElrQxFNFL4Kgu
qiiUhOv1mMELMru9uuwDXLchraVpi46GnI4VYihFqIw4znqfsB8P2jxpc7Xy6Srt
3vyYbQuhxm6ARaQTBmw5nsSnVNiZurHOOvebUTarqNb/Exa0JvMql2ANLkHTVH0r
lNnTQE8rteDWCI7dEiiVNuqb7e3xSN1svjtE0zV3dY3eGQDbAX4QyCpr5JghPVXu
WbftciRN5B7J6b9whJ2QksNNXO1RYgtBCu4oXLUL0Sptfu8+INKE343cgRJIAr3H
6Wl9AWDdp/Hyg0ys8wX0ZkghAd094tyDjIunHTCdoqkl8kfIWEhIXQhAEYeGaSLu
mtIZ4Q/r2I27zxZkhNBFh3n18kOBVViqDQ3weUsHGHFOsCi04NCY6rnMLbDHbeWB
gcXet7y8tNrZgbNcuPc+4fedd/U1CGbiXoIaL0ZqyiOFxFMqGa8MTGgYaMnrRLg5
xfucjtON3F5Z6hQwoHoj2qfKl4ENVO99wmQUcm0Z2okC5mX2rJU34JvOAR79ic7n
Yk1C4ZMrbqXZHAQAa6tOaFKuj1TMF2qnWq992eiqEU8tVSIKt+v0p7/t1xAETNWK
mKLyy2eWu0jUVAiD0GhZ661Fn+T6Cv27n/EIOWsrsbEZV8ERyH8N+KdK8+emKo9x
klU+vy7GXSgJpZaX2/H1QfTARjlz8OsUJSaWnEMzau88cUi/xx9hdv760XrZHnv6
M6jrw0uP20RjPwVEPHmER6nVwbvzroDS190gl9y31gDaCmCxaMYbLDZxP15+0jWb
mo4XNEV+zMULacQKr/SBDTgVHYx0Zh6Pe1R8tsclwsrabMnKfYdC9lVjXY6QRQWt
Hff1Hkxi13Rib7iwlm1OOXn496oj1410WB3TQZLbvcgL6W4x0XRQajOzCLArhpQC
TabYJeodGIMmMOwCt5Yy0aJGWu6+jzowRZB9gpRfOq5wp6kVh199zizwa+HaI0uE
BICIHSn1n3FOI6Uhnq4yNKYp3h+5hITwRMwWHXoZWvU7czwuHvAOXPBGEwIw8FUT
dPRxpAbZMduARVV6Uh7+4wwzN34SavztZmIingp0YtEJkvJ1486nnRHfS9v1MSUv
byXRxR05HSMKc+QtgtiyuWSO8OUrI8RYEKoq670K+E10l4wleYUre346Ftcsi6NF
F6n9YrAIBWfLdWuj8ougN+Npa0IDdbAJPtZmY+hCWXjtOhxlHlMhoV+EO/ho93Ft
Y6OOtGj99bx++9iOn0XccmuyHOyYi4wqDsk2UIH9hMwGsuOfDPVETXR1ft8ZNoPt
RthDbAMP1oGLhRQh7otgJTpL/cOiSiPchGh3nDX71zUUmV+Rvaux83UcKwJpk4LY
H7abxHFtktyHWQMUY3MbYaO6ySqlH1bPNmFHcHh3KnnPn9wqfGzjlDgbzwXqyucl
wMR70Q+61WpBiesL/7QfhQ4tWlHS8JykOt17vKqU6zrVBiW5nsg528PAqg6UnyRN
1OJbdYUHAoqW7O3/dMVejqq80l3UixVxk3i6VvlKiNQ2mobAN9s7RpMkWrvzFMic
lIDmGzfuQL1q7M9muhFir1koq3n2ygCUeUcp1QtWA7Ts7ZSp9GrkikgGdsPfth5f
rhST43ek0KSgNvFA0OmK/NBmOr0L4xxlIQeQhRvFGYgcsbPHhtNYrv6D/jNkZrVr
CM2axDW5gLI8fC44QTx9tMcvlNPLaU977FtNxOBsZkByejq38WO9FGcryzALmf1s
ABpUZu3eM9W7ysNq1YTM7DdHP5RDTJdKdVmSgYIxVLdVQA1cbcJJUx9FLVs0vpXy
vhMZSk7duIbH5vUFkH+xmrU6H5owTcFZ2wzHJ6ABMaJYLyWOCiRy2DfU0al+Sl3o
2BBrHizr3pdNdzu2T+ThljSUYjD3PimPfkqWcXTF+msqsyw+MsK0bn6wTGKQCFU8
ygdl2j4+ccmG18dimHa6xXWhNcMxCOXvir/AcGqJNonhgV7LrUA9CbzwV1oLNBUz
XGXABRVo7BXjJVKu+K4QR7S4tThdbQCMmwKtm7aWv84DQ6zAkwYIgjx2fNyhNYHb
b8cnrlV/IvexUWQOwEkxuf3zmPV7lleT8qpb08kcikYzoWATPLAyKqCX1yQ7rRRS
DaszyHOpigaM307fRct3vcTomVEufsIsaU3zaxVVC/ZIIxRu37OhHrxzUi3e+CsW
PqleWhZ1Ju23HM6fh12/cexNrFADJXn28LRwPXYAnydJjtO3VAL4YSVV7SoCCIDR
saw7IhzpSac6nJ78INCotqIVFnxgKvvF0+ZlCwTmusChMN8HS/WaeaRZao+zLDYZ
1DK7dyQTi6rn9HSTLPHrwbsknQf+lJRrXlZIoNVlZ4FoEm8aVuWfZLtXbx/R+Q7c
WfcmHphitB5niXi76JbtIidGkm9nq+EEl+R01wkeE4ePaZkruVfVAJIirvJ+xEh4
WboGZQ1b3FzmZmrLb0TMdVe6wjIZxDnRHu5nohvp4LLhMM5W37ARyqdZTyFssLl5
qAyj8ZJpwMpjls2Ghb7mfLOlcr95EoIi9IHRXOkUsjIJt42izO7N4onYiN6U8KoI
X9a1aYFtv1NIVMIRUU3tRMWgSAcDpz7NxFP5svJXQ0ubxpIAPlrJ8yIkmbX1xk5O
UsFZXggOrpwwv2Gs+yU3Joy2FxWCgatoLR1n04LAcCKrButWwdeghp/cjfakbubd
tA19tpRVFcjOVtST+rNRwbXuS8mUkeDO+PwF2AaUw3df0xDhchHFNwfGBL7kSeRv
Ujsqa2+jWSbHAmBJE0M6/j/Mfvha+xQ0Kyvwg7nSqlkgRvF9bHM1Dc49eXeWXey+
jRzTdO0FlommZFFVdk9+Kv7p0TzMQ83z1B2NkObP/BEDdc+gROsQFdcaDV3lDreF
mIbLBoHaPx/qA2oesPgqoPv595KH8GOxuHwONVfiY2jxZsw4KHSNz5HARuzIJxnS
0/u3Y0NBu5oD4LkhS0P38ttugvdoP+12qNSkXKZoeBdTyKWSORay6LfA4kz9D4IK
2b5pZyWyxt/XxHnFGvRCGd+IWFfI74GwtoOFZjPxwHOMZb9RjYJbVynu9V4aVRUF
AlNwqJEDifV9XLFVX/9IwWr4jYJ6+ULkRUzhMFPDzYjCejT7ti5yvYX2EoY7fVUS
iXxv3Qx5lHTG6ylMUvGtWW2RgpUt08a3UH6kCRuse5QVPUBfgU0BYVQDfoPKyZbw
9YVrvPDybhO9HB2/W03FVBcHXJ6R+chmCLelMqRjugrWdiDjMRjCxHKXG14N44sl
5Deoe9fPNeRklxBKR4pbrLxsaczp43ejuuuGjYOfUrbTSIldNGMA2n8RJe3uRnJ2
hCQcAllu4gXLNULkS9QqbF39mEdDyXQsttU0MSrk+cplCfvtmrpjwYcTp+k/Q3UP
s4xGEWF3hISfMiCiCBi9hZFHF0vEv+PK7wk+GvKzdAw3zVlqETtO25HBAjV4eXLz
lmVz3CcXeb5I6yqEiW2SGEo5K96ZBkRrRpnpsh61EokMZwlEZ88EODYr4y6eeqEj
XBEJiurfof4t31rKEFZA6jvH+vKXDQtt0ix74q85fnFUxTE9PLQMOWNN9xlMc0FB
ILh6JC0EOgt/9mVvS1A9CDpFP+oz8ZdmdkTkecUWBlsXdAGpGPy1eo3g6ScFQnQ9
Y7bDRyq6swY+WmYo7xbzg7FGh02vHSE/mvXItvyvaV5br0WIVRvV4WVacz2zWJTT
Qxt0DiDY05psTs/my6Hv4L3oRInM1M/bx1z1cqp0na0di1dQ0BrtRYe3FfQqOmIX
7//Jgd8b+jdA48sSTN1cxEBILadcr7eSjdUA5R78g7pbomNjNnm7HOzrxcvi/EoI
vsALcAC4F4WwMk6Ae7dRAzOUZY1YMCN3t/dBtfNAuyvnIaV13XGPxMBzjBqKBvUT
5ATX55mxD8YGRy/UUyG9FstWo21/Nfr3vxcmX5AT4jaEQCnXx/qJy8LINbRSwEtN
L2fd+3hK3DgHHznMBo/YBdJb3S5/aOSiaQGlwwuB2Rkg64ptdZRwgJooIr4OCdP8
xwZ05/YoO45DiVu9lKRhka5+66iNI0o/wvNYUUtm7FazYEjYalAn5WgHhhyXjbS3
in5C3OmAv7vxV+5B4R8Zoy6unv8uRjFPkrMyU60W+687xdHimDuoYhzlMxckUVUS
/p7hkgjpEIb3sYCt9A3ZsePru7E29TLqCjvstrouCQ4iocM5sRzPmh7Aatewqhuq
afdecNU7AE/Dc1OUdbhOtSKsUiFZXeFQnZ4pXMRcXUmWX1VGQN5+va8w7msiA2zV
nVT6IWcX66oCsXa28x67WEu/OWACdjFbGIB5Dpcv8DBjMcCnaAjzPQiuDxlyoOPT
zxoZdq1EhAJ24uP5aE56H6SMk3ghyYRtUoqCrBK9xVO3K8/NKybnkn04B2v/vVFO
7ROX/9Xsrt8hWOdKmwvd7amT33xquWnaJSi0nUPcNuWkPYgzZwfwBEqHq8qFIqUa
gvf45fsm84FO3BHcCmQgEzv+ZR9D6XVwajsglaxGsszZuXHo1tkKoyCus2U/qHGi
9Vf1iW1hobXPIY2vIkBrnjHtyafUxdwy9756gdR6LC0ouTHLNEpffWHJXxDQBELQ
HtmOtyASYpToV14ALiWtcv/krSdIxpB64QTHENbv4GV/H2++5J6YIY7U3FYRsM41
BsDfsDrvVGmTSZ4CUdK2Svk/STCc/zdmmAbGaY7zZv0tx6czn4kM1CtX38V0YF/S
fwO1r9b3rd1X7skIBroxUr3XzoDAZW9GKFakHqCAyaJfWrLVxo8ehIkofPwoN0vc
QQBJFyrr9/NrblvgoYcXmLsDS3scz69c713lxmY+O9+voZbL96SP+o0uxaVrKDjE
XucLBSOpES353SxRvce0qQQ69hhr97ijMr+sjDEfEsSIvnFQh+P4UPX7pCngHhFY
QjbJmLKxuJR3RraP2zCryDn2a1FCeAbhaZx2MlJZckhCTnDEetwW6yDiX1G19KM+
apr2zncbxYfYnazfW9wsc4alk8CbAVb8u5A6oB+EPDHRAKxI5B3RtOJUZj23AR30
4wjoJJJUL+JX9COIn/TJ5ek9BKTjXRQbxaNZPDBRoBI2W5hOhCZ027c5OhPz5NhX
IWx39jiFCkLiGeZSaEqx0+xcQIRzlcBK/rVCXYIV3RqlxY5h4JNMJYReYOt9mZYK
TbKj6BamcAmNuVdVTEdTDKgwaNuSoO94dV4Uvgv1wQ/RQYyB5pAgiqIPCJJfGoos
5Jmr/Mva32gVFJTNKRQElNjYdqchdpOpdqqBsgZKUFO6YI2Y8A84dC1kCpZnMhv4
3QFxSY7KC7JVv9TC0GJsGqNZutSgc593FfUONHPcuCdVeuEOWF0sTiA0Wx2qgrY6
2f3hqISeo48OS9qFPfXmzuZaULrmPxa9N18j3ypDOns/C5llQUY6VRFlOdLU2LtF
30FlglWy7elPjYP2ofALzIv9p3z+Oj4jAv0nrsEyqnB8atUWvMd+n3aruQoPPkXX
TQATqTgyrYp1fE6fnTKYIdkIg8F4yEp+wbPbMJUjd/TnBEib0eHwsCKA8sBfu3PW
aievQehhVD7mnyZ24bDEz1v6dbzdmZTtOt1pFBjTcvXPER1gDKs+s4+FTJpXHU5x
+GA+lS33FzTauaNpC8eFCoSV5Z5DGrMhKjclgn3a5gdtIlVIqnMoziHkPW3PqtN2
jXdu8fxFN3bQHjTXw8K6zvGgA9x35FMjmNfLIejJiVkFzGu87I1OBH/HQQ+Vr/C2
qFQVjfq89CTIY49oO9p6wb3mHo/IIZ7nBWVTFkSa2LJdJGss54I8k9p8J3lclLSR
mr8AcZ7kx5vt7k6t3Mw9z6rIKGmzy4e/+TkA2fbKY5HLs1zFhh/zlbJ3UywRhnAe
kQi9A+bXQY540E3hHnt8VU9vNw5hxD+JKGa7x4oxNVzJ6e/7wwY1tMUol5lCz/2g
0f/Othnfu7LkUsnRTi+Q0Z4dch2uzzuQWEzEReAjwPHiJt8ohYqsjH9O6cg5/DZZ
Ru5SxmcVRqc1IyQzFsOwYmBkuxN9uDa5pah1A2XZJshDEqH9IUbIf18YPHuAdBux
JWgFoX2rbAoBJU1mF+jTUIH+Vq8NSlYmR+d/k0cs9GUwNBkRXXi54R2uXJO4iKw/
gjU64aaKS6WAVCevSKVxW/ioF9ZfEAGkfiqOUN4oSPXXfd8pPGuxgbl6N5lnSPDx
4n5pubVhs1zgNrMVVP9Tae4wfSVRmc/Kzm+VpyStvD3mndnBn0dUqmD06kCnF3Ql
6sO1iv9XIZC1V6h1WVs6mujxegDLIkk79bTeSEiEwqt8qRA84J+zXYIg3ldte3+W
DMitjeoJo+8nttAIZyliskA9zKOK8PlluwNXD59X8pFvYC+/xI9u0QN3u0qdmRaL
D58uRDGlBhjKi+ygJSnoNFanjeHeEzEvCXaTCpXWWDMbs+FDwV3DFigycOv7KbhA
H1YzmtfSP2aTfPWhtHPBm23nDpbjyJm4U8qfWyKA1tK56uN1FBmtXBWyrvY33g62
30n6lYECZOe8aVsYmCQ5lf/DDsk/CSY9p4vM+2QxTjfpAtaov1JiV7jabOGf/YZ2
M170jEag3IeT3B6nKMhMS7tTIjk+grYbTdFc0knnuN2FV3lXActywm/7Pm5u09PR
yu6qh4jLuZsUX3mceSGq4E8fXMhlpphCBc7epwQkioAevksmj7YBdY32l3sibEay
u+KF5LUY18zIgrlfTcGIgznreKihZuoAu805cocSycDCROnlfZxZlhRwe4/z7G+q
sgPoQf6kScVTIxkz015rPgpAB1QFwm3imfvtVROzLAHmvWVWiu7TB79CTVBwMU7T
V3nM11EWkl4nMwC7V0OZkrhwIufOUf3R+QqtLxa82z0LqWkERbpZ5UrwJ7IzlfUx
YypC1xwDuQ3z8dAcXRl7jlq4RJu8rNOJ/XlFyFeGYqmGP8nKkfYEWEKrBtK8wtcG
wdDJPlJcbdM/sY6sBQIxHJS50w7yMiOYdm2IyyScwFCQRY9eGzOM3oa0N286V451
ECf1Tr3W1xmI7c5g4zXPGYyP4AVP24uLZ3tkKwY/ZrPuEvekTphuo4z1LN/dqoUk
foHtOqVz6eJLzt/q2HKrYyWgMRX+CcGp6KIFTAotUFa1V+MQ2PIN8tTJFWwblp5j
A+R5ON5BdiXdtJhlK5d3u4e0hFbrI+phpCs+Nj+RJSF/MYDcej6AFCXJ7rbewk3l
w8ercdgg+5mnPReTuowNJdUjGjZacjy6wqPUILdhrs2dKqM77l48gG3MQBHlsKZ+
7FA+faQ75bh2iMLJJNfsKMaM5KD5v4Osb2Im7NWrInLw0/loi90MvMOFdsx/aBeo
sLnkHMcpWadNiqGWt6Xp3czvEZZkYQdLNQw1rW3/34ahTWu38dSot+iPXvRKbYaN
YChatrc5WoSXeW862ezmIEMUaHAUd0GHipud6WEs/Eu6KBOLus/QNJscY5w8Bylo
NZPAZpBkFD+GQEUtQZzUJt2mHagQ/IJdt0XptfnQC3BSUCRcmGUYS7DpxMzDUJ+7
BZthVUMIlGnCt9sYv+owPWFsiEbs+9KUmRo0YJvMqyV0XJnFnu/Q0TQHxLJTl01x
0YBsRq1VULCl1Xt7EJdI3Ku/bXMTbxlDtFsTsZ9Yjppy5xdGm+BgtpG7nurSIB56
05B6OB1IyVxm5U+kZlDUoHOV6QBmCK+q/3k4hVLzmjHMumHmNR6c3B/ooMN95FsZ
eEXSpwho3TRuEvCRYBJxdKmqFQ65zVe1X6ZTKn14yBedcrgWSPGJLVGGFvVEQUXX
/d8Zf1czEqBzo/dNV16PtIRfLMKMLN4b2MGIqAwmo9YTlZaa88AWWx1v5JASU82A
h223fPK+QSUkyt9VRPeWNcoN+DW/Ex/3+0eRB3rv8rR+ig+4aofcxl55Zz8T7ewu
QpEGjmLN92U74rLP3b7k4pXF3T3O16P4HIQdGcYENsd18qVLbvd4zUETvMD+9O1W
fXTE2JdEiSj0MWHfAo2STYw4cSR1ZG+BM3wzKaWU+04x4M3/TiQ2RdM64dNdNMSY
cufIDZooIQ88LI8vhMPhPSvxroZtEZkeBQezsZzPYRGgk0MG0CwDvHEyHvVa/maZ
lel4K+KReGvE+hpj4W98rE7FISTh4AgsNwEpxj97W5TBOqRiIOaqZgIC0EoUbem/
YXltEjM2R36PZmqcr/mrq+rNjf2Ufp5Qb3YIsiJ+AgBRDN4kySjgI5oGmCh2IM3g
5qeYPKBdBRVa8FlrpxoaP6vSSfuo0jxNHgoljOUCDttE1py1eLW7FFCDJ8BPI9mG
pWgnq/bSXizNpYTya3sgb520cpK5eQn/VMrlJ8pnkPn3Vm48lNHwvNujujDD6ZWR
iZ1QtqctolFhNu7U8PoFmnM0VV3zU1KSqhnOI678RwUekdQOV9SjpcyYVRVq9ztU
qQW0hVhwAVoNm+aBpeEbAuWIJRxRthpOkJapBANVEyit8jwsatu2RrlaYt5/7Wq8
IniejqEL6ceWpco1MBIUgwThfcdKLGLpvYUhqpkBlAKt1eNQIHRunVyodrpDQdNv
lPGtAaHM5yT3RpICpaouWLDEaLCzG7z63J9w0mBEYHKvwyv1SSA7UOV5SSwPLcse
FuWbJLCKI0x0C30mEEcQygEvUgv2lVDZ+9HYDkBrA+45qLFCODkOM8AYHkAHxy/c
fVAJFBwvYN5BzWPVhWe6muRsD7RY5rqSmsAdVP7woIHUmuqVX98/xB7hxAAuB8sT
WPVWsbI9lZ0vGaNq062DHcwRRjIq/hztFmBvg30RQHlVzRZO9w9MSkVQFzyNlNJe
/qw1WN9zHAp6fMzMtKFluamrMzlpc57TqS9HIx33Wkws/TWrmVGkmQFFYpIs1BcZ
QVPm+qmEnr3qclvzkQh46vRqkBem6E573XqCLMErTFKSNyWOdrArRjlFTbTaXRFP
2pu+roqpTPnC+rm5lpb3DpDl4f/liHCGmWyKbZ6uMEX+eOek9dZOMiS5xZnbQ1Lq
5WsipCNBthakIUvorJkzoCsIMR+E8pjxM/a2/qs19PZ0Xg23ystbgPrMiRBpA21J
5xfihejpJr+KC96e935ATzoF27rH4aurDC8cUviaKwwWH2WeLGHMcFvDe3DHmTjg
eBaWyEX/TSsXKu0BJljmNxEBXDjOnPZGH5bCY+4V8KQpwJdjrz0WhQ+YaV67iKKE
8y1K6xyRDOGg/oEN0wvr6zD3j/84rbswN1ZT7GbnJ5UwJy6MvOS04BK3X36qnA9/
+Kdq1RJNjrYFZ6SFTMXg1cDTjTwVMbk1Uk3TLEKJv+MQ7FJLNo18AxNkqhNWFpId
6ieUygAJruQRhlFYqdUurZNPBSB2pm9h/lCljYTN/YFNbwUUG5G+wpzXHL3f0gtr
dhsJlQAQXgrq64eUlFIFj1mMbk9axg9qTKT28HhGukJJ3NNIGj8SfLpRSi/9sU5+
A/w5tXU1aB9uintbQmdG1FlraPoSuRhyRoV9lulQiwlrKorKRJtDTRVqu/elLGzY
F8HXVJ22s2i3KYDr6yE2VSSmdOThzir0PK0FSw4E9t6Mlcep3AMLCBE04t5eqTMy
F4a8LU/FfrhQFE0xAnh5d6CGst/lH7kgy5XDhZ3z2nRVQd8KJCkA6KdawzN7dCfH
7nmPuYim/vTMlzhdhW8oQUDE+VK4JwhNew6iMXSz+bGylzUOwvKwn673cvzVQDTq
GIGGjsjyeqXtmzCjkm+iOttQdoFtfOJA2hftHzoh2t4SVXawD6tqdLaQ4Y/+dJEO
248a3pBng767PKK8ezouVPb7jy/7+iKRHbijeKc5yQH7WzXeeoHSUcodsSHqJ5Hg
N6dD1itnQD1S4e9oIK7OJ42bqNc3ekbl+2eZ0wHRpHaagFUgSWXnL4zVGFmPjyA/
cDcJcyPn34jfRh+qdeZEAexls2rGx0obvBJPA+VkZGt4jwa5IjGrPj12Ee7EjtV3
yrQp30GmLGy+7u2o6dz+KWS4yB93YuGMHFpJsCX7L3uffJIQ+P8/nwG0Lsh6ul2Z
2Z+zfRGTaCg7td8PdPo5p+htk5qL7/VPP2Sm2V4jHQtw/mSXijn7Y36f2H+9VLkf
6MlUCsIyJodcFz5wKrLpDn7YJ0QZn3YT8PgPNzpSu8CocLNdkMMS+ooUY73SUKq2
JTzugdDIOGwtHuWss6cYSDVTFW5qUR1lPPc3D0jr//tma9QCsqdZVL3t03AMporo
p0MfeqzottPOAGsuM9HzLok+2Ts7OVkaBNzGBUEDFt/iScNQTfXxdGEBz3mSkJ6d
/xi63IDMdywoe+PrndNvcphNTPIz8Lb2DDNN802RFopPJQe4XwbDfrLSChvRaJSJ
fWnCTX9bAxtoPY2Po0O6OdlLofNT9ooi3SBLHMyQ3mkrDXUSd9lK9UQOC+0Qh90W
0yjgkyJJ5CO7oOSsEUg8cnxPgpHZMu67a0zwLZzUUmKZqLmVOLEH9CFv8k5RG5nj
XJLQtg5td3uq6FCUBcziWZ4NDPPIwYIEPqZMMcPJ9iwoqWt51CKGBtmAu4S5HXKb
KLT3LTfeU/Bk5R433Jej1dEE0cLY48FPE+9RI6dk1qPNnD49ec1I/osp8M11CzNM
viRDlrzKjV6kLL/ptDl9doT8qHavDMq6nx86S5nIsMW65ckPyjOXa/DH8Wpkynme
vRAu1cQrzJMmRvDDRhtpqJ0n9PZfBjFISTmSO9xOqK4keYJWLICXXGaAUuOH/TX2
nbdxLALaz3y0vSZRu12//FVr5M8laXaBBZE40oh0jncQrK2KckpJ+pt/FyVxXrxa
n72MAoeCiRaryWbHbMBKERwQTLmrvuTlIsoDFUi7C2aLdiCvyVVxqAO5i86xWUOH
SzoCUCF1fWCj3JpEHFeitw7XiVGnpIdHLphgL0KlyO79s47Xpezw7c9bdnD2tiO4
FDSX+WZjpPqIjoj3fPCrxHFnGjia1QuFJ1pFv2MX3jzulMc6SDcLqrjpTcAB9ew4
Uz3lwkY4PXY2xsg/3xFbSRCpM3l+NWzQ0ZMKyiNfwIseaeDaIHbE2jBkM5MtlYYt
Pos9coQO6pIz35gKqah28m1SemVq4hrYzjX1voucu8ZVZjJhOOr3TL/vviHAM83T
66run24TIVWH8lWMwK0ANoUclTCsP0e+XRACH0zIT7k9Hz8Nm2if+g0e2y9fldvJ
VxVOX6A96mgdxOe7FRbZQvD+tVQA+aoWQJUW4ID2M1Wh7VbKA8hmyF27ztcxNTre
VhoSYgexpD+h4ZPPZFUMNLtB6GxpXJLs0MrAGIAWw1dlidHe3IWGXPkY5De0zREd
51jey7yQLuKrcrVrG5E4QX9QW3XDW8rxKLArijgMEe2t67fks5iky7oVYBNTVHmN
UnI6wfKyeQQWikZ2RmZAa3ZpSFQKjeI82+4cBND0upoK5fxaFmm2C6X943ASE08Q
nE7nzlX2EPAML+PefOX9axkPsbNZnyEQRJyTjksW3Vd5R6nkgFDNMLHzzE4EB0/c
AYLo2gfyRTjC/keBZc9ixUOIimsuj7YMqrP42tYvZEK0IQrwCdrWtZ8bmlGlkqls
OdnCrNDE4AC6QujS7dVEyfHR232hc/kMPhnFaEKolFkTtKIGwEc0UZCur4XR2vFP
fRdkec1QkyRXKKBv8Xns6aqs2RgXWhLFkwzKWYT8CivZsGHgzUVR2mfKo3w7XtW7
uyxpIjGWbQ6aWLcLjlf3UpNCfuBTEv+M2+mOnK+F14fRD1X0dGPCynhScCR4us71
6czLa5BMxxkHP7h0hNvSEEHicRKZXrqAhSHfyFJX7AChryVxCPwWZ7MEx4z6l9hE
46wbNKDOcQibOBaoIk0gxJ3UMnnlO5km160D8o+b6PsUNI2TM3CaUHImfdQj3ii8
pm0gpzja40XZ92YZiEuJVgyWGBDyeLYm6+7jSRLoISc8WHChR/Xi6eief98uZ4HP
UqVpGjEa64oYUUZqn+tK2djPQsy3ds+VIyf/wxk/D/f7QZ57i+cMafe9WYfitWCs
bLYfRARzJ1bfiP+wORgxdv6gAPfdvj3u9UVoQzn1mulb2MsSVXb6kPniSxTSVtFE
L63JDZXzlxCYfqFAYX47fa3MKM89bFS74eSz2vLQ8PlfMX3Kp+lbTRObkAUHTHQs
50e8VRqy+K51kf1t1SxuymupuLxvIu32/cRpeF1A7ZnSRjaDAJmQLEcSy3134rVL
sUN3NRKoTtanjQvcTtuiN4ml09wnpSGgL0gs6YSkb8dIrlTtawrSBxpvILLGBq2s
mNBesSeo8EurVBYLHJQgFf7RTjpIrrOVcXYYIsDGny9GpaKanN2nhL+DtQR7YV//
RSHoxYqQD38VHDg0liWDZwLfpi16N5a1KOfAypRtKTJLlNm+14fqUS1O/WYP4XRn
Lc1J3ZEO+7osb0cpqgMl//QWhOEDU43QSXo0Oo8YCaaFvfsWdhkbnQKw+rHjLY2A
SMc446UOmxdZ0+oZXNvJPr/k+G19KmxirZTVa03OBuJQq8x0nSKCL4BrOObaCxwy
2D7ItIq8CcbwpktHgfHzxMUK+22fpwBNCkU1M/Pv+8+MWVuHwLQvqg3VXAQCz7AR
9vRxKyRrJQZ2eZ1SPkB6xRlTqdGVnMsqTYHWlfg0vxlV1c4kbYBmvodSBslWXNy3
hoBerzWPFdSQTEiLkbFrBtncaZ+WhTmDTj1vkBDW5KKc8XdR73/5+yCNfqZPkhmZ
5YJB967lKPygZeNBGHOMHMb1MX9iMBkMzLY+4fDlZ3anXoEzAcXZovGqPfItWgvS
L3Pk2wjblQ4e4ZMgAetSjNALdM5ZdWMZtslJUKkid8McFCIzUUt/kumgnkhMUwwm
JwvInq/eJ1vE438LDBYurkN/KnmdP4s8ubFan8obteshreFnXAILAlyqQLsO4Mam
ya9wMYM7eBm9RbwqAO68FotOPdx7FJ7Ksh2oJSGnjbt2cKA6Lx2pQPPAn0WRswsE
SLQuzI+uGnuKQqpDw1QCMP9/7LhtXGkFj8R9JQEZ7SIDvP1R2QuRaI5HD12svfGU
HXvqRoSnCfhdBtN5iR4AtEUrrcVxVmOJj5mU19zDfI7ZUa3OI5RIm92F+fsWXdeX
wcIukowcXmrN3pn79ddfmrRHf/2O6CnP3Oal1kS0CRHOLPQihTkzZ2XjWNPKMhB6
CDKmwmCr0/OcVzGlihrq5yh/5Q7ZpaZKEgAgKwQyr9/rwDzn29HB7MqN0B7l/MFh
71HjQK/Ja3igRUw8BNeeCE5uJn9rlRx1h5xq4S/e2rxvQ6XBLqs+ZiKwpQRC05oF
6TuXRscFlEVhSupOm9vmdB072HPYToFjWrDM92uSHcAkzIr+OZihIQTB+vaaX90n
TQbnn4X+DfUATOoJPkMMZvxRqbrJr52cNMayGbQTjNdfX3NuK7ydNO9v9HDMUim6
YWr7INP3HKHZZjhJRPQMxm7ppN+XiFS/cpue6X8SorwCgR8j9vFyi20BDhsUI8qF
YDWZTgC3F+vZ0FRpgv5U5flGP8u7/hrfD6s9hvyDS9LzttyQpYh9SmZVlmRbV+YK
hynSoA6Pa8jdaxpOyiVzIXS83H7Grdzk+suY9CA1EfZUSIr3yF0h1hRrDRYjRElE
7fw8YCQgm5UWpwNsdOXjyIDs8NjxaxFLVMW5txwpFfG9HQUWxmJCko2VrjEU3t1f
1/hEsAoj6h03/am6M74Twy0lw9RXHtYJRFltrryVTi5PpoeoNN5hskoa0CvRkfMe
OZSUbbDsjFi1O/xZ31hOeR17tzdUCWo3iYU39xm3UeKu1W+4YaHy9YFiwRcjAj9N
5MIpXGZyF7cvtohJcm1QlW0dIzsy5Yg3H+KqlcNjN7YpwibGIWOgsfB9pVwwD6pg
zo0EtS0oPPFL73ShDmvmJFzUuRimap5MjAGmygqwN5R3RZVRH4srV7bspRn7y0yK
SxRZ9dZiB06D6k8gsquXBdnJsTMFo6NRX6Oo/yIG0O9xf+Pt2F4O9ThRXD49nQhR
RVThaWEpe3qd46gXH64aOIw/jm8fDA/JXN3c9cn3x6JIBdInzIidvO0vvu3kY4zk
FLgRRJe9IfPGaWx1goERMvLSHa6B8X6xpuJNU29jJimrJ361uaSAY2xF+nTgsc0Q
FsLUZGIOWRBgHYTQZh0rgjv6M1h6nTCSfBcQ5ey+b24ysuDf2m3V/qTZzBUPZ0QY
GH1TgmwuQPpLnY/RFae4tJQOoUGd9sbIFtrv3mpCDP0EzquuSdWfleLvkw5M4lO5
OwrxQ1yaMfX3AFLkw7mi9V2Xh35Kytmi+XqpGgI6qwuaDgggYys9jMnOAEc43svd
GFrzDeKKikf9bth0NHxjUbEYVlFSbOUjQ2vDjFPBP2V1RZtIlK6HYut5912yuVke
6fZ/Xqem/28TQC/zUCFX7jypMHjMPW+F8wcFih25hrcqKAwpTvW5ntta+7LSLZuT
bVut17hWvcv5c0ljQPlIN5ToiuddZOuwX+XvPdYOT6bUWnWAjuV5c9qiMHaUOf6/
1kzKaNjICi2fnv9g17F8BLKeQ8okgKfZLV/CWoFcL8F0RBgtWMtO7CugnfBO/QeL
bDRIIQ7VbKCVjBUhrYPDZ5nolVb9TOVqJZEG2+wEojejxyoHsiC2CUzqzcyvTM/B
XYK+jKRXAM/tQg7EdgtccVxWv+MNsyBRVK8vwzqoDmPHy2EnxyBLj42mNOU6H6jt
9697ziW+vOnB/iYsTFqb9k+U7XZG9UzOMwxJT/josHc+akKW6QBptT4inQsUDbS2
rbngZ04jS0AesDpXGwhPLaX29s0jQDAFPsINdekgLGX6JDzJhfOjSJ5gjrqgr3QT
6uAZTkqACavwmCG5esJpnpV0e2TtV2k7Jn9d2weeGzFNV6Ch2wDQx0PHFBK364vh
JWJoWxLf7qy67hoynHHiF1WFTUsz1ncfjebCGNNheMEWotKCJktDHW41G3Rcln6v
f02o24iMaSnjWrHQMf76/kfmzIHfIcqFCyqN1jA1wYuTvGxoemWGTjQM8wSBguzr
n6xImmExBzhjddvI6znWyI7JkmdEKOYAqTuslc9Jd4cQ147xRdTmvtryDrpOk34K
kt3ELXvvKgEIrF22XWC+fMqA6dmkfI0zP/Upv9nhMT+LFKw3PssetwYaEajUOrWs
5qPMWbjCFNWmNVvz8Fkqgkb4a7EJKvQT+EtqFkQZKvwiJHW/+UU1zygaHTlHO4Jy
ChIISjJqWJvXcE/uXOu14I+nSnGPpZkg5LJ+rGou0POwRm/n8gDFbGudMkCA34R6
GvSPLyg+NPbCBmzJmPmuG5yio9S/LZQxYClvXgh5mQs5SQyLP5M8/sZJmNykEYJs
QNQqAti1uy7jfsL2spExGKa+J4Vmml+OamO6sElwzV0PyxP9+kNyzTBMcl4l8ogV
uHZfiM4eCsqDN7/ujFbGhlsr9BDsHAw0TnRUFuebLEkBqKyHBJrUY7yYZ+v2tvo9
lnD7oxQ0OHbStn8dbGzwG8oXALNt6F4dXb2vO8IxrapIQtxtcNbJ3tN2KnIADLY0
DbratEc2eNATPxfgnFSZ1efIEbvCqNoPSOLjheQnIjL2nPjCjvmKf4rACJuulOTQ
WubLg5nQbkgf12pm/G/mR0RWAjd/QWfpX225dg2/y4gXoAz+841IKiPty8cUsWLw
++6ZBp2Udr9qge9ol/ezcqAX6Sn5Y5LzEJz0Dm7z1TL/B+EQeL5Mc4RuWD4m1aAl
9LGRJGkccRxBYZWdqBw0WRTL5r4FnYymS7aqo7lN02TXxEjjyKRDEL7qJYa9Hgy1
Kp4bNMzepx6qnrFe1v4txCylg3rm5kGox2bk48yyggzIEJHHjtiFxwMeksjI3AfA
MH25uWEXd6pGoBGr30BjNe7WNINTfy3adF0y5pHR97k40t1g/1Zj0I7Ve4/HUaGs
Hi9ioDsfeRytQ8Wuad2WWGT/4xo+Pu2bnAqpJCYGmQQeDChnFcXJjZm5rOdOjq8e
t3UaZuqMunjwUGWockCOHfZKVp6GhEadRefA3QlPE0dn0jim2CUuAaHowiUV21o1
QYpKZ/ywNtwhoFRmt9hRd5efWG8WObfd6BnylO1/j5ugrUYlPiz6aRCRyTO3RcjT
yHCEwCpTZp7tDQbMOLpNFDIXuQ2ZDizfux7hmcuLFYmMGRjlucW0vR7fmsh4XyVI
yufhcYUDGHZJvSg7LwOPpipArQ7vvkF6lFkClzBDwRUceEdkeZwj8Fhax8fBwycR
9UupKB8JOsyhf86g8gu3NqAktwtBOAAxew6aB+yhEXST1r5UjbjGOwC0gGIBezwP
zJDT/Z0fUsSp5OezX4dF58dmBj5zxsDFDg5CoFkhQB/NkYiFRY+mk5HAMQ5Z8NuQ
hQgMfgeM3SR3txig1nYqtefOYnzABVu53AkybNpCYe/UQkT4OV4nYUqayH1HmoiY
a7iw2SWsdJxHarms7uHgBE8WV1K0HvZuuBybztPFWj0ohbfiwxJ6KOL+zYXYrXqZ
09dWMqjWF4TZ7CgHAYKByRTRaDSAE+bv4qUnun7nYxCH+PvcDB0ThRdbXDjkBjUQ
Wz3ZrbRop1ToFurV/SnGfjX4aWJfGazqU18zQai/8kVCsH9ICrYq1y2Rrja5bZHK
gpcM/TeGNTekxl+CRAQ3ZRy69HF7hPDJrPhl3ZSQafLYAIKquX8C0/pE5+sHHnco
ZZ8d/ggPINWjj2PHPMiiB0Qq/sSk4amtAvH2SCIB1n9ZcxNYsZcoU90dKVChMdPm
Lm+es5uiINQ1jCJQPTa00jRD+nX5oQw6prvucuv2wwWgovukJVRPdgNDgLCVhWT7
+izHDcWSZxXhu2hVV/LKrqiaDFsVShLFwsC/igR/VwaRcgg27/2+5FKG8R8h/6cD
jje0qFYvFKBdqQAyb8v8Gq8LvXndnvOizrIbtWssXHA1FdJO8eAqMBku1Xja2UXh
Z41g/rAIxzvz1dJWopo8iS0k4nXHQb+quF/zRenxKw9q4OZZOKZxP736Tkl7TGrX
QqiHa5Jh2f2h2GPDWQDCxt9DtZNTI6BVIGJAOYxyP+AHvS+/RmtXb+nstLvv/SPQ
YdXnKHKdNzOHPV8t01n6myGy6YO8JnC3bwekTpMplLPR7jWtWDu9cwRtsUAPKn+I
cSMbdEdgKRCxADaxYcrO/Q4QthFEDA4DX8SIukOLoh0ORjAkgOBA4ngE2gSeUvQl
WWajMEJ5ZR56C61NfulVwVdHxpJ8wV7gSlC+H0Xr/f+AaKiYTSXSfyrPrGtM/Ce8
6Dpqw0ryI5rnRctt3v5rhlugvOoeVgtyG3DU8sAPAlilUe7/bOtE+U6SwC3+bhz2
Ji5O/Z9rXsuJho086xsofqlgllixMpJ/6gjM98FOz401YOmH+YFE3OJMwAKosSgG
rcRQ8sQDa5ofx1JfEgJwbcFS+ovMLoHhQ7iMfEq7yQxLLsA+5AsjUkfXAosvITSD
Sf7T3JV+wTRBB15dCohycMKIyn5LysYc9IUVoSVQFjTZxxdLs45FQ/j/TPasfdL5
5PQlK9/Rvt7aS7ZHQdfdfpuBnXQ4U6/NM8wyFYsTuUZ4/rad1IRw1JlRrhtNxXPF
o5030dor1t0c9Oedgco3FZrR3krZpWasI+kFklUuZox72gXH4/FznSm2n6l4QiUw
on8HMkBD9FxNvoqQGaGmMSfijVOlTQUaCEonq5I5oSZEtZQ0H9AS95culk8FZYCB
yotxi7bDANzSBl641ZBa5oTOvZ9u9Tcv4N7whTHkGn1AETH6JVkJSpCoehXfxoHj
zYc6gr6EEYsImw65cD29yl26lIVbCHAlVCFkgf4ooW6X1hedM0Y8LNoIOfUNpZW8
PXLLEx2rJwCtfuDWwPTrhOEJBIeHnu8UQ9xa9voLcJQHFLoYMnwbn2HwUzKzynkE
dA/3B61j/noB43JOLskgvewasoFp8J1cAvK1c8f8HFYftSpo5aGnZUxPdzat7v9S
l95Tb2TFdZ2oErXe+RmT7rm0atSDCjUPSqt7JsWeC2MyQa+P6Wn1+Z0oBbMzk1M6
IKxj60vfdq0yweWTi5DUB9xHp8J4cUcP8NjotUPZERqTyHGwoQwDsveF0LcFUh2v
y9rdacDqpNSlS9RF+qTUNI4lvcU0kOen+AJZz/2s0Mxm+JC/kUP4kN+7a1yo1R0T
KKY8J0p3qnhgLIzHpKekPBI+UROzlFAHavWPQsqvL8CCC2MIYjfnJlIWVvf/l88M
Ox4xsMYPJvz3o38ZIeROP+4iwxS13CinZ0VexKeWkeB186zL3Hqd1Gs6E/0MJfdr
2E6JejuFWQNWa560ndKAtW7j4IXPAWUZMkAHmLQHSWgugr4J186za4N+pUyDOBXS
lMK31C8CsIq2YE5pYXEPtQg8bjG1Jv1Ga9G6zpC/SH+ik6NEl58jb9Q+FrjJ5mna
JZ5PGrK99rgmIk1GTjI2moDrxy83cwVtpTgPC8I1889tm/0j++KSyctfs1XHNvSg
FQvYWYEDAHq3BDkGW/FNzM9doozYEoRKlfI+WECXMeiRCvVLLakEnkE9uA5gWk9e
/1poPEtQcaS7Bj17gqvBclvGMHRwXcDLnIt2M2cscloHzjaVIyC/C48OowcmwK2C
Qn7YM/C1XNQA5ejSfLj9SXrlVZjC5AkVXB3UILVZvmOWN30PCMve+/NujvPXrg0k
3NZxDPO7T5xaqr/96Fd0GVCObZgYdAho/2LCK53a/KDOXAAz+5bxaeCQx9vjPqHg
bxrYDFhzGBqeblSvbdORS7OtPEacwmeDLDhoMMsdJOfW110xgrP+Xj7VTMHo2Xxz
f5+P0BAmNfAeL7SauuIRVB+/iiqCR24sZEODg6aoneHgpP4YXG697/G5pCR3VPYA
qQKn5OPaIftzwtOvGaQZf/nmTf3b1fOYaewT7JzaHl6dbV2SVTDA9URL5RB+4+wC
F5P1doHEAdMTahgecbFgy9+oo3lWXTi9eb3mePEwuur/UQMt1QPAamYGk0qKTJud
Tr0GAoywxtX1Hk7S4JYEVwythVXwx+1TqOnO3k3rLeiSC2l8KegrKLiqDERwmrW8
RXCEo5YtN9pEkqYrO4iP/lavibgX2I+SGGehNcapwgBLr8mKxg02HyUIaFvxKDpu
FK61J8jbpAw/fR/3Nr/XGKje+JwD5KF+vabAdiazALzqi7xwvLa8f5THuzRz2a1H
Pfws1oN94NfIjch1VfiV3NQVEwh6MIScIZ0fHLBzU1cqY7snYHCrNAqaDbJneFKC
s8uEfLhEVFxu9cUSgHkXFb6Qsmrf8YE6DyCDW0jmmwOAl7OOASaGGxtn6VNtkw4A
hZMgsYC+x4W+7rHKm0aUrCHAuQFdDP5DI7h6Oy3OIwOMUt/R2xnOH1iEUp8G80L/
K/vw51i07N144KHthL69nBVcetsBr2KwwEbk6JexbPR0Il5/NIlqEsMst67tDOkp
4Cz2hatufdqEsaSW2517mpBff37AbZr4GqashUgsg5PKN8TPZt7H4r7kXPVhUufh
r0NjuC9aIaWwgIEnQLCPnrydbsUcZqLXze4j4tBn0Cz0I1iVQAzpadZmE278jvW3
LMXIDd7CTJEgaKpP+sWXpRG88IbO8FSqibBQwIk0ESkhjexyMJ4t2+SjWUG5aI6S
JWw7KC+V+deHy2PrGiSyNimKrCKefkni/V3l5r612r8IzfXOuxNWBp58m67NS7al
FQcqpTW/+nP1FVphTn42sxWZ5T2jZivbHIJrF4t5RpaIkz+H8YlbOmfRwCi09DeK
0SQpFfc9ruLnxqsAaVOSpme6HZ3Rhrh6EiublsclOXdEhU8dzzOeVp42GMynlcFk
U7/pqGZ1kEs1ZkvgaGzvJqAs3wT8taSfzJtYieLOKIPmnMXBy8FBnq1DF1YlWnmC
rG7irVbdguYnL7mLTnImYJuCYFwjSj4VIu63kVyQwZmyhOrwn4NauqofXZ6ll1+2
g4iZsQBKHMw9bx6OZd/kYRg0sSOtt6JSF0anF04RZbftr4B4BX29joNOgpudQus2
7GXrftoih6eOtdGwPUFd99x//97SUni0rjdX9qEzP1GjNFn9UQUKlSuQWxN1Ie3o
Y0KK+NZVGFQSIaXCxU/S3yw2xNk82XlLe3SkTj9mz897m7xwCAyl5u3mssTuS5rg
xbOmWIs+iPl2WVGXx1bpdR9ayc5msHnvRDx+RNFBqp1zCXhm52cGmj7mDlNDIf7F
gZiAt8OvgJm23K9L/XpQk/jwlfoA8zSFHBcou4aMnUZd5BfXiMvULzYb4rFJVSTP
NKZ3DikI0MuyvM3Hvq/4OduHxumo60wmz58VTabHgVssrPD0N8BdliLJR59MKQTj
ptaS9DaC62NZOZatLZIX9P+MJI118g7aU4k2j+nqhL9MMOjtVOgxaIM52BbvboEb
vSmomof+X/icC9M/XSWzJgyKuEgFp85SWLPmXBmuLkAIg7AdWoD1UCykzDGMJWzg
h0+ZsLeI5UxjmeSMVGNFEbPVKXh7u/D11/VkATS/dHPAHSHotJMKUEym5RX+VhsN
Qx7plFMREOz9iXcgVzJUkG8ZHipgb4RCnvM2c0iya/pPwx9h7BZmv9rOkJ/H+P8S
o0pdtj69NGi8XseVFoYmxw2QBaApPI8O+3RlWODRJDHLaglO3K0Mw0r41YXQb0zu
grhX+e9AoX6s7hz+wMPvyZXvxeRyMl9t3H0XspxTyQb1jzrPiGDQt9bAsb8g6mPF
8hZRfVo0IBqWo3iDzMiet0C7HPE760JQEyDyXr+LIBWCiXsvprnPzm+B1k7F6O1h
TgEvw6sJ47wsnaFinohIInh9Lifrc5XwvY72mLMwHVvGiMVO/cpZmWREYTmw/T02
KYhcATkENAZc+5UzVc8hG5z8PiR77yC2gxmFNwF1KbDrTl0rme6fkzSS0dL5wpPE
8+ofir1DzcEkslZsTFm1T8TxivQZF6aP+/w3iG0i5QkAAZvWdnLhLPb6ZsRNtZja
Gv/fiEi+PsK6KcSO0/UO1H7tHj5euFuN09GBqRW7iR/DMzFTLBxVHnoQuSUWbvrZ
0C/ZD/jxCC0F/KnwEuglG8tI3afzr51+fCB4dLngOWL737DEz1256D3MQxbzixe9
Xe25aA6ejffaeGTUxHtrqY8zK/6Nf2DGedIC4gmzYxc9Phsk24GUIX7GDA0F4l2z
7hExUDGQoM3L8eMz9jk7wh7DyZjiFiZb0TUesupXqEwrzRe3+6rnbqNWIoolDz+c
gRCt9JmafDE0j58mpWsY7ilplr6Xnk6bMlNfEzoal4u90KbY52eZAtvZ82qGWHCl
rdWX4iYVyyNpcWDHfFhPDU1Pv36ZDr++gH++MGBHTS2Ssdp0UIeR9yOGI9G5Jaa4
V2AXpaXR61jYNAVF0iWsI7zhB64amyKzXO3c+cPeixU3Ki52aetLDeur1ALPdbTX
eZwA5gKEZhjZYFxU3q1sILtHtHNu6Yqxe/ozIl3wv5wCTrlzVVKYuCVK0wMVzjyw
RwJAFKEHSTD/dlDkSn/OjUdJxnjJJ4Io2ZpO8lggd1PGFtoHaLQwDv9A/8Zzgo+O
0FlIsmycEAzVDs0HbHpDuBq2UXdhYyGYn4g6IAxc4R+YOxQib5mQyfjr/GO/6F6P
/DUtoOe9ogG1cMbhEQkd7KAfxlNjpWy2HgV9wBQ/sE2wXrxodiHIp5VDefLSJ77M
rsnBFY342B8LY+3zzaJkY6lGMG5+Gen5leTJJrs9YtaWl01etmn/Q2aeOLKQCpNM
vfDSoOY+vtI7Nu1HYV1OWBb5yEY3a0HVZ8Iz3/9Xurq7qOCJyJeewkpSQxqQsSjJ
T5VD9NVHdbnPTqMnTls9YpEnu7LyTt45/QoayYewQ4pc/KLhuyFHsQiahXLfj5AJ
bHrB8W8QhhI6Z/VVpSefy1gXXbHJh4HAEuMIwuFA73SLeqSDnblRdm9w+KGy61Ev
c/ajWk0N0NZ/dFy+/kT3FBZb/PeghrhEevB3IuTZYGKfc8Nat+AeHAntRBvyIKjA
Ueg52Pr6Nr9NWeop30zIa6DZpSmBrYVGVbdjKyJsVryKRb0PBX4eCjIJnmB2RK1C
JlK+11TsiO7ZOdyg3kWUBVe/jVwQhrznWsEiEzrO1qS1qhrgSHkQpJs9u4b7v75V
2jI/nRatpu0IZG48lzKxtcLwaYkFsnLBROlorXiQgasUJghYSgWw4BVOJ7iDkehj
stD5g92QqOFd8Mmaf8xCmcG0R4TyaHxRRbJZfpMaMxH9DVqgl5ocLztkOKG6thO0
A6F/XZPjLVBvPF50+1mbo1v7i5+/VUXn1c9vYxS8Qx5Ybu0q9tXu1lnprWaX0H+1
//4Hgt0W2FU5D0FGfvIlVqHXVqWXz/jNZ3+hF8po64crIUhFPkjcIWQBExGMXIlz
SUOjNPd/7g2UzksBWqzG6IPfXM3UUb3M6xKf09Yq6iPeZsevvfbscF6TA3wtcjTo
ng//J2KlpSKSYfE+EaY5+cioyeJnmXa8VvSvOhnWkasKiCZwWnrpR3a8FhD+iDCF
x67E3/rwitLIB9PvVB7wzvf0q2F1ZoyeDmTqRuGkvmUOT/vgx4dt1vQIgNHlvVn/
HSQ2sbkSEZnrqXJBILbtIgwlzARTiiPQUCYocZ/B7UjkM1igKbUpEhxyxmRqmdqz
CPOC/WDUZCu9ug/i4kQ0UlTAlPdUcd9MSahw+mKujK95Zn3MJEyxNR6bSELqW5tY
9bEm6WAjCUdYqnK4JHDKh7xGddzsDOip5IkNIlI0eH16CPzDaYjpQyEYBgK6zQpX
gBmAmebsLFcwf4apHbldXyg9MQIaHAHwfYMJSPbaknSBd/beByBfcGGPOZQoGgXh
2RmSjhUJf9soZi1cRPlwUjxP+XEccMbWnj2LavQoEO6LO3gwwnmF+LtBZzZEMTvW
d7BC1199+YAPpO3CLNZ3yC6tfFFTC6NXcCN2of6I25ErM4d3d3Wlvk0EVpYAzt19
SI+dSqHm6xynxrIiVAthXvv/RO2qDiKK4w/2f67Cu6nMXNwbVjh75Oj/WFBPydiW
FJ8D4TWxX8QqpPxLepZuZ3Kla6FaB2Ps25l1ibjiVlAf5SMuYQ3r67p2fPiORv3N
yg4TRf2QFRF7R3i4AXt18dFQlTQj8AoATCdyAK/ebHv/eZB19o2AYurARhSrLe0N
twwaz7KYi9e7OGVkN9neiBgRfYZs/DU+SrwxOgEZ4mzoGwOQOBpIhTKNht9vL/ha
rd90H2M6LL2UET2G85UqKujgUBhxxqMjEqW83DlyXUvOvixZplF25zlGRgSaKgWd
x79gKJJPHY2wJILHv7aIQyLqsFV39y2fms3/dDqctG4fF+XKx7jfcaOvqRQsMb7D
+0IZ0PaTzCAjwLCG3O/0Qm/oDJDHF5zA0lnAL1UV/3+qwSepk8+1wQLDRvPiwjit
vT9VzoDOT8oovsrncL1vaCItGORJcF+RJ18sZU0tpj5h2qetUVm671eODuqgBQlQ
HkIFi38YmgM59jIXJZ7FkFZ/0/hOB/yqhiEwtIMK7XPkgGxkyCHyOgiVjl5E3/e1
kCNGeEdjVLuRQXrsSY0+Q49yXCXLSnRluLGrSK6U+yZERFX7w63Obb+m/YALiPWO
Z1XCH+Fbpz92ycqITQ6k7xap13wYMOT04wyAAk6r2jBWfL/ToVePY3MTgmwoCTEo
3b/ARWg3dTCnvOoPMeFmN0m3yQbUWzZpCK9/LKZhkqMWxOdv+yxF41eaXPD93+PX
nhGVzwh6Wzc12BWxYducxRMh78I5QIENFySoomcyUxgFx+vdKN7/Mzsp2mCeOt6v
EHNXGvQn8I1U0PnHDnrRwcRUxdh+lHfPitWl7HXKy6fPCNrNkLUNSeNPIufG3yzA
iyuEWwHdjOmnDP8W3TPeUPiVnW25NOYpG6NRFu37jz+wH3BeXgZwMgJzkLNbC6Qr
eCScZs/9LvMYQnos2yT1Ba7GKnc/iFTVCJFduYv3UyhHhG5tGoO/sTjpOHXfJ7MT
6QABd8bYTDZ+vrjZ2MKLOoa5t0nEQlGDoX5/BGZTWZhnFt0+GTxcnR0+d2XPB6Qs
bVMEImVJ7Uc1vBhUV3SHQPlJIV6HaXRiOji+E8zro/4at4xbZUroyCpwXypbJ54l
B9oBXze2dTr9mLX+8sP5X8F4/05gs22J0paic5/JcnRjucXPEGvwRHPtqBnSl72D
JzYcbz9Xo7ByxrDXZAwCvuzZ/2FlKrSPvabX77FgdMuPJyzQGEv4nTnyeYLn0E75
elISZkYqXMkOJzOFiboDwsxj/jv1ZsoeSKLh3TKkm94M5X5fYT9ys5H62+HjOE9p
aD4b1UyN06tetGawqI6vqH6drcnu+bBUtiekWeGk1GfInmt5bPeZF0WYCBDnOHlw
FYc9NjNQWu37BIE3HsHdDzL/iWvz+An1JsuyK4tYipu1pj0fJJ+tZ53AuzR1agd2
wQM9cdOtZCO8y+McJHf3F2EQPbkDv/6hGbvqLhpsbYh1ucAUj1TXU4wj0NypWadn
YujU38XvrJ718/eM+lWYkPUkUVhhN7lK/C/+BaDB0FzTmgv7Oa6t9XTL+5SZxifZ
zIYObeamr1wcj+t9uaWcFOPk8KgtB0nFMPxDwyfFDPkIg6gannnn4zRbvBnjwD1/
hczoIHTbPDEu27eLt3oE/M1gOv3Nv9RLZNEYuScCmv0uttnxYQZkWgZuddEEBpa0
rPfsJjDCC7ACzWXnFF28FbWJKLhwvggYWOeUyPzxC4EW7sL9sAL3W0h3sVrf7fxv
xIQixO8WR0wGTar7f2dxcz/ee7/HBdFQm8gA3aZKijT14sqt/nwwN0gt56WqfEqk
TF9TFzi8x17Q7hw8EG2hnWH7NyaugjU9SnLikCtNPef6zZ6cI4+3awPgYpvRTzYI
vuyrofpoNZa8bDAVM1M4oS3rZcCOn1kfITVFU/HVWRuxeqTli82AVhW2hdbh+SNR
LUwjC27rKo95uqCEdoVpgo5/jtsrou7c9GsfSViNoLDtUf+repGRfddv61DX0knw
Oq9Im5UOuM9LfW9K0u+12xH2HZBxqxqCVFkYSEw1PTZHQRAlP2RDCmRpPeH028Ys
um0jXklUTp6O6tD6Ak5mmIwYNhh9y6PkKUxeW7kNuUwKgNVPukK8k63EwKMnxTcM
vUzAlymsUq9lT/zJNy9yBPaVbbJbYYHUC3WygGSn4WY6LTEBqVLYcIMqA2XLO5bs
7A37JXLYk8zu1CiDLY0+awCLivEaXCwjBCwaIDO8R1fLV5Pp946YDRqpkJKacP9F
krCvV25AhCek71PTYA7UI7oSQ2orSoGZlLgSQMhwzEoP8EclUSApsUqjqTNW2YY8
/wuKm7bjV6EqZnpuhnvP4dkXyqO38R+eR06hCap1lLARCrHnZgFgXlZo7tJIyGdn
IRKeXLhiwMEF4vWUT+7XtZc+0cOCGNcv8KMzC7kIvleXg3Wj4lvwVbvV7HKPoVDR
awdtukfP6KkrQM4iTT/PdHLzS+eHV+T4tULm9fKn/YvzTUnJlWJAXEQB6+qmGiUW
rMwLeGV7DvJGGiySPcgg7Nw9cPsAx7S18Y+VN9wlq2OozPPoK3k8oH8jVT/o+fNZ
joxya9ssiyy5n8e+z0kujLNDYWpBmo7X+EVm1Cj/yVvBjxmKbywdktT/UseZTHD/
EVJp46fMe6+jXcq5PICI71auHKqgpmLzVZN893bwoYLPR24Zth2662/8i96BFwsX
qI7kMVF9lvh1vxMy2aXc4XQvLCjoRGDf5yjq2SvSSPqcEdYwxS4XmK3jhClZkf2r
MGyvGZPWXT4mWsZCGXHglPfKbIAju/bcYb6Ttw+AEgkG2ekZSFDhPpO4AfNvQsGs
7ysKtwiWiaPCyqhvI4U3N1ufIa8F3bJhJSOLLRQqObzOA5EWfKLBwD0Y3r5+5LfC
EqsF73Rhf0wbnnvy44I2JV3QG66eAOHFl02EBcGA7RkqOmhR5Xa1wXBgF9K6Jb9Z
gvEOe7PnzRFTANogTa7jNOFGtw+pS6DqCUQj8WTIkRvr65Aj2vaUm/g+5rO3t1E1
McfHY7gJCQH/Z9PVZ+/hCc1Y0RAq6/mcDpNnUSjimh1qRNWXxGUSJJ9D3lFz0fcg
0EKt9+obA5iLJrOt+uAXdAqo7RP9rLUdJ4EqCIeFbI7bD49yzj4enIyy/JST9sLv
CU3KzGcb/rupD4l07Mbk8HsxUePeiSXID+NUHy6XJZdOLeisNERlyLsZx86jB0ZQ
mctR0EtsEg983noHOSl3HtAyk2rqTY/9pDKEVEj0HyDDiB6suLX9WpJjf8fKcLOx
RBU7Pa8HChbMQ9wLrMcOZo2JpuMXmi8CvjaEEKZ56LJyeSvKB6i+6TebW39VAKKK
s1HIx7eXemTdwcwisudbF9wIcKaEf/B6JIZJY8rXyByxyOGc1YM5NXx4HWWilBa2
E870V11TT677sQjnKZOIlqBrkHibKVy2w3L7+wnxGjT9CSFodws5m0h0WeI4iF5E
Fr+XJFN78fnXq1x0bRKuRK8hfN/nOkFS4/H8+sWGW5m9IozxfWMSRO3FBA1FTp6j
OA/iR+CaGNO/Mqo+3b+hV6EHnNqxGzoUUj1Kt1Smm4h5wSRmWkIuJtDAQ5rvqB3F
q0IKWmKg6bqPT9ToFB8/XWDHNIynFt/9gPKxcxRvvU1XsufwkDudE4xNvOJkc2PL
CiZmHj5GXy1QOBYWDEGOqEgycvyyca/RoEZOzc8seCEJOFj9KeObFS3cB5RsZIkj
b8qEiFoANQs2jJQwMwEDDOxtU+VJ6fHfpoqiATu/ZayYVTdlRXQU/u9v/SOMZUsF
hQJDSuli0Sc93D43J1hWFulOG8530B3FQWRcxfiOTlANc/OzRnbhSyNoZGqfwPgR
dlukcN3vUdmQob2v2kO9YAY04yp2Sna/46Sopv0xBUbAxeE/TK1wszEZAiKj8e+g
SXnAEaADMeIWMK8P7mcnq1DIpvpy6rXYlCIZ3cOGXlQ2yCMW/sSxzxBqNyI5ihPH
B0A3bInrbEIxCdZTPWLmvcsO4aTM4cTgllUpQg+5brQhBg/gBzEGNkTeWerfxPTE
0R92JdpOiHUja5bLPHBshjiexjqcL5my7/2c2yz9DfUoaMLiYFvLiNxMvGDlVjJY
VnRqPYJtblktGa5fdCXzeWnzSI2/XTXvlJVRBiHrFz7rQGygpEV186ze5+I0Tik9
F3FlDmTQC03PXV1xg2ElrxGhjOBex+haMIEccRsFyxzcf9tyusmjL7qR3mkWEvXX
NZiO/vD2tJ1nYuSVsHM50cSHoGVM3qLd2V+4niisCI/9SSYE9hAhQ2JKFX8mjEa0
61jP60RWO848Ml8MPdxAxRj6Pc9oR/ZfDmEAddN62VHC7w54T/rokIdH6LZC7AM3
9OCB/A2QgXXCUU8snqsHEXZ5LdGPHkLnZmMhs0457vMhoM42YEbR9PqzeuWEq205
L79k1a9/wqfZ1HEypWXzXCUaaFQL0aG9VzytkSCdEgSK+CRKPRG7y9OIK3gJ52kO
Z4q9EpTgex/6gexpo8R8sbDTmis9kUBdkNc5UmPe9Tv1rqDAxcwVG1v2xPjTfy6t
mtWDJROdp6K89q0y48mdDAMHjrFtLuM95Q4GV87qzSo+ZdWl8RAjhIvCDGeBacdG
0v9D5s/s7bGYM1F56ni2OhC1VZSvDDc+Ap8SkDNwo6mpsTp4go7ZGHNi3Th9f3Sp
q6Hx35rMmUVITMFF0n6unOc/mVO0+pA+tiQ7zAQfkANCjCPH8czJD+hUyrNqntgv
H4P3eJZADKCC3IBetf7RO0rd/r8lDPD2c8fAFZ5gFCf0ZQdqurbJSOr4opBMj7Wd
EEQGA2g3nLmomUDw8SKj8JmfTSzwc6No0HGPDxSmeKdCkj4z4DyZhOaZbXa+k+EE
1HElI34Cjc2LZczdWnfvfCLgxjiY/2+owFSCk5TRt7EBsvySoXp2f0IVmR5bdZld
ziK4mYoUEFfHPjrvjwy1EN6jJCr6u9+qDz4RELUu2dk5IT8B+ub8yVSBnN+WKwpj
TGL537iAXa3u+vR4OLGdba7Y/YGDu5Fs1twO1z2TGpC8iuMkfjS/IRCALYTfnvFC
2LUxS+lWtht8EED59eLiR+OoKQpRcYtR0YeKnB0m+V8sDFxa3LcsB1UFK8uwA/SJ
YBhXO5Z8X5yRkO4ZM3/6gM3Jw5YrQFXAg8fYmGwPPaS4wjgpYebc2m+BzwfBz2FT
dJqKd5UUTUeuvqZMM3EU4mKlkVMcom8dH/6/0LzP2qXNEc9UmhCLzLnt1LGOOvWf
bjSPKxo9TTWLBWxMyImA/9VS2f5mEaem0MyZniaT0uAD7SKnWNqnV1uKJ/n1oXog
1vFwVkIiqmIpCsUxgRGBUjIJvRAkoH+ziOEvNwRJvd4+GGJTmNMg0CkTf3Ltl66G
bb6Vjq3pBc4+SN+0oFgBxhQmEqfFwkCHSEMtHYWwVCKxaZxoiLv5RDO/Cig7A1so
xfGQCpeRHLZd3FcSNfoxZ6VAefYA5XfGPiY70GyLfWBR5GgiD2NTwzAeeZ9qhzRE
/liKN7KDzaL31FGyRa6Lc8YzrFJz6ist7cNHFmtUQnU/2teGAal+VAkB8YtiFXcZ
bFd/7qJywRIJbv2w/4p+JdzRmWrNcPeG7CtpVCd3pdcUzXYQXajOu59DKBq8DX38
ZvAgY/iF5qToky0CWi6IOIaYRF0/Fin0AgDieGeLDqElOSr3YpxeTYbPB22aPiar
FND3ycmeQEEdGW77zXJQyOyg2FWKkpgAWllGm/p0Oh+N+XC7PtZCANm55dy/cWGc
nuZnpttXNBFiZBnnx1SoluUuYrHCgXdbDMaiUABowzmv8Fe3kCcK3QN+V/E1IDGz
yY2S2cJ75BxiRqM36ewKKif5TUgTQcF8lSbqW/6cnAoRdIz7pvygG0lGGAVwUNBh
Z8dGdJbVuC6/68FMzT8Q3wy3KQ2oLBerO7NZ6RG2IElc3UWP62UuUk6dNbxgkpTt
pJYFrCKXe5bUD9zbk8tc/P/y2OtBsx9FAEezg23Nj+x/xCYl01WPez2tiFf7YqZd
6gSVtqIWT6+XOoG7b9abiK2i61sBOsWAa0dvCa5MkTVZz4P511QfKD4yavlG1mxS
sOCKuFIuMNxJXHRmAygD2f8M78QDWl+UWDw6gazv1FEyvogl82pq4Dz+Yo86Eic0
IWOmNoeSL/fxvGnGN/1cXheNorekOmanqcoMEkMKMnB0Cqty6Tb4m9l2frndeZql
EyuznJn+WYsnV1Zgt2CPK+DrGxR+6tQD7IC8w/fAaYcFexVxBtIB10HtOImRKW5Z
cJnhGp4MRo5Llb/fTIk6Aam4bFVupGuuij1ti+/Ct69CX5OoHLrsz2+dr2YZQIGR
cknlHkkkXUzvwDBMkq7ktficWjHqFIa8eqyvi+FdIuUuG25H0xbLFLm6UjNQE6G0
2EWzxsVVr3i0ZWpqtnolA+TxTsw0Fcff/NZh7hjrJd6y5YIceAxC0/XsAlJbgRZC
tC6ka1/5sG6Z3cDMSraZ0VteiZT7RvWQ+RBfdQ5uP2o9qRxiYKbzR1oNkTf/S4q2
YsTo0TzHq7ChD3vKgaGXsSACua45spZWpah5Po3GHzddvyhWrb2bXnqHLPTI8NKg
6X9eq7/YSXz/t3Am+1U1uC3OejohnqLmQcn0XzAq9dOIam8/Fm1mJycmIJIk9y70
7s2oFaXc1gSsKCyW/6/fj+fYJgHXJHI4FrXYi/aU0zYWbDrjk5j+Fe7DWhXUznd0
3Zh8EoYl34VTWADfsVwgTzv6odV43GOTdj0jbiBwL6GE6eIhvdRtWrVbXBWP+9Kk
VBk1rFM+M4Q29GDTHVA5jnb5AZQvICKSxh4y0KNtdbYp+pWLLpWg1K1mat7AoOY7
5a3WezubqptvohFCL+ckwo0Cc6U0iiRDauA8HJ8rHSP++IPRkjFo1Kqf3zV9xbXU
seoDSfz+T615vGoKnZcbD62L3J2RKLpEGOGNUvFGMUX7OHgzQWrMDTNHz/zd2Qx4
lFWE1P/8EHolAXsRkjR/nb5q0R6WIjwadb5RiiQvCUD+p+xEh7bbIuO5xvLpwWZW
Kgo5YkJNbVt39QoRXDHnnKr6ewcdeo2VchSaFYGXg3LWzRvb8tyLGnyny0UTA1pF
bOcilONHbhfSC5qVM5ZuUT6ZL/VRlkaiWofwgwjnW3Dh+TUJY1vawFlpFyASOhal
5VFxXP/+79ELb6HOjMJ+hNorfriW/t8E36RR+arxe+plGuN7mHjXVIx9khoBKjnP
6TH/TaZWOpNL/SaX+epUs2HcB6gltn6JGicbLzLtJfgJcqhBJfripJmvRYOFsNdz
va9Uv0Uy3khiK61cG9hXU3YrjILiRdFga6AGQGb9HANrBfvTtmZpOfSj+2sl8XOt
GZ1wKlGzkVmo91nvJHUNTFFunPoJQDBY3vURtxZRWsYSMkFnyts4Ws1WtWZ4kjRx
fGGCefZHzLl+wJONNYsAAIOPtfpyQms1LGfqvs0yu8jwIIFkzDr9ccLRxTtS3gic
IKMwLrhGM6dcfdi22Uez869dQ5D0+mkJhJSWi5NeiCRpZSJmmdt1/OV6xvtcdvyQ
SPaywqJe1yga8A0ax3Jvi6K0wmPK3krz5+hcti5/Baq3vls0tUHaI8B/0/JUEWLu
N91I30E6+4Z5xZpxdOSFp5xQ/SFJCG4AsueNf+iO19jL2Oxk7MzimsKN4EnSTPbL
Va0Z/yihM0cOajCM6yWmd2MbrPpeX3b7aueZrUyv0PmkxwMr7fGEAc2ANQRaXfYP
J21NimPPIZD6CRHpr7hccqIBRNoDIuOt+w6nFjluwJ5RgiONNBdZqlmd/qW4bPA7
9/8PTeAHcUnCVCdN+N0smV07KeYUiD3G6UU9yOs3FqbZlbQ3nuIiGA9DjnynJEYt
6jNIQdnjKpHPr27MOEEvjA6VGCajkpOeGTAQUGzp++1Bz/H4BnimR03yMa97fc+6
wDsib+mu9AjPFUEqvlvmcX0TzR/MwzLkto6XGEjeu5s7tltGg+wMNF+RDTRe5rEO
y0pw7actGWQSS7M/nMuqQYi1lRR0IeA4+pFy8Em3ATIbnsAm2Xr3zh2YO+x1lJ4R
Ow8WxHXRw6v+Twvt6l70zuzKQybHPYI+s4PuQaMb/GqpA2jxWvADqK4bpKhPP8nn
VSAvj5m354a0NqWu2+/GeU5tOapGnbFML4XInd2bI+UWRvBHOZjto4tCA026Uuuk
Lwy/oUACt2szrLLRRtq/V0oZsE2BQezDNi1LJLyEKaDfPBHX+WHOe1rJte+IBgjO
1bu7LWxEbTjJXohVtY4Oqb6CiZ+e+P0r44rgtr7wvuG0GYpOpSCbcKavDxgXkEyZ
0g+AubLHh2oJUnRGZE8VhmcUTXPVlXx156iRS4uKZdkIA5MgeBDzKBQcucWGMYst
PYZW9l8CkPDXOs747cfXQp+8f0WDtR2g3SiFNxXbk7JBPjCJ+WHkY/tstmfFQ07a
Wo9decCJ09XOZnKraxnd5lRR3Tc5/h5ZuKmXVzI/FSKmuOiSvH+B4RgyKy8tMBT6
Z0XXDtyZmnQLJakDNLb93C5QjAM6qu3I8N3LVPyvHLQdI/fhz/kc9N3HQRxC26h+
MxmxPbF5jYVtRIvNSLTZPuGj3Jw2MlQkV8YZIlLreGgEc+h0kTWRmBSThAEL+jub
AxBKt7wvJFQpMD+lNCCSu7n83ZUJcH7b6LlvQdIx1xF6l9RAlEQ9hr5G1k6xCV7g
NVYc2dwmYPXFcmImhhRxoXONuRC2sfpsEQs5M4YpjLwh4Rgfrcfg8OdGG312efxB
1WthEWveP/XvDYSGghaXqBVH8hks1XQRpmLD+VBoo1R4+PmWFP/wjaZEK1i0Gc54
gsP2BEWzCO1KAcB5nDkk+FybuOaDEVcxfJnMwFMt+MLzrpcIP4U2sEjpDjxydl6Y
QDbaQKNSXU0pVoqkdpBqTSPjPrCWzDykV82UZkzZEPLQRueZr7roVNWGA0+hGvdu
2qw6Y1M/JVoWSm4jBFTHQEYVU5L3mPF71Uc9zRui4DgDscka/vOZXVUSTTT1cfX8
0QvWNm3eb72VZL6FqGqZ6swynrOL/yu7rfZhaY2dlEipqxtLzukXwGbEkevfBjB4
wJTC0MKmG6WtMA8ue/37yrSTd131XyfkKHBXrnIKiab1m8PdXuYrfgcSWfkZAeZs
9vjJ2bav+Cj0Qq1Q1IfgWpG94ihh0UAOGUndkDGqXmOfsjnFvX2fPrQ+YRTltneb
1VkAslhqDxxA56x9UtMFDajHUvh3OwMVdWhmXXpwDJJzFKBomblFqy71KdM3Pkax
zOQaSvZWDLxlK/G0Bsgv5HS5qHETX5jIuo6e653Qoo4PwAbN4Hw7XrEkwOYUZgLc
pgpcsp5mVQv2OSqPC6HMo308OhyEOu0OvF2I6Igk0UOCOLopEYH7vt9vMFJiF8m7
GvFgLgVSk3Nu9s6pLd3egtZ/+Hv9/o6VOons9vj4klQyvMdv8DXeH56nXomso0eK
gXl6sOa0lw5fWquRFN1qASpIOsEbQ9FGhzPATdTpYAZ2Oovs+9/EA0asHCgTW3UO
dQ/m3F57Jgzu32cJnJ0mnTPTO0UDYQf6LYojPHyRkduF9udQimlweX9F3jToBaDo
81QQZXqeeIC9RojK+sjbGqtJ4z9HGl7v3VQXHDn0xR/A/ZMiqp1whg0U//43toYM
tFYVde1V8EZMoygksGQMxStQd32QX0jrbJwoIkcV0/H4qV9LQ+TxUbniXUW0zQJR
0TjY65VhDlPFw9R2jMTrQwasEL4E4shR+Xg+f+F9hA18Ejn7FN9QFrlgdqo06dhu
SpbWJCcco8LV/4ZVfzzjk17jST6mS0hU68Ea5tj6vyHYr6y4obQ0vaYZ2ArzpCFU
mVLrSPESApN6VJ+D+vMGaMeJzjsGpPXJTKki5mPC+OznfGkuUlB6l9WIhk3NA0V8
MoB2iF1GqtxmM10D5dP7MBXdnXsyZ+42czAwNuCT/MJzBPOODU+ufhvdxMsIlS5r
ZOs+XTD+N+UYJw0DKXgRcxeggZRcinaSEwqR+3OzWwbQ0ZV/N3s+let2Cmf7mArY
DLE+5U7xiQ3vpo68WGlcJ/+6GPoFppj7otthSoqrcKV3T444rXxUdppduq/pHXaf
SzBiU2FJiD29ZrjLDTpIKop+dpDmT6fKc0M+Io0swvcexwpcgkEUOAKSLaCxMQz7
Rr819TuL+vy4adGMHaq1768xctTKp9owUMmzZZFdJmHWYBRFb1c32dE+ADNSNdgv
uM9sGob4dAKo5LrXeYwu+z5Q1wP+Bfve/WEF+excTmO+WC92nGe+9iyQ+rxpC4Rz
wBlRYq8wmzrAsMBBfj9ZbN2IgW8nA3bBNnKwa6wzrwY9LkfXDBBe9aCgoSzYVxlZ
/8MUdlLrFGq97VqoF6BS5EdssL7vjke49vuxWArlerGgDG+s6dnc6oIOEol3Cm2/
s7pUwVit7hEmSAn2NE4b+hxr3/cZivtJGBbgqIccRbjL8D9lyXf7iQZDzhSYdh2K
HjeLrLMfq+cF/gHstph6dZPScEBWTSuNuF4TFfKE+NZDb8H9dbR0VUhziPmxLh13
3ix0qPpEvIP2VOPm5JQSPCm0CEpj+NvyF19KQAuHtKWNiLiK1tDbUu6pCg8MApSX
VL/oznvF1n8njUDKbZ0FOMdrZeRj0D646ks2CrLxYeY0pp+QfS8NxR843qWtQD0W
OSbzQcDjy4pzC1TenpoyVUzIaBbMCufu2PGUcFLydgudobhn9qZMZD4Sr6RMbB9j
lw+4M4jVxVafE0+5gUEjhvoT1q1F9gxscCmVBuShBfCzSC6+oCQFZFgS8v6A7iGJ
53JvkstUqv++5nfVDjKCx24ppHbFCFZQ2d8cKLzgDH31mdEf6eHYkmzEnRdpM+sW
2bfqDl+DUQICqHXDgU0zucs+kmxqgT0qjGYa7cNMfeje8GSYSLMJ5FxdhUX4U452
WMC+GOTJBMXcZLtgcXyaSOFcRaJz1c8hf1hT43AoN59De3I9hzpXZoSPW2AB9WyJ
VaxZns2ATzC59w/fjmyPIUBoSfMsIahq48H0l/0vTGJtPOmOTqK66N+JyRi7wp4/
oEdkghbYEEOI/NIQ8KuCaHCXrk+4nUzu+akSJZbI6xfdyzJ4UFg8lcOyMwM/RCXw
VBcjjA/5bd8zqIn0mBhGx5EXYMX80o5NsvmGbrukj3HmdMQ5HlNh/h/c0k1Cgv7M
eQMFa2cZeynZp3ZZzhCtmXGxSTo9Cs8JbpRa+UtXmCPXwlVbgOlHhIPnpAYuI+10
78QD7/BXZxJ4xfEqnHNJjcJFV3CGwZV1DB9q+Uqcwl2S33jJKhbm1DBw2D8BcPij
LEVRM3n8JpZ1scE48y+FMLw4cUzqLyGZjNd/8WpleVkUU2D6bU2D49yNvmHBXFoy
y/XB4/WZoR8ffQOrOYdRlSlxx+AZD1jHNBE+NGc0bVidRpL+1xT27eGBXJ0EJlqI
qKupVUyRbi5yemlUId2lHgHvzFU/C9n3Tuj22n6590TksHp/E4UDRO2I+iD5mUmN
zszGsZodHMP4DpShmNY+J4fEZQA4md63zZ2/wJwAp6U/kwUKfV7BMY9TmDg6K4mq
BX41Uc5QwYdeYK8Rl/8envATB/c0ybsT6ch8U6Ls29LUzc5cQfOa4+Map24S5J1P
2Fptp4JiLgLkOe68mCVi5N1OOHuBg6NJMWqhtlzaKziAJNP1N1EuLrkaIREy6eNS
ABmvDZak2CJW9qt+UCfuXJvdwh6whLJ1u0XEIwtQ1gUiF/z+nvFCdP3dczFGhO+6
rW6a73XSTgJKDQ1usMwAszjQVCBNhctXwQLHfA4mK/wyoTzPWpDO0kowqvNhGNqp
A5vIsUA93gKBXm2o1ONfptG+0JdBBRYZkeEsg4CW1JIy4aAfRYuD6wkxAWzUCxUK
yFsRzOdd0mhgayU1Qm74++n+wXKruhWfFLeFbY+YTbo95TcIIP+x7TFpl+ONn4oV
jpToH/Xc8uCuGEMiwFLcgtH7trZBLE6mPvBiSlJNA2pd4zQV++Erxjt30C4JJbUB
x7tvbiqpPKFspzYDq7jq6L/1iDhqvo4vphX2iIAIVI9WRjWSQPXXTJQw1Nochs67
321Yccy1PTqVTaKWWZIV3VmIt5iN85XzGePSwQYqi1M3zvtBtokrkuWG0rj1hzte
kQhsd8yZn2LFjrVm5X844xs5xx2BBfEqAwulRwwU0g9QgLDy9HwDnwBf13QpIZF+
d0tR1tZ7khawfclTf4oC2L/vj5sZsxxYAr9uy8ZHQbaDgyadZoRYBL1o+mzS+UXJ
xQ1tWtQTHm43oyvz9M7bgD+P4MVJpU+/f/A51Yc2Np+s8112fiFWgIFdlAclRz+3
vKs2c2jxUS1Z/fIHdzRpqHSrFW7h5uHecdqomdwRHXXt/Y5CzKwD3kGzCaBgkx/4
9qbq6PGstdz8XherI4i+5oPIUXisMG5YE3qnHQHpptBnBp9CSZBd4HWUZkaOC2ZK
aO0KM3KbMQ8mOeeAiVWQ0J4T+moKWqKzQwYA5vPwvXLMk5dRLN7dkkLMCBmTkrPK
DCFzVP799iKxiwkHbSQBFANIweDYxmjci/w+Hx/rxr29pu2B5jmvfIlkPpWkdzhv
u/4Nqsb7a4For7fdlUll1jvK1yiRUg+Nctr8yBiTUZmwO5NBEzHwxOt/p21Nr58k
wNfhHQwv7lXdT9byforoqjCR9panXeKPY07XICYYrMOo8HCYcmxTJ4fWM+jrIIPi
iwzzKcgUPEPRLjpUmOs5wg9BWgajuGJrbmdgbJ0XNDPg5QsA3MNW/U6kx9qS7NmN
yrEsJGEJ5+3H6E1rrjPfC9HGXxZSTWI5svwgbLdFM+IZSO92G3jiTdLcUArXVc+c
Rq6mJII4HbMDjFQtVkJuHNlvGq1ulzyNSIlx1npAYjgG6O7eyyc51HqmsOHCCUWz
nii+n17jooe+Me1Pm/GbjcmqTodoR6xhtHTxhTFYOaPj2/jFGmFgqC1n3jYztE8H
S2tsgn4konzXLc/tyGlODKB/Tl/Qsq1AOPgJgb4GbcTufXQQ95g58ZvOBFSFWY3h
V0/lZ7alOfYa0FvgAO5tqaFtmXGqxfRpxOwx3wSjFOVSsEQnFtMp2s/JKjeyfUOr
AY33NXnknBDt87POMuxODTstrTs+pVMpQjLKp0t+phj+NWkyoey4/6Sg/DlKZr9V
uPHa/ipPtzHPFX38ab9EXCCyl9NDaQDmzB3gZppfnGgTMGlKdA2kUXkkxVmaEVLR
RCTbrg6J//IgXxyvBnq18d2kEV3zzG0rwdbePgNyAH8Xm6TrTUpfVWAnxcwcsxiS
ODokk91A7D3Lgda1YKG/b1OYrl42cOWZkkpvmQxLhlYpQiIwF89kxDMTGijqmhcG
MlW/cosBp2NMFQX2TnTFSn+f1CBswDbitM0MD0zUmUivQcOZekk3HRmugUdvbS3+
4sL0HXVjpV6HZs6+kYZV5KLFFsF1ukYwUNgxy7qNoCxjYl6NVxdavL/pAIa/nR1C
5qcEf4Z0ukYgrcUNA73wQacXA9hL5/75WmpG6VpFxILFyuA4BJ7BfUk0jYywPZ/A
vjnEvglmveMOe04Bjk+VndJ66Zr2AJYIHFb8CH/wJ9rAzssBleowQPC0XAkAEN7P
OQQ3Wd1Q2JozfTK0VSfOFizUbKZsmSI/gt1EeG+QrMVjpMnGi+r2pUdNjgrb9eyq
ZIQSwFCUbHUX5sDDMP3vymT4XeeKKxWRwI/5qe9YNgt94XIjjyeNSlpAjnx85sVi
n78tTR3t4MwDlA/7OCS9reudqaZdYMzWT609mYgAmKgsnBZ2BjMUOMM88CJqkAPX
kY1QmLyDrIYwDHipjKC52XfiTOYvl0rEcgbZ2xw3puaW42UOwGTD4e2/k14LZnlv
BTaC0rB4m5lnV+VzVWqLS36UUBh0WxC4hHOPKh31xUDgrfqPWE7C8fZRvz6nHcDy
pASlwOCxE+veb8WNX4TvVtFIZ5kZBz1tyNYG3iagZU1gYWG1KlgaLdmQx9zu9Hqm
99zNgqI7pYLAMgflfgSEhTzsmqaAAnBFEv7ruDD/8k0xdg2c2pdS27Pe4W6H2Xe8
1wfqy4Lu+NXwXsIDWeg0O4mUWQy4H45pNQFi0vPwsk1tkKKC3ZLd6wFR/XAwPtRi
Fn409v6XXMZJnNWoOeOqKGcrD2p3QB3FvKgR0pkzoxu9FSLcvziWTJYKm/7KJxlb
Cy1C2R9TOcnI6B5Vqj+6eCZKOtkvM7oeRYd8F1wEIyDllrTFqSCBUYULiK0Ox6mc
gCY7gDqGYzWnoU3isRMTLBXEDYE3fki4KWZt/3FdV7iGPTjL8bKzqdPreELwLYfM
EwG/uIYpNQRFEH87PG8AM6UzSqixqqIHB2jdUollC9BDVHVLoUfAGcptvvNtwyko
WUKaSX16+bRtnPKZTctq+jLaNHb+J+t/b7+tb0RjZh9Fd0vkuSJ8xqZcKeA0HVm/
Nkt8vRCiHJ8fPmzRvtms6zkgzl5q8oGpQqIN0zpyt/Ey8DcPWoqAT+v5P6s0jHH1
XFate2sPcfosY4yr+FoSrCxtjvCUzO3Al45D5OlLM2qpmAa0PqSDAmoI/Q8lB7WR
UBAG1eKu+JxlQQqANxuXHYDxLzGT5UbrhZLeokCvNbBwkyAQx/jE4PrmYwI0Uwna
0+qMhvcK3JZz4SOWfVHII0LEUc5dutuJNBbWbY/+5YNgX4DwP+QfD/KyknWTME21
ocgoezqVrSAeemJuv/sdLc9sAKBDVV61ubGAJfUMoLgjE7mjSUUWHFaleZ8TIVRz
/3NjqygBuTXFslBuZQqeB/OGW/GSy+L2FZrO1XyF0d5pMNJqwkasSbn+z7+ADnBG
S9eh5zm3xR1Ts4kXSqKNI8W+w1S1qEifseTBCKKwRRfL/GVyQ010botDDqXIfKo3
joYCtnMsDR3m8k+Mmwvk1M/EtSrWhcpwOwyZQSqKQaHIVylWqZ7KUjKKIQWtFxyT
RfyJqD9slz2XsJikid/ELoBO8P3pjsYhj1ivoimOxU5HLEiFE96MI/ibr0N3fEeA
MJmoEceYvHhE4WQoxSuCKlDvGilU673FnXb2aw9/QUyfPWgATpVTkXnotF06tW0M
yfcpkgOzTE7dcA5FE4fwTQo+DvDGAhZhiXpTNLeH9w899lRw48GEqeQAQfHhMFdV
ME7EtGMQA6FBrSCGlfeHUcBfaR5zV6/xpMKDCBk4EpHHU+9+Qci8aGH2D4YtVEr4
13/Q5nPhzP7NUad5gvZnhLMhUThoZfik8MV/rR0MSDgvcLgRjhr1zdGI0dEqQzn/
TRUwNpIMSkJaGNeiu0y5shkbusnqDklG9oV2pzfXQEInM/zmcJI5uwYUjIV7PXl6
7LtGFO6j6tB149QtkvzOOBMry9Alsnk3wPehSfSMQTDSmy8Ml9gtav6UNMsCdJb8
S7eGF7bP7MiqAx14lx7tSDloTy6igN7gOm/us02rtl1YH50M1xRE3IB/o8vI86UF
INmtxP37ek2SyAW7L7mRcpVY2QFI8EiGQgyNroRBhy/1Wqi1qrLlLohqZW01a5XI
/ZoJfk7BzqZ9gxulVGC1rZ5SnE8lU0cfCmAjxmdnwL72fM7sKccuUia1nyGAY99Z
R36u5THRMFX/YmtkhyZfUpLjb8pYPMTEW/E1tPkT3sD6KvsFmR7Nuy8BbMJ1K1wn
FPMa/WXwR+gBlT/WTDTe+8YUIjhsY0RNSMdU1tWtiGbMTxZ5BqW021mKum8wKBP9
DgXr8kCzQIJtN/L8zJLSpUJsqWk6nVQ4R5eMrfh1nUqV7PQ9JMF9GW6cGey257xX
c5YxlLJvE5ncV5wBMgpbmbBj/JyJxPQldWLDVnHb4k7SyilxKjIXW9A1tdbNE2T9
LfUgMipu9RbrEZEGD4ru2OKJY61I4ZGylTFTnJMZs/lY6PfNgC91Xo0fvTiJvq2N
FjIKKaC8eNqu8cPgcDVuj07IkizaGDOhOzNchIOgY+uTHaxe6uakwwP5jxEoJzcu
Fns+I1EWYtiaDrtvUcI0jjN7jJmhKzwM8XXlgf/qOEWXPMSHNtvvF8cqMWyWCXiZ
W0UHISSRaM2ZwfVf4TyIwnu907eorW/heGV0Ce58j5G0ktb7s6TFKxImZc2SfhDO
d4XBe+pgigsZqaePwAcyZcakK3po3N3nFPbwlugeiTWNRnzRK8+0lQiPX87I8C/f
CwjjLEJr1S5wV/lHwdHveXMfRAq1xDLS2Q/p2Ct3bjO3noNhWpMY+tm4IcvvDrUz
ndZoDkFK4xdV0KIcwZu6DziEIPBQa1PkA4jwblH7DJ98lW4cAsGXe7TnaH917KLA
sqiRJHbPoeBCB/ZYpmPt7hpcnzW4Sc+h9ziOOtZOxWF0G8pb+bKuEMfLbRm2rUsa
ezT8wuqsB7vt8V+Ab1lHFKay5EqMiCMAIy9XCLETCrl3vO8lpWfM/NwVjzJOg8U/
ndIaDJk5KN2M5t60pGMTVhMZWn9nPr/hNdCPs0UPt9v9cvCI615wHdlf2Z4njEmP
zMzk6hcAFx9/nFSHxw7vRpxfzmE4daI/c/jzVZzBGh0cbq+nLY0cutwZCXU8SZ35
f1wsgkxQNg/99giRlHgisXpS0gqGCRg6Vg5IRBIRvIHJNPl5kcVKRC4C5FOTnoxM
ppXpiJdZri/vsnGCqxBy550LRun/TcuGwYJCv6ra8Fe9ivRoM3j80VgEmz1ZkFKj
9dsBdNqUneX/CiYOQ3vDH1UQSEdWLDIHs54c8ILD3TD8tJ3qD9KShfJWH23EIwjn
99bi4iOT78tqTc0lkIJdLvbV9HUnN3yLR0my88xZ2RpN7ZMlXjnZrs9+44Ysbdwt
VohW7VxL2OmP9lESKayLzYK7tqgU1lHPMlc0Bq6V1qjS+YxwMx8f/yzOHTllceRt
U4rZmTNt3se0uZShP93qpNsx7J8jixb+j6gDAoKvi1ZYPeR5kgQckPEpiYa62A2N
jJJMTlhwv4U+6iZL2H64yFx+D65z3X7/nskamaSPulhhPU6Gje7hoTdUqXagYJX9
rW98tABwBa+Co7xiXQWpbebLkkaGgeaGPlSdqbKuxSYKkxVXxhjD6YoNi8PMY35R
TEF3HpGsyjeJj6eU20uIMGji/88kO0l6FExVzp9cK60nal+28s93ohO4QPlyDLtE
Cg5lZTppP8390l7DZPTfZMkbyDUQtvptQL/eglOq8Uu+iF8VkizLUxN/bKA0t9Yi
NpKuuIMJn4Ob4GW7s4hfVWVXECbhoc2EhrluxLDLERC0hCTScn7VGopCfEZMPTQy
kwcpiQJHjDwgOZD5wXQ49XkvD0fLJELBe7RLzqyHalUtM1NePHxefGXCA5q3zsrU
BieYE+/NQlwQeHYmGt3n5FAWW5UIWrmVj0/oyXkZ86rBXB4LnK3buHUzVjJZkkdh
KRf55w52dmMamnqYqvI7hh+eypkTLEyuPySxCtix2g2ApB+JWhEbEUzwzkVcAkAj
cfaS7EecgD888fcbyxMqKJIa5+uuRozScCkC0qtLBj0AUAGdR4o966uUOI5VXHpf
jPiuB1WbrUZJplpa2aXJyUlUBu+dXcKXBk7k3p93PIDVB+d4qNcTjH1/MGK5qmzm
mTuPz2YSvfL0yzDF/kYxlO+w3hbrttMSsR4dL6kljcXLWpl23ZoBAQB8d0xomPze
SyiDutimH87sDvJGwaRJ/7uNHMSWXopzddOA5NDHCFbBJ8DzSmEgWHiYaU8zbALs
cAcf0bOENFf4ZStoQBRX5j2O02DHJvuXZM38heQYVENiaHIaco4z9gT/tH0bs4PP
VvwzTzdBhMXbYeujuNRv5jHiTZFoqMj/aSGwbzlVFCkrhS0y2sd0wyRdkGFu2kP5
os61R4OIwxH1h6MexjqcePI0syNeIRW+FF4YqA9Ybr/z32EtPeEga0fT+AQ6VsBW
cTm5SAjMZYXsx6+otoUA/s27eOitv66GErWVIlAPNN7mhUu4sqDQw3IfjkGw2pNu
9wnMrvvXYekXDrMZKm/qK1MrwifpgnEvl6xBNAWvfbGqA7+7XVEufoNv6+qPxZKQ
OQoHRszEzM/Q85LoU4VU+6ar1ItVjGZOtjPYLJrwxMh2lmq5rKEsHJ/q1yUzjYlN
tKOa9hwk9qBGXv5p1k5KVH+DLfhZt4L3ReT8ZDFeV/0jFZcemllB2fyBAeZP3R7F
3jkKvgKx4df2X6GpABblooxNZCUYwqKDEGh/2sJzzsaQ4tErhWXUy6Uq+hIJMpZp
9fn4TP17WPeUfB31g9R1krtqQrpnQxUkZPl6xAOYzeEqAU7UcF9SSQzSy/jzZdYr
mb2qzu4UtkABFpLOCJ+ps+cnR/FCpEAd8XMjBufr5CkDGZXSZgjEe22eM5Nhhe03
be9aGG3oIfTChjJw5rTHT/IOJkt6tm30QnuwQo1VfyipZPbJUOoZ1qDkcPimI7Xj
lZqHdP+twD8h61Hr0v4+j9/GTOhBQEKAiKFxyf8F+dyZgDLJbCRQDhrdpZ3ux3LS
N33z3QexS8+knq5PlYSiWP727vTIh+NQkAaRPwe8bDkQ0mMgOjbrzVuoTySq0H1S
xaNNH2Y6XUr1QVJVvBIYsF2UkfLBLv7RUB14UkHbqwRPc8sMdM9PeZQR+A0d2L9W
MnTAa3dMaeRbZrJ3P07BdANVhcX2X1aDcC+VC8WReEKjYPYgH4JrRL5yFfEWWMJE
MlcmlfjBkcgqCTkM3UPMMROPeRVdbshxw1Aa/GF0hKaFdINpi5Z4TQFt6YEQz1c9
LIX+ajdmBjPiDLZqLwlF5gbdigy/Ha3h/wIiN3kry8jCy4Dv1W1n6Fv50mXJkEah
QFHEggnAIUIFi/Wdhb/u47xfXseUs9/JiliWoURJyZIIKqGz1REhxICMVESGFo0S
xmHV5s52eJE5zfNdrtfu7y1tdtKJrOONmWDMBYrD9QLfQjBgkjSbG/kRiSq9FFQD
gdcCD+/Oh8MXCaqZ1agXutUFN/I9oOJAcQJ5ZzFPVVPrUdWfU/AuN4LISgokjtwB
V8UrauEXlMAGW++Pq4m3wDKCIbyjSRe116Gi3gF+j9z4VdRRtRdhCJxWpROx8y++
UtYlZChrfgm0EJ5aPYb9vEzBZxkaZcy6IwXv6DNLeCXKgiZAcgWJS16N2WWkXbK2
LEvugggRu9t6KuRZjypfwrgAATanwpUgq5GW7V5nrCu7DjT5o/MtHtgeoIeVPHrI
D1lk6txLM91sjbpXBaNLWI2w8BVupWJq0qJ0uZSI07JyQIB/M/yaQ//A6J03AU7G
N9rtt2byezyQ0vimMdVQwlRs3RNfOHEbIFRY2MGxEHK1NYTGA/YnuNS6d7V4K59z
+DVc9rWVQCkNYBBFxb5Luliju0ErrnbX/fWOCwR7mqppubU4Cc0HWIrhyk1TzKAy
F+f7JIBN667DygGMaYnckpGkjdBe4s+gFhV12r5RqYlz6yQRUWDiWVMmfNE1hq7w
sbqiLl56qw6uXX4kATaZ0q1MNXIcuTTuulFSebMMKA3Jc6rY3PUjTsJCq9lWnVpS
3ph5aJtF6HzsCB4r1N+KiVhD6CFnvEOCh+V3uzeS3tGk+Vwnx66RF8QTiDiUt2AB
fjtvECMuIDiImi9kVnSTWHiNKOiTBz/v61ge9TTlOMwt6TcJ9hJJK3Kp2YX9JSoa
1RM/vqjOMSapfMDpKRt4QJ848xla4F+cHWGsKSgcDL/uV82RecrTaV8MSygRHryS
vFjE0Jqkg6yj5F2mqtWkVi7wwpJiBO5Lpq/TfINlmqXz77+bcvjvlSIWf0ubWCO1
2GyKkxnTsQtGyWxywyibOpJA/CSkrthCUcFapZjGgFM0NqdduHzeHhGkMrAnoBR1
ecEQsvBIEO4QPBf+Tx0zHm6xl87d06IrELclg2mkwlPjiMmJAsQxl8nUFw4oRxg1
l5bJNDyJdXlpCbf6tEgH3u92v2JbKdr6lNN4Xz04F+BCSimyT8z54VQQ/1Q6AMpv
7zUbHiQVF2rBYjvrwbM3InDYGRkR6QIKJgijB5GnAArbddvCc2ksS18xQp56KVMj
9mZraxBtUJOG1VcQC9lzjQhwwfD/aa7B3G6gRf7u/tsDhLY90YBY36LpacqltmZA
e8w5eEba+tdvssvh5Cl/o/uTZ+BApMbjwAOiYR5O3AqTXhmYvF9kXrbtk5mtWCL3
PjZYlHyfMLtwcAr1DRqyhC5SiFxW/VlLEVwjt92uy00rDvji5PR0sKvuN3JzGU9W
pHVBp2q/InheEHfhu6dznpbre4LgDuq0pf/GIJCNzDS6VEJw8tkV8acmU17prBtp
Yusoae3vNMb2d8g2q9UEhla5frr0VrqpsX7J1mqTZojPtXROpevDmnqn5B7/5pYW
WDkwtDF2Kqq+4nR5wyh5eyquL6CsJtxHfY3w7QdzTe75Y/dNUXpq816OA4hgHMO1
8BaP0d48BN/6Qn7jTL9+OOPDmvEBvB1FO2Ey+2f1XM4VmAsxAja7b3Dn+LYxsRPS
MKopEMyWXRyfs/gCSOVYF3dqrH+r121A0J0i/3JxarVu9gj/5E2yrV9oJELBRmDi
YtxZt6G/2OnGFZRTdZCx77g8c/k2Ut/7XvZksaHs23hzXEvi+aPUQhL7YCmJsUiz
hwkrHU3+EnPHUvwbzfmPO+eFNtAvQ86YzhGYyqqRReibh/unuSccSpOAoKIpzpIv
bqhToN8XrpKmREJ5ptUwud5f/nm09nP9587HeQjAiTIcGXxCO7FHIY3NoSoLSHpU
/aRiMnTD5OpOeeTHReBEnAMrrwLjIgCkNWM+ug5x64HfKq5eFy5kG4zQsILKmZFH
NE5LsfbyiVcd9E2gSyl415i8Jo+kNqiufpw4W+8sWh0GUn4vTcpX1aiVLvqK0yqO
VRjStDKJJNavHGVTISWLPZ5w516P0jv3msZ5AumEjIJNctdD2A1IKm9hjmLPUgYA
Dak5jsfywyOgZS0no0rMnNL5eYgXmVnPuG43eFr9BEqpJJxBe9HDnq6iN0pAEt7x
qiFfe+eAp7XJmp2WaGwBygwlDXDbqj04y7p1XaVmF7MKBAG/FeYzkkzQ3MZ1pRrN
SgQ199grnZmOIGFEjjhl6z85zzmlCkU2hJBW1AtL0SElURl7xwheYTmVTzTL5wUd
uRIkA+9HI/tiTvEgGWfPoBHxel1t1h1PQ5U1rnTllau/SWuxOKQ4NMjpff19Rnzj
XquPkSJvtoIOA1VhU8siOPbMYS9cre2U8RV7txMw7CQ5gYMeJG11owm0ryYjydVS
IsZF1vzPNLDlBTTz1EBcZCjUCu1cu90RVBhq9p0MKmfbMXGkuUl0YnwtdNVD+KiI
b8qUu6S5XDjcbHPXBko7rE8dbNhgJyuVqVu8IEop1wD0VO4vIAdDKLJEfANdNKDY
Haoryp+57qmtSimkxKloEi2UhQRb0pzY6dfeiWUBgifVqZ7ruWnYxBgbOWLrWdvv
7PdJr8b+tV8U4QoFtqyJYpCYjb9tnWPOr4L9G9avVJtoekvbEWynbb7GIVOPEzcZ
yyXTEp5jCLKj+IzQrtaLGJK1e0AFIgFaGS2knHrGEbTh45y+QO3UURnh+V/N0eIK
6ghPSg0falS7Y/Irk8JA6C9fUOxeKlXLCgHTH8cZxsRgwY/sXZqmWRLo6P9Zy3W6
w/CFETqruze2oJLOswy3n3W/vlACe8lS1Jw0MZ4Qt4oNx+0xYHUZTrG4yRbPMGkP
nw0xqxTer8iY/NjvY/ni4MPsmEi5nt0sOulduM1epyoyqwzcbLPLUCBb/n1ZnHbc
nH2x7RuEo1OmST8K4KGSN5Dx3zbe9DfckxJENoPyqz1pAvmq/0PkgNsQv1CQZnJY
WCHeoNDPsyAWfz9ijVHgBNgzRZWSmZOMzg02DJH3cdtsNAYI76muDDDoRDPUKmAK
RfxLyiG521urufSZgeBC23tsaxoEQDJINXk0kcs9+g6ZzkTZe6t7gkzX6+yXHkGL
gUOSBkBvYvDjA21pV6ICzbDBAYPjBfli14KghnOwz7juWrTO3o1cPwsbnt8umOha
AzdzvDZ0I8x1KYKdk2gqq8jcQxivPIWXWhtp4X4hyAEQSe0lG6ZF3mW5Vu1c6R7w
6Xd4IH6EEn85gJLfvpuZi0FcuBbUCcazpc/tQRnGLwkDp3wuRf6lizxiXMEXRTKo
inpfm6GGyhwfQuTjhs+flKM5ALUuEwzG/7/CGIwAnAWYujJKM6Lk6RdcIm1HpOzZ
DztBs3dof3R4LNT8SgS1fJqhQBwb5YIPShcHBAQSdlIhm5Kw0kAIkRtWkTukBtM3
Jp1QwmDlzJw8b4muEgho5tUC5i6UJhZFOT3RsBFP8tiM+h0UnSquN0jE1fdab+w5
qY39/0J3s41JY+CyutVUxlzV6yvCElaylU36R0P2aaJDMXNgor2IMaAb13rswVm1
cZcZtRU+jy5UymQfyZKePeZKFRZrZapWH+6W4383gw59t7ln64kgKZxckZY55JnG
ItO8xYYW5vpsVC2SVVqE73krNvUNwTJnElXiGVdhPccqfnAkg9lpbgsxjWA9hmJY
gSg6UNXay83I7kPmsz8xJNjTUaNEGcx08n4eIbDgkyA0gCKzMsvghZTS5cPRS34m
EMRqF7qqyaGVuv3vtY/LTAsAxlWxtufXPGAuFH8MBje7KshDsD0nJ+iegQtmX1wg
NdnUIYmB1jybthqgeVIKdT8pt+28vrbrcB0rGRRTZH53e1nHfz1M1eI50wN+DOc7
4oAOeT24jcnmYanqK+UkDhIlhLjGRoi2CDyUYm1Nw4KUaY+TzZJzrs66fufhSHzk
k4so0eJITJDIMBZzXcKR77T+0Drc+hpKHlkQhkx0i5hqWgm+bGzq4nD6g+/rrM+E
UdtqSIjHBlC5nw5UKyLF0YUmtImJiXANqpZaAi+oPL84H91oWkF4LAsKwII2HhZV
eZLYOUZ7EAS+gw4vQkxquSNLxyTxGgEHyQeJsfLmzzAJz4w309Hc/5TShTuErfkR
BrlZ2IdK6LdRg6+CF2ZYPDI5/frfpKy8DugAHh2Dc492nQydsQY8M/3m5A51B+gv
oedme2nbjQWThsMx3QIh6Bnw8pAyLXjIQF49jmZ9W8DjpIu3ybKmexN8LkZba1y9
xpngrrMF2EH9B167Bj1OVK4MqekYj8SPu793n/MJTUDA40CnQPKn9XS1Xe4upyty
5kHnFG8BKMZ6HDFW9uw+PyOEZ6SW8pTjHfKMZw0SzX/Jm9zsSD/DUp1F5i5WAGZj
j+9nJQQTcYj8U0+DD+N+Q0yECFWF/wIr7v8QLpzvUYzUHFI/lB1MGh6t2nFq4Dt/
PeFoPZioJ1OMy0pAlHeIwGQSL/iyJvXfT7u9wy1w2UaneNW0n17gDNoRvSFJzErR
pMLfXg8tv7J4YY3H1m9ZBLDBIs+DbP820LSKFDwGxaI0oU3SF6KaV8D45O6l8PdI
rhcLJrbRSNlvP8n7B+ICF/UmV9Z+E4H9Rx4hmhklOg7cyG8AbJW0Kvxs2wtK62TE
vGkorXbib4QJq8wx3FRENZWxgowQ5YYegRozeK4Q4bKxkyeqcEs1Ge6MQutv9L8H
RKDo56rLspZNXls7RcvsTFclkwNTUfajOXffkZ7yX4GcMFIaDxOQ7E6xwdbmt/fT
ylFbvGyUQqHnW4z6KF345RYxakouBO2pq6dB1I2JmvjBvj7CvmkmEKM78wraM6wf
gTE6VF+1+5Q/AHkJPgJX5GagklDwCtyQJIq7mVeF25J1bbw9+k1LyJUbUFP3r5+g
gG4i2oky4ulVbCtqvUUXdKMX2/wFGy1Yp+/39pF2kYb+zCTblRxEOqOvlfgA8lAY
iQJefvQL1ieNP88nPhfcXitxg3g+nSMpxfJr0XVoTJKpm9hCa6VKZH7A/dLiVRiZ
ieT3TGh5QiGV/Kwt5KSyST9wi+EAiu7QR6lm0p19LHbZmiPRd9FHw79FdzhlAAsR
uGIH+fhuCF62KvnwtOsV9b8xlu1VJhsQfV9+APwY5LGfrpGlUjlu3o/DfrgZS82R
myUAu5kcmEH4EKjZxFCgZ8fUZdTfLknCxRunhRN1fiQtD0cFxp+KUwdGFC7kPqmg
3Vjy3S13A80gVKR6LGwOFHlVbQbKe00XwsypcKaqLylDAVSRDw44qqDfVbalwsrk
QNeHfMUFIEG+5UjIOt5WsvRqT/xkBHLFuV+OW16G8VHV4SCxmYHkiwLVLAfHbPNX
Om+Y4Aj2kjiagrTVQxTCkFnGvVkmH3KGN+QzUY4sir1gS7+XJE8yH1vY/GzOyL3P
BSPtHf/GBckdSN5w6S25jDRtGcNITE7Zkv4GKVOL0WoIM0hy2rayOZGengPFMlMm
rW0WIHx8bIgV38PfXU5r6vlZUh1B8u/XbwsoKqgOINCexTzVTHlUQChtANubN9Yr
4MjQIYTFS2VtaGdpmwJrAgRbDNEcsG35JOPZueHtPqfrPTRvz1un17KU0DuLBONl
r+2kPdMpUIC9vbeT2EimEK2H7n9Lix6c8H7gZYFAPmA9MVJRjNuR+GLPmGlJ6EB5
As0hJONZqXL3NIiZl/LCMJHuL6olrlwjRVRMFfIHbhmS00sXLFgwCVGdirTt6gc2
Sai6XL1ZSqW8KO9Q7JJv1cboaGVjwaWt7wE77T2M8T6f3BaPk3z0YT3W9KyvFSLx
fvV06ZzCyU5W26uJCKOBIAMZyJ1W/TH5uIpDCNML71Xq0AfYNN7BoI7USsE55HzD
9MeNmptT4rpoNr/VS1pV+Apg6iLTxk9UhBN7FBdmC8Rgo+UHmvTtBkBn7T3L//jt
8hwwuYcjUfSnLMt1+cFXQA4G6lW/SaWk3CNlUd50Fp2Xz1k4hrNV/jGc3O47l3SI
hvV5dlIkzgiACFqHWhwqjy/2hXhqDGB5eIAZUq+a0+yQMvb3Cjyl0IVQNWimKkLc
sVxZns0NyPSyZiDzufPNT7/xBcaPZg6xQOtbfY5UPVw6IXBxU+4CDT1W+t+/qatr
DQ11xDfWN5SJsME9LjB7o4+zgPMgg4RrTRgEaJP9XQuIrjLI79RiTAZME/LRL4h6
733nyjq6NDpuy9LV0A7l1HLykRQsVwEna3l9qBxa5epVegfBkktzJNfJ/XsS5sOj
ChkfvPNxDLpFpCm3DKGiglprvuxyYcgh8wO3IIT5n4FV9bsXM5QLQGWDT0eKLv22
XCFRz8+Za4PF9/t9obUn9X5lHJwua8mUzwXRYzEisE53pVGFE6kC//3G/3Y5OQUN
+u+t5H2B6a/7QIxPdaiFLE140UsFUmpBCCDMnv03Px7n6aHxcjwCBeIdxzl4fcl+
nKVj3893AXlnS5AaCYNgtUXUnXL6Tj1+KylzVOR8cDWIODZjzOgCi2e8i0zBihfm
3FrVqtU7nF+TMhupgkWwFVeluCqty9hdEj8UUZu/Q3Bq/qSYa+H+MUERyjJV20yR
/gGgdyUbAqhJ1jppb2AnksgaQd1asyIUNMVFELfJWGEgql2D/mT91z1jLr03AQ83
RgMfmgvF8I3Bm6+JWTGzBN2o9/eWVa2xzUaCIS76zboX3T6N089zn/blc4PLUTxP
G9e3n6qNG2MazEzOqi2nn4hPAbCu3nfRd9SvQoiqaytzDkcdeE8iVH52bKnZ4A5e
2RZeOxutEG8hAiGa6olnGEpbWL1xhMZokiZpWdLO1BGOPp/pEse57+PeNQBiLnJJ
e/TUJM1MvIWshXffSB0fwr27sedKe7XPYkKWpMLMbKtr+XTFWvdRI0fLMSrib76n
+/7bPzinYZd9Lb2bWOLOB8mvlsJLVoFXWBkUt1mEjudtSUVaHU57cEwWKOFLcB9r
aaiKsRBdhmyEDY/Y3qu+QqtWsZC9eN+k/nSSFuqW8gFO8j9HyDAddzs8RNbTJm8K
4iBcpGJoF0935RWxnK9K3uZvzImhQZTJwur28Q6wjqb3QrMBQo8NJrZojdaH4aBa
w9GkqRHaGy9VQ4uk3ItwZrtomcEyz8nXMCVrOGTXvuw5nqClLXwCQsdDl9THdIdl
fRMT/UmkZggr40XqVqTPDhH1FMRv4RNcBoIh2xLLYeYHJ1YNxpEiNPFbSntjWzsm
wRWD/+qdyKwdT06o+RFypGSLN/DWELmneBoNBb0drM5Ff2dLJT+FV7zwaVcR0wLN
UMhwIel/MP+9z6IvB32Hd7n8Ju1388mFDbnnhE5M2UI+wu/w3MMJon9zQzuYIwNr
DExnqxUviCdKEPeR0ZnbeY+vfWlQkiPKuQI1YB6kkrHUHyGu4fAM8uiC38HqOqmx
wQ2+zbJwRPxiDBNO0NM+KYVlqg5pAE74eM8z45kSM1sRtcOaJxIfSnpy9jH9GCWf
9/hHqDg2/IgRSYmZDsZG1REEEWSIA/h2bORWc51DpJTAgrvbgothdpb4PUEL6xd3
6ONGI9tS1et6XWs1D/sbFEgN/UHOr/3k1mn2ODRuRR73pCP8JBjykOKOfCF7iNSh
dVrj3G0oUbs1avXhr6ltM1do/2vJmy1ZizcwVueKA2qff3VH4TLvYcWsySMbRmdm
IaEmmZ6aTRScprhbFLOGyrBOEHR7htktNg93OLPSjZdI2kUQCf3L/uEjnVH+Y5YS
wrvXNAFRGi3rY/BJQ7ZQhV6yPClJHxKj8IMzkhPiXKWuYDZ4b+YJsbFP9sZgXOkQ
baizj906tzVrdKgrdjmR8yfQHZH11T7vVVn2PFnCUE5Rvu7UwBZIEmj1sk9cIvby
MyNgQXK02lJyjZhOC7j++5qi+psXCXScLtuzmrZj5xkPMXNIeq9rvGc1rrMUHOak
pe0aqdbAgD29CdaU0nJ3qalQ8ADRYI1QCmRwA4tV+LM6y818Dao9Q3gW3mLClp/U
8SJK7u2GW8f6SIpNmZkIOFUQMQiGudx0EHarYClilz1elrYygyFwYv31fD3A5ySW
B4wJPDhCqz/jTATmD8LQiwTNyLn4BglFx/QdyhaRvxj+uLECHmWCSxFh3vBtBjVg
Z2J/46mb0auAU4HaKFe6DvVgOElCunTj7Gswfi0L0K6y5vKEDYPpYngPmtdf/MVQ
v+zgC+226ArINWXEvUxLX9RDppsY2/ze/hZwPVYOVr956oi2a7lNecv7qeFIXl15
MrFx3xSNO2cvh/ivXrON/rHfkxKJ20hZWGykTWbc51Vhd6VPW70gJOw2gEZRQts6
kU86fPkOcFYWVMI6mfjIF8TSEFGYFszjVIGLDjaNbDwwlJAu4iuDcX4RkNX//h4w
Hqdn+/f0IDAzAQ6+pACQBGRilZnQ9cVGtYtKn8nBzJ6/Stn/hwOAtKQqEma1K22K
epNjDxHjoIEc3cDkZabcBYtwHNI2Df3FHS3/eXGhTFQCzxAh087WgC8gx0lSQWH4
B4Wd5+NCzXxn9zHPTxcqyPOFWxqUUEfNhycofwsfk4zSs+xjR9EZ7oqqEwluUhqN
btjFmnyIt7wtoLELt3ljzZFDKjjQbAblvb+tUczqQfz4DaVpFCISxWK2BTwY1gN2
514AUUrDy4y7PEbqdpc3/RblbE1Y+GvtuB2mVa0S75dW3N5yCV/2d2uA3HQdQWQs
FFtGleOy9tuqBF5wwiIz8sgNpQ7vYJLiHLgz/QtnoWk9rIUOD2GDZmmamMBCxXoQ
8N4zeptosB69aAi6quVKnZt4PxniagTO6joWJFbmX8a+LmTpZgiq19/C8EekWcxd
8w86mdXcoZMKBc1zlQG68k0vJNVhVYZWZrlHBWapPGoY/iTNu6GGv/SiiYUvdPfa
h5K5U6pBSG67AywJpe9tp1Ipi2LjjHFyIHLaNBUsC2iGWejCQZ/T+cRyGuKBCTr7
TCCe06cMoXgYSKj6847wFvpp4N0lCiJsV/YEw+Z52VClF/l1aRwDoxJ9kwWWF6xZ
gWKmiN5A8lRFhq6nPUK9A5x3unLLQ8f5e9LeYZ+1Pjx9VOpH8BicgC1dORHMnwjZ
MlN9vAZ5yAL1C/IusuD7BqxUK4JO3uVh8AQk0WuYgS9rL1zqipBuYG/zHgRzGsCy
W0BJcOxfSrQzgtNYtXnj/7VgG4/ojYrCrH0qvbIwuBFiKn8LlgHDj1BukoqxnoLI
RyvZYE/Zcbkp18o9AswcytKZ9uS2vvqU0jl9ppo9gbhvymXzeOALLHXTB5tsipqL
qctOJ0T8AOThu1PtYzTrsnKOxlc3CVG+aCIxmpezSCW2oFXetEKVfEsFgns+aufn
aI8QWm2YA1mOLZaZaaItXRjpQ72nAXwoWs1mS7I2tMWCeSoldZBWodMy0N0xLLkm
xe/L+BhC+1z4m3d8bpN/PofEXf7ha1u+tInEUggv9riu846eYsTx675p6tba/cXK
ZFLj7JY/MXDlcAhWXvSFW/tILrBaJeNZ8GCU6+k1DXoFNXgOxNHYbvE7LG9dUJKk
tMKy4tVybLe9KzPgLuy7fndo1whuwxJ9fY2ibLb33mZmTLfNqfKtC2KfsdZlBk48
EA4abhuWFFxHxE0tnqcyyrqAq7RGPH4pEk+hXDPuYTtMsO5kE12uJ+u88lQSmnqE
p19RP+1kFOfvPEg6ODapQe+FR70zrHVE7KnDUYewMh2RbCmCXVbigeDzVz/7xq2d
2GJ0pnab/3dhU4322Kmx/EoWeRqEevGPQMt21vKLIfvGQ+660i9BVMFjN5GNEUWk
ABq2TegR0BzOKYyCT8wDsrC3Tx6l++d5A7V1vV5q/NzGq4DeENTbMoy1iWtsCQR9
FuxwW0zirE3TCHIexZZyn17AT2r0fZQSzRJrVYHpI6LH/M9jfjl2zYv6lXgcKFR/
GcT+utCvRUuUGLvdYLDEII+4OW34sdlm9S3eIJg4xav4Eaptq1XlKbTpERRDIXg9
5p7s/RGGYNql//prLBUSk2vUqkVLCSvEZ6U74r1qCTvecMg0GPxPaFxwQkzinQtY
BlXL56fgPaQvtrWQWQuH7aNpyfkZCJ+qAZR2TWpjYvrzKlR0IQEwZMRh6KIjHeg4
UL1aVsTPhO2dV6Y15Xp0D5dKtXzqntRvXQ38ztiUeYWDr7txKBgsAChwJUZEC5bC
7oRQKF+ThTyq1ilZHqeZuOOHhFum9aKQtxJdihQ8doNupM0E/r90D8lVyCMXti0b
SFLuof4WrpsMOfshDGNHXT3azMJGmMPlDZ03mQ99bvRYqqhQYt7n7ZFtfshGCgsy
kpTrtd85ZuEkgdRpYHHz1R80GLBvUWWwV3ZfQyNlIVlaWieFl95qAzYBXoIJZYvC
ZBv6iqwy1EWLCwS6ExdRhhQn8V5q9F5GODRGGGCCZ12uyu1bqGUS8OR+pf4xcf4s
+u/W4FRHyU33IiShNyA543kvjhgGwkGlQXJD9T1TEk1XMzP+dDlHaFzdeVlmbAZu
E9ja7LQAtFEJ5defI6xjeAPclZ2xV5KgkDf1zutdoYGK9sDKGZEwrpfPXipcwMwx
BEzy2lK/rEWNVQe6HJHDdBPWD9oFTyz0TcI/0IzFrt5eAkAKhayoLhI9o6/m4TWx
28wcgT+kied81giewEoD5T8cIguJLPpWpSqu7Nm7CBjAmygjJjINvafoblA3DadC
/vx5DC/F0aE2iDWeUz9rcqv3SsRdUOelmZgTDXZfEPBAYFWE4NcFMvSkzzTKKpa5
ympwNqM1yHrKbADZI04OGf/V1i+sXyEe2/3aAdo46vTMJCQmHxuJV3oKeB7xXd7i
bvZQv4S3BD9Z16LCUHlMfPwoIOUVwGUnWPiETvFMrfO24oEkPwpLv4rBM5/kXrHc
IoFPSU/kWJHDgSJPnONfmbgRkbWxv/98xib0CsxfYZdyPB8hk/P08a/SjjhbvnMC
HB+DYOiPZ7HWsLXl3Q2/2T7D+yN4gtA7+VrBUlsRaP3MAYpJWvB/3UVqVPr3TCOi
idQ6Sn7207AFzNx+di7xZTPb5JH/eus5t6KXpNRqJA9EwaXtXHeodhO8kfq5txMp
vWQ+pYciR/7pg9z4ecKoyZC99xO5+WkLAH5v/Ne+ckKpR1EW5djKDjQMXEMFiDGE
/aknwArdXOUEHeSuh9ZtiBZmtQAvojvmXu9RPVIajZl0Y7myuryoB1kb/M1yvYai
r+MCUnaHeJZr42XDNydJI6/dqYwrtHaR2mepmwzq2xkHcd8qWNYCAB4ie1jSQpJY
Jd4J3x5gz5lLk3+H+zgzjiM0L6Qps032mw4veiy2mLkY9QzKtMG+elQALo89DxIm
zmlpA2YZOrxnX1CavsFNhKRKjYguWWuc5f1l0o8xT0TM+33glgh8oKlbvrWj6wVO
TfSLpTXOuKm+me9EDcsvHXWd8MDP8jmBHoDQ+UPP7XwHumA1/3CMUe/+5apGUwYs
MxebVaqmd2MT9KisD7kJ+C/SOXKOnGS90fzwr/jyi7GSUMQ5RO8yflOjkiyutmFu
Ha+l0DHyohTW7lEeYOt1j3GBWEgd7g9a3e33nUPf4118AZZPlTD6w16LDnOQj6GJ
S31VZ0iPJAyi2Y5DuHcmzkU/vMPshI4Ng+aykRE/dzy92aaqo43PysGhytQlljoO
OloN8g8QMIR6rIFEAei+0eV7BVOqtQH8Kwfh2j1T/DL3I21jq3RWkSapt7BlzGQF
rOBgXqkRBvuqcds1f4Mf+YuEJPFrRc7rXpSoMwHEM9NMnQ9FcBr4Zd/wE0b586u6
lLwjdkp0LQroKzOSwUdfCYBUDYjNBEV78zTMO4cGdokIqTQBaa4b4ggZ+oYRo5Wy
xsTNZ71VL4yy54MGYaYYyHBzx5n+SmvVfEpJvq8dcxi75S1sYLXJUSRzl7+UW+D8
MCAOMPl7qLts3JoLq0Dep0Ajt9WXCMYjretae/9JTY5jiyq2Kik1npWUUoZyyqc+
K0DOkNu+bDdEI3WfJB8a0656A8P9a9qcW6uAC43WNBJJvkJsvucA8PyGHrPiEyGe
yfvCXD5MO9v8cvxwMBzLK/+A0Dyhb1tAXXnfC/dNOxCAYASmiSK2ZfsvYcF7X6bZ
FCyv++I3gW+bj/MpJF/GGk7MRlwEA2pJc1xrUq3jUQsIbhMy2EbkFJ4JkbhL+1LW
IviZeW6R84PpOMTPY09y6SC1gQPMssAKxhpyk3yX6ho9CZ5dWSAESQ11+inO+I+a
1V4BpUwQgItv+ORVSCfEA49cM05wEL3KMzNmR+OohKt+2WLc7/OYCQfuJzIg3rQo
wDNON8OrP127TKAPrxsAQD06RJOlP4A89JMycniIAxEsibfEeo7rV0/UnJdPf3M/
cy600YGVUOUHrQa+aPDmO0cnJRKJgRDWK+jVIzjw9E2nb42hgcXB4ylGCnq2bT7o
JJ+X185mpHAI36ZdN1a3b++fWo1BjyHxPEPCXNtrier9HF0VB6iHLxqG8Q9eewCy
9EdEHoTu3bBSBDwdvNua6iDfO1dEIC8olx5F98iiD4UpixBTy4jveeVUNFoazkQF
wZ1ZpNk2Qo+LFih88JMZN9h8Bw9M0PyEXH9+Bzc2KN6OlbF6GujvOEQut9VobBqI
3FPgmaWDSjlSYjS1Au6vFPaM661lznFGdJb4wp6mJnH92nRDuqAduUGOzRqAW0xB
cLJiDOgi9ihCXpIUNi4oI3vQmihofFzQhSD+NLmyVxQ6rdF3r+YNxIf9fZIq7PdI
IOz34/ugqP1RBLePRn4RKITTiP3z8pkWA1l13kTZKubot3ZJMXjLPMGEaJ9h7kpU
76F7rARZroH/aOdGFXDYkCPhctB7JibFqFPi9QucYOJB3EXfaVzykyzT2vHpYVQE
GYcXCz4T/QtIj8X8GpnHzqghcYlJC6QK0oKMXII6JIA/5u3AF+NljVDFamx9dCo0
tlfq/J/3kvixHzNSiN+pQuS3t/m5P8zCpcUOcU3P/oy3/IfT9UXMwnaMw9MW+5ND
fB8WStLC+B5b2rxCKrPYzmp4nQTe2FL3OwelPCfNjSG6QxUJlLsk02gnRYqZa5hr
00SwdJzwBECze7EA9IgKZv8+bEVgrurNU1/p7imO3RszSoBXRjqMZiY8Hh3QUXG4
gtJPKagYcy8DiiMqmdvCFSDqBtgTRcARGIJUrFIRXDpTJ4wjPUwe/6YJUP+XnauV
7tXiI034VeQSpii6DLRktmjQvoyOUgOgHgH2rocwkQ+hFFq64RYbvpBsynARYYSO
koMP56vHPH9dsGEoeqTi+l2GzOnEAA5ALHHVYPNGncQqnvLu7JGzacYNVo05dyT8
CRzIt+61Spq1LXU+38XtzfHLjcUFSdbdUDwSjm0kESTc/rPbGSZZrLn+yw4nMXRC
CYX+2NvWBB19kJbt11KJYbBYKxAMLpBgFYmuH6KsnoyXduOuPG4Nl3b4atZlBzrF
tUaypEjKZyQJnDBe9AjCH0f0QOjAlr0F9TihbOD9sH3aRn6FZIBoXJdWNd4ueplT
B24513osyWh6sEPrR4Mvd7ntQYWjQOgrcNZL0ikevj9CLGH+QFxOwVo+c/Yj0Gt3
XETco2Jl7rMvWYGplZPsKzxFM8IvA2F5AIgu0MU+xEFUdwWH98MWHeqlFOLWNE76
kRsl70tMgEr9Yi76rsPGBnHdJm+2JhQ4DfjiTB/arQ6zIpcaGiWlosef1Kza2xWS
xTHwBEduA4WT/EW0Vw2E6oZJ0djcO5XOQLLEb5O5aHlJxTwS36rRjtouWCFvP7BV
qgJo/cBtXgRQCiJG/ZgFXjffUgj2vg8OxXf/BSSWnz+cQ1o2DOlsB7RsxrH2k7z5
vbNMKO16shNx6dCjSdjG67SHUY+t1Qw1jWdM8igP68yaqebm45LzKjD0Fs3kK6JK
ejmu4s4koJ9QPk6TfoNL4xL0btInfkfQcU6cmpg4OE+CnFsxccDiebEELKsVGR/E
ydGcSrmqnpPJhDxTnI37iaSSr3v/WIC+nAbX/p+5Ooi3sQmyX1UwF4KNqvRmhLak
pyEsVWgCAFhIx41BzoHYhtgDL/I4dwSXBE5wCX5nocED4dPgJZbePXWL7oZjrhf4
8ZynPzCKkbhkA0C6sCB2lPDHGytexKN8b30VLeB2/LPxDgyo64Y1qWm19GfvcdbT
1meKZl9Le3yRgDe5iVcNQEYBUmssxwnLudlJAtmApp8gEXSFjy3c662l66ZSOFsJ
ZNXNb0iUENyKIhT0q+m/mrI+b6YyI5kEYgsB7qJthjOCYS3iUfL8WTvTRe/WhpLr
17eYJoixA+iqLWGlNVW9XF2tgHTOtXB07CA7UzXPvcoHJcmKRRiPa9hN5p4w0pSh
odhUaPpYrwRTwbVFY34xq6MGpG2ZAWkXLfJCuqqXaAMyYwyMMPLeE4SZ9iCc2cKt
VyTLkXaa4LseBYTq9WVWbm83pJBILOKt39ggMdiTkRgniGPKYOEohAqchMNR+ExT
0bg44tf65DmXGOb3vOZgA3hopBrjdmnccnzvzq1tioQyz3X9BquD6C21el1cUB8F
ypOuz5oBza8jeZxOOmWmqeLslbQu4U0qwP0Z4ZPh88IJIZbJWJv8c70If7emRH72
ZMV7+rh5h7PWam895cGWX0xY7LNh7ZceBJ1fXmu5h0eMfY9o22G9bjgEXvT0Z9zY
nMsbsD+MI6fxYlewDuSeVHqoGZmI+TTvYkFwBXev0ZE0o4aZfWfJ8W+wCG2FRiof
gsSoCOXwEeW4FdIMKSc7BLxrO4fPu4SnPdGFyMX60CBsx7ifgOSUdPA7xQfWzqVe
jd0aWrK0wJrHYstVuoLz0xOS8RhlumCdXSDiO1irtwBMJM1im7UepVZDO+1x9mRX
2KfcvP4H23ee/9MVNX0TF1J2oIABpIqwKI7hnno0FMShZWc3aedOGxqY+0bSzXeP
DtY5h8Gt1pGzY6IwvtnBRTHvLv19wPuEAH96hIhEsxyz6feRE75gInR8nB135ySa
/nvbBfXypR6ieldnSCuUlvZvouRBWYUOhIDjNiSm/ILPMm7NkKfGM26VbeXCmTQN
nPcZB/4a4F6vhIfViUrwiTChBEOckIB7mIEhseCA2v5IKmfgdikb4ySAcoZfx3Lm
Rr2uyKqWvO8AVFHnS2KxNNT+BI+3kj+q6cHSgg8QOhe6AJ4kTgBS/wUqxAtiPyGj
Q3e0fLyTmWVQ+6zlBHuYOS7LTmQLtzzvhqQwkWSNEapLqPNPbIJME0CPWCiSvqt6
UUDVus7qSEVEaIcsqKV8mmh45XFPSEbQ/ag5ANLDUIjbzxrsPr6W6W2y/4ST0LVS
LZDtZL27F13+DB/y8GKofc0NNcicsrkd1mbwaA9dizyOiB/fKNn38g/g6miCFJ9F
Obl8shWYttK+o/i3xTA64gI1cvzM7cgP41cSWuCSwo0sk35r/VkThJ/P6WZgumTV
a9D1I5cb4AWZoYXASB/6JhY6X7gMQ7tMRa3znIy0vZOOArZ9SejAMriEO0diE34A
IOYWNfbOMe32GHhFyfOMB56M7qfA+dCgFMKCq43ATdCqAGdgmc/l1bJXDlioeSTv
Slnge4MZRUtPOck8xy3t6mVlI/eox7mI2/+xNWR8rKI73vZN2GJhRIEBaLs7I1FI
lNgjbQbeqfsL1RjBtvvEwMhmrNbxboXRZC/pj11FyfNniA3kpFluSufkBMgX5sqz
tqZohMBa1Ddb1BGT+3bLGp6tuC7gjt91fO8x5NbseKf+1QpK8ZrYcS8SDz1zdxQq
50wiT532XymlfWnTImTrt5ZGuKCC1gLmWM4JOPIARlrtwjo+eLnU6EtDFDktvySK
QPCtadSd88bvceUYssroFaURbslPD9O3btTy7swcNCQeBt+jGRENk5N/Nabk1jTd
8BZoQaK8u77RAnP3LoOTfGgZ0ZTW6jOz7fNTUCFi0/T4/fled2geKlD9iCVFGk6l
pbaXepjoQwS55RiURNhg94c0fr3pjDZsJXWrb7lQcflmVl95u3/VEC2qtWx/PNoy
ElRhrpdtlToxlspP8DPqvN2AJxd6NXZj+kumY8QqTSD0YWxg3ywsFCzjin+u6jaO
9eMqtNMJZR3JelYAGsjY8/4fY3gXOi5Kqb9ffdpixckOqHQaxLWbYXAYC2LslHXJ
e8gXtUwRSgQ9QlqyyXhaKEapo2pZWD2HzQCgc3wR63kY67lRKNEyzfII5n+KLZVV
s/b8crmrsOM8nvHOCqEgIJ3j5I9KNq4byYHS6wZbNS0WkOyhf08woostqaNwS6Ur
pzXMtmEJF8gDAN7H9QNbBrNe9f4WjkdWymHAxWj1349E3NCU8h9r90oYqZ5HVnue
+kUuN8olKZy3ow7C1HLZOYZb53FNwV/yStJCTp8L5qv7YlmuZAZoOw+ETQKiOE0f
tm9R0zdyLeJXOLsKThFX4U1rPRcVw8/HtoiQpqWLuI85VAw5nUi5UvAMjtIKF2lz
0uput998UizvJdb+Buc9b/kvqqHUFX0aQ+c+VrlvEbt+kw2erGWmE8Btbt1IW7tO
O2NqXFsjdU1RMmCOdL2CaeWx6LNWPcZwGCrvTvL2D7ccnhzX+Vz6e/UVOc4mY94e
X6BOekABMpeLJ5rLPdfdnSKa3x1q7hXToHmaj617hrrFJYviSysNSt40yG+HrujF
YIPW13ERCsK5fv0E7mvBndrIhmbSGQDAh6Tdi+zQv50+yiR9UwTdHJ3l9oWJWd+f
UgOAa/xOhp6nHiRWhUGalbj5lID8XiLT3MOQbp0MdNtzJASWEVXxeFBh5CqSmjP5
Jc6Jd3rpRCHiMmcrWul2i2Nbd34hW2myrOgtekREbyImDULb6duOSdXB7aHAhSYj
CDpydMyDI/gIkum4eIhBlS5hat1JRk4S+lbvSqfbV1RWMwEE+cp4597SpCF6YzCP
dPtAhlPcJOWlrArfPASugNQihwAsiXHy/bKCTedFY7Q7dArwsVj0sTVOneM6cfe1
5qGtPTNIikppHuDGpbMP+A/4GRxLNn6pslzEKK5kiO3NC8BocFtZ3gpdMPv21jWo
+BBc97JpyszeQSdBWz6G3xl8qN6AS73lDXKXqRvMgNaZMeUbUWsdvOx6Kc1169rl
nSvMhYXtKRhiOkO4ovwpv5RdG8ok6Vbh1z21kOgRb5T+W8fnC59sd8hnDTr6f3xV
yya57oUlmxy+Hb7l3Of/hafTKweJADtDfzr42afpGSh9ZKfyLe4YjGYs4rfF+8yP
2+UROQR4DSA1FDLAkNE1JJIxPKsKmtmqer+6FOoB3sH7cXM/IGq7CD/t93DQBr8T
U9+AHen56SGdTf0wVPCFmR3JGVufIIAk2l6aaExByjt0IZs7aX/6fgN4Pw15lbxI
zAJ9zG6XFU+hzjsszVf4jwXrQaX/yZKybtogOADLOAzitAbvhdg6+o+7l9dAY212
QlISnA5VpTZhrwzafg46Ej7sy8AqpyWkPupeW9mLX1aOk2M5QVf3RhclMOf2rxG2
bPnrcQM9rtrezPIA0zjo3AhkTKqsrODTNiSQAMShENywBesoMMVcY91V+km9FxGB
r+aA75TmQcIm3lmXXqpqyFWnHZ0RV5H6TBPSkB6/yI01uXqjNLOd/fE0pVjg8XrI
FRfX5g8Ju8GJa6CXsdgCJXdlFaGNnTFBS1066K+upIAYhVYswskgEknOJ9e9Pc4h
cWR3S/d+aLpApnY8MYmmefi6pozeTd13yOHIKUTEfkOzmC0ArKFxtoVafVG25B52
wUtX/NNY32HZIUcwSI9FsW3BGw/v+WuypMag/tXYM8OalrVhUpozubmfMO6o5pmC
3LT3dObWhmmnbKZb1EiWI7W1NqZNrzJP2ZAenVtbhuPEE/1USi5dPj64n2QlVJWQ
hpd4eA8ZhDXWB/IH0XKk3IqFGU1V93Hb71GHg3OdxJL6pEfHvElWZoWBN0MHsbyi
i1gXqkOLXPiF62xaZpnYx3Xbr7Jg360qGCYB8qBPjVt7lug4YstEE5P2E3Ho4sW4
u4Nu/UcVijQLMDRtd+GjtDuNnYeas4sOA6xMcE8BTgbOqblhpEM1KpP3yNYdWKLk
qdlXR4De3Glm5y7Hw9CJbFcx9bmFwLwm/ax9H7aaU4a6TR7coE1gWcroGGP3QJ7u
fez/AiKiCY0SfwI7eWkszXpW99HBScFhOMHFIHtWirc99GcE/pCvAJW/uzovTkk+
U6lyarlYFGyf8aUJVhlyYtEL+oi1o1wCNzj58+gonclb+B5uiW1nt2t7WNapIXus
XYI2nV3h9Ms6IbmoNZcGunR4BF1vdpxmVSl1RTdgbHjUSbp2ICub2uzoVtNbeiDs
itBpVSzCKuhWVuoW8DJPDd6YssIT5pZyxwKRc0an7wPl+9LpKrX3X2/MVsTQjzaz
cdAcd+TcZviaP9Ll7k7ZaRpoWWRvSKPyhbJ6vEzmCyyHg4KYpnoMeUwmEK70Cbsk
DOQ7ZmB+8/qHjL1odu8aYncq0Y0qGbrikZTtug3616z1xA6DSwXQe1ISSKKbU1C+
mE4T4XQFIy8i1W1vaiuzWwUxZf8ddSX3sWv8Jk5CIkLI1wYoAJF2ElgOpIbrPoPV
4HuC5PwCuwany7277XEWr8qAlJ/H963wIDT9U+YiOqWO12Egk+Ujv7VcRLL+GGaj
f3uC7m7kh+tBz6K3eS1vB8m3DG7g6GAUlSBb8C3U4A7QCMH2BlaXETiHsqQTfqOh
J40/HL3uaq4pFmSfmkqkTXkZmpTkLUIFJtphJI03WaqcFot1Q2yDKo4b79rslwAK
2v+TY+BV/Jf0rbMFm7v5l0TgcZOjU/Ra4/OMsCj5cORsDghwbrgTwrZklds966Mx
gU13m86CJNZMPNOruxpBgalJkb4/GE6/DTlWjfdy1XLPf2c2Bj5m4zo1Okt/XBEp
1uK1n67oWJ8xaggqDHkgYmGLOtFIvbxzSCOSj+NItQ56eDZh9ghk+A604PTYEwyG
4rifjPrfLxiZZ2kx59XeAIuU03GzGq2qFIcoy6+RusjdH9VpR0e4X3PE+ewwyT09
sn1b9t6jcUdmAoNhAKEh1QPm/3bGjbmdxi/D7Knz+Iiain8WhFv6z/WXYVLbyZF2
T2+7t0AnSOW6IqOGxFy+68ieTz0Cw7X4EmcoEyj2NI9siVvm8CODjvaAqQjAcKTb
hr4/9XhWwM35r/ExdnWW4HIRncyeSpkXI6nLrzKWvVSx31GTOMqkBG8RcOEX8yrm
UEoleYd5ZzzUq5ZN1AYp/pdshvgXliwR+xMNJVk0fH7hzOyR12opyK8NNvq7f5ZZ
Ng6z5Dy0JidOQ0GxePXFNwFO6aS7kmNxFqgET/S6xt6SDQ3gRhB3dEmoA591F30w
85eWua5cmhALIq8mCMICktj+Qk0T9qm+Z8fjRiewiRGtdP2UHWeBf9mL7o7Lj0Yf
4FAnmiXwW2/WBuBrV0c5mZAqBggqhvg8fXXzM59uLwQYGSdSgiL/bClgj/0ovk5g
OqBinpOAwZz20P3Z6oD7iX2zsNo5Jz9XSbq0lU2QKFvanBodGFY1G2yzvhCE8FWn
mFlxlr+xSq47E0Hn8HMjxapX+NMhd+toWljO7KLmAQEA9yLsMA22vQNdiyt8vcSo
v7lnFngMbyLNqz2JgIfAnT5HC1+xMNtnwlUFwo5zJqWc2bT6qXTmGvEtjJAv+4mD
uAhv6z+HRpGbH8oAOTrF4LKwMJfw2Bl71N4qAr3SY43lUfmHqZ5Zx4QZSvbFkstp
n+UbknTyVLhX6fn1atRAIpWLYJmsyd0vEc6pon71gmniIwH0qk165j4hmXS+YHvw
YlD2i6U/mrPeBlC2I0zAkSdgeN9d9cqYQCEQ0ZvGJO/LJBsMmI/zYcXWjod7z47V
paGaDMnvFPjljxE+R+qR3S+Q9aiLLQ1VORKQOhBLiyEWXdOsKEuCzrMW8Zycusgp
OvZwXiLxZdurMeP6JSeLoO+5fNGhSs48Bq8lMY6E61KwqmREi03MRXR0nnPszpOQ
sdcje5DIodsUD3BkuwXO81qUgsCuKYifD/wFe28aW0XvmgtoYxPQpeimnHMxscy3
J1xeI2v47wQJPFTdhg8hoM/ZHNUlHKH34BUC2JImyB9O2DpmgNb60qPzgdtLXm3Z
PNzzqAykWS3Q1rkM36ngWilIjv92EPAc6bP3XZacRpFh4DoakbMQ1+J7McJqUQZs
/q3TEgqMj87dVf9HtWFRBnLjtbWdFpXxl9ZVTdLt3bj2UYZWj8EtgkHGcMWBMClT
fZZuioKFLeX9Yw+ec22Lv9iOLDL9r07t5EhoICwO2hgs2O1JK7yRtbeTcDr5+Du4
NEPH/FBe2ts38Bns96ngb+8FGaQJBbuMIpu9uksP5VPWUB7Tvef1vhveTICY5iTm
ovWzuloprpMYwVAXSX133GcZ8BWnRBcRUime9DvTIT6jsJhoaUiMtW1M4LSabmHh
DVlP+SuDmGhAMx8IFCZjOMVcKr/ouf5RI6qwDYw2n2DAeZkj/ZPLY9tpwyCr8CHr
RdrdItzyEHwSCJT82Nphm3fsL/8SmY+PGduYpDi1qsIuqWk01vedZOGRr1FUhfnc
6O4kkzv8C9sIIvVfXHjzZ8P3cHIPAH/bvC5GBVAg6YXpjOf6Ne9FW34W6k8X54Mt
7CVJP4KEWVY/uz6sLa/Kyhx00DYI0/LK1pJ7Ac3+JbdsDX0nDsoR8Y9Nq02QRHyP
NQSogcIgg9+Nuv04PoxcjQPNqPYQo5Oq8pDbsIkrtiiJvFbp5XHu0DRRoyy/cbva
TyRGM7d0Z4+aZuoEgjCvcGtGucoFYw5jEnwDznX2iRjF1KuPqQ8SCDlNLy6q/Qeh
spjQdT11IGI8ihZGA1n4WXD/ozSf3Wy7pGdGx4/pbtfuKIVUJKLG256M8MP+dYqO
mLFKunbYB+2PI5obZGYBOmkYQ5t0rFoePbNGSyGc7H00Jpop6m9oBwIKlhiBfdFs
bzAdmgMmSojkPFX+V8eUZDXdoeA+IQkSjAgPTX55q+J0fz8tjI24yQ0EoKhmJYOZ
6KgOX1rM6oV6snLmirnlhkvX3b/hKHDC2oshHhnKjLFZ3J993s9+OU6/lktxnh7j
sJvWb8XYNq/KxT1JLTZgb7mdMRHNu8iUV0bwoaD96+2KHzYEtBt/d55O9+LmbDD0
ViCL1qYqqK2rYv3iMxwoyKF8I79Y3gaVcgnSCgoCSxzf8deFWRNzHHec69IjNdf2
QlX76bLQqvac2vglWvDAjfpONaSRrPcLYDIsGlI+7okvdDCnzjVZHHxgnhnoTQC8
8gsRezsXX8DLFxAEJoLn/hTUOg+0Yi3Ou8AHwHcZjPbY9QuY16UKtoV1yF6FL8j7
fsnS+Dp81ICPsO4uwfkDW2G7dLCjexygFJqs3pM0mr0gc3Oy2fypw8wvNa15N5Fx
oPX7N2tJooNspOn+cJQmHziaaontf18FcNJXculuPxpwZF8jxPajcclw6elMmVpm
87U8A+952E1YR1VZGQcFdmW/Iw5dY427VHL66r8TcEc0DHYhTeAb1ogiMrFqHC3E
bGfihagqQqZhkxXmrwjupA/MNdKc8zmKjGwA4ccTskLLocppJtVrezwIkFu5EFVc
CJSGcO3eUVIVRDlpVhSxEp9FGvyndENEUY1EqFk/GWW6oGdqbc0KPWKZEzQrXndu
5ky98XG5ZywhNrIS2ynyQ+5x4Dtp1lT1XXClRdKKaX9a+aVlMC+1Ut0rjIUrHYVR
FMYdoWLLO6mPRWq0pqEA0MvMQOdqgnpodCFN8rITERn+lg78W0XOQf+3bJZSU8Nh
9wCHsc7ETpcwmLdmy72QZC7KyB8HUCtyp9DJ4yhx10B6ASGJdz2JwKe/idakxf1X
GNj7u7s32xIu6M08L67S95HX+h10kvLYwIEjHMHXLY6ZBRkFgK5i4QBjBoD0b5aa
5GE0dFLKU7HBjPmChoxa8w9SRkBcJu3t6+MEWKna/k6wQ55Uo1Txhy/1N+UsTx60
Qu9p3JLhsKXZorD7g1z8iVF9iM2ObetFeOFrxCPeSOe0CVov0cUbX61/Kg7G1Cup
ZZWX3yNbwJAESfjYg7g0NbOB09j5uuPHJE8f3kfNQpvcDoR7bdYBg0ZjtapUqLwF
sWDIlH3MuVlHaV/TmnOH7L2+Kx9+41qq4sk03mhF/BYdiet/GZ4+4+BWU5Upp9dB
ef350B/aRpC5ln5TZW9ugvtiD4ILxb+YSbAmeF1fkWMQ9+K/tsreOQqbna6GU7pN
aBpHKRK9nTN/jVmLmS4AVTO8br1yZpZqwErQYOIv7wKNSadt91E2teTQmpkKYunH
slD2FuLmO3lusesU04x2m72zKttrL6VuC5JRIMcKjwT72KCA2AyKpardV2rRriKU
xBe27d/T19s1GwchudrPO5TvmCu9va9TQ04XalSBM2uisVQY+SuEiK1m9Y+l38gK
4aDaPId/o4vLSPly+f5ajaEObi0XP7CoJqRZNpu5jB4MvBhukANg7uRwk8QmYy0h
tx4ejAdtWJ2JV9k00E0p3A31ZfQrzwhBZvl040DyKvfKXW7iLWllAnEARofnIYLk
5brz8BKjvmH7znCPTR/4e5GgsYzNklsnBGFSZ7reIatFTYg5kgI3Lr621IV2r/FE
1dSOyLOQKq7if+9Nr4qOQRti9dtFBiWk4CpX8VElbF7eqpcOEUO5UJa71TA9MEQI
JhaWBqiZJL1Wpjj38bmhKJc3mbBhlKaED4t4NZRUdjjGrtisKcrfaKOFgU1OMi29
rjus6tstzGnTYVMS6ptBdZGeoZRRBwDoLnxQglvHLWmjQ3YP97YxscV94F7qTBmn
eZbBjbbRegKqjkUNDFQ7oDYsGKBiRBAH0Xq3vAppvTL0w/t4xBQDiXz2ssUWtKPn
uHTnMjmAcpdEERDT6anY3/gh4CUu3v/6In1t0optKM6rVsBfynEH28rPdbm9tpjU
jucmiXdv2GFpdYJoizOBL2KuApph5nWcoA58dh+wZTTIogAkpTaVYV8eFBHARfux
5I9C7CYEGU0OuMOEYe0W84eC82L6ZZGkB1dJ+Iw0kgVcakHG2qChZGAqWSCJOACz
3wt5Wqmg3SAD+ptK0cI+3Cje5L9N5GDhqV7KYCqsfocvactaSxmiU1YFFtIpNxnM
Vcb18xt4rij+FzUsBOK9sLiSQDFUF+PLC1EG5pj7k24Ltcs1KFUyqV3e1grhdHhs
H7JYUnGONLS8Nqn4dzVpkSr91PaUtMkymj5FZIaL6SwtFWHoEmGm5S4mgIJ/m55/
NtbBuzt2iWOqXCXk2Y844dniLfEaP4F6QNNCv2Y5LJzbpdHyegQ5JJQVkXqjFyiU
5w45lC+qkh4beLqBU5n/+/KOtmncLSckKAzA8RSn5cJDW1CVPwGZLa3svN5E8jS9
vh8XbBr0W4l/55Y2yoHk87ZgtPxjlEvs4av4zjNEShvSkf6j0iIUOeDJiXcI+lix
6AGE70ZhJujgVm5ZzDAp0zbCthsTpZFuNNIKdRMeFmvzuMZZJVaKa1eVUb2x/rHE
+nd4nbBomnu+IASbp7UHjURvYTeUkqTlIIkRkT3Kcr/0Ou+O7E26dBB7Jex4tleb
2sn9rDJdWhPB8UebbwhajFYfJoy3lgUp2KY39uvQ+E14ARZ+MvLok+n782I/9W7U
G6vtjdmxhRVTC/cHPr4L488vbXMhMpyrwzL+LuUEuwnSVP4+KHBAOdaB6QXxQrgY
X3qD0qMFQkkC9fNEiwvAEU/ToU2yUX2rIM/+hlcy0v1ltkVWkvMSbbEFBAhxhq6G
HI2wzN5TDUlfGajl6mQ7ilbUnzD3lJH4BNp3TZIXQzt0uVOi2BdR09OHMEIe1mMg
n6fj5g5DwF/XOy6MpFTCS7tfobmOV+rlFchvslZiA2xHIMHQ33xzJkf4NF0LvfDS
7yioWjb3AdFelH9EN4Un+uZp48uas7W6zb4flmCYOskUquZp1MIgm36YckenODMd
7aR5o9ZojoeSfr0xdbZFC/MR1ROMGS8tl+VGkUmyEInvYWo59DTCAxbKSPOirDrX
inMb5l1knjS9FeZcwrhjOZZem6wopV0cxpNVcI0tARJSiU0LPuOAHIqmRgGE6jUE
CdLsdIHpl29bgWWxjkpS/2qphO/WRydCjy7U9rabNy2/FHP4Hsr2NYZVVhfv1nF6
Hhk1i/WdIORPyumQb5jwZsBqJRlagsLgi8haA9Xp0sI+rhL34lMqqb7dUvM/zTK/
vMMQEZhScUrZfEKl2qQelpPXip9Y/0dvYOJabuMfbgyrDqhgElWpzFcWvZ7AmMIH
rNMbgFET2aUevUWj2qPg8UtNFmHnErHpROSJDTwSdf4X+0aXaTEaHT724SwrTOdT
kchnh897F5o96wseMJUdPX11X7z9UchUtUDqklwC4BKO0eD4m4U/+myKRqJcLh64
1itsPSXigNq29TNLgiQbaUkjpSnKoEvkUPnuAhD5rsslej0yoaS3pcEm5YyQPYUu
KyswVj1+ekcKL40MTliTTDuCdVap5cLQtwJG8DhfNGDOm/l7cYCDeHvBZ2r/p6J1
s4uN4PofE/P84aKvjfHQxL11FpHdUJUvXfJGnNcgjoQXqx/xVA8m5TzvNcR64fyf
7SonA+mglZj22uCkCdzx/IGJD/6igKlLYAme8MNCf8rxHQgPzBahkWPvqAz+/dJ2
Uoze6FmXiUsgnsXnO/7jyfB0Aas0egb3FxEt+wT/2WRxnHpNZCvWAxGmgHgPcVUo
4ksDE1Qj/1hj7i1fLM1Db/36wVMHs+yUYIqi3wudV9L/RDR16YJKgzFv0l20XElt
e2aomg/v+1+xCbvkw3RIbXqy8fD4BbxMrbji3JWEKZu8jqKj+x9k9hEj+1T2Ujen
J5pg2gNHNga9eRNFK70DMdqyq2cqvoZ/hSFtLtsy7U+GgO9pC0nfrOJhyg3IqE0M
eXb+mu1tLgBgYMzAKP2RYZaiUHSFGqRDczG/7wunPG285xYvnG+jAiiLJCI+RAcM
O7TUmSYddQhChMEzU9MTDgwcqNU6bC94dfGofJCkGYdrKrRig5pVTUzkgmjiM3wj
6hOli1HL1nHW9zbDbu/8U3Pg8QnBHxpEvxHD5ZIrExjhQow1wwiWptC5eC06hlsN
otupN1hJBDGf/353mhMyOzmBCRbgJazZX5HXalWWCLndFcJ3i7O1UKt8fQ0YmMll
dAZbgwJdf/b7ciGwhZBzWh+iL/dJQTKSHBXvSdKVEEGwP50hwCI7JMVz6tKnfRR0
OD5uy4ew94WoPjVuMD67+6Iq3VrEJxNGU26ii9yJDC3CXs4hVRSqJJVScvXEN4XL
Sf50auWvYMlQ7oibiRxAVeJ5vzE/S7FgH3tICoNeEpM1dKBxBl7YsTos/2dQ0jCl
VjNBaLIecDD12UGURyLBw1cVta4Mq0sw2Pvx4aF0DCeSkILmZw9t9AwV0g0C7cO4
Ta+Jxr3JtwjiQUKl8GiyNyIqER73XoVgIXB27oYvFv2Jmci5QDLV6SMUGYjm76f+
E40NduGXfoz/spAoIuAkT0akFX6d5mfD8WN5DOBxTyA7VEhm7WWs3T7wMB5AACq/
RQu2Un7UrfZSSQrQOIzJgVrHZNqx/hRgQDFbmixXYmgSC+jXyG2FbUZD+5kKYYfi
jJnaAyDGAmN7jeHPf54/OPzCSH8VxiOTikR/VeAFWqzrK9PmPFIkstudHSwQNe52
XYMHyCYv741WHbMgKcM2v9kWta/sx3pZhnsswv/4MZ57zjaHKyo62VeFIHUdqG8r
3wFNLPsGgMEvu2YpxiaPpDAA2XKAmUHmqVuWw7EF+2cvvyQ68559DjQ/LOBH39wX
g8xXUENfUBbErq/LJUX2uHwOYU6himD+Hkd2LoDAv3TO9KgRIy1a61OMLZjrZyxc
8tepFMedZzpgjYT/zXGXsbaWPU9jILg02eTFVvPrJ4tR/hw1FgLsHaSB4PMhxt09
LXwQa174z8VENXZTkac2d+eTqB/AHVgOM9IdIganDwA4ou6d/R0vXRce0x+QQoyP
jDHIzbMecFKt5ug52yBNU2wmLKAvUdewbFKx5zM7oZ5LnFPHgx3uCzfcqq7PPxeJ
/GW6P5/4N9R76I//kdX0qOkyBraeSEeme1LlR0oAcokZfMKNUd01cVvcIOMw5t/Y
Osj7CWPY6/IHnzw3qV0iDsxzujzuQ3Q4o1BwbvO/eXWGBY2BlO0seuZIdNKctkww
F6XxGcC9yHGEeI+ahVjOzDUVCkA9ziKej64xtNV4/of+N2NssN9LqqKumyL5n+HB
237ZBAOFRL7tVOvmNfcgcbxcFGRu8a9rGOsHu5AbO0CsuIPd6hYLf53qww4YbYXU
+pM0HIa96ou7uvyL3qTHPR2O3FfU6VZJnETL0FbTZw+vvGbEYTXCDPUsNzyh+I8G
EbWEZXw7HRxVc6hTvgguT9+OTmR+sXo0gAinnJ0wtT2XfY//Go2Z6FhqAifTWl+d
eHIaBZquFdas+INrqldXhP9Asc+uVNGTyzVB41W+tsRoXG8eDwfdectjlyw58ds5
C+Gnw/J8p8jSidusKORi4PpVb2nc4U3ECUL5rMhQ9jcYe4rADjSS0FauAcnauzx7
kV23ORuzW6N+1cYmdnx+mSQlvj5x1bM4OX+LejhPzRqelZEDeBECmyLCnFq5lyAv
0bt3Zrok+tDEazhV2GiZsXUf6fLFEXGerd+gDXCA0kNHWHNceLCy8/zGAi03Cjtz
YqRSCF3opnHwRnYvNftk774tfYJOXJcv8LgC+KGELlcYAJNORvK3cShRjGMH+7aK
m7ZdiJyZjw6wPwp43isyrSv9rsivyg3QGzQqQADGQZAXzBc4J7uFw7XvDPv4gl2a
z01QOSyGqs4AztuUQD95THjb7H0S1vv8LYuba3aJSY+5yoQgprovacguEjKYRzLI
8cQoiER580bCIoXKDLLRqlLuFn9a0CJEyUBp64PYNitrAO2p7PNKi1fbDSs73bir
y316pinuuHy9BSjDT+BJMPaiJC01BE/r5P2LDygPtIb6GkX7UMeAldcvEMuf4Iqn
TN6Lyus7CjbVQIUPHinXiu0ywUvE3/s74cM8U6Dzf7id+oi108/QTDNFMV5qw1LI
xyWLHNVuHBIZdhtVsI9sA5CpLL2+6uh5PwolWrHqr0FhntPdPuhG2GfUKBD4v143
p5Gn0hcpNU+0oRekRo/ohA0JOWanhhhL5FFuzDt2kHC7I+kptEuZeLDI/ntb8kU7
UeoVLBQ9zeSgXi1vJgaAjZDB0aRtwr9PduRatTSJSECaTFPC+isYmaHJi1GebJyx
J2wb3DqGeB7p9esv3iPjMvEVaUtZldZLJNwZ61ihidiMlpB5OvZ6JBngz8eGCeDn
LtjAMMvyvU0FPRHdZ8Kg3nOYelqIXHWX9nfXy7nZt39vuyY88fNdU51Pdrgms7PP
cPz0GgtGFg6T8h1cFZIiGrPTONICtqNSrzKAHI3IprkkTeYI5UfyLMXARolEtqa6
llwycPQ7UUr4yvYcMu46sHijszhStbERO5FUeDl2ntKEcAPxYWZo+h874g5TRpl2
Ki+7AmX4AXWGHLihuw+NafrVJqibgFOzS24URpUi3L9hw8XGD8Lok0FxpqLnLOtJ
zQzQkzBaLkfdm5K4dj3RihP0p8RbdPcreXLBjK9xdbzLTIDT14TSbeODxNQFRJss
EbswhO+kSuOS+7+LAyy356pNR6QN5oPGY66KBQT0FHb6d9UIQoZAcBcL/iFNhunm
Ck58pGJYS+QkzRWc5kBSeLsaV+4gdlCbO/+vcqAoTQo2bQLrfCTGyOe2d8yLZJ6m
Xt8iO+0tMdS9hW2+b9MvbdvozxWsg2Vt5ZYM3XogUVUHArjwUbLK0GSALkh2rCBV
Z8msLo1q3wBt7HyqYxDz1E5FQJOPwfIIM9UPtOxo4Q/wmUcYg0yBiRE+LKBXBCZf
edUb7/PrmK9jMkwnwJjltLnYccQJth8CwYK2GzQJyVMEOV8ZwZPOXoi2rwipf9ZS
3dz0655G9LI3SSfHVckaaJcwqgs/OYAp0CKNZTNuQXVHAujdxymgIe1ILeOlpXn8
VVLDxrwPjLuMbUN5S8bIEF6Rx4gY/l9B1uAixcxgHL9szNEprhqoHTX4qEiGa8Bc
DxCYrU7eoxRWQhVHDjXTA4s/P6umLCbNpwmy5/InKDuZWqetEHayK/stUXvsk5pY
LIIofpPyytHZUZKuJ07I/gewXccQ2X0ioWWsU0DgnlatlZnaprAdWutNYUiJ89A1
db8m9y6O+1s3GJpJBM9DfiTaB5T0WWSmPY+gx6gorl+y/ZCrZMohEpUCUSAPhzNI
qAAEJ3IL6xkA+7mehhL2vEaLlZEceZoMArilkGHXoCq/mlyxf2AZvn0/ZkefU9Kw
/z9atg1TvdfIjUCHwgdiCOuKQ5k0dOReey3PdXhAP8nty40/JX4KWXxp8iE0NFFQ
BireRcwBrKiQqpE2bbO7JeJQkJmBmnO65n+JYjlco3HAKbtHbFUfYYsmTyNVP2g2
XfbzsWZo4TFbBLQ77mMJpj2wEvbchz3GGbG0HoOxyTfGm51YFODtkx2naMI1JAgJ
Ld1KNB2w4MmpiOba6OQ0bvqAumAWygHrMgFS01O1rcN8shcavn0KCRMcsh4+UsTB
TYYecVmY0pAsLeU7QtjMJvizBpJv+BqH7QICaikgzjGvREXuNwi4CPY5hOtRjbp3
BGVzxJxUcx8wM2ZLNJn1Rkd0zXjL/FHrzlSt4K2pV1BUS5gYEuaaj2/qsPjxUxFJ
B8FGHiY2RRHwdX0gfWThFHyMx5O1O8m7T1tmDusHjw65mCmmgKEdJwA6Z4x61Ila
i53dmvHZoowXOt3soKdlJb2Hyz5dnP5c2oKT0DcTmjH/oNkvRnPxrNlIoote6BRc
VzBbNRo1UR7K4qyQskXbCl35YjhIGvedOkuhZKynX1HEo0fPwTh7UPkWZBBKUQCF
+E9lZAsCE3JjdVsYPLYo+y7Emr5uYLN+Fg2rcCdiuULASnhBUlu0k7TjlxBfMYis
RKh7YJ26YzTUpBwjs9fuZxR0sSP4LRz9uI+1DVpuPbm/CI+1ViPj6luv/MTOSFPN
sgtq31GOSFmrWVqSRe+7IQC7U/CZ3ffcLWdD6+LdAaeyMfut3xJy6+bOepkofV6J
UiLf4bboAvrocNUTZssreVWVHtRjGRZoTcMU9lvHXzhqUAjOGqnkhgTdELKZhbqr
Co5Mv0dz5GAnwoTGoqssYf4NKkGiJ0UU9GYolF/qTANcbdUB1RD/PYx3fuluU3R6
TapbWE1eXPhxKHw4AJM3jLHHNjXObAFqO67c6p0CmKsBqIxRUqweoZXAfPD7T1o3
ZBhowv3ZkJXyPk6SWPI1tTV2NgoIs26ep5ZCM617QzgXzqriFx+R5SSrR120whhe
fiECyjoYN/fHSEEMnAmX18QZdUcB37lAkvMHfI9Y9PYVmeO4ePey9kFnV45mYlXr
NodopVBNA+QSZ9jBVdWyXJE6xgd/7pWb0RhLcfexvl8l6EsbsbjowYm5DWDvafMq
jF0N2mHxw7OA/WDeYtFlvJVMJI0fo/ZMGNUcKp3Ne8Y56d3B4lAifMkK++sJ2bgE
mql/9Ot5Ffi103HiXRjQxonD//Uy/k80fFU4aJMmiHsLN6tHAa+Z8sYxvKOjPIuF
YAJm+wbWC7i3jdMmz306d3DL5C/YqbOD8BQUhtYuf1Y8yJEcBObdFXRznKSN7a4y
ONBVDb5v2ZWLJzYBipYrGVUL+8lxtg0W7GgZc79TYHCwcX2L/gHDvSnAKRW3uzz+
ylzmxABbn/N/kBpOAEA6jmAd7M0LqgZM6o72UD6WNof3+w32++eBUb0hhXkKJrrt
SuavFPYzcMDPbWB+2XhRfPuzUXQm8k/K8i7vWeLcD7R7F/33fMsiQmpLIIXnEnrX
tepCOo9MDA7fZDz+KsoLEDeMXEQg3NsP/JYA+83yMQxAUFGJPlT+3808iqDXXYuu
3nb90RTl6HUJtddV1JCUabbYzHzTpxItH19p5rNuA6m4SuAiuNfMokLFpzSiYye9
DMvESyaRqBvcttCt8gRHRrbztHGy/1x1vvQ/JeJ6e0KoWPPa0hKu62xLUYwtO4CG
4IiM55GPNKOZyzWHjQxX7UMZqESDLORs8SoZ84tVwGsA1E0Hj0xMU3bFVB2SEa1n
7LiB1vbm6ZoqUP+/Pt7RO5jTnsvYNFxjLo5sWWs8+9oW356DlBkgEapUPGWGdZTg
ggha1newo0npCVgk4d5L9MMGyildirBz3g2USab+uSBSZI2WCMuJWONSY3XW+XHb
wvrRXzFNK03S3WfGf4Tg9JsJ2fcMQjbP0QQadNsYDFzogs6XR5MxqOwaP5oA39Z0
+gC+mdfPugeDNJcpWrW2MfcXg4djtm2zPjIGfTLPGpCYOO/6FVRAOLeTvxm5hyqf
7ivrhYB4qSPfHfXjumFDPJsGn/XEtqtUnjmREr+JJur9a9EWS195bwQnxs+3b9e6
4V8Xb06TNF2Av90b3MCOFong8aU6fssX3eK5ck2qtAOcue4S20ivSb2ikrD5Mia0
7iyBBBg66tctWHuwVNXMwamt1Ub+gGQoAlSMLgN4mtVvbMCTnjOBLkmUVXl0sGOW
N9MUHBnLPunHErgjkXRBj/OS4Qb9GQ/3ON6cNzbliWcm8szKRMOq67CoqbByuAmH
iWwgwt3olTls5rwTl62EvnszA55qHletLD2Q1t0/iDqMY9RODZHu+nEjNcrhRJDv
NP14lgK9c6zduq04lGuujv5YPA58T8Wngn9N6KFKABOhqAo8Fc/SllooGuGFFr5F
6ZyiAMLLukU8b/1MjCV/Blt/mvR9msJATakXJyX9zqMH2bGkNPa9ZbWo6+pe4DEq
h4/kgvwrFPI2vCiTiuKUwgP55p6QGWxWo0iFXep01Z0n0YWFDr3pWmS682TkRhjJ
N7IFrAnpxcdOUEZ+LadtUOXMdlXc5mZERdgbUbr4IA8PUAqH4PtITmwxOsPQFiZf
uGjUsr1vjKuJt07hSvLHB2VwWBEKf9uHy0quVNU2DqDdQQCmqJCqVtjB/hKfgNcZ
Ac9PaHKiya4GbCqic1wjcrmMime7FHviDwt8IFPXcKs6C2LeXjc0IkrMG4IQPcAH
Mophmp1QUdr2kwgw+BerVnQE5wj2XBTthDmmpWGt6JrhsAUCplauFywdFPiZTnuR
pt15AN4mfGyDpqVXMiGrTjc+wp547fnFGBV9E/OMDZvpCn9qKwyoWEsWLn29wUnO
TIj0DK44bsHsxx8QSRbVrVcjz5EDNTPpSawXdJLLotmbDAEQSG9KuG/hRZlw2igf
KbkGEOJbFEGqdelDBAhnnqsmVOyg29HVfHH1MtXMVewD0HfKqZ/49yckll6NtF4z
ndoogz11X8ANdaNhqeQn9kFyLq9TuJtu5UTEs//bzXjyaCD6GatOty+Ypa/zazs6
ZgWw6nfLXtQcmQz/ONP8BPB8IK617T+lOu9pUkoYIqH8n6Mby1Nag3rZdtle3468
Cny4QsWyUgRfkZM5QXZHvV/+pBlnWdCJp6riXHBrVMpMQJqxDu+k3InR5TK47788
+UEhXwjrOvKKa39tHaDGL/TyCXg8hUmVVY7owES+aNOwqbvghMo8V0TJ3CVhsrIw
MxSVG5PwbD2yaHFl0fpA+cNEq9/+gVemEZj5D0GnPPyqS8ege2KcgUzbk/91DVRU
A7YwgGkBin11epjyhxrNeK3Ii5AKm8nfv64viKBz1IMJlKmVruxRfnE3oN0wAvOI
6kJ3WnWYpa/LmFgA39axFda7P9LHDB5lFgfOYP27aSNXsWkhYTLYMrcQ2UKJ0XPk
NSC0SuPAnhDO/GetWULJdSV6cBJMu1WpKlxdWgkltxe+DHnTh+ffkKaPfrazJAIh
TgG0bfuxcg0P6C8mrGi4WNybNz+wYfBeGw44qBK7ezgS/l7RPM3GWSVI/zbXbOj3
iMTLT6W++Br8tCNWKT4l31B63R72KbvmXQMpP5jwZJzwiO9Q579CwWIrGwL1Ih81
+hUEuYeMIZPtDvtZyogjlIBHTwlKHEyOUSE/LDdsco0GblIcc6uUg4H3t7Gcrv2N
tzAG97FzvDVCwbNu2fA2m1XGv8TGp2HF+Qxp10xn2dcoBrbS5pCTw2rYAWpiD0T6
ZOIdAgKLubrbIuma2eKEjGm4O46WXQ3wmfdrhmpszcnHNbzBPUwClUuz07ouv2x9
OWCvGDpKt7tm3JrYTLkTXJr3YrniJUBCzNUTUBajDb7MwH5JMlyAVNPOChlTnMxV
51iVcxthtvAWfUUCSHaA6WPLlcKb7dTdigtPn+Zxq7M/ke4L6sjnX2RH4RAZCkJq
O9xtatk7T+L2uVQfeXRgckUXTDJ3X3gEYDMeMucajoXSCucz2wmPi8FQm3KmRR38
2nNdKJvPGWYAyPKf/8VXExTGW2a4lCfcX7/NQ7+3z7mhwF/L3JRc1JDh/mdqrXaH
+4hlmKiuFFKRfhTz6AJ/ASmREsv37z067/vI1MinM7Y26909ESH2wzKIvaH2X1fR
WOebdE5geHZFz6ktFExZNX9lXFmGODDXbt2WFaK65CYhUq9knVNSaDyWwvXDD7CK
BwAoFacUMqzwCZ3mylyyRplzewQvVjHTyLp/V3Waun125v7T5DVdaSsfRRdrMPHi
pI5O4P0RxmpMvNnhZNZ4Vya+nWWkOQM7ePRdba6QyfqbaADFZXFZAzTKhIGPzK8V
gOp1bzqQ7NFzyWb4BQbbgfpfb30xU9ydajkujqENDP5FkwagcWbGjlEKSYDdORba
hm5/8GyC1RycBavF2PEXQizSXy1aCuezSI1eAGKeF5bo5U+BssFKuHkNqO2U3brW
At/G9lGP8o22HnGYzYbA1BUw8lflQqh5d9N+WIDg2o4i1a4LjB8qpdtgcMrpoSpf
mTK7qVK7m4fFqDwIqRgAxvvgu0Isa3zUz+6wsjPnhk/1gkWtrdR+mYRgdqDCQZMD
qkbDj4zhgltwhXceKKcTN3dLVmFb4UHyijDe/2aJoLEn4CoFptkcHFYcH9BT7KiA
2ugBkyu7vhoFQAlZxcmwsY9lzDA7PM/cnyU3lszUaCibnOe2lAeowMWsI5EHLoTT
KMQK2LLPd2eJ7W3mUkAxou/xnAdN25dsqceMD6ZvmJ/D1bH3EcRxPezk0xJTC19F
3P/OPVxPqC/YitFjiDGDJq7VQ7oJG5F28clj4j4E4vj6vaAsvQ23VRm7sL3mFWkO
UeGDwirx0S9h3VrkcNzMGaXHaW/Bg1NB91zfX+VdKdus+90n3pByvbylACDlqSSG
bDxn2klDKSvTQ1DDHGmqeWr6OFJcLJPdHPlOGmd6ee8JEHmICIdtJEotc4HuvdNB
LDZtLrcU8HfcU2ApeancwrCYoD71yJvr+35vmm55gh0ccf27aX5XxE+rWHv9KnFw
IEHJDfgHVmeILZ2Bqa/dNs1oY2v3k3iA5D3HsIH2tp5wU5/BAjfjI6aapJ/wyids
gjRtXVxFPOf/tKV+9wqCcKpxnwCC5WZcmeKASFtkWhMrRJhO/MlGh9YcT2sc7X10
DUFehF+03RT7cNtpIIal/mTm5tnaL5H5HKYnS9FimcwZmRe4133sebat26cG8mto
Yw5GWVSU8xO6IjzbjBnRl9Xb5B8fKJhyQSZFVvO9mmR/PLtOfhLn9OrYYhRHvXY8
hCq3TAaq/9po/MjTnLOzqTJuFdZXkF81aWiHxACi8jchjh2Hu8BiF7iwbj/coGiO
luycmDK0ftT0AVcht62UtHcb+WTgsWHv92oraYGrtYmln72on1GKQ2vH6LI2TTAl
g5RqtdMyv/37P4Rc5jkhs7QHBvT4SiWyz1YJuDGATlAuDOy5fDrf/kG+MvT2Zb+h
bJmren3+zlc0PjJLp1+1/lw2+JHY6k0+qpA8ezM5G678EZP+akx2xQsoY1+qwVAr
zyEWpOQ/cJE5BWDq7uRyoYzo6yWiHMj9+KCyLV5mKPZgL2fHNYotSOhtcqVp6PAG
1+2AV9v2sAx0KQ14zXyQ8s9nmi69nShgwCDkM0MbURe40iHdeB+GX0KaFkyqUt8v
a16PlOZxHXpZjUfIqUKAbkMxoP64BQ6HV8tCI++J/5I/292GcVyiwH+W4+cmkYDO
fxxvd9cydMZaXF9RSD781MfDcbr9UUQnqU7hTZv66QNgbkKDpMAtW7UWjHLycYWA
0E0LNj0Nipy2aT5pqT0i8IM4MDyMw8BIW3Ma9qMyncoPr9riOZR8xYYcBCfBj6UZ
3ZBBakKyyc9SKHDecy3kXcxNFm5I2oYBRBvo6h8JxcO/Bf5bITBLXONTszq3vMie
KBANYWVesnStsMRMaGs8Qq7QPa9Mcmm8T5kCap8mg3Wh+/O/O52nLwCCwuu6hKpn
boND6dZoAOJqdJGqaYANbm9cUD60Nf0dXNuVQ0Pc7msD+W3F4scDfyMNToVxAavs
zNQQory+ndeV+3K4R2yzQx2hy6D8qt1t/4cCLEJ5Ag/1Mnrbjwt7cbZgVw8aa7Dj
zcMCYakx2fGu2n9gl/V83PdqBCz6p0Qd8dDKeDy4K/KRdrLQiZRA6HGx4FMvM0mR
6B1/tdxgHoAlxc03w9vRta3kGrOoJu5iGk+YSNZTbt0e7XATnv0/Y2Pmmjquz2DN
3c+3JDfsUGL57xAoPysZ6QxWONod94zkKJDvHNVy0BaDZLE/ft91ewvpLfON4Mx4
yde1rDoarIQhJIeuA8gyIh+i0b6en+p3iYUQotiBelfQOJhFLypAb48JQjTx/+JS
rbALP6vBhQomWvpVKhao/FGrcosg+hFy8Xup8dlTFpHQMoD0CRbaYx4EmO+INGkU
w29TG67kJ6PwLghyoQBgjnh2T6ciqbc09e4FAdElqABsUbJOnZY02hR9aIfx59Zo
dmDKRStvYIIpV1IG6wkHmv9K+Iqr9fQngNpUI8prB2b7qegsEAnBANmFYR9qrWDQ
XSJGyL/0FKvocN3bpqb+fJ77QUZFgKbMnyi/qGY5USBtaJcBw1amNMLByd7sT/4p
thiZebrzt2JzRLXruyXmA5eG/3MU5AVnN+AEGhd4DedfbdBdG7VClsuLwX+rC9h4
x9zNSNK9AVUfAjXc2z2z1HomZoLW82cz0iwysGtKMn4ELwRvbwEGZvTY8gZlBHDO
OX37Dmvf+7Br9ECVnWFqU0tt6xtN3CXOSUf9iJMi3bltyzAm0pJwJ6BiPKUh+vTS
2FIi6REK5Mdbje1y/yxSy/U2jUiKd+DjAh2eoYDkmXuJ3BKMQUjnf5eLY4U0Pj6c
0DIbFl7eKG1YUebzUSxr0pqGOCfTE+rrLBhRP6U4hdz+UlLfaPWEinz7JyjCFEOs
qzE4KkFwr1Zwy0orcalQsr3YFyjbvFulZbhZUDtlNsceGuzaM/Zgle24q9Ed3qbN
lFkcKB4xKZ5cI8SyCTt+d9vriM0nT7MKp+Tk6IL1fStm2vKQcwhMDfUXkBw+pwRP
3kpZgRRaMd5b35INBovSjs3ZvG+S/+Bca8DEFEvU0jj/gw7leKUlSNJCficXnQz2
GdeCVgxC7sdYQbt+SqaCodhqj/cibQMFcWukuKl1/DOZu4TCM3ptI5f9RR2W/+by
SeswEWzTsCsjSPXQ/4zIZ4ssNkqPB2HW6SMKxyHcBVKnElx+zLNjVYvQD5Sr2vtU
lEbDh5lYIdL7ig7n+qrQ5ZKJ9l2gYAlXW0muh+wVquuW5OIiZjGNOYiGQcEd30LN
ylXVHageIKiXclkpQXC12H/2HseEuYQd33LuV8sLZBuEQzsQTsise4eXI8W6U1Fu
UEQNCo/YsuDFdI5/FGdn//WHIxUfTjoNrf75v0RVsBo5a1MmVvsLmdPdDv2ufNFC
I/LJWjqtgLdFdd9FQq0oaB61ejucVlNvU25BRjXdJqKzbN1PCmyZGDoUkiEMLf8a
EhBmdqwGRc9uA8wLO35bEI/tx2yfz0n22jxuPA0XuWZje1XKd9x56SjDBLHWXB56
V+dQAPzJHhUEmLwdEBxLt+PQnvq2q/2bmejH073VjfZB7DOzPQSUE+JgEASOQYyJ
PoWjohp7V5Se+3j29BCIX5ZSkXqNh6f4pdZuFkrEw8ppG6wz7V5+yrPBYWLIm/OB
xkp/jJC56aBjYCHUQdgYbPxlC1bNoMUAK+mC17fETsENMxQLGLONx6eS+toj334w
Nu+YjzK5WNggV9/tMmME09ghSLEOCTM+5olfsL13oJVJWToHSsufTb4oNV/Nh05M
QuEl575XufaTqOCSmK5B9zYr1kQgiwZdyAoKmIaOJCMgghmtPosYhocFsgsIUX7N
FBkhkw1q+9ooQNyujkJy8rIw/GB5qx2hxuvRkjh32aITZsynoYJ5brTiNLs6fyO7
kB8d1wpjl4kHvDbb6ElumTHeNpkFte4L9yrzqt/6H7QJ8opdKs7+y5ggpXtZq1v7
samdxzEwprP4UXqTsMozAY1IQlYdUh25H7nvwXz3l/q+xpKO1UtRxpIlNk+l726W
XZtqn1OL2M/rJa0qNKUFFOsolZxtgRR7mJx82ofYCaWl2P23O06zJWtCga5coZCp
qaUvNlAYOLf2qPqzfBgcLHnDbbd+5eYiYO4/IbYd5otPwZGF+Mlk/mjVg5FujkHN
2jxa3Krvb4nsMlGsZ8hXYWkxFjQ5VANOlymmmMy6VJmu58JRd3IF5XoNCqNgz8t8
TQyxcmxL0/UPpMuCCbBldgYYx8b8+6Q2jBR2i/zhaaaeuxMX5cHjpwDxCS4a/v+3
KFfkqVIQM7naSykzLNxHCcMKnWECXTrOa/0O8zJsQHgD54XJKEers5zOtaqAt2uD
irYBSQZNgqpruooeR1BsT5a08q6UknlqnX2Sgm4qaeESY1dSvXniDBe7OmGlwd3R
br1tCxofWWF6N/HxZN/AIIu3HsVo/ZSSumWGfUf7QXehRoLb6SDJq2O1xvFkIEmt
ozgmhbspjqZs9p9/nyi1Gvx5r4EP5EsFvGyWBBiLh2ltiBQzamQoIXhBFKH1Vc6L
NHiWByFENCv5O4P7IEd6/Zb6DF+tRKH+2j0rlERUQZf05iLWA72NB7aGxV5be+yh
tgwx0eqTtt8wnS91pEFBR2KXlu8RQv3cRnhHkIQKKlpjwex+GLmq0G36DJSTAZxV
HwM7PbLczjGsdgGerj23WeeIAisZtdpKzdL9pxg4gxto9Se1KMOrwpfWsiofIgV0
9wjK6GfXYj2695qnXGw56ku8/IxSM082GOfoo4Lh1T7LeMGlJ/+8rhVT2tuJDIIS
dDzL4lQyEhdyKo6iEH+coenUnbPrw2T+B+sxQV4BvIhAbpMVuoh6ynvt8mQ86PeO
78qOi+ycfyQugY32aUv3e2PGVwQZgM+wfYprwzdWPVAZIMp1LmGtfCOlozZcOoFa
E4PDRwuaYFlZZZvQAQv7cfHp4h6rDhWjhus88cPV2GkRyqKAgk457ImL1UdNS2f1
riiqe2CeB3uiXtvDNzpXBjrB94AkraeQbmDoPkKJC/jhClFImmRKE/iswxolfxum
tQMqUsjDiGP6ydf5QiQXFzEmahvaRS9aFHHkkkb0iDt4uGhCFmlG50U7O/V4l4MW
4MMhb3ZFpNkpPHqGJAXiqr61Owmp4ksVM0LBN0KF3HLrRknCJWQ5tOpm57rwAoKv
wiL3Qdakfftmuh8ERTYrzIu7GccUu5IK6I1YhseS62TpkuPLHu9aEMabcuHdpo9n
ywEH/jRYEijFQ4MRMshuz0/EVxOkUWACzQnnkZLjKt85kTjf/zU4QX6bXeW5iA57
JFpkadz+ZxPVXAu8PZ3B8jsxtscShAw6duMwE3aHaASioME+idh6tPj65ClSuJJu
w8Fv4hITCD1gzgpZ8WCIaJ0dp1xz2Qm9mZ2sNyc8gdf7zNExx3OJIIDS/Tpz314g
XNn8myLjkBl+5qFDCaTp47Eu3FpkwP8ABWfLPJ1W/GRixbkAX0Jh9oK4o5RkfTG1
zZAIXJjkO0ZjvDjr2akpo+FTX4z+Hcj9+bXNVtfYHtsf7SXW4Hxp2GaqOEY1+1am
jkGspMOpzZMDOPoUz0x4uQE957vkb6dB6ANCIBf27nZ/Nj9gk1NTvEHFZGc8ZbaI
Ol07ROvhTeuqbAkVIUP1g7MA9BlPevX0+aiaVlAcUCiq3bQpMYNPku2sCpfAbOnI
Jumdmg6f/hlB6lqTodj7pV+ndRWCN71eoRpjzpWhhwIV1j9DCI6bmT7ngT31odyf
zoB8TlJF8zkul04WiRJKTucxpUNEgf+hOl2NNUqSnDZN7ndpweSS59ZKO83Sx2sc
CUtfzXYoNT5qSbSvgbMWs0qG8Fvqlmp02CBdfelj57LjsnPnQPyPJoeS3U5zUow/
Gxx8xBOFI6gS6xuaxj0czlFzbHu8+82m/0SLlS/htB0SgUFL8jHewjW+HBJUlm5m
eHyqqLRzPCQEY7okBFq/hRjkfvvQtkGd45eEllhy7mUjeC1LNIxp2+MdkzVbI1Br
T5OcT9f7rlWgHFCceGvPudH/z3VMiV+IPHNjUP8LMQMNLGy2I7pajl1CZ8p6mSub
zCj997Q9aZgne+05gPAWhTYbBA3y0H+kMrLK+PnJ5wVXbsoGhowxV2XlAS2244hR
bnzRCCbOMuZHVbCKZ6q5J2T6IuGOt7aUZKaYv4dxeBgvZUpVZE9+Pc1MGPmB7n5+
6IfuZAiCf/h2ReigQ7XgoKB5xAqvEnwkCu684amXI9jzdPwKmCscsTdzhMHr5rDi
wDoXbHy/TbW14N3YgC137NsmuhIexsRZ5u8er/BDKDHpedO8BY4n4W2eK7eqOE57
WSC+qHuKW9M6YAG3h1OpcwzhdSOo2n2/WJ3v/ywZyHgWBUCmXg7QcHi8DRppIik/
wBn+V3XqWwK/Ho2P9Y6dUC7+hdnbgU1KFBH7UOdFRGMlU4PxxL06QaJeDg7sgfPv
2uK92gwcLlb+hAIcjgwXAjkcQyM+I+UeDokv7gas94wEz/RJMLSdAtSRmrPez57l
cU53oxrLlbb7wz+ZTBHAkpTS0YaAqwC2WZmLajY8vK3hww9aeD1757WS1FQe9j/h
UNGWpqasSagco2S+i4aPTpriXV1Evbtw9LZja6F1/5LBIRKi/hiIl3f/wuUEH7XD
8whtVslmb9hyC710gpHITB1bfP6ujFzPjUlUYnhprvhdYiUk0gwkePGlRmM++p/p
Z/TbapA4smsd535hy7kIJPdfZQsSx6okFUdApK6E7icrkn8KwRTj0WZjKRtFB33q
8tYWq1YN7pM7GF56DlNiOXobCnLEdEZC5B1yg13YxsT7/ZHN1fq0AS07Pc0bAnGX
AmTECNgaWQm2CD9U4ejuha+vtKvMltoS43xOXt8SdTNadButPKH3dJzhOaIjVZ0c
Zsq5cZQKgtftuOJKWu7OsAA31/O19WJNPDWiOVfP+jwdnmRB3tUhkPjeq5T/Gaa/
8MXlvCtVG7xVd1YByNW8JjxEmlyWvYUqyazRrM9vmaF5h1UuGgRFLqgcWMTUBjjF
yyxK+Wbz0kianuXR4XbBcveaxMXZctQBBRwQT+DqfbCX0/erGM+deLLCHwMDa8x0
Sgfdwhhes7ZhlasQDBJ0zBgrshJrpALH69c3kMPor9NAvXA3ETX8E/lnvJJcOexk
gzc2XD92UJU0RSu9jtuQAYO+ahSi68Re9lj96c0NAqn5IjIeUbf1ZXaapRb/VVrk
PNJ5iTirS4b6RohZ6hzGpxXkhDrRoKJAk2lZ8PYiX7q9xH2Pz9fbCLduhXOXqP3M
sQwlKw+Spg7pLNsp6oOZy2BGEaBJz7nnylJfWl9TRA8WfmRxiiMTbphcnagr73gX
rpxQlewTcQ+KWtxOljECkHWNAhQ9suay2nbSv6rkAPogkfRTKUNfkal2JlfM2/hP
ugPEOsT0bog9Aeh4Nw5g+ctBj5BgOErEbrMMv+uik9IqMp6usWlioVoDaPe5C6Ae
nLq4LbnITiiN6s49y7Qm3J3dGmuTlvjIyov/pfzSx9erVKPCszyDVFrTfDGngaV5
ofbWG/X0gix3Lz/P8AH9Z3A0jDyBcc1XQWLdhCxN8p1EhELY0Dv80GfJw+bLhmnr
gaHnkz7vIckcDDUTYenWMXVuwKwEOrnWHcxwSKi4gdF9P1NXvhvyJjjUfgRt1arJ
6bYwkGXy9b2MLk+Pi8jAuPhTc3yf8oNEo27knET9EyICJV5l63DkKyKUVsDs0Hm2
6kVRFhNye1bW9SZhOdd7fuYucRGv0OyGpcDpGqRtTvIU4pfHI2vu7urMZmuZGY8b
ITdO6t0AzsshbBz6uwO6KcWClO38xND9n83LksMwU9LnhZvqaByz+pi5EL5UfFeP
YYNe36cgPMSbLx4VGgYIghepT982bLIofyOrNMiT23tuXWF+xcgo72136IvXkjrK
v+ZzXmqkx44hk+HfQThOyiTo/DR9Nju5JSB5B8cagXG2bt/zUW5R0Kc4Fs6Mxs78
izFZGPgUnX7xkOxlX9jghb8AfvJ7ksR7Sb1H6GRjhTG5mCMbLPIj92wWS1Vk+wRI
w9nUFgePXGzDGPlv8epeyZ5ADb0vkD60iGHYawGhguFqLKB4QRA/hnkbXY/MuLPx
11k3uDh6IgFEsYBG7IdhwswdKJ27JEEClRjPrOzzbRgJpTCO/29VJL+9YMK7viSL
Z2MzXQ7PNhLden9I2P0KJeEiFEtE/qzSdhNq/lqQXv9/uL/bIb75JfqN/OBp+pWR
geOsJaDHNkJ77eEfgMSgiQ9s8qMlBOJUzn84udK64IggWdkyOxoE8NyMM44HVD9F
2ilaebT3z+gWS/0F9mET0CUW6P5NhoifLqYN64AMZnP7VYI9Rb34gdY+mY7IyG4b
JCSbH2svU+JR6a5gtv2E0xwHLRysFStxskItz7w8RHFKgeQ6NZIrqBtNFgYV93Dn
KdnTb77CYqEQEi0MaXoggj7NB7ny87+caTafNAXbTF3ij7/LxVKGO4bcMc7MajLE
6XUsoC1rwQ972JlLMO9m+UEgO5RCh/U+hftjxaGtC2jLY3wtPP20+Ur1hwBuq+z1
H8cnyr/rRHXQa+oPT2+gXgjPMCeWbWUp/ZXWNYnuEr79uXW8bY4pVhXtnlWSB6Lo
MYHXfVy4WdaqZN/EAJiDKF1tVRK6XmqD3SVLREzkwnnK5Qovwp+R0r0deMOwWd6+
58X57UUwuGZjUwdiN20iziPSkEdzWzkeRSEQj//jwN3rLgCx1GgY11f9TaKSApvU
WbasszAE/HS1By4dbjxciNt+AupStV3KRi5qCH6u1SSwz/oDDt69VqU/BGaFPP5J
QpB5xaQ6uUWRZgHz0KGjyWxWDEJDyn2kRWILZbH2JwG3Z5jHZMaJvQvk/O7kIKRh
DcwPvRuPlMu/mte7sa40X7eL4IZVNuEadihvEU3ZteriZGNTqdlQGSkSsXnc6J5j
x4fxA+Zx2sKjA8jaYnDXVpoktd5d1h9tae4+2bJRq1PIbR7rStijXlYWh7cs+9zW
nh7fFJ+x3DB+txZhUYlNfVkbryYCnjUYdTj+EWUfs1d3W2AqD9bR/TeD+tJhcq/T
hL5RpP36U/AaMlT11joXDQgoHvXhOItQyr/8rZwMmdmNdTyMZ3sHGn/mIR3LSrmD
hZiPjGxxd6MbkZL/CqXDtwbXWy4nGA3eHOX+4UAEzcTmPqDXeco8ruom+zuKuBqN
LwKQKymkfKX9Eg5SxvNkQWdxUDWYVRn8MDzRZ2++XPsXlJfgvuInf0jbxmy9DAyH
9M2o1E3Uh3CoI0Vl4TrOoQKiO6d0YfcM5HfgFW2grcJjZUhIfl+goTauDytazMs2
oOlbdX7Xz+BkGgXptRNBZwTrNhonL3gxPXo8lH8XiHodE4jEp1yoNryKh2BIunCp
BkyIi9lCJe/sStMKIKYTNVEkDv39txSyOpktqbeLkxK9pUJzAQce/brCW3W+XTUP
kNt+py492cLgI3G3n9NjvlhSxGb/GZM+TPZAkMoe9iw2U2Ogf04fKrTSUKQ8GBd+
5aO8/nh/bFpIEl0MRtiHscBvybyBKMEnwfb+5nOZHXryca3eF7Kg027843GjH87U
G8urJoMmy+hCFmAak1/kQMzooUWx/JuNMkgDMs8H8Yt+HW54xCGLhE4M4Lw2etc3
SeEiOaZqfpfC+q6Zt3LVQ51skx3uosXX79Tj2Kf2OG/J+WvT1HAi+UxyhztnB8pv
ifhwYdFDzHp8CaIvFTr2svwCc2YjKG++t88m1iHpdB6ePj2YhYmPzSLOnXLIqB5k
e7kNJyRlYZybTKeP2kdi4N/H1YTTo9aWL4dfvmioNF/IRC6SxmRlC1sS2tdaFskh
zcjuFGeYjfa0C5wrnc7xUKPuUoRwDMctmBb/a9JtzjiDPwIYTWtMjDJpsAP3TWTv
jr8uqZ/nBqsGBafABdk/btsFp9nfe5e+5g9dEMvU7Dqoq1D+uzt5jthoY3rF+jiI
wRvGuI7bGENzp4wfkKWW6hnbg7+LZ04BypUKKNzh4X2XaVTswXv8SS2xuc26ejkC
FWy9+rHLwD+i5R3RBSfyfD1j9PAM86qnkdDZfkTV6m5Ck7E4tOVRMGZpbwI0+JCG
ptAz6LtGXI9aG0xs8lrv9E6/jkjGrx7Y5rIdB1T3xDrdoJOgOrHl5PFNYtDsYVfZ
zudBwWxEl0o3BK7aOvKZ8rxpJ8RS2xsYy0hei3B8FFs/D9KJfuWQLlwoIjvCIEC/
UCfX7nLhmKGtJocry9Xp/xixCReFXXIywlgciEihv0Q2Lp2m+LUO1qab8X0bQvrM
mKCQQmUj4HP0FDJA181aVSjjxj5yqJ40bLQS3OPCjkz5UrXfeTgIxHGZWIBYXVq1
iM3/fsnbRwIUj2O1qSo/cRB0vbyRVm1IgeFgXIHJ+v2h+nWejIYBnvDYyavi3FJ8
jAoVyO/wfWtIzYrHvuoAkqtRcujE6w+yz/ZdV5pkaTxtFoEzRiu5FmbNEWb82HsE
MKWpANYLrNIrBDyUbDRiAOq3UZWPWjCViAs1Va8o7Xm2cBEATaSX45PJ/81oCO13
lt8C+wg++GkdSrTLMFumhOFvqREi7xXaz59ewD96507YHgIpB9R3sotyvoFXs5bx
3QON97+ORXijLs1eYqOkMMiILevK6GlPYnrIlltpibJ7zC75N5ZBKsI1p+n7eIMC
yF6kStmGkk54CKaMjWbdzi9+fTZ1iu3KxHQC6wlNiMoEKb7HQx99Mc8ZThE034MN
O1pszAwO38yQ/UYrfd+J0GNrVGc2EUNo14s6ZT6xKo/F4njakOlOu8NBdhd8Daj0
QuOmmSmvGs10ifPqCQqpmHTLzZooMVYRYBVwhN0zWmTVNmFQExnSW8kLjzkZdklw
IDfUbb+qmXTgZuW2jvjyJw9jJZGr5B7VMq8BmX6vb2PmOzt1JOw6Ldq9mwhTcoqr
FlMCiBL1j+nXsDB0iklPEw73sKPC6/fdByevaoVhThPlU30fzJsWr5E1JB5sCPDB
EfuuA0J0JoA3eleJauHMq3EqOEYZ6dqSrRVpDHhMPS0hS2Zkz81YAN4TAbIsPrIg
cf2rrQVaVTH2uk10udBCBusz3g4Bd1O9gjkz7osaPExFT4fa8pzsrz9k/RqVHdOO
Ls/6FLjSXNvqSoyVyKAYXxPtJ4ayEiCu9lE/dqpd+QgzKGwVZujTk1DqvExDOEUo
xYPt0rRagBAl94gMiUMS/lXbyqzq9DERrC5lyUNfr++MXczIrmyNS3tPZCiFmtHn
fjF5h1e+HyJ59+zknr6fVnDrwjhUSnBaU0C06T6/sTJ+2ZR0Z9/CwZq9bgrgpKhZ
9m40XhtggYwLAtoOO8yILk4Ar28mDVUiG8q2IVh+gCB+dvXc2ALpiWwpGOB8cxrD
7i+T0cMqjMMiWRJQozMwVROa3nD4ddoqeWFRH7C9xlRXJpmgniunpWVoTbfHC+Gd
h3L3txJMY8m9DIcTzZEi5lm2fDMCfwJGEPTqFoS/ssD68LwvZTz5ffqRe3yskquK
9E5Pq3bzdxei4S20n1k2S+qpT6vQMFuajMikUGTePexBtg91jhAKPxdMV+8lNtAE
+VTB4Zgxt6jywxEGWb9/42ObeetfjNLAXW9LBYtEFlytsMSJ3s661wdrSiT6aNaw
KVyl02sN6OEcEKmvQUhMqTo3HFfMTUtB5VrTpmEL+zWGEX37l71yYNokoQdoijLA
PRQapyb6Wn5/AV1+UxWr0kXXvH/FUCPC0uocnWlu1fhnkHa2PSl7uqeFbyKD/lpR
Z/XgdcCcVR9PG1bDJoLiUSacK9YWS1WO+s/Fy/BfIoLnEpgfS8iSMo+UlbRAYZGl
bkXt0yN/7FrjNyhbpb57GVHWlf888IUvXSKoJJbWVpeA+LTeJ6R/PHXGsA3lM7gE
7LuDeJnOpfR7fG5MS8kgU1Ir+g7fPXU7anEVAQgqNU3LwkVSaOGD6pDqLZEI2Ywt
J/bW7o8dLzItce6+1RhU1AbcDqizfjgwdyrUsU+Csx3Z6bFilURtSevgo6fHWAyQ
Vsaqco8U6SQVBqpMt33HIv9V4/trEpd/bndTiqPYLujJUidGAp1OkBTVg6Jhdck5
BQyxH33YIGWvyRy9GlKr4ld4gXAR5FOFj4MVWsu3hr8vCwQOqPDGnipVg9znwhJi
A8XIbH/I3OgfQppitFnQsHu9QyEI8uDT+I/RlsGF5/7V4NjnCMOK4wOxwH8+1I4T
nLN02I2AswA7MRYHfwmMn/rEymn9hZkjCvAjuI7Y6KG7n3lIlrEOvwdMnCUi5Q8v
fEZXolWoRCrbcG1QISNeMHpJ8F4KJU7QXdB7+mc5XIreyZebP4z/56YpPlAeJ/k8
Ccfi0PtKz2lq5KGsrCYrp55y6rkl+hBfVE21MNVVoQ7ToQVF10oW/oDdq9/0+O6s
qeF6go0A6mdHSYR8IwRTXUpN3wFEKNTuFkWGuIMOXZchpOfmZ008+DKcGrds4QTq
Ml+qGiiJC1Skd+GZvYb4mE2oZ+a86Ou0u6d9IsWwWKENXbQcrKZrgHhAUOKFjJLf
py9hZpNj/6ylsLuOav6FYQKpTONNOmo6NY0z8+8Bk+NJ2LDvu0pZQJvzCRIaFp1z
6/c+Mkox+YJyJvYBmbf49vQmEfQbbFtDomRRwu+ZEJCmR9EZ0+Gk+pTyV8orD3wG
R/UkFbvCNtSbdrWwYcyBu6VESqgoZqFRd21Oa+OmwGz/DcgHouGvw9x6Fj1/rZDQ
XX7ZqUIF7hQAuIPK//0kHdw3U7C9RtJcmR7UpN6dcQxWqKeYV5IuW2Mks4/JAgJ0
qZ7IFl0yP+Qoq8eINcCxOPJ4rNqx470tTq4GTrRwPyMkgNBmu3+suXPFrqq3sqy2
yYn9ij8VWSXFPQl7CNyxEHiPrWK99mX2GERskrccFJYqZpqizpu89Pe0maaeh3kO
U47WD3S1xyEjEHaXjirQNIAqeyfCkVtejgqDRF3LacgbR8pEyEP9N+6GrhZryVn+
2SJHjAhKRsoaHuFppxldeLqnCGqA+AEmbAnEfWF00ZJEJHeEr1YTh0v4yER+86Qg
y5elYaqwMC0RkY0R5y4aznT9FRJfif6tfo0GpXSg8+OKgtGpHyt6HRcjevMjsxnt
f1sh3xcV2R3GDagWvRjflM5tErBRnONm/7Lybhe4vNTauuKetibW6JYfzl6Ll8c8
CLEQC1fYI8bqcrZlWitQqgyktg80MMMcufM2PZXpbZn+fVYviE68v+gVMsWdyBG6
OHYD5+lbcDYrmEPNGZYEkyBbCbv5yyPzvnFNjXSCIE3AuIcl9ReQ4NmKbklFhNt+
ED6EBXql8uL+Ib9tztt46jgIMkQjgWeSMIALOIVzkoUr8mBKnRuKaQZCN0jiXma8
ZEBLKMvpMtBriWKSPyKTKQpY8xT3xmH5KQq2vsFL9RJoWpblbAbmia/Ppa3tuVqv
oo/PobOvCkvxc59IwGtXa5+NMvDXPRiEP+ZX5+uB2npkdUTOMQO+DN/ygPdcdF9U
wCGOQjvPmuj9B7GLdc5257XFXmUX74gFIDfXq/PtJPUHdNPyi/+8WGteKS6l9LX9
H7LClejFcKBmpQLWL1RbL9bX1pc7lyfIJZ4R/+S6SVioP6Wqm6Dl+iIfgjCTrtfV
M1f+EB3WkYnnEvqZ8gqrFzb8nUdOFhI7LlGGRPf8ljFQgTIJXiTWGywIBkTV3TmU
DWFRgDRkxDznYSYtK6zdb7ylHEo+wdVs8mAhChfgK8y9S0XKHstG2igFMJ+YzH1O
RS2/XUR+LHg8dC1WLE1wpZ4fY2fW4UrKz4NhA8vtpP4Ia4N4z7XaT6bKMz2rHpss
vexf3ns9v/3bSIwRK0vGR30aHxaXphBF0l2Q6EmNu+gew4nNscfhkpJqbf6rDsMn
0Tfv7LLd8qTk4Dh8l69MPgxyxfjyyS/S8tBy0Rz5ayOwS77vISRmFB5xzNmuleHt
0eNwf1MIenBSykUV2vTMa1sN6WTB5cWJ5X14ejNnaTeq7YIk5ye2bJAqeYYdZMFW
UFaSgDOr/grEqUyCGFRJmKQRacAsesMuIDlEG9GkxH5z7rsNcUqIoKzuNIXhjmIr
zQTz64Rq2RbN+vuL2pH3z52dIEVNrEbw/26FzHhs5AhqNwxptggHXzCSvDm4BISq
3xmplyJ2vQRbyWcyr86JTj71P4188+c7jdQNJoI7b6HUkXBEVHdKn8LY0Pz3bhCY
+/JFG7Cq/kVlyDbKZZdbXMJFtCSzdALZ/qYgmN9DUPFe1kTZJuZtAE+6pv/0LAIG
+38IxjVChvV9soY48sedjc0JZdn62ql37dwcdbKjvuF6atowZPwTfI0h2uR2b8uo
XPkFGw3OgMxLq6TNgVvaKstirIRjo7omkI0OgBqIpYf0Jg/QHxBE00OmeTb+MWQm
XZhoF52KB8jWvNV1Bf9H5xTiNaUcZ3Rz67C6x/UMXdYoTewsbsWjcH2m9XaJZx/l
gk5xtwE/a03Lqf2f492GFJ9G04Oli3Mymf3Jd9W1s7+KJI+yLycYqp2gZpjpX+6L
MLwGTObR8TuXFhX/BeT2UeFUm6426+wlQkCqF0JVDYXDIw8eDss0B+E8uf83+qFq
vPHuX1XjY2Yp5W6qsfCTzKfgb0Ii96yCHjOpbwU497Cs0wvvptzANbF1fd1BtYhO
gejohLS4cqtsMM2YOUM0/Ue4qycUpuYX3IUq2SPSSDxvcE1YoJb/XZhzLobdaLYA
VtCvUDNBFFbmF+NZH489a6MdtZf39DtE00bg+UVYW/21bRlmBrH1gJPka20vkw28
3NH6ielBKlIDaVMiKbzeoR+w5TUIeRnks4MnLKtmtyGGFWZE7snkCJYHPJH4lbaN
u7KAJzPY+C+cMybFvM+m8FrAVnwQ4PA+fmgsv+hJvCBa55CtnZxyTC2C6x8JQa5N
gC09tTJ6w+Tvr/kMJPWBgGV+lVPZguNbhihj1YQRzDh4Znzs3SRJPKczG6zgDJSt
ZskKymF4LTeHS8REctG1Ai6JHbnZqzsjrK7IIcRlz4Ezz6+P9LbRSI5QLBPADXyq
/p3CEntzGdrLr/vyri5Kv/PsmB6/xPowgwnaYWD62VCnUQ2EMvM6baBfDfW4hcFa
KaJLqz9gpUWThVs1kKF1ScN9irlbpppLiNlJPot+shYcqz6eOxT7e5LRF+/rODYX
B/QOi/s8R8dUeRLGHxhDoIy4sB8NjmrFZoEYbL8nN0Y+7UQlHOgGK3fKp1sRqRhY
r7A2U6KugxB9eTZaFo59FhspzmnGWcmqLY08+1Lko7DuZs9N6PMze85YxIU8UIXC
LXNExmYe40NzzLjL0lRccHezLxiNvSM5Ybbmh8Ci4m/rR7LiOaaxzKcqT5coPgIi
AYdWAduHMjnqk2CaBXwBZZhMGiLNyxr+QBH6Ye0jCQoZVkvjgNM9RnJaG0YPbaP0
7WGx4bJ24W95Pxia9fK50AvxA777iR469k5/ruAJFYrge/7xzTuL5DwDHIgTRfSr
PZ0X2d2U75oNjXpsi3qIVzVqP8HpfI+sFMX8iSA7Gk1+yjvK+KCpSoEIfIQ5onia
/kz4dAspT1SbkiuLgK7CRH3jNh+ZlTP1VQ5DIaX54ztZOcJsQNiYisH+C6TYY5p+
TjVbkdReo5FMVzusoDbw2BXDzxCng4VtiMK8DOaUVgVQspFB9x4ZaX/f27Aku7Wg
7rShhb5FtxpXrr+QogRTascmVZctkNCPWswo5bp6wfWbR3A5tNDeq8owBb5eOKZ0
E0vLYBz7lreUIcMY4arBa2pPs4ss9Hhi2HOv5iT4yjZkSlrPc1u1nEo1C6eFdSNd
tZvqwBNEhpJjprB87gpmzQsh9CNw+RiqPzRdQPlecsOCzKLQIOwTA8xydftHPsMo
aIHHj2/L8ghsTIiGH4anIzA0sRHzZNe6gFkJ8SF9UyI09fouS5XwRbZOicF8HpVy
zfyKePMKSk78WxoIm4xcQiSBInV4D20FTbiPed1LEe4Kh4KJ3K3IWwq2FAjKF6cH
OPF3ibVnFNEakdM/8nTZoq/Cebb1Fw8vjSd+9kXEnVsueERlp+aVUgZHphnB0bMi
GlacLozfSausVxypmiuOSNyzViShtnSFOxptUdDzOMZBDaBAIUBZgWe1irRrOypK
Sdf0cp1SV6uBn1OrLZFrrUSFJRhBBgd151gqHi31cZt7n+69N4nH7fRGNmcNMomf
SdShtcw2hTMypryfCdkUakOOobzwUpKmFvkMLwUUc0e7EG2r8DqkVUIwaIishvA0
ZJTKHMrBFgOh4i/HfKX50QjNFlwjZtRcveY+S5cn7YSWnfWnnVC9YM01CMDjVkzM
4kIzAWc3ruYwqpt3YYiNQD/pBTW6Z2rBwRfFka18/LgLRF8xfBdQHLx7+kMCW4qI
8rlXZf1l/m8ybCTlIhviGXAW4ZSGdnmXTPz4no8pCHMAU8nnNpyNN2z/DbG/qIPP
tLcc7ZQS/a5DzIr6POp2B1CwR94drtWHYOkm6w0sasbKIpsfF1soEc/XZoy0nALw
cp9pqQ069T4fPX/6xJq61J2R+VyB3V7EoHRyxpqGVamwwz8EpRupUhHfZROPEf9i
utqbHDS1AtO3Oi20lkRzCOOJ9cYHmZN8bcLRrSkfcqEX9myLIgMQI1pJdgf8c/dG
HdEDB/eBptbAVhbUquXh1j9NcwaJDDq4c9CEEikYG3iNr4iwRhCK7auvtRLhoxlD
ptV8jSEFrBP50VVg+gLpNMRquwse5wdjTiKqSyUK+DLGmI9toQ5yq7tt/nJIQjV5
Ug1iVkRkW4Nj9lL7bBQqOTZ8PLAR0xTSl0mvZ7eLnbkixkBqT7HLnYN4l1WK7tFt
YV0sUsLWkXYtE7CziAMc7+b0Wn4v3KMTa1yIq5F1C7d6gPiv6wURixESMG0Iz8ID
vjYDqJRisziNCZxwt1OXArXZtWJs8TnzpxvD2Htave4GCdc3R7yhg4bfF0cB1cKB
p20CBkgJhod2V20xFxVaH+aLYdTayASyH7vVW1c+gDjqWpMk4oJFGaNRJPhWk9th
Q3ivkNTOR6znKDQY5RjmIZFrc48kiBoHLGnz520AAvE4nbrDDZC8hTRjReF4A1GR
On2IkRTfxFjvHD9mjRxCDVp8aCp1UOGhfL7FKqxfbHXR8lN1Q/4IM9pajIqWJ1xM
ZAihL14Zsxyk8QP41r0faV7AIf8uAR9TfdY+gH18ynZjd6Zt2nSEq/VtJtEag0IP
msgs1De1X6b+8ZRplx3Pbjr9TPFXbTuilNWvcIo59lkhS7oxKTr7cudrWKArW5AN
OLm/2bzKb/27pzGJc8TvriD3/Pv5WroFCYm+ixtobjNZu58rS+wM2AsEDS78vmja
Cmfzn2/zs34nyIF0qMe0Cv5DP/9Bbd25hlU6EhhgVb40jWYLQneh6srUD1ezdQ5K
KRa1Eq70fuX5RzEFlkGpDlmh0VfcDwMWLcUnuacAX1jiIJbDQ7g0faJd6cAdh/nu
B9hXT3gzPSj/X33infIZUHubJLub9FBUtNWNibnciRwj7qIKBzh05/KAkL0JmYfy
3CY+Fuca9Dc5h7sfRvHBvDoIUIHmriCq1YasN6g5t6yjOxyVeHqxYb7p5lIfsGS9
dnU7gY6Wz6oY2iQngGkc8rfiOVWPGz65Aix9RCC1yKN1B3q63oIkFP0WgYBbIVcm
WjS2BV0d2KQ95qRdIdU4/GjCbC7fcoJaeqazIXYl1uAgxLQNZ7m6Icg0Nwo4eWeH
yMI/nsvhTQSVsR3prNagkTGCZwp03ADkA75yQrHuOJn7bEOyiykwrh1QylYwBQH1
kv43ViKlc3lcZSWtlGGbnlAIg/DcEa3MWeWSuEi34SjSp86Ph0cRoiFWmJbWwQ8/
gY/a3YjKPRPkkLwNrkbTL0ry/YnYbEETCADN9o/MiAjKnE22sMP1G6v+/3kq0F5u
xITx5kOrEBd6rJR2bSDeDCsvzB4ei0UH//s7UHyj7C2uKgsfYhyZ4vngvn3mWOA7
AdK87SGucwF8Kx0U+b3f+qL27PqWd5yKvII+3pFBbQk8sOMoSOn9Nqf7NjAUX/CE
pu4l4ocekx5zsoIPiWxRiM3UvMxUXZCDAXjICUIGLFs7BSFVEvRfeTsxk7U9Q8A9
9Cy2Ztm5GLzTdQbe9H7G2+ks9qATyJ5hIQSFSNStkymFerGzFm1A9cKVnw0czrAJ
HQjPzW1uNey4zUTsogW9q/wIqkkJ+8b9/SLdmnJu+x8F8wUwYZ9cSeJHsPGe6aJc
vWgx5slg8kLpKoBsN9tDgdaSaJlngVDu9+g+ymhANXtbqOGgAzp/iwWh4IsOIdgA
tIfXiBMXgo7kBHE7icnk+fsxWw7CTUNzgZQ8ypBx3I5mnyZsQ+JWzYyIqRt/hdDk
uL/sqpz8LjDZ01HYwOsV+KoEwxW+M0Q2NprkQ/Bpq0uXjhYZ/qOZCvYjAkvkHQvW
/tc5jbAi4RbXhM6nODP0ivuFOwnNTPYza07sxME7KLrWzLBa8E+fZ2EojnfiY8GY
/pNN84a2luWFNUGgyoIHziLWMv8S2Bg2lAQyPD6K07CILYJ+hmy8qmn5X/xa+1jV
LypAebxn16RMHUn6Jr8w01qynVsa/6r+s8weDjYxj3640yILqRH8KEBBfuRVUGCW
qVMSXa2/8oKMBdvIJK97x03Pkfc5fSNhEP7L1A/pAu32aBbvWicbIKMfAayXlCQX
THhMnHUXJJQNNeTymIU5p/UEuLDBD5ht7R4j9GMTr50Yqxq1zIg/RsPW2qvl48vd
FWPimzyB3132qE9EGYIrvAFgGseIifMWb3Y2J6mB5qVbwyLrfyQ2sp7LYeeokcSV
dzXx3P4CK5rYjlxOKtkC9dmXB4Q4fgQP/52P+GlmHDBEBC98qEi7U54jR533byEO
KE2OL3Z/gsbU/Wsm/T5nxP7DyB4biDWas9oJTDbuViVHhHxxA461oTgrea5vJ77w
8vznnq8z9gf+9g+1i7xdf8mwosrQADX0QR0VjSfqkkt7fPl8kFDSXP2XxYld7bKH
XF0nWXYWNfINHpT9uqEJyM54No474SF7dw2wdml9kNhQP8hH799/yZdQnS9w7ug/
SRMyAlIpJP+N9ZctLlClEEG/J0QOn3l10QACjkU5Tv24I378+u/l/uGOr+zcq3Ny
FCa0bUyDt7QjiSQPhq3KZzvD54y7neZzb3oByvZPLFVumAYp4yHm6zVinGWR0mea
v6/+RnAX9GlqSzwMa+9XqxhdQ99UzKSgaNyJEqRg5jFFeTCShC2dpRBSJVLe0zvI
JzvzTtuzT82TR/X38pWHgTbFokEegi5tM/6OBPOfGxo440Wp+vl8XTeo5/waD+xM
HN/uQgyEEIkWEl2lVGzX9KuQPXjkKKZkeRMCUQXCnDYrH2iv1kiEhE+yBavkgq9d
XYJnO7Hk+c1po9Sz7oSNEVWRXGtpr2MvZNQRRx8q/zxrLvZlDuuDHWcUfacSadx9
j11ZGV++1uB6pYtLG5DxrmXWd9zW0bddCn7KGSe1OwRDzHZLa3thWbcrWlWPEY5g
nAFz53iOX9kjyZH2bbgel091Pf3R47x+o38t16CpQ7OGrfzwz4nCRMAuGO8XPMW+
qRAAWydnOVX29a7Qndfu/c/wBJpiScfUz/OaUduGa/puI+PfOo4owZ5SQ1VX14IC
pYTSKYoeZfNTkPZdiGi/viPtyCBoh/mygasYX52u6YStU9bcF2rHWVzop+i/F7Cd
TVFImUy1F/1dfMhz0rZhSzxgLhR97XwUnrrCCynD+uMoMio3jF5xL9wUjrzc17HA
9FSXvB3VtH5H6Y2Ns7ac22bxJJN2KgTJIVByMTvdfOad+8b8/JD1RGmNvpxJjMfI
o++6fAlyO1neh5jMQKKDHwJyMAdtPLX8skb7MIhBOIWuc0cGLGfvANc86DQymZWi
yNy6j6YAr6wI0Y6/kJR8Jvh+iXayDkpRWAHRTe9sj/7ctqgux3pMdPhHPEjI6vu+
b+ihKGpas1H2gbZDZMSDH/74shTe2BxuL6X9+DCybv+57jJ0yxAx1Wu8s6Nw9+1N
6QptMYcikmRUuNi24lS2Rgw8A82jV/6NhVzzODTAIRkqsG8hHEQeFB19wY/MzP2X
aX1rN9XxmOZrqzYrN9Kei5ND+HZ9L5ZpL+47ppzkFoNyCSvVspbY9AXdU1J114wv
MNKwj2U+DRAQsHTeo2FPwpGEe4FjurvTsErHWGyWy8AUmKc4M3EKMhzQFTMTHr/X
Hw0eeQd1HkwftSr0C+fCE+ReCTB3UrLmBlJ45rIkeHQ0je2knCJC9jl5VJD6Yu8P
XkAH8OJVjWtL+zCf9PW/2ryO++vhy67uAWFzk903jdgFPXyVHOPLi0+QETeFe9/M
3R8hDsP5GU22JDVqA4K4gcLz2Vg2e9Q7ubNJL2mUoZOmJdrdy7fGDhsslNhERNDy
TwT6gb6L/0jy2CjK6rfEotUysaJTaKL1Vz+ZGX1XdBOnSmxlWUDmQqHHe96443Az
CxtXW/gjrb+FZXg6R4MwZ1OizPgONnIvNkU2FWUOuu6KvVSolOEwf7YaSJR+4vH1
SSNSgDUyspavgCVPNNvTSwhQpzXqrxTbWZiWeoAb+PzEK/Tbmtw/k6N4F9un0WYy
VhxofykTJQMReaLqPzZ2gan85e4KKlW7H/LMlNSlYLtEXT4N3kj27K13M1M9x6Uv
mFaONKK8OBXdNiAtqfvyICSm6KzFVwbdSd3zOzcjbNrszbiXoDhi9HuTS6V2QnV0
BSeoFFT2rgZaHRKrLIuJeElHLp5c9q9a8gHE11NPoYEaQ07HPNIdKLiogg8VlhGz
y1nhC9Y/Hxw9wMj/iyM732+Kz9v+paQ0/FIOjz3PYluVNpAoA7u9khsCvs/y9xhZ
ILY+xO7NbgZIjh9Nn6dDz9hOWKrA9Ob08uMQYzdcBp2G3EUB73rucOtnuaGyUOA6
qFuG9kS305KSODA+6tIE9HRjrcQyn635YhNDiKWVVizUZ0PGJ4O8U5DPQ4c/C6of
pwOqK3Ne0VqMDYpSEdFzjymx6H/36H+UhEEJyCXEhGYEEOjHobNKNIJfTV0/8zTp
TLmmzdop60x7cq70Gz2U/mkRdUa2eadDLeQVpaHeI+NKHGWKTEDZ1DUPNQa6Pte8
TJAjLkNfcUt209qZUE17mqqKNEVphgJL7A6hEZB8n3keriDsCtgGrryvzg3X8C0d
4Ip3C3ZYeQ0KoH/8UKZq7QOHlzvorqAlt+pGFSI+caCZanGgWlhBobUbNHxqWriB
jBzQlM9Nc0d5smX+dvAT9WO83a0dohlL2y2Fhq4cJmrN4llIEir2q+1A3jBE1evq
kZUhe6ilSFi2m7Cnbkgd3FM4hPMeB0DwteRd33uu9Fu4Cj4hS5cYrxImsygt9eCP
B7SBl8tdzgh5m7yJgst+geuUP62gnZO88UXdzXSatJX0B2/m0QjV+jqNQGNd0/FV
aOtMPq1d15lrNZCUi6Cx1JBFbv0WG49xtJ/HloZfBMXREiYsqYxquVN9WXyaZjBh
lThtaNuLj9/nAIjYRhUuP/A8lDXY5NC0M3DeBaxrEAGx3nwHQR1cN4hOVl5dinCI
TJdLP3Y8Z2rUuqUj7bs8oYr6MZPNzkU2o2UwuHPUfrv7xfu7rQfomWJYRd/Y4HcA
ckH8j3AFwat/eU86ySy4ubrbBg9l++VtwpggmbrZFam3SAjkpr+Xxsc7otiVdWka
DBZSzK0V3rMEhsWbX8zsIxM18dK6FLKFIAq6zA8nA+FxZaecIavYJWkB8gQkufoM
OP0tDcvgC3m3bOPigHarUoDwAeszl5IJdW3qIQuvAmJhQMXouNF9e4xPakGU5uS8
NZZBeLlBOiw7iqA5lTaypmo1T/Tt1cxX0nMxKjgc4+6H6J2FKhomhGZ+KKsZSltP
VY28WBGSBCNRuV9TqPp4PpoVaY8eBSSRyVcqrt0I8axBWdqcmzE2IT/jKdx25lhY
G6+IniUM9k/+fi/1CPhuVwFVoDNd0hIv6F9tNIqx2faYrriPmoEQE6p4QhyGlaB1
t1dVfQgDe6WBW/X+KxyYQsWwZcJInr5LTdgpCth8zIiFh8+vYB8tTbwtBxH69zlE
BmuwE4yJPvODoBlOlOPBxcjPBWW+mnhUStGE/rXQcCx4Qy4yNxUcTgoOvGPsNUZV
VJRci/HrD/qH/UzO9sXhIUn3MoK1eaT7N6nciC+oAtSxoXMyu8aByY00t2RvLiNo
OlowdwB2dT3rHqD9Vv5nueYcnx80XmpU879XAI6vrgGK/68H9Jte/xcZTbk16kJh
t6xPxxItO+YqF5CUGJpIjxb4TeZiB0J0XiyeOhLp+l9grCmGxFttM17Bfg9sfxj+
jdqlbQHD5CJtvwQ0awdUqN2BdWoQytAfnwGyM/Ct+Vt4SooJFGVYfm1C3PfCvd59
ob37n581zrjiGzkgtbHAKCw32jzYT3uLBHpGCdTAsh4IzBT9DAK3fvbXT6/m+36o
48scfaFL3AlTprFWe8+ohabGKwcKpHipoyeOpnAIqlc4IULgF01DAyVuxfZ4QfKN
kz8XEowfn+dfMv6xyLCXmUM0u5KXMcK+j61HVk/xM7jzqGJvLkMrrd3N5Id6ZccP
TrMaBp7Iq2Olkzu5ee8cA7bOIbmAQaqTVOEMs2UKj8+5vXwRkL9GVo9eJ7/JBq46
RqYpIADdynOt/Et6vOX4dWXUJT0oeP118Gz9ei3bLu40Ba0hjZjWcGvCZL1YWHtD
nXZXDGgzmM3IYdtJdLCc/nGEn112twrPla+QtXUvIhqqMtsHE6K8Wign7ybgWsi5
fUgTbET3E8nFhbQFxEv4+PLcEtXNAsgkoV8Mc6y2JFfwjq63bfONoFNZOJa7srm3
DYtFLgjBgSn91GTRh/Td5rN11fDZyjiWq1uevqk4cNJQxL0bEXrRWkpdpNZjLgfm
Al7l08he8+GDjrFr97gM9BGTH1oWFEveogGjdoJPMbNlBhvXV1hCU2lTfigH0mVy
XhadOeJKm4uaNqHpKq5YEWeJAl0vllmGBtMiPJuWuvxtCSqLQzKow5rBsIwvaS1h
RigK8EHalUuC+da8/hruaLu2SbdMAJjMdnOTjE9ArDPMACQezWZDBYIEKpeR7Bcg
Y74WazoE8t+XNdQUTepTvDfMQJuELV4FvYt2U0HsTMRDcQ0LcDniGW1JfVrSfxhR
ujmrp7BGvP6dlWM+tp2Z6r7v92hDGH/idwezqTvbK7j1R0JmMk8Ctg1yXWJk/wKd
gV42cyzG63uU6DgUi6gd7usjACYxpVWCgmif5tkUUR8zEaB7AcsnWZ4Q1mJZ4SQN
oQYc0aMykQNnylM9s0Qotpv2WMpPXMRPTGrljtQ6oUsJT7/XfZXLbh8lHps4tvmv
WUiAxG2RIQCenZYgUV0LCGkuBzV4fqlHQZOXakEKEFtiJkSIYqEmdrFDCYAeAUSh
LgP7Xcp8s67s2Gy9cmXGSx6F1PObQnGADc9qafvPce7JrYZgrZPJZFfR1ChcLegi
5QN3WtG4t2wpHRxFohi6X8ppzEt24VLXQKqv7TO1EyBrXLEY29OOYMsm7J2SICBp
33bfGh4XCuGc7e5gkc6vJFjHr139QmThlf+yi2onEZ43MD5MjW1Kcvc9GRKGU94U
W6VWw4dQQRB98iyRwIGT58cXUPCVZO60FSFHZlOxLmnrVvUwpQz8w+BBsZwIRdsN
nzOjK+55pARbGotTXy+whYMsZlXamuUGf8O2fRKnm6qDSPz3bLlsFopQAkMXaeHj
SWejimS6DCN0Gzj2nIVYlBKFYUOFgwycz49bA2jD0gpV9mAJKMQLY6uKjTOuf9xe
/ZVfLtMIhuM7BN5Tss8bUfm73XTq+aRmR9l7gwp3EYO2+Ywc4ToHqRzR2xrDGeXB
9MsBXvl0+npSI3i+kW8WKIZTF8KTrKysWdy98TF0c9lhNny6BoDUc7TtO8FNcdtX
Z6uuIIkuR3KJ70+3o85XwysmCi0aeRQzeBQJETe2/vkOR2LebShZ7s4mJoZAin/H
kd2dRDrD/+xJHYHQam6/3r0wxl/oLLiQvKUF8oh+5pB7LHOLl8cQKjstGd06Z24S
bRHnC7nq2xNCfq6CANsbDfW6bXgTIMSo+to6cJMNHmHWt+8q6R3e+w02GuGklyEz
4FujA+xOLFohKoydwuiiblrmjrj2S/I6897/esCGBDmCd5V+tIJIJHAgv8sB3691
xWmGzJ2cxe7IHyq8mq4+fjX+ioOpos1a3zDCFmJjRmuBCv8IbOhoNzAj6DysgnSm
+kA18HGHeVAC6ixbhpqMlLqjZbM4geJncjN9FqTBi64lARzcHO76HPl9XzrJvz4g
H9rCJejbgGt//wBx7Ssr1Dc7fXaZjts7f8F3X9TZyQMfiOA3KAYRxA65aK8Mwos1
KrNNoIJqs1Lbsq+Ue5PinOFTebueCDFO/h8Kl34MoHrHNydwEdTIKJxbJy0Kdu4Q
tYLj9IMzmaWLwZcj3PYOC73lyvhNYXlAkFee1wqQFOiMTvDMiR0kjAEzdwgMjlvX
zivq222LlhvOcvbqgYBnO5m6k81MKxauTC+Gq7UlgbAM+q3MWOjC7tgSkhkkJ9hf
yRR39UBUa6kKqn5uvTRhjUBdjBgCpgZUjRgaLZgPIiTTxE/WvwBzH545SakxA8qR
HYs7Pi3DX3Jih2I6unthtbnkE5qdPiZwCcguHj5OYqvdVxYUxPkouFaOU6BK4Qzd
atCg3dJwKAc2U6wl1aQw6WeCzPdRKMyOGk8u/88qWxv9RvsMO/U7KWAsh2fxTt/A
mB4AG8veYITctoRPGa4+3uQADhyxMYXxGfHF13zFTBKz5l9lLBLl9WbgmWCy0k7F
cvo2n52dMt9JHJKUWiXiwzxyfMBiSigg1Lwyt3ZSiQNJT6hEdmd+H8agqnvPQHyD
+J0NnXMG26fP/xT9Mx73veHQkkooAweZKisjdRYXAJWkWDR3/rzWMwD+A3FE/mpF
imUgKb4V+KXhxwdkmB7r+EVO6+xr208ZpwSmBb/Xh6UJ8fJ8/+56R/zzXQH3I/Ma
DAQ/7DnPKF3xizjFVwRh6r7S621QfcVc4gqHrpoulS1P8yZ5f1ibdsTJ3R8zBDQM
fXvKD/nma15xJDPMDgB/89n6ZKMeSLjgJZK6PtV0LgcSRt6f2d7s+y+wG46vL1re
o+hzh7dlIRhoQtdHkon1QjcUmwtg5kQAwQxdA0wY6C6P3BVEEXbno51wAaIxOWMU
Vj58NN7R80rwtg3YUUOC6iB2H5ULzS15SyRlD2UCU1L8IWnI8uOyeR6k1OoBW+yH
FPTby3Wg4HxkoK8nJsUeRSDpv/LI0kbZAdjfJCHyIqyHrPCJJ1cS1qJHs6qkPffW
WRZWjcd26DQxgjq5fNWPUb6fvwiVGuRpFiCyED2GHXzraXKZfQLESEGDDX4BnPbo
lTB0HPxitU3Z+l3P+W2xprkGB4LEOt0hvYylyEBgcBUj+XTAc38LhpBhJ18OojHy
9GTuMRYe2xvNF/dAmntnTwsGpwbgG+5zCPST14m/tAWMWR2Ej82vmL41ezrkPHDR
5pFtIG0Hf6oAJsIcPbg05jvfHvJDNN8VvkzMnSHete+eO8CPCEaiFY6zbvbm6XIk
DkMeAqMjjOpPtb0jA817U+p8+mwzWZ83ejTiYbG7er/zpHsMUWj3+Ef7sNetz/CX
tlv0HylQ/7GBwqPl0RLGAmcFDdij7Hy+8a8dvaiFrzRAyMKbM3Ov+EPFHUXZKrvJ
LaS0EsM/lC26ud9LyvdyGTn+L1MIRnO/UrQhy7JHVvi70ukrBtG6R04UUwmh0Gml
KttCPQolPQUbTtqN7yc/ELQla7ar5OJBjOKCOMwI/XoQep0qrKUs6mkvuSVoPSIj
XMd+GSOP0R7pQu1rc1SyrOwZ9Jst9WyfUSnucb4sIPscKy9fXx1/8eNBG76YPGuH
MWOtwwycjXz127/WyqtlzMYHXN6dvOGSmPYOCjmav5B95pXraZCHtiwyD+FsFUuz
3mfj1+UKjvnh+gdv1z9ixcYB75AV3vjEc0L5x9aIlQKcFerD4DCBD7Vekobni25t
746gLstdcnJZwT0gr+xVa6Q6XcUsUKQ4jd7h11v+lLYGcg/q7ucmo1i7LG7qR1im
BDCUBDGF+1jrEDZAgP/9zjuZDh73mpVoUjOATgW0lGVI0tjEgWp8ilUPGj+SZtUo
5v2EFWdU9X89UaqRsspBbqH4nXYrsskbEsWdbVnQTgRTDpytIgDHJDMIV9fm187r
oBSk3jhmYMIrzKqDW1iseBkVttKEIL/Qwub/4+jolKlJSYNyUarN1YmzW4yVIAdj
1VMw5acW+cHOHH5NOIBhgq7QArMFxUgGE1Shzjen044EA0D9vQLCPno7ewg5t7s2
x81LHmkBz/RKMbuL41EbfKJL9tvC8r/U4G0lo5FSuKRhnF1DxluA38AmzhLKWeOu
94c/h9cjF1dfdABdNIMiQd5zSJ4vbNaoRXIYz7YgPB84aQz/7vRU2ZfITqi3NJUA
ynStvgu1rSV79enqzWdsrbq177HRFLJ0sk1wKckyaQGEYZsfABZ8nS11rjALJez5
FibZjQSawXCBpl2Cz6/SzkNGqdNiphGglzOa3OT/YWQuOdpchXk69C3+cGL8lxPE
0Mv5bppyf2khKvq+mdTFQSQruR4x6QYw/9uGdzJ46ZahuEiZLZ6c0svEfCQe5zNG
hGrhQ44JtSpECq/2cyha/OBUGoE0UC5jkmyTUFwyuQ56HpwUO7mnUBhB6a+bUOow
6u8J00uFA0EYjdXoem2bpNISeba3Nj/wmK1eVPuWw9QIoTBp680jnMPD01OWXXjp
mGqZVuO2cVlL2zCSZLAN3sgQJAh0WgGQ+fdALGZk7ByoaWWOQ//Dogsntj7qU8SG
qi52cQVGvJJWXwEk/wiHg4qAWb82yv1Vw6w6dBmvwRqyUeBvI1VTs6Pu32NgKuhB
vbBPnGM7PrFNlN33AqsFpXR6Qdq+yIlZKAFd0s3J5yuFVqGakRbJ9ix5wlTz31g8
CY1D4SVL+75eFCkGfGenMAk51IQiI/r2/Br5hj1XjSkl+hfVupjwHHgXo5ALwfgU
fAlyXa9wrPPg6IOxTW/uZmT+hodicXiSjpdUOXhTUXY3ZEEMAGS6uOmeC7OCDVMF
w+rD8LzJ64v6lcRNvXyyrPgFAFJRlKiBNfW+aZVzgDoh6I6+KZXTBy/3dpiAZKw/
GrnKJHHn9Ggeb9ZFP7BpMusniwZSsJgx+1j48HqFdMp5kte9Fxm7XbCWXBnBj8IN
PK7CXlfD0v69KLKyyMLmvClU2Lr+QPJCk61xOWxhpiJJr9v93vH0aY5LHIkslO12
+zDjCHn4PXEUxmeDCCM2UGJzDz8SBWE93gg8oUwGYoFmQqs22rKK4htTiBkD5PaK
NN7A96TGFQ5VTSHiDIMCrAi0sMRFR1Y7CjEkO2BlVEGWJi8I9q5zcDpb5tq8Go/Y
HHvshvRlWfd9J1J66xtqGZOgC1FLH833/396nJ1CTTwKZZK0AmcwALBlNpIfxWHe
ubE1e5mnIC4T9ruL6Avg8RxJvw8P/4W19KkHCInDdwO0Y/M459j2nKHCOOKqTQvh
yv0+GOdzxgYiETUNrDZXEgiD2h7Y6UonKa3WPyu1BeIHXmduRtQ+syFAqUkwxA9M
DWT7ENrHYIrFiX9K9NR0PpdE+wKeWfb174oOmSctXOAtUDux9QCGr+wIqq6r1Z1y
pZC54FruXLBPKmN5isIaQMJpRtHBjRrZo52iTBtKDm2LdJkfdz02OGLNATxTUi+d
uhh1EZ47SpKzd2HR0NidYfYBeaLZXJOaa/XA6Omu38/I6+bQTazRlnXGOricPuIn
D6eyzgazXMdJ2CTHEbO1w1Y/IJcQTJg+5YDV5vefVVU1MZDwPt2gjUY3j8e2BJaf
3ce1VcKs9i3co7PexlA+oLybtWl6qL+Gfu1vcnIU+OI51CVErVZ+TT1FTR6hdlHI
IbjMLpG9x9BMsqPfrB+9fNwZAB6YfiYYeLnaC2Oil1kr+vZUatkGmo3dVt5uG3I7
rxGmudGfeA9bLVi/WNlPs0+S/Hw1HY/s4vtSxKLFLDAHiZ2E+4jNk3UJ54K/GSVG
rb/bnMO9uccmsDizj1dfz+s0PmVUsGBbKGl9nyI2yd9KlFkXNHVOziWwVzJh24Wg
mL2HHIbzGF0rrllV5llSWZ3Mr/f9XfImZAyR/eLeAp2vI4qP5dHtBAcWBuP5JbJM
yN8YTdvvQtar0vVQ8AYJ/iAe6MMO/gqQSpu7bzwZKYDVwm9Hb3jXceE5Fw2N+gjR
T2fgQr/nxGwKSzaR1xMQpXb7+hi9KYXxLkZ0DnPdfMvupRZSdvX22yoI66FR6rUC
1LcoAEyUwWNYNx2GCaGLWuEvKW2SAfz6gk6sZVQ7ugDdOiCOZrBexo0b3u6NOs5I
/PkzpzBb3lBwmwGPCH0erjcVFkEoTPzQZomIPFG0t6p+I4chlXgfreXCjShlig0A
eeeFV08xX6Sv20Vqn9/aRCxukavWZdIsIUQ570pqKnetMFNRubqhXP70oA2ItHLi
8sp5nnBhBHkRBPqIYiIvYLzaL5H0hxBnDB1MwZxpBI2kz41piKyHc5AvjEdUdYvT
aDqjNPdwdmoAGNmvQDS5yb1ISaRWmWdfRnVjzhINI+veriNfnXUGPY3Xx2SuDqPC
kFVtE1ANurqNuBAGMSGkdCv9uJ/ggHjhlIac8+QIyTE8Z1wzVYRSnmkjnSf7ckYH
QpXzoff3w9HlQBSruzSmFP4hbuUw3/l+vd2Y5hT4b+L5gA+xd2ukwjj2UONNlyMD
RGRewBu2WV/+RcUzcyDbkVAE/BjImchKZdBEj5KCskAHV//QVC6Rwvv3N5OZ9iOl
eA5OFGmijj1bJRlykZbRptD9ie/HuZYWEYLh0ksrRu/m1+GgQ1zBTOicfwMf1R50
4j41La7BfDGAwXedbUdPNL5awhHnRF69ym3sRO3yvNAZe9ssNNdJE9yfxc70ebx2
dDTq+rKbX//ChVDQEZCB+J+m6G1a5dC2iJEbBfHV09N7iF6QV0QDjw3oTRgEy01z
KIFOg/B8/EuILX4N79wT5TOF6k+k4LsHMEqFA6+bQ75idCcswqZpu7nL/8N8Jey1
LChmbxQX2xXJ/wYZn80Ma4Twq+DDF9YjLOuUtgueptLlVfhxcqPDjOgZ2LxdZS6c
pWHVR3TRZg70hb5cXHjUS+gDi2PZb4K36IAchMvmZ71d3gO1TBbBLZzuonAcDvB+
F42rKP7ME4quaaPc3Q8ffuOQnx/+bhxSJiYGsuNxQpwpYNWub0xViEZMZgdSgt5E
nH0w2q4DpCypabtw/6ZbXBjTdlqK2sCeaVFmyZNUgETtCGfhVVH5jhn4GYoNJBzU
VT02beSD722GZ/bU8zbQj0boZnKCLoP7ASykmsWTEAxzGPbqKZ+4sx5g885qiCpd
BjMascRm4ShgrIXVVNGkBzrSaS+qobM2Eqm/9gCWwnVS+Q60EBDG2dadg91dnq90
pVOffjNdUFfBoKJk5eN/O2IWRZJsce++6/RYhthDuV+AtlsnR7l6uEuPjGNrv7YF
YIJjJ3INWBeWDnRhVaJtAS8Mtn+nL9gupbVmBv3+SBSsYvXIbdib+bbcNQkwZIDu
gCvqj2Ed486DuRotPtfp9pKIp2KXL8cS7PnPXp30V/do+agUVJhI6bRE2lULzpiF
qm593nJd+voCas2h9sbynO9CnbnqmwsxL0PnGQXR8yabKKn71mWvGFaIl6vOcgqR
pzKYZXlgKcIHCjMiUiWvP4DMUrgrVWFJEtFIHY4+aMr+vk6zd2/C9z+LfaJsKvXF
tXKihbJ9yk4vbPT4/dYPHi6UwodC7UcxnfkoeSNaKUNbwWI0MynEHLN+56gjGEWU
CttGRURSmowGs8L+zv5eZ5eQj6y1xqY4gpktd25F9Sd854KjTpAtOBkn/smSKjRW
Ge7nKP1V0Tg3dC+bL9RPGBAHR5CiCgaB6MFokWEhawIISCzRVkJefksuh8SKE/Rj
N8qtsauJnvk10pLEj6oEvW8gtR65KFE1dl9N6wKBRGUYLsohXmY0aBRwm2FF95pe
T+CXSpEHCTjXhKYZ0xROlgkyo5l4g03riYCq0jAH0fUxrjsAbaWJ8GoZsG7idzFN
6iQZAQW9/HPDPKQLpWC/6cbLSSLi/41YFmtKu8Ml1GVTUJNxzN2FN9FOZruiaPgC
nFVUIydlB2gLj0q60KRHAi1l+n6Y+0CLMlGnIzjBpHcr8E/nvwUzRze3Aa9VZ7mI
hI2X+MFA9NznX7Oe3+IraKKSKiiFYKNojLOlSkUqRGXHZSJZx7kNGmfLidIMKGXx
KmzZJ9EMlTjlqqcfTiQo1AprlnfOjbrqZHWzFQy+z9CaqAFWCbSnn4vh4dMjbFsr
glpz2g28oYNCvANjvXfP5xGqnRbYj4L54aa5oCxVGVETjKHqLV8i8+clqQ1P0Pvq
WCXwnQ8rqGBXF4inJTHrIag0Mm7OLl4+n+d+RoiwL/K2OeZd+N3/z/rJSePv27Yv
7LuPwryvL1edKk9PTtdkRiuEEAk2IkYHmN2A3VTYxH08NV7N2ivXj5ZZVI8ezB3W
WJd1zsBDtvNs80NO1X5Nqkd/XZUP5Nq4C68XtqNc4ixUIlre1/SPHNp41a9vXZE5
8IBMaslNEODGCgjd/fnyoQflY5wjY29Wh5xBI2tjhVm27xTrKXBskPQ5VvIdw1bR
umHFn0IdFk4WJI+FB3wlHteCp2k6g7jJb/GkdoGf5iCv8eScnTRbXKT+uK8/iK5X
IZy9eP2uOBuqK8FSxzIa9aYMnGZK4rC+6+7dgBbRChalMmhQAhg7C+LYAQHOc72v
cOVgwXIQsOza2eriwUTGQfUBFoDEzDDvhnH+4KFt6KZ4+gdsF/5Yhti7z0XPbNgl
LA6fw3DLVnH+LzN3HL9ZkZ2dmygvok7RppP/ZVWXrHHmgyiuNe8tas/QqYoq2x27
bQ7DNOxS0UUn4Rz4CIpKR69FvGjmbrBD5ikt7t+FqXcYtQckJnfgrp/0jewXLrV0
fd0hCCOvGIQ4ADICB6IP2c44VAZs+UTVM9trMK+THpRsnzWL82V9ix28D1pdYWQk
uglH+aecpqROkbKy5wLhVOeSkeYeCjH6ocUsn+MxNd8ZEn5NwMl5oiKbhFiawjaX
+O4Ix0pxeD/82h0rkdyaEW/m/XNW611OF456Gbk0LlgS0JcJEnXo/ijrWKn8Kz/G
AnckBh395+XMk0YtT34YtSMOryj/KuhNAJqmEyMuvS4igOjdypFnZjHiNpOSNcEY
xKub9s/jE4rYZCE7fDstjE/oiOiiWcdnmHo2xqFmrgYp7PyKVzmRxfKAaT4ARtjF
W9qERzBY1tRGhJyZ4wRsj3MG9XvV3Iq/LUq1LW2jh8enf2nuQ63PRYEF0hzxvHvo
kjFhNRflzSfTEkurydtXlo7X2Y1gmWKJvZexYIlfDLLTCjsQ/xEi2sSfDatOdB6l
cLhAVY1cZ0JZ5SCod+RPOnjXq85xGwegNuKqzO9KeJDv1N1pbQ61wgycHmLy/qUN
7Uxfa1v30h0odU3Nor6GMT5ORXYGlQQ8f9SoqUSn153btOB/vnqQHHAA423TnXzU
EyeBCBgLeNAH2q+1z8uqMbJUYpgy/JloMkAj3yNixQXdp6mY4t8iKhz7xJ3wObb8
EHUaMxp/jdLtOWDrGkPQpLSdb8GnWofnmDlcdY7H4IIM74Ew2sS1AdO3NhhK1IxD
Aiu5PpAPU1tHNzCcedYehEMRlOzPYvqXxGQ+BNL4+Qf+T5XGEkZqGcD5TTiKNB92
pqBUwZ3VXj3rCzJj7ZvMHPMbJy2UWUoXVNVnR5xh7xibxkuiM8AKC5OEMvl87XUX
MNragpglzynETXbOFMCoZJRuteP0RiAc3g8Vlyk4+RzAhq1B8NWMkLM9oh4bvhGv
2mEdxoXYv1SNn4MSQI08U1YkDcaLHERTELmTGTber+x45VofadF3OdBQm+MPQhNK
simI3MEAiCxdXSzP9wDREuLZFSaPvrwGcAT/9UclH8quYXLEKXbawGkHnUIZvSOY
ZJik/bNQJ8do9SYycs5qNBnF8by9dN4qQ4eb6Y8iE50oTHycPLvM4C41FT5GOMjr
4vzcD1IRCLyVPdsaYt4Ug6G+YCjyGKK9bxW9Bj1MziSgi7X37Tvr9vZm3/E9zB/s
X39sxRK5DqBj0eF4dvso2Jllf8l1xZfCvuT9Gsrx5bURPq9agh8On09vIViuwAVg
2Pr+/xSlkInIqMln/FYD35xHlJolN4X1Zby3r/yGKVCJX9AUX9yG6NF7qmv6iJ1x
sFhsyl/H1so6PiadcRls3VdSoGD3qHLiPfELSeN0CbW3b8b9H5L+MkSknXAD1QTy
WcXjYv/EBuVdKVTeacxo1N9qVpEi8+oRwMVT5Ny9GbJZ8hsnJHQElXC6e+KHHjf9
wr2aQ2/1sEPtuiGlXtgEWrVHWigtD2rSAzIIWKr4eZ2h3F50VpTmVdt99q8kapPp
dyFniBM2lsriISmJ1NKMd3PCH/iIYuz2o20EyizvaoO2A4/dunacSSZnis1VlL5P
BiHeKwp7mEO9I0WM8ZqjBGzlV1Bgzvzzn2YWQrLCJJTq2f4eKzmyPmunDzgv8Wwl
dz+LaSWy5ojvMXCxgIW1EV2iU2ALtoX8j2ALYzToyo8qH+EvxdIDQ6/ktafaeNdb
9PSQZeid9XWWQRHWhw4NK8kaCOgaW1xTkIcgfr+LRsWhJt4MH+20ecXzGKJbf0lh
7CWQB2GMVdLz87BEbSK4XlvIQpF6RDYSjMlhMvpbEJFzAccBBJEHunfN1q5Ui301
oCoG8NuJ94y06BUGDXXK3Op1l/sLXQoB818TFNmQpIl6yvXWIFKDesC8PiLcp1L/
gWlhLSi5PATME8MGzHw1mhlhKv0PG+r1t2ZoJsiFOTsJ9uPZzvU03cmx1sCt/bm3
zDPtpi+1dOqcoV1J0EiOohKP4/qnFmCopasAMNZGcPXGDbpOmtG2c40DwzcfypFE
y2QhyyoKcOjNJQqTeVQ4VEwJbYkbHHc9niiP5aTM6W37gCSLBY0xZHoeqNFIdOj4
327Gv9f12RLut+fgDWxG3WKYSO+iRNcjBvQ8j5rPUv+c0LMNBJvKKBRxm7DLPYh/
l2/0lwhYZk+Z/upkGE+f21p+45clRfZFOf17QBeRMN/9WHLSXRSUFJHe5G/6WYD6
kbdSDTCH9XvLNPeIEu/SMDkZRBHqHdYB54LrNKi+Kej7fDDwL2gs5WqZJaeiAXYU
6dUHn/vdZG7TDoaS3OBkh2fPYtXAglfDShu4W+iKKEihGP3UhAVwVnRwyB5OtiMm
kEw5s0K8+DcdZncJL5ekgGbsfLRKgO3OpPVR6JdtS8rgPvkPYWWEw8A+7lhpC1Qr
074Ze09UwHKoL0iv3I8hpeKmB5ywezTZu3Qh5brxz1/ec0oXCEpzz2bqhHFOX0RS
gHZepcLZRZ+JeRInq1wZzRSv12V1AvXLh6xPR5bQ55sy3Jnb2JMiLS9jztsFJ3qO
NAVDrG+ZymtnH7igvMFw8taY+8sMoz8i8iWIlCehOC9rFBXT7H1Fq2k6FPv+4wiJ
MBiOvUgYOkPNo8asrmaaFMQRYtCNybceuyUEvzhCloi4rFBVtpPsyMZiQEodkxBI
rp5OSJrkODJX54Toi5yGQNw5gr1jG1y7PsfBoR5d9VhePcgqLI4a8J1LtuLm13bQ
xFPMr4mGvaptGsZUURpcgG7D4pYlq7lFX3idnaLW5Ep0qlix3lmgB67VNcSmR6pI
YGRPbdMSnFxGd/I3ysrfR07G9MJexDIECnT+Eq3ftMhwXykT3FjyApHUrOazTT3o
o6x9OTOxdCOoB6AJVmFUJ+5OzNia8TTDKMVbjmDx/jBmP1wHu8YsqUowIEVNpDCV
pQpYDlFSd5BubXaaj9x5dXnJzLvnTYVxa9fgO7upxgcynrgAUtxTzyu4Taim7+rr
LjvOTqQBGjmS2HHDK8EurSS2uZNXMeCfA1o+CLePJ6pdaCrLz7NCfiSS+c5oL7G0
MjswMrcgg6BhBlz9dAEk874qpKBSXqwJeIhfx3JME5sACaZ76HX7EwDUpdZWLbLm
TPP2okSSrn43JdPIv3IeYRJktCFJsOWRuJtIRHamqQyKZvHqSYcnwpLCW2Cynwz7
xw+21Cw7RmLC5MJhcjCUipTXjpMhtvhi2tvWsGswLcV2X+iqd6mP3g+6LgR4ZLKk
PB5qwDd5uSI7gaGZNx6j4KknVq2CExqFwIo3mZjxhiRgOTqCLY1qPybPIE+2BGTo
uV/yHW6LkE45ywZNf9+6FY9fUAmwsFmAhBbEuGBSpvSm1/OPg2elMPtn2LbSy+gF
X5MucsekfZVfEH5G0qyNdawW/eiUlcvNqugvxBPV0+qmZzinIBCg/JRQxFgyV1V4
pPqcazbOHqszPvTot6/b6SjsVVLyvFExTvDGkXoK0cLfm6vDeCcvodNoUttTiN6k
Vimvk9OdbbqNfs/I1Muo7MK2T9DxekUJwB+7Pqsx6aslo0H+dHvladSz0TFDNRxB
2nOHIzC6wQcD2NFSI+1ou8ODBpmz2zuMw8+6tLYIyHRDt55f+0qzg4iscOmQY9D6
tkXzlD65tIdEONqBsG3grbuca+sNkdlVblOs6hJ81MiALeDYnj9LXFBQj5NEXe5e
nYJPrmMeyFDImv79qmV0s7z0MwSyoGUJKO3icnI7AvsLObMKCOf3ncqoDnLRlNfH
MG5YDW2n5cQRSRwakbWukM4ochD7N1eIrdfRqEJzsovWF3m8L0pMC+Xsw0sGR4Wj
c18qbX6kR0UTIJqhPdWs0Q2oDRwVGqvYzat7F/hBlQ62ybZ4JX5MH3uJFKd6QUb/
BAS1AesSfpgd1DGtbNR9zmsO2vXMCBLRprRH9z9ha8xhuIP3SFdZhyiAKNFQeowE
AuH1DJ/DPoi04JQGO5aepXCwFYWfic9yJyPq0zhIQZMQwQiNEaBMoI4PizPmLqYF
1MwOgOxyv1a1KBfTl8mVsdgIaAcC6u5mk5i4ecyy98Uf6Bu8vFEBD5rSjrYlEjHU
s+EsOULSSoAcvr+tn4N2QNMSoJIMCuGUTTKA4pkyJ9iyD2bNIo7qfRtyvlk99d75
NWTC+xMJh521Fyd9waRHeXvjWE330nrp0Zz0z4FG1Peyhhr/9lVZmAGc/cLlCK9t
9NdjlAwHJQrPYDQ9/0P6pCun5KTKMADyTpKeVkv9LVQVcI6TTnrOpOITyHCXnStQ
0BZV1KDNqMLg6q5aGMn8o1ovBYviVTUsPsxd4+UTheedhumcHjLNU+eVfMQm/qli
aTYjzOG33NZcro9TnrmFC0AwEhi4MDwabEBKC3vfq6AX4p/yjYjlRvuozVbdLh0L
vAp2pSFYXtXXYT+NBv+9DSvczA6GJeH7BoQLD/oeM6zOSbgxVIB2I7hGZADFT+dR
ERRghmHqE7OrSblJ7dhMCjxHfZodKHfePVlY3pDHDR72mE1S+a2bcOccQv5pPZwx
QXZOAAasn2AovMTXJ4EUbCQkNQ576Ykm8cm/fuJQbabgG8W/qf9Mf0ou/HSlLDBd
BFAPEAdGSHh9jWGmdQ6/hQb57MhWYKpGmidmSi/5jlKETGo+b/aFzSxo7+G5UXRP
B6IigPz23g3ZsuAifYms6OLRZbTbKefFQa/qePm4Ehhj6l4E1niCJ+gkEl4K3vDZ
MPyk/FgeDqwQ1g34dt7mFu1J4fy0pZiMvT8EfF6nKho/PAnnNS/fk7q8EHlpuI9e
D3MCVo8evbJlo2NnM7fnx9QUEfp1o4qYlJnIdH71HEcRWHhB026otjSIDrAF1Alf
fMstpF0JTg13X00yPX8pobhlfmDjJOd5MxQcENJm8enZV5LSMSVSoQLygTO0IJuG
ieDOCdVeNPktNsmm0PNH/0i50Wxw993RGrgmB0di4LmoSoE8VX1NdYrZt5zq7yWR
fNJs1Bxh4d2vth0CF1qJKrR36EFjRGhqE5HzdrQCHIiGfCt3Smp9DtzvthsOJ3mx
9/7zehp9mYfrdxFXGcvMZJCdLUfRJt3fakiqkBtQ8TCZSFx1V440sGcJfjnsxgKU
11/m+WShdp8uanHRW20PJFkKoK4pXqLg31HSJojy7Et9YHkcxDv5ZDnrD5Lqn6FR
RFAo2AbdmhV0uxHc15c8SGxKzrKSNo4UofCGxuuQzxZMW0N/xMBO0HORNJK1SNM/
0URIq9zGgREQo6vMC4l49Ztk3Htq0hjodnn/dvx4DPL5AQyFEFUBNrkxCZKV9Qof
VFke9VZSfBiV5zsE9aMtaKzqUc0wTPfEFybR4YdHk//893GGwt78ugJNwCRfAuOm
cDJlPA4RL8hnSq7/CcvvcOsqQFQIUypEqfGdikIC1LBgFdNxSQz2TC5LiGuIRoCI
qDLyIyNaLS7yaPy0yGmgutl9aHhsGcGC4Yu7CiBC1VGekOJwt2yU4byslj7wCKtI
m9Ri2XVDObieGAVtaNzm589CwOWaHLpKjpLtu+qJNwXWmNxxTfFhqknXjil4n18G
V64Sffkm9N+Fbq3bjiB7xpWcU8zdpy9prw172V7AxldsxMKgcTa9HV5P5A8JDCnC
d7ghIoKt93Cd/N1kCWT1BTOgxouwmpmNme2TUG++onuF1EmJotuWsDyfTbbwTc7V
D6JKZCuigbW+RN9uW/4WhYjxJKiVorQqYAbI3xlcf/D6B6n74555SHsZR/Upmynw
l5W7uotsJYXFGrPLl+2QfkOD+IwosUDen0+/yMdpLUcAisvra6D+STqmX78cZy/f
akiVNjBNlobt2MX92ID5hW/JjaoFlmFuwIxYx1Ybm2SAOIt/v8VOQyQWxKbG9Cn5
fg2ZkGxl07XvZd3QQb7urnetL83BLi/79EqSwIAU+QDO82uDhczI7wGW759s/A02
ammB9f7T674MvErIssbg9kCv+Uiu/Q3U7g973RJ4akiPV5Bk0xlgH5f1UmimnozS
eWfN+pQP0YsPVqoJ/e9dZocBsJWZm9FLggIdBSxdc15wYcMD02OycAi4kdGIur41
u+CP4qbJICoYBAl4G9ViwrrPur1PoWRkjx2uvpUFVzPjKwLJzlcORAmqYR4AgyMU
dKvVgK2HIh34wuIVlWsDllwjxzo/gue35NoBww/EbtWV58rfxFrkaClU+cCBjG2q
3W4jwMKoUiML1VkaT2k90uusH0smQ3JxNXvHVRCvZOVTI8pNBa4CTJto7XcyahLH
gfJL84lXYveFb5FTPDmttFyn07v64PCtJUR4OMhcySUYeYJsC6t/LOIilWczHoUK
OjU889lOGlmYEDwVuSjZ5DMEpvYXmil1D0T3MStK+mdeT2FNBwTaP+1mM0rz69mr
/BnXzLQSjr1KV9n5Dgg0zScFdvZjovTMJGugXCFb7bDKpnNKYc4zUHe+Wgiao5S4
AmDDMQ2dKuxyvmrDn2BDnbU9oGQnw/Hq9+0N8g5R6OY6IQx3Xoa1kY3RYnnOclT+
FTCh7pHMY1nR279No/IZk4jZgWSDhwrU0LXQan1f/8c/IIi1f6iSsl1ZgZxQp2ig
U7mbKfhlXT4o/nOpsiDHoMBJuUqPcpPmnHE4TRm/At7iYKrfREygQq6EJ9r0JHiz
FvyAVdRp22mhDzM/Ns1JQQMLHc1QDgIY5vFbfJ0SybX6AWlUliHbIyBElFs/i4v7
0FYfjxPyLG0FXOPWSt5JOO3AKw5XupRS7ERpWYexLV7JTztqC1kyYQ7u1aQ2G7CY
+Omosv2OnHMpSWSFs1ev+/nf1JyDos3s6yndVGZhR5I3sGBWqKZj/olR9cZUsLKA
MvD4rzP0AS7BKcnEVD6tjZZHK1Quc2dBBGmSlmi1dj0W8l+g73NyCZDwj7bxarka
/f1082PM7C9vmur9OMoHUv4q0PhMifsmtPHDmsyZtnpGwobO1NHm2cqfnFZWFdu0
DNFnTn9hOdTa5mt6kUDD7wgLkreKjztC72LZiHunw4806D4j5NRgchXjdyvijkZ2
xF7pK4IvgIKv9FpnWRFXBH68NhSG0Ymh7zdfmeZ0e6YFJjoDO6R/MRy3P89mfpkx
nqWquLPWfqmlcQneBuaNZygk/tVgeavohCvkv/pFup64i/0u5dY0HJmjUXSJoCY6
aOSPQZF6bRjUuWfA5H0Wn/e1o+4BXI8/soB/+3I0y/8teMpD2yVuCQkz6HaHi1zp
YfNuvCxQBK7IfR/JaTxiknAuwBDHH/PjtNwx6rXNgRSvAPCtylPtcsjqz5Bsa28+
3hoX5ZRKPH6LzMxFytpvqRNkcRN4qwqYb1cqb/m6P6G6cScPG4xuovAPnp+Op5vx
EffzxfAGTTzOFSLprFZij3g4xJ9jBXCIaRhSQMQFtU9fTq0VNgGEqNE5Dq17T+0F
FuAW7CpEqwTHD8PkTbbwJHYyaE3b1dqUwbYeTNss/iLIbJtqkXHlywUgokoJlnHu
pq2fg1FC+wzH9teAItNv+d2uZFoQHbKu9xvDzuw1s2mDJQLYuLeiaoiFYr12/xOi
MEbt1iye7TVTWvmDhnXBCWV9214Jd+WKcY9eRigD/gANK2xCrzjv8BLqKGluOOij
MzEaoOOniekW7qPatOkSz9seFfS/o0Xd75Ue5XICO3uYrvM2VomUG4Xf2DZJN6DW
1v7rDacLWWrmFK9Y4BceLxqJU60+JgVkFWYj5uXAmyJkMrM/XiLLuFUhjOOs1I9W
coXegtfThDcL0lQLo0SiimixySVEH1d9uWXFJHPaC+jgeG+HALgGi/xD3e9vkR2n
ncnuu5pIzZQq2the8L1nhW7ZTmTv47sOY7yJeUt/rKEexiJX1hvwn2jLu6DjaCnV
LCGx3DdThzt0feika+N/Rd5M4q0Lkxd9IjR9gf+2sj7+IKrSE9PqJ1onruvAT4i3
i8PyWjlg8cFz6HDMzBGv2uSGHkGH7bJv3GAOema4jOf7OLDaE/Q6Z1toMupczySC
KKjYpl7oYJq7oSaXyRMFO5Z685usEj++aYkmtKHtTWxJMepISN/EuWGBfW+es+ap
4NRxAI/QoYBVCh11Jq0cpYMUJbDz+OBJeFuIYqv/moK/jk0k/H64cwVtZ3Uvzepk
/1fuRCM03S3zw+x/k7BF7ws69SBwo7syyI0CKzkLjFkEVEbKVFPgh9cpkl7XAHMK
6nKu1IcLzoGr1jIzVNtegAPjMMwRTROu9KaEl2HZUpdvg/X1ERo3as97AguW89yU
SzEnEbbXbtX15WMBw8B8lpO+bzaRM4pOBpwUfC2JVwGbxbBF7e1XcZvkAWSv8jHx
hebzeqEsSkvqnU1uGZ+mxFhNUXLfrFDxZjK5TrL3+D2Jec/WXAGjYF6EEfFwYGZl
LmXtXgARWnCeclFSeEa+eQ7YT9Ne4eXjU/FpM5NLEJBYt9JNLo01/hELWdwCEb07
urGTogdDLQyTxfaXN2+XzfhVFZxLbUt00SZI/eOC0T5u4gtfVbjVr5B9UIUW1bgq
LhPNksYCrfNUPwOEH+jWFs2LpCrP2WdG7r5bp5dEYHt+hDvah5AKvQXea4QiDXMV
tS185XTRYk9jtzu8/xaLUkcXUUvMzOKyXSWa68ibeD6ou/YzRJgutK+h/jNlfGHw
vevnXMpfzzFB5aLqUQMtdnT1rodG0tATUHCZRpPBdWkhE7EzE86jy/wvGMMG3Zj9
7U3AgOke22fZurYMpH7yxLE33x+Rx/xLqdEAfSu0cOZdfhhNCpCcslzAyvlYq0tY
tzuRaN2wGD+Hi7KGuMS1o33SO9heM6EIDFzg/CXtJfhSZF3X/XzEsrbQ0PanK3lE
ibdSiYdKkwf0g3Bqs8PlUehqUfvyo95W/HQ/HWIsI1akpoTnaAJnCCfX4Bivkkj9
bYxAJKvMhRcqvdW7Oeh6OPGfgpssBI5cx+/aBjBGl+dNy2oJOU0aEYtdbzUJHS0+
TuASstsq15PnwfN8bsoN8KWQM3tDo6WcHLC8b4GSC4p9FgLBKmB7VnTqe9IIw4bZ
u8UE4IJFi9WVoh2WEr7qpoRveGpDjAWPWalIBaNbo/dFTvdh7eoWeEGcjCAUE+RK
N04Cnu6PqzP0JU4MRXGRDbat/76YIQxgDNLGjjfRS1FoDslJQTbwC9603S66x1LC
gfqrII0/7o7pjg7TNHE7CAlkGjGlj0G0Tkl9cyzkxNjDWxMWfcQ8Iw926unBMuUE
q0qr0z2BxoigzNhYjBFYY7/wwC5WXHzX208O7VYCW1/IuQ+b5OfSGj7q0hIgo4Lz
js7vQO+jAslVhvXp8tRm1aelQNyR67v9MILu8/OYggK5wASEdSzcu6ZiEvwtYTMn
5s+31JmwCpLhFvj/2K5fdDVVkDZATqPI6M+7deBc3GJlAYqAZh+QIZMzCZpZN+3f
WIyPEZ4TlAAbKu/uiNMbKQ2FZffWX0GcFzxoat9mvNbTrj1cnkqF3IKE0nM2zAte
6ZrwY5GMUiiHJhLYl/TD1btKNOFLoeqEi5i53wPlR/mUAdk8bBEBbOcwFd/Pps0K
QHU5Bu5c+WjK8fRIsp/bwee3lBSiE/Hh3DEj17WxNN4dnxDiTPUa+J0L81QY5Tjv
v41lCzN5ZRSg/HdS8P0gz/ItJJROulHlalHL/euo5MffVeOtNPUckE24c3HvU8Kh
9H8QDleek0fYSqq3+FPaZU78IPQTaM/StDnTCyhtxD1auTleEmOxJeLpeig30RoO
8NzvyGqo4gfbzMqN7uVWJy/1hqZVZfHVvhXgDgY96df637KvZx9rNbCKa5yIZGI/
JCqUMx+YTcrbuYL/1W76/AZfek4UfDkz48YJGjuWiqSp3CVz2ShiDqJdyvTmFmms
vYLnXYlsSh/KP96W/Lwb6HgWZJXNPgpz4PuI4YPvkeoYHCTCuO6R1FFDtCe/7LiC
m4frxCqFc4ubTebvgGhlb7VLZf8JhwwJwt9XQ3I6I/oOkOq5Fs9OKlG9PJp0ANYd
nnLRgjLMf4OAPRYDCIJk7ySda53j+C3aEMBvYrnZgWYdyFpW5EhTNYiexJAk6WAE
LS3XNBBk38Fwibv8Z2uEy/PpUIn+i4l1koJF9Lkz8x+6KJpaT97HmBdy+wHCEq1X
IOIOLNb3yCXL5JMYZBGnUl8EbGRkFBnLvI2WQ3/vsvfQAivUtn5BBzW0ShAT+kRU
7qqSaQROrtx8XeJj3IZz5S6Qzax3H4NZRKFA3rplKERhyY+ruFnmXVzL4anEF+fo
Ao3rSdF5nDQeukAjBhoytJA/AArNLzpbOPsU53hc3lcc6IpU+IZukZQ7Qr6L0Q7Y
iv/iGpFEe6/Xu3kiWRB0KB/tflnc7nANpPRcc9yji3fHPViUj6FC6sxXbO6/BAwQ
ZocihxuQwKDkYCg0BTS8S3rCpVJTttAHQYLC5SuCLPJSwM+IsDV03WaEUzy4o616
K78ei856cP86O02DPZqzjVbeQXWSTJLI7d8OqAZII7sSWOqkJVaTgJfWi9fG/HZc
Eb1xNdwsuftCa0BnqIxhRyFjEhJGPvoGE/7y8mhHX64k8+MIwwPAcl96DuTs+Dls
I//WGMVjPErsCbL+u9e0c/cyU9JtCMWVYXxRK30kIOLFV3drCCOrXr73oRcdXlca
56cUJBw7+mR13IeUrSlbvsiNcF3X1idkNrMFHJDm+I/vezz4cgrhV/Lqj+ZuqUrS
1/HmE7MOF61EEjCH272yed5PGeCwEuOm77p6ml9OofzfaZF8t42CwsLBYsrSPvA2
S227giXVpjHOSxcwrz5yj3ILuLkeaFebjG3Hs9TH6esRUHw4g8Z5SfmV4bRu1dv3
A5o3lOlZiztU69PF9/D6nA1mIu2MWl7iZAgH7xj9d4dr9zaH+rVx11mgGoQkdBRS
cIT7WzUq/uinzrEDOgZNa6/+U6PJ59hdlkk1dOUpAUJi0uvlG/dCpSgsOWUAOroJ
gxE/eZic11WI4ypYgrjY4UHkpVnF1ScfdvB7eq4Kd++se4bkYfdmguvyc1F+H//1
m7yNDmna+fxMye4oI2MjQTWbSRdiV1H3X1ijgf4x32C5aok2wN+zu8F0LQZGN9RC
HYo2s2bzB0tCsQTAwm+SuSA01joyypSkfNC55Na/GI3lfMbIkfGnFp6s6u+ceKgU
bD/Gh7ZzGlWJuosl6xLV78L/XuqdEhBtlG5c1rkcUKc6g+Xs0dckELKMRfm5E5as
r93WWTXbahf9z7VsHpr5XHJastQ87Qc7+nX/3Urg3EgZivq5WrUlmWpxyK5usIxb
Y8JdRcvM+2Xed+u3XQ2Pmd1yCLnLviTW0Rj9CLujOCNbIZwL5T43j6CwgRmYPWfc
QD359FR1D3fObkbhvoieJhOqvA2LGsXDNjfBbT9s/aF54OAakeS2ZnCpMq68NvH4
nQKN+LB//oRlOoggSGxc+GuC7Z1cWtSgzzbc29p1DdSVJde/Qk+YQFDPnAIzq6AS
whgZBAKPTSWG3b6dzjn8j026foN5pxH4yGbB7sFGwkE8wSo+6wViXzJTEjslq4MO
3o49sKmooFhoHaFDS5B+KR4QtpzDp6Ye5LNyuLSC6TKqGTNVsidXDHMqLm0pOpH6
YZLRLMgTVyQoAio4HlzfQNttgnK8rmg+K90IgxvnEs+NOktF7AIAXzDD2PwlnwWm
aMKpRTm/vSkuWgP32NcsguDXIyW1aDTX0cKz1CsUbTJskH9TIXVam+1n6wFi5xdO
hvV/zBMpUpzwU55F7gnEwHg5JKrIeq/6XFx83/h4IJQEad82mqHuEgh39fTcP7lB
6d15hAaWytEMSz9uV4NJlinnt7Qc0cLXkAFUUMf0NstCwafG2xhepv3mx5fVg7qc
CyfpEfmJzSqhhassUOkeVJslwpQ3QGm1UqwI7HUkyXJQHWuBbv3vVHv0vbHCexIV
qVVcXMflHjArBuTp/mBpmj4whoucF/tq9A7irpa3tZUGU2FSQaNayfK+6Fk8cK3c
4YUpBAowlJIuwotIZZyF0CHjQwnxBCctBEluKE9R9tUpMwIaX0X9veNA1QgIcFdP
38XGTj1X4lwSP7wLPZwxlwLdmDFD5D6D+R1aj6oQ4sIMUjqrmsYBqvIDrykCZLKU
im9jBv5twIO/lH4zbO4OEwFDaOwWNOEMi80fL0/kXilQxTDeW+HE3gGR+E9iDR6n
a+FTCKPsEWpHLZU08ymitGHGzF7C06zt4RfhzkEZV7qXxP2RsYu4ufISQTkaKOno
fNVKVVm+0jCcXeTDrK+X49qNzvuHO0hv1Rs/r2HvntPQVXect21p1tkf1otqgtes
DWb+akliLP75JOMLo/edKX9WREHSdBptsvOU09VT1nl1UvrHHHIAlNCqOCiNwq01
gsh0ifygWVJoNW1fJ/qffzjw9HB0Dclz/XdWwbSPX/lFYTaQ0dW5FwGk+87so0rr
27qpiy3gWEyXE9w8XlmjO89nlIkTtR8Y8B3sFNJS6OkmmlSIbx80c/Lee2+m9Qe3
M34MqK9KxZvoxUI1mGi5A5cp7s2EwKd3Zdbdxknn15bdyejJHBxRni3zXAE8Y69A
XEvHzQwzIww/JeukbmoQwZ5QbjF8bFF8WRCElT80GtONOFWHIqBXzL7ONrXLwwHV
K0BNJ0CXsH0/69BE9OORDLzVZqh5U+PV5HTejIVCkQYBNKz884qEUogRQ0V8Na8d
WTCW11e7KDMUg7C1MjCZIKL2XzQZ0ko86WGCO+Yftvx+ctuK3AOCtkQL8sSkjX23
6ENn56+Rk/NWHrMjQcHGjV2TnILgMelMeRoZGP/u8VYuwwBLwBj9il8sqCf4gMjN
ZbSCjLWRyohAE3rI+g/oP6n8LvtfE/oN8OQobPE/CbNi3sXc9hI7OgUkntnh5NML
iMjV+hphEddZkc9C58Etq/RMSRD0H1qGJ6JEC7MlEw2dXTfy5K0qiC+aBMjuaIvO
5VDHroeVnvsJ61gbeP/9SqpvW9gF8vhUjSHgcQU6cPkoey1NdIvaptjua6PKdIFq
xn46kcCizqZuv2Y32ot+LcjC16RLLJUisvQi5zK/Dbx36OCfFHjjbAn5UGMWbBsc
NjQBqeZQWgJV2JXHVsiyYieOX3cicU/rGgPtdUWl4GKXxQArprj1xcqWECQL62nM
tALlFWNcQTjwo1aHctABaTBXAqEgdd06JJJ8FylePaT13VqTUnSPex+tkklLFTKp
ABHuj5nJ+TpD4jpa8bhuMn1yqJjreeR3pEJYNNIfvdYwQWeFbQB3sj25kj9octDK
sNEmR6WROCKCQva1Di754DXsTBlHtJ/AF5EmttyUsAVtKTDy34p8jZ5jzOTQJlSP
30BUmUXAi2nKnAeBR8WfJx6PxE2n5BAg1nnjQN//nnbpySsKkZICo4BSaYoMmoXg
2WL+EIKDo1dEDUNBL8+Mj19r7e9dyqo30pbZWXQO4jmpe9sWBvagePiqhuU6FGHj
+zG526yuEykU0FWpbzkC2wcFn1EMFn0zSEB6VkldW9hL2b5+lpf1V/Pu5B6MpVOs
xzPrBGmbXHwi2PKpfzySy2luVrD0MDU6tG32X8DEzxv5eCoQZa+K89jHXKjQjZvo
PIrphR9fd0DmyE+VKDlCF/tcHuKUPXCF+Mm5KIZSmUSyT91EjhEGcCQnqTmucQzX
QrpXO+kJcZtg0UOQ+jJdW3zj6YufS/WaE3YAmlDfqRHCyTTxg0ZlClJlhGKfD+ue
GsUmMYno4sTBQoqB2XprmrbS601mr5ngtDsgN0ia4U0FcazXGycTsbyPHsiQ0tnT
NrJNOXa3zbT9GoaHVLz14O7Vm7B/68zvC3iThcW31xky9+MAeeFZXuaH75FRw4CO
WT27Bz1Vd0vPu6p9Lt4v2ty+OqtIPo1970SlcNXXqtid5W5+4avAZqE4ExlfoZtT
Jq2pCelGV2oUMijV1Wohj0SVkNrLHTvUz3qPSEUUXzyR/CQK1gQ8lydRUUNQ92SO
v4K34ANcFNX4N4hQ5liREHPgXh/iBm+6xHfN9IA/MnERl3cAmAlwjKRom2UzNm/x
z7Dn+YAVc/6lve8UlM3OEwNDIMQ2QCcfc8NZOv7FTb6GY/bZl06PAo62Ea5UkVjJ
ZEgjo2RakI5pT1ooEDC5oE1NlWrSv3w/1qKBkORg4ZDK1/qQG/9BM9jweMD0MVY8
c78xHTrLUD4BKl4FgJpsW9+w2s+VnDIPw/wT4Bjxbg8wyh361CL1XMTo9qGFs48C
ABDPC92zqFjTToYa5do6mczxmREIETyrRhE08mtHLxjJjjaVqHKWdsKwNbWbpXPy
N/HRmypFc3ygeCFbLvOf3ZF9uZP4CjrrlXDWWRXUKq4Wrf1JcJFSbWO/H8YOU1uF
Vt6UICDUe4kVFRSHvgSZw4QmIGn8fpFwGiTZ5J/X5psM770zysQoxOxam4J/NmcS
V/vK6YTqwzl/7NBF0oFirjo7ItNgmBE5cRRrZU+IuMTtw6KMuEsvpqHt9qKoS691
e8eVO7Net6NrypuSWhTowgK95F54n/oHDmDpUF+FulpgRN75htBWUpsaUZhxl8x+
/LLNTJNg5FHBgDl3kM99Qrc+l/P4qhtg7I1kyf6B3zIcWZHUQJ/XfydJ9xGgHc7k
8nmvVRvbuP71RlAbGROmY6D7pp2sPmNXDNetAfS5fmOCIjnHNNLQlts8pmQwScBD
QyrtTc22Cg2z0nSMCQ0QLV7AxeZMEpTK8q38JFYIGlPazV1hDNaMaN6WLIVKrqAR
LiXYtUnaGBBhe+kIvc7J5+IRYWjlJCun994RpWnXaIgXKY/YhYPp5tgK+o7Krti+
MshWaj4cc9InC0HwuLTkVBVd2TGtIHN0rDWuvceTVCigbpfYiQ5B6z/sNquooDqC
kerlJarR5/c8RBAinNbSUOSiZmxeLSYD9AFlHyxI10qFl4eBLnLx4tlBo+oFtUAp
sODiQztgMFFkUhF8nnLQxIYlQDNDjhhUjC8Z/kdBFhpjxwlPSij6+K28SJ0fpeci
rizUKl1gQyqMdikajv7ZKtmJLBE0HZRsfMwdEwfrGg3IQXc+WY3IST/Nac1bPh0I
mVrfcARtFEqUdQ+kLxLuo6fgQMye/hPQPlziDowseDZ2jphYIDdjLXaqiQ64BzOv
q2E90yrHs0nO/CEKfqJlbCmHfxAKJV5Da8oRqSVGUBR1ogs0aX4RM4y41wg8aFxY
Y3Wk7sYP7HtC/JELtnaa1OexGTfXMrdAYA6KFaXGtgnEoyc7hyOeCpE+YJH59EVk
spdDJrok5EqwTTzY4oYiZKeTgLcUEkhr1Rq3uflx87pLNwDPzRPkBXOFE6S1rZUO
1LllGR3m8fqRzxT0pRcGbCswlN/phqfBJ6kzLMpxZ6ZYifqIb1GlygKkxrhZMO39
Xg0XGbG7FViYZO1IwP06ONEWq59eSii9LhsmFBph/8t7aPDlc4btbydLdooOwqCT
Q+Vnojhs6NUwyGyRzlyJ7gdQoGaHFGp3d/faq9ya/wO+FRKzi3lrZAqbut7cur5b
vB5Fdcw4DDVU/gJCheaC5qcKaiicodAUG1kB0eGdUb6+B5yZGRILGPIJUy0Sth9c
a+mfI4rv0gvYi4C5Vn86ELLo5Y2ci22S5HUC3ShY5TOhOQC+hhgAXza01rdSf91G
Pu90T41QK7RXPfO+b2TN6RFdukGRBUJZmR27Keku9iCeizRqZElB9EBrStfABNRH
Wkvrrn4Hw/w4viqAvzvifN6KInPNEM5aiA7VWz9sc2+HFFNrmWUz7k4RUEyZRHND
0rUmevPP/phPDy3iqyNXn3IfSrbMFFe24W1SgFG7wAu097utFNFd4OIarRnSQTxF
Gs1P6y4yo+Z5Lt5e4imMuDBUfi+3uO5lg8fEu04AQdYjv6UxzT0I3fz6UNK6LN06
jBDCM7IXnzZPJVeLt54Y2vIHAEW8Stwp6pbWvKRD24SWE7tNqXZ6oBxVXqe3eyB5
MO54ijkNL8LqyCRODsz5YXZtyuoOUh/8cgchkfauQ/1R/QhE2FHP6kvMsmBEX0Bg
qTpY4QxgIVGE1ldMvT18a6PA19ZaQLcjMSyHgOidSyrzjDL++CqxI5lce9rlcInb
XBdeRm0JJ78uv6GR19bYZesBrFPzTqnCC/dKCtg9eJFv4ofb/sxlgrGDdhS+3XBt
tAkbxomSSulkSwmDXyhVMwDvhjI0eliopbR4rBA4N9u/tZVPhuUH5udukQ8TgM+L
geJB1ii4VLAHi7WjYOKwlT5wPRNnQRXopOS1020DFTd5FHkmqYNH/5BJ9j/5TrhY
Gw2+1otkLCmyiig0pmilC8uuXBK2kjEhxbI7E+nRezQxlhLfElCrrkxGnI53g7e4
Ut2jaQqQiD3YZbvfhvYvpFButjtwTKv5dBG9vUDUbutSCt9EucSspUvuRWSzxrSP
tmL0DHVyS4akxaFBFxHlElDhIgm5kyIOkn0diNY5o/icinRzHXtpFo8sVw5VVk1G
u+ZAq42fSQgYM5nxHMMnH+snCpfvxPPtRuGs7JLKpzUaCr04ozdlpT0sqBr2yvZ8
PlrdgrctwR0X8/dPEvI5w+3fWTO5PkaaIoBcEj64POi1yssRIoqt0r3oLeei7ces
R5i/9npE10tOuqrwGoCV2rBJuYHiYSOuvU3Al+xyP2robRirQYVQ/8/nCnOv7vtK
gK2G24jOiIws5Qy+Ic+ozMrur5Jjsu+Ha9qOz4CTGfh+EgIndWK4D82gwD5bffcr
2ct7YbHfK5c3vV7q5MICZrL8aOfSabvel2JxKlOTxn7mz883E68bX3b20sUMEmIy
/rk55Cfp1T6rxxwYf8D7of37ZAHRzFFet5VY415SUEHTq63Dec6duo24OPUHGm1P
N728RhiGdGbJZjrFtzSNGrTnlUSa8NPKH8lpiX/oeatwM1ETfQ7SVLvO0CxYEXrn
z+lulps2Vzpi75ymEMdZr1aONj7thYMyAaAoauyVkVCpEzThN1t1+3Clgatj6s92
NMw3FbPWp1mP0c67/gSBNRK7QIVAzdU15aAbo7b0qPl2ABpSW7MGU2X+OOVWoaKK
ydy4IezigBLG9MhpwhG5Y15ClTzxdYSuDo11El5Y875sNkZgWJAfEBasedh5EdrB
CEniHGv5QpSxIAhS6p3QbfqSVQ4cxgDWN75FfF8QDBG0uCcBSqteiOzI5UrpH5ix
6LjA6T2Jvtpjbp5pYkCmici36GCaufYTD32qRYAAi6X7AshY6i/68qMyN3zR8z32
vgL3mvutli8fEZV4zbEAj2hQjNWPk7eAKIPq/lXSy0ogE/5WrzoCn8319AdiPZVe
ECuwPgjry+76EN58ioMGHJ2Dnasw6hKgUYfUPsVQ4QJBVPw6LpsGsMRDk9aeDhLV
SbvdfS6xusCvKCru4MSThGsGQQktRv0OcWEikv5jCXB3E3ci96qvlszgV/b7DYOp
Ta/pbyVbyRtBTF5g+Ii4vNDX1wV3ats0grT5rHPqCN2bVSr/fVzkzvch8t51ztIz
DtxtecXgleOLjZYaKSAkYvHSDToeZTKuJ38kuWkF8JPFxgIFGaL7VEVQ4e/KAKUB
xQ7OGl0b/vrB80UNAbq8akefSMHc2YN0XMx50rd+JxZgIrr6plaN+UyBZXSZAVJu
9Ge7sQfcOTVu9vxc62IpQeq+IYoEQ8pc06Mq3lpZ0WExIib7N90oESubV/TANb2i
sEZnwupPkTdmMABafUGzoSBBTt0+r5xmTAbJ//M3tl1n98ozfovuZjkr5pKXMG0n
3w2aYdHNkyd0ffezNT9T2Rrzqc/oe43Qod3/K1Ko+Ymea3woLMhBB6wYGu9ChrLV
NDKC2himS0GHWRXBBnKDlOf2c4rfWzIbnnigqJ0wkdV1egMKAeQQtg1Usvo8K1hG
dWx8y8JAPNmNzFDJL876RlFPyjvWZLpgvTMHEGmAu3iuGzzQhKTPe6qgWubxYrOR
Wl6/g5JMuHKotZLsVN9knlmDb3h7Ky12QMiUiht/vpXwyDav4TFQPczCRYEP/gXG
nRrC1SElEovZwhP052idppGgxkCmcoVRGVfX1LFno4KkAgMkOPCOuZ8x0iiNULAS
DuF/7cEq3xvGnPEN/0DXWxLcCfy0SDn2VBomydHSz95A5qYP/A77vHzeqGhijdUZ
0NIwiR95O+hrX6y4cJ00nbZoQ/xDyJLt3slgSsEo1E0EJYf5KJmtolQy0t2tiNAz
Vdfr+zbtECaaoOPjEJxj+bW+FgP//GlkBwZwYTWdD2vg2eHAMxqgF7qLODrY/O+y
VzkECsf1zc64qE12Zp0otB0hUhlI+alhQM+AQoAmnujjqFWJsd7RZQbVmoP5v5Pa
twJN5iT89g+YzVX6kYGpWKjokw2wFrDhXDKqDiQqbQsP5MLawseu726398pGGOBe
vQOWHhGu97r/9sbS1B2yrIcSmbdgESKo0Em6Z9oNsp2wr5lkqrmHjOFV/97q7iO3
9UJKBbeeRO8ZrMCTQ2tQ0Lrer3c+BHnJ4lPAatxet3TmRrV3YE2V3P82EYtoE5g2
GX/pRvofRae18ohk4yqjtk/nmXQ7rjwCRenH2LqNx9TZu2QcsznRtkYoM6b/MGjR
prORd9IRU9iA0K2B4eeXbjUXt9KiGDyJbfeEv8tCg6GTgEjyKOC8CcooHeQdx8jF
mtPRy6CXd6l98xaQdr+ShnCBS3gtXdbaEVXCz2Jwvb3lABas1gOSUxipSrX21f1H
zf0p0Bf7X9711ji/mVhH7sIPwCUfzeuVcfdeHPD2hFILUEb5N9EqmXTwdnTOd7bn
riNkd+bO2KvGPlBtH3KuALdxxls8XTms4rSIeL1KtwT3PB7UZJvzyAz8N9NNMNUR
WUmLt304krdd+gFf6Ip4oUiHMWxEhonTrXp6NQi/ovcNAI8+UP7AsV6DSAsER1Cg
VlTcBg8H2WufgZZd7rNgLIZYQLnZhlkXbQawH72CSanLyyLJCefGZNNDvjrM7V/u
t1Pb3XWQJ5nm5oa2Io8fiRUyBOmbQ6nl9C7WWNCeV+sYDNO8+Fxu9lChUV5bamww
EumR8AEVJGg08N12+qRyuPgoBOFdV+fP+xxfyBUWEL+V90ELE9xHTFNXDtPCGp+Q
X8N0SZgxyax1Z2RRHCKlbQqmEshKGf7A6HP0IuNjAbWeppGWnXawj5j5gbkK431x
Hd4+7GcocsORapJsKR/ZbHAu0/Yk83X8xbiiwXHvcH/hjo/xRbmMhwLV+8sa+sG9
4XWSPUEVTdfSUf8mOkcONrWUspV96wcUTUnzNbUiUtzdK2MKE1ft9uV2/x81aKe5
0Z1f+PqsdsIGY2XirS1uVB8t3xygGu01cY/iLTicjqtxDKlJAL0fdKLhoJ00ourf
aoIFCixtWIHABULu6PfRxG//8LhbSC82YuqsBxWFzdTDRrPRGguiTZ8opA/Hv6dW
aJgfiuD3QmdbbN2EmFvCm+LRI9DUEfnwXYw9fnEte03Ek9Fk628AZEQFIaHtVznt
aoOpLV4wbFlMwoa7g6oOxfZdV6SJkFDIgPWF2vlQNlw6X9iI9058WsI0VVGRNSjb
qatGz8YdEuCwp0LuPKe8wvWi2kLe9SvdIaB+KjsDA+45b70FipU0tjTxwPjQ/8OA
lHUPO0aAzq9qEC+ShK3Rx33b9dua++VzZA910J/slBTqfGbyS0xtP9O6mg7VOGEq
cRl6DHNa24+eRPNK1lDS1x8H0fWMfsqiE66yat5iajrH/d1xA5XDzaYhnOi1Q+n9
gzjN5+YqRtwo5VK7XrAT4P5ICZYEZb7vFHOWojca43LeR6M2kQzaZK3Txu7SUBe7
iE36Zhb7vBL6G82H5EQSd+iZovxjXAQdky2/SiZVkRVp6nQ6DwPCKKwFNNwoXd+L
Uj1fT+WJvjxQR5erM5HluBZHmOoBajV/pb/GZ19wNjgXworecfZ11UXZkb9TIpNK
47nid9osi8pF3KFpTEuSHIUQSaL2Vk0yV2rJ+CLWtR8vxlUd40nRtgM4psPXWv43
Iky6ONaTq4gysGmEbDNWC4xj6eHac+eYylHdpDYt/WOvu+FOwW/mdlkDFwsa00nE
HI/2uX6knwpJPUg1QCoYqdhGnFYn98/x5/kBSXwG/MuHCuXUY9GeLxl72PXnxa7o
d7sLjW65nmYsrO6u8Aub/mCaEpNor9XiAMkqUa7Ggbdx2ftO2yGLUs7V1cwbDyMD
ctI8xYXTAArWjpGegcdCleArweg6NiIbuZnDE1we5Ox4BOjE3VKs1u+huY6z8dty
JPql/t+pv+NwIfF2pD2bwi0QBD5NK4qvRuj3tvM3Tpy3xnrSiGZ1Z/pJFNO2CLeL
mpcwKHBx8szutGk3QXDngQdqGr8NeOw+ug1L1YtcFDph2v3TAKaTG6Ad14SlyIGv
fbze6zUJ97RuywDMdh8cfrEhReMnpiJ0COE9zYoMHEeICMBpSYcfiIxunOZiYIEi
OZ9AD+73g90TvrUXGHbIsr4XxOJM3IsibMZ05nuGF1QEaJ6tTAbwVENBNbxZgUxg
lqxYoq1FksD2R+hQG3166BEH4ejgNH+4VUzcs+mrxBdCjAQkMyG8uLQvuCJGPdxx
BO71gSsG/oAsrkkFj9bnPA/4NWQV5N3TMMUidbOpTuK6THEKLFYbFgqVVBnU2Kxp
ugxH4METHS9Fvv48mbzDVWLgS+QJYr6E597oGU37qecGeGyu+aXJaVzMbCfttu/r
paDo7Ecj36KW3ayfe/eT0pCMmYZU5A8CeiUcYuR5K3PkpfwWhtqlSndsJGRlQkFH
uu2KGpg46+YXSZx4z9i3c0cu1eUcWgZ6UqQy5b13DB4NruPxN39xSly1HStTJVKJ
hztumGxAuoMl12/FJeXUDRnKqbqPd7LF/WPcYTEl1q4c46peMWUUDQE/FJCgC6Qs
6kdC9ahjf73voBl9QrE5SX6R36EC0bjFErjo3IxX6HWVdPxNgdVy1oAgqoWPU8wH
WMMNCmRtlptBRihFtvfbpXtnT1mZRhKcYKxq3wC0h4oPiaSnrpF92rKJ14Cytwl/
7wyYyVCal7jPlboTxxB5gBELAPzPOgYMSLq/HgszXFiGw1sBwcZtrNv89USV0tGD
+ACi4Rm8i+xvnLqChFdDIkV13yoHdDNN2KKdkL0u8sY29m6VVMMm0zKc2yVw9m6O
yE0jzq+ZOuE4hamLBF+ij+jSukDL72liZrsrI8Za50YUcl7m1WPo974T8T1vyoWJ
2Nwaa0v7V54WkCDN9+KSOA4z07YXfDKi3iWAAdlbfn6dj0XDI7mW1R6aOtvALiJX
Nu4h6dtuFyVGKqfGSOJNrn7jMrCTQzEKhaU+elXz8A1lLwqM3Gqpctj7KJ3RHplP
bpFWbDcwgfnZXKbleAnh1QCMxJDWlTMrO6tDLBQMsPLxHRXm6arDJwlY3iM/T2Oh
NUJAWyVMofz/IS9X9dM0e8y0t2uYfFXGxNQZdE++YC/hM5rKL0tk6nL5zbiTBNSu
J95pTUyvO+rZ/9OI3vbFNh43DH5myq7kz77fH5Y75oK8baM3/5+GnXeYW3c1njje
dnj1w37Lcx8IncNMFVrJjfYXW9kYVQONT6w6J/ud47Q88rrXAoOr4ctkeOXZqyQ9
0Zv4K0iAEyunzsNzS+2RRg226DWfGKusxf0JS8w0OZC82BNAFRN2OrfeufboWjjf
Ou2dB2Py9tRjbVaKj1F428MojCLkpTiqBUld5rOE6R7h2CmPhpP87lagjj+A28bF
SNcZlEEvHJPPnLn0gfoTVi3QS8QUFaBLzgEs0U+zTQ5iNHggX53B0H/IXGOTO/Wd
1Pm5f1m8XITv0YFH0x9dhOMKDOkkmUKRlUQRIqlIx1NnNiWP/oojagvqDo1vFPkO
ci6HGQzaK/+T/g9Wx1DI/uFz3/p/X1FIhl0kcQW2bRVyu/Aw5y8cGiSxT6aWIDRr
+JcWJKCUYcUapdT8EFzWqZGTNAOuqP2a5TOV7aamkuQGRvjTLlygUqW3rb0yec69
dsuqFaOSgzGbHvv73xsRBK7y8Y4ZQAbejf++R7z4esDRE8RYRM+F+JulUeq8Y9J1
Y8iLttUm3ys7I4WCEq4gBUmr92I26/wRcJCPPhVmzFNU7EJYcbMeC7kniaV2CIo0
JMEK+rzbXDnjJGnAU0uD1svz62GS6rjtwup5IbYt6YTjsfYglhvX1A9SB1+6jszT
cSDIlO0A6p9AkMGXIXjSlIvoINzMcYUKclMSnkXTL/jxgrJ0zCWuSp+x853MHS6t
wzaPbcRIIBpCM5oMIvR7cVIHmG2SohrvDLWCJau58Bfb1Khg4fnse7kRmP6L3dM5
6vQ6x+3dD9c1jpog29/qH3p3Uyv7miOjkNOzOAYdZ2bLG6TN5/wpe814+W2t1EMz
9x6hsg/ymQBx8DY2zIiftUqSNg6jDjvbE1eDttVj3yUbzEvFCgHGWBT/MM6XYPfs
iu60xV0ZSNIj5mJjNecoS6pxzzM7Pa6xxAj2xSbCArrmzRfDfW9k/0AKHgfXHSfn
ccvN7bl/9qnctsafVE6PZ6uuCCkkiiMc+7TXapMhAOZwRy2QvfOXEKFTq2p8GkXY
0mF2WpjygouomwlY4gNdj7q9CcT3B4DtQVkWK/M+fpQnDpGiw1l/N8feTLe+hqBq
aQdDJLKDJH9N0sEdbQZ7npsH/p3JEx/IzYalww1A8rQ2CkBPRM1NtoOlBM9Y2qH/
JuCcnHjDY+JbgmxvW0Hm5vcUljgdQ9833aP8icV8DnKrcHPjy9Gm5I94ieXmr6i+
OB2Jm1T6u1wpon8uNJOBLWqcfyvHZ6DzTWYE1Q/IQWslpe2uBqsmcSD6Paj05cjT
KhgNv7OrO54vHZpAxXEG+3yks3eAaV55F6pHYkg+39MYoYvYtzqU+gUZ+8LhAv34
pyLzKYqTOoIW/687UioIrkD+dNFT/PqyEh8N9THFUXSp6qJmkXyOsinbMJojjEwA
2DP/gMl1g8AHnqEjU8QZWP4TuEMK3wvYQUWyrFfjhDTZD7h3h3s0Vn1OylRSV9df
iWcTp/xxXYgd9QwOXe/r4NYlwMPtGYzEM4nfV+GGugkHLeC35PTPm9ajAfhSLWGa
wJj7cYf6oFy7oHvkOIFk+jZyzx1wgzyVGY7SsCzIiLp5Vto4cn9pvfz+QsHoTY+v
SG+kj1YL8BkyjtVfdCw8WYpe5xQIIpat4Q7adm5it965ROS5A9vgu6nLiFcPHRti
QZfQSs2U7oFcY+C3LPABEuvo8pqA5jkdcIANGOG3h29BfZ9dKXnWQuWTMm/57aGf
owptCCJfQ1N5qDV8Jd1A10BFIQ+AbjnUclMNRG1xtlXKc1X2rj3oVXYGnL5McA66
kOQaZUwcken9oeZXudQloOVTH3w7YW1uTxzpEgehbkrOvpVVG+ApUFVLhJHd/18G
H7j+VGj/Zkwy9+kaNGWl30fo3INGF9K9e8BDDxXLubFIeBDh3kh/G3R6qaz6okdg
Mb9XRlKzPUqXesEgIpxtVrsTXbxgArV1AqMJD88LCtepG8evcz3r8rMATrZ2EvsA
umMYrW0Ai2gh05sPiU1V3v/LF5DfosESCYTVx3PPgfNXvOLUj0xHboPiGkna6jjM
8w6mCRHkjhPSYLHKqChc3LL9ExWVC0WxPyiHeVRD9oFaFyjUlVuZupUX1LXBA0mF
ldtk5gVgGsVCEHwVzneR+bYfcpzIsi6A+Od8gjEAm60dvFZdWqdZnshkdNaJ8v/o
+e+8pGurjf1YP1XWVAoSLdaQDPrJB+1E762OsxVMr5g5BRn1ROfAUhY8WIS/i2NM
BYHAGwjOKhwyWYS6+X78AC2SYfBge4TiRO5XIPAAR/FbOtK6bSKiPuAkEJmNLKqY
tjcXke53hKqpFebq7Q4B070kA8tQ7XOzKRLaYcYCuv/uTQCCYJ2EjZbPagY+l0f8
tg4g0Woqr93oo2chperBjc+dUW9E0ttvCaWpWNFN4iFGvmotBOnDR///1ivMYTiz
a/Auooi+WNuXtV6mOONRIVQx4eitN18vBfq2GpSy1rO3djdJZZPcZQxpmtrSEx9W
dYxUWIF7wLIRS/P1NCTzAmevL/6HDkKnibkjyHcy8x3jjarQ7C7OR0Sgql/4Y6iC
vXJ6EWy86sTpzwevqS1MKmrTt1n6Aqz/i/Xp0YrfDLraJ8lsUq8RQ6zmE3FtEj3t
pzyhppktvvaO0vN0kSfPIfGXdlo2CjMu2RFvbSpEViuWjLmnJ1Kt8BRwtqztE7Db
DWDbtdHtenUvgboNoN3LQ5IZL3lzWlbTkYkHI2dGnkqiL1lRHe37bwfar+CLPMBN
1kRPbonENt1IGkH8i/ZORHF+gnQ5TzUT3+Cnk114/mfYETvJWungasIJSVatiiN+
r7cmzRzDwlOc0+38+1pDmxZ3ZlKEfjh3nbwcf4anv0kJR3JFIIPvdh6IM1ymbQi2
i+NZxdV43KoaYIR7o7Z+Mq9XyQTM6mhoghWVYZo3+BH7kMcLAm87WBNDy64hDa/P
l4Dih0pCLdZZ0g7KsY/4FHz5O9oik84AwpqEyhQATBrSoBqyGowSTqCQ0+BwFr6u
PK5f0hB7Jd7FvrI4rxf+dY2erDh1U5p9wchkkULLqu9O0+n4YTXX6U1BjnxCnTkC
JHwxQ7vandUyx/hSPvxgpdeMOg4CN94JQygqmxUdcvyqGv9eRrdOzX+jtBA8qiI1
5g+fIgaowh2z0dh+qMlBKUujAFwtZXQ8hdfm2JYybLfX6/UPGAYPDJBIXZ+Og+aN
xnoJPWZS52cylm1tWGBUvy6XV7k0Ma0a0TyCda/FOcQPZ+tJ7eDS0IS/TgxmP4TN
h6XsS06ZqMkLctHBI359hcJMLsJPrnp9BcbS8hWxz9Zj9omMTCqpoYAS2UuJM9IT
VikD5uVsHBS40KUO6aBv7qVL72zESEFKJs3UsgPksiS76F7BmvP9576illpiXOjh
iUtH+qAJmTQLpe5laVknBSbZcieSsS4RLG1nJ2Qg09Ctvc3X/CILr+KdTupdqaIz
cLI6noZpB1RbhWiK1B9Dkc+fyKpQjDbC6ILERkqNjOTyCwo6S11rKNtCsx3ChLWT
rjJZaYNxfuYKgKkl/Ar8LahwV8dd+RLhf7XbLHl8t/ifAW3k1KzwjGYaCESuGsFD
ebzaU9GNhYe7S0kRXMk9tkqIyDrk1su+Rtai59d4r585USlr5PBqHbBuXV8g4g6K
T1/4VfDYBNc6+k1vDtX1eSZwObgPdZLasNwHn+y/myv5gbk9Sp1j8Jnpc60oM1av
ZfxdVw6k9UVtjlJMLo/8NjqzyV5KUCAdL+SJDawKmu14SXk61XKVp3h/JJE6nZ5y
CzzvIgP2zsW8yhgepTIrTVnRv8pyWAo97f6cD/BuVjD8gj1ZY1RI1f53zuM0Uj6/
JY2K32yLFWX2IAby5y2xYu38YK41mv84Nji+i6gJzSSDW35EA5btd1e1vHyCWbIE
Br1CBcew5MUncaFCF5f+eMjRnfvKVbYX28vSPagzKCG2FIYCbtWsaf5MeV5ZGQNC
Zvr7NQtAzVbxVRwBiUL4ulLur1xPeBjOh/NqGlebDEE9hARbFJ46/GFlG1pA+FL7
YYSUAlp/cI8vMRrM1vGfRF4qHGrGTR8Z6ZiQ3U5uQbVgAkghVPnN3pDIjkWLrh+T
Sx+LlFFjA7TEo+rGvF5dVIxq3fZbck5t1xNIItzx9RKQJSdNhkLx4afVRolHYcqL
LqB+sq9tcT+bKP96+wUnnTjBOPcuUsGrAu8FiY2UvfUbzDmZSfUmV57mjPMvUwkv
KlyDmGQ87of53vi5FaY3INSu8ro3RFPe6U4d7hnSgbZoOuE3pAB1UHIX2mZ6nWcq
e5JBvpcHOMaZa2ILbXBog8Srqc8cH0qf32ZmhVAvGHXDbG9w/8it71hHEx7Oh6sv
8S0tNdpu9fBTj21jNG1nQrSb8tN6ONvtg50eJ9UxeNPs77B1Hw7H54tj9uucxR+c
EmNfJkwEYdetoMDEmkVIF+nWoSXl/p5pBR0pcrIXXTGc1ntxVRxXBE96QSboOsaW
Evotn6Xoq3L0KKMyRcM5EzWo7bIM5AzuNevyk2X4tzyFfwrs5V8gve0WeuCK2oRs
TDCivLz2MwJZdqHHix1ZHy9JvonHuu64AKPecir8E9Wr9+cXzSjsoeTbaxJ/41m1
atxG7kGgzGu8POPV6ZC7ZN9xi4nNnNct7rH7Gqtv4x+kkKSfuVon1pJr3hphNXvo
3EblC0zlLz2ibw8ez9DIVuJIJ+/1XSqyMIgm3O32dc49wyrP9sWrqbzij+PvC0Dj
eFOYy3yYsCX2koTlr1dSClzLGIOnwVucRqjTVaDtnz1TmG6cauTxrEGwk0ARnWRr
8qET74h9dLZ519ePFh6s/ISIEAwTZgg6m1CGVKpKEvTHC4LGPH5cPdjd71awknX0
u9dZelBRmuxUxFf9EUedGKnNE1djdbezAFtyeSrE2tZZ3ceODOpaIsyjJA1Erw76
KNwnSMn9gQZ9eO+6fJdrXR1X6X4AECBrODzf2mb6UkvM8WPSEAjcVu+pyU2A8sxj
smtQteI53AejUS1T10ni9LD7wfmKnVElistWQXbAB/Z10O7biTl84FEznEADnhfg
quKu5EWx4f2ZaAjv3TQEHWMsWv4+87+dLPpnZNcPhVh2bo22ieLgRCXUv/GF+h9V
XMSIzOnKZzKTpOqC0dJu0dSLR/9YYLOf77yhYDyQ2ivczTC4NrYpaGEXqlcFBusV
MvqdRG+yHZEtZQj8UDLvI/JHleIr6tC/uODSHbfvHC1HrD9+uzeggjxNBt2KFLrM
ckTYXgamkbraUzfHk5oiSlLb/Qjo5Le8qTxK1AKJLFV/qDfdXAuMCzR567D5Gd3I
cRVSSbjap8RxX11r/SfERWKtdArSBBUo3zT8psJw1x75Te8RbCr4KUj1diO/66Xc
xKwEXv/wxfjLIJJs72XdAviGhDm2R+JWNEZ3EHE17ba4buRrTolrO1XmSJSyuWq9
Xd1tyODmV8gXlqsEzys7ikgMV/U6N00Ur0EEtj7G9xoy9z43mBh+RU/t/S4RwMaM
+uI2EGrj+hbnQO+c9pbdhDaDSxwIIPLeHmdDGaWNmD+FGpy4Jo98M+S+xAgLkk9h
JUy665qg3osM8fnlRWl4yorgAl7ABYjjcO77s1ct4E0TuV4ralnbpEHC70bU0++N
x5Fgs3nvIKUwgAu2Y2Ol7dj3Dq603tHrQnd3LZ1c2uUtZ0rTtovtqEno2lIOUGUi
U66/uM07cKS9hyMBaMh7FLkJ9PYqVXTFfFXERk2GY7IQxtohTKzTuB7Ux7npAgUr
9Q3EDoCDHzvu+9x0XWs6nbkeTOq+e611i34+jvDBpsXm4o0hJ8HvkrKp50gqQelD
B/KKVCKhAX3WWgMgsR982vZ/SC5c1CD4L48UGpA3WUSWSjuhPaISUzGop9rlo9VY
W1K+Zn1Xr6KGwdyRTLNr/ZZnyyr2AxPu8noZa4Dy1/OUTi4Jv6WaQ8KMWnn6XNWh
qB1nfE99XAh3KDn30tsT7TImHClbaWmoBByeVU9Y0f+zkfiFr8Rszti+UJOErgss
YY/ycL2iEsW0vFwUvhxEK/5PpJ2CmrLfiq8SCzE08axZZkW7/DFkIc+VJrdHvGsd
KhYnzKN04OxVDFBszaYkj/CLj6iHHt559pt0wHg2foUdXJYFc82z9BDhnn5wp+Og
mjJMakkkYNANVM45LzqBcvHYLSNCdiExQFtLjO2C2vV50BQlo6t96ZuY+Vr3mYIn
FXYW7RYek3CVJcyAWeNcLepcQ2NlojyJaUXfVApYMEdRz9AvRc2rYieQFzoKRyGl
YgJ8ZwFoqqFXEe1w4S0bY+W5wu0e6epkfwoMZokbqCJHO6r0fUoyV8K+xDX2jF+q
kXNEIkvlXfCjM117UyZGK5II6jTBfxqceFJJ2/X6zO3sdY6jlKTSr2xuhh9s6zQQ
MS8ioGeGRi+cnS2iiVjTr7w1WdL61rzQQFar0lPoPhb/1cGQQ8H7gqeyaKbqIvvL
MSCI2QV4/aEncqbsYK//Hw23247i1sSvPUOCLNF9U/VJtEk9HdeY4LVJR8qpdSlc
hLTGGO/SWPVK1kMHUTJD5U/QT7X9uBj0ruTCXbTUCWsooT4bq1JW1l/D7LXN9i6R
1LJpurnpEol8D/KIuovRRdln3JfTSdp9mom5/Wzfv52Ro0jXxwlp7ceZ0BlVNMs2
IpIaH6ez/3BEM0PoATPbDEWGpaTC8T2yfzDXh3/gGjQ5WWGtLZDfo0/h2iQraMhB
SU4MeeuIx5wxPya9pLQo3oSaZNV7jvekfx4IAmxo/muIA7P1Z1PREF0Yd5cNeQUd
oWVkSp6PvkibCjc28rudgfp7oOLjuAZn44My29c8XfSlYwgf8QYg4AQzU5zkuYYo
PzljdVeAc8SS4Wnmwqo3mj8n8xmU1C6ZDhvi4aTEOH8KfssruSP8OLpbQMSvKa06
tsoTIqvTDBnbsLiV1XDNQaAtNupSZ4560UlJD+gd1isNXBXe8lmOMhrqtUAzuXpG
YUUWBLBzAwE4wgd52FXl1sSNZtf7RNBgn2i4kjJj5U90JMs+XB7B5xHQG8TVyGXd
2gcSVKOJsZRxVrcOhRtBIypE3OdZsnUwRkP9JzmhWEPUKmALqDKZ2AI2KQYTzZp0
53sb0puUllTFASwXmYuhY3hmXpS1zSBz5/nEPbz9kM2za9ATbAIWpxp0053clu9l
dBz9F2MAHLtoguFmgMVPyPzjZfV7xSpUH2gpzqvFkm9nSnlYG+HgzvQkAFUz1v+d
dkIRMw2mbZ/h3rZy3DGM/I+nRN64zQz6vhYKKlSXxIAnCwAOA7k/oGMd16nyZF6O
88Sa+BV4PjPxtX9dPvN1anEdr2Ea8/aHu1PT4P1fke2S4BnUywvYlBUkSYzgoEuf
r4TfRRDCzdvHGWxnipDZAqtoFaAiid2NnU8aZ2UQKRxWerlrrG1+7EnA3RpXzSHh
0DWCssIpr4eVa/YcppB36vvxwjic2H7CeYi36eIPBZzG/xMAGk13Nq6E6Gwb54Oa
8ld2cE5WNErjLxjQgNxNhAGySg+yx3cyNIIY4x9lFGyGcLVi/gvTzodKZ6smyHhN
nlydd0sWCZcjLNLCi/ksge6rqxiQ9s3W1ugs6HHlQnCx70B/0x527Ojz43haNRhO
VIR10//vtgDCurBjAf8lnPxpt9wkwPKuO4G1cWC+mdQr5O1+ApTkH32nP2m7FLeM
y9CSSArRr7jG6Kvd0jWlBId/HKbi70q6JmWpo3NxzBmg0cA46s/DsfOwwG4PGqej
M5NO9xknsYwHLicRzSzXJpBy636ADdzse8kl2QujS4ps7oumUxYmmuqcO5up/hVd
mhHaAeGi7LzkHaZTYzhjUE5dKRI3FLZCUCXEAEcszMABq9rKFp9LXqpu5p6gj+WJ
uu6xbLbfjfSULfZXPgl5G0ZUd5Bbmka+LsJuniM14QBuLPq7ZmFKXAtSO/5NVrSU
XpDxqfDISwv7SzLQcGBK7sDI1XslgrJijltP3mh2cawGsPbyMgvlUSlTxz+rviIN
aczdYlXf8c+pjTGZ7OyaZyZfCvb+OmVqjMBP5kWWvOxb8xxJtw8fLoRGBolFvWe4
Q6lo32dXAc6kzcYPCc+vl2h4vPkMr6Kzui3EmdeS1aQolWjzhOG7Vs6Tu+MT//ua
gnZIG7tIDcZU8evYjyUt2+wBnQ1vKP1+IzMImfKXd47RPn/7uqSXSHyMrysCuKxt
9TOvimqaEpMrBm0UAckfT58mtSBg5n2pUYbkLN1C4Ebm3hTkuopwvSfGMlSs1L31
UU6btTuMAS0wBPyM82Gi5BFWvB3vuD310UWPayOIbdhikI7NPdYhp71TJ8kZIIkj
/CSX/NOs01e+yM2oLMbKnyhsofY3/sIhNqAX+8Wxx1YQw3ds8YLKORvoYU1Uf+rA
8GETF4CqNPBK5PXdiKkyTST00NiLSAa/xR4gnr1WpTrOT5bd9n5GT6YpWqHO2LCE
1fvmJ8dHWxya+G3X0aJS6eI69fweaWlL40O015MpH1KuzF38BJcyCDpl3Bt31B02
2noWsMgDutgXGpgIpuIRc6isNNhxoVyx00xMseAlxv0/I42nglCO+fC188X38rjN
kiS4W0+A679s3CunU8WJnba2TNnE2K2QBQFxOv3oEMpHk0u0YlnvFgREAwdUts8f
nYq+HxcnstaOdFGMmlbIEVRZE/WSQH749/tNRnTjNNUZcB0vVZslU4i+ZTtO+jtQ
qTDven9oXQxoTQcJ9o33UDdRWpg69AOoagE3W7FIXsfX+BTSkFpB/nQ91eh0UGd4
u5AJ3bOTwbQJRousOYaGMsskD5UCVT252u6RycT4MnNNETpTwRsO+b+pcUcHWU1p
tntN4K2N2vPLo9GEjsgAoZ8ZGToB1NC6wjHDM5xTrlRos+LCVjg6b+Wn/WGx2qoW
4dcmzLU609Oyga7X2OpzRImcdUIz1K/kpengpPq1CgD61cU2E5IineYDgnCiiToA
ROp2Rgc4iONTtH4IVVItbqjKoAeok+ziWadt+24QQxPjw8j9r3RbDGg0LkPA9xWD
rXFpGUGdrnlIytlgYqeXPN9pEM4a/b1d6a2c6qm94qsYkWv2gSmQRuGSF6NqJV3N
tOH13NjUpmAntOp6P6w+oc1mNaa/ko/kwLvF7d6S0x5h2tDlVNVBXU6KWDIt+ujQ
GOcpDi7uvVBIy8eSCPEN7S5bWY2MN3mP4eJ0QTYx8G+h747aaGxeioLQQNxszVZa
HyVPCsrBi0Ia6pnMmyya2/j10SbYdoiic+YgkDicUrawe6r6l4kxeX+hbgntNPWC
rvLyE8YXhZSXHFP95B8g1DkdiNxu8nhPaLB/OT0qrdjAWy4NuT5JRX5D+aQrQolN
66N5y+EXW6HKSuS+/BEo88SqBTTWC43sjAQeQNTSXb+b4sLTrpqtNTeypbjj1tsL
VMoP/tLeTM3gsXLqmsyqBxL9WwetIxxmXkzjX4G4VRu0kzGnC2fvCQahMmCxaNlZ
XiCqbD13Q/Xz8n0vgJktvOhwrAFpSQqRSrxv0iz5u1r8LgDJcZ2+3/9onnzPvFJ9
1KzoteZpsYradyIizzLdzUTJqdiHBsx6G+RtHeuNr62ZsH544j9qWmg0GhxJn3vj
99EOh7m47kzp2CrFWxBbCXpdRl5hTSEqGwlLUqUn9yzyGa1aTbCHEd5Wdfv6NgOh
6OYkqsILDU6rH0R3CZVyBTIu4vHyETteRW2jTqsETsQefqDhKLOOjvWzrYklJayl
GjwCIyf8IdQ3RjqIlOjeijJb8hcYLzfhv/ZjON6mQkcLYfmqcGZ85a1Xfn/e8oGJ
Irjgn7oDa/xcSrlYSmewzpHsBuYk0ELCcs+QUFiVhZwuVwlP1MK6WL5nKE60APxR
darBvSZA2WEtGs+7KzHI6MX1/pvxNAJJgy9xCV7LVvok96xC1a6f5PKcLWkkLIR/
mtbS4Tt5LxqCKKzzW9IHbwlQy3NmziMXqGp6uriHCKoJZI6ELxOKAfGG5bzr87eS
dASchDcAfaf0fJrjylx0i1tdq5kDrRvN28gs43HWPHZn8oO9HlhLOf7u78IxDBZR
rJoAdtmwUgs/4dDARTeEtqmINxe13Je9ktrXFMb9BTFOEhXA2mi2JlZ39bBTcmi4
49ctDeXN5S1v9ANirlkOj65PEyfBsrgfv6OKax28pKanZ0RtrfTvGyVvlFM/T+J4
mome1P/8D9XEKumbN9xV/7tY3rH+GYyZQB6TfJF4bftmqxAJK6su67dUOE2ign4U
xnOIqRm6zMU2nDGxwgXiQnHLLOANChdbJZtSVWR9vXnEsikcUZ5tU3Lt3r5tUhz7
hF88JNc98k6om5jlOaPDy0YZKLVCk+3ug3WKP1T/SjW2tFbtc0WhYhLpFYMErvtl
M/WArzx9swYyncUqwPRF+SFoEAek/WTeEUFLF4FZrFTEPQ2OoAzV/ecsWRh32vPL
6tDclX2OHejJYWmXb/HvlS1tE63bTgx4cbVnU0Q9/94WkRl7ecuLcQrJ4gn3jDDb
c4huJjIqWNfxttelszUYyl2af2DayDneprNLhyCBFn/lUm7dRR4U9m9vMmRPVzBF
CbnWAtJoYoNuTXTqm3+kH8x5MLq/UBjP9EVwsEOy+uw0pbWOKur97+dgC4L7Z3hI
9QCOdgasAjZOBg1inkap58GlWwcnhXmJFatWi20gsHEAXqKEDvz5dVS3G3RzetDw
5kkNRgtvfNKRHFX8QuywM13p9t5zRh4eCIl7Qsp4TBG/tqRMpFXWeZQzz0Uupwoy
agNo5w+IYqebGmaYST8wGMfzQMHKNtN5RuOmMJ8MqzcGbIX3xMG6g4TvTDAKY1vT
CxIYclbVLtAVu76CYQysLgqOyu/gGxGHpg7d7H83Fr8wpa97OdXNkkXuy/qFShcp
AEzfx+KjonJJKzeZsx+sG3O6Ml6oZoEm28uFG/JFCK/UIw7lufGvuKGTtxNGLKRi
MxGzwYHZ/pdjg+mGxSBrI5wGcXIv2zlE8koKLd1yjW6l2kykK+NvtsGTu5+njA3G
hROwBX3XABENZicV/wf5H9ZVESuFyM/fgWRIDWbyrz6EewMpghrtXJX7hv7OwtJE
AVlVlZXv8xcknpGR8Rr7XLaVqWwQXUCvQ5X6gM4XHrYb97aUOfMToCqHDe9BxzIb
XL0YhPdrhhH8CaRFUWnOiXo24uoSFy3wVypPbHq4CvdIRlsVCeTU7+OiQS/stFcq
82HThavleKVj4b98eiIOWhpsFeBvTTfX5630OiftOTNUSJzh58sm1tRCHe9CLadi
uUdz+Qbiw0Lrax2hNiH45MFkhqO1ym4CZh1s4Txg9bo2T2U0ekH5W8gDuyn+BnM5
0c9KAUXW+nJpdPr3P85Px7nrRAYeYHnaGoEWJzgL+Bfq3sAvSMMU9COGhP6kv8hp
SGIgAHlY6iCjnyvYa8yd3WtEnp887/mL4Jnx3/u8Iu0BV2nbsc0pevqBKv/BbzAi
g2TvBXD1li/NRxQi6nyFSHy0jazzXlMpTKagygWjiR5mp+F5JC6opt2yRUn8GKxT
N7QOxeLTf77HngouOGDk4rTbnnx3lXsML6CeXbYUB5CthsMOq20NFmR3nE+3y41D
JUi6c0JUebYzYkss7f4/YPbmJWvpIdmEKQIsppHAY+yGt5P3QGRfApM2pvM2YcQm
foh9gb5EljMbDAOkUiB5K+pct+IBIgkYJu+D3nfrSQeyJGjNS8uG85tRIjzFQXWC
CosT7ReLv46ibV5afCD7ybSoAq8NsbZXsMZs4V9iuZoOiK0Pe2lmdbBBBPwW7f5Y
ObKoCtvmVlBo5Fxg5hMrIOreaXYE4Pm2qnB7bNOE7XBg4Z5Hss2ofsV0rdYd0eRV
GOWxp4uXJGnVkU4Hv19wCjTGFZISAG3nFK00Ywq1BwMYREk9bLq5sf/lEDGrB5zs
imjhhh+/KlJTsPx0USt0wAKqzVFmPFeCb0U6M55WgEt35PMl/v9pQbiTO2ytEneO
Nmv7PaHw5hSvql4SWwAzdPB87HY2058zANUzWZ22EGYNM1ec3/5ZUoaORQkvfMV2
jxGluBv5T9zNz/9r6LZJ5cKORT4YpNAY0EocQBwrRluxyedmsYEgInHoPYJGE+x0
nK9Qa8cNGwiY5N6RAgLw/oq3DQ2rTSkn7OOw0wCKWL5uLz4CWd4nDTQmd55hjk3I
Q7X1XKpIqQH/xDCSpWYlW0QZeK2c31M3/usew2N3L5HhmfgkT7H4/3j22uhMFnWy
3ayM66N+8bGYu7JpLdGchjY3Wnpv6Ge3E+t/GxrBw2VqZbZEB0jDfXHAhIuMyYNL
ia9w+v+THqGrEtQ4SEip6/AKF5/xTnNlDNDjgORyFotuyLwvvtZZjlVPJrinjlFo
it8BnIGwZzzfCvc3YRl1hkkCBOUQYww3SDFMm4N/lWjxuILDK0FWu9su+FWoOWii
YFXBZSab81RuUNiIBisqWbhBaPl0VFc2E0o+8W/evsbUWPLIGA44I3o2JbLeKeud
3KHppTjK/c/64wEszGwtAcT9br228p6rtk92YnBanjbkp5700hZCAeRFQ7BvYYg2
/1AcCX5qK9caqOaROjKWJivdXrzyb7xk4fiy/7q4gl7+BlbYabMCRAi4PbM//SQ8
ygo7GTPzCcd2x8ACUbV+++q9vRYn6kUNj8jYFjEgxkvmJEVucVBGO0piVMBZQwEN
ZyKcwTlIvfDLpg9CWw+AzXDygMFbCV7ZZPBSAHI1nbHGhd79JWMOcTdK0l2IeqAY
S0U0EzmyEImsm8+sNrWB6y6L/A2mqxc+DSbMmIvyTM91aJtXTwKbUePLjMqqnuUj
SLRs4SRONgQMLICCTOUeCRRC2y5MttgKFuBpjUXOK0WQFkyg2GTTWUxLX8RWJpL3
7WAXozAmtuHmrUoc+aSzt36bDMaiDGK0MCyXOMT/I+Be5MMu/TRFO85QFIwwSFQ0
5qwGUwKQA3grgdsbB4iJueVkf7QRKtc/ixxq7uYJjwQt+H078QmFgFqbQJtTs9mr
Z0LHiWy2hM3Gk3B79mgHrD11u5TV2mNOb6mFMdGBPxhVJGRxSediMEqLuPdijB9d
dwFG8O53JA0ksu8dJDzrb+iQ3w0oxvvkxFehQ/oqhik+8Hq+1svAanZUSJhMZj/2
RkcTglKn8has9m2zXH9vkUxNjYVs/2OldhoJQCuTa+72ON6en4FcEkuTUJLQiosx
WqLk7Cf4+lFXgPFZZMhcun6HhebLwf0XDuO8k/Q5M8xMoswpU2sJrj3RjpH1BCfX
5PIVFcuRlE+BMDk7FmMIiESak14NNM0FKyhOJx5J7ABoYH/IzChzeiaYBQFZpWVO
tV2INjIIJWVSGA6ffZCnRwJt3DNxBOnTTUqTldJT2TaPMvuOA+YOl5dH0Gmuyu+s
xmRktSTN7uuYz+oLAJ99c0g3eKqnGinYqbrUbXMFekTnGDN1hPa4bZzL9Gj5cDVu
TAabJ5onwLajZzc2ltZPLsZvJQAqsYh/+wnzwS3MJ2OEqtdoA1sNFgIYqZFWGHHf
W5ey6594bV9M3jd2EWvYqDj7qEvdQiwcx3mbSwvvD/zAH2xINJmZDPBOpL0zQkiq
519yq6ke140yoBZPi5j7eWbg+fyc03YjpkQa8pDzToUisNg/2nCJJKqdV4OKTlsL
GPtN3BsZ+t0Z7DoUhg2IlHl/icSfppyH0U5QtUBuwPhOv+FTKtifPAjrc8wvjdHQ
QwPLSFLWGSkyUPowpIxQ7ugs670sT+7QHeiHWIkCa+N/V3iSmwAdBTxMHb8BUcaN
m4PRNvrCz4YdOMvoiadwA+rqr7Osw9NL/U1oCEU33/qO69NfDPqnyPYU3bRgSZiG
XP1YMyR7lprgHFuiNObHQid61Ml/InjJpPhzLUFOmwvIddCrdWrIdOk4Jrijyj2I
aALF1cAxkRGZoU5KBalEl/Dpc7Dy8JI1Sel7qMl8zK+QCzPNc46fEdT8b3OnUrnw
+fIb4o1MqXDnnbn+JjzqhZAQJ9Wqj9FK573yj++eZYKxFuot/Tlsdw+lWyrNloOt
xUYSnusIXo7rWBPGM/BSUmGDqtn8ZUlyCeOvW8RzDQ0iS51knJk9+dveRkVUtj6h
CUSsct3tJHY07nVIQBmd5e1NgfQj1P1rQH4SOhEmpoLUZaAqgUCWBxiconsSJYsz
qWOtd6I6wbrtP8t1rrsrlzQ4TIHTIKGXx+F4ynazsdTVpMmSnqvKVnQxCiK7wPvu
wm55ab9ZbsT2P2O+hkeROf95z0J99ecdiZ8ixekznUPyG3UVhWm0N8FyVlRpOTOK
/+GhY3grMf2HI+sTxFUbQPIGkkbmy+vuLgDJ/ixGVQ0sQ+cNjHfnUuiC7suKdvvu
YTIDEHnHpwKxo0bip/etljy174/miiVef2ZucY778q9+gyBK14g4sRon6x9LWRLH
C/hZeIGyQaetvT7k1cHBiXPwP80iuoegAzg9zOlIIPuHscunaI4q7wBih2ZcuaCQ
Y6MZoL4flsQVWSxEUcK83ept6pJnfS87/mGoYMiGj78hjDaRDC2HFW7rRen21Hm/
G5O3Pa9imEOOWDDtsUAlNUl6RaGLwm4oHd9PR84e2kBn6RaFNoxOAwMfxw3Dw+4u
VV7ePXhhXj43hs3h21jkj1dPBQDIDVBBhoeV5SEB22mloX+g1A+r03V8fY/aMpRh
ribAsgtLezhSL1eCxIWnEh7rLYemW4dqhA2krYaSw4KR0yaTFuBrZcZ/oTvokAm7
e76HTLgvLFa7Krr1mHqFyoBVMwxKErPoor31cjk5AK3LH/AInTLOBIz8HdoSK0rb
oWNf6C+avJfje87oKaja2KmxfafaaOKj3hONvRnEDVPgnwm5SYBMBMl7W0KPpsEj
zB/ww6+CiNqJSneF3/3PRy25qr+tZedUM7INCud02cgdKvahRiJVpS3SB44HxjCs
xHqEsy/ggtO+AaWzkyhWXUkJNY0gnaGYjUwZiBZ4dp1zFcP1bm4uJjkpHRhOQTKV
f7jb3lb59/FecH4c9bbD21VqJJEdvaT8mFNSk3rQPSTeKXVLToRuvTgjZKlaENdX
84PjlcO4A8w2KHeS1U8+zWjrZs5s0HLDSvn61rpvxoeMGz8xSnvkA8oG27Mq8tnd
BWZ/AQCKzcO7HTJ7S1Haxi6JrXvxnH8rdBODGwup0e+vRnIneRaYF4PaHJz5cv6H
0763nQ0gW4wVfHenrgge6qn+7C6VgADv0DL2iWBITM8huxmuWI9uEO8MnoZ5FHFl
0d19S88oVtkAzrckcPbjRxUni5pcpBlU39JIxOf0kgOlshQ/wBmH6kkQugY5FEpV
Dtl+JRyZNoXNhsCOBAjMjX0Oncz5kzw2NOtg50R/bzYshpCwhmebNlFEQfPXRS2x
QMN2nbQTJuU7xhXUt7JbOyMyUMSiYltlCHKD7mFtZw6h1KzSRfSNIlG700wo2Uel
xP2sL14rlHIrvFKugPs+wNctGGsetZuphV6hswcvxy137f3YbabdZrJ0rmLXIu1e
NtXf+CCEP3YigrPbA5mSLza6EGboI073ZGWASZRKZ2PylGms3FlIGr6s5twFi28A
r33+aOnZJNxzLJmELU1z8Q4BgvKta9x1ziMJy8QMuFz8TAmrTPU+aRjAR2g60BPQ
ZDlnqm+Sn8pd4kEcCE8EiQqiqObSsqRnz4Hk6Mc4w3d/5zKrCY8QWBd+2WnWBTpv
Miq533x8zDvZ5MLEfFXp5JosjhqaXo8S3WNbMnGj+4JlONi/HcMyAKDZTvmPuyAX
0PLvgycKDe+XBJVi5CsMoywpaIqbvMnixUfuKEFlyrNyLfkZzKDp0RnMraTQXZXf
XI7cKxr/6YDaIdBQIeKbdn0sIPy7yF93UsjYyH7LkTtkwEx3p7UlqNLnzF/oWxmD
BjY+ZFCMRZdB0eGTyyv4INJwt/VFJz3W8Rr7293793q/m2/cPzwD3mCvcnpr4CKC
gYyHBUYvuAF/yuH/YnCKK6eWZd7nFc/qKmL6Du9HmvBrcRLdMfgQ7UmhYrrJXGxi
EqwtqKZkd3iWtxSBoPuwWcGMSUvNEjSJ2t0rSlegQCYF8tRQ1k3+c0ix9rLyobMF
RzrLTJZhQaLawPuh+3Xa0SiL5t5dZCqbUfrNh+BIQKMAtQfX0c1Kp/lFdysc8t5a
rJ0DV9pjvXeFvJUTEnPUaf5lQ2CDatXvDSR9XiNp78r82/ZJqq67YCOQxET4LpBK
f0rga5WTDbeIEoj1HpgXMxO9gqXRPrxjzWbQBPzp5CPrOfwl/6B0B5FHXKo+9tuU
25vrChgheWovyiuqkNRnIOtzC4q9D9uduJQ9L5BsIDGbRI53aAd6SAeGdqGo2Jkl
wraYnrPyc+PCa9X/tddmUlZVYmmjeVcKPxrkOvqXYzUrIhVdhfZeaZ8Dri9i3NGp
lTtfTwLzOGUMv4XkFqXbdEcXI3LjUTKk2QT1AH+1frnfqxFuANnLLLi3Kxp4T0X1
QsGFAdJXL8wggV/lez2JxSvdHxLS4tvhX7mHJvoWJJtZ7ZQVCjkjTIZCJp8dEeDB
868dixqPrJ1PpmhbESaWv1oW9A86dQEjbmXBQ09G4S6B6C1Taxjn3e52os/F3uIF
vji59GglDnhsV33Tv/VbhPIAU90rmpODxqiUHYSOh7vWfCFZoqkSDUWrSVT2rKSL
nHzHi0DmSvZSaZxVKArHho27jpzPlEuvDegYe3ggaz9k5WUaGahy+iNNbyXPzfEN
ztJp6+UiL3JYCSAohat+LM/wtRhlolpOSi7P7GuqKC+v/Li1vUQU5r0q7Wfe30lL
vdg7c6zpFcdhxdKq4G7x2k1J6vz9HpQSSw7l7cRd9OFrXzNR2uAy6BED11IEfKre
0wC9dF03SjUXQRam2USAR3fhwyA85m8Ze5+RuP+WiYkyRGoW5BmSIc/ZmHSNrILs
aX0Y3rF9gIwYbq7RAVyI3QjdgmVfSGQU+Mob+3XAc7TZW1X0Ab/bbUzrMCVXN271
UokIhwUqM2FLIFCp43ycDM678UasCq3E4TkUWJuIqWL9f2OwQxvKvjbeHF1PLQ3O
nIqCEhnb+e1XfOZCidtRdte6RwgMUK0RJeNU7pjALLcaj4PylGYLvLP9XloV81y5
6nL8oE1z9q0KiE94Nkv2jafo/PW92FZPl/juSSUr2maPYpVXVpd/KT6YWI5GYJlc
GlTIJsONvhrIoPQcmqFWggczCzkw57IGKP/YYdoMXLzf4civpAsq/2NsvMFQKgDS
PTJJrYl1SpwJfCp4nMJ+7PRqiy5S60AYGhnjSoxFjGQHH6w2YH5IgOMa2hQfs5PU
zDzmCSZvXyQbbDIuVKb0aEGP3DN+quaQjSlZPWIv0lc7M3QvpQ1DOrTCZ5AzugLe
+FmA8W7CIFLlP1FYADuCv1CRQgRdrN29h+CKElUSRVXMujlZwJnUM3J3j/qE+kxV
DYfGhU6/OOpPMdA44kynaDPzUngJCh/w//O/t5Q0xTHyQUHkpi6b5OfZhHYJ013B
w6rO1L1jtcw3LFl7GE/ckgxvXQoEEUcsv/VG5Jb9Av0VlLaKOv9KVjDgzF/TxOrM
NRTgjlPsinPFbrSrM0BCg9XSSupRTCwb+kwvIPhM6ZkawZwcUynG76Ys4jHC3uun
f6XpulMFT1lGxAcMfQzqnFB+x2bfsY9hh+U4L0MJNIhwS49yLJIcjzY6M4+0JZz8
bLV4HeUD1r8ifHId6ywC+jSzF8EZx+KD+k82c5Xvjjdw6h1lBFO2PyV4fnSHVN6y
PItTQH/d2BqRXnUFbhEilbCSZsWblqNvzoawIaJ7yVH7JNJ9wlnDNFmiPC4JGaYW
IY9AfggGPnqbkOe+ScZthizP5qDC7zLf5unkv+vrLd2tMEJ/nT5HNOa0zN6yw19K
67Rf2Q/gI+KOzuxoioLbOfz/2Kt9wjJ1tXQ7lr7ZN/pMVRJm8mXb64SgadRcDnAo
dZKohlV4SHOczxY+jKpiKIPRrFFLo3oKMPS9hCumYRtAz/kJchRqGCvJAIZLjfQL
yBmA3aaBbPzE+qCHNIEmQ/xCX+AMY7IZ3Mptx+eXhV39g9O56dfuQDU6jr1zmNU5
MpaJ1DG/J8I/Kdu/DYq5EeMHI+WcskHd5vcG28VnaQBHtgKHZGMxu9ZJxZ78qTJK
4EWkfoLgz5RTPvsAzBnh9pEfVYJmXTR/HPxYCtOUz/IaNQD7kX3S8Fl8Y4s5Q2l2
lamDv5QZgI4ES4sX7AyXrZymf1br2SCxOKua2xArLHdMX3ORKbNVL3PQlAPMG/zB
7vlh/kB83Vkt5D+5NaW2mONTuX5kod4WC9XCmTnzN21Ug2fMsH1YzB3Ft7xRbhda
lQGaGtMp0BoD82AyHwLxhSqc2CmoE5K1qE0udGdOc1KX6X3tOqBMNToEPhzA628l
19+MIUw4pVwsQ7jFYZyw/7n5qY/wimPIcqkTxsYrGcClExFxrQP7owgNFtsnao25
LGkBrTsoS2oCiXmaIdB6Oe5JggF7wkmgXBIiAGT9ur0uECaY2xZm/2eRfV6ZzXDy
byC4b14PSUWnJ+SqmtbCwaKGz41UpOvzuetqsrhO/zSipYNw+RI1wCAt6i/7G3ut
a/iF9ENJXWf9fTKvm+FKGezj9rbz/5/7CaXIknYrfNxFoBzQeAyidbbDkr2bI6TI
r8CWTMZTeyc0Gu9QWKqI2RV62US/2oXhCzBfryXE4WcbXJ0SNQYvTgsFAdlvu2pO
pGddF0hn93KLpFiBP13UY1oqRZo0yUrvKbk5hUphDDvuXrUewprXnR9S3WbSI3ES
Ew4oRpEjPPOZnE7R8dhX8x6KsXQCxXlgfsdwTMYNLWdizeNibQPvM657HF6iFSxT
4GSAe8Spl09WvaGopf73b0vJrPga0VqsWatZy5e5/5Vrqmwic/F3PrE78nYnJbRI
xcerIXS6kQjtldXaEqhwiEwxFyHPokZIzB8Z6nKtUiS4CwdhHdXTqi+Gmzclqg5v
vxIwBX2h/UMHoT2KUlTuKTpIttxEVYhasUsxmtsYZMk9si+svkCTERN7RmifsARk
Mb1wOFiAEGDxdZH7EK/e24wu8pX6+7lznyjn0eMgh6qfuqdW4ERJv19DQo7nfz0e
LRMKwRq1F5c0hA6wS9+ehITpyr+rqAEARQDPuFp94lOhIppL41a8r3BmevLwZ5ag
wMZELYHJVVuxKTxatls41/h3SV9JtOqmpvOoDdr6HtBdksILhswFnCdborxciVUi
lUybbw+7h1qrtyo6oRtQfWyZ5lVna6YjF+DsQ2LX+QZ+Ujf0kFmrD64KoJTC87IR
O2upoCkdLb5df9qI7jXZNVFVKUNvUNj8t4FTd1swq+/sLtLrnJoR+WcGhAXStHbA
O1lcoTuZaSpTUl54quYG37cw4Wi4XrzWNYK2w+V6dJoFYn7zogLXdeZZtEEbBlSQ
8PLkB8bHkwg7AZmeu7Oihx7G/l69w9VYn2DGlhOqCeADvehr6ERaf7Dr/hOU1lzs
mOjPqn421F6Qz8EaShk5DvLwHr/bSK1TF7FfNTQ8LuO8QEdSDy7JCiJVXyz/IL4F
n1BJGIhgh8olP5H4us/9qSq++ggYXNYlW2KDdNqFu4bNGMmmcKjTES7/xyndbCBN
nq8yYoBhHzyBEiEf3AgtxGOYEWkRGd+zsT48jhuda8BxTivHU4AyitX0/GrxAIT8
kIy5Vf2gzHXoSRYRGzdWaTDoct5eZ0rK6GCXU3TqWxNKf0W1l2Q0sKD9cO4p8HGk
usAvmZWM6VF5wKoFl4mDKfiluv6szeMgvOkCvZddaNBWmmBPeteXf8P7mCelkF4I
7s0/vTnTwnC4zPrf4aHZT9qNIXmK4RQOwz5ZYJpiTWSBnbtZu5k6yXKYPBV07K+F
ZHNUaNtW71Z4IchGE2+B8RjqvPIl9kxIP7KPp6+IjduRrWJoyq8J7HSUmDkCJkE5
uP7qaW3afMF+qGiZFnQ5CwpK7TAD4a3eYxCQG9t8OIH3uGkhpmgnhrhpvOHDpsda
FNLIZXair3AM4+BADYN9e0J8rRCqko/Q4ivO5INv5Q9OmGFmu5CLauDayjXcmdwR
IkWFU+eKtVAYjh+l1XmhurcCUUmghCosO9jr5jO3TWmH46rbuW0BM3KIMPjShkHx
+PdNV5EjEJUUvk6Hw7iuRhJxtwFJBsXaPCJvM10PmpoRPt+8YTTqXYvEdspkxPDt
Wi8e9JF5vKcoA34c2GIlf6kfIfdu6BYpF90fMwNtOoH/HSdUNlLrJl5aCKLkae1y
0aoWV/EzaKHaqRCPesxuKkdETKOAglfbZfDqWsqBHX/hy740Lw4zOsZYSEn1XNpR
SgCSF+bxIWTG1XZ0OUn/EzBxl8f0PzpUy6gxIBewkPSvzx4gvF6TdgkPibd5pI8q
CP0ENDImW1OHeyWSSUE8JcEFWExjeXi7l9xtVZKo9+Z//OG8iSgFXUTQnENbhBHL
jAl5w34COw6iPd6hbnYRt5fx5QPVvU+7+7LlRM8eE33zn6LdNVI1mPpzdbW3sAcX
sr5KZUfbnH6aiTV77kUIeYlvJ5xKGbphNZcK0VD55097O1s6yJUa0FrGpvehJ47s
s28lmiqCUjgKdGTWCIE8t5YRQs7VMJ6i9Iq83vCcMdXb6Mh5izBLdehqT0j+xuK2
e7CH8zLIhDS4k8PaJK+baoXpNlLA9XB+e5mf9QMvrxByUG3opbnlq90UoIVP/YXX
f80ZqK4Fkdw+DI6HU0gu69yR7HJDFPcSZI2iwEEhfcKPFhhbsTLRxPR9mnid/xDo
JZKhi3JY76pVlwnXysxR+rQnBAqjwMxLo9Na//gLy0zaqUCnM10OYsjH/v0KDrsH
X3J0amJMyFfLM9iIcXIFHyqn3XfNmyYC2aJDlfjUR8lLnBFMkYXB1CS8IewjViMq
ifRvucFTM/EDwRRWsZgOPz7EcdlludGgoPcwNjFN/R6DU5WKCqzCQs/mIF7zu0C0
0cXVxQngR2oeqabt6orbu7UJo1KB+XtNus++R2TYF2OUgxpuJq0RkHae6vK9Ll6o
k8y16NzmGRNcUhTrhKwwAsEcMg3ORgYlAyf3X8nwf/MEvzFQN0Bu5JlFkzyecFNQ
pcPbv8BiDBEpbr5YBi40Ey46XTOiRCIIgUGRYOELzoA4YHG2KxkWGOOnPO2Ehm+t
4OvIHS60dkwCRMw1AenzRq4t+CF8+K1g4AovgklopzPWEhtVj6TUmQheUASrEKQ0
/l7B63vnlW8n3W1k1lQTsmOv8rxbafzwcNkC0nA28knRf0fS9e3w24OrGN0XWBvH
2AyO/vJeSyC01r2FXkQpnObbH/pkdlRTfgXx71Az0+xpR9Zk9dj7rHI/LTR8lZqp
KLOCv2r8Owqc4D+T884Bi4q51WtNEJ5wfc8NvSL23iLaGnOaNDhMWm4kDkUdzxOr
pNWlXggJPUx7vXXTJYF7ydOZ5VSOQCV5oX6RLzJdrpMIRG7ElSzKX3xd3kHVXsVE
Gzhh+qQaX8u0mFQ8tcO6iSuhB0WlUT3/tbDlPGOHCGf+6NVBAd0RyfgnisX9n2yy
M85r3VUoXvxwdFnVwa/NRFAwdhZzZd6MBW76pGc5SkNzMXfZkvL1RcC93PPwqrNJ
fv6Sq9KqL56rrffzzSwPznA8fSq89O/ArANQlXXFnH5lg2kjJdbQRV7OwUsYC7K+
8vD2z1lgUZVos9JeJXPLfi5I3Vrgo1g7Ypq1tWsUUx84M7tq2RFZMNTuNLLkL/eu
X5TmRSh3tUrxqGArZ1xD7SBFISml6fL9vNlj7xrC4l4A75QJpsZ/RpyiuGxbKN7W
ctg3LKCaOUxAxzPrrWjlgxBUTdJoA4cZF9B+Mek7t6RVWL513knB0tATVVDabFCv
IY7uOBazq2Uaa6gEHEls6RXaf0YIrzinp06mJ7TWiFyCUrE06HhqqyZYL3xXxiq2
lq1n4kvPxZBBe5r/9tMNLIkdbl65kHuMY4YXGaWdgvqcaJ7gAJfV4v0cWJoQ8BGZ
0Y6jF5VvRDTj5kLHd7fIWVq1orDdoDb8XyJKoVwvkFe9k0tSFmHmFx7BMFOWCAr9
QXwHGpncnO+rgUPv/6LbUZ1X1wb857eihH86rLX8iFcyCTOAagQhajP7jY84yBKd
3dnd4SmjZBS6MCGZXT5aghuufNLRFhSFXssiuDnZZNGR04MG66YM4OEoKiuhiUwW
ardJ+O4XtaDIQxoOgNGYTKhfvnVVN/0kEWBVXTX2IXXscQ0YgdAa6Aqn1c4bcp6g
xBdwvNIbhf+xSndba7rMud7m5bAHo+4k6SYmMbnQCnybvHdUpLEdVvwbHy2G9qC5
wdPMbVpYFvWtYmIW3P4oEF+cTlyMJVzhK42hk9yg/6W6o3w0EODlwg7rDdsjha3g
U9gkdCl18VOG8IsdE1e0eFatUAB5r2rBbF+WCkqT1gm0Qg9urYyuJ2X0y++IGMPY
9qvMvZNh5eb2nmzT0jD1S5tiMWtlWrvK0EiSp6Ea9xOrlQVXp0EYkbqbbNhJtEz2
Fw2LYGGyX/WaBre4w3UbUUjeH/VUT1yska9hfgS8xfPvyB6oKFicZgVoq8Xf9DVp
UEGs+AR1wYbuIMneQVn8gfKczPALJJ7uYudwp4Zq5dwykg9eywKPvC26tPtlC/rR
jnZq4uZTyd2DqY4svN0gIvrTo/cSVXtc7Khz1qZOVGGGG4iX2qCdmufZipHxWHZ6
RXoAKkr7vVjz1iAN0LSueRGQeuM3Ex4ov4ZM7he/i7QJCiuFetN5ivsFsMYZf/kP
SyYT7PlPmDhvQgcDUhnRZLfnuRo7DhyuSjeVV9NCtl7439o2JcXVwR5oswxMsnFS
NfvjgKLCp1+GV0Qn/CaXC04pPpmoFPu1DYNLr8KStktBnOrBvGzYSTsqsGztAFcG
GK/haWp14BvXxPBQaQTeqUQre/txvPfIq+wvFf9Lsq+dzVrJemVcz4THfcD4Od74
Pre3jDv24zWTWuwB9HPEATFp2rzadN9jhr7RljdzaoCK8Kn5VJPiwFSKPty5eULa
cv71LuH2VVx6Zf87pQ5FbrImXpprL0nHalNdLup/RIioxBDIVYqxy+/GpvE1571Z
ldTDjX75x4oDW7QykSkQcH061OL9EPTHchSsNRmyGRkc3zR1JY8i0+4jvp6a5H+S
N8ql/kUMkpQVWlzSDNLlgQiwJZ2X95fJZz3rUTTZH9h6we1QXJUObHo9RPgWOGFM
C3k41zC59Qlc8UwhiZcEt2bNY5Ti6HI1w7lXVI5txgOUpnlCr+tCFNn7x0jKFPus
oPGO6nOjLV4Hmw50of2zYJIbypcTWpK38UcHrIJ37ahLVsxstDTzHDPYOpIZsu4B
G2hZGWiOk4vylX0Yg6zOifrm7EjLpqiHy01unUl4hjsJ1jGPOU/QVvil5DpeFWd/
dsKQgI/xF1Rja7RJySqxApHkLhu0hfIOd1say65uIr0OPnVbu7Yve+5RjchYTTWn
FEoXnSFbU9AKKeXGsMLK2H6aLGNn8mK8kDYvNjIhmtJNlZjtLzHaHmtt1P3rg8a1
IW8TPRK5mQUpiy9M/M/uj4ylGW+PrMWeKE1hneCysiLRVvBTPFOpjfXKGBtaAyAO
LRQYCOLOCa+3NQbFrEcFAKVAKkIFTtQf4WBVzYF0/qIx4M7EWpgTAhZNL/xYFDXj
pQ3vb8TE2JqJShxdC57NVWlcTJv8wEfZaAuaHZAB2HnQicVkbGOZA2aLegwVQJFM
cme69XFmCht7gxMxqJiq0b/mRIK/b2cIilstN63aavCpLtnFZDOxbrYfTU8UFTSu
SdzFy7LJVO9AP4eimAEzmZWEDpIrIpGt0zTKY2TiwxBn1M6y3HcA+hnIvH7QauP0
4b3lqeSNlgrC4IpDxVbY6YSKnrDPgnlhesatiww016UMFIQ82DaI7gL1Jb5kuzd9
YQZAKEz19o/fiKuJGRoPDcBx/Hzaft1qHK/spbmaM6eq6ywslwImYAOAbx9Laikh
NttSNoa/rHDyAxyQ5W6nnhl7YQyFSE7RNXjrmgajLb7C6AGstORrWrIk0EuKndWP
g+EKemUVCNDPgi+6wNGYrFkdq1TD/ktRkVK0x3oy2d+3qgynksiWsFMPrMMCCJA8
k6IuUymXkRnhHq9Hl82rYmF0Z3+IwYRXru27pLkl5+ocVgZtWhw72ryiAYI8vwDW
qtPo+PpL6jOClYafzw0NinODVBJxyp/JKuZ+yjaQz/KZ/AaaEtuORnQfa5u27uuv
hCEmtaF75dyoAVukm3dAxrVSP2/4OFazEK2G1ITxpRcQgFF77XecW2cf1BRYuZIB
TaR/04fEDT2sTmYZTaRtyidRR89R14t2rKl3EWabbJSl35o1TdmBvwVIddCaG38g
ytJnrrzpmba+v8Zw32ht/e2EwiARg1FLGtZCkDhfHJvs30NMdaP/bzimngscMABl
C6EWNd1VKVaOWM2/38xH+FUYy5nAwvWZ2emanqlhj3ItHHjiRmFL9yGPtKHJlprp
DO17k0GNXrzwAOr81MAElshhBDF7tSL7GYN4GbvLaY2rOWzR+Pq0/uRATxniX1GD
OhOLf4jpzlDBW97+QV9JVmsbnZG9tAAIlb97zEZjaN49FeUTG7rhPklreODFK1IQ
6aBoXBm0/jY240Q+EBAzrbm0FzrkxLAus4A5c8S1ted53h4VntN19TpM7vILqatJ
HF4EK2r1zpss+z+goe1KdpCIMOu8VODgj4WEC+X+ZSMxdyJbrioOQu4PnJIzLBrR
pxTgU7+gOVEfPVOUmlqPtIK22tyYl2tfLN2hsP1NZ8Qfoq/pkBwCVGP8j+ntmaxg
3+hnEiPmUFHL/TNhDuidpVKHvKiAtOERTTvPAMUYg8ktgDQERVKC9YfHHoyC0wnx
+bEmgznbtvOo1X6NE+sDXtw5fA1Z+PmzYTPBTREFcswt5RgTRcKIbB/qu7PSh6EL
d3Oy4yrPxQbOAAjbGoY/hoCY2JvygDCY4EQxgcn844MoOXTGn3G0YEacNoAfw2jD
zKHF3hgco/Rn1X2iVPtJs0+kEY5N+7G/32Aiw1NGI6SSxg46/ghBrNGaEMcL5D61
/yG4cFbvqWx9hKMRHFNyzczKFHLQiU9OHXYdtGCmJdR9eONzHwpLMiR0xZssKL1s
Mw7m9POKVkGYlVBPRK/6GgfkVfpdgqEs/pZjnAoTeZJjv5LcDAzJQ1+u6w4i5ik4
2byNj8DL53Bin0CAXpb9iyJyNumU7B08qi0mi4/UVFGN+65Pvt9MaBUWrOyB4Qbs
yeYKMz5BUh6n5F9vBzPJ6wV9axTk7vWLALTzzmVFAvufC2pVzudx5Gy5wEnptPv7
tD5NyKAu/zY5YuMcT29V1x6BRDq9vs2fXhP/AmLqNe0Go2ipu94BzQ/dQozy6N6a
2fAP3SoQjPadOpMcas5nVXjdMuA7vdFc1aOrR0xVkmzfew+I38fQCLNmxO826okW
qP2f3thdx74JFs0YWxdp0SpP57uhNvhWKchb3ZVDkWSmuRF4cOcS4zjRYPuqrLfc
cfhBI4LY9uQTPCQlPH8E1ZlGtHHc8vhCJOF0t5q64ym40VqyznVO2Mo8m3V0a6uL
TbbEH1QgE8CPLlfqOuVxpkjKks8LwAXYWNyxSCFHyR/T7YOxeCalvNfH8KpEjdUZ
BMDGN6kx+WUMAC20bcNAt+E0CSXionmjBUnMuyBrYmWHFvPwv9ybLYCUcLXIt+SY
lQRQ8G7liCZzFSWgq1w6pQUu4BbfoLkOSdgHx1jessFhFRPQrIeEJeDVIKVyeOwI
1z7uTjdRYBIiLslZ7sVzU5QPu4jIJTtvnDMvSY1qkgPBlKUctOBtMWr5l+nMK6cM
UjChHsboaLH+vKwzThs/TxI5BMLuPnHb8eJa7J8/S20lHq+yOVJeTtcXD3z4H86L
fj5gMOY8YRvUOt2hM6w0kurtnVAAxSflDEZo+DMA34ZjEwdOBIh0PSpVEc0yF0yb
9AxfQ627bEbokicnYvHs6L9kdnnSlIrTCQwHWFzWSBUjVKrxM04qghF9ap17h+Hl
Vkf+nuDNNDy7ZnWyJg2dw3zpas2bTNW6B6p/+DSxIyIwj1RSBV07jCHJp0kyIOKi
YY9BL6AT5SKipPre04XKj7muNsPvyFjGcvTtWt1ZslDA/NrO1cdF1+HNi+izM/h7
YxUNSe6hGrXJahpVFDA9KsgXwL/oGc+OvmwQ4zzUc1VcPTVJ1AR37BFQHKKw4vii
g+c8mFahjTQZO1u4jqjjq0IA2c4wQFN1NsxfoY09BCPa8iPPCNecrNxLhAMTz4sC
hw03iit3GDm5MumVLpFWaVqTMtXG2aaqIsVEljt/JCi0bci0DbfD67RdUCyK4kGP
6rymh0aPQpZlhDMhVDu4cyU2tyMbr2jkduVrzKQbpsgff6cm+UIjo0kgvlnMD+yo
vlo5v+D96C78RF9ybmNyyVBFn3zkOBhLQzEuGd5wY/wMjmUUHesnS9cplwMMTHUB
2niTCMlqPBJVXRmWuTCqkWPpm6/r+SU+7CvkH3Ccr3A4sUTIwVqI6L1QLVlAl8tq
ujZKkYiGil9peL78y+Yt3wiZc/slHD3OfJRkVJ2PwM1613VWjSLR8VW0Glj/jD+T
G8AsonivQiEzxMvLFDES4aQDDJ3xmn0r/wWPXauPT+Bat634NyelaX8ZLWyukcK6
X7F87UnhvZ10LOR6SAKD1ErCgsK+59fFI9KPJcT21a9B3VK+nPSxuYh5OK+6Q47e
wyMGWDU81rQKsgBTJMiNs5ENSzfUEulNvRg+TlVNct6MZSrU+sysLFQZmzCInDvw
uNK+XF4EFOFMalwol9U7F6c31dt2KOYEexdHJxQvC2xkwGFRfglxZHBxH7TSm0Xq
BSdz24T3NVNcHFP+vB2KNWx6w1RW+PBDFxRinBICVdZNZF84G33mp7b31Dy4nJF1
mQ1tMKLsP0PAHpYMS44hs6DdUAv5GXdVjp9yRJP9plKBgabIEAIJ1dV8G3OnsJrs
YhTzpJBjjTel8Pg2o22h36HS8MfLe2PHUOSt//vH8aX8WrJJFtBYSoMaE8NlStjQ
x0au1MwQnU/zg9rp8pmWO5w2Nl6+7/zuYTQlvn92FKToBWLm2FQDNMLyZdmxh4Md
zjdJgxaRonM1Vpb8zR9QuF8jYN1mwoUZR38XJiin2YZ4aUaPPTkL0OY/IEmITTUt
VHfXJZlptO2gOJmh4lAUbXgaoEWX/cV7R/vvRin9HSfgkoOVKblSojRuEAbu9n82
AlO1j5sdqEO6szaE5r0yZ/irpGpynPX26Xky+oP2tjhKKxs1sd2P4BsWKA19lbnA
3FwGionLi5nSxEEwgNKn0K/59Wee0abws1l8CyhaZrPJXfmaru3bq3oim8HuKKnu
rf/h0Kb9KyJOSNG5rsGxZqtACeHvQrpeE49935Xlx38irxONJLjpd+MJ6eUoJAt2
sRVYrTQi2vXWemQXe390mQnrGbZqYKUU1knZQcYIxYw75/rbBWf+Y3LOfWfvCwLT
ulnd+HrkhmoBLsbu1CzIMzZzwLtOrYkablSzN0TrXr3sJSHlyVgp/nIW+K1P7Mpc
32endRONdd0Zbv3jyT7UK9DoyFik7pROZOf+mOVFZPaE3f06AauHAmjZhBUps6QA
0ymLK16x3dFOD2ryxI9XxBk+qJ2HYDkS3mXObrxCpQHiC7jIz/tHdhMgBEf5Q4dZ
BOzxRb+JSjAw67C68u7xftOM7Ly93M/WAnOO7MaOqVYHhQPn/xYAwAiD6ntyeZjN
zeJBnrocQARg33nGcR8S/zHh0kvVArGVWrcu8JtUb6lhBY8UM9omkzyRVOSgDYMp
e61EBJnF1LuBdwYCUgsnXNaBLO/5+BpFciojk4QP9W34f89V0F519JI4FXvGUCJ9
kmKLEdG+4kcyy2NVRw9hMz0reYzAGZwpdLYMvTFJFx1b62XM3f9Vu7y0Ht8wAL7w
wA+St6koM23ajW+EuCYAVJT+aKVV0iKTxCKZipss96O7tAKEcpPKwxw53mNH8SwM
nE4JQShsQu0okJKeMUbZIRy9UDyoQDlfkogx8G4zKHPi2zjRzIJiKov6SyzRM8eR
rmx4xDs6BhyH5kjv2bUfbSRb4/8/Dl0iMBNoDvBy2xdhUFOT6WhvtChFXVuQcQGp
nucXBQfpq/EZ+QVdcKOCp+FSP5iDpguSZgdefAOiPRfTCrvJhDmlGBpzckuctgEE
N7grTxQ7ZTB/dOEpGuor2/dWsnxPOdMr0TbNsl2LAmjAz9fHMJh4zvF+RoX/mk9p
dObos3hznTIgiujR07cs9YSWvNUNC+U6Gc6pF18MF3uqXpS7+0/cVtNYYBxpwaqx
jheaRWV+SgJN/Pw3gGw1qzWLRRDtc7T6hxPRfOE5gpDxsSwQRUCdm05G1wEjiBWi
lU197YSkj/qsBBG4qeqTKYMcfImdipmvm9U9Zy75Zd9cV0hXCHm+9X+dBB+A86F9
AtxEzVV7ZetcCI+e8mmb5g02OHP8v/UCTA5niVI0F/Lu0mHBUjP6/L+Ec/RoiMVA
RiPHtvOlJw26hO96Hlx14io8VTELNVE1+/eOHLl8tk4L3Nb589RsrAqFzi/QzboO
PHgEXxT8Niy3feDJoCam9GcjGhqdeqYOVXTgESY8MnmzeZPMFqBYHiPy6tLAQ4iY
wRCalCPXu7Z+D39rPveYND4bnrhwQcqEpLC+KAVDpZAQrRGiycL4AOSSDDn1DanL
hnPkUpoQZ/pnFNNudEql1KcqVxQfXIx0inwSDRnQFl1pOoHqafZY7gYpGbZE5hSR
mVOJzwEQKH0JXNHJGrId7IY/nDdNPs1Y52KvmVnZgy4zxNoBPah2LxwMf+Czb6GS
C/mf2S0Q+Q8pZFQ/7TBo1mN3eyZCE5ItYKP8d85LEC2dEUdWf77q9KZpjhKeRUDn
47Sf+EbcZxVADSS97V5z1IQ1osEn44BUDAYXmm7RHMl2Jj9f4bLIPIo9L6t3xCQJ
AEVtbvDVMwiDn3qziAdKAiY09mPJvDWX6qQzT6zGjPTPhVQOxnfLYtL3nRh9cqmf
0vWK/X2y8QWTBJ8cTXBUseBFf9YixWGDlKn6M8CWidb3o/iqX0wPSITYQs4AkIws
zk7dHsJbGgWeH7mw0k+7MoaziqdeKgpr40dLWW2drTtu2NX53JdivlmoVGu5Lx4K
zZiBFgfbFvNTU8oYPjj9H6uvrR4NwS/fUytBecpm3Px3hu5GhWN4H0wuULDDh/6G
1R/dYYAQr3YdT5cRYCjbDvK6WjOtlJ6JJZD/rHABZ5lqDtEcJiUEsdlMfc4IJbXG
wy+V9qlCEHo2yUBFTVRpYy5rTNrhDMvItmECni2g8jjxEf7SbZG2+gxxdf4o9tJR
TfWvgDZvVN0K+oOeYUdCoH4fXLWhfxrSu39juN3QUxO3mSG1KhqYN8z9G35x2TFU
JRKarqToJBZqfjwQPXE33AwJi/qOT0e4gimvZAgAlBA4rha1lKY8gLj/THqTtsNK
q71IHzt3St77YDz2JApxaBYXKo3kdAMw54VnBC46TkmKhQEIdmXnb8lw1krmNGGa
8pcLxouIEii1VoO4QI1JOVIlrZxEkxhzW67KGiZTAA54pxUxsmxl+apfzzAbvvTp
C0TH4PsDdzXCdXXIYVfeJ47Go+vfIfd/eadyid6FQBzgzuJfrMCoLtaoeIBXlXDV
R+Qjm73DNQSueRrxMkbOi8n5kn3/pLXurau/mJuT4GmE2oRYtDWqZYdSbv/SCajk
bDTNVGQWkHYy+9c+gMdXu/mkhz2l/Z6wvDJb4bghRaVXikvjy/sfu9OAGQl1gMVy
GB68PEhDIWGhol1XOeB19sB/1PIhmknYtrGHSNQMqqFUJCLAJdKWZp6wW5nWKNFm
SiFBmFtvJNc/83EPgOhojWPhkF2mRfBL7YqnWRleZSOAEpSopNsj1wwRv8/C4X9p
w9EHpsn8gRSJATOLxmOhJ3m5m39swHjxx84k1wxOI6cpLwJwxejf+Hjv6wkYxYa0
f8ZOykb6cCSGKSlptdIxdzWeTRa46+M0PYEyoCuIBW88gNW7eOZbkBq2pNr8e3/b
hdesYyEIFm9nGTBIq3/grOXpQ8J7yVf8uEIcDLXq3B9oqMXy8NaiY8QSJCIgbegx
idPN4Hl/Si3kbJlgi5nkXSMsqNFOkdNaJaNerazGiCyn0nO24smm3nS2GDhi0N9i
ntq3oM4KsBDYVDWIEL3QFejL6pSth8HUs3pRjoezo4MDukPZeFJQ9tS7h0OYj88h
D0DIYOxdfQuer6Ow+KZaPGLr9O0o+0Ga+HERQ43rQlgzB49/C6n6zn9xCy0xOus2
g9Y+NOWBrkpYwUa94v8BObAqLbsIO+aXUtYdL1CmwXWBVX4tqjBs5c8y1xlmTwSA
LiKxNf55i0Lwy1nE+HISDDJqivmP5qqWERVpALSsLIdJQFgPHd/ODHu0t93cdpgi
Eh6MVszfeYIFiyt9/C305kYzrk6TaUtbyLeDXL2D/hIvciI+RQ6FKgImc+Zz9kAr
XMHUf2VQrvPWdUG9jf42637bwJcWHlkSTcC5dmGH4kgHFi+vgzBOuoO4l6fwuGMZ
XoCB8E96wiFVj2NisM9nnuqGkvioU4o8WhbwD8rsBF2hBttqo2BQH7XWzjdN+WeL
xZRHKx/F53ug5qGR/wKiFsg6NF0JJr4NuoIjhdgUAKuwumJETR6kWHQp/VbQy0wD
oBdlvcNDlssADFxMtkh2Vb3epRDcJWUkE6ZJezFA7FwW++4OJPaE9JvXO4uqZcaS
wWA0TFPpyJFJhQwsOuU4GTPcOuPmRuP+qrTTb8+kfpoiej347t4HZdjFKXMLjAIm
vT5bk4vPCxCya+/euMJsnFD301LNbbcULJf7yp/F/tKUMJMF0qP6a4zlh9EPorXW
jdE4tL0P3wZZ6Bqq3X5Y34e+1Aei71p0KkKNsVMS/I7laEe45qBAdqYaNIXBb3cj
LQ9D3AQH6js18dD/aRBYEE0uP4f+Aix6Ec4ckylT1jrfWmyCGLyCxdwSVgxOfvnw
VuFXKzOCghVk85mSy55VFLw4zKcyt+FR4H6n8DWcoAMFOfg1ChtU4npKT+p7j2rT
/eezXIGqwaosOgg/BottfD7GMpB9TAPP5soYaozoSrQmpExkPfk48787AIOkJdLe
1jLmHyLA9s1Ku7ATI0mBL7Psd1YMZn0H4A91jzsSgEmXh5KqpK3RdSWwncd3fb7A
w154dZtYETU87QJDkk/QT3WGblcYvHI5nO87IYkXJKZRbdDBYdM3w0PAWx7W5zsX
GhHLAFE7z9BmmBov3H1B0ZmVGLOBC10W3d6TUuMrW8W7eUMFzImYIvtnHkNaDehu
LFiHH3plmFH61uVkcMX11gXXmuGAT6FI0RW3olfjxyfcr20u1BQjPikaALqDkIjp
LGDA827SND9Is2pRRdgHBikjZitbOP1UNNLAf29Hg9sYVr5K7Hnj6DfQti+EfGW7
0ndM0bKmjonVTwcznq5vaA68XPt+I33VX6+zrqNGMD1hzn5DoiKVPRF41YzGB3uu
2j6QmwwhsNHZKJ2O3Tg+7bvXedl4JOQeoQTmv7pCZnLLpVBCryuXiu6eNkKOMdu+
FNHdC3Y6rIitPju/w0vay58zrTb7c6z4oURuhrtqveETUWLb/pG1WpAaj1mY5Khn
7rg+VBvKnNBRHQ4hcCHJCptSdSPpdVOXYj9XREM4zDSsC4XwJWt/FOj+dnNu8Ug6
mcb4BchNqQrLNrqf7p++ct3OASd2Uw2gsUJfcKA2PalVVMWVKvVL/I6jau6od+ZT
N/Xodf7Pi6h46d9CNlACKChpuGfmkZXdgtDi3vO0+oCEQT6d1Nf9U+m8cM4xeZUk
h0mCEn+zTorWqE4te6in+B8EV3qM6u7imbIKfWwijHHXYUHlqszopaZVuTlkearh
/92WrKER1ieaDCm7zJFAxA82AFw3+2QpSdEi8xTXKvWwC7LrynoPikkdMtPA1aaR
ng5ROLWOqmiP/RbeIqCkxGiVFzmKzwG9WQztj7Vllo/5/XYenRz5mI5WHtlcxwzz
u3jJX90OP9pxMlcyHfQgKB65+w2YM0hm+BHEvLg9idqKoZEEqGPRIDTZGyI0dRQg
K+QBDOd3ifiSxDbHw3wBKE+uvFpSv0IkoX4ZdkOwa4t7xw79rzfn2H0CmDGPcSVV
xhWfBeAZ3L0ZneK/uePqvol1Z42OAsEvdZ9hCKWsrMnNrU+63l9QkzNO2lhjkBHg
gfL/B49BxBhT61invbhSUJgpJI4gTEo+4cW3YYwLql+Uu5ahtRB7X+bIHdina/oc
6RU60FPwbboxpK8H/bzKsf9DQ1zWpFIUoRERPeTfmfe5E+5NcMmG4Lt6o5Ky1LzN
nqZ4UFO06/x5+x3XcjrOCr7m1NLw6/n2mT+oS2Ek1Xcc5VD4AI4JK+Au10Geb6Ob
GFPVD65k8nC/W8QoJkGYvbIPCR6fiEb+4XjX8nXrFj0I4kuV8JijO+YKFL4ifWbY
BID+BtCUKj2QWAdIyErPFwJyLWGtq1Kg7qOS3lwlOoABNOigw7Xi1Mnb29fJ5bLg
arWSJ+fLKoAKlLFoBm4G/jVr/XE6N5dyRkCRYHtDqyTMGcbRftItn2PE6qR2URVt
LI/Qda77+mHbC1+vRrhyvJGhQ5ow2vxZPHurB3vbfMArR76O/S9EG3K5jDy20W1S
TeDtXwhegihe+PvxsXN0LeTjI+VMyInsOxrrH3XGdbPkoLnLyoN/YwRnbOIqkh1V
BmS99GFu77HIayelLThHaHqVsyz5XuWh3CVK6DYQdrlW84YYUcsDc3cG9+zsQhmc
+n38HWEdWJvdFhk+bRuD8ieOpa5QOhKPvpcVmo9HWELFNBFfKTO4QlH2JAOg77U9
6ofnWWhpCaEoKFIFZSUijNx2ZmLjRxPlp32GU/+orJ0FbdTAdoQUnGWGjsgTpKhE
h3N7vbIyIwrixQ4iu0GcVK3LFtSF9Ol3NsevWKfLTvekqZNigs+NI/QcOFqOW+cV
p8pFRDc4TWkMksVNSzyhr1B8ZnEyNAyEeaqF9WA+oJOSTrkghishViBosPJwKawt
kBrqL1WT9AewCUkPNXEeZZm+iRUOLekT89bVxgH0yLY2uCJU6wPgNQtsFCx2Uht1
iPpKcdXXWSrM3R9cGyiUWX++1qgBHO1wrfkJjo85qz19CrVaJoqDdonbI84IP6pQ
KdCt3+aESItGtfAsUvtNeuZOGjQJZLa7SVoPJhMaT6DTI1dHBIOrtVwTizVbjG6h
a+G8eMMcwZjuQBG8notlEcbgIKAOOCc25bMwERUORG61BILPMpGltxxcoweCVciE
8271u/FMgGpKlT2NS/CccldaAfuthhSijXnfSZtS4aIU1a/vSNjEBvQnH8nkD4yx
X8jEaug9MhTgh3ZfMz8eq7c7V9d0/5Ehj1SQV4TWiGJf2oJPP3RKGH/uojH5rRjV
s7zx0hy2nh0SbG7a9POidd1dF8eW/m7A2v0I6fsaeZCN+1Wg5XQrQluPB3crOOWm
G0OBcpfpMCE1k7JUWoxULFnjSns08t5TUW87ZbxBF8VZ7f3fsZmoqDXsPvn9U/uC
1yyUqVvn6DvU/684zxqNwaHUlXFM/Fi37yJfrkR+hM3DHjDDgZ2WJ/yL+gFMH3ra
ytnFCEIowssSJjUmbWvcpEQDcgxJF7lGhJSkqiGEhUJVnY6Wg3surgiXi32sZZ7Z
GNuYukQAUez7f9KOCrFrOHTMslZ8TtcdzcRTAMcBHt9uv8dbB09i0My9gXAT9CCw
EiDTGNoT6IWBkMroWzsIreF/Piz+6r+l9ymVFeF8STaW8g9A9BVFDdLPCiz7GQdA
OZfAoBh3p10dp+SHJpGxYEzw6NJ6MdhcEkGJhQgJQ+5ZtIkyQGzUkGLYR4WJ6HFi
nHK5nf6EWVymtM+64LdFG0WKNjwxLC9ZwZg/EnYfsMzeWlAZ9Kqzcert6E26S2X4
oBqbtYiA//UFHxLxOA4Z9aJUbloOzekh/yeU/+zu4XsXGEqwV7/Emva14EzWoZ0z
lhHxW1sCpVV88YHyrtU3zMXpEWz6vGFBRvf5AcepvThCB+or2kQscTxn3vp2JR2W
iAtdrywQ98QnwWK3vl0/rRV9mhtVsZYwPT5OQrd0xIo2RxNp0KbTcF0SHLSN5mFw
G+xyJ6IYuHpQnNEzp7vzQePY08g5DgaVyRIWfpcz97ljxYTS4jREb6jVb3LHuAOF
addWw1VkRtAQwHx7r5EBmg/dx7S1VELtpDiRW1iGafihwfrWFcVTMj302Gnn6QUI
mhw0mxgUUtqu8GRyz8W9gw2M3FnYecaAdeIFwkBjg+mpjLS3Lv6sekWVhln7bXRa
da3J1jTDZzi3II6T2MzIxOFWOTKdDkq786MoWF3P+vRo4ediungLLRkqjPOlZ1kd
TmcxUfDq2+glJuy06d/m13Qv051nfY1cjB951CBKJFueqffW+MaZVE2yyYm2dsii
gGf4ESFy23qz9sCoh/uUVN4wiMsotS4/8xNkaxhfJt5RCF/a/oP3y/f7z2jYlVyt
wjhlCUZbYnzfMbAVPLzZQD1FdzjDUEBYULVadi/FX72uJIAl5dzEI/P2vLj3MTQl
drGjG8/In/fUSeO0RR18JmzbzVlNiJyF6IHCTRkJLi03+0S2l6Jk2IP//wGjDZWa
7EF1YntNrn5JQiBWslkuzHI1BWXF0gO1siGy8R5uAct3W8hKzobofzDCS6MFsyVH
Acf7Z3tNJjMcKOfwxmPmti2P5nl4nThwWhLXlAZB+tVsq/kRGw9huELHh0BT4p/D
pPrvOfYuWtVqyoqoDE7OOLH+0qytaz/MaAFvtQUNc72xSfE/a/nsoHODFYh7iyKb
VJSJ9sVLImfqcWsI9AMzqG/I1olItbIUdo3scbqbB+d3xiLCGkaFPgUmnI7nM6yS
V8fLnXLrI/VBlVTFdWfyGESdFeX3MGT3CKI6n/6kXfiprBeSy3Tr9zvKU12gHugx
85HWQRB7UaSmUyiJXku7hWVetDewL6dxCUNVvBIo2buavM63q4xyTC1X9BsCPIgp
zaSZMeWBqyDEh5D1ZUfCaKeitkQL7ae4s53d+fZa6P6oF35J8o2X+3DV68w3yHCI
vQwDUA0kmVjWDfy+BtKA4aFVJaQikmRaCQEXKf0D8LozphA3DCzT9A2n4XKQd7Lv
gAizfOGhR+LoybdQJQwoJUEv6IDoWqxK7IbRZdoWCIVapi7qmeLd0CSfFm+Slise
L9hIlFu8TAKUpkqmReU/WlMFnqpVHIty5+yqEz6xgkX7Ar4tv7cZLCbpMrNMVyH1
efSd3Ct4CSjfzkFEyjb8xxPb3t7bfedIbhqzqMisaqgDuslqPSiVF9GYXW/M9fZk
jB0yAt22mJeBRYke+6nKcT5QVVxrEz85tlefOj2ta5koSAq0Pfx1WsMWTweaZ1yg
aJvfeqLZ9tjJ7NPYeSuCLIenn/tt0mGakyZQJofixicwlLuJc+pSpAL/uE318SQa
r37MLtjHk2Iv3kQqoutgNbfVYz/qPYkOSh6HifmcW6WutPneYwGi4wXUrEPQ7use
ILV01CzmRGSZVtUt9/FQB3ZluCmtk719ZlEv/D4CEVmTPz7eYclWEplRyT4WcXkt
s93WNeSCjn2Hhr79SalI2dl+YMdImW9xB2uSXQzHd6sPXLi6vAVOgZGJtCMxUGDg
kZ+SsnHQ1lX2s5BYxa6KfBqovj0f8pLky+aB7LSpQ5G5TQOlYl2BWgabWnz2phvs
5MjDgwcTPjz/905aEXdsNVrI/EPRZcbZELtonWw8x0kXsjiqc8DVje8ehn4XHFX8
khLLQGQeFsZACrH6hw15MedMnsSF2Uwv1NjWgkMGlqdrrYf0D8b/DF946kThkOb5
xnB1QNgny7tWtV0Bk6vJ28eE2IfAPhiousDLWQWHDtk8v6WDROHfj46imV2G0bBR
eEylTyQGrc7jEW9iko7s5gpJ/42aYIkyUFL3XwcYCHLE+OBoSa3KYRZ/Ki1SFx0h
OPIv9jUKMS/5d7SSqCo444MIEq5v73kkIgDV0oPJfp3WtlYU2cYrfNVO+tEQA22L
JelIY0sSt33ULobry1Kjt9IjoTtNzJROsTU/CdpZJ9bcfKi5I/Px3BLXYhzujVO7
5ZnIFl3JgY8zFONJvDM29nKttdXQ0EB9Exyoneq/r2yve/53L2HupZthagP+K42k
CWIunC6+YGB8/HIzS4Ia1vmCZ7V8doJugUw56FE6tSaj3A1rPYPHsdUu7c0ABEtn
kW1vVCLHR/onul7DNalIvZfJy9jlsDaQGytp5EYD5yD5aSqzuPca36/xm6MPVvQx
hkpyWqkYtDHp0chHQoVTd8ZUdfgg2s/VEkKsgdTWeWzWAWFY6nzHpDqsWq/XRLp3
h24CKGFQ8utWcOOgQ1+q3HpMohrhx2qcAbqcVlHZ3algZDrFRGQldv0iKV5t0oe9
4J4gnF2NZQSEUqtBb2LZKtffXAjNKFEKCLAW35saAnAc++tsYu8hFNYjumieXztV
6/GP4tY7a3Jc77eFgIIK03KAUTUZi9ZukPhDnCwrD3QvXxzLBa+CQKnB2HbkLXVJ
ZmKjXZa43iYiV100YikneqLFJK1tuDXSw+RIdJk1EZL4fJsRxxBcJ+TP7wYUvWi3
EXgPXue7VUKg3apHuvogKUU7V1K8Vp70vTIdH26jIz5FklWHQ8xRhwYHtZxqiauT
h2ly2iG9hfj3yE4OM3b+pVh5VjfBJTfol9Qna2p+YhK0fuD27GL7o2sNg6wi8QjT
f5FZA5jfQn5kNHdUpWQkPL2sRlAaBt3tGgyYOdatOjMkyGoVOarDLgArMp/MTpx8
opBCmtfpAnMexv4fXGZei29DCCaAriUMihuLkpTkuQuX2Nqd38HDrGIU+sYGk9Wv
zvRVZZ+hUMlllFKFby/8q0NPEKTbZF9kVev55AUQ/bcauRiAWzAaA7D47MoOr2EV
gFutE8OMuo+31eTi5PMPGFH1nW0J45E49Zy1tHZluKRW+u0k4IxLlPvzeEqZfjhP
ed72NBX2YHICBJUCeoJVK+6ryt+KLzRlRD2qpesIgLGBFMHKB0fpMyUSaOiQiVEe
qtwgHegCRBI1ujYY8t3/jzPfm2sYQZXZ5naZepQ98ZGUwlpyfCKbIyEuJgwu6CNh
9V2HWdKJjcQ7YmqdwSLTAtdpO4X3Pumkb2tYiwe5rBtWImqSEJ4AOPk5rGTbCqxG
Hx+oco8kXPIA5nXuYZrkXituQ+qfRvpNNuQzWrveLxEtqFaMAd/ayqCMj+LOiRhB
jMqvUx59n+nGoZ5b781KQkMvCQXkT5aDBgCvjllBqH7eCAyVb+vRDcULD+F5zIrC
1u02RudJpIr//cPHZXEoI3jQsmKVP2AXiTWWCo3WfvbVOykxc0vzm7723DZyLTKA
rRaThVpAlc9LLYC2Qei/k12SDe7JBcBEROoUdNNRPFjT3YmhlSMx+/YicsLPHxZT
YJCJ1/tAc4K8XJPWL5Cy4cR3+7kB3ZN1c40OtIYuCETushh7idnkDVEv1vGCDSHi
BqXj+xqhs0tZ4VI5hC9peTD2Nz0i1iWpgRgcGPYjIfLPaLpZskRePBXDoUFntLSf
qCkiTLxlxElJ6H40t5mW5d9F3GFu7R2fbSmiXL6ZjCwDB0YqQvyE0qjC1MfYNp5j
rLqC7ulBatCZF9IYL0x1tbZQTRbopg+1VPmSkEBQf9JUj2Xz9ykU9JDc91LXCZ8V
nOJU6QPvNAdq3lQoUMTtJnb8Q9qaD4rbziTdkl/8+htan1rTMadsl8QmX3ZbI4Nb
ffJ7x18OhBq++OWHxhNF0r6IdHmVJ8q0DMrXFFmwXoR3U+RkFOSM+oGurlfktZKz
rtyCYsT6rxLxMYSW2IqKntXg6tG817bQfW/oS3hrIZeobBMaiSMw9+lfMjlgMZeD
vPnrR01KL3qm6/MhQQt4OHilii9tm/sa1pWwPTNPLCkBzOmC5SDHwaLygPwFnPyX
S2fs0+RBFNXJokvOqQ0YiiYUPy1na979J1bdMtKKlFLxB6L6RWouLVAzmZDSgYjM
o4R0r7ygW9cMWqDKtyJjFi9SNOvYkZDY8CX82IXOLdLz8kuM3IeHcmzBLkxe2sbP
qieLIqoq5HZgq4XF9Pu/DxQu43tKsjUs3rZQvOrsgvtYkG61gTKPlDra0AF6CHMu
8FqvO+CxcsvcJ0KlyOPT3HMEZ46CR1j//4qqQzWF/IJMYI7U7QH8wKlQ+GwPhMBF
NLVGncoow9Vm4e2nIZN4aj+XPSACO6wx5MQ7wVvXzwccg/KVxvDw5V8Fwcm1cAnu
YDiVJn5ZH0o73T/g+gWMs5SCVhoBWMRIj6NZspMmTDIoG1quTzLBz5627I35idxU
YNcOglMLArJDmtBJteXUjeHbV3VhNebCvEfgOz69SfaFN9vT1Ev0XBw8FojCt4Q6
aB521RD7jw7PuTlpGWnBQCGqb6RpLEwPytkCAcXBMWnEKr0monSVJIRSHPpamR3V
1qa04miSH/DYtrppQ0blS45KyCdCWWiTalFtuKU2dEL5R6HNZUd5WagU7uz7Mo9q
nl5saaGtEBGZgFpX0YXNLL/f1MkhXoC+WI6AWH57jjBl2qQ1qHM6uy5CNmWnYMGR
IIqXbxm5QOkF5ciHK80ZuxfrJRH+PMq2wnevLilvNN/uSLmroRF1tokE5DJbMe1f
608mCha4mB39KEqcYQeT3wDFfQsQ4cwdNuDHRXCDzMCf/B1qquSQrSBFEMw9J3f/
UTEQyI2eMgvIsXFXszaKqbI/ieCEXC03FjCGMkoJXNX1VlgG+N+yvyVi1oChjRgq
nBS7BKdmMGsjqWFB5AX17CfACiEn6+oe3VApJjOM2oDUvmt34Cvb2+2EAPhOq3kL
0FOSAMVXLnas8ldYyvghFXEP79Xb3GJ8gLvsRayJ2725gWHrEjcuW94kJrkRg6tJ
zO1aauynjMuYSKAFGjUsGOi+gnhQtv225pYeL1mw3gkK1O7q4jarhDM45bwxD6Pe
bXrT+cvncuWJibtNAOjtMOLRe4Lv1wybCph1YpTUA44D+a9ses1zpAhIgumfxenn
M2t+mq83JEaSEmYuccX+A3w+ghYgckyye5s+kAf1sKfHu45Xs0Q/5oTlNibZDAs5
DkkOSADY7pz0gS3RDWjf2ggrCNhwBXnxaGbIQUsRsKFjeNLharvppL0I0wDnwZiq
X8CNCWdBYcq6P0wA92XpabWgRUn2ol7djhdQCrpz5UHHghg/QNr8sPjVwrHd+3c4
LYqBFDFIgAp8sVecElQCr149sk3QImQY6JigPFMd7QzRUJUcIR1k9hf2PofttguQ
1iul+qdnYKTbPW8q0N5jN/WQBIwtpy6jhtG4Xg76ZxwkxRndBNnHarWLuJ3QhdDR
Sl4+1NMBLiQs8sZe7ikvVwEZmDYfj4hTjINRcxhGI93KuyFUDrjrtmlL3g6TcgxI
AzcElCn9oXxQcgUvnzYk4VdPJFIdwYiYw03REbbJsdIengX+MqjtHO5MvivMUBsz
UKH74TFtNdz6LMSlw7TpBJ5mZencJV6kM4Hv1yutDWP0Xh7t/SlwHgKGHqjHt4Wf
f0v8IxjP6Ryi2sV2TcIYJscT/3wbDX9sXYXLP0eexfq//Esv7yIeady0dKUDeqXr
pIf3mZi+iDnFBlIrBSvglGAAoEMuyZR62gEDMXsh6Du3tfpWI4y6bpOmW3NVXuqB
5jVbBlT4wDxJXyxuVtXpTzwsA4eB++JAuB/DGYLEgmQeVI55X6RW3LzDW75R3o+j
yA6x+Q5fzPrXwGw7HQozFVdt+V6hjUHIqHAzk1gKs4eqPh1On0iBA1iAqgN519QM
xCRcIoB5Smz+wNq3Q5Cp/AT3rY9BL+At3fC0xcOc/n5MHdr4NtvAKH89TZ9Q575W
BvAAGAgsSmGT5Fv4o7aneekBdL97MJ3LkAE4gpkf2iiojITGO9yrYGpRwo11ujFh
p9e026zpNfA3wJwOA96Va+vUDxtPrHZIo7mJ82yr/Zc9M/APtSZ1dJyG2igTjnWx
DRmDM+vqEESOmr0uuofIY5UNJCyMI7E2LKhnnFXDpqKsv91UWvRGcaQtkxLpk8v9
8Gwgk1d9NareN4/HVwHdaIcuRcKXLheUjs0zVPTYE2wdk/IAGbK0zUySVd9J7bSU
z+SPt69VCXoYGDYzdMbn5XHO/Sq1e2YlMNsAnSvn1lzEA70AJNi3mdUU12GJXrUC
SuRLdHicJAtBFr8RC6HGSOep5sFx6FQkYcrS/x5WQRCJpycZUZaoDk/tc9niIa33
G/REghiLb2Y+mTteCvYl/DT2q/uk/vhLPei0NDzHI5LCsrDNNhqVXEB+U654reum
pu3Q6cVQDEqaUNwHDnM80AXrJf6nRCgXUemEdLoz9HX2qaDq/ptD9ZyCwDBEKL1t
rC553mGmAsjJSLC1E6R/xbyUrPo7mt78GQxsECiI4cBRGfx2OxKB46j3VnlAz1ZR
R75x67WtVp2pryGVm6BKmsiVc//8EtRyjMJcL6fRRotmLbgBgrEdtKIauQfyezkm
lsfwt46LQx1A82WqtnZ9GuTI+W1kFmDrb2XVcb3mEO717nMNX0WvwSUtZK2gakhs
UPz/G/ay0BKmliwmhoc3K0I4/2s+eXsrFb48QhRcDuvGDvJHG7KS4G6RO1QutBtj
FwhJgg1rXIlWKRK90B+K2hNA0gsUyVJN5EV4h3uJRrczBPYXSXaSvXzmEkIRVdNM
ZX9sMmcQqB+50wgVvAuo0xz4xkI9pYsMsQVfvSikxHRGVP2c6HwgdHdgDeihHjs0
eFgEXlAtZeYgs24XeVVJ+iMgHuajVV8FqJeJLZ7JVfR8b4/UajGcP5PyPsJ42Yk4
AXXtCaWRy4vGLXB42ykz4PCeqbNReqAA1KfaX1fyvnupUnhx/WYUMAl8FFGap7zK
RW4bqZWgTHTb17DfEYsBGf1c9jOBINEnXcfFeINPeVXJxpPUQUkyWWC9aVE4L8qS
4u3x9Z/MZx7zpY3QhHtBOemN5Xbt75nmYKUa1Q7Dl1Rb+IlYI0/c3uxw7J2Z4JgA
YW3MFy7F/X0vVgX13N+10xuMW7KVxiS3fEHtC7qMI5S8emfxtnQQk5QrwPBk1H26
dnBJum546KVnR84lh+M92pjX2rLh/R3fwMtLAI5qj9MYC0GErlZo/k3cvbkQ3PrD
b0Jq2oJPz0APjDeOxyycXyk1K7aNQrCdNAs+RjnFJ7vIGdYDk3q2j0PtRAF7S8/C
339e52ua21oNMc/qNTUkwuodI30tpdcAZNfkyHH4wyC73fGA9CGaWgGuJgHw053W
ZsF7GxNZ3ovnIRzLoYCYwH0GpgxQZQhefWcOkOKl/byGOnwEwUUWWgdHA7zdVIuo
6l/tJMxnmeDXpL8WIqvRSH+5xbCvc71AUvrci5Cc97dRO8Y6BzVP5Zsti5CZjLGb
LGBQciXOZXTaJa0thMHMJvfY+KgqRmFy6kXmUVjEwnTGEkqyzsp5zhuYJm+3HPNU
D6stBywnwe0epCCpQvwHeB/Os/pNwYvSDJbvKmHf/Wn8ft+qlsL7Fobp6XHRu1gZ
xfCX02Y/oBmxxwV44z6Y/dHMY+wMi0V6WVX5OHl1pos9dNvcFjE1M/i/jR/P//Ra
8FTLtCPg8LBF1Zn1y6NP5mpGtNOZ5bm/mtxtITz53sx9YuGOLw6Q3l3KHraIAlt0
/l+RcxgILqPMJ4XuGBmRWeRjLOWlfTn4ALHzG79khF7l50Ou/QfB4dJh8RfYclgB
/mteF6Buu4d17kpmQnbBIRhVW0I6e1beZoelzn0tAWWHk9TibfmPsOrWeoIz4w0t
xeAwVJnpKOPcPW3daqQlniyzLdNSGWK1jPTecrpK2g2r2dutt7hmtBYdU9TJiGHH
fU9PCKiM8GulkMcAnpf14bDbm4zgTrLhBJqpDpXdDGz/+TF7GYYuKQOG7PLmoCSw
DpPWHZhHgVgbJ9q2f1k5NZcY69JzO+y0EBShtwJnteb930L+m6l4uare5hPNsWVh
Vpjf1I0tfjuqqNL4j8+fS+0cZAV0l9lMfR198LD/T8WoszfKCH6JZQUY/YM+dGRM
f4rFjFLLMT5k7Di3mECmHVRnvrHyLbv2Pjc+zGDup+s4t8iy7ejbyPRt1vwlwxrY
aB8E7p/RxyxdMyrXWND2+d49+wcuqvWvhzI9n98lizUHV16A0kdazMIN8CrdDYTT
xjfGw1H4JxzvqFEY7Bkw43OZJcv1NqCaArfnKAKthQr7BEriEBeVqZJfC058eLuG
8nFDnPoFxeCK49DzxTrkGn+kqXMirEjI4XaUEiahYl7gC0l0WDmddVtJGoKiH9Si
e9KIm1YotUaX5tob9tk1zyYGV6lbYHFC16muZvu2qHeIue/JswZvt03/kUp7j5tc
JUrIw7h+iNqflma6w36zOQ5VRAWq1ZSTPBWIbspvrdZ9F36w/gxNYW39dLMwWCBE
BbdmXmpJWq0iw5EY7qxIIckJ1bHm5vpBeLPrN4WyAAvFDVzEzSVs6UsNEHVivjDg
+bBXWThitjy5dEt9EcUKvbsClnYN7OSGLIuN0tVeXvw6sxJT+4ovkLOqI4qrNqyj
A3mXmzMpUiQHc9QiNdrscie87saADBi/yWzUyjQtcI4Sm+m9nmcCNxknS/8K0pB7
7JQW3P2V/5BhlIIEL2QDcaSF2g8i0aTgyJLxN0OdRMamw4/SKgp1XRPiIpIlLIXX
5NvAK0jyAF4y9VA7SFF1qqBHDW8RdyK3e/YtzKF/7Dj9e8tetKhTEs/eG9qV/T7S
hci8iRCsbI0t8Bd+LM9lL46qNU+LJ0eHAZhMwOCE+tcBrDRKDCuENlng/iovtLmR
8An/NGbKJ07tfWwWYLwtmDLD9Ufi7TwEghcETPKXIqqd50MCv2LwHoHw67dLMS0r
Evp3143BgWiYxR1NDS8xxP5FfG9+ic9aGo43aBJ3jJi5glM2zzDHsjZsIgGAgMI2
q86WR4nxsxN9uYduJmfIiuwu4zcI9ogq4JxO7EH601ocBPdwhTR0Yx7U41uDXWCR
Y4BA40vccBECCGuH7mSEeuqWegapEauO8m970GJtv1q03zQQG3N4iWuuEYkcVSY3
yF5KefNRBCGQjFfoyiM0KD+cUapUJNt9CiLyLHSzKiJCSTEQOI1UBpeVtC3EjjJX
BgeiIfXHqw5dIy2whH0rk1ml77gDIZWaN2Yp40wD8mcYfFp9tTEX03UaIruxCWZF
cfMRCH+ltPnjYn2m9jJF0fLghZ5PU0IJbFbKBWorPUufG00E1rj7KBuAhkIYC4tB
1PUqjmWxxhAxTaU6Y8FZ+novEE58n18W3hd/Ch2qoA1ArjrRsQ9ZkwRLKo2xDplh
R137l7X2q1iNYTktiGjPMTINqVkhNq6ULmxj5XiCD36ISjUBoVOUZD431dn1slYc
kXVx+vMMOQ/yrnqPiQpcH1xpg8Fu0MnjoqswrGIjERINmq9PYGG8G2i4nJY1kkUY
q9BjFRcaGd+Wwo2gcGHM5uFtZscz8M3eejcE6jyB+OXT/ElAjMaontPqHrm7SImO
IOT+/36d1bbA0KFJUmq787K0WTEFbTlyn1qsXSjji6PVYQYrMCDVKp6ayoZmyC+l
WIpdyvDAhTXwj2g1WtLa0fcquuHZz1noORrkOshszd8KlMs/GZseBGRaIdv7scC0
JZnuUuwN3Za6AwukwTk9smjfKtWmBw4h3dD1Z48BU67LV88UdacE+1dtGXlcFkhV
+LRI74TpnXK2nZTglfcBqWCy7A+wXdiGc6sWeaft6aknfX0vuag/ytQb1ZMh2q4D
DNfoDi48FyIWnnbm53+N6g6c+ATdDuNolNybxdnmo6e4NEhAHjA7/bSvG7c8utIV
wwEfaCy9QiGwpchOdlnQU2YhoEJveQtOcLT6JcCnhGsnZYsNvaxj7E5Xf4QqN6z2
ikP/9SvSZOp7TqjaAgUL53SrzQ3SX8xT9Shu1Cqyu2DFFzzDGZWoKF/4aE/uuR9x
Bd4ckEPvj1839yfbYSXYc7dArdYZOPR6Mfzkvm5nJFynBorHZnv+XBGy+DDgMmLm
rnMDtoEYnjlmULz1hTn8cBeAtg2s8VIJLMrMgvIJSWOmm7gYilW65wvWCnLkcS0g
eUF/yXj0rFczmN8H9YJ5L3ouRBZp0At6K24JfCtMgbfITOvCcTF/4quRCsZ7+81q
Av/tBfaxPv17ky7bkhuLWjn1AwrKmM/Hfeq272ZojzIDrfSa472O449HQRGSGrWy
c7S3fKItaN5Xh2OMsa9ZFPFOHILx0Kt0cfJFpkAJHRJZUBVyGTAKJ0+zgx3qQwjv
N7/DLxZbVmHkWdU//wRWoXcUf0+WxCNi012TLoyBwObXYk53LtUkMCSxQu1Wdp64
tAmC7IHmEb7lnSYiV0nFNuQKEx+6wjRwQWNyfy8R0oCvds1XEjXR8USIn3u8j24N
mC7AM57UDDkLJdbdm0T0usaDJEmS0qnZlAImgRauhP3ZoAjFm6635I+B4Ql+sW6s
IS0S64KvlmMaJtPa9Bxlz3OjzWQZtK7WIhyJNoWjdU+O1j5ISl/4SkPCgFvxJkBo
zau1E45c6M62DgOA2ZkwbjxDGjqoHcjwyZWB3CQ9bUjgPeoQ644nK67td1JxI3vQ
VrmL/SKVxdCfPRvB4PSsJW2ilUo69lAw+WBLU/3BKSjDxW2Lc8akXSt6G3woAYFt
tilQewCgCrN5tZfkz+q9TJNGcK2pkOFIxRpyLaIXRqLzUi0znu74c5rgQXFQkQNy
zUkqkAKzuFsXdHIX7gkhg4CIlaPaIGKO3t2zhnxeDG3EI1LZAsuon/7MecEA5qmH
bK6BPf65ELE1vcZck9tGqbliT5RlW034cjI67lNP1M+Q+R7Ga+z5l0If018QqDlj
n92Nt1I3oIc02AjkgZ9pZj/zXsMogJXf4cS7B75gm+ol5OvejquD6KoxSyJrTXZd
OLGGuZU1/0HZYvAAXweh4khXd5Qj34MBnz2aRTVycg9uhk1oBS28mtl+jrMnglDy
i0Xt0TVZX4txDQmekB1x/FGU7ZsGndrC890EsOMg6A2xccRjsNDdT864ZQxL1aFA
wuFC4dcptqX1MDCjFE6gGmsS+zxAwl/kkSVTY2RhyXeiYocc+E7hsDqqwqUmoK2A
oyj9Xcr5GCy4tD4iSPElvDQc3Oz0k85AFo+Xvabzymce1rn2HPa36N6Z6x4uDTgR
AN70ZDeR5xbdh76KYAFEL9vI3qslpEJ1mlgVmpHS9FoNNkqJGlPtpuy+1JbCMeU9
3/V6LOjW3q+R+d298HwIHWOJlilRZu61RH8hAdZB/Y3kIZO2+HlAj2k0t0wk/J7D
lU8zMy3UFOKXlgSJiy6zNnVEoURW9ivRwip5UFHWmELF8KMgRwJ1A/kJK4+IZEdA
70rgUx0Nbqz60jZdQodlSV69w7X1ccoDE/UyPE/WyvigY+Aj90C8l9s4ZXgzeQLi
6U3u/fccOX2eAY0ycdLNc+DSgJpNP33yVaX/gt5XEfctx7iaV9G9DALK6tAHEfIA
y0BWOcgstTXy2nTs1PDq0sOSvI0cFpDSind22z7ZnCpDi4IXmx397jfnMtjsLAeZ
Zn6oUie+orps7xms9EyAKm477hheQVE+UuGk1f103ga4sjgCMb8KK7KUeUFs98hp
IwE2wHwACqNWA7R3c896Qd643E63fzn0pZEGZONNDAGeP9ZM+ptJfy/wcA5vGkex
vvkSmXrqu11DVcmrqGABC6Tk8wT5Z2FkbZLBh7BKOJGVMrUgDkbfWmRQWJouQ+pT
Uo+J6BikFshYYrv2tG2poOQlz7IOu8i0gTbf9pM3MKnffVQ38Cadz9gE3QASBHW4
by9fF+Ypx0F2nPzTykHBVdRsmjeVXzT3FLsx46ZEPI7ZAi0Do7+smUf/yd9KGSMF
svNwoRnCNOSHXhMf8SZ1pGVCtHm+8oDeJ8GqKjR2gWYGlCeryWRj76aI0A+h/paP
Nznl58gR2ndF7D9nmOaVHlc1Zuwhy2YLDa1fU4yEj+cZYZ2fn3+OgTLOsmMVJ8iC
VfxgLm+fTzM5u1p5QKM02ffsmRgOB6KBrj2KLSP/Dpm+VWn4yjncskJcNpROLk6W
wHs3l4zFf9D/9+WKvc8f0nvpQPMEUS32P1kxj/3dJUlRBgMMiWkC8S/1w5AQttLx
ESR39hoXiKEtWz5EQ15IggwTiOHg1LgRaSNeMF3qRppRJhhPfYnCeiIDSO2mjJ4w
moTyMF6KXcUxmymgB01Bn1Tvj69EemSCP5cqMu5QQWFm1I6gg6DQ84dqtUe+Pbxd
uxo8PZqTXQCMY14DxzKDz8Kjp57v7KkC/eBf0E3npuF9CNHncOSyv2ox5xtXvmAs
DhoyGCG8MSeQpAFqxR0CG1X7oU8UzcsesOrY5SiLEXUoKVZ70Mv5a8dwTBsih/T3
AC6UUxt79+9Z5/WNMaoeHc+5yA53B6muSHC+7ixoz/s6RdHll46hZjSw2vfeVYm2
YWhATPd9qbY2jXmQL0e4aOeqfwCmPc6ojxq4kFSci32QiuNaq3sYEys8twwxVpCW
tmlpqw7WHGTfkS1wQRN1SGCJAO9yJZUUNC9SVKxRzm+UsGDtmFcVgm2lk3//ofEv
Bd5Y8tVNat/ccvzLBs5Lt9Qb6KLntgnDkG6TYzIx9J4+SaidpoTQ9p12pgnzDHpu
ozO2vE8bnUJoQ0qxba0ut9V+AH0h9hC2VyHmEkkAImV9ElCxGP+COhAQT50St2eQ
FjmtNPz/k/9ConAOJN2MIPFOLogaxVMbua1IiVyNolRzD2DA8d+Kanw8Tvgwg+aw
aAyCPbJJk4GPghXU8nf6MvZmUINVkE+EFhdPmY/5D2PMsjTAO+Y4mSdgwF5/+ppM
nMv+nb4eBnKQo2dpdli4Hp8iUrCWL9aNBdEhc3kn9t6dFsrHALa4Ggve508H62eN
jTmSR1NXoGv18tJTH5fCbkoYWqmyBNGfPXotGgSJuBavupKJoM4vTNPV3jsaOGw2
pUq1aHc837OWOxP9DfuYgfjR1Sd6/QwEUM5/6XtR86oSGbpnMZA0IOk29hqNCCHj
/rzsm6zl6jB/eJkK4S6oIFelQMJZyFPk/nwt2qB5nJA0g9baNGh70P+NOPmJ9Zdh
hnoYOvf4EPQ6W1gY9UmEqzjxHmj4J3ab0oSNfstPX7IcWTg9Pt3yTg9W3Si7pjtk
BMO8pA4NG+kJMXfV4XHNgDlpORHmPVNInHzmzs+WzLfih7wHbM8gH1HBfEkHclN9
7t3OWyRBjdrNiqN3RhbNZL9nAVTy7+aJzA4Q526Gm5zqsmlL9oIZxt4bgKVuKUdo
A/3ymB/7d6GKJdoL6qQ+CSPOpSsyB4RfumzF7dlL0Cwo1pWpp5kEcXNS4Qxl2bRP
BdUMvOyHScH/hhbOH9IO8mmonSDJy4m/03+yBMVRG7B8ZY0/8dLuvfPUMHJwDwq2
FJJ+Yho9QKdys6ZaJSK3oLUgcZntIudBVTnFb2aB7lHLQr65lYGuu9k0pTjPhbWg
yNJF+yNFHMwjHKdhRJCr9yOF6Z8Y1zKycIvzfqrl3M6Dq+4mv7QOHSi+ULAvoDmX
uwSzMkPhhyAScSwzs6uQkwmqoXf5KTgFkxCVU0O0kF0l/RMhCMUMJlAsYvbGy2gR
SY2ekLUxn0JbQ0hVDGChEqv3OgN9BmMYIQFGMw53npY1khxaZYtf0Na7zTZoBodI
DqOBad9VFJKu4UizXNPChk7AOc3cn1xqVVakF9tw2Gs2im786DAJM7vRhhQQyyjO
aP6+mQ6ut2g2i6+f9UzNooOo4knJjsjxULsNKrjYYbZTYzIzfzq8yKMK1/6QE3MW
7k43G8uSamoOOvK0ezJwITHu5YbmiGdql2+//Hrd3HWOoy/EdKuds3/e1GodwBxd
BGoppxywAQ+zZQ0rjvgYwgHl5GA4ngCKHtuwmdmexazfRUiXWXUPZTMGKXZsZo+Q
SW6KeFRdgq3nwhhpX6FHqTHG1tFMTjqBgKPsSvS6NQVFZY+HznCcGz2rW+cZP8i0
xE7gSQ98vgF5MgsHTtWxofTR9Bf3auGE1ybhsU/xD6Z4fWdt+SAAEBCnh9CKZlp/
I7QB/h0I3d9N6FzKikZUfwrLHsRlT2BCuC+XePndPyp1b3JdxoN4hOqnD0P6DqV4
8X7F85TL4udleWOAbkKw9CPjwWWqtINZwT3Apb7Q/eE0+weSJRwDtDH07jD+RPmj
tUo7PFbfjO2kyRFMXsZBF/7DkMfRDiq8K5z+7ckJU92tkWZ01BD9tBXsu7GT4ht3
E59ZBudRpOZcQBZjCaHGlz/SHy9IneWKq+QNPTTqeBAvtEAzWq2ItgDt/GaOLGn5
FaJUMZ4y/Hwx/kpP8nt47SbSRj6H33R7MKyeAZPczAWCsVH23nX8y3uLBhORj2uF
iBzDuW0KCq25u4mgKt8eIPzTOx/OxUdkqZQMyf4XP9PLWlfyxJ7uthtIOzysVoNh
Cpm5eCBT6XevVgaMfiQDHWdYYUjrYZzB9/n0xi42m0wIM+HtbjPxoojOMoBNTx/D
e3SDrGZvItNvn7NGZvfHDB3aH/Dy6/u3/p+D6YglN0Mb9WvLkPPjGsW5Uecq/R+y
Vk5hXrl9rK4yA4h+BvSVwA6F7ekkNK2k+0uAH95k+i9miScY18cqwUrRebm1cnem
QZX5Xojc4QDmkFCA5QFsbJA+D84UPdwFGxq3yNVYP4cJrYXc3b4wY+ySfZxpUPyk
uQ1Pzn1WIj7+6uMa68VPPC9deYXon4800IP3cIlprcHdm0LblUpGvlggHNcV5Ull
fb3Gr2ZgUfmfucNxpc7V5e7fJikA/w+eJPw4mJPqTIqQSnPILWTMt5ooLzleWGAR
+c0vK5pX912Fq5LzOEkWaI+He1cV9MY8hDCqj7/urYUM26BrRX2idP29MJk7vl6K
SZab9QTAMUPPTqnMpsHx9RvpzpMghmm9zmRA0z7yld0dZMonjV0RWddZpjsCHEH8
yQ0RcceA49gHK51TU5K62w3WDOmj06n/jdYR6rfKTS8iombxeLVzoX4ZlDO4oJKI
MD53UsXutMh/dSFw4hH5vt1BYi/3NA8F6JYIQJXi+vsuLEAnTESQoHrpPQPiUjmq
r8ERVM+g+Niqi5DmZgohvWDk/LIlH3TjM2gqKnl1ISqmnAPq3P4bgzU0/qsEStPj
mshmdIYbDcGGZEANiDebSapConPyNWJK32dCMJ3CAyYLbyQcB+oaTHjBtWRM8c55
WMwNBXBXDDTzNeKd16f0lrZRWAQRkB7r4LYXYhw/wRQFN99C8BsJVLF3wwpXeKSf
e4Q09ZpxKgduzG0WZSkDOobLXzZq8ygAIb3ESlCQgJFW1O7W9YlepYQKXUZd1TDd
ZgWYyDWbi5FtZz1N/wxVzTDagndQQjY8UnAPvKx5IgfK85W+ydTiI42A34dA/cUZ
9p1SuqqN689KY9IhimghOCAHNGeiJVAgDK1sA498BydDpVqJg6bjiuGimpfX4dFA
GsTIpVajVKhMWrW5yx78VnYCc3gythkxqA5R5b0LJuVo9605DaYbJIylO2B11lqQ
RpplZEVN2FuL/Iq2qilpOPJY0ccJ2oGAFB8iDcza+xYI1ciTGG+6oXDAqg6L4FBh
H93rr4B/4NQyDjMP9Zr2/KvDK0sQXxiruLgr4j7xkTFAi9HTap2a4y84z6YiZZQ8
rcF3sRR77yvdHvaMT43sTRL4KdWM0S1oiZXOGdIxMyo4Ux3yLy/arYJI6gJoRNWe
evkJgAUN/ohtEhSyy3KvDLS/PwdStruHfso31T7fcVOVDGiLF5js4p7r1Yf/J6YY
vQbkje9bBx9tGavPZgesKVCumQB8neYb3yiG5/mK0fkZFZ5SFLQ+N2Qt2SjoPfoc
PB/MnKHp6Gz1xysR//xq034kKow0XA8CgI8yBEJ37zT5fDK0rQYvR1FPlx1iJzo9
leK/8s8JgAuUCyFvnB0ydwP/FViYOCz8lzImKDy1TG+lxXQnUU+1Vi3JdckaCdjT
48HwOX30I+wKOcBoxGUicNMrKELyyotVzhctivj17M63XLPeghTdp4g4r5l611qD
gWL8pyYYaMGwa/TE3+qfMrylAiLAG0JCH6TYLBTAPbVjxhsHCfhEdNl47Ya/9M2f
ZaRQ+E9EhXhQ6M5V6HHt9l+jI5t5iUTznSNV7ZAKN2kS0sH+Bmq0FydVU1n7gpR1
OcU2ZTHOCRpAjLfX4Sy/TSXk0iYN+oASPxOf8mWklsaPw3RtrREz9azv4OHHGk/I
bx9dwvcKYW6bvLaZZH6xdEYTIs3jCEAx5auCGHDbROPyRvmsDNPUrZCmYjKbZwSl
uS4736K3JIrOnfrAqV5LmZvBDOZF5VtKxwELrEKJEUZSo904AY7eyqOdttRV2Hs3
99VA9Xr7UQtufZfuQAySQRRP1//YjtBmiJyKNe3rjXcayzF/3g1AGu3aWoh86JWp
PVeNQ8jJ36By6/yukk5G4pTBjkNuqnavL5iE0EX3sTPUAomnIKu6sYIpnEpjCigr
iTOq0DNsBxuhnmgPtLHdY5y7fKAkuul9py1giZA0wm7PNsa0xGgp+EMl13a7rV85
WiH/OihMYKehXxmv6z+sDmysPOs5PzJ+p9X/YJ0JmIWM7/AsXsVcmrYKgD3FtAwU
gUeVjymQnaDtiN2/QUKn1QonzbmEYpfGROb4sZkxyFqPN2jOP2Vlu2P2pIsoY6Ms
jAXpy1SF8LBkGLdqIDHcJspum9FSUdQBaCCXZ+HZdi3xNB8Cn9miYlxP7K1zGdNA
m5I9rUwm7eDchqky1mZjyxblbGp273cM0eVI6ORlGdU6qUH131UFSCSUtikP1RwZ
aFH43YzvHhFXsZBUP2LIBmSeecUxMfMzk8yJH3JH7LBpCFDOsSzYdMgBArIfbRI6
VyYkSIWyf5FeP4huOb9e3tMZhaQVbdTusSXX/gxZtEIOtMKJtGCNm0VFSiuKTZUF
PnMxQl6j4tsC+KUPEqL4qooJjxKs0mL3o3QO4fyT65ss9O1q5eGCzBeYAimnuLo7
Ip4Z23l4kNcCe8NrZPxxa56K6nSIt9nOMOxDVZT9pDDm04YWpINYtIDRz5hDK0L5
WpWXLb3GhskzIOCeRFSi29pg866yFbQYMKfOauksrg4iLUrDUcQA/BV49M+AKBml
qUDWUj5RokMKCjmBRT0NqiyKIPmCJRF2RtKY4a6X/v1fKVX/gW3X3JjpQt5G36ea
W/4KGg+cBKWnVPJ/rzQYhxpc0JLCRfbG2LBGMo0Qw8phKQQBWdS5Xq+eScj2mhWE
jMk2Dq/j/1X5LJ5wJHzViL+nUUavfSZ7SKkT5NPUmn7Fs+f/jHGnXPPD4B9iuSjn
WEbUqL4k8ZQJszj3OgViuJPi+VKZjW9sKp4Zcf7iXkM7PTvWG5mf+cIclqufEajY
jXcupllLViZ0JPk2ylsw0CMPjtaHQhVzT889Yr2K3yYKgA6oQM8Y5HTJpYhHle4g
1+BJQReOGs2pNPoRPGfxmse+fTTzefRwFGJPQsZM73gwdZNf9Hc1/7qZR8D6zyaH
tpVMSeHgeEZ8KETrR22y2kQeRcp+kWgaZIzKFFxlPmwbk1RT7Dmy/8Lz58TCuKyG
MOQUZsU84r0W86oY8cE1ZXADWBxWq6DRL4wwdvCmG3OrG9ct0oH1qXiKqYk3JX8I
62Yg0pfocCkc7w3S4QZCuzoKhUIjW/GTzgwU31ybwSwH8XuXJBN1QqiOMzhcyCmR
ryDlsMxRCBnfMOYIReq1pEPFfpwxuiZgIOyNNBuA4VTfqwef9nOvt3Qk58O2RTfo
h3WKjZK8YL5iRvW9lBjZSgQNccxH+naRGxEX5/WClfEl/24x+plQPglZVlP+F3j4
gJq0+LnyfD/tTFcKB7YzR1qM1X3AKH4/IuqVyCOxED+Icd1MtCBYS1eGLF75021f
YfVXK7IYTaqeaZfiZ6Ok48zy8olosgiOBPLzqMRryUUjWxPeZ6jD25TUwIGt1l/m
TfyfCmKJ0DoOrIsP8u4/Bid3935ZK+XGC9OXNA0x/hU/aCJ5636vPth9aLUE63Pp
eRAqQK/oPf9oMLUU8FcwVio+PA8cYg+RibcOVCLCbN0Qtm0UnSNMUchzkYyTdeJM
0ptIRlAmX974bRw19OLtmGMoCcwvZHykUuwN99v28nPLgP/IvWJCtkoZL7PajF5D
7NLZUvziUwm+DM7WRlBr6gF/KJll1oOW29+lJKocVHyV77A1qSiK8bXlrCjRBoJ4
vkO5hJP6nd5431GBcT8n489pVWvWzT3t4kLD3EjtvOex44d5csef2R5YtfPUN6vE
SWARZGrD3d0xLJDjMt5iLuqao8xRCmxHOgjsddQuCldva0FXIz8YyzHoRPfuPb+7
ai84RH19jz1ZoJmqE1NWW9PuOh05g1YLtVbdDn6L0rhYTvVthCL5s6XVB+mqLIKU
0QRqGYTAv2ViSu7nLxze7+734kaxluOtjXPP2Z6iEDH7KBQCTqtxxbiCzUy6YuTS
pTlpobzN6pA1Bl4ndLcHe1YTg01P1DDObGJaU1FA90va16rzVYSqkqtoCtOiWT6G
rEvcZ2VQzxMbEeM2IsJ/J1cm/e1PM45zA75+LLVXKunoDyeuKWk/kCSUgaGmPc4y
euP4snXmjicFjh7d9G4gyXorv8DcqEmHN31gxprjISx2fWmUZRlJQ1uO94aI/Gf1
uQvcQP+pNjVvB4k4x9GQWHMDs3/tSldNuvmVMjSjNV++o+7KskvLWicmwwgaYQK4
eIaqR+AUREaHxRmY8g/lrsQhfabtO866Pesjf8JEJ+SEqg+nR6OyF03I58Op69rB
I6ms1eM/JU/OWixFO5oEo0NyadmOCc9eZuTu5sn3aNKKQMDeSGi8tRRNu3F0HQsA
e2qtcgvQWlLohUo/wL6hbF0r7xbBoI4OtIEn3PyeafxBbCPqDqFTPXOR1VIcubTF
v7tBqJXYweOUsxW2ZD3D+iGrkrzWa7PKpXY7cxidu9JGvXEcYTesrRMjXntacQ5Y
oceFekbgTBlvIOqrFJlez9OGvDGKOcay3jmu7MNEmbXg3M2Z7jSaYfaLXiLbHEsp
bj/4co9Dage37AMka0qxyD5ocpVDpRSkKYXXlM+t8nu/Fmxi0TFPLpJpKNmkjUFi
NybPDnds1yWK5bPzGk0cWiNpAa3nQgtAhkKrWk0B6IUw6pEs9BFlFs5AC+a2mvi5
nqU9BZUUpSkUd42lHuvWGYvhsBTyjFb6NRwlqWKR0PVC9lItn7/zIbIIy7IKmsEO
8UHkKokj9+/PQFe0VFpndyLDA8eZnV8Xd9d+L0XvQRZuFfde08unf1bpv4mh/TCR
h+DnYvLr4dnYw6EsmsIUjeL6RZMetYqP/4Wdgdmm1k1nTmHjfeVoXlPLcnYLdst7
D8xbY2BhyX63yIP3wkOdG9wiSxYwCs5EbocZZK6JhlmgmdfwOHuhGE8EmzktR/DO
5B5kLHjW2GAUoxbpQYBd3oNYKDIcsPVS0CBMqeWJ65AJV8rMZY+aS5VMS2bkIDBX
oLHJH6FMVihkoPQSvwzpF15sqI1jPEjPtDgwDt9F1Hz67pj10O4cYXpKyoYJ+G2B
U88M9gqwe8FDUajh2sKs/6O4S/siQ8IERoXT+THZ5cyFFJPzpBUJg+bUtEmYU+DK
dNUrf7RhcgztQXq+t27txklD4FBcM56BkC6Dj7ZyuSyypHTIZhaYQHUxjHCine2X
oxCEbzoqYvaPYdy7pymS72cE+xb0aE6sOz2a4nCTLXRHoJrjYJ8UiGJEvw+56qI8
j+MoEeuRiUVqVMug5Pb9k/xG0lQ6YgAzNcrJiu4GTTPHnPXc802IFV4cDLqzsC1G
OfuxNRrIQvq+NJ62PoJf00Tr+8WKcVNvS65BDGLuNduEc32KoGk9AzmHZGh8opqr
ohteOTCY/mjVoHaC84SWIhViekCgjhwadB0gGQ+Ef/ums7/F8DDZIJodEROuLRB5
EbVv631Tw7tINVk5byi6XCFO4rnT54x0fmJ2SB4nL0OTtTb1/FmE3NhDtO/cU3xJ
KEjSNqWgbvvHFbkf0VTZJclkQQXXHvgL8aPXE++YwXKcHGMN5eCFq0p28FrZJIhu
ep6Lmar+ngmtkHl/48xYkB33MP2z/uFVqZLmCY6Pd7mQjV2qfhVoGoM7QYuYyRFs
i1FL9FtpqQqs3L2LpJPpYy51yt2BttutlBZRHBgaqzeQw3kM9mYEjcLFaWEP0vRz
RTX8Uc9jVxrymF+O0+FtfMCbuxHyFmbrEZDSGWapVKT503j3H+vI3Rz55v+oBDLt
BX611/5C3L69V8VU+HS5xO3OpAZGmB3a1BDTRXhi/dI/IO72W8ilrKLuhFkjT2+7
01tAnXhIVGwrVMly0pk2D4fI53j4fKdN5BjnvgHBuZixfBFD8JZTuyX1CvxHAMrU
eGJvHFQburKwrzrCrBhOLA5zTBjSHo1LXPcQOBHkfcV8Ur+zgbeOb9KnP347d4ds
fBIUfH8A+skySQVulch5caXG85AeaMj1NZNV6AYbtLHS2OHmXvIk6H2b24LLSmE4
xYy2gs+NW3LZfBRMvVJ8iMYyfvJ4Xlj13BO0/cM3MD4O0w3HqMoUroo22aBy089r
Kj8i0R2jOsE2RV35ZcDyemtiVCJ3v+GGy3qJXcl5ZIOzxUMw00CedWH8QKjd6aUe
1rbcPR4TAv0GEAwrgcjnlrsKkME4Pxw1HWozXuil9vzxe20r2shZZmZypyxlSsqy
SEx1PpZv31fwo/4IDwS/hNjHoRx1DvaysmFNZLFavyUczxK8eZCbI5fV9AFDuJu8
0PooB5znKLBYAQEsliqveWGaTkpeARz4fY/I9kTBIcI7tK7r2BYlTjC//OJcHkdq
iEH/41jwbncLrmzrKhSG+xGXHxAtGcQpu4NGJnnUUj/WA3TND+Tpg78NQV6FsXp8
2WebTJjRMyVzzVFg2ZWB6Vaq+jZ48it0WQWpzWB8a27NiCFXHAlVYZtpz+7gCThB
envCeem8cXVf8KfrojR4m8bWbEObko0ctr77IM903cnxQBHQKemNeWy/FK51Jmc5
v8j4npfun4QcqGLcFiYUO8g5UdP0gQEpzM2repH5gd4Cpd+zckbwVMN5HXIHPoaG
NrRugdHRV3turvXsCo1BtPdNrSXdUnBaM/rLsVRe0gUtUllsT+RVcWHlsL/kHgbE
EkAX1i57kKhiXCgocY9symbKqzABg2260HTqEc5dXzTmZ4BNm3wxIC7O3MF2lwNY
IbE7NhgvXIigt8VSVNd8nbyuas332tfNGlxFu/w0occ9d8KOBE6nWb/2W8QyWXkB
7LCi09yEs0mgFxGrHXNbm/epOMf7rR15k0VylHUQuoW6RQOTEFCIQQubBMRHUDNx
LeWIpOAnUd5CgdPJ9lujWtwg2KCM7kcI+5Si2sUTCvPn7ja9B3W53USyQslaK5pB
OS0bfMrF8NU/mDJha4S7LBLxYBVJ1HLlnDCipkV3ADPLor+PGIuVYqRDIXmJNkyw
n2CwCWzMuQtCfEL+9bGDGxkQIU0JILiPYufrEgpduGOXdveIZHFriiqVrRj1a0bD
P9HLM3dDX4HWpCQuJeqDlv5J5TXGBTnpUV17DlA+QGiHf3GuaVm+DHgjiVCpJkj2
d6dQ14DaGVV5JhP0VzOgG00k7VognVEz8Ns3TOEriLHitn4P5WPCp0C9DXDZZjlk
4D3pBg+M7a8FEnDQv/mWcI8mG+qSytEUSAzPo+/ZmnjUajnEwSA2qLmorQ/9XOqa
XOR6utYW544dw1T2rgYLPqOmZ1JSL6evPsXKxI8hp6yAOQjxrrYIh6ijc3ImwT0X
S/6KgWm+H9P7zh06BGyJ5OUT1RD3304/Zjc83kB3DU1UyOIopk3Rx3fPQpFe2a97
wXD26NpzGIIeCW21jlT3r4Y38p6cMvMhhdajTnjqpyT2ZwZVKEkWvB8XgZqbERNH
1ZVKhqU/5p00gwxjhNp1MAnBg+ebR2cMHI3SVhP/tQcqEAfAO6VKV6+/ZnAv/1Ib
sq49rufvL3bWDzGblalqw/csOtw4Sji6xEnp1LJA037c4frMkOff7UYH6etotAY/
yCoo0rhQTltOQNN4behuGKVuv7IKqLpeb7v5bgKbmC75+33NkFue/h5/tmQnAPrh
BJ9IeP5XOVMedfqs1DkfbkKBFE8oxrzAxJ0Y8CPg3zH8nunm5RF+cAc8a6yPxOCf
95X8PiQ9+B1dXX+WKyikMYHbwsdND7TtVNOKYgk2SpTj1FjFx5IkDI7rcDe/Aouf
EXIaMDMN9zahV9h+ET8InPMUU9hauN70o1RLKJWT4c6LzQIz1blmtoGJlRlsPl6A
LKY8GuEWmy0FJc1lvqGI4duwIr6lKuw/aTMyzEOjX6uWN6HEOAcZq6NdDbSAlor/
HM6D+H1zhHHxIdJwU9zzigE4WNWIZ0OG3vs/yMD/G6qH90Du9jrK3gZsbgCXoWLM
FJKpKUYb/epYChFav6Owfik/g7WSwS/GczwtUByaO3gw1IEQ1oVzAahKIps6M7Aq
AiPg5J6jH3/n7Q86kpXAAFScOutP5v4W6ua7jjgUYxlLcDxFHAllDIN31GUhfWxq
8vvwyTliG56ODdsb1XCo6Oy+7ttZYMUrGmbJSD+7Q9kcNgf8Jf42JnEJYf8Jk3HR
YanljB/hKvPCv1zpHrasEI8BvAzf/6NjCrhqpmJ38SOeVtQYTC0stN4iFIOSWWAe
htLinvcD1hS5yGRWYWPD8FU1pRtdG6qVHQQQvcqtj70od2EoF8gulXHSwmOO8PJX
STCweLO2KaAVPz5pYMFkTE4ujwf75voMgtDph0LsbyMEAG7LrMksajttQd9T0Qqy
LJNfeo4QJzva/ZWiZPYz7fUwjdLUMJ3w93vm9NxlVJAhMyjy1byb00vj08uWpt0Z
wg/NS/UEL25+1q2c7M3cMWnoNWJy4vGK65PHRtkKvX1DYLVgQ1fT/uOC7U099fsr
F4QkRqA+LSQeJYWcq5jWUNbpTgxVGHq9V51Bdb5ufAPZXbhT3h9RPMS/E5ILbo4/
YQSzW+H7gGRyxXcMqjvfYt+p45+nl+mnTcBqT9bTMVVT3UTHQzOtno4wcu0Bgcfv
Fk1OCIP5s2eYcxrp1s7vIrMdLJAXf1Lfigjxvkykr16YgEbiqQLrlqJhg8Lzgrpp
87QdaWVrhJyi0d7dOTY5tecTTyykbDoo7Y4Zi1dE4e+lxGedaQgB9tI/5ZiLpU5o
2mxHFOrfW8iCveLqeAKFKiJMD9fDxNJPrHeKkd4HZYDst7y06UaKdGnAZfmSHNIy
k3sV2eSrYJut7DMH5m/bUf4Xk4R4NVpG7bIuqAhO3BBQPRTR6F2o1ufgYgAt8fT3
QZ2IrDjt4qoRbjmUAzj1XjnJ/2/km509U6fnK8zwYRLL+JIO9mLrL1mY8b79Oy5S
oWDcfp+WYQdjhUSLBPAj/zjQvD19SsCPFiVed2TkWSHvHHSi4P9WawfzjWO37EZR
ojYlxGKkcB5fKT1Dp8RLAciRyS8MlVeFVfcJXJwqxwoIFXoTW9IkqaeMjw0uNazv
A2KWi+nDvpkc4Xn3vVAF0KnEuh91WFuboqvEUjSo7FDltECl2Kub9veOVydN+wBU
aLxb//cVIYBJ3YXWBhuTr5vvOyipHQvdeftWYyX5xH+pZXIc7vFTAO+dtVGd4QZ7
TxIIVAMQ0lqz1F5T22DPbEwqGrprejLVZ2IrblTTbxLDDh3pDsAqar11vsK/Ld/1
g1lLpgy6ogdtF/NZE7i6+7hMj3iD0P0RlU82o2skxkh/jAz+cZnZnE5RhrgJnZaE
mKyUA54ArE3GJizZYEp60V41XXbIEBaFVJqL4FNXLXr9sWYawAQYPhyh6U0zUC/K
1AkRN2fgFP0W3RbyzQLmf1GHaTBkCS6budT4a6MittlBrex2UtgIjHvxM+NwbxWv
CKc4kuHEbDEYwCYVEQWOZucdxAjRtZkkGlXwvgHGvv/MN6q/AP/4q0QeKqeg5ar3
uKbwhXU15Nm4Pp/lDt356pHDCw8bGMjVHxpSQoCUDspJqqRhOLyyMbpeP4zTyQX2
8s5tMCqKbsUnq7ZdrRv7zJljF7/SGKfe964EVDulVPbZYfTr2PM8UHjp1VG+cJkJ
hSGQRC+yELqO7iqBm0LTn30tfx1getu0OUc9JUke+gJ0MgSnXw5hNotNvbNUhRPW
nRSj2c8Toc2E0vnYpqSlc5Z5FAVrj8oe0JQ9Fp3qQ3HvBtCAbMViRMxcDQSaaZkb
4o7E1g4hL9ITcXug6PWZiS/jEwsmI2iaIsJsFg3JwkcUg/6kFY5G7haIS2XL2v4i
jCoJAuPx/RDE9J2ZeoiWDX2BjTqGh9cz9KDpVhfpaDuqGplf9AIgCCrB1ZshSvSG
KzAd5mEyF3BvsaukCgekI+GktSuMA2dN/JWPsJ29/CYSCmNEeoJ+IuGhXRbqoIkF
eJL/UvwjjJczcXNq+4qqHwKsi1Pu8fJermp0yuf0xCkK0gLDamdow/S0da2awb7B
avgExNWvJC/fXVVDvmEHKx+LkH/AcllL4iRIkhNhqBayl1rEh1iZmpa73zhIarbs
i9UWPEwYMMiHWqfBigMz5ytwe3PXCe/3tc4GOu8LsEOHK3I+nKrCB6rnNKHpi+LA
e5TSK+YVyjLxvmG5uAss6E3mdutNpErmxKc1JBYtA7W+5PPRfBxJdAHNMEt9/5yN
yWOkRf1yFFLImsxW1IyxJnQ36M/R56Ht884FoCnJF96p0NbD11Kf2x+qdKecDfZS
qryMAEYQy3k0CD6ILpql7nQKptvr/Yby3X+OkdgD4ecys7d19QohHy3MmF5R51xG
wquST1NvjGdtzEcdsgtsImSUCSo+KuC8hIlJXantSQyWxZGV2Fqfx67B2o4yK6ZA
E+pv5Bo+gljVlgeyI88f0/gMdXOFm7wEcfanwDSdP349zq7NzaDYw2zctWSk7k/6
TaP7HBrcgsBhZTBxlgjMYXPrx9M6/G2zGczUF9Q+aGxtDa2SIoubELZT2UeXm6r0
kdkbT2YHRXXgNy6i398iCr5nZbHRBYqDoTP7tyvuMiyoasQlxHaTy94OyXrWbYaw
Y9rwhqnpqFbsKf8ej2iBokk2yZpVF154gdEukLbIkNB+Y/nqyBx7tPiBx0Huxtqu
nUIWdAmmQrB47y+53qssxsnZ/MeP0w3fHQpYJ/ABW3Zv4ZWo6VQNXyPKOhX26eA8
eCV/05rtNh8nwj2efmgU/EEAKjMeDkMyuOXDzWK/EDuu8ilBIzr8T22zUvJZgX9z
OL8r2p7HcBOcFYSf3PXls7ik/V/MxtC48obb37sf+jDVmfeHa/2oZFHqYe1pMtWL
0mGvmHO8NPzts1lDnqMQavXWBZH0YNkF0sPgswaxaPEapBkNuqMkab7yLiQViPUY
PjJiyKV2RKk/yS+9ROL/3mUHMdLIJzrT0cCyT11tLgQ/DY87wMiQuiEMNwl7XUEm
tKyPhBCaZWKkycWRup1hl7hq+ySBViXOS5S9ZNQRt4kz70i7ytnyzTLQqzI90nEZ
ZZNbGcLsHkF8qjH/EEkhv915DZTgZzx4ZRRr1iwGEkp9C0pasyVzdFGTXmfEbilf
wiMNLIzLJv62ILKKSafJDZNFK4ymYySkrIIN97qotU4/S4cu/YnIWotlsh+AwD5B
hiiSElJQ1yFGq78ig0ZgLGHU5jbXJQwPm+iksRRGHuzZ9d00CMRh+wFjZq/j1EuM
5VjRvnyIssLSjmH04qiRPZcq7CbXVkBYEmezSxebYJ1yXhry7hLqad8IPx6exsfO
vNRl/u1ZRF78/5clZAqYZ9QB51ZwDvT0fXt0jO0XPNdWOZcx0cx1gnuDWci+b4j7
NPDth6wnLskE1WmxO8sj5xIieyWJbquJpMqa5XtXqwfmqGPQWpfXfayDPb95x5kF
4Yl/L0cn0LK2iNGoQvqXx/cOF+GSueh0S6mHtLJxEjf9t80ig5uNrtb3sYiBsNpn
ENPWpIqrFAvtCIRdhaeLi9L6ltU4FlHlh9M18m0Cbh2XSa1fXcRWPh0bkeI0FTEh
GyU3I7v3nAyDFyAIDfoY9Ccm3fzegjYMZ7oSUw3Ree2UfC/VEDKiECN5GdTp5nEa
vrxiYn4atdStK9tFdWyApteR5TC/CtyQ/zI8eD1HJyM7cM5OKn+9NmFi9lRsyJns
8WKpmokEvnUFy+qFoJnoomwHHZLAu19zpLFPF6SIp/n+XP7zHNALugKLs57ZoQ5N
vC6UeIhhhy875n+nzEBi4IciL8xgxIO30pknE4RqcVCukjlavNoTcrvw3SUw/RGm
CD3qtcOi6UtZobk9EAX5Zs+jKDhV2sC3guO8wBhNbYjQu7NITClhrsnkfgjOjVwx
+txSKhkxGgZqAAIn6H/hvNiCCWtQ3K+27x6nt92rrHrT5cmDiw+e1WcjWBCzfUxh
yqC55+DEnpykcvTseKk0DRiHDxnnYQz554Y5qpb/qv4EqKVfxXyVHV53zSE/LlXi
H50R6jSZ4MYD1+BleQqBNh3hD4aD6km7Ufn8l25bhBlNdRZaLcPBZvoLp6n85kH1
zB/hBd1q2XJxwLAgRCur2WBMnrdXYvpqJK3X0GTDTxJgVIrlrn8CmGckwFx0f+T8
SEXFEpOlIKvF1UxCvwGgYC0SOUoma9VODY6wuxOggIAKMjScXNykal6jtvkoRKiF
mjPUSqPvq+O9+CpKoqaEGwcJkj6kgzIbEwcEWvGSwDjlAHaHt1H7176/jIaEyTLq
TKLp5w/usVpIbtFuPhGtN3Oi7xl+0w5WSegwLW3wJNmhpMCPW3dphgcZImrQNGnC
JC9FhP8PQtB5ehoVyw4GhSq8xUqqMayEY2bb/y9kOzszRbqH0L63i/Q8HgV/Ibap
7D5aQ5hntaz8fhORhOYAZburOlZZg3qmZIomlO5hXHX/tTiECUnd2LwpFkEJGAoy
2KebQWe8wb4kItntameNW87HVeskNxS7MINafeJcEGJJhup+oJagNRG2olqa8GAr
iWrNY5nZQZrzuBBaLhe6P7V5/DPElnN7Jz4K7gjPHDkNhqvGI2oUNZm3HV8+2dpu
dqolyJjfzegTKdl7yVOLYgK8y4oXee55Nlpru+7z+JnIiRopOpKo8ZqyFj42AWu/
2mKehIVbqJABJEUncD/wUGmYYi41DZpjZXlsbCWbB5ukuWyCcFfJTOjdlauLOvVo
hWkI9J0jsu6z03d/nyCV6/aZjaO1FKlvgPcurLf6zX+kqNLqEYIheZamjIz8Byfe
edKSdUlUP7+ACi3VPffj5QTSTi/1bxo3bg5eIiojmorc/kRgZiIU5uvQ6Pt0JE/9
gyIRwRGHkm04DmEZtUIF6u61i32ueETCHVEPCJsCXyF7qBs2m9XOI4EMEVSfCc76
f9QGZPppfJyGilz8mwAdQiZaqNbF7z3aVZjd5sE3B+Jv84brbhfCNsF1NP+ghBzp
7OErUfjMR7s8IWM91jrXTxllF0xpIq+Tgaf6jDVaB3J9ZZeA50Q1VWUUV92J6HCU
xB1TW5tQ8NBYpEJcnd1k0i5F1+Qgv+SoislP80vfmBVaP9Z61m4gsbtq27PrrDn0
3kNKduj/XQGo19DU1TLCrVrlZAWQNVGmOoKjfiPbuZ+v9FUDO18s3s+4Em5UvzRa
m7ihSfgbvrk6TPjntErUPYDUKXvrYUh8UNV4ndrzewGuuGfXJ6K11dAshLQJ2odj
O3xi17nd4bUVStF9+0/JaYXGvSGPfDWOBszwJLabbRrHq3HurNovO6TojSI4xixF
dv3N5sxScuVFeufWzUtYrF7CgrAwQE4QbTorB6KP0FLY30Oy0HVWvI64kwCKODrS
sDY6b2xZGmkneJUi3M3qOcmnrzffumWdul82Yn3h+RTknvVoNz7uexgaVe7RK3Co
HQsbP2IJg0i/UDfb73M+nhOhlQBr7Sp4bgUnC97cMUMCdTqdomYjz2B5FrB2Y5BL
TixKz9gLrHeNkGmCnUoe/dpgaQZ4Tycff1yQnhmiR86dLZUASOmtZUWs1Z7juN/Y
ALRwQRB72cjfeUXDTo4Coaki2QXyS3AKQmaft604Qp0Li6lohlT3lHBtc4OJXFjP
mR/BCWD3WL6r9wKWTUnUVDrRJc30WoIg2CZB34Fv3F6H6n26Dd/CoKmPcpGVQVRS
/2gM9a1NMW536zfC0jfxMdSRboTLLXe24e80kv/CySQs6NaqHmGEOLkdVN5rC1Sn
ZmPvp19jiLz5mrPjDi/pSejvfLn06Vzn7OHyRHUHuUMb/sGMKpKuIWzI64FlWxLP
IKtJgILe1/5OsdAFtDWbjJZ0Ml1F/MYWRBn1CqrNVze3oDq/zxcamzP1zIuuLu9d
z4zIYUf7AFQ75Ul8O9IBbdvHucwLxhdcPIhOWU1qYV45+KejTOC3cF8OrdQyar5Q
QogOEHzXzPM9m3DREHWEkAGpEL71yL328ogy3EC5Szl910r1xhOzs0jbEWOMNoiZ
GnQaHTe7/yJB8cA8meq90Qc1e0WTkPJIkYHN20MrXimL2NZurpAJDJmFETzJnrMb
9vGJae9cNMponW0gJ/MySvsiZyoMBirPQdJj+OP0Yhes3XHs5MSv8IA0DNKgsNyP
vFdWGVE2o0dz6UAluPr7LV8JMaCN7FNAHY3uk/WypEuPpa4wrISSUZjL8X1cmk9p
uRdDv78FaknTFFO7kc++j3N2acFhbpAKxnhGYMrmVy0GmmkqEr3paYdvxFksV8aW
Yjoe6plxnwfCO0lwsr3cRQoF5k+zcfN24LR+J1nwmsJ2er6pzB2UBsUQb17ym552
8a+rBfsESCH7GdXkwXy4fuKO95yYpvQ6MVWB3v7n8uGGx2zsHKBJ1V9vAO4lrU0d
5P6dvTt90ElNzIKJc411m1miJolM9vE50aWhlJ99Hzh7g84J9359UFZXY+1yJphk
kNFhPC1taP5IhO0Zl/vhqiZNOhhCI92QQN+OUzb0XQ5WahZ8s6jl4Ahd4DEPdebQ
alcDLhj7qRIc+t3hM/Kx712mDvKmiGDnSBJmBglOk7SW7ywQPZ04QZVJHY/wpZv5
eJ+uCTrR4JozDA5zLNmXSH4apYnh6eWtPEuWIJWKhLmgcPhguRwnpCdsCyfrVToa
e/KOHb4iJqvqyki2n6RYnouXFkvGMtmI7YDQ+BKDVp9iA2/PFC0lSlBiDHv6DVIY
lILtliC7f0/dn1MR45LRQz5bCJP4VGmaPZhM9Uoc2jKrsfQfvfv6qrAt+VkcOWpC
2hj1XPvcZFwyMlTwhrvbzvomS0IbJKfSxhMqEXdVfj8cybNbmI0BiDGdhzu2Ccho
VF6sCHP5ZTEbqwDu72aUyahVnrVUQvbrq/MHd1WpPtvOBIyDQgdyO+jMFqgWViVq
d2uvfQsFZNzvxoNIl8icJ29gp1o0siCzxNbLZE8k5kTVzd6xBWTqH+Ylg/PXPCP/
vfmt7NB/YGdzWQyMkZxWsem4bbU0TOgq3HImll2LFR6OfUSJPGFmSbnQYO61nYub
3OrEsfvbsiU173OAbaE7nijI61yvbkx1law/Kh6Qsy9iIW5NoiPWK8thZ/aFxeIk
KEKegYFvrC4XDzlf6BZ3pnhJn8+4VpQdvnFqwH/M5DOTDy7KC2ZP1QVXPZ821VzM
7txtf8VZtVv8F5uJmWJQZZmr+tBMcOrWWC+IpdYXRJdTReEUMjMPpRnxthAVDE8Q
itLyqnLwlsOaIesapSqYsZPq1OGqxFrRPbDgiNOQGcKtm83T82ENT1bfTao8g3gL
kjCcUVRy82+B3Q3bc7V1YFj47hYOcaGGgF5s7h4TJ4oaw9CXUFMRcnamYL4REvGH
MsTdbItPcuSwSllYDDuI4OyARhOzYqZhZx4tMmE3hGPyZ6DO6u54mMgyZuziNquG
/DSsn4/y5najVyCcdq/bZfsbHkbrD5QEGnbK7dihT+vryHTQY586DcEZ+GAqLFaU
SE8Bti2ZCzxfGjmbBYtsvPkuZWSWfB/HMzghkzVO18fLOtaggULudbix54faAvYH
AKYB3aD2Fqf5i+4moa42072Fi6FavWczS/E+KuNhbMqStnypfVzhCqeM+vIt+58L
OLuHSrV5tfgO7+O1woSNQm4gvHQV4gC6RRFMxa2/1C+34J6VK2DnEHaA4RqjkBnI
X3w+rxun7iZcskW6ZhTtMRST9FntBIRJCyaPOb4qUGMG4BBBv/riVNBUkYVNPioH
Vgn+Bu7Wje/AqF8rOy8t3uvWUN2BMoMQIc/RK9uU+87JjNSBZ9+pIKHlF0mXSRM1
RGe8ztJrX39z7iY+CwtO8y8BD+YTsvDibMxoBLHmdbtJHnk+RzCw+7mgaXFxgTYA
3zRYZUkZTQwIRAfvkCRNPIuvPHS6mYT2lnyJCrLmMa419URciR4tOcDX9jRHWbDy
6nrnKmevmOpuhvY47dsIGEJQiE3dPh8n5LnPvr6nT6qOiTLpeAgwAK9UbjVaFhIf
v0a+Rm4oTIKUjYSHnF993tGX+6tRnXLJ1OvTI68kOuNimkQH7mmBendYW54F6Eu4
U5tRVvXKbPgk9yGPMk1qkDaFiyATu4lZWL7eehM5+43z9aYB1gqgo333yBc/aejm
RLi56c/GMU5Zwuq8wv2VObUCEokZLWtJb2ASjxPeIGEJuvmYTSpCZMkb4qYmB62Z
tE/yM5uge6cXYfAkdjy5d6ubPHhnjRXJMh9h7rZn1qxKaDUqX9gJNSNi9z2plCt6
ZHuOSTzAvTl4lfo/QVSNP3isbeOEmTMcwOhNfeFhxIVsk8nHiZdMOGn131E9b10Z
1ov1yQVXFVDf0bwlHsnrmcgFtoRpZIe1IOg/lRZeL8D9GJNbC5qpNwL/GHU7+ahV
GT0QBdDYvlqjWcj+ZOTE2CrrhzrCZKYz0HjrmLhf/OBamNNnB6IMCSoICqq04D7e
42WM/7RmkppgWp48v+7emeHfQx6Y6J+vkCKLeHLPlGK5qe3o1HQlqxQBFS5xi7aU
ChE4uUOYbsSV+IocOJ37O0rvqODHAo4Gb2fjC/Nc+w94k2KLrqQcIVrHoosUrpZO
mh19PEW5VNjDv7Gb60WxzNeBy/6zkS/PpWFeDc081lDfTmv65Cc0NGzO31f/XC1M
Bar8AUhE03vNe+w7T8tR3rgCQEvRDxo8cxslWruHeyZiewH4pMJd1BanxaTyJEvT
lDkFksLnj6XgOF8CJm/mr5dQj4EBFR00UZVP7tOn7qiii3T2ZwOZajv+h1MRjncM
+GBlRWoNqi4BIFE5kXDrjohCw8SW8NrFqUaAcIgLodM6RCZ7lr5Y/iq4LyEba61z
Nk1DV6DBquRJN66Dopb0VfCyOMp/odjXP6+z5QY6EhCL5wwX6rayjUBuhK9Et+Co
0LXxxpCd+JIEtLr6yZpKqHcPon8vnsiKbk6vnyvXKZC6+YvHisHW6H59TEySK297
Tq6Erf/LbkIOpweNdlc+hRyKyylbx1k0zJsgd3BurwANnNL07nOqgiMiKkvQv0G0
PPHGX6GRVOPQjl1o+ZZoM+/FZKGhE7RCmx1PKWhrhItEorPsxMRg/WaqpSErurp+
RNkdq97w7RIRdkgQA9YE4HMrV//YYm/NmAYhxD7A8X2D9mKEEXCZTJBpOSVqRdfN
+AiG78w82O1+dmkq+V9zuiXU13fVpI4BRZPMQTUdZI/I5K8slsUpJrA6A2Tz7Zkg
4Yecj1xoYV+zxNo9GoVeFCHvU0QRxP1mL6fsxsVyFkDjWSMHA8N6sLi3YfNPg/El
G+NVReIjRT1NferFpCmSpm1CKuoH4KAd9YpYxTcbDXaapb6q4WWcazrVfWjBsys0
ZTuDrrVnGwkNq2ap4OmpBuqhBiL8uHUZJPO6dPCrd51tn0TLLq65l0f9E05DVcUu
Krc/nUzQfGEhezcZkHDEng8a2ua5jwEb1/6zblz+zlIKX2mD5fCBYewNTvVOReyS
l5tYH+VtsVMqr9J3RCN9s9UcCn3Va32kbsmL0ZNojF88Bi3QsJmcxq9ggpqSBk4O
p6naUq3aWkvsfJBBrq1SUe4G0xD8BDPAYhF0IxJ/oNp9pBW6OLhhxNaWPiutKNaz
tLJIf4OqXmGZO8CIGYlHlUp9y2DYEPVf9JLn2tyMU25vqBNqT2FJxAuyZuP2ZQgN
T0mFGDSqz6aLDma+CDTYtuHQd4wZoQP2yoUSsXYwligMv53+2EWD4LiOnqk9FVip
8PN9SauxlkL+ZopWTkfdNAeovzqFGu+pbKe4xiTd6qsz3yTP5OQPq5hYduDl3zO4
Awe/z8lOMY6McA0PcmdrlbxysknubiMOlYO63fsqhplpcdqBCW0ysT1f9NbIqldC
YxTN+wzH9UvXOZkwD4cQFhN2hCDi9ylI5/SA/7FDm2HMCdOawPN0G2Hh2Fh88h16
gkw1b4Se/OTTOJ2eiIov1r5fzretOaitEfdAlL0fksa/Q61tT5h0TBmr8shLbALn
A/JvmOfs27QMzAiklW6SM48RlK73exzkVANHL6gzm2oldLVAJ1KmR1b3sAK6v3zq
ewFC8ycv3RPXqJZ49Rd5AjP6cA7xmk4iZSkA39oy+b9DmPfam5AxnSD+skbfFlQ+
39cYoIAACV1SE+ExdsWhxfOCaKjHycYOhypHQuQzuYkb+RRFDyYV/tsi2kiRlJxv
2v2jjQ7GlcHYum6C9uvWI5WZGPkKvXcCfj46pKxSWQxO1F+t9EpVTwIms8SELfek
tWi4kTVctZa1qOSeXaSlYsdTvbPdMq7KErFkjzFxrwuZivNGHkYL8aXqqZOvJiQy
uj0AXNnfsTzDKYejLqIXVVpbCjHOpW+5n6hycnHZgCz5OnO+3FWchFJFVPZNmnKJ
eGFxx7bwlCyEbm4jcVovR5RTB5nfmtxoyGxycD1xU3ojLPMkanR2J/1tx8oehcpD
H1YYThng2ZLVFOtVFLJN6ZtQFJEDNZZN+f7dtnctSQzhrTd+88SR9T4ZAyT11mzg
5PUi2ZKG92kvdKJ4Ks1I1B9fR9qX55e2OqLBK2y2hU8x0qux4mq0qJ8OxMXgOEGg
OMOrdwoiP8hXg02t3eaLKjUT8ORB+3c4fI/2gEgLrwdBGaqsoNdlKjaqEYFaQVbQ
UGUZ1srFFI5lfbIbr0U14bwKh0axFUYzn8WgUtaccBFsVQLpvk/jH2+jkkOOa+Dm
U2Q7lY5QCS2jjciQ14Fag0Ymi69IQKSc3YxjE8xctltJeC34Z5055BXw+36ImfPj
CDx08ZEayF0eSlBHeiw3/HEn13smbZ2+lS4lnSlu7LrhKc01UIkrUE4JHWCKlC98
UZSXhEwlT+Yqguem5QNBfyu/UT5XYgHqTxS/U+7tipraHzg6dvor1/ZJ6KspUNt2
c39FQjYAbkTTUgWCrfXDdQdnQ42ullAZqspjHQF7lP3S01g9Hph8OWCaqnSv1lDd
XNYK5Oj3SL3bTBI9Ew0Zoam5WE4fI5j1hJwiXqPJp/932siU/XeO7mecLkucAiLs
LVQgM20U25hZEL7XUwJKZIXtegTiSylURl590QAGwCe0djwlYynZ9PQ2g8/vl7Lk
AXIm0c9IJ2TkYXTEYLNdS0qrzhIHG79NaVd5xdWZ+kaZ5jHbbUqcWUMshrLDgRTw
1hGRCW+k8bau+1c8+YKED9bVwbf2GASI9AcA3iDcer3TByI5MGVh14F8fgYMEYBZ
BUX9kIpOKs7YaNXAON9m+XWP46imyraYzbIJ+PmB/5lJSOzcVem+K+dRMIUd8Fx0
gT9KSDhPcJdhezHCtc5WObhjYsBODBCfLGkl2j3jlNwdt5rin9Ysa1UDeZgGRPk+
MpnhIhXdzdA/Q0QQ1l4use0RcbfUUThG6rrsQSymj3vzX1XP2vtCGyY80t/zhWhg
jjhV3rDiyoLn+IyoUm0UHKRuD5JR/bCKUZ8D9CJWN8Nh5bpYjIp0Fwuxpkrh4TxE
PSONmA4ouJVqCubM5tcNu7lUmZGcZ0aAt6152RxOn6vKlDmNEU+HG2OsaFw0qQT9
0jii4QgdQjehzqWBroe/VokMd1ZLFykFm9D7QTSxRL6M9gs2Krm3w6E+NDmr/kfi
KicAzsCBPyDKFdRThkHIDqcS99v1TpaeESf8Y1S3hXQiXYmMo7Oi/xFmyqEwCKoB
abAJuyznAbA9GhTXpe7ws9YObT9lwSWgiLHNgINfAoclrMN3L0rjyhFZ0+U5C2nO
Za13YjapIRwuCealSzNbZysKpm6kxqCyG5Eyv2YBDwvfpxCeTgGyuYS2lnK5QNBu
nC66DrOo/ynHv/f62s9i5w5vD3qTqRSItwafqzWOAKD83La7suM3TKW2UyDnkRhy
qIO15GiheTPLc/3V32xEwLc6aVpoJSIbOIOb1H0dBglAqMFfNtPZL5P5Tuha8iSk
jzrv3C/A5IjV5wjQiSaEaJui3T4I0TqaVE2vJmcN5P98LAyrqutB+MBcNBp6a7uG
IFn21km8T1PqTufD7sF0LZxigK/EjYLFPp6HhZNuB54EvoU5aRcfTHq+5RFnwV0d
bcKQsqGNnPBY0AD32W//+KBH/ktkmcRWj4PyaIYj5S8iy5YM4CY1BdvUOMJJhPnO
UuR0BmBiFSZi60gzT7bYzNNTmvtINeNnwwVW3m5t48gFr0w9L4XBQoJNhctPM5kQ
JYwGfeoMSXesGtpMwzLf7emcqduCZ6dhY1Y/uonv2cm1gvjEj0duwv26A1xA/jdd
ivrlxWYSpENPtbUWffyFG5HJw4xpG8oVFkCw5GHWKlKR8AAQCJmoy7ztewqrxAmC
5Umwmc0Pl3D81PedhvR8cLeFHJnmuOt9HLq1JNXdXZkjDdrnoZ4A8MgHMrnpChPM
D52muqUZevkWMiQb+qHCOEws5gc+f7sBphpdPcXzPeHAUuMlNpK/K80SqsvXSC9U
UcvKQlJcLOK1M5isjlTyIikzKSVU4KmAHqNMTtHNg7qgH6DmhipQvg8lLi4LvsYb
Hea2LNn3h5rsjDgR0xXK1I/nAslLNT9C+d6Z5PT82xHqeP+vmExoBdYQUGsiss1E
oJjyDv3/ple2tLjboE0wrPCkJvEcXrfo6mi0Qw2ujo9K/NWN7lsxZJSEMr5cwats
1u46+ef+bXrJmjdWQ8gMJF50VvYHBqDaFU1m/tzMrtlX71+xxfPzpNoL3v8ggSUV
5P2AfqI3zdBo04Ri3pbJx2PmjUo/KjbjVoXw1BwM5LUcNcBCzW3GX0RYcikuDKzY
hoe99hpZbShKQaab+PK77u2WlI/fWe8rcUVKGtA9qL9pMbftRGPk41iFBfaxk8q2
oke74JacdAqNuoNBWZIJD5N/s/3ITAnZ+9+ZblgG9UCMNK9yvrTJBiysNnI2Oh6U
Vb2ETiBd0UESsmujUtaZnAzhF9AQY8473E1K+edVp9QWHKC2s1vspUKTMxickjXt
Le/TMm89PtxoRTJOilhItUccKDVxDdkWkaEON85wPV3JCflnYyDzLYxVsBB4kMXa
0qBeyh1JtE3oljn8FxQIRGd28fP1EYpT7lCTfdkg7qOLpturw9yDAgjoCQV+mfWQ
JKGBMmVOLv85KWCDfDO5Htx2Lrj74CbgUYhrtJ7ToTZq1tBtkpExT17J+ad5yeC5
eXdoAuNM0IWL1zOqciho4X5pM+9kJBxNvwg4ITcXe8huSWi9dLoTcUg7CgtaZzDv
8+vaykqc4B10bQ3GQCFw+qxw9MeqTSWlon4WA0HvrnYvpaRPlKRT8GSasjYra5BS
ihZiA8v5kt03fRAHTUGB0dgvDKB7r3FsB+jUniPXfc5CUhbLITxU21kiwmXOX0Jb
CzmchaHXWhGYwSk3+i8kCQ/IURDA6C3/DPmMaUWlOK+vZxuk0y7v2vrJJ4qXiDfU
wf2dibl5QEAHuvruydJ96I6tgjj2SJvjQWHrH2jVOuqaV07uOO+4uTvG0qTl8Osq
AxdRMeC54aLT7h4eRtwnMKTSUWQbH5WLNSSao2M7AyPtpK8a4i0ER1RwWwvQMUGp
rSIYiCgzrpAKc7sUKt833jDYGwKSBOuuotrU0CokUAKMrLvlxTtW89M5WJAFg1et
pqm5hqNuzE27Um0RMlFtlgsanZCoIVKmCFrUEgSJzPof2kyBjV8tIgpVTW4GaSuQ
EKvIfUDHlrWB5pe3JUvnOBNRDYARvkBlGKDgAttVbAb8QGm+jNlFovw45TQuyQXB
4eCNfjXUGzi1yrxwKo5+Cws6aR0p6XDReh2lLWKXZBKqFrLc2weYJMm0bDkC5mx4
2hiVii2K8eGBWEBCZcBbUHwxRXujCP3DfH0LspKTlvU0CwLB0FZMThSnnhGYQ9mS
qWTPk48MgkvO+ybFwt6JaBWmg+Hw9LFaHP1UoWG4N8epUTDll+Mammu4eAuE3TLG
OEZbUVlpwmekytixzztc9h1J5lsAQspNdyydERYKspgImu1gyCrkc83PrtPMV1UY
GR/YqgUpcR8jnUXI+AxNqOTXcmScb8a8RbUfglLAQHYnXB1JO6zynowOsb9VO5Ya
luUld38ejiWYHK8MM0bJpnbHgHfWkjRKg9uUG4zNav0i51JexObmVc8mQX3Cx+Uq
T1KEAzwdIEF43mH+Z4EtNkJ91sX7J0RDJ34lMoGd4ssOKvRVqhWoKDkImh2pB6Yz
aGvBr9fQLf2+tf8729M051Qt8eX4tYWMEPEMvvN92iNincv40PIE4EGGHUaGtxyD
pdeGzye/c7aqMORWhAnDYjZL3OQXyj5YV61RURsR5WOvhsFd1mPnnZXo4z5F9T85
cvRfo9b1XK2fYxKeCoxJqh1kgjLKDmtGhm8k6VHPaLvOMDwNLKrjhfAVZmyP5OLV
CJAjV4uq76E05K4h5GpBL6kSnqw5ix24lArGOk4oJjh4VdA3KNwLJZFCdiIKjY/3
mc5lvlEbge6h8Ne9o0wfwDFhe6HV4yemRItJrfBT80DsOX47DkkMI+ZwB2aFt/m4
DF88hZJvOy7WErPHkhMTxy8l9IW6wwQlibdcAEwCa8UOMZ2b3lF46A9Mgrv/MsRa
js8DpI+g60B6bLbbbNH6eZUpWwFN0fl+8k9tyG3hBk4d2RI74l9EweCEBBzbNSyV
A2a9LfkuxD9O8kd267z+VJQmusbhSTnO2ghDVh4D0QFVbbs7OoNXc9kiTNPBSRPg
oN0gZ7ONg7QJTrkzuq1LpAB7x1Nt40OubDmK/XQElQOksfOzqF9vbwqlllXEfhet
/qGFIALshTX5BtVPrqo7UH5ihLiL9D5akjbickiJl4HLC6dX8kzwAb6KExutIAl4
DG3RMiXghP+Fo8iXhs+oxeErlHg376orOnUE8H1wWPZQAfqlZB1G1MpcL4Oqski+
/xFmZN0oJSl9Zfoou0VaDFaQzPlY74DbDBX/wwuF20b+eM4yVRflUNK2shUis+6v
cj5wCDlq/CC05Hykja1NMDbi66jYddNxlkRQpXPvOU97Q07bXso7LRKLpeL957xs
A3awMktb7ZZAp6Q/N85+mcpME1uIVKrl+1D5ELoQeoBsi8x9NYqTYNZhUJqXkE00
1XFeFwqEowDAAr7OQESCNHB5jSPIeqdmdyR/4pF6FqXmvrB0LUKJwE0PSmlMfDyx
7WABKG6pIAM591BEpnJHVdzKMd/Kddl84RHQ9TuQ07onREbKdTlS6iwGc2X7/gAk
OF6HpAu5StemDTIbk8i44AqTnce1BpNxbjFaxJMNXq4Ila/zArFUafG7tuFYmd6I
Ta8kT5cb/1BFooklrUbg3/TQXnwLv/d7VE84fVm5XFqp9TaLM4gOzzEvSF25Vol4
/73KAUq9c1CISfNYO1Z8UXYqEADy7chZlPWnNAEw9brJMEBBbFSjkCCe3j5pR3dF
qJXADA2wapU+piq40+BuT7suTc3C3uQb/ztbGSMWRiOHWw2bvqB9kK90cfO5p36Z
Oc9vok+86D8dc9YPVbb60ygCAt/783J/RjGr/c5dzZpBOI2iM/8oqiA+Qe3BpYRu
3nPmxYnYrT3DQPVc8ZRVBIG+FtxQLOGQSNLZx2GjI1ILUPRl0JpxlP6lzAF9Se59
e2VWzG0I7haErxYnVoa8fCLJxKbLFi/Sq8J6n0IuQ14JC42eUSm+Qe9SWl09kSv/
fdBsvksuQC20yKapIk/HnmV+z5Ebq9tccCP4PGK8RbcdpZsyljSaFZbBLC+jsQRb
OFParBFUBaQynFOXV5rN2ARyZ/9ZIxBjklUP4ZrPRScBR+AXgoUZuhvGZZmf4/yA
83SSbSRvlf+r1op5VQMoS4ZxxOjR9yhp9Fh8dKtzAXCQUanl+bTArXeDtqM4ykQ4
pmkfVzTg+XOj4oYjhq2ih7ltYWWXB1fYN+qTNYrBewS/9HsP+aEfI5o51Enq/+CF
wWKlfa3vYD6RHZHnOSWXhAYGpF2tJ7P/8K5+7+/csqLBusawWQMRJDRkCMpxg54X
TPjPVs/ucIIyFWNSG8PZZBs6Hh0bWFWYv0Tn3CzEkidcVASI25PHAhsvc7hZihnC
6F6JUwMpTyCD1m8z4XdTQuwndRFXKw01cJsGA3HqeHQJSTGh2nieUzqQoHxcHwsk
J+h44EYboCtVSl8VXWLZI/jMiYqkPYxd6ukbnsqoSnIY+j3bC6X9HFhifRl47JgS
j7exagSKhxIcdeQCSDV+i/rNMNnbJMTt2fm/Vv4yG5b3++8CsPKSPCFpKoPHvEH3
P77xwOM2gAbrO8x6BOhrddFFIwjXigLetU6KCKpLA045JyYHgnUy1QiQX9FSkSVX
Z2urZKz8t3BIYpxHUIg4Lhlqg01astWXgcm6PG7AcBwjnPx/nD32qJlPDV6WKyQH
kFuOUN6g51uooG221DFfRKm+D/BA/3ch7cRc/E6UMfSDqSopdpy2mXMIPkqnqWwX
zLrO75fLcJromhZzVqfltL7wwRrvUrypNjrWC7UVSfrM7qE6ZxEMBpIOjm7atcqe
cBcasqZi1OvzQeEfIGMzJb5KZ/YQxskIkRr9z+LtE78/F420PxPywf+DebQkyJ2G
dM35a2OK+85jPQ2C+0d1+WHBmtAR0FfUZ350KAw1eVEAC7ghM1+tNnA9vhC5lZSW
ymT4j4+X6sc9zaSFYj1paTGgkjVWRF98zhzI7G3Fws7+YugOVRmRlOi3KAJMalzC
yAAaw2RUUOblsO5H0aLw/Y/rQhCehtvVSeR2q0y3vwu43WeBl2+owi0tpgJbanx0
swYgCHZiAP4B23w223cN+myaJ5fWuJsy6uvVJntFGGsM3QUZIeyHI1lYxY0zfHH0
lfAje6VPhboNfG9mA6IeiV3xEsrvOYxqDtJECDFU47VN8yReIvzZjZKkq9dcZKu+
6ub7lKHCBVaD9q6KNOXo0fqZ2IBsN9u4EgofiokdEeVQI2p/lnOiyx49Jm1o6R6T
zFlsWcEBA06vOIdmyYDzhi1+rIRKWY71/2xe1Vfd0lXezIQiAUZO68EMN9QUnF0n
Hq/ZP8WuLRelVMXHn5R62DY+ETrQ0kcEgImTkdebAk1KnuBGS3AjVfaUKUJKaszn
PDii7ecXmB/D1A6b7bg1AuVEtVVPw7rPhjxg67d5EWPwIN3SeBnNrUB/jJIRjf6w
1edFJczCtWCgKiJAeUA4fWLo2QEVgltMF1p+iTTSrXhz+4qK5Lw1GYpyvbW+Q5oG
ikb3j7uMng17FuSTzoT7jvXjKBDDrvfQgw1fWoLsooRonZHDVrwEd7QBM0y0CoZw
I4yQRrnovf63wuoXN7Qmg9L4n46z1NIUiXx906qFN2tL8oZ1fuAVmWJlzNro5D29
efDw4qfC6g37egJclBDJTU1Xb6XiK729H/vJidV9Pgf4KxbG2K5YCLLShRIvTD9F
ShILPHrX2RRwbLvZaL3nXQ==
`pragma protect end_protected
