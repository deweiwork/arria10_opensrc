// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:03 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IeiZuebyYQYmnpZYaxqnZNFeIaQM4WDjqtrvXB/KkEvcS2cGLShnS6Xdw2My6p7u
u1Gkqg426K9b1RHHofYebNezvu4bB4ibwm9R3AfGMf8J4TEHdFVilGVTGBXXHCl+
W/fg0GDkhg8Xvcfhb4/FC6AuMlxKeLyWaBt69n0CcZo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 749616)
+oRytLrhepFY9Bw5uXRAqAQzK6ZnWHEDWwW9jhZXVi1548I5xoXTVvnfxhUwW/sj
EzVfwan455C9Vzt2WiERtA8PJBnrAw+UmaZJhU2DH4pwR8m0my4EfzqaV6NfcH10
JJEnFnWppBUpH3Dy1837w/9MxghGZwM7NsDbdGMwJi+alt4ey8xonimg6e8RhMfq
reZ/bRb/eNjEAfeoToJ5nvWpbozMB7hmXV9MuzELwlwT55TehaldFikGqWOY37FB
Oh7pEpZKlDGpHPfuXsOv2S3yE1jKIU69uNLZ6DFQMDzfIoJQeXqdsY3BFhVM6JQl
F71TzQxu+9ALPDl9Gla7ghsIKsaql4aO1nmeTyLP7Pof42m3MPmk0j/JQTEk0IVX
N4K1Rp7Hu548EZlsFBtBNqix3zJjhvvx4zTQrvxIZDcn/YwlFRbjN6PLhRrouIp7
T1y/Zhis9WZYvbltjTpWgUIWLFSP7EihH9hfAiPAZ7uVzArOcSo1STlEGv5ZDU1U
zGJbVVScSYK3DpIwYqrepI5U7edp3MKAFLxx9PwhnkZkmzcgAwhFz2TAHlL0dfwE
21OMGsU+Dktu89Q/dUIQxY21ZKGA0RAFWti3tC3JVsZWjIBM6majLm/3nDLNr08Z
CZgLARJg/icion5HC0yhxOL7WDH2lN6M7POvHMR1DBLt4nplaQCh87006ECm8GvB
ypgOK8PY+UpT9P2Zpc4mR+IkJEZzuVDbQYveAFUVwKUFMOyyHCGjxirpbvwF2P2G
6bI0M0lhmuQH7uya7Dzp0gqgPLe+fcPSERqsQgP0ramXCKoL6U6mgD2FX8fN4ZF/
WM8J3l6Dc6C+LaboYa5UukuKtpto+KFJTePkfVMxAC6UyLJUal11rb1wCshM35eN
Zoq/pIAws3RGSS3+ieySDDo6pJjSLeFWw5Wy1vdxqDmWJvD69WSomtD8us1Dhri8
vwUhXWxOAb+7H4hoiEIH4Nh0iUvHrGOA4xKF81wdkdM+UeeauzLwcUOyE9hCZck9
uPSmA2przQETDUZKmzoqUAVRjL9vOuhRMbX3jqx9tTS/zXldAmsgTY1GONt4MRJG
SzjEsUn3T/fhmy195nOt6j1FWiqZ7jmGxwwEjtlnYxxKwQNzHzFDlzPbON3ywW2L
rD0uD1qEBfLB8ZIAAm8OHbJ5ZUQoqwauiOFB1fUeXRstyi63/FmWxuSW1xphpv3l
i3c5Z4aWbk9fFZWFGnlFPWcxGwEvs3lCGUg/Cn5CIl2S5Rgi8RhgVQioaQ6ReVEO
iGapfK2yDv2/3ObtuRGGaFTrl/IPsHsWJ3WcwDm/uycA4ie0PV07kU7ilq4m0GB1
ZkjHNl1oyRtPkBmjojSlgUDxVERpyTajxWc3en8j+dZTpGarjI70fhKURGv9/GFd
K04lwv+mS8ImGxyv6BF9KJJwuhDDLOw7/YynySWHyGhPYkQDktvJxCqN/v3iuaMe
AmEwsWDDdV7iyNbRd92jA+r9zvNCrHSjFtNd2AzrBRZfv0cYXWut1AFVxOynB3qm
kivInhYzr/TMVRRbPyxJWJtQnI4GJisBb2RVYKJfY+NAT2/w281qnRPAMLUTQJd3
47OEQl40Ja28mieTnOhQEgluhW6FnXSIXjcJAxPkrod7mkA4KK3F/GNCBOWjoPRv
IpUneP3f2+MhHbVYQL5lo4W9VCmlxB0UOQfYiCEwUnEuAGxxXBL2ALMlV9DVf3dg
yddEBCQHc24Bt70qb7V53hxkBoDvKB7NBCpQFZerVx3DbycxijqNr5OnnCaVQQNB
5l7KaxyVvIrXwS2Qp0yWSq1w90j/tzHcSeJAQZkQhQnTDVlVOl5itbldqBo+TspD
wOqKTBWUBJDXrIEiuYOUbfOCnMxUVK+C47dfOJwwodnF7SrSha+637+uV7zKiauz
tV+4bAEkZ5xArTK3ksgCnUfIUxREH9W5L58Y5dsyGjiwVCZ82dw+kT4s4RUDv+WD
yQi0q7ZselYfbLvviUoAzr1ndN/qO/va/i7uYbkrH9020Z5u02QhpCOShReq34bI
rrYbE8EE9f9WPMlA2nuoOaslshFzwsfOFJjQvt1AaKfveg7dk6B1JBmq9+9c/Lay
Trwcwb3qJZP7+1p75kRhXVMNGAAOnJndRTK1NkGOzPQoFcvmVIF4lFJDglHzWdiz
rhtLsEOnc+NRmkYw+2GjmQ17kFNb5Fb+xsP9fJ/2FSC+Cgz61u9MNi3RJCJx9gFG
Vv0DED/HWuFwGIsxJ90JJXlAitJd/JUZ7QuxnyndGienZ2ksDk9FJW14ByqUjPmq
pIVW4CbzOhzvTPbhUZeiQ2H493Gr7NH3KKCYFE49/4jan2kjTG3wbADkA7bM9Ds1
CEUfLE1LmOakUCzjeOeVxKa6Ja9sgUKZ9TbuoMJv9LRR/YJGUfpDrCO3JLWQnyhV
dYEkBeh3rHlyznFbURTqJtFgOlmo7sz5e+/ysAcOWvFt5HZgkN+S9FABHmjbodZQ
iOqfqJIOupR6OU/w5oA3DARXLRrm/s+5mGvLLkvho23r1spxNfZUtvSrz18t7lky
sJ4v3xN0zMS9xw5OP2jPqe+aIdKfZ0FMSjrqCsDPbvwgystytIJteuWR+pWaEVuM
V2iFVHcqhDbaA9HkxjLtY9W0wE/NvX14CCsqGyYb1Kt0m51XD9yUXCup4Z212uRJ
sr4WBZpjYblpcStZpqIiVWnncnY0uZPnzOrazdzpgUVTWJYPBaoytMaq2s3AD9kV
1es6TiSKJRZbregJB8oqmkKWcClWmkuAcwOCZScKnuDJmTXEIQbRMcJBa4S7s+48
eQZ2GkURzcmFmDe8NwO6NCRM6+b1khq/xMFXkCpT40Qx9IiqpiKD8JZkJFS3Ly/F
3ssvSLQ4yZQgOWvgWnaxZaelj9cqDq8zvO3v8LcuJg67/oodA41D61ocmNOzTUDn
47izb+Wk/yFPk8kL7x+Bar880jN5ziW87a7u84F4LRemfKgU2/esCfrtr0ZPb8Lu
8JRkuGtjJOGXuGAAMgS8i/aZsAh5/YY6KwcHu6UR9kcOcRYXi2uUvvduMP18yUnx
kKnerjfdjyRMAmkKgiNfFzI1tv3opKCAtdURoPuS4D6CZsiCVy5z7IJnauOikbHJ
IhNloMwD2qcqOozWtuhHT3vDGBzraOqjtrOxa/AjAucbvbd0Y6GrssE6/ptf3GT/
JOLlJw2GGjE5Xsmr4JX+k2cBX9Js9q1lhvYAdUFQZOXjoUmUVs7M/y0TRFvRxm7R
7mnRKegzdMB60lqTJnnIKcN2EW2sHRVSUAboYSmv5+IK8gIG489+8uaat0kEmDrB
GfLdEiCCetvrUn3TheKboKvcAFkusVSxKoQlB5Li29p10sHSVlEGH0LDM91FUiFJ
bC6NckPxqaGoDnqhCXqU7qMLA6i/oOYq/o0mdp/LsENfmwjSdAUURINbHbfOly2F
9Xk6DQEIl1/vKMofqvm1lR2t18VGkMmnc84PqJRksvg9VAoV+GNFrPb3djtXWOM5
yHfauT+Bg93K78M+hI+kGiwb7Ey7Zczx2Yf/6fFBA3Ss5NrWzFNDEYKAO9Irf5KR
6bVoxP8t2Vd3PSGRWMjLKVebXWcs43Gk1GaygJm1ba5Mkz4g9+yi8myKggeXOoY/
F8haPlclpVgRomxdIvb4h2IYEsum40rz/QjX6BHXw6I1MzLzS3UlzsGPsSoPuIMT
87G+SgL24VVO1jUFHe4k7qVDMwFkAnyFT1SwLF2A2utJ3bwzaxlLhOzrYhaD+1Z7
HbSniw3glEwiEOjTGBHC23R6ljOZhSl66n1yraG1nUqqmHwMYxgyvoUVY5krcora
RZ/gtPf8etm0aBQgPJVeZqLTNaEtqw2l8UWi5gKQ22evTwcBkURzeLhYsE/07A5i
ciAwe646TE3XgdNRgloZx7hdZsx/fs2z0HBB7Ri28Mtcce7id4t1MQF9JmtCt90q
X3f2YfJe5TqKOWcALIIeYwO8kZnpt00ETXmhbga8viYcM29fkJMF02TlkCNUx14e
do7bLtGe3Z47lNWRV4t+MtmesFjxeOM1R2IcIx1nBgTK6OO+JIYE13lobonW4Ea/
ezXTrsWyQklgGfUnO8iSegke7OnwJ05Am3l5mby21r+k+KkghQqFGDpu0w5fjVHS
2qzOQIzuBvmAJUCHebgDe3eSv4TMfMkwxnUkY6nH+9C+SbPMyrxAfTYTWTwJvBtG
z3ZLN91Ddp9ETxvb9M1v55nxT5Q3c+vpRwmd7to7bwoV574O8l76BwVs2maif5du
wfWAv3jsneuXCIi4/37WyMv/cergYtnaHGGY3iMKLVgogxd8hH+B/D5FP2nVI2my
72dtR5Zn9uq8Uu6r07PrJXzE1nyX/ZXYycHIp/1q6NxhEJOifYZwvJ1IBjPIVE4T
VPpPSJdRcJuLF6OjiNSq6dTlfN8Z2VcEwToQ8CZlAllyWhIsXpOmHfYYHzEe2I+K
djJQzFkXMtIIDZTeGYGlKB0a+g848rQ6InMKKcE2dt5DAO+19nuAKr640N2dYjvS
Bx17ekkpgI2qolHH86lIJJz4mH4BRLPDWp/O5COMrXfCcjcxeXNSD8in1XD7zCPa
xoLnI/8kVxbLH7XO62WwziT6qsnKBrT5segGIhdSGaeJ1YBI/aJ1wDj6BPUvZNnD
fh7b5CHDBo8sO9Qqfc3Wvvosb1sFquZOr/fOxg7TAVMkF4c28BnZKWYCBF5J4VMS
CgdXNHXVImGUGmLxGZA64i4jtUQUEM0UFES5mc5YFpaJHngmCFjQ+PDgl+Vin57g
aHOENf/nWGCgk9SCTSfR4fSce1/qWEBbju72JpMCdpZG0UWlf5CNmDMCmldANbn1
2A5LqVmtQocaK9bYUd3jNW3qKT0o9T5BYkSdCUWdkaQoSS+3XCpuyaxlUFmbzxGe
fwj7SLr5p8m6FuH0Q+BvEQjuBpdxMmC3mfU7hRVzIXRn0mhmWOtoCW+nIlP9m554
AENHtlHzSPzlGs1LOicexWvz5IK3TGXrsL0VNKk4eV5LdhCOmp2OXYZVsFFjDADs
cAL/93LHZkyxhR5SFyAVliRQFxPI7K7ClvNwX20PVjCnJd+EcqCNF4v/N0Rogpg5
feYEKyID8ilSiyPULHTC/6T5Dqf14Ft6qKrkbRYErjLZntTGGXlfMMgSnmR7bfkq
akzV7w3bUGnpXRMR9l2d/Mwk6HTQmlwLNEzZ/ctmaKtMsm1mP04T6gFz4LpW/nTH
U7swlAsDJP093/MtLvRR1tzJ7luD4BWRR6jInAGtqVtCtgHYyye8BNUzZbHcq5r5
AfqVHO1mxXQHmwvdTPTGXRygRSS2+JUFYD3JE3UKChV84/Yfir7w8Uj0nffHnCRn
XbG47xcvCTE7wvoMO0Rzgj9h2kE+nAlmC0lVX4sACyrOMkU8d+srzpv6lrfDpHca
dB0/UbM0+RUcysYHELGlYmAVzKlzvkITA5losU52JSIWYuqt+R+rekegizwJaAZL
y9iSNDp2Gd1jSilQSvVWoBY3hc7IqRPGascf6MrSCli1PX7WTfk+2BJVTQdRyw8r
QHDTAFrujj7ippYsLFMqEHc8RPPWq8HAsWGpGol0/soUEzhUSjHZGbzGASsJOPnC
JuMR/lSBCpciZG6e1OZ+3XZYwryupNZ8bXMC8WD2rKNtZxabvApKjl+Z3AABdLoj
eW1ueUGqalTQGDT4uerznXOLpPDFTwCL0wxbZygkcjr31cUWHxxEWQGTv6zzKgHL
E+y7k77aBnXQaMzT8PHlCiLFuXPX0MErP5S0bIUqAEoivBg8uR8SbqOwU7d6Fics
lECH484NwZEdsDs+99Y2Q5lMgvXYDt1K1uEx3mxW6WQ36TceACIu/BKfy/oQFseC
sbDBHziKqV05d88DN9wstcAPh+QTVRDwIBkzDKPz2wCeV6tpn9RqdhdIqA3ygulr
VM/HqY8YS28Xwyt1L6ECAqNVV3JR2D8dNRXrs/jPF/4vd3Jbi3qvOjHU+cyvcWFC
fCBsxU8dJt0rFKBgh6OS3c3U3gI757vEomc6lI4MBN8DswzEl7KkRN4JBm/VHij4
8fhZm8J0aHF6EwppqToOzczsWxWtPfhDAXMqnRhRn/N0Uf3TPrUnfSuIDUBHIi9C
mZaC63FPyX3BQ8wTH0wjLffyVvQs7RHN41IFrZHM6wKW0bnXYD059KBd+6xuTB3d
zSbbWs6PEwivEjhowb09HhAOPnnxebSPiHY9tSpk//TQAr2T4pB343lCSu8+F2Zl
+NyYH2+dixyLBy/sPEfJDAk7Gxx91z5UaGXdfh6e0G6PzD4j/4x4CuVBB0gg/l++
f7WcyGkQwEva8Zu5IycGS9wfbxZPldYw6Mzh4XB6e1duI2I6x+xvm+K0P8mvwdw0
lBUCTECjx1c4fR0tkCZ+3/rX/WCNSOYiO71bJk6kAb+4kPLLpijNL9ZdFUFPMKYC
flXFMnSOz0xYP4Gq3EySd0/C4Mxx63UUHW06P8mnZc9lgY3+9CfKdj9y0frP7X4x
b3rRX43WdMmzdBmkCk/DhVD93O9nHSPWyehYsBnaE4bF1uSfaU8dId429geUi+ly
K5XeX/xmWDj1yXzh5n6c2R3kxJoc/CAk8kM7b2PmwsP1fKvkngXbnB84o4DLg30p
mDDRHT38f2agtQ89pO9P5n91CUWxz23nVzSNKQ1xkDhkWzeMS9sPdoHCqcbbbhWO
5UHvpLMJQmKcawjNHImWf/wg2ERVXl+7sNTucfMaFB6wxXPNOS4iP+4WRRibAc+D
8PR8Le6lu6SRWqZGhKT/iroYNYUPxJTGApgpYK/gs/aqRgM1Htm3dQ+csr9Qbko+
VQml6Exp5KWz/LjnHfuzWuoYEyjGMa50xR2cGRrXsZsYK62b0GOjea86wH7fMdDX
cBz6cQSPPxS7wb8sQQt6CEEJGcDmPCXl1sPKPqNNl2FGX8uclgI+KNsPOS89WfDk
hMX9/TmEX71MVww8YMdcwFC0SwCx2IywE1vKxmDANvx8xDHL5K+20NSvGoTgX7qR
n+ZYT+6rEpWYkweOS9g7an6nP6/QyB8WrKmUJTs6h0daKCkdpHKm9Y94PaaVoFTP
+HjaZPAwgdK8pKGvznfzYzsFYImjp10P915fp0xy1nHim4HQRM2tWEnkYqsnjeJC
fjtgriy9MyMT/HqBBNqVxUoIxti00Bm81FeuaQXBQRYsE9jRbrCrNG/GcicDwiyG
74Pdvwn4KpYeSPI3o+bF696XZWdh0nFVCU55vD+QpwDqNMlbOPO27e0T9YJArGlE
gQHcKVu34IOwkoJvXsmbatjHJBo4NNecWm2e50vJQWnA+j+egw/tixfd5d7lv/Mq
WM4HwdDj7Q/iNcNt1Et3aWuIl4udqfjvOQVZ/kwu0+ANcd4Gbsv65ry0iMjnn/MN
AvydORx0x6m3aErvfZePresR7qesV+aJMS75hBYd7E26lhYqIXzD+MjCKuD22TjV
W3p+eXY8+/fJfWF01U0BEeqAADwXysF9r9smYUY2X5zwnsJa/8B/hS8bBVIwPq5y
DXgabIiKwwRCnHS4LKkC07OASUCGgzzUH3hFcjWj+Zhm4iFP1oe2Y2VqjBk6alBS
SabaTZSKUBcnX+pPiZqK+NNWKKO+P7+9Y48sIbauazdD+HjGYCDCLhh18R611PTa
wDAUcN+Q/EsKup2ovFaPK5h3IHHsFLIRBmf0IxSJGeBUuygWSpdQSHFOsUdgRUtV
E/OXvvYE/s2LT7idfvUL5YfW23HNyWDTsy1mLhK1mjPgfZz7GcdSqdyzCTiKQ76g
SL4GoiC/L+mHbopQBiRE7AZyXvSsNKqJtkCUCyIRQXGyZOsz7FOWJR8KPM5+r4pY
B4iinV7fSkn3ybZzbynoOIUea4OjtjS+xaLmQ1bV5IMblRMY0goi20CPaIvW2ojZ
EX/U5amYbAk9nkRQ9ol+aCwIv4jc6dZU3nBw1COwuaRBfgI/jxYp3X6ocgUHyTPt
P8odZRtKyVQq2YSAq9hRAlDO/RFP+U0rCbFmw+2UrQqgQqcWNsCjkMfGThblNs9D
2SyxGOEH/j0PryIhAC4JiZO2skPkAMiciy8qFi43K/OzeXcPLYI5dmb9sG5pRnth
bxaacqKr3uV7bFWOnVisnH/MbEGN8rD58dqhOY/Mc7awzInjQt4juQOAC2qS+ysi
xWOqvCKrLyNGlzudFOYJeAGxmpJfHsh4a3zEBx2Dv1H1Mf++uMD2oxOmYxGv8sJM
n3EdnK2s+E4zw4WvYq7BGrYXp00vSxXI/AtHYhv8RvgjdL4A8yzLaP2w930sCK81
rWgETXqB3lH3Sx8Q+EBTlwW6B1cPZ9zycmiNfzqsVb98H+4LlzD+gD8FAY8LpNKO
MuRH4aO8mjXrk5sFcFuGXlAqHGY54bikkhKvZlQlEdm4kzDgbB3IBRcVTyQUHSh/
u6esASQTSE0D9/uhz8CdLdqDlb6HsAjNuT9ASMnyKRhZzwsKOCgWKDW0poA0fFGC
r7JYcGApDQWV/lIEjYqI1fVc97VpvwBOUx2P4EXdAcivKtjI0CDpkthN3i43O6uH
f3YPtNvuSDYbYhtBTtPZyESeJGQo2+mnmcUzbdb4ouQz1vPCi5K50Up41DIV/W+Y
T5bKdrS82L7jhrpBwSz2djDxlv4bous7aRotjcQwbGhMEGuFYnqbJE1Otgr51U5h
Btrnq2w5FUVnq4HNFf6X/h6/XjNqMV5U+p7wlBcHzViVC1ROQUF8Xc4k3WBdSjWZ
FvtZei+ZXMP17EqYEXhZoOckfmDCfn1rM9nXAAsbxa5Fm8GTGsXfGOMjJ8YV9rP9
zu3gMegyLYRgEjzZxruc2INCX1lS8iq8GNKvBRg49FodNtyA6pZewz1vexBd7snM
9uqE3S9Yprp3zrS4fBkKVdTaRcn4l6RaW4IIgT6SJAAtUztvgXnJ4VUTVb2/8YXG
is8Su+bQY74sZmIdiNFLLmI4LOWY/YUJHEoQqrqihUCNTCFdHCNC8+IhXC6MFkq0
Fb1QavOW3DzCa1HF82JtmzYLGaq87MuilwIt4vliWScQPaho1ptD1/80cfrr8tbG
pfaJIHXWeSrtV1V2Bx6F1X8ylCwwzincN8sNE1OhVwLNUS+kQsu4UDLoMxlewBDb
bvegSr6StsYiatP0M/nvBT2nhvt3rEOKu+fqb0X1ahcphcDi2a5OKnF9dVuHJ9Le
+RlbJgCfTeX9XrIJtvyigDoF3onVBwKBwel9JmNBrwuDvdeGYiFM5wPCoQg+r9HI
2u8RdOpu1sq44d1PrmfpNq0jcBmlf7IEDwkhz0wu2cI57wuY7y2rlENhHv+rX5ve
VuTfMfSpggkMTDxjCJqOcD7B4+bcmHOKYosVW6+fLDjaQtrZjAZd1WSW2hVdiIc8
wL5XKW0tZhC+9J9oFHe8hEV/TvMkvx6zM9xOpVcrTQHoA2E28CCiZ/nTPcmt74hQ
wVwnZR5wOguV9C8gG7TSz9Ru+B8S/I48j3T610opU+28ITTrMxqvSGlSinWPue1R
LZONItL4GPsAVWgG8r8ygfsRgMDcsM79gszUByE7mCwaQOk+jvYWOCji4lULwpBt
plEEa8Kkx91wtub75GadkHhba8z1xNt5T8/829fANoLpPb32YIaxAaqHhvrynC8m
7UQD7x3zv47RyQob7vqO8aAWA5dBYDj3e1EadewVs/YnJdPs/mjMazPhqOTZk8O+
0F6dw9yVs51W00MiplwKe+yVRnCXksCpPw7DCzf5UteZYREZINeQX+cFVICyO+6Y
Si+7w8r1famGKMDC5eF4y6lbC0drYBGLxmUOubWMNDTqD3jW+J+6bBDJvJYc2Tpc
in7P6mTM6NasZR4+C0JrEc57xZImsighzsdRKhWhWJnz1CqVa1m38xJ1K/q5souK
QQTJKMz7eF0WEx4mYtYqnUAteYwA63jmPyOW+bnnkBW2I1DvT62TGyzS/56KlY3C
JymQlugZPxeWl85rCDNy9a9tqYypLFmuWoI6+iFw9y+mSV5M54vzjVujCjMpQl5a
SGNIfCGE3zEdLBXWe48XFCcVM2vzBBgTJHndgARgCdgbG2+qxDOGtknYAhq4mupg
3tlmKNl12EgCY1mEqmMTUMeSlc4MOY4s/DxengbUmVn4UDlFIG9ufPYnk2sVro90
zklNdN9eWSPwBmKTRa8WQv5G0bYqkISW0LnBbXzN5ptICsntXZ6z6UAgqIm/+aXo
KKanjF9XMyDJvTSav9UNRY2C6Qqc9lJHs2lZA61NFfVSlGl9mXT74LZ6ybRoKAn2
dcIwTniyOx6JUDsxPHAEARXph51KMPoMYXxLByysWkLGgZVilwVioEb5yPjSvDs2
To3zy1FGgdF4NqfFUOGcakRBBZg/mbTLTkDzWIbGeBUV3feqttQrOOTQBR4ktaqE
YjkMJTuoePzKRcGiDiNJXg1fpOCpoTjAZgXRgXYd+T6eDHTtfQvk/bjQ6pCM3zNi
e3mlRCRvtXkUqw0+41LRrAI7FddxfywVVADHa/n+/UdI67ZYVkOYD9YYN5Vku+WM
UoJasvn6N/kKap/4cLoXNlZTHWSM0gzfPitZQ3WUNJIfE2kdsOxexNbe1K0Bdwrb
iNDKnapX6xcyZLyX7uYWQje61FioCeU78d3tVAL4rUGgfMYlwSdghbCIqaOith/P
uHQ6LeCN3jbPRDv4mg971LBeJU58hl4M1P8MdmkQzsRn6Bp8UMj07l69QyA7y2hO
QXBrbHAu+fWpPRGDXBZJ7O8vvrFWP7llrUcLLZaCjrCGUomh6NLVSkaUDHKB5xm9
ozml9KgMWu9HEv6e6CIuadsA5r+OmErgdX6A2yxGn4nJgZlTyCOBvP7YQaaXiLcl
eeW08apE/MaIrkfFpkHkkSadOmK7QsZ1+31lg5VH0Lv9GPEeXZWZg20W19uCszGv
9S8vEuKte0I7oubwYP8vkR3O2VYiypUhqDSxyXEE7uF7gDWegJwJUcJAvN17BOtq
a08QqA7KQir7jZnbCAxGpn2TssCldZa7HeZo9f6OXK6eXX37U24hLEfJv5h6pmXN
h4rGwaPhgSTBYqJVNwis9RFTmcnIVFfT/nVUM3fifOcCP74qPjr/z5BSgfP44F7m
CvsabsLEGozqrTlieYSA7ax9VQlZ/qh6eYu6FeomeDcfMyPBGgwvPyarnRcd+uZw
xDN5BaC3HXMhwKCycbhwDIZEKNnMwE1GMjJQskkahtneK+7LVHSP18wT4U3yepDD
WujL1dp7B/nTRnpuxKsrhHhIzGfC8WdUCipCHk9R3FlCEfpp1tuwcFNkzVKgfWUd
06u7Bskupmyr6N4Vq8Rrc8XS0AKHa2RFN5B35dhDr0AvyxFEQusLXMaLRjJLJJ5a
BTw/akVo8Ss+zqtQetwAJa9v1lRUgq1Aj1Gx6CoJmdZzEQwef42J/7k6KhvEidub
zl47zGjp/YslCja8wBAJAmgWJZl3tpOTU3gkW5iURkGxtWDvlPHkDmQkB3gmGFNm
2KfHNRg71V8fKGTS2sZG09EMnjDGNWtbAjWBMzKa5x/BRkrTzJGLmHt1KHMgT/Or
VeFoTM9A/rYo7ukOds9sR0bF4fUIylWJHoqm8HBKTn+/z59Mu93CPIP3iw0NlrPn
pCdvABvZgZLsD5t6Jn+T7OFQfQAanyud92O2DQTdG6NY/dL3Tp9lrFBc4zcy2Bhj
aM3HDPf2nFmEkOzaRmD4N6daFtqb5fUa39xe01b3ptyhdMpkpncEEjHuqs5u3lBA
7rq0HfIx9D0m4eZBB8fZmTwWu+4cvWUG3vbRh4dc1l3/UE1BoSSPiOOJn7ZgDvT7
z5+kQc+NMGKYHIKhM5SmVp0wR2iGXYezpeuVsg72cddjItD1Z3dd/AYVNk93s8/A
bEgmwVDfBXOVEJw4wtmGVmkQdNbxvharxkMKaObD1piwNXU5oe+CBvdoOAGLqaQN
C0WM2hHRhR1gOAZxzSbCbOhbtydC5fWCLMTjnv64Wf819tXUR7lEnDWH4Yh+W0YD
t8geXdhx2s4D+wiZ+sWHLzclFqnWHhhYbLs3v/C+AMuRWedXaTmZ/yeB4SgYtWBK
Z3gkDCK1wFYP2pqwwgY/+NX8vqLxmmys2pOPjSELWfkEyz81JtINPFGrkpG5j+mO
MrY5fVufaFQglNdmjHhk8jb+1YK+fBjGJka64Sp/YYt7MEaTfcWZUeLKAnE7DVqB
zw0X8bb2CfD/cQeyHXDdWZoVx6aluhQdSLZFxix+KC3WNangjbguyZyjEEvjsF5f
qVPT4TgZqfx8aCVaSxDR4TgNj25IjtyP5dcP46n9gZd93i2jy83HPdqyevoHcN17
/rIxa0H9FQ1OxgHhJjzkbTUmvnDTrNjIxAz3UJ5mTjKLzvyZF8s1U4ImynAASD34
Qx/cSYuRKuZQjGBvSAOCZNwSvPIsMSPEPZRGcXwmmu0F7gzOQpB1okNzrQX8l+bD
FPMXXuJh/gfODW76shLlf4GGugJjvM+UfYmK4hcoe65m4GAUJ69lzc50i3/nlnjh
wr4aUorhgfNLnVOInMjEtq9ksvauyMcjtxemNkGfCIlakGtM9HdZh744YMqtxlXz
06v4sB7KDAWXbKGOSLUU4yZztDjTMjnSDyfAXsZ1ZeHvDFLa4HUKEeFA86MWFxw7
MOxyCCQUBXFS+H827l2+77ucHJ+iEZP9Olv3p4CkPNKIM0n/g+nDyeR5zl9SQrI/
PEoxFRvYRItg/WoAuAiY7LpSao5UxHsrCQKP1m+1nSSNK3wxLt/weGDfseUEokz5
NXHH3ixWXWYurQ83fk/a7HHZty17niDNU4GQkyrh+NePpagAU1srQiu/TQLCbuGs
xmxcJvOEBIGShS3vEJjjWhWJoz+dIm2ObhP83WKSBbQzz3tRSx1bCZiVRZW0E30U
fzQM0cB1+YW21Omys6Rp01eyF2QunNelmaeBTP9CXHjppSh/6x/HRA2BXMG9as1R
LCISa+gXkSNWOV7rLTMZqpiKcoRbHZW2Z4svtWmPSYIDGLOq6FJ4XIxZdciIv+nB
CNStzX8XWp9EWJcbd0GyGvNMt7YXCT1/Z0qQM6Trsved3sX1lPobhdLiqCwf0jS2
czq99CId5Rt17Nhm2/ufvcAE2xA7fkjuBGWOs53/gkdIPDe5M84HNyEVB070FkDr
2H410lEk1loW7PRH9xQg4PpH/LUAeOJ/YlzvOSUhyaPDPU9Aw94wWdfu00NU5AD5
W9b7z11I07i8IqQjJ33hsT6raO0xxom8AfJZO0NZZVjvi5aFv6aI3kZ90H4aDeKT
2M3ryxaH18J6ckLn7lErcs94NTd1Q721ppKDgUuSPELcXWVajrcXii92uFgubYef
KMKMol8GNbGyM56w6bOBMLKhQRdQ7eGuQB3EujpksTqlluL4K569Che6iLbYhMNN
9FN5w72V6KtJI17yzdRESLiJv/k8OhhJavOHUc4mi40TVSszlp1DxFxR4waLGXoy
zbdlBhfEYEuvlHizYIHYdfHg9fMDEFDRCOIeDJu4Py43tke5A+oKDTNZNWguhSnj
a0GUy8d+I3YF2xf/KcrnCydsFhzw/JFMO5IAyzSXCI6xgEDnjd/qzePYVqBqCUbj
5McCtLNG33UsyqFxHlONSJrq+l3qQIGTvJ118tia2aM6aQQbxFgRjoAX0VuN3Zix
nGBaUJ13qgA9oxjOeK2PNoik9/Zm55KQm4TsuVBeCGuxJnjaUm/eJdt8TMsXGuR5
6qp8gsRBsEPHQCpvoPYhOi+I7rkeir7hZ7cl4K3IcIFstX2bUpA1vDMN7Yvepu+f
acAW2cY3lOAohagK/SoNrKijDRI5eloOmqcGUQo6nIilIbE/Zgy8U5l+KGXsIm5d
er/D5NrGEQywucYpYB0NWKB+TWgWh+scSWoAFGchqf+d5hujG1k4mWc3m+q04xo2
GHnCP5dGvlqLZGtCBiQrd2c8rcDPOrOUII1Hsy5mc0sXxVXUw1FO7gsuEZBQPt3G
xbxpQf4Cclpwt10p83I6Ls3FaNFbWR3wU+FLDBvFzx2TSn/eorEKxObalCK3aXGz
+ooGMNboXmahb3MgZns7GmZFGQA8XZN8XcFEKqm0R9U2XMgG3YAx7mjFuVys0Gf0
fgDit97z7AZmsXliEvZN79KB+82bBBt6WWkHmHHJS7cMPsygNqyPq+rQQMuIILLy
ZuJJEXSFNQ9Le4DLmukWvpNVV6pJI6yhuGh0QD21DB4eID7Z2w7w2amyH4RhDn/b
wQaErIp1Cjed6GE5jqhPVm7MzLSwZXGsBlsB9ZcMITMJbs7y0+UF9ogNoD/nrhFK
zM4JuGmIogNVrUBKnIUNrdb7MYKIAWguxR4sl9zh/pKlWuJZgbE1k29j9/Vnohg1
68Io/+07JE2fXEi20heignsCFjXRsrLDyoMFEhgdoLFRr/GdK1e3uK/nrDBHtv55
sjsegXH2NpBCr3fOAsBrUSbNfeSyrWfQa6NwmAsdOZZrO4bqruMQb9YBmp1C+1or
4MNV/uNg+6U1NYbdYYzIRksXNnTiwiP8YliQf6+rs+aLfmxcmuFrDUxhJIS0Rgwe
ERnOeYMZm16ApYNjQbbQVRnMYWlBRs48wAiEbETUeug8Mq8W8fnlx8XljXTG1Ite
ICqUOYVJuZyGMq4IWfoMiLDYbJ7RZvC8czoZGAqaXIAc+e4b/rSTGsvXJsdlnBhR
rXpV+UaM5LRWVDXcgyYnTS6ifK6Vm0rG+eWw2cSBEgqo8sJo+xxkpVreEcrxArJh
jKV+eRr1iJXllX/5xfTV7Z75T1RRYVIayPuZfadrYmlOE5bL+hgs6tJGaDFgmxR1
atj0xUgU2RNjEkjopIoSpC9r5hCTuPQTRE9ISdvtx9JlVMZJBFVwQKLYophEtSlo
SfNa6pVTmP8feKt4PlowMnk3/lqeqgdJOxACecNCFmmimZ4ac75Cx9DkZvZ0JLWu
+txaqzxZw3Hsa5Uk+3LDBMJjZTyhN3sQTlkPyNskxSKMyKri+XwTJ55/pAyXv0Se
b0rL7GtDRysYILV3iEbxziD73kP1/kV7ezoGpTRrZSqgOOI8dTJCDUcFzW4WiT9O
pc7XnWRTrth+OnHfuxL8EFyBhRCTQAAAtoCnTmP71yuOsQCYPKnuyOmHK3AG3M1L
r5+UCbhOYwTC6lV+rOWa6k2xm7hArXdyBjSJLlyauMvQxDmB3YJpW6v2LZ+/knMU
YG/CKu41W6KPnR92x1Cu1z4g/K7tA8dvnzxmfJfomB3lStrCgUkvUfRscGwWj9ZL
vtwv+8ZOvfP+cWM3fbtHq+erVjNXYOS6+t+z98DSAPUZFWFpeW97PvpSf92MrqY7
WWJUC4CflSCWVY4rcsB1w8WfSdJp8ofiq5fCVI88BFzMYPG3xjVQ/Llf0RBcW2nw
IwSYqUFOoqvVTc+FKS1b0vQxVSEjBS9s5rJtA8FXtY5Ub6HaLjTcal2j3keDVNBZ
ZD2CMSWlxbclTQOpUtmoGzdBPA0MFws3GTy9PRV97pKR86lQbbT3X9Y6hfaT3t8y
2c4fFkcHZUwvWlJeG2Xobm/PJNoqtclIqzSCfygVNpYMR8NyGwF3qOQc+xgYOXSb
RgnAlL6gBN9IhlHtfW9j2y4i9qAwx1MABrLgi3C9z84RNZrQx2NDN1X2pMCnxJEL
siFfP8fRxqz22MOXWYTD9TtHBWXpSZqwbqJkS2Rxx7fDJBDaqVf1zFhHd1Mg1JWO
lFoJg60Ub1aCk7XyjZV3hcM9IIQxNgHDlDiU4dAxLjaBDFGf6z6mCDP2SBRAyu7/
Tr1qrhbrZwBi15TMzQxLAsOZ3cPcWgJhJc43hIQaC63iiC0Rijam36mjHSqB6bCu
+e/oxbKoK2ggdIDixiPjqinbbRichRafMCbfgRDTzdXrtoQdkFnY9HfiWnps2jg9
Oc4lR9sRizYMfxczRL7ZR/uDnlyEMIYFT6OSzE8gMYJRKjHw01Z5itUlWtVdqsDJ
gxsOVVq6AD/vLENT3OLncTwJoLXVDHy7Yi+mBmMmlKjncu9xSoSy6+0/hzwEXtWc
+R5zaox7c/0fHI4zCxiFTYVYmfqzGM2hW/A/I1elcbwZxjt4bSFWTh4fsUr9BG3L
o0ZsmQAXzZirhHZ5uKAJcVQ7oi/pEVtrL7NVC34K5rAja6xCE6yJPievrgCh6ROJ
4L6RXoCaXTKv7uKWvKeH9lgjM5S+aAXqFr8wU+AtAdap+HZaW5GUp5aTxybkcfWj
ManyZC5am/Mw1W9T6TPAAFh576qYKZKX4TIKDpbXu3ObEYfnYoT60+2ty3yqzJWw
17oHYcly5chttNQkZoKeW4Zp2x2+RKMaVNZ3gVEa0X4qAK1Hye4krmKBnFZ89ta3
OQ4q8Azylycppp65aQF6Nimz/IT59XmraneZAYSY5GbVj8FPDd1kPX+zJA5fQG5n
kKJ9DUsHyKLzDT22tLg1oVgrs+ewv24aTNr75gJfsqABkutDJcM/vyyopI2ReQgE
59ZTVnhsnorD5hoHuZL1IOoiBP0HxUmsnLZJ/VdWCf8W7rVzoznoc/yIb7hDQeAa
X6Fi10rBIgu2wI5hSPoa0LdWaKM6NTtjXVvnhtZ4mIRx0nxnqVd4wMtiofHAlSIt
5PnEeNPeQmQCwHcvi9711Y9l46gAClf1WFTvjtgAlipqFbKux0wQc9owe0aeSLhh
CrTZGx2yMX5OCORplSsQJd5JExLfegW+SezvcjldTAvg6ZRdvKLCoWPWwcM4oy6E
2FNM65MFe2G+H1UfqgTzxowCF+BLlVKlqwt13kiIvFAI28mCGGmpSHJpmLJYNs+V
1k47SicJ2wUUEHQCogOGKxM5+m1fsw2h9efWNb1pn2Xv5GFpr/Y1bKLwa2YINTZ/
tisTg9dyr2PPac0o9TVKwtTTKNsxTdt/qZYq+qJmiQlauIQ/Gu01h0ROlkKyCJSi
q1aZrZg8+lVvLc4qMayfA9jtDxO3T0BwcEcWxTggdookf6UPjA3MEMrGMln9D4gw
IofH2R6WwxS020ygG9T0EK3mo38i4a/4xOWSvrFC8pv/YXiLAsbRqEa8qaqxhRpO
BhBswEPY4ARKFDOxBfD+H9OI/1+6Zvg7YGYe3euMXQ1/+DraxE9ba6FyGbr0WG7o
Y5KCxzjglMznDKgJM+TC0EbpqmhoBP256rgBji+MTqXX0K+fqbEl3Z2b0zcDTWtP
vuf/yzKuSue5Y4uZZR9n4+fxqOiYK2/92oRipYsnN7T46DBtaz3sbBupyX8qc8Kb
nkA+TnY/A9mIfhEiTunYAe7SD4+hKgAVSltsORtzYsmHypoL2CulkChuzKUuwHjj
jqNIYTPg3PXKo0Q2Kbqtos05lXCdDc9kAaeobR+ZZfm0xSElyHDxuMAchUIZQWUG
nH/1SY7PHqPd/nsYep5KvIrTnwOkSbI4qYcZbRadlkRWY3I2oQ1rmJYz6fMOz7ha
eSZfPZAD0trBHz84WQEOxxRXR1jbUrV/Ztzyl+vUQNTqrjRYY1wG+V7bamkcVj22
Vdj27BOdtlCf8soAiz+n5KOFpc8yb6SNzkmOzO07pwszSlmrl1S8JM73UfIqkuZK
Hr/LE2iInC1yywci+0imo+mC65pIPL8g054AvOMlRr51yOJU0MyxXL3yvF3NqvY6
IEu5S7crjQm3wnipKV0PSkwtZcAS5f7z5jg7uDYttFnUtPCHhewDcfYmVHMpI1yP
ZG0rPlmMWUVyt0kC4k8Fsm0P9pwnk8wHtX11P78uPS7vsRAlKpulKMxYyL0Y/cw3
PUE8p5X7QsZC923v+iM7D59b7aU8+PRkQDwrz2mpP92dkVWN8aFOF61EgcKTrxzd
R3GseRUZTxFl5VMtv81NkD3f/xcJFxkgt5lnW6KYYwEtMpxiOE3UO1VKgsR4ioWD
Oc/zju9zAN6PG4jwz+9UjlJ6O6xJYKBNBUATOPqFDjOitzEZWkXefIRLsxJL9pmc
+z8HA4f2EaGbrmqkqAIPdjrB7upRjaXHBbuPAI9DhMZMeubw7RrnPoWIRxUAM3d/
3iyx6sT+BOADGKB0fVpw+x5nwDeBMUsywhgVgwbQ8tg35CUCEh7Vad5mKYca7PEh
1OlW25F8iwwg0O4A+X4D/83XKDzwlsjTEYm20PR3d7+tNn06gjtCWMqGSMZe8KWW
20y0w/ykiX2Y3WYlTh7Gpz4dG9FJF5JCqGseTQtc3nNAM7tPzTPaVQBwvqHNcYtM
rJz/3WZZ139YKolFmqsPtgXg0Rty+ctlp3beLaDj/iPGqp/4ELWFkWgnqW+sWBva
jzLVJ7lfD/4BG/V+e4n8Msp7WmcUKqVdKRSsZc24GGqKw7Jj141VPTqh4CqcKbfq
ZsD322fQD06CjZFNo5VZXkevN19lJgIVx4vMg1VxkAO/X2QhzOkA3E/PTgxce91d
8XtjH1m4R0grNvGo8CKiMIT3P8pBXhN7p6E7tgHYm+4FKX9fSZerMXQlu1Arrd5w
TvHJJZfa7dLlyjtSMxpjAnxV0kcvGB57ey6kYW5841o6PpB1wxFJfU4uW+liXoAC
+6k8+r9sNJYxLyjkG9r7Ei9DSwonSLUW+CF2iX23UAFkZqTeOiXD8//T/NjyehoC
6YU63zw+XL0dL+a+dsEcLT43SN24xBH9T+uJ6xhTP9riIfF2lvMqoY8PZ3o2ZjPp
CT458cMjqRUZx2U+m1dt5LYjD80h1PVsstfncvPkl/6r3spTLIaKMVlmjSj6gQQn
9gD3ROCOz7BeN+Q5GT5Trksw+f4egbPVbgB9OkSjKxlGk0HvekciLSmzasaXQ3X0
9InmFL4ZVwJ2IjBUCTPiICdNgQBErxX836IVEEcRkJ59/Q+uohbvS3QjvZr1yF5Q
dCtnupkjcPxlrvzQPKCMLYoMkrevS/3lmdiYrgneXXZboCvY3B2QXdeKPdNBRzJN
oRhJdxKQwJGtsIl30O9bBEbLYv4hM30X9opwXUphjDIb/TWN9yEWxJbrn5yH+Voy
VB0nXlxI7/mpj+Z53SKcNoIrodF7HF+cCt1MbxGfnbtvigfdU8yT5DV87pHKSoTn
EFQ9GErBa0m45XkWWFFPwananjT/lCa8mifOjIPiyI+wRyHmnrCh9xXGhxIrsvcW
5tCHhPM0RnyX1R9xzMSl116WUT6mXCSd/GNes9Vg/5e1pmfXfJW2z6oJB0T5ZjQw
SZhE7QkrfX5dEAjF8uMxueO1dk8KyO9PW7d6ModqYqTGGjuhylJSBYZWMnhYxGd0
cQxCZYXZXghfq9Q5xRnqa/jULaG4ppTBw0wvlrI/aER8LMgIqrkT4axfAxqGmiCo
2gLL6YaN/QH1U3HYM9j73I3nMUqE6t4p40YQpXhhWzcebevS9N6QnPiAG3TwlZJ0
ln+6/P8DOJNmrPB/DdwkIE7OqG2TSHvGS/Y14lx7CQAr8QKIQ02g3XF8OTqDhLaT
O6wNMQh8W+YogYmz7Kj+6xFeHQXRBXCqJMn45EVe2xgwrCGJmw0PideV9PBNMH8t
4oFl9lyFz/fAgIwU8PZjwfSWyGuJECVYTXVW+vSvR75HTkM5wQjVyo2NujgoigR/
TUR/7m/VhbrRxP72EZTr7PNIogvuYZT2OSkYcA8JR4aymAFwQ3wzD/E4g8qs16qY
zMgnF3dcYmGbX94x8bTvkcZad2pAgx6vaW02zv/CLDnBVxU3dv3+bDdt5huIvswA
3y0kE6vYZxwaBAY4vkI2V1JytF5lndq+yUd+kqsRmbsQ3OVjbByVLNHE8AmUzS2I
xiftJ1mT5K35WVmdCTt/F4XF/NOD2eAgRtbGYleHv1CuVeH+9sMrxaJew04BZomq
EJdyNgtC+cz4Vr6C1snJsnbb6Qq36kEB01CPNSLMb06YVyDIje5ViT7LGuGhwtFh
3tqoqlGRjH1eDmN9Owm0iHIGhxff7WIyNceGnA2FCNbPB/E4PjZGKwweYpbLR8AU
nujBMxETvZlHLPC4LM7M2YCgH29bD3oZU0Y7ThgadDIY979OPDQMFZqr/Scw2nVZ
N9uPz4EP2UwnN1U8rP4oW4LeZF6DuSZLllv8Yz3UbWBsmrUjhWlos0rkhiOIRzUz
IMwY/HQcm3iE8ivjdrfTf0uA+P1p1Xs/w5y34cPIDoGHDriLDf/zXMFb8ZvpFFeA
iYeJlRJKk4S83HJ2fQQnL6xXlNeyk0x14oC0ntYlcn1sYnb32IlphPGthgQrAM0S
P+P1ufy8dR5TFYp/Rdqib4WqiRNu16ZNrySRmfnJr3Mic/I+4YO9n5oC7s6h+yEp
7Hv9NxxcsZTIuZvw4xOBpU8t+8osr+Jbhtgdpv1SAED2CluHD2OxP1jhUhL2f4Rl
2m5a+nTBN2R1LeqArjqJFM0KIOWvLHpGBg95LNmHMLyeYjqUQ1DAmv8+1l7PV2gB
ybzyAMU5GsRCSwzrJj+gZlP/Y5ut9sjlZoTRt0V61geHhdQlvlk3mGZsMVYRp275
KEkPMUSqkzemIPaixB8s2gYzhkoJYd8sw16bH/+l8KujOSlSd+Wp5CcYtBWwptfb
AnYJ58gdmj8LSYFOQ0NAnOLzj16US3gvc5/S3VFDktj11Njf/EKj2ACbeELsdDxC
i9BbBu19+BMzDZDAlvoSbqB6GPv4SeoCz2kaXhc9ybI6ZeHri250ejL966Z2cBsK
xIrWsE/GWMCm5aDIp6ALS14dhyKhsll0g+Xx+xbDNYsYfhHgON4gMn3am/Bet3Qa
CNFiITm/SZkIDQJckfejg9I3/g0B8Qg+pnJNO1WP0B9PZ86dNSXBqBMLYFE+TZKR
Bp7534Q/sn4uWSwDg9lbyf4SKw8E3Hs8gC61eTjCyjY++JBFgb5V0oBjXnZ/tv/q
+kEsRv26XK+rvW4z718GKh/3GKD+A7p+vrOn3GGr60y4Ih56Ytqf0VLIDKupxAxQ
AXbq61uP8cLvkjF8mQEXuXLNYaDxiHG4hjqIRXC1GYdCnY0Bl3JyuOWvP+n030Ca
6/wtpIvJ/wLEinXsMrqkUl3eFdp+AMDNtWRX0sdG5/6OKo6hwDshTTE4clE5vQXr
bVzdFuP8iLkLe7MQ73ambrE3XzQGrI83ubjd6hYECqoZRg96FqkfLxYCMtztJ2gk
kq8ZrZ5ICNDrC6c4ql/xiRSB74bMD+x95ewuALZ9OQf+64JhO3hmORsU2go+4fn5
qNbc/Uzayc8MzEFps23BLdoeKzGRtL0K9ihKr2iD0M/yJR6I+LnXUbpWcQjxbyTK
RXg7F7X2+0RV3bjKekz0ZDX5k3UbJD/cubHX4EhWMmm/3srd5YXEgvBFxCZv+8OI
h6/uMvjt6jWd/CahtLn+0Tu1rBxH85qsOJyUqkuRdPb01rJ9xjGog088hZ5ea8wY
ornwAoT2EoeV6VEeRop5xgfejIK0N85QMc5AcjjybKDmSVGmJiKRJ0YvIEPgDOog
YnHz9jRAhVYk4dBbo6sLZAHq+Cb111avaKoC16cSuO8btk8RnLV3+dy+6JFg44ry
eQEFv7fjAsWkeElJIQ/0uj5biLD2W46b22SRaCTcJBL785mrEC3GXS7Epd7XNeRr
Ezizmv1YxR8kgsZhcTS9zJef1Zk/mIIoN5Z6xDtJQd1vx4H07BtzgvNWOzk0tnKE
Bfn8hsQQWlOuDMUzOJ0YCvXvOaHx6vUnQisKVvS38lSCSTzLsjEFlSp43AW63dKV
TlBoVce1tWVcsdqM/D2HHOzEF8Gb10lSbJoLNDYrobe3GJjCP0WkJTmQVyeSVWPH
EFhJd5flX1axjo4erulSS8VG2clUgKvv2Mp0KsK6NsLrH9xZPHSKxlQ5F69ZGfTk
RSt3L8lWDqaPoR1bGQvwGjlwsimJQ7T+SfIJ3FYosgp+/YiSjU7P2eyZHkPmBza1
9BHr4BBUZ/SLBbFPFXhi4i2rfW2tZoPYJlVY4rgA74hlvMFD0LeVzPJNMsly2lqP
2NyWsfOHPreC8uU2+Lt/ikcJxzBv8FRjDYwbCueQqji8dWERBpygeDndpSJsBpR8
MXQ+cLDur46OSV5RtVUHvwFyv81U50XnUKheeeBoBHLmgFffNWE/UrlN6ruTBwqc
RnPeWtP/yHfAwM3J7l3DCUAViA2QHN8EbWsOh7LQvgCKHTZ/bdsZlA9twiA4g6p6
7EcUihbayK9SDVHQAevkiJTbgvJ4nKQkAMbkRuKVZ8auZeND6RI/F3EZQhMAhkDM
lMeD/TZn49blpR14qDkLyHrXSlHC5ytOSVFXQgpdheUKPnaFxqO9Oost68OfTdvX
vtTDK6mJZXq7ap3CUiCqVR9zKo/22IbuGyvvLlCYcP4BlQFzmtCYkoVCx3MY/ctf
AW3EnmeB12tbGw3W/lrDoYCxM4y3GIAvawsntWw67I3tdHdE+4JP9AX4v+FIVXw5
dOQp3Szy+uzLri89n7JNS+/QlgkYWvHqqOPhdbtAlk0ToAXjB0ZVdNLlIzJ5eSFd
RqhZVZVcwTO1ZTLDcgZkcmNY0S7MNi91lNz5Jo+NCljp19TKuAS6y9BKZm/B7PHl
/YxkSg6mAQQY7MQJmx1TFqAbtVDnvUBAfy/HAhJO19mIpG8sO3y2GsmkefoGCqUg
mYL7ZB8yC+SPNO72ZNcPwEUNgSm76PzM4F4u2mH7JfRmZ2h+WMyDOHZSG1YmWi/F
R+YgwCklzPPO54SD1YfdMVZ8h58RtOjubkijIBKRjgHQpJkXRdFZC25auArmREWD
8EqO1ebZ9YChIpRJf1DjgcvjZ0mGWiPlNz+NvI+bwccbpbIZGEpYPuhTLsrFkZlq
aAq4Y9wGniPxk00zKfb7wijIxJJ8IMGrsMDkiL5SfqgKZ1qiNereR+sLSmoPpOoJ
C1CFJZEo1IUT4vtIGtuVLTGxDEIl2jO0pXrnD3n6TjL/e7B+fIL+zsMegzKILEP9
zW1+C/o+YqWvyvzpZaNV3UvtDplPSL6cV2Iwj33+RjcGrMGzDCQNBeyAESBLk3p5
UKuTcc1voYGu/dqeO1PRsp9MTxLjVpIEMtczK6PnT0ZjoLqtJiAt76QH/VpRtP1u
xMwau0XiOCuGNe99KHuyfqkspn/QRZKnca9Yg5DcA9WUtN4f6+rgvgZ7Mw82seqf
HFbVllmvPlg9tLrqmwrcD05wlROaVrpHPk+yza05f8BlyOUZ6E8X22GyufsyzclL
TRFHk4n3zLUaXezNSPgziw9DlLW9inX9a41bBmyLxqMKsBvxaDyeXI26vmC/+i3M
q/uIGN9t9iKDqrxOJ0odmd35Ai4rqLIDOcgscfSRMpVt4zgf2LcLFINGFDoWexty
yf64Qf6iy4dabu++FjmbdQa2MiM1NIIKN/WCGMfR25+Qu1xGP7AFYjsLE/xmnUC0
oK0hd0zZOhwOMiWpBdwmSmZOA/56d+RBB82WrfvpqnW9tBpVzjycMmuiIDdTi7fS
s/PY+LJa+Bnl6p/RF6e4OaECdaJZtXxNKphmrX4Zu4e+g9yN0k7YZ3Uo9rcYAOZn
ZDrtSvnUej5pjgqjKYD5bFoloLct1FsUwfSx/db1xhLawSEk+vNUChIDofzv+rrB
e/fQKwCBPENP4WiXNlRsUN1RIXFd8h42eEF4Aia1j/k5h3tpeBX2gWPJF56WjpPO
e5DHFFjqWQYhUBPo6JiTd7i0p8u4jXb8zq4nZzC8Hmj3GQnFtrj4iK2IQhDDyqfo
ZNirluoXtedIdj5Z4RkSXn8njlangbW+00zMoTJFVsq2XVd0WWcuVPJZt5j7OKAU
AM1DQX5CjoFF+0zPQXHX7Tu5pVokRCCm7QbOEn4XE0a3ixWkYqiNNlpZ82nMz5A7
C0xrG2DGCw58ibBO4oVow1ujl+Rx50DGcFHZKp6xBh5e4c7Xqms4lIviXjxonBjC
JSHPbGr63loHTx0v7mH+uNQZzv35AvTxXp/dB7LjWCP1Liatdgsq0BHgoOzPzhbz
qP4NsTWZoCX1gRWmICTSwNLlEelj5kRMRfsUfQf+fLZdSIyNrBZaza4L/QwAlKrC
yFcF20oIqZvjv/3ElVd/1TVtsEseRhMEd7rzysZ9eBrsGiefIuvzsjp3B7lsc7dx
FD/v8SOku1mPmU3/MAaOm/sqJ5Sj1+boct2/CDIEGxWsjsvUF8e8dyozPpy5SipT
conSwcEoTvvoKs+nZVQx5vHXMcWXUqlLtjldfNcWdqyNKRuLMt012kCv/4PcK6UK
oJpFtxG1VP4b0Kjxxq+6As3HyooeWaVZYM3eQKCP6EU2Q56dB7Yj6PweovWYC/Um
ucaxSgL6/vsV4BzJRBNVpQ5bKMgFE1X7OwA2ynlbalEBXJi/ZPtvM1WgtFraFZnU
fEsgKcFJVx6G3oWY+hwhjOZ61+5oxF20dkTOWbefqlOEyqYrXCqRBry7qGAaJIja
uY2L2s+zCPotiIbn1pWqdpEixAlQMhMBuxUssmvNafU68LBc372YsMd118Wzc/CY
7xqNCSZ4ufpLnW8SCwAMTFlcKCPM74byv+G0yGKqs13fM5Kw3x+7QQr7COyuuizp
PYk5gWSe52oTYO8f0ZKqK1lO0j3rFuH6h27ZBrwMJfAlImmo46jaEfX/akK71b7x
febJWSK3dusI17C01hZKAd6YZ6iSL+2D7AmMg2EZFUcpozu6p1HCWF4GaGSXV2Ko
dzwliBVvDNtYWKrlfdPjWt9ajXwseqBk7GwXQcKtg6+7rXYGL9XR/+QcDYJeC2+p
AicDOlOzc6OaKS8kPp5wxGU4c2zyalHMaIQ3lMowP/eu99d+4kaqSL6et1Eu6v7d
gbsbzXQbWpAJtXacP8jPv3ifOmr2OJ1bQWJnC0CQ9DlHWe8wg3g48RDkpNrhztC8
qqlVpeMGUUQddWUSR98CaVAvi1raviZQAJPTW6xJrYsnBIjsPNAIOU9hqn3CgA3F
f+xdALeeqWvHOyjkBNNaltoNgK1sXs/wRJrjQJHLeggX7TpJNfTedVYy6SI4N88S
ti36og3nkoNMFTS1jn0uD/cpmQNjkwF+f/tcVhx6G004khBddzD58nmer/+eU50S
xtc3q43JduLS49g5Qp5tb/llPfhBnNex4lOT7b7fMu9im52hPMQ4oIDdBpGEEzrb
w/wv7fWD9jvgn11QVnnKFbJuDnUdR6HpINOmHeYYAv6sGE7tVGnsxqYbQyawUM9n
PCVTZWVmA9YBjj9Y04MM9/5gkz0ti2mZ+NqQuV8/gfqSztWm+eg07A++KhAgAY1v
yAaUXzH61W5ffZraLiRNQF8mVc/XKfP6cZ9E2zoeoJcXul25vz9r4vgeump7EGos
SBZmtgG0pq0aqklYp1Z1KPUxFQzWZSaaMDoE6PTUrUD9nbQN5papt4OseGY+2TNj
Jq+2P/i5HjbHPEHbB2ETx4M1TX+mxKpe8v8TNDsb75V5vhmt3LxPLO7ZuU1+NyuV
nLPWrYk36eaoOCyoj1I6ZCRADdcfTGJQpk6xPOj3Mpm/v2Asn3xuofJL3FrTOWqY
fOqu2OehBC1l/3bgpfr9F5aofEvb2ASD9zd40hk9VOJTvUtsgLiyIaia4FXqDpcR
g7BzHBvM65cs7RlTRUOyYisN8brDdX9GIwi82aI47a7Nje7sjrbYMA2dCVVws0R0
ES4QpyX++/6s7DqVTlmge0JiILY4BARLlojTwuSLnlZRM37m3/BT7iO065ArepJL
Az3i2tACNssj0pxA7DybBKt9kTdyGcVH7pCPX1BVaNOaQxGgp9WU3Xc5YGNX7qzs
TJdDxvjwWP3r8NM2iOIbbb1zm0hF+sYEGnQ0orexEVLENdBacY+/hEevNQSg4riB
pengGkXWt5eTPqOc/6vVlevrUvG+bxr4cWCegQau6udXqnHkA9DoRYJh3KwDGvkV
vGrVgeIqXg7WXgyl3VtEdJPMDMBpIO6jijM0uNr4qLdEwVosbFeZvB2+pxRGiUX/
UD/03rUIUKpYFnL/+wQuzb1QeB6o9vRnVN8G112jf2IKiwQqI2YoKHRZjQSliBXm
1fOUGhqWuUNivTRuyB7Q4y+NjYByax6EVAlDA2nWH84S4DmqqTyxUldwsdPi50yB
0WtJuJpJ3xPpf2ayUctbIogl9f8LG0mnfDkMPcLctfyfBoYU+ZZ3WhDq1RhSzspa
nB3F08L/xILaWFwPvKJILd6vxMLpxSQWXPz+86S7BPdPv5NUAYciZ0VLh8D1YBDc
NCNe7GU0z24PWSTX4Z5zK5YZZQKmXu0T56EkoTNALhB6OYwMD1auhNfM4lp6YQ6U
v4l2LZlwGpW/18xMMiS1TvrtrjF3hl4DVVEVVaZjW5gj/hn3BQ6R+3BmwVv7uQTN
BwvHQTx7BsTyOoKPGAdKhsF0SyTz0JBRTnzTgW8qVzNmlqYjXpGaL1ZKN4shbScJ
beJ+HL+gztwpjkK2lWo0IohnZxdjBRBQylp+yVosjZYOY4Xl+NBspE2TitIXc/As
Lf7MN5a43etPqiDfpUSMgJVbFPvgFLxvHvohoRrnriiI3MTRyiwml515g4kRw3Fh
pF15/Uei+YEcyEezQEJiw5sTHK8n8DHTIGnIzcyEzBpFeyJiN4VsaXIvCSwsv/YW
3mJSjgY3Lm09pqsHx9uhUm9/ffCLkgYhCQJsUzTF3X+H+fFCNRUx+UCKdPUJZ6sv
vc2YqWoNMl+vmjpF7xhCmOz8atH8i27XOK2wqxXl76RYeffov7axHKWvHOC9Qtu1
s9C6SIYbkRFw8D/eFsyXU9zKzhAulvOKNHUf7kopI3hLSaHoNq/pZouGn2I7lajT
Dk1wTwL0VW2+YJVyquTkjkuP0JWAC6rAjjD7RWSS0Ih8ihkndh/NFZ7uZil6oIVi
vp+APDrMywubK7/jfNJJS4KiLFSxpX88jWQMbhsFMes8RP/4XGbWUnsWtkaKGom/
wSpguzIdck5PajTofPBTCsXfXMWJSDadJLfCJ4RHkFyv0nCXSejdiKc/+ofxFyFs
hBhF37ZqZpWQJjK02viXOTa7SHBUe4OxP/h3YonMZCsiHWLLFn1+PODRxcQUyFHS
M0hqE9rryCHbJlLOopNXsRn6WYrSN2ThDEzNLk7XHHbN4KOjKka7TfAqxUxpW5aO
Iav4Vh28wvRddbUU+XYL16COjJrYK3gFYzWF7PIssoBalb8inj7eHj0fIks3dmYq
6vteQ4uk22vvCc1qJsYlg4ZoW7iDJMXzkcUZNxUIEaHLxH8EGWBFcc5o+J2KCmQi
LnItfNEzTbaHXOef/FjXbFPzcN2yvhZ1xdr3zL7aSQB7qiqT+QbFsQsSfUKy+X7J
UeUqbkI56Q4UFBzH7KWJq6ZDQcoWC0SFT9ITNEzTKQLFkLP9XLDDO67jxxE7KfYO
3hiM2qEZK7pWeV2OR0M2H73lMf42O7NhCKVpBZ3ilWwziiwO2IfTlrMBPXGlWsaG
YGQTJSwYP+n8oKyxF5y71eCze035AOMd0VBkrU/yvLCGs9xYdrLwwTU8TLKvvVSw
Nte4grPFsGlwxzMSDeAwmR9/Wtals1CnOr70nk6wKQYwJPsdYCsVqATezMamSWUg
VLIEU/HY+a3xmJyxqhw4C7HnApRN36BHoLL4gjOvNYgBfy3ug3tCeLsCVD7iAHHc
XOQOO2p+cSw+uxgkEEhFK1XyKG4mw5sD8/NlvTVDWcD6HZvrpQjtobUIISBzCS1j
Wkrn9GaQBBVIVbb5Jjpkbfh5ruonvRBIzuiafnRexFZapodiGTJBVMI0Qm8baOgn
zMIpO7+YgrESt+Q4OoYi84RLaIrjE1zoLcfDAiAmX7wzjp9TINNarN0EnSjSAmaQ
HLJOcy2ReKfcB7336QKH+eKzJNNvcyjbESX4TkeMnJw3HBLbAcF52Mr0JdsYY3JJ
yUTyFggJP+hAjVT4u9HqSaZOtvrPaIq05du58xrbcZv5vJq2JPVACf9iM7Iwg0GO
oHAQBar5RXRABLU6l+3WDO0HqATznRcfiOq4lB2txj26Qv9W7Z97mEqdLbPSbbFW
dzcKw3ReX7MjX9i8tN9hgaVp7iAnemjszkSYzK6uVGDbx7qJYVAMpVdXUxakcpz6
D2Gf6rdNU5NGWEdIECMKjmNZmoMMOjAy4OBtZ3N8Hw9KeTw6+PfYnjHlKaYOWv2f
vhaIA9q2f9juBQPFVRQftNtI8Y5jem8nzfB1O7x6eCaL6VQKljL6Ld9AfkMonbvB
+mGp2uxAEcyWf1W7TPg9bLvIDk3AbfoNxkT45TcChR6g32xI9F2sELYgkdsA//em
R75nRF1oRp4L1RpN2HqeX4b2gpyCtzRJlM7zq+5Iifs69ZVcwzqETbkbez9InqJD
TjpyJipNRURKWlDZpsUJMUSi5tJT0N39L3+gp7UJSSDvMoa92/QEnCWseV7cWrS4
wHcFyOKpsL4ZtBxYJM+gnw0d/OqpigEqo3pDXaLkEtdu7nWUWPlyE5K6wu5Iq2Rk
KxyOTRrE9u9CuehqqQzAAS/7UaQhS9/NIRLRll1/mbaHWleTFdJ0b7Vb3aRuiq3v
68okaNKKZabkUMWRD+c7iXJCocmVAElLqFp3rETNxCvWcOyJrRdDJgHUxFCigDrj
yVnqQSRkhXeNygBd5hH3V9mqFAV8nP8Z9twkdb+Jy2abjj8QJP8BJAqUmGW4ZVER
uTSU4iXxGOUNC6gDZvpAax/Yfp/UI5d9L0DcureAbZLmAajQuvHYbmh5FVWJ2S1b
PDL77EmONnQ5ialtu+JkHkK2qrd9lZYqqcD7E+4CTb2eycJ2A9wXyMrFcd8xCCOb
A9zw9ezbNe49xzFJWu2pEKAqyfxEMOlzRLZmror0wIyX9QdQlswasYZ5VdPkl2If
46yc4zAKJxMoU+nyKyzy/heZTTAwm06CBTp6E/BvaaZBlOyE6rhWHOPqcxkNQdpl
hlZaxLCAfj65xmkz8151CxTHnNxhW+2Ego2mfS7+7EsgwrymuUAM83kiGYOTWHUV
N82iYwTF/VPoNQE/yKE56lL6Pz7Ynm6uaddj802KAvL6T6+YPxvohnhMH3aGOX8v
lyTYM7RofkbW9gfXml082N4jP9JSjF+znTKO68VqXlhX/ZBZsdRd4Ro4TykaR5D8
6gre9rnwJ0ApJu69Mv8aNs5BZASjDaNRNXzS97fxR3/LvUi3YHgvAjVNVgT3347h
hy02Zoy35NnxNkMVImG06SDz3ngDJVXJZ+9NbohXFAUVNrYCizUkr1iCpZH3nAPY
0egu8xACFUekpSuvPGPXsN/szkdxycAO5dd3qSDVoAarWZBmQc1i6Aafdo5CTElA
B+lHL6SjFxXF9PDod7FUPua+fpH4Gzux1Rt23i/m6jvhMZeEhHp9vHx2Jq5X0jL4
3eJNw/3J2lr97Ruy3lt7SLXLku0rAXvHJDGvjY49EDM0m7VNzFxAIrZ92Vy1vQ/2
cyq0tfqMXBmKK+bhcFPLH3Ta96M8EsqElqMieZB2q0SYbTvErGJhYpQ5FhWjd9uN
bbJme79qJL+zNa8EDd+vI3J31DqvyGebS/n7d6D+t6Q/m1tfq5iM6CIVKzsBEzfG
zIrMGlRuy7N5f76+Y78cy2n7Af7Ysx1NWWnljAVE7/AIS+PJw1X626drFHcDJrUm
9anvkZJSxB/vBe+2dntu28Mbep8YT7zujWFDVnMUcDLqVFKTBWV3fKZvyeIccyLp
6WCo1PAOsQn8/Wk5qmhBujypHJTkbIns41kP3/0WTISCHnSnbLfjj/NyJttQRTYn
aigN0Gwd0UmToAm2dr9dr8bun2GHFHQpFUoFGJGkSw3V5gkXLYwrN1W2hH4sD6L9
S6WPtCttUCykPLaQxs03FnZynjeYcONWkaut7DG1skc45vC25/ZBWM+solx7lTH5
sRPv1yFHZiUtlyUruZueOAkp97Xop0Dad+d0OAdIPL4tABZ2HbIzxBknqAbS9YjT
0Gf3AbOukuZHpRE0X8rILiy6ZgA0FEFvg3E0l5iYHu2oMTbkRHDE7sC3Nm15OurI
fK6i27Y/DOYWMy3HeGRRbR5BM5hyXg4mpZMewSTSAfG9mMQPSr3UOHi+8HU5h9Qa
+Gc00Oa6UqJjI48OPf6gWzl53X7B92B0s6O1q466sYrAwS9IoPV1xPcYEKgneLcy
xvQvIkzc/Oq8+e/xux33DpN+s5ScCxZBen3Ky8m9mVpKUtxSdHp+YMJOP3b/GTGA
gT19TxG/q+9TaASj1AY9tFo9AucTPRxAeCD64hlaRf+m81/f7to4XLDfo44zvobr
phwD3U3GE5NddQPucKmZqfBGXdNrPOiCuwhsZxKMvxXFllplbnWT/GrpyF5kXW9N
rSDtlDFqqJNWQ/TWS3gtQlAUE7sc9iL1H/Qhgu7jSdvjYjvS5BxnsMIeyIApY3cG
CPFeIeKsGgFnStmIzamf93JIBOF8NZu6qfA+CDDK2k7k2JENQ9oFuTAu+9aUoG0d
e709bvvaENkOZ18rEyTR03SKliquKVCSx3RXX+Q0UvWx9X8V27DUiicggVk/6JkQ
E/plCqk//1pp8KrcvPwKUFA3qlhpnM4oufDGar3gCnc7ygosp1y03WqMW2z3piHx
XsFjHXVUoUwuwQvQ/v3NFsmKGtOALSDuq5ce2nYzAUhRncAHBO2HRM5W0rIxMgLo
2W8wZjJf0AGUozaUSf3nDk0vRSh18jrtGuQIml2YcltplDWStvu9fOv4CSW6L6oj
u3DGXbZcDWrrrEc02fGwbTjcBgve0mfjdib/gfebyid/plX6tRxBDIPwaOe+g4eT
H3zPRJ9zQNlJeiAgj96bNtAffaWvJo/BcXpOpxaql50PmxH1IMmYRTmOjZfJO/th
NK5RD4COmeZUV89NoJq0TJfx4wLlDDeOwzZLPCzWt5JS6mhvUe1fVTk7nrZT9CEu
x1SeMM6tDkETfvJqeRi+JtaDJFFLjekyn+y92+79aJc2MeD1yX1IB8mGoXIaWFZw
Go+HuWSht50KC0D7tFcPPNtzR4jxs4gsnwTd2IJ3ECEHp6w65OWTfG7s0L+Kg3ab
W29w7qpVyIcRUk7eH7neCjE9Y/zOGreOpMNlgCkQCF+KRW0Q3gL3TAWV8rbQ767g
cGB/+/0/Qh5D8Ge9qjrFcI6idlWFLTfRF+wULG7fUb5QnbDFVnl5LX/ks4KFiXeg
5gwwC4qDdLMRtdSiDF2TZsQFHT60I0J94UF2Wit/bCXDaoXE0zHLl7Y6ZHPH5sSy
nn2niD+w2TsviJIMLK4jJbK6vnlEW0bjlLr57ulrq42qetar/s0PqlLrKoi9DOpm
JebE2wuJrblExMkpcJs+1JfPzVKBIIJrVHZzYJ2zGHPBeUZKCj9z9CQA5C8+IXK3
esF0QcYg8MpPk5Z6ZJOE/XX/fK8xhaicwZ5JOFbvHQEetznMXzryfGQCIy0DGJsF
ZjhQUcw/+n77NmmTnl6rUM+5bG2Lo9HqT/ka9Iiacuw6JlQnWZohxEnIgnLYXnR8
yJY7INlHOy6+mq+mgh2iRMYca38LiVSbhp8xULKA9oX9FERhCcG1DNdPi6HSiIyh
g0Vq3RRd3WDc2rZPNmCqwuCeE6HBC3/oaAUPf9WlXBCvOwT/+iCeZWTJ3GH+8QIO
/4Mws3LcTPxRoP0eOdW+IEwDYcjlh1XZO2cP2o2tcyb3qR2eX54Ztm9hUjWZX5zp
8pIxnVxSEu/6tIxFtF0VNAG/U0aiDfUnhdatgtMEkHAyHO/WAseuuVM8nzvQDcYx
/gL2Sc3Y1ASuw9liNFwjonpU0MoQzBlVpLZZl75pnpDzIwZ5xOAw3r2agrJz4xl8
ba3pVhgUD4+TWPFY6vVn5pY43XKeAuBZq47fHp05kMfukuoSbB+kPdZhjtu+InIK
MKhvQciL3wiJ291UoRTvsTOQ9+VCOiIMpUhTCen6Xx7a1i2olLwhXDwBE8cFHU7b
X6HSkJxO3t6uLL26WcB8gxrM9R2mO9cUp9y+u6y7Ly+CXL1HN4IE8INCuhDc3GHq
ev3ffc9XBfM2ynmqcmrmk4xXY49PBBlEBnju5FCnEX0yHJqh6PAXm4+EOiPYIbmT
QAKecLzBtRp2UcZhs6sCQ7xuOLjLqP/JUXxx9vMczDCMJfkneUcrJNMUNZSLDFI3
wNufZJj54c9r8mSK/R6y7pnnf1IKST4eldlAP6F0nOWOsnxE/I6aortDKaK8YfSl
xrPV6VWSZ+LT8ltifjthmBozgVDx5iCf3AP8TMuSH02v7kDiM9kjOXdpIclRRKfb
xn6Ft1CnEdg+zB7iTBMOr9+jUB/btfbK3+esqEmrvHbgcnhx5T7jlCNjF10uD7WV
2AwIgJmbV+vGISmN2W+HCu5uAYujxjXGqCofiFJIfwG8YU2OWFfM5kJoT4vKi7A5
SlZEerXFqnT6iJM2QrK/TRbJyDCvmI/eOdndFuQHyQsWAC/gPlMmMvsqHFyRxtgU
rd3A1mg8fr59Ibq1XzRaS+DJ30+Y0u3N2PtlHrx8j/jnBCyXOLnke1+M5F0cuJ67
AcZquJhjFoAup2zlXc24lx5XRzxltZ27y8/Vla+YrAKdf1iDGiuzZuvpmlqfhQL/
nFuRqNkTwUh0PL63xpUOhDe6+YLdztbDsV6+tHinJhC4/i1v37beYnQQTQ2+MPh7
5rgCY7uLongsYS6t3B7KDBcmcwgYcbhCe3jfz0Yg3cc6T0usPEekmPOgcuak9Glg
/TVMmDKkBcVvxX7FQrdf1P9oSU8fl0lRjXnMS4tbQug7GzXzbbY89SzrMXRaXldo
sbbSQyzbcfKgorYn0+vHJFfE0bO2sObmrppxVE7JtVp1O/LDoFSN8hFCsG4fxmd/
StZpnaKqJ5i+2bBEDcxmRYL4CKBKAKk1/QvEsyxDhLgmUc81UJPVaLILLeSETe2/
w1ZEabGFH1jto3I0sUvSgprCtxSL1maz7XYoSlu6MrEu055HSDABH3Gcc4M6zwgD
WGj9XsQ/vnd/8qg15XdQOVLoZUmanEVn/5UiDRGyIIVKAGt0gc0y97BeaOuSWdrp
EDMx5NjghuJ9srEMe//AJlvRyt1SrUtfQPQ+Bnj8HFADY19Xc3QUQ4RNyiOL5yNm
kRU3mBM4141zpK47DM5WTM0saiH4rLS/X423EjzzR+/2gd50HC+4fRK43z2djXwL
uQhGOAKdKcTboTgmdENxznwj+wluPqsbArkdlhp8usy6v7icP5nGKIaQ8iF+uh7K
cZC6h+/UIzN60p1EIhF+EphPuUHexYj6WYhwv1+IbrT0j0+zFlRwmVskNkMlpKRf
Rh7G7gA8yH21wZaCMKC7u+7xkhzWAPn3xhsEjhg2Fq8NqtR5ZMv0Blhgx8VVOaoC
Qh2s8qiIvM0yjleBYfAkITVB7qn6BSauK7PiGdRK2YsRiJVjVnb85mcFIGpPuI/M
/8f1hvqmq54DDJfbJlm1Y8ddGCG3k/Wr/Zs7ltZwqj1Skv8lQH5PWSo+UQr4wSxL
I+R6BnkpKdbUEtr8uiu+8aoP3VDpAPfL8aHTayldm4RCVTdvTazXEkgeR/9cmL45
wiNk9AzdRoEuk9ygKmed/pJdOc/yI3BaHBFDOaQpqwck3QyHQaiXDf87U1On8yTD
wOhlIQqly68x6IP96CLlMRbWomSheOsilbwsqmw/l1ZQ66VscLbzhocMZ0yiUrPq
pM6IsLqJai32q5KfbF01TAmdT0HU/9+ByqiY65FQi3V6/cy8zVpqP5nsO9j/Cs55
wczE939B4vG9sGvMyxOUF+oA4YNAOyirPuOAGvuAmRcVGCS8FUgNsWHzsGWlLkK1
X3eVh0JnT2sVJq0X6P+n9kJs8DC8MObjYGvgbNbaDCtvEmi+L+zKImmbRJ1jmsvo
io0iV9mUMgiAsixwwNgrvVsXZtaJiLQSipRgyOitQy7t6LEnOG+ZtnLZ+IM5a0ap
F50KvrDYYnQv4kN58QBVNl7IwsDuC+mfN9TVOKI3LFim42RxT2r98VZrCo/Dn7qV
sVphBrS9V8v/TU37z1h0d77SismT4hSvhmRyWwkDye8WIVi1/AnKeSLpCYnmog+6
gjCIIvMg3dBlh82zh4e/qqvZyIgGplbNRIvzaMKVq7EjaAVtBya6pM2qj4M59EmJ
A9Wev/i00gaJkYgTK3lWi5zgdptX6UjfM7+rZmFcAOgyO1uzovCgBKYBEda2qQbO
uhTGH3k5ZED2F5M5+5q7q9riv5Zvytt5Opvupdj1icVHFL5QFA7MNyAgONBPHLAE
xzys0IziOg2HyOrpbp4igoI5zLnQApFdzqLXOTYWjQI6bQOL/0ALGQIMoNiXu3dm
GQcRp4s5FIEZhL6fv/MWj5tptBi+O/FnsoWRsrBgHR0p5Ck8JmdpsDWPTNMuqRXj
TklVoodqWtJdOfRlVnQD5o50zczMzrgQmDT2F8K5tQwwRlyZ4jCoM992ufbQj9wj
23zyje+CyF6XdYSyCfSOoyxrDpLMPW7CzWFEp5JvAH7rahkzmrPtgMQVnQhO0Jc8
aGummlLmeeGkxfzY69m2ZIHhzsZ0eqNct4BOZtrxRtMo3SSECPPbumV+gRupHMds
k6tamB7TSTBsylqGE9a9q1YQtAYUIs6+gPNaogkntQhtPYM6JtkFKxRUO6nRPAvJ
vVgeKiP6atOmgebghr+TWiGEDuUabeIA+a2Vgtuj57KCIRhzy6pwT7Jf23s9nuiT
sOB/lhHtrkk+ufFIRrd159ibhy1rtFX2f7L6pUOyqvwx0ZshTLV4l3S7GE3OTq+C
5nR/NVBWfaq60EkmLnjx+wTeAXHjYftiPr/YrXAUyfiXL8qg6cIIxY9rPCGDiCjF
qTnUNgEHXvH0jX5UfPp5zMZ+jN7bHZbIkdgrNhPlFYH3fwv625QrDzjQ6RamSbjN
h8d+okgw/kvR1aeN20HGikZdMpWBwjshVEqrYSrMHX0JH3/uG5MRWwxsTFCuPp8v
sDxEJQvvyl6IEmqlKm6fBHw326d72BZSliDk7Xvd5M2HEuudUHgzn/VC1um8amPn
67GbSg+shCeUFmRDCyr7fWQ/QCmAySZbZyInDY50eF/+thdAtV5M7Agl6syl2kbE
l13nbd5UOBJl79shyX9iAZlGDjzfaSbR1Jd2MXuhWkvheMmSYsKk55PXNvBiHmsZ
yvnCVJ6CyzrHNMWVMqElLaeZ/6VO0TQz5ZMAJAO1kfI4cbPI/Fa7GM3exahTJdti
TZmDsCva4suVN4KJVbYnM8C7f00lu20tia4ypDM8plEggpegbe6Qyfo6KGIbozYF
og5I8TLZUz2HVKvemsrul+ZCP2M0iVXIhLkNji2Ku74EXLX6P+dbEfL9TgBveRMx
gcxksoxk+uSKolo/BaPr3yFAkLb0IqVvaL6QkRtBdhHAriE2JSY+K5AyCp9X0WgH
0afj9FnzJgjOwLnG7VrV0UXZiWyB14IY1YTCNmY9Q2/oBt0bvcT9gLcR75oIldv2
Hzkqyg3FUOhJ+PaK0UJGa5Y6vUq5oXA0RrfxYRb0ZLvq9BQwcv2i7IB2GZqVovZo
qHdKNhYS5dBLoc1DDXUcV/C9yz6zF1gAOxTRTnkFxEw4CPb8g9QDZufTRGNOwLww
fU3JK1mT9v8FPEFOzLwbalZ3Yskou4JkXBmZjur5xRccAlz2NDCrikJDb/HQ3M2U
Gf7URXkLlYzoGNrW2DIUP0QRSQmCcc0sYClCr2xKP6cb0FO7/a5qippSkoBY5S6s
pmfPUxC+BcpBtiW2Ahy1kiT24UeFxMvWK5FMXEPMO0//fVzc8j7CGcB1FD6H+H7m
qZuvsu/WaBCLzH9/iWEBJJg/53OAfSIt0Lomv6PNOGmHhO/VfLrm9wOW77KB0hz2
jnOVeLF68k9GJZsI8J1qpYYEdKaki6OLpseN+4HCrpoS9NtgCapg+vX0VbFulQWS
tfJQe7qeUq4C4YUY5l7CScvVfTOEQhA99n92tJZ1i0cl+/0tNKAlTIQFa5xRIZ9o
CbiAEkNtKcq/z5My/6WIeIDvDUJb8Ev+c/eSDEtXCOIf1eiIPuZo3S4STF8n6+lS
FMp2cz6+5L6XOOiBrek2kTSP7Zbe1XPq6ISnShRGsHvlTNZEyDto5Rxi+n1kT/dk
gdCiAQhPJ4AgTkpwuJwkZFxP0N5JCsHzmdbW6JJGdPM19sbIfQWSb6PbXSdK+F4B
i2EPD22PGK7PkoiW0r3sHahLzmJ7kmKWftAKUn5/NnLYr0nBtgzv9teMEAoaX9D9
q1oMTj7mYFNH733uABcz99jzAzCPF5Gee8iBe01Eyf02P6LEcpr5IHVEmwMe/ORG
qoxVzVxU6gcphORHjPJ1/xLYZ9AEnTK9rPlXRkOEnSkQWauDa0a9j6krqS1DXhfj
69jDc7wzIaWtWqpaKlOk3w9b7OfSBCMsdOkJaJrgks/KNfbxg14qhUGGlZ3f55rx
3XjGSdKsi1bUMaVOv/BSLMbQRfR1n1hSV+hqr3S8mXl4X+bIZts8KwxoHhF9HTir
MZIBhc4u3lNMUHDJ06pYcHoExiQiftx/bp4Jx+eU5uQVXLCK+iruv1RFRhfGiRNZ
/dSA5DcAnXSq5aTNDbQYB7+dc8vNLW1mG4rm96eLDAGsDrwHsh+zJnbLkjrxCl29
GKQp/6kR4kf+37L7KU7Yy8SsxzHai/bNemktVsd4Ev3VhytHjBghL46AXSbsIQ04
TL6/VkaeSKZI6HCgMdcLFQqjYIFowkdkRXTEg+mPc8waw2sBoBizQRqKKMyxvSGp
XJ6pWvYT8mtb55glsmysf8xEu8pktiaJC7CGBIVd1AwMeZW1vIQnE1EcdPAwfUYi
2ajubbEN5tUHULqCOtnOYIEQmDILEg8AZkhU/xSCVFzNMMGs0kfbFD31w/vE9S6i
7hDtim/XJomlPEUxaTai9H0UZ7jQYv/w+usmGzaNjNlze//EvsL114iRcx15Twa6
FsO7BvtyAE4IsByH3nXdY7T74dK9G3Q4sGGaZF5zRtvighREVoKc594Jtpz56fU0
seZLTPeAHAuNDs1beGSlCpSco+OATlqwNMnP3dpLeTu2XAfpruGA9CTXhNVkkmHi
TfDogWTDjFbhgu1r1jdo6Yj4Zc6XAuEUeh+oJuQwBiyW3J3TjIb/cd7PstP/BC/5
fITzq18FOEW5yn2EOP95skNYAhijx/ykhmiKOux7ji/PpNA7fiokTG5v9x5vqsuw
6ZQXniNNemZ7+y/o2cXHfWr4eDhAStU+JSxcDvvjqmlBMjhhwkwjkz17kQzgZXG/
fOJIwDBvt5NgyLiCeXukObs2LQn5JnRJxsezCqdEuQ2zlVfzERctJW9CKKMBx4r6
zteKcplVNNEYlol1dOWWo1Q1ZL9SqPT/I9kZP+jBX/BxoiSRoKsY5d5e3jfFRQOv
newrSVc07ExUr+nlzG1uJk220ytoxikiL98Q83gQW10ZAwrdSAO+gRhVBUocdypj
OBQaxL6QBpVBgWeqo6eDVqWVO5f9RVfHRcPDPX56kkfU9Aza4LbeQNEE6n/69ZDD
NOxsvLVG9GlcCT+/ecPUXJh8X3GypS9mG6k/LeaJOWc+0gVJIfLDvpLL5hhIJ4pY
h6tiX6f7kKjkIsy8hB8gqUY8N3mULaJYvjnF7xFub3Fup9vjYHQSvH3R3doYc/Ye
4PjW7RY3YPTkQIF+BVL/JZMHDFyh2m5PhiW0klC8r1JBeKS4bXrU3lzr64yzxJtV
+AuEWuXdd82JnZK7gHpcskvLtgpHFVmEoGuSjx9PTdUUgcfJRkujs1f8pw3onSDU
N+hndNE10TQBQ3doY/G2/fs128AUhgGwMUp3UGGvbZjcR2yeyEUbO+gKeXOhgfVZ
MZKmvJsd88JfSHwGvQWJNOcgC9mIn7sPEloxkFbH0H20zq0meDKhwPNskQHqLQDd
NEdLhXCn12/Dc+aHWNAsJVaK917yUGns/DruKS0BiEWWB6C8tz0KgF4QOxmvhaPI
ZArGYF+FREHKlRHQ/UGoLDs516eO3+C4Y4Ikf5yF508SHk3qB3U2lN/xEk7oLfbG
fc2y/C2X+u5YdG3U2ev/LuqwYF3h0GBPplbFLvZxOtVvlP00j7bMesEp7P/BLyxr
6DJ/shFOuFlGCFdiZwC3my/yJO6hX0U88F2uRL7hDIQ+5lnCmgeeEmIy4UrxT2x/
v06wktG7dtPNsT5dXOA/WQTTT7qMUC4yVTr01lh8t0cSUYnYcqbdjQlJDhpeN3M8
sBiHCjJjsRUHHygyNFUtjIGyfox3jWE3m1wYA7jWixPn7XYHciXE2MFOhBTYilyo
LEOMwdJm2EGuuWJR+REkfe5/H+zSMWDO7Ccu7uOLjskcelhHksMtImDkzt/glO92
xDAFWSoZ+0dtiSekh2VWsGGMGNgdM/mB3lXGvewGBsgEplBRe5g0qVzmavPrO1ZK
NR6pzbMAb+R6+pp1QIe6YHJpWt4vD93ARdTf3LynzVKGw28wZHAfhaqcw6NSx9Kx
RXukjyydLFoZ7ntItdJhXODmm+JZ/M7oF2kJJuCCbSgep7u6JcUsxwTpXGHGaz5q
OFszVkzzsPn39hQvZ6FHWJz2LSazCS5VVeFPUDH85N4yx+FisUmFfV2gZdrIQQZa
7Dqxvh+XDX57D+dvCUMd+i3iTbvSEoM7R6pcDqRJN0mjJZFwLFQ/hfWKyIKBlusW
5DQatSFQ106XtUkCVCKfZEVEp4kzdzB5oveQq//GOiXuKxS3OUWzGiPM98ZnU75o
D9kikdN2Sf9dxTN/VFZAJdf/UU1RqlXYo4YX+PLPFdK/QafGknr0Px3dQFSZEc34
hNZpp02LgI/uHpcIaFpJzChCs/U+1qGrh9j66ECHrp/7DKN3zZC+lXTIXniboOXR
XtpbK01K5TVr+fms1Nsb1kCW6FL6oGvziQzbLr14kIvcebHtDadjoRbq1L8HMGip
enUKp+dI+Gaa+LFwIdJzZ6KOT9fXbaQB2UU1QnKF+c08mLSoFWpfykJN8xgBabsz
/GiYvdNgU85ZJp74nfQYVMA1svk68Vt7QljVKJKIRNihrVOCdvp5vmrIv4r+sMde
6eYIWFBwo8ltkDxxMHxE+SJC67jsgnlu/BVl5OWjeEdBM4AEMeXhqjTH+GDKavLz
npyaWkepIblM2j7886bHzFaCUnJrq4TeebnB27IlmL9+KdzRNQOzXzoKXXeuOu+T
12i9alfPv0+a0x9MdfndrBDTgtmmVIHh1VzkEIVV1mLu5gkuQ3c4+y2XVtOfHmEy
wptWgOhQoEq9Ba6/iJBo139zki0lkJmwMBrbWqTn6wS5lmWgcWpL5/H6dtqoFNr2
/o+Sv0wBi1gCs8j1VRjmbFeRPh2b+oSYd6XwNfam9EnmKLBNhwzi9eyXRLuLBlEd
ID/ilqvjfD0odJ5tB6Iyr23Xjg07GzyaDYKLW5ynW5bTh4DlUUVwW5as64NpJj2e
YsIVzWWX9xGVGjCai76QBJHV8hMtr9FrhJsYfp2d5tuCRb071m8cyoypEoQF+IQx
ERFqoh3URtWCY8X2xc5B+z1aIJtrIAvno3oWHEk02sAM6rQjw+T51weqltep7oVF
L7s/3eoGtZWPgPYCOp8U5sjhb4vu8JVGCsUaB/m878jgLg07JeOYj84i/2GKYlwG
raHkDHFrpx/FiLcU5X6JZYglb83Q9aYgK21F+f1pRNBZ4c3XFFYsg7O7clEAHZXy
uE8hv6aEiXP53bAyyOzj+u5JSrQCXAm1Ylc3hOh/FtCgTrH3TghSFxcGlt9pGSZT
6nP4sLEgFwjXA+X2jH4/eWGBETy2Y37xaPWZFX4Vf/YsPLbblOW9d/Cp0QhjT1I9
IEsafcGtg66VPD0lYB3jcYZaO7eMGCd8EIxUCqy+zNwJJLm+MmeqKWfqaoVkxR7f
gh3M2ZU2uEdKqaSuVcxNXI8t6dKEFhgtrJrD9pEYZU88cVY9GrOuIdlp5i4UrIIk
FvjsSoWFv7X3Yi6sYtvC4FhC5wwuTWTIrlJREoDzpASniflPME3v6BuEuL8zW5of
dHsrWXbYWkdDzNciZeKfuVl8nSybBk/xngCTCM7xI9PD8rPKeXJRmq0vS90/E4Qh
x0Qau5j3QDxh1eiqLPBoxLH9c2JDxtEpyBQakY2ecsan7x82w3AHFVDRNjG0aBfV
4k/jsViJgjz20hsj4712E7FKjVG/xN51WriwhOeDHBXT5dMek5PeoVs7F58j6311
xZZMlwSFCjzBciMdSTE6qHP+MiWkf7/DnIpjhlw+K1/iTCJd/hKWcA3V8AlGnkrQ
Qq9O6/SCS7idq9mOwVz6OxGJEwGjQSv0yq1FVneXNndVCkTFvqIbI6vU/xD7SOq5
OqgYL5t4liXgFSRmPgm8JabcifnA08t4CakCkHKaKA/8kh5j/U8r9wW2HnILqxR5
aWB9lNxYIt8YNAlCAL9gIpqXJufSBYFUZv+a+pLyyqS+5vxMv1AxbThfQcfHRJAA
VQL6RuBYGk0EwicpLIjsUyASEbnbF41AriXU7yEzzZfZlo8GHd6DSyZzCoTbw5Yh
wHznxSzfkjs/bGAYKgeV7R41d57/rOPLuTTujUGXrWiGyFaeGaJRPPIUQ5IYTgD0
7z9ym8tR5BBRbAuXyrQBJabNDZdVXnMXjrfrq6xBVJ+CC2MgmqNJv0X9yK3DIVAu
fl8dYG2JMBH+XysjC7v4pU9ztZwOJ/0iUFF2rBcLDEv3XTgWT3OWCNfFDBWA2Lqx
8+LfaOudIVC9B2MvfMl58cOkXqOXBMvs6qlpS29eWWxRZRsQwOHZJl7AsNnvVF/r
gdZEuCdWhkvcxEJazcXudzRc9QJTh+ITZxoexQjKbrkNOWZg23kkInqikdcVPbxN
p2QhoNJq0jDyxktbzRhd7FxdHXMIc5pHrsCGtp+gR/gvM/IP91ANGHyGIq+OFPfB
Z8itSeZe5DsP6TUHrDYMcWoxiyAWa8Cc5ZRO/g2itf8CBPdgF4LEQb/blkQ7KFQ8
nqunecr9G5v7k1B5qwNH8f73Dm1Eqw1ovHt2JKJuYejS2VgD19A+5uI6jLFffKsS
+3DgnBys99iqdf7yKaIC8RLJb3xFxcrlQKOOnVwggG8g7Tbc1SE/rHcP671gQg9l
iy6GLb+E/Tp7Jc6uJMF4TDc2fNCb35FJhlydKc0aykblQCJG5l8xp91Azsp/G0tw
1DK53s2WnxFLuwIh5YAXKOGDrDmkm/8SKSogzzoeM3NUs204tw2E1FIYihJY7itb
Er5YJpQtNbqL4C0d43fyMMbLuRhQlX1mILgCU0o5XZ8UmbN0J9VArgk0QWiusLal
LvkWQGcIb28E69JFxvsu9yrLXvnbbgw2dCsMLtEkM8ChOyzUpEdEEIrL/dTgm8JA
bf1sGTpLa6Un2iZjyUlekD/BrNCOQTprwiMfKcEkzCjbif5hvm7rm+5UaA4cjvSB
onfVl6PgjT7doVYzmZdnk2/jjfQ5g2f4a/A/AzJGd+30QcpJyxYnt3+WD8bF9DdM
xNv9ni8+c4gg68geoRv3PqxKBH4IZU4XHAh5rYmvi2nybpwzaNuSQPyCxIECYKWs
jVgK8dF4GUA4cs7aCm7mqC0pZIoAZU4fy8ocHOJwGroPS59pXl2SHr1/s2F8kyii
JbsgtkEE+TKMtfrevF+/PrDrDQpHmOdCGfxyvKZGEFM/Dl0WnJlpez3hcYUyFWiZ
YwBrgH0LnRB7A6QWRwk7Q7GYnEhmkhRoxSymaExYboYIeTgIxynSFyn1OJx8EBpe
qmhC2xqprYu6cZiNQo4uo/AJpPklp4OJ42p/w+4csXDSU61N+//GKjvSLxkok3Os
oCpeIVZqpWdnxic2EZfT2rWTMOZ3PKwDNmX3qAf9zd6x9S/8mX3aCRyea9bqi6g3
B3LMPE+tlZ2U7cRGAtVVYDrNjfmBq/DretCM3NFW7NRfs/zi7ActmkZ/dSfjf7tV
GWt1iJIKXPS8abHFnFY2kNp+vO5Pc/Y9970kXOh88kaeb+OIrn1Z7EmObsLBr2dH
DWcseUPpjh9mduYda8UBlbj4v7Z0keYhzP3zFv6xNRG5eb5r7aHag29HiffRGKjC
on3N//XKjcqb9IcSNa6HLOIBv0318XAjK+kFomJpTiOL7ykhKN1BHxSfakpTCE4W
VKkr71fWtqGhSmAAeXckJ3JQxVYwcVC9EXACaOOi2ZDMdDVUMv9PFW/GDD0A0FJW
xeBrE0Vk40UN1xsUQbdOClYhIv9DVc+N6s0/YnzpIERoYQCOzMtTE2+26MyF2VMU
iaarNYWwPfYVYPkoTww9CsBKhXiH4L2Hz5zYm7VAGugbtxg6eFKm/vG4nq69jjdp
uvKgHMsvZsDb3MLPnU6i4Yp777ELiy5u5aI2/pBtE/jwdhzrgtFaeC5aTA4++JBt
r9m0oyifGdaKZuPxdaDaGBJDosjlRTyzXdn8jpl8irlmtkySYcfD8S3tC6H7AHKW
7Dej+RTtgpG2EVA2j8G7GiuudNr5Kv35V02hjMaiSH0Q1BgfmIIqPNSXMDlq80oV
mq2WF+T6xwAUeFwmsk6RoE8TB8UNCFSrw6POHCPJ67tciplSZSeL3t2PWSz25Xlg
sgc72o5Xrc6uR5quETApJaYil+HRvavITy4O6fKeDCzEJbSUic79VsAzbJV1bw2T
CdAFRgXS9g3FUXZ397wm6VeGOR4AjKadhV5sahdq4OF92EWUelLPOF0HWD7r3fvx
SB4xagOkqpNMdeuutF+pFCwLoxQWN01/q/sFqFGNSd6dkH7trGb4768mKJNCUKfV
lZnB/lFq3r2TVTEq+ZhfKOIqqKWbdJ9TEh+4Xm3pbaZ5OmeTcL+cQ7lvtcU2eepK
8MB0scCXlBpQEsIp+ulpzTaAkk+w08nr0xEjuT2/9Cwhr35G9p4hd8bOsXEYHGha
NkxcSrhMtTrvyX1vlOvjDTwVHCZmnXk47Dr5dvI/5NSbA6M6SLiVphzw/Vrkr/QI
EKLQWQbhbM48kc1IFC6F+CM2zirboPQfaElv0H6ncb/8h2C49t67Nh2YVPkWmojs
6CTuCL6ssdZTZ2SdTEVm/e46xXYcFi7ntzNcGoNKRoaqnht1ouvIb+Q7RoymIyH4
CARMZpUsJDVouF9oQ8ntxKykrpsHmKBYMtAXJ1phfU8Ofs8w13VTc+Y9hHerO6mc
YwRLG7JC12dquS/IJ+dyI8SEU1FbpVI/dCnHN63Jku9ZeDBI1tSKzGgwfudOhGRv
ZPuGt8I/nloZUCEbs49Gqru3bMU4XM1FF0TNkolu514qJYO0nhgjDOHb0q1/qrhu
9TrmA9zYk8K7wypouJ+n0uXRrV8evT0WnljIL3P6jjN6cOxvwOw1mo9FRAI+BEp1
ph8a37j3omGhULGwiLiANx3/HF4ALBmPIByA3OcEaawjC0ylIjBAVweTUyLjp26s
uSKYtFaDBfKQap1TaMF3WoMcPazheq4M5sMrhk6t5BnzOWZLBiQaR06BBzJAOEqT
MM95D8B5P0PNZM5H8k4XMdeM2m4qBiEnPvnTmy8DLyHvmYtEp88b53cZGojVTuOE
zAyNTIlUhYnhOYlh1wOYeJdF2zxGOPnBSFLPyRIsYg2fS440DFVfPkPH/km235US
YlhnNTC1o/ktQh/6U/PwwrL8r4xi20u2yuPAk4dthGjz0DKVIpxgM0MNP+l95jR6
SOOt7Sm4NwcNVVnGwR77UCoid0EGOJrN+oudR90Fd4MxNUeYCCFkc9fPHkzl3ntp
HrtU+tJwoHDOuRSG+F2q60ZK1kzFV0eBqbELRpPWgvTCR/VDLgfUvvGIf/g1VIJF
8mD8o7kPevlSiyX36f3GYuxxqkXLKsihyM216eT/HlI1+l/f3gqZNRPkrMxBBEbf
YYwbcer/Cy+3lPmrceWCaPNklES+wrDFIl2X0II6jT0zutmPjNzvWhTIGV11bpsy
9VqD+9UqnKjLnFtYR3+txWdN0gItXdj/gko0MRswEww46xCCAcD5ozwUJ0ooGP+N
kQymQuQpJprlEJwCShgWmsbAg1/L9NasS/P6kqBRWaXvxJ9b1qgQmPpUtoFREIdi
H4pybupfr8KxcJCLLYsNM5KGm2vOVsLm7D+bfu7ZSAawB8BUHSG+24539zmyzmRz
ccojSSbXAezhNRadPis6ysUC3snNkHdDajkrFqHbpHUv4seiV+JRgK9j0gGgA8hi
A+soZzKzt0+1DKGduUPFqhD912ldayakC6LsE0knJutyeu9X6qRNHXUixftqY1of
yU8wqnQ6cU5AsASKAjtCpitotBv8CftQoZHsh8/tWg3fD5kxkIe2z486Zvg4bU2O
9/w98ts3bRkVvGz0TWT/yLcs4uuzMXD+Q0ynRsEYdGd3plydeNZxsBRSMRBSTnti
i61LiuL92iuSWeXWvcUr4y20U+mhNgFQAeNJnkJXap7NNH+sdyTUzEwqjpopmPs6
Ei1Vkgr/KEk4kNpKJBD11STuRxpU6HboZJgqv6+nbQSoMCUiCLp6mwT5R8Gtx4+c
zO8avDO4E0roPnweXuYYgtFi8Rz0pU0APthm9gS1m9zeMC01SMOKS3dOV/drq48k
qVkvoEVScj+0wgTsAnfY5a+OyiWCKbh3cgirZHbK5GL03kGTo/B+T0if8t5mgcvM
qnsG5+RyODZha95Nvlbc4vnaivskR0OVce9FNgaYUT8u4eyAOLhdMUCJw0fOZgYu
24VzUtuKnBORC+lYWb6YZ2tqWoQ1FqPEuHGblj8haG5pszsYnuJ7gTLYORda5PiD
JPuZ3X6Kss3YyB5yUlpNJU3h+O0gYdcRXb5UzBxIGLnki/P8x/S4eoYh35AZV3ao
I4YElggJomamWzvdsCtl6ALu+L3kbAj6t+QWwbm6jzwMdd7mVVsssAjf/DPUjZZK
q4aBY+d3L4GjriCRhEl78OyK4gtSN500Sz6py19hQDSLAjWkVgL3o5oPAFhjZJjy
Wbf+ymalQtehj0YSW/1L9GXsa/JM0Bcf6cFlSHWBoZNgKh6eZwRm8QpMFUuRKrvv
z4LZYjc3WxdVuWUxpSvBMArbRuibjR0roDNVo3smnbezbD3zDT+vrHspUfga4z8z
8pF6PO/5QQ0fMkydJJYbnYjfA0nkMB4HSq8Wxwqxu7U+Pk4zbdLDentbYoDRlq3o
kLydkSkDO/25qKuZgRknlU/mgNvG7ktb4HHsrcDT7nQWS3cF8fNVc5HNX/AAbjEB
tH0ehSmmAFRwIqEHIh4f4p2fc2RqpuA11ESxmrqC3amf5Cr/H5axVXqrRbNjkJYS
t3eaAC3sLsjiIKy7M8EFowbHfLUp1pIN+CR8NeH3BTmDFi4h0+2OegOBNS98efD4
W4zA+ZC5OrqvnxnpmV+gBPGtr7K2N2ZHBALha1CaqeeeJ6Cy5l/NwbAHICJYno8l
65joQHtIHNuEh6hE6RtELqM1txXKyBFqag+oAOX2IyvuwDFPyXtlzppFq09JIEzi
JHLKn0mn13EGJBjq6cYbKiEDro8yUlNma6wFy26TbaqsYhIitZrVwrJLQ8s2u/rD
8xd8mk3F0FIeTOnZI5ATGddqDDCfxiaDGKt7mm+IGf1kLaZZxfh0tCiXSzOhx2q1
2V1SGm0ExatqsqBDxX9ln0ojfMOhP6CnM+Kkb2Zm4pFpXLWlkPdc4rkcuWRQ88Oa
1/xPT5YkuC9Y2omJETf+9xMu7WE3CkpXNf/wiGU+8BhdQndc0gqnFKtSPf08Te/d
uJpK/aO4GYdDRzLdajwD960MnIBQhdiwHlsaw1w92nPnSSMP9kLXgnv3NTJcwhD7
0qDFQxBJ7wYqiCHe6WezL1pTfr9Zn/uErnxj3/4XYg+4kPG6dcjNJ3cpyeeQMtzU
dgDJJzWcA5MtUjvFgnK3bv1GAWtCBxhVDE9KlCOpv/ItvB1m4WDd3VwjP4ZqYbg2
deV+zLh79/YuhY7JOAZlH1IlNlVVvAam0fW8Ow509ReOwQtxLE8ohlNebubwOXQf
eETK34oPYdxA+3Hg0wW/n/qSssrvYDBYQC/ZNL0Bul/irmJ60YSCyhux8uxaNPPC
bPWz4IYYeoMJqXZp/YRABeaiI7AdOiamgzRJyBYnglQ2BQ9vdYpyeFBEHNYr08wA
WubgYz9uRQLJtqgZxjrLH53iLMi3uGN6h9s+xWvfhft0bBcsgs6cZ87VJvhoLLr1
hXvChuTDqKvYen3nldnQqdMqlM3EaAtKFkadm+TbRt5HlxnI/Dh1WE3NrhJBG59u
MGcieDc/XHj/nTFLCOQ/rq0AZU6Yn2NU/9HSrAe0TDoVq5nXIsZ3gud1xzNNTKHi
TvNENh/i5Sgv8LWat2aW4Q5nOqcGYjFCNBD6wDznIMLSopjpf/4Pa50aDKvfeltU
rJNEQLVAd1Jxg0sZkbAeFVGpPAPF0Of+RfotAN++uPn6nOp3eh+gXdCLm6TWQUc7
tmNWqgxHexy2OfVz6vm5qZEHwzRhCu2EYXVgsvgroOuw5iDn4NRZgmN4fQOThyWx
i/j/7KdYcQHlLgu3F01qyxz9Buf4vO2ZqbLyHNkNSZ5u9s8IWlZ2MEONuhp/ju11
JhLpEFd8GYQVb+PFnfhsF/KoJoaFB9IdK9yvFFFWV5NWmISHxv1fe/2E0wNiNWiH
6EunnBAJJCKbIUAQ7jINo0y0XC36rlaLNUmhs4dMkIJysxxQ8i0yV+e7W2+z5ZJ1
iyeINvjyetbb5Cjmr5aNBwSZ0JpMzn/NUFa6BhcdY2H65mMp+uwjyIoFSbJHOSNY
IxhfBXHscWaVR/Gr7NWWdm3pS29447nbBpsDKxl/5WpefRkXA+C149AT59GqQf7Y
9NX9sk9hLyzMI2DyImLxX0hyH4TXtLKtrC0LqgCeZQ279RWB7jgG3y0BuwkzCciR
vbRq1v/pQWGVM2KSTYCcy2AoGEBRxwYi52qFDsBm+2JB/vsCOyW4ee8I229RDBd8
gRJccmYU9u2ftyWvECGVf+lWHnkywErVLy83pNp14QaDA9LQNamzmDFPBYo5NZXJ
wC4Q1LVsZOJRtduxJnlE2hzvugWp4vnEufr4IFvEg4WFx9CNGCzjsn7ppLu2yYfT
rWjnseoZlhDyRZjnDTMNovvRAdfgENqGblGbkUmIux4CIfrPCTS9hY3Nbiowhgsv
3COlVrisaH7NoiDfcwb9MlcuyldwaSmc3o0+s7WicpxZKuY4HQXhggIUx1g4KLnh
nHsAyAiOBv7l8aIaxkh6NU46E8f6H6N9R6wTcvq0FvAKYyAEIjvBiCW4iA268ldW
QmXSOI9zlsWQv9qxgr3xGXpWfn1+TRQD/k27Jgbcsj+8BwsxRbFLAgvUQcKexZvZ
79MHD/OJvAK1TaBKgM1PqTVDArhJyJ3dYWvlUR9fJ0Jvc1msuwnsjFy5wI08lWs+
FTv1hrrPQ7g2p4m5sTRDTAxchy+6JgV1HWlFlFT2nbCmJraeJtsi08606n6dQ2pU
sdTLUz7D/un44n8DcFmsaUtxAXONzuTzQAsOee+mS20HcQexYQZwwavDRXlF7usH
PM6450qQe/hRHxru5wn/Y69ymkni84kgS2HmBjcUxlOH+VUqyqpWZ7v+/Jtm7zYU
tiJ/LXiLPh62TWi9oPxgwxAXB2v8ABalCfyb/G0YPUomu8uGKzzxcfw+/SJGFSYF
uDgSghB10BbYJb/0Cx3nj86IHL6dS9aXA5rUDMTM07dUErWmaD1oPXQVDkxqUQ6R
+rZ+iGK5vk8sCJwBDNxh2HmXwjaP4deiwer6LWeMfAxZ+YSJC1Q5Oz+AxcwFrnBs
vquU5LgxKplTftIplxTj8am9wXWW88PL9SIJGu+JKzt+jysl/P2WT40bmE9Osp6G
04D00etCIK/PJVroH7KZiF6l7qAvdyd21FU45fJP5d3i/YnAXRy3T4lxPzpD5OKM
DsxLrMoJFYPWwhBqwyspS9Ea/WIexS6EPzguivcHqZGdnn77lWH5MQFkwtNg038T
Oq+Q9Ab6mQZVytFqxVOVmbFi/dWT0U58/6QqiKnVsjngDbH4KCTMNihYmNo0LrG+
SwHBMl+eMcP4CmHrOR0lJWAOB41XP27OVUtrZSGcXPa1MdHvdPr7JF/cPW/uGYo/
YJ9ZkoodKzfAuUOzH81OL1JQ6HePCj0Do+57aABs7JYnurAqiU+I0d0hEI7T2cJl
xRGuL2eJKDMeLlRvvBHzjrK5HJmWlH27Q2mvSAkrCfhei2g3mwEYWPDSj1mKyZi3
qWtCS/RkRpBfZO4RveynI8p9IH2xa3F0rTlGJMo9Qzqq7DPRcUaG8ognogsvjaes
hBo61/JGbPI9/qitAwCAMhgzDgX6Z2XMHeBy9wAx5VqrT8XyznDCi9yYL8YZQtYT
elQ1fMgrZT/ehUi20ENFGNQFnWPvgosFxMER210B15iHmLd2RDVWh4NCKrwRgxLR
eu6Nzo05budhD4SHB+hdfWxp5BKzMJyrKOediQpnDPi0rNpZIpFQqc5dTWt9YZsl
mpyxeALJsZrqSOsUxbXIOttA8NM0lIilChmyeitbe019TzmRR6VRJS/RaJOGzQzL
UXyq1fXLdUhq66AgPZuobz6Vb4lEwDECycvr9q/j6FORa6+7cpH07B1b6D/kCuDt
fXZuGcJK1C7+mkL1c2wXIp3rN0plBatJQFPvn2nhS2hVbSGDLx3kUJxvziEX7AkK
mZLFAAQGjEcM7osc9CK17AfLQH9qOVZk3ufSYKspivaOFT/Gl+M/QSL0ujOs665i
GCLPpYd1dqxLjoaTK6VxuJggOF0wSTaoMEZuZuIPrquKpo3rYr5RMPzXTMUl+GUM
3cQ16ngC0Ozs5i4ag+Qfd9MZm3dpKIYGS8bLjm5OgkAjHHx12yqBD5ZjAD8wX9gR
sty8xiAG86111P03YoaEMPTg+GR6OU7aC859/vbgHxjr1cFjNermu+I9u88kLi7D
My52KyEw6cgHbUPy08vX/uPVA1rjCsv1+W6MxGIuHfW0sYoerzifi1UmGMtYO/dO
amMc3HyYk4mgZeKZ/atp2egoC6Xaei456p9dJ6XSG2aldRQ32LfZRgzuJaUuS34B
P+d3V7VXC5gJhuKmwW+Hn6fQ7vYteu/EP5o+AXCsLCZHtFn/YcF/tpCneSSQ+lQd
jEf+/jnrr2ctkV/9blfPWp5c5So4jkJjTdg9quLhcuLJYAANTamxHH1OqoMWHve/
k9/18cy0cnlLcYiGIcosCXt9CwHxq/OgiczZ36viucQeQsHIgHbWD3AIpnMmkmwo
PAKWM8GVGvRq9ZJxg5x006CkBX/H657ubOeVeSWEJ6cRfKi8GdkBXiE124pqjB0W
x5RNfe6IPqP4olQgq+GBKXWvfKbh2Eya3repmcX7QgtDEAM1NxskVduXY2z6NwbC
XIrKuMVv5qdHtvPG5CiesAT3yPR+54HIkiI7nCxreS6qy6hj+ZG5gi6GDCREte24
3ebjoSErwsWZZ+qEoUZ+nhEb7vnwoGMH2z66ywY5/RhiMICPw65Qa7yonAs9KHQC
3nAshu05ZcP8CRsz39bTOxTYvgY7me1cRJbezUqQcPZKSR/B2NR8hd79ebijzZz6
kXeo4w1dycgogHmBogB/4I6lTbYPRrJwkurr6FxH7zqW84GYoistytnywJ9Gyi7/
Lh9nS9zxLq0RzxzgMusDmRBp2YAnbWWMO5PP0pR+H3u8SVrT/w0nZ0AuwyIPR6wh
H/Cug491gGoL9WuBmTE8E0slt81nrXeTCP7Nic+ltE2See3cmvXldcvh5fhJnepG
+Bs4DHPxV1TJPcg6NrWgo9RThvnOXJWvJbXvhBRTwjM53nEOoXRhI01svk/4TyFo
MZPk/AYkLKDaOBFWaLdPNzpdyXleuHgmzbQe47YFvDGrj8w9v8cacCBhLniE/yH9
/YPKUwc3pZbYy22cKs1hv+YUZ8xeaE2ecGLNw8PqjzY8KV7MdI8ZxM8MBJIfUAJf
IVMGexYPf9Ep4xuqQWQGSEqjS6IDDntuu+K4WR0p8b1i5qY/aRFUI3aBc0nj/hEX
W9qtu7xYSYW2to/Qcmk6Vad9ret+2hARGm3Gju4BBev6dho2kmXcDHAeISSxwSc4
RkLBABhXIWch7pE7RROuFEy0/GHiEVCECUaHE/NmvnNpuA48z1o1IhhwGU6g0Z0E
HaRFUMoAAJ+hWhfsWAl9NnvqLv3KhJeID545erlvyEP1O2GV5aKNYoSRj5TuQV18
u0dPpPJFQOgKo6yALBtza6Wg5R/2fjE3yM56lkHBZFLioodZMB9pi5kOiMH7uQ18
i9wYUmpFK3PbcKVCBSiUQL7MHL8kP0807eCjb48LAYlMaApYJmK0DHcg0us/+B/z
Lb9mbkYaUtPjXnbz/fWAm5KOeshAvdYxTg64qur7PTT1G3dkB7GMJPnWeUzVo0OI
3SzQqYN0dVr7miOGx3uSOercLuTPqSvEIp4ysJkASR7ECOqBQdZU8RKRiLHsrng7
AWiRQRyNweWN0WLfF5IV+47rwyoGqHSjmfKQi0CPAcFSAO7SyliukrnpZzkdpPfJ
NffVw1ZKxCRldi4ArkdUTCsqHqr0avAITgMl5kXcGO54fyh05U7XgKqgaxMph5ed
oUAGe7xSJybj1l3Xo84Qj+1k03YMdKqhV57AvHT3+3Uxa9jtyl2VEnK25oswlv87
l5eE1A183J+V0hn8jNFhQRxwL1kY2zVsYflS1rMDh6OfW2aJXhquuDfMepQ1Pazt
j+L+JHVjC45Jsb22ER1MhktdktJKcq17KXQWjVxG+qDhVLfXSiig0wyBsvdjG+YN
QiLrFUQjzid3i4SjjrEiPjApMv62thy8rt1MXQx5F+xFzhMCbDpysnjcL6clDLmv
pNka9vdR23iPDA0W96I57jzn2wczN6sCakcL7bmsUKGZbi7XTTXkpnV05SKskNsQ
zB9RjP5lGlNkT3uipP/9P+VFRkrEikICGunMnztTY17hccLpxTUq3mwqn3cc7fId
560nHmDjYzhL4Nift3v5UPscM8rZMeqQ8u4JIsRbiFjL+6TczEJCiXAVf4bpQNeL
DSO3FNg9Si6hO6jcmrnepE9d97NuhYBPtnPPaDYAQzVF30PA20cJYGr0QYmS+S1c
Pz7bfygCd0EcLJQFMsejSWO9UfHwWu/VhorIp6kSnfWiScbyMpdZebcoAzs5OTG8
vMEAakSdlJJUNlNAsMlkeBCBFp+67525IJ6QLtmzPf20SA+qAf1Z5h4aR0NHrjjp
2Xx7doTCiWaYindcP1qge/bPxegOFy6ORGzE2LL5KC/m3HrArKZmeMtEYA/+c9W0
Kz1podK4iLLmBZIjVBvEccxMJBXgpjdiWvlAzYlEVG4im+C9AAmuj4e7o1tfnsDK
GJG1lW+FPM19uzeCvW/ibVOmL4Zhi7FqT57ULiC6xUaq+XhytwPh1HU/yGBMraYk
vlQ4hdVmofVamfaT9jERuFLMsc0DWhGrSIQH/0LlYYkPwsq8AJsoghchVu6cFgfU
o3aof2qBbUPBmgDnCNcjfs/vOJdK3dtLbMNzOCunWFHg06j7ouYWb4bKin6+TZxJ
dU94+hR8raEEazpeOoH+UCjPMwAYWtx4OLK9sJmVPoceifGH5mN448Ft+Lu4Gfhr
ZhHXS6RPKA9HE3ANDMwmt7Uug4X/uw5ISElyf739GKgRWrvDpkZGYW3tOzgngNDA
MYgbcAltK0PBI3lNwJ7rGZt06DfgPF5zuWtAiHsBlItOC/YD7rDAhhJ/XGyImKwm
Zk48ZWPpfNG7k6SH5CrL10xqvNG6DPeXE9Emmwr7zgrxAFFY6BQpwhtV2ZO0He/D
mN9iL2Jf3NeAbyFyQY5jA8oPrzJYwlAV6pkCrzolLX+wMGSt2Vb7t3wZn8owO7zX
pHNNKLkcqOXeTDh+JOL3F7C+VEuZGaCmhja2ymsvfu+6iZ6WGo2lL91M3bbGhJMB
Y27l1dWQEfgRKE8+asAXLtvGUNOFozej7M7uPlrisQ2R0YumYp0b8P+qY8jD8qf+
LTfzM/S2cOrtDbXDHVIs13hAjUsKFrgONpTlNuLDGwAUjmrP4wy2Q0NGUJwgYj9T
zS6Y745yP+77jU4yJrEkCjmSu7TYtQCxteq7R76CY6PXsSTDygEnemKlTM7uY93S
owtblv33FOFCgvnv9jpCM/wT7mmFvFn4gGWLptUMg5Vxt2PvNEmOKtofsd3F4szh
GyDux3v43kGzN4xdwVVhG9EaNuhw7hCRldeethKbIK9oW69zL5DSGSGmXHWKo6eh
1jqazYskjs1Bv9FCBA09/oECmMc7gMeVAOWkkqGxEBfmIY2QAVZUp2BUmHC8Rgmy
O1eCr/l9Tvaq2OrLaKSS1X2Pba0JpO06+ClnV98xZ/f4Tltdgr3VSOmpz+d90lif
CfCzfsh05+dx81QugR9z1QUUMbvTrftDrbvZEiYZWU1z2zrWeKh+N1Fe3YCzvPt5
7pkhcrY0rp5NVHPCrDWudKDh+dU6o9vokbGZlEubhPvl1qBUAvJiHIcA72A1oAzu
CiCX4mOQYeKhUdbELEGZs2tA7Vh20WL4XUp9lIK7xwDBymwwKqJiqIBcxjF5WZbR
3gT3rsXvlM0aAbP8kiLxkg0wqG5dX4yLamwKMsNrzUr6JBxUXIot591Tr9Y+OHjD
Q8R9q3gyNv4vqGCUzgHf5JKFFrA60U1yWo7jIZ0tJG9wEjvVY/1wjRkUFYoUKFwl
hHoQmiPUgTK6LYvF58NGxObyo3cHpmW7zXstNAuK9vEyNj/11PridWvDDFDRQIyK
T8avdorJDpPJqfaKbj4KiVFASW8glVh9eRuu2qs4UlXHnP/VAKvQ0vgJxXR39Uyu
38SPTub4IsD24deBdw5lo2u0Xm39TELSMtSWKGH7cFO6ZB8MZx1JM+pR9A/JNzNz
iiujU6HfOf5jZwecuxihvz43u2p7CRgk+eq2dRiAe7mN9OUq9TG4MGb7YvBtVla4
4hPSNvYQ63GJzSSaiMp7aW8IhyQQMV3HYVpnUGIVgYMePk3E6g865XabK/iu6tGD
V62MgTMitem7QrYrsPp/uhYA/XkHWtMgbtXLuGKzAMaYPF2s9cCQR3VIgznRs1Kd
tndrzLPKkBKg1hH9KVyxtE3IM0/G/sX4RktPHm1sXjXxcfTAdL9KXvthdBgTgScC
N8oXH6YtYC/XyjGP7Hoj0TzMqJvtD6EV4kd3OpaNYT3IalaSCYqRSNNCpCgrDbFU
dSy7+eiQ1oIBSm2Nbd5TQO5g6ALgW3fbfIa3vluKspVX1hdNSB12eaJ8g0HZC5n4
uVdTDR+GOboRbb5us2IReeL05Rg6gMiyLDMq1DtHhQeLsNd4XtRhGoGkd7kFtwEk
x3+1l5mG5CYuN1o29ukiHjkYEiQm4CH2gJDqoXcUBenYMSTufeYMDI5Sk0CTxFer
NX6GhM9xjoE+mvUgvCdHrGqZPz80vCCqcum8O62Sdkxrxygvy8OfikeZgn+flZCr
s3Lvs5BpWP1FL5TvYEDiHhhebKNKQrsPRR+GFojvsPE/O/KJWkrOkczlsHChwl7P
ASvOERtRoWzyU0kSXVUPVW+zgdTlpRuwDL6h1sY9rYu1fdU8DMhSx2mrKRxIFAyR
vjSVuZYhg/m0kqCC2QYUsgePCy9G+nYGhVhloErqi5Z4E5cKazdAi96+EwbA/L7m
vPd+cSFZ0Q/oAHjIZWYYEamf/G06i9dEaKfuBC7LbthjzPZn9A1viYj8qIIMzK2J
2595QfsyxXigrKfSRsE+2TOyVG6Q340l1qjAvp4XjAVYRribH0unEdqfwvvAO3R0
RjUGePBoAfO1LGGaIqph9VmVi9ltnSQs9ofJr2TR7scTUlXGKYb4ETYhBdYpuzWA
1oUWD38LI/tulPjMEpHN0Ze72uPzBvPHxxzBxja8Zx/7QBk0DnrhGVxKQNhOV9Ro
wmSVETuQZ+BT8yx5SjmKQ2M7jfejrv+DTNKpzo548s+NJGAl/2deXZYVjl1pYKfl
NgqeWH+8Qg8yJmy9DptHwYITDbKW30fdetRRGHbajvkb0+Fcs4H3MOiOvpiSyiXa
T6GEqFgKQz6LJWYstXqMCJPL1loth33wlImNBC7tCi1GsVuRxrQqrxF8MQZK65s2
SsGL09VTL9WgTXt/G0EmV3GYdxtxjvSQl8kod49vtcV+8L9vVFpu2w6ALUR56uay
4HvOR0DjkDxP4FNgQmHLjHQXl7xX+M7OiyhbSfiBoU3sJZn4qQbnnwzbxBm2/q/T
CjzgxVkTsJIcFK2Wq2Kd2AA1qNystvoW3vktUa1Sa3pO/r7l/BZV9/FM5R1VWKX+
dkLiDQvQ+xefOSy4PEnymCtGRrazb9jjCVHbND9KB+DRDgsMA+EvQz8VCeYPOpNU
MPewgGnY0qT8VVc3C2Y0F8tdFPcQ7ONa6ihj2Xn3mj6FBAJOyHTi0iPisODjjP2e
bGZ1ZScFzlql7dYoEMkTtiIF7CLJAm4CszynxlcPwKZ/FrN1VlnBw/iUW3vce7M/
84NGTUnOK+K2VC4oyQEfknxVrYbBKk3gKQB+DqFCTw8qZ0w4vJP776bKp1ebmRav
Md+QwdXV5ysRfVZmgNsV53P4NomF/olXUh5itJgDW3UUUkAC6G5A4o+7PsKiBPSU
b+7jI0SqA1yJhdPVJQyChN74bmIBFdpc3LJUUrX9yyomydYAPjvRrMVDbNM7/hES
Oh5c+kNDF2a8KNa6IqziORmFkY8inqqqbUuyntCgyjDzmYtOhWr3D9nZbAeH+p7J
ZpC1sSrP2QqeLwbtVOhNgVycaQEtBgmeTIkLM/+8JB0flpedgS6LPNDgODrJivkI
WqvXpDAsrXOA7zYZk56h9sOUwuuO99bEAsBv5RjCfWsbkGgcN6FU3xvSbtpIR2Hg
TPvZG318uZ5oW80JJnvT0zCdW08jAw6iFYaHje2MhziYPP3VLseULHcuqiCVL/C6
PYoT167FsSXrVwMZpGyPxIAz5TDUCCxTJmk1zbrf7Tfc8viTkNNzPSyA9bWK/FRS
+Zx74Xzmbg6TwUVUpYEcPwO2yqA1YsVPuz099HUmtI0h0fr9TEvwLizeY/j2aAO2
fW4YufVf7fRvvFiV/62PQPFMFofKOt42JjXe5pxiqhiwzgzEqHc95Ow+B5w9n64B
vftNBc22LUHZeiKDlYfyqWw66A6n9rO5suf53x+htznb4NCtNwlKgaJ2n77waTfU
z/ByuFgPpRggAnlZUbe9EwXa6atFvlPaHLV8FQzjpjE/eCviBV8ikiGTM7cK0jt2
B/mY5BoG6vKOr+7szKpfWAvkhDn4OvlkJ/gMyIwvi9AUpE2FFcHP08yCMw/XvisR
4XeTRJ4peyVGKfyy0+D2C442bQ8OjJVRCi0E3/85y/7ZoKKGtCKwYsmQGd3J52+n
6GG90zP5x1byK0qEvb6hpKDH3WXTy81ZQez1j21qKRI0npMSgzdSRDxvvrpUPeJI
t5JK1lw/O3VjymPlOHi5JZAPNpRv8iX8uUAPqOx3AMxiVBJ6oGRWBV4u1viekdo3
qe2TWjeS44ZBAl6bDOS2UfLOd2Uc723roG0BZJVygcgxxnEoiXjiKsYTWIosXto1
Yynx4JhzTkLSc5kHX11CmbhMUlmqH945ew5QJ/Zn3MVk385whOYcrJFaKUFJupf4
Gy+1Qh+Xj4/96D2PpnIk74s/XwCSA21uVFN9ha6liUrKO64XYZmZ+Y3bjZlh5qos
0BHrBdhGiMkMzbS4aBJBhh1KRTrLjK1wwB+Txvm7ypJd85aFzCKQlODusxRV19Px
ZN8mCZ/xjyTA9yGmp1jhIoayP+t25skKHvHAI94bs7IaEhmsbxzkKtbNojjq9/HK
tzLlPwkVP+loXOdFFNG4wdmIrCaalYXUM5bMzcJS2+lLdZisXcGe8yjNxu8ctIN0
DyXiIo6xN1s2ESPSJs0730UjqtSZErmHyhVeNyn2ZZp/JG+DoL1AyaIeC2iKpjlS
0hv7cXYdU8Icws4gGfEisTPFjs6/KuDZ+FP7or5ii6jRLn0jPuJtvNUQrNtAesbs
IMKIlOAja6l/MMJ7FJ/bnzVRdwmOGUI879b9d5Htp1TMizjLah2KdEAsikOEZlPu
BgmljaCYx7nrMaxnKUk96tCW8KNbHC1YCGbCJ7m3BirVYzPOTtvyWN78RqnPVx2g
rq6noI+7gp30Meb3YvoLJEf0aoG8aWa7Acb1BCw/U64SrdVDFMUbIN7XsffNLOqK
FuFVcnLj8rzfnDRz9T0CmXD8egQ6N8pejGJU21o8nJ1XIejEa1YeClJpLa6ZuqFb
n/7qIaB9SzKuoy8O4axRganZI8geH2WDnbkkAqOxXNGOuLcP0nhk9KgvBCSpt4oj
e8Cwe2cnpQV4/5JdcuPjakBHRqui0v9mt/7YiqLFKrQQAdXXCAOAM66cJEGtUtU+
+GJcmX2dFyfUUmMw3KeyLZPuEKKE54IAN/5VVlkdyNwkCl4kx9SuRwnCEvnrbt4c
2KkEyezg+/T2xUm0+/f965ecIWW7r7I5IkEGv37JkFf6McS6RECwa+evKyJdBWiF
cDkGmoLSsDxtnoK446dw6cjIzjbPGjTvA/CMCiSqu/0plL54aZS4utTMrLQXgvq4
ZQ2U0crZGSXuUYc489/pdxmCF5aJBcMtf5Gf3/ku2vbU4R2WO4LzQllShbl8QPzf
e8vq2r+N2oDsRH0Asdaxhfyq+qyH1ZOvrYxaJJ8sfhI/WWmb2peL+hJqAo7oMoYN
ElEiSP7kCp5n3xSosaftJ8wZZeE0H348Bc4VrcyZTyDF+JRHV8ztcfvX8iUo8OTY
YAUYq7UKxJWoL+NNjwm899Ho+UtiD8rOZhIT3PA1QQWtTNjC5Ah+sda4NOR5loGw
vROqfLZDjzeC+bLbDEBFfOkY+W/fQHmFxZ7yy+LS7UMgGDQG/voG87NKjz0OJrqJ
WNwwYUTdsHTbpfPir9uoWLh6FVufbQONknCydsVPlfCs9LFX3Xr4i4lLMP9EWhN4
IIjd2XTuWrdNQu19PFyVBvT5i4t3S2MBvZw2OWaRQOzs5YoDW17FH5AXzLUWZwvw
gkpzSDIzVa7Du+G+aeVi/78mG0l2dZ0+po0V0slQAz0PvSyhp/SMf/RY90ksskcb
mCnRwazUMFUwmYUhe7cflHI+ahUL1WEeb4SY100HeZupJUHSJGckth0k4nOSRv4W
bfe8vHWuJV0ccJ6C0RM+WGWYD7SVMM4N2FRYYfMvHOh3lJgxUu5jpaJxZxl9psbG
FZ7wVbFXeK7pBjSccia8JaYju7str0iju9sXTbY5t6etIxPgqqBIYDpKW75hTBnd
PMV0b3hlpysJ+dze5nb0pC7cyRL6LyHjskqLXIF07qervUZfZ2UZWyH4Hkgi6np5
bjxtkBdMOSXJI5P8kmEeCLvlnnkiJC15S7g4eOEr9URaCOP7aTu/hpkc897jHqy9
rrDiHpEazs2Qt5Ce2v1DL6mEdZKa3fDkU3yDMgNqDMci1oXuDea9SirVwbMGGhyC
LlIycOAxpNuurlzPRFHNNfRYEDuhKMghLABN0TpiuuGc6GVBK0J7hXvYoMJVmkvC
VRFpa643hbMogGnlWwd2MiQjAoAcdnEvicvThEHS3gWa9B4bQmX0fe6Aez1Q9b22
x2cddO1hLUrEDxXedaBlatb48GVPBiLG16Ztb92TIRsbTpeftws65a4/mmJQEbmF
OwX1uqe3i162m0zxoy7+fmmfXw5TscH/czd9gh9Cezm8nPvQUyv4WLbyIFGcaE7I
bAmnnXXjqGHce9FRz341RwCfikja2d6Mg3+rEfqjAcP6C+eFvGAgburfaLYIsOcu
jG8L2M1/BJxoM5Wd6go6xOjHMAbgK2JfAEfbYhK78apGMon1ZQb+HbLBtdbTy5SZ
vLwf34EZCQ1rNXPtcZEjb/PhDMz6vMTDYiJFtdCE02XNMfZAmHirLrajcQlLXPhB
+LyHezIt32ukSy8JMdgqI7u4jRxE31/Gb5GAJ3t9to7/a7QmlNypVQQbm/Znh7uF
tTiQalTwivBnvZXBxnHQOP1Rp4xjKgt7tbwiAExDiaHs5VVNWAJh1GapBrZGAKBd
+sygL7jO8oRlVqbIVIEDtUD0xgfDTMdzCn6O7gav2ucm1MMiil7yYbS2VNtuUblk
QGV0QqjcCIUKI/KmqxElJQfK9Z2hwgRotW89t9mZkHQLqDLAZ2LiFggpZUTzovOI
hEf9qYSJZz5ZczTCAu+814GO/GInh+a8O0GKA8/DA6teDqbsJd7L2PIfrEJ/WuXE
hrT1aWuHIY54eTKGbTt7xgMbtVu4ovb48v60OPOAx/78Xnyr7gtbsOJ3stgHprc2
s5/C1FMv7IfFsuzppc6DpQZw1x+RXlICOzofF1EWXHlYad7EZAEieaPQvysMTIaA
gdJRFmP2pSY6cnnVOr2Snpa/ZIRMluLig4oCcxg0md7IbV4mDie+UbwEcJck85d6
wEOQ8xeXrDkq91IC1Li9qjsxXCl01dBjpjt5N4rMmoRA1qmKZxFh1yYJPYE6vSfs
ralmVDeMh9tIsik+HsSJErVZcON3lECcbWv3fKGj7DFAgvDJY3vyK8KtF6iOphBs
zNxVwgYkoQVL9thi7Dp1WYqzluyq80SJDC+2ClkYYBoJ+iTqip1gYMqFxwLs9FvY
9e6bQ/TbXGmDkSfVlPRAcfIo4R/QvuakHV/G+JK1xxNXrcp1ZPFK9clDTX2knMf3
x3WS8ThSlieW+AZsKwVUfN34a+SinXVH6Z7PSv4R9a7vlE1q8w8YGuPrKxT4T04b
ArNNzItzK292SWs+NshLU5nHRjNKKDsQ31jEGFnd81lJMAa3hlZ8q9Fkh4Wfg/s8
JNLhYI/QTOBY0EyPb0DHtCbakbn7p/wkyMvrdK6KvXnrRUbD+Kaqb8NMTQjdMrIL
U3lc824e/0ZMS6UJTjiS3afNj05M3hTz23R2RI6qlzTX4osMUEKJI46J4/bCRkXY
HtfPsVnsfavPqz2dMAf9BZlJRPtKNvdrcuVIQ9NVq5f8Fsj7VYFdh1dfuVPukOe6
iTp6Lmdfg3xVBJbqV2nIwatfFkR1CKTupIS6nOiA9X/h3pek7vgapFXL0n9LlIEo
W98EKEVkoKpZ6IOSTlfUYAF1cuJ3fLPA3946YCYC98Qcfp61fISf0djdBCC/ikQz
w8GqChT1dovfnN9fYSDyURVur4Wmtfj5LEaGciZDW2BoE/bPK2VDbS8+17H2BShE
wW8cUxK8NEAP2tUDjRVD2j+An9Y0JpxXeVZbjGL3xc+HavuQOwjtYHkniDbKuev7
+OifSaVDbZQvf+AXmObOx7/Y24dHdD7j1WSr2wDktBUXcCck8ZK4l7ha/IMW4uO2
9DdDuHbnO7/CgTnQhBuLUaGEHRI6kpAHrNbWYGDgkjjloe3EO75EO2GkxrH8c4Qk
nzIQ3/qQ/o5qFWpUaMALHQaXDLv/aqusy6JhcLvvvv29BPsYMm29f/J9p+9FLFdM
nzvGIEJEB92gH37d9Zgb2uDToKt3wEHTfm87ytQNhyKTRZj2Um0VyPoLt2Fnt3z4
MeOr+kXXPy11IIdvGLPMOc65qKl7ZNe0SL9oh1wSe4jnpmoziHjUk65Q6z317ltI
J6CxUFo/PBjehISy0cr+eQA4ZLi+RZ4COHlsDMXsRSotIoKgxbVnNy2HBmlYdrKV
3V+HgOn/mgnaO3mVPdsPQsd4XDIeO8cGOfJFZEr+ZigeaQUayJMbg/Chbo6cfgK4
5AwdDEC1tBK8pQSqp/bO21bSaY6wXTgTSIEhuNBWzwBVyn+FYuUy3wmKf9or/X1d
Beh4BwtciGt7ke4B+gzg0/1tYN4sf0XU0r5dEzxrL+wXgF39Kw+JzcnzyHgFlrl/
EAr0Le2sU2ltTzjOVs3tP9N04LaP7bWk5d9dmgdOn34Mem1nHXehy+piQz48qEKf
v3b0kyZ9gbqxmckgCmxSpsnK5T9mb6RjWb6gqOH/mEtPk+NLJp1cMvwyZVALjJbE
yXzO4Td9EH2/yzMNnQYiYv+DxKDRsJ1NaUGISBxCP7oMdsfY7HsIvI0jAWT4Xsda
rcfknY9F8xUAyZr4G1Qh1T6TB/nvdGRQsyzRxbirQ/vL0rAcfroazZVjlivuSzUz
AwDUs1G6a0n2IHomAxDNT0C14UOUG2u/wvFRCrpDXRxVcNJxomqgBFSo/9PDAoOm
GuS0miIpUnNL5hYBWvWTzRGRdvCC18eBat9aQ0jK3EPlYWNbN9HQXzxA0c7DVKWK
ANxnCFL8oUO0WksWe4l5A89niBCm3zivHZvNz2JsxInTQhJbvGq7GpKeW8OOZmej
XWcJ9epZMmDVW2d9xIWB59XuKBxwahJCp9pFuLFFzRIrPPH7VSjMiBgxM6H57Scc
Dn9CJW4zHqPrAQOi5bqpoRZLnKVBZQ0jwYTMegjVQCgA3ZUmMoEFN39sTCSwh67c
gFzKs21Vxe1pBeh2mZX2TmGWpC5WYFyHPkyjYmnpaP/qOQlBkEi6jrliniZh0qmb
0B7x2pd5iL7MjURxEXayYB+rU0/hDPjMsUBttuYB/bI2XnHce/S2Ax/0bdyWf431
TsaKbel0zfNX6pwnl3SgPl3PGoG/+RXxFiXx6jSwTvhJhKanUCPz1oFFQECYq6Lb
3Sfd45SBn3fMABw+ppFE+wV7kSb0lcQ5Bm/uS6sOFAk6TwagrggwJb3zBYe5PPn7
+ZXSG7CPkFqxg3mp4tpJYaIWYT4l/I2tbWfvhqF0A8R1lZqK5j9DmWsRfMSUfw5f
kULjxr6x7kMjkj6DMsK0MwD/8lW630ho0A7oJ9/PuW5aDif3zMGFWIaA4ghYbqsL
4rVvO+UGZRcyEeEdjYya+LBj8gd4tHQOrwZd6xmsruptElo5/NuFmoP1Veyowdsu
nDfQ2jitAecsv6jQF4dWt63BGG5yDpI7sND3vraxtEWeBNc/kqzLtsK8fPrERoAh
2SllzS97SeY4uYxpv1YH52CwQgAQX1jlE2nmQQhkOmL64zd5I7Cm/qBng3ntzmey
kgSomFFnqLua/lRvnsgUXfiOfVBP+2R/iGivMd5JR70iYW2840zs9PxKZDdKqRxJ
V983h85jYjCZN68o6rvFcuANYDpiFD978obuzrMAvMX2N+6vAoqMAOjyRZbswOGf
iq1JrmEzcQoDSdiKlioEhUmMy8iGKAphHjNz76y5phijQNb8M8m8dzL5IroUPDDc
6jfEsKkd988PrUEIK5wFC1yzHYj070ebSpg97RjBV8h+wf/Gzu+CYuQ5u4QpX1K6
pApxYtnY5OTaoRa6XEBNC60OFYbj9OWiEYq+N0reS5YH8d/fSfUnVaKu52bNb2ry
Z7XV67Q/zN7m7boaaM/+h85elFnJpSy3NiEyQQL3lxRIP/+wCq26c1O24mxA3VyF
5xHvFHZXj5a1s+Q6zPSxyN0hFOeHWzHoJRQOeclkxa1cH361H2HHtF9I8/t5gleS
4tVLmUbskUanwgsCMfCEmCjZYnNmaaknuugHJN0ZOLDZIi2MMb4PWGB6iZcJwDKV
nn/8QbXPuGWmUkBRW5vyEwL2dFtKhs4QsVzB1pwjIJx2HYN1GMmwMeClH5feS2Z1
Vb4rBZXKbMihfvYyDdWDrh0Lw5QyRSsn0VF4lUKnc8Au308TGfQ8C8dyMBeN/UeF
jhG/nmvQ03z/1LMKjcK3TygJtXgZkxN/RUyG7StyPgfMAvl8xAlyLVhNnf1lyW2l
uFsEkuvS6MsrX2q1YRrdJqz42PhNte+EY/cct5EhotmWoKMzewajtjItuiNiZ+/6
9pRBrW7XlYdmMHEgFzCO6onRgI8EDB23VzjrXVUl0DGyaSbkrMEjYzztkQNoTFjb
6z+15MJ044WIbwwRSFL4gG1tj0J2sMKXFYmsRBVTdg6L7fiK8twuJ17m9SZ4rZpX
fGwGLli0cTa4md+7muA/Cun18F1YW42Pg+Hobb8sbZQqNa1g5r/L28bAHMgmpfPl
3nYLrlWgPpN9VmG00ZZ8/GcFLm6y/elzwVZ1nTU8u81sJbEkslhzyU8aFuvQsIh5
0eNUmjG7VkqM3PMhp9/HQ0Gd1wvCT99S4ZIdMHr1wOD4o6j8ftVvaozBdApHnBU4
G94hhupnAVF/cOiKlDPPYK45DgTeK7fhJUmElGm8KGsWlxh4VDRIM4H/PvrxDh3/
7SVc9AR/BDPoWTNS+lTj9RYaaxTcT1vQPgZiFi73ujyP1iE6c14GQD7fw4UPzDOY
xvTFshMq3m8nuFxosRBY3Ez4pIZsi90++5kBc/lxfVSDEM9SGDOhI330S9XWvUri
eCXI5f0wPR8odYfqsfs1yAnDr0utjP8MH11IuRMpa8TMIaXjttadONe12whLwht7
lRN/pbq9JyNQ9pNWtLYiz742FIUzi8f6RJSv+5CLUFr4lGVwKoIWXMu962segJL/
kboxDYAyRLamzxIt2o9fQ3ZW9VSgtX+liVXz+IEti+ZDwXsXx06mjJYqu0bkunLq
B+AAdKbaJCvAhmSYJ5si0lszvv9EgVEnfQLGJ6w1KETPLiS7C77LOHTbY84N9ejU
I6VYS8PoGnACVRjcgIwFCj0J+REcmmT3Md+Hg0/zSWeCW4TTvw4da68unr1UjFms
O9yHcs9yu+hppu4OiaoBqSbetZyPHpBHil1XLyIZL/eSQ45VarX37Huz7ASe+8h5
6ffYmMbMc1faCDXgp/0sp/4k6M6jpQTWI3XfXAXStdiJW/Q+fcY8ZyeW8nQ1DKZM
r8wnSedQN1j5Vk996+yEQe50w7x2DDz8ay2gP4SNsW0Q2gQ0lzbNYSIH/JqcSsId
PySG+b57N0p31yykmP/QmvDVjY3E5LWCojcWEx3MstP/dxQlwz1iIhMiuvYTXWa9
w5Hk/6SyktACiYrNTctUCPNvmrOaTO5kA0oVKA/T6Q3Rh8m6ChD7BuxzEjo56Ibl
9y09l1Uw800fbzQMxjlZhnJG2v4j75weOxeQpMJ23IkP+/apfbt2v9fCp7Xv2Bkr
xkhAODRnM3sheQG6gP3CllxKhx3qZTM7sBuwUXaNNQ6YNBbVDHUIJEZ99Q/upgBQ
56aQz5wrm4tWGnuPK6qZqUdB4uXcamhCZwMQKMmW8H022aGbMAYMdL4N+yJXqATo
ZNvgx/Qa7UsCTuS5JHjkaN/3ZZ4sxP5x+YD73SbrRih/h1wUYVPo3uA3PZC1Jw6Z
Ewh74/FUdrmCgmHbPRCH0gd1oPYB8ctOT49gw56JH1TBtBwhLAE5dw1NmdbOxAzs
ZTqEu2oSUkn+DBR9xsWA4MlJFNteEgagMww6PJhch0FXzhMHbmXlp7qz62/fprPz
qz7aDRGopJZ2zSQKaW5K2963YLxB3JztMG+mlYZq0v2atGbvKu1lVhyouVE4E0j9
QXy4mUqkiFLwqR4PcDGUEe6tccpkAP/nHZO8ZBaAFeETkxxvw+mdQWBOb8oHY3K9
sQaN4PiZRSpV72VZFOTCzGnGybJpawXn4zSObCGTQVs/YWU79b8gIOeh2tl9NWie
Eb/d4F7OENpNXVyLQxkBwhI+DalvcTKIt9PiXkHsM8IuCRb05xEWX+Q4Mmd0uhTQ
cIvI/VvonDl2uH16WRIMaTb6hhe0FRwoeihlvxkg/ezL400FibJndxe2mhP2xl3o
AFELQSc6pDujk8kzAJuHZVNeWbTSSLCJnX0/JJYC79R3t/mpI6Twhy3JXk6rHjNw
6fazRIS3Y30wXr4R3HzuiJR3Ve8DBvaTAWub86bnEtqOtbLVFYPMqHoojkiXwaN6
ZXqq+fmVuov/NTXwAG1gZ732OetHh97bm8Wxv2nc4tNKIiOBgJr4g47i1+e2W2jA
fOGaeBVkQpWfZ6OUE6q6lmEyZ9ErV42GEd3+CQuvYpv5qtjdDwUUG4L1zrS4stgj
JJfxaFs38Kh1U/HMS/p1jvfJwHlSnPko4FXw8NwiRRGsUbyjqnS8R3bwt00Old3R
LROJ3JOJsT/GA2Fz9W4VuNu8yaQMOKQ3YjoZn6PpBXK7QGr/quR6WLS1CyJ+HIDI
fVLReCZ422pDGnCC93UEEBk4IR1q2kelXHqk4WJ9miNqh1rVRgvUb11HVSt9THiP
P8KJGgbxVi5hlk6vHPqKxgwQ6B6tXD1J2rqHAwEG5uUkE1KJwgfkHhv7hExMkwh9
hNBNB0RXresDitAlKzWbwptLtod5vp3Ro2LCvCFk2uiljiLiUCtu84eTmevecjvw
UeFe9kA4kCCmWUxpK32v4i8MjKjjQ3NMR+NF1alPTB+2zWtabKZK//jexZ0lDMi3
ZCW7G5TtF4MkKXM0qEMdbLKxbSd05zbnocoIi7cOOjR38YqI9QavowIv/1AuCyAf
DblBtm1nlGXFk9TfKKvsUZAgfdnR3ehulQ+KYKGZNnvXHXvP/WS7fZzVxRANig3A
ARdvFK4Nm4VqpG/o3bOZ6z6pthozlRDLA5HMz1MbIba1tApwBMrQOqII2diwse2E
wewOXHmAGU2RZQMwhJc4D3akz2v/MXJqvTS9fn1T2KiJXSGBBLYC28jGrePi8bPT
8Rkvv23JHXlflLkmQPl6nUN/a7hfWhF7+E1yzosRD/wkO2Bt6eQ1tBceZcjgS5Qc
omef2jfAINbwuUxZ5Cal0CewvNwKQe5eFtsbkPkFjGjgoVIdpIqWeq9NYn536G1b
zR0+0Tv5sGfDMChXEL/CmxQck05YY8xzKvlZ2wtE5wYzDHKlT6rRzDDrpKfhyb6H
Q4yNNKzi3TaQTV2XsRVOZJvKC4O1MYTjwCjmu4lCu8RC+zh0ajZxQxoPA1pL8BDZ
aIHpotnBNn7yzSZKlZD+ZqkQzcsozrG34S+eRs9rQymgUUkku5r7y4xpj7fva5+z
F/PtP8b6Y5eHWosa4sdxjKxKmm3WhiPtA0DYdG6WgxhSbzBwECPFS2dhjWKLrI4i
yPWqkgrC3Ciq1A0Im8kyOxyhr+/gB8HdXHGOlgfCHh6qrJO25srY1e+8TX8rkPvH
P5ffs2zh16wm7anOmuZitIWUOFFVICOP9sdUi9x9jxthLG0tVBuFIYsgsFUDbbKJ
uDlMSCI696JpV/gn60AqEE9FDaOLwa+MWSLUaJ57zT1HoP5Ah5rcUngB5RW5qtKa
jX2/rv1ymqcsBKHMaSgri1ynXnaQ8TTwDA9xvNO3bBDz914dpYC8IZAKGT7tKm2j
R4R8M3AbxxGqZeXYE31gaIkBUP4AYNt7oL1hPXRCuZAK9gHz7mQ+oDaXcxSucpMZ
0ky6uoN3iggEz4V3oEvRCA4OzbHhz+Atu6Kyvvustbxu02hcskb5jIF/56FScG3C
pCOfQIxRdh4oU2jyo9yS6mrMkmvJvcKgcqwdWOv0dtOoKxn/3KBMvCGiWwAFfpoT
E4iFf2/fB1494oOKiiBSmiMldKwhoGcSCpU7BcMZXHRtMIS4stNVb4ZEgV0roiiJ
bqeoKecysJQ7h8j3SyCOGXejAJ4fhrYIcHFZqWVPmhmKogywwqQY85MGtf5h4BAk
t7eITzv+qUaKtoMh7lJu5R+cHtzPrUJs1yV5KBxda5OBK3tsmN98VlCfTacx0ZLA
zPrdMyn/+pip64bIUNroPSADjVi4F2NDO5NwWHyMWOkh6vt+a79p/iIF6+5Cl2Pj
4swuyRDg4lkJvdN8YWWfkdpzUeBXfz+DGAaRPnNjQxVF5WU3JL3y5yzqsppPv//w
sWYzwJoXzyQp0fvdUzO5BRRLDqGx1O7SaK8UhRgn31/+kZyJy65TXb7pg7SJz/JX
m0wEeKotjWomIync6ZQctsbehde5KrkQ3SeextCsOFdovrh1f3pqkdOM/rZd4s0U
7diVXEYuJjZhAfc/p2nlFWyOj9LbORoD1MbHJVfFHsabUYnNXmk10wVH+2hlDWEh
V5bXm2tV1YSgy1B1VEGOYH0HI4EUGMJ91yS3peQW2EBlk/NICsf17R4P8HoMIazv
LoEQS3rkOAiDjZ0A5sSiIK8FNtiMqvCl9IyXkuZLNic6POjCtBoXMiu1+O1GYklo
tVQr4eqKuggXdnQwM3DKj5kHHiUdU+ivGe5m8yHWpLqCfIW+1HlqK7W2Ts4w/xeU
OXek7InkCnRg0aStwiopvB8nS4WNzAUi1Vqa6nlCqspHb6S0Hj44v+79DVvgjWHu
R1Xe2arqe699Yw18g3egjhhXE0emo02ipUvBetFFkT1G9bDvBV2ezZzOT6d/S73X
3tBZotZ3INyrqhGmLfjo8P6wgbEeBrK8xWaiSmKJO0Y55yi77p5dStBc6SdiSjww
vksc9+Z3KOKNSTaTww1mkdO9gwHncXkZmn30GqdtJHF2O9++25ZUcvcUbfWcueOJ
SGiItuEYPXm9pzpnIIiyD1yU7kmovJTlBHaAI3mlidohmL1/aZeobMWziyxNFg/u
0iD7BxY/G+S+zUOUE6Gxg/xFDWS92rHAIznnc7+sZxGBHZzdotVTBNR2kxf109Gp
AwdCV32VWk8Kb9wDRoriJaQJf4usPwoV1mC+apHsc6/0q001F4OhTK9q+cCnDV80
qIlNqwu0Vll3WA6C9yJ3XAIjoK0KtD8cqM3dBncdIW4zBhqC5yJOPPtTn9y0m0Fq
vH2OCGToRUaQDQPdZkkZ13S6T8USTagV6UYERaNJz5XmTU9A3vWYP53EASOUSpbD
BKyzKvoAs2QKubOgYC6Aet3MLg4woX2YhRWIrhYuzLUvlsPTwKnxMPSQelYpjQCB
k9ah/MiLoLadeFFXf0QhSKaNAhJr4AJ9apUZf+SToDAb/N7h33Ypqb6dmps1D1dx
BP5Csa/+vZL5gGbVxfWk8qJIfaylPeSZcqLL1OZRd9ldKcZ4/WZ1AzEolSgHN3En
Q6duF3l4oEy8a/svSs9SILP3dVVGGIdSAYo7dJ8FXZKZQCV4/e25aIogBPTKmS1t
O4DVDljf2LgxzjBHEHfLIUqRJcApvyGnqds/S8dYRBOdGxJsqZl9BXX9JC1+I0KO
1YECh0HCGrEBdJi3vB8YbddzQDEcnmgVZxCm5DJbsDYvmsxNbe7LBCr5rDYQuztI
ML+xKsgKglrZfqprgBMz+21lBBwTXnHuEY7W6q3lcWW79a7ZzLuwHaqs0auAgUL9
dx8ad8v6UcTX+gleSKGQZRFSbryKhrDrSPJk2z6P5SvG/NBbU+cvDR51Wf1UZBbQ
Bz4BGHbRO7yf0SrPS1zVmmEKcqosypqjz7wXLtuxeaYnAtFlLJab3B121Ndj2SEY
otxWbV8yMhGNDdC4At2nB4E08+aYYyYYyFMgZ2k8shm4OMF0yWdPXovwJh4sjUCT
HGxiHZOfBMpvgqkKtUIZGsQSZXlYsSSgCSNmBfASlZ5CbK4TIUmGR8klqSxkmz8S
1gPmBBsr6y/ydQGCQJ9pyteoVeO02a1heZg5AAjCSS/vvJzXnI+0Ys4/CXaDBd8k
haYADue2hLso+8ZgNQaUwb2Hr3VOgAU/XgLl7IEDiuYIE/lFjWCCfb4wlVUesS2o
bE9UVatXklKHDGCjxJRqAkuGGSPJpG5pppufClZjOlCBX5d94tEIOWGNVIbsjdi9
qq9W8AmLXT9QGJ6cp6DJJBebM4paVh3eiuKRaPw4HPhrnbbl72ne3mbGRG/VB24i
WjfEYPwUxuvtsfsnOn6i2gaVE+R/Padf5CtVJOWN1HPNfh8WKn3mc07lnvoSOyCV
G3A0Z8WoEP31ILEUyWNsfR+TIz+eINzPleTuO7kr+fI3ib8ortuPX7YmmRnMic/P
fTTLvC5iT1AkWfBarlDTvQPdSfMcgdjKiic3l3Jea551Tl/Ot9w93cse4xWpRNHE
vU6P2tIBXvE07sOgEpob8UK9Cuz+r2EJmgKXtQTtieS4+c5T752g+z6fmwEfsDex
rOz7THdxxI30999U4HCBbJiy1tPy8bYBwWtV3tk81Uz0PGFYCsfwGqnduOO6NMqX
UD6CwlkkqmMAjx2frcl3pOWEKLDzIs6Rlu4ZIII9Bz8vKKlJfZ0yU0WpyApQJrRY
MU6sdftbtX5LlWaVWOC2rMNs2Ln8ny/zlXjfxrXYTyDUGAT5NdKYBQHmz5oggtjr
ZvQUg3Gk1buOHDMk67dvAhHVo7ZguePKzNuZlGSW33bcLb50RYLwTrK39IEvabp1
/lbjI3/mXfh8oXkfpGQprTykJYwObxKn9M5z3VUqfymmhEnZnphLA9i9elZCVHhe
X6Bb9TiCv9TAx1v7xy0mEeOfTqnE+LaP5y5toMz+dP03KbDXxb4LKSKqVIWJLMVQ
Ds/7NqmzaNZQe3LqqBDO3RXQxZsq80kCOK90ZwHko177PAAcUPZdeSw7LCRnsi4A
B/UUFJ4ZZzJBrPNk1vIoSSWlZZIjg2omdYtCRz5bLZnkQPNHZx02hKT7H6bqQDYQ
Mi+06jUcuv/ivXH6y++LGTBfHxA+ND6fRjVz9OjG0VKwl9sIhyGX5e2jQlJriMyh
+nb2XduBM4NAKyeZt0l92XGge51WhdNh33AoWftcwrTJCZ/ocmxlqQykLYYu1gN9
/MFIZPnBb4yjfns25P+tfjxjNAmajdVZRDc1pQXWzCteTQzVbZ6rFIsBD1R9Q3iA
RSV8FX/1o4EFq/akVlnR1J+Ljvg3v5tCf1CDkhj2UExdLYW+dBWgjBOlFvR4IV7K
hYm5o1ujCb8IGI/nxaEp3kFLcuSENVFTvLmcZG9HB3zHKRumaxhj5Nku4ka3oGEF
IWFRzxeoktMMegwHvd++6lh5swE/hHVOfpGBRH7vpTmf7ugEtqz8FxKgxmuNSGE8
Yf7i+e39bJPS51HohJ7eKa4MA1X21mkdlARd1dO6wWloF6K4W927z9SQK6q+Ywwd
V+13F/wiZA4eDSfIkjAPle7B8CqxPdcr0hy6haYmjoT3YJeA7yVSfC4wcOWmMWTo
776jyjJridp0ZgD3VmPaPID/BsHcBJuTLHeDChhvBjg6+S/hwGSWMHaIXO/uWxYD
1XZmZufB9cvr+DxLj+ykOH8gvPp/CtqbT1BvOsPJplDHAyWj2LSbE7oN5IG+UBf6
M6t5Ob4vDlybUGr/EfHJeNkSdhoLNJZAJ4bU5RPddbDc7WWdiTyhhMCIa25As7Am
QrhnU5rt4mMQ8WwqIvPWBQpe+bZTy4NagXmaRNPikL2kO/hDwNeQ9N1n7yRxY0LX
6PftQU1ylIPbDv5Fluk0KzFl0axDqZO4N3mLDD4sLM3i61UtMyGQxaZY95Z3Dbb8
H5xWZgtJmpSZM0Uwu7THCwxBR55IuE8IvfQ71XypiVWJBFfjFEDayCPEUpnyWXwK
b24Sfa+d+mFMMxzfmtRmUuYVXDKW2f4alyva0oKrrbwnZ4PiDTdtmJd21Bh69x6p
+lwjcqmp0Psi9oJ2XhSwiOzb65aUHoi6Xz68REuQwrCWhg8AF9a+y0XNGNUVuh9M
fqZw0KlS3JeMPm6C7lBODOpZKcYBguCktQOjUUeSsxrU/mHzz3l0jWsZEOWE8kZ+
cDPgfVNLjAt5sr4deSdKjQMaZ3E9VbODZNcxhuSXUz8sOR76YBbENaZE29k+024I
JYMUhjI4PtuFfA78KVjAiYKz8S5kigaDrOUHkqpz+Z+4UYCxvrhkb5EpYZQDsmpd
VyIFhHRvQJzlXsDgF9QUKkRlhNKTiCDqqe96QaXEuv5GpMJ3I0dbzmezkwFZkb/C
k3zYgxCFyvJ2zDMTj1HGnfSCU1m4exOiQU9WJuNdPasQKuIu+ezq57+TQh9edSvR
wi1Kip09/bRmP8jVRuUEZqApWToa4Tsa5/t4224pc/VDdYAcJ4fDrbrNB5B48v2T
zyTpEgPSjhcoGbH0upj6VQdwZB/7wx/oAyIHyKQhiJCDHkZmo8zNXHKrbYVjprLV
c2gdPWjzYqVUdCDKUNIYB85JP/msUvckHJV8/Uky1PDZL6QZFe5j+NzCseblQxmG
BmYL2F+JWphnrlu0CesUrslC9jCmYu1UOBiR5VmS4Ilo11A68MX1tOdCUYhU18aX
cm7r8BmLapvIxTEtSlemDdbVUx+5d6OO/FhsUyxOQm73yApFug9TvSc7qMrr9TWB
QgGrnLWJT7IGQDOjur0b+aKY+fCEIyBS/YV57RJETNxx1YmDgp+2eNg6T2ZC9xUm
RDVntm1+t1vpgZbQlNgq/MqahlGP8GcJnwKFl6dwYM+bwHfEV/3XRCv9rve15kgR
U87UX8CTvjpz2FpYiwd2ogFZY8eq91vVyz854y5UT5yUUE6cSoU8xxK1RRJ8g801
C1huYhKoOz9S+V3G4pwforSWP8UXTwdqcouspk2J3heeBXCS7dVGIUplSm6exv7w
JrfdH5ThQn+bxLBl+kxg10pzomWqZhqTJVzTrBySPPeDhr+7Qnh7G3chNb6H+ldt
4qAYlYRX4rPPpXZ3ycmr7SosU72E49264qp3o6SE29wS25qy3QN2sjGIcF9eb2R/
8Usdm+xtEZrOuIe/oqiBhWdy/X56Ikh7e9e4u85kzi8WBy2Z1Ml80Rkep7xx36E7
YOGHEnJm93ab+mBCiZgjb3W9ujzLR0ES2HQlSc0psA07iCczwAlJIDg14kU7NSgS
ZQF72jes4oIeBzuxAr6Lx2Ttrcm1V6kcpPJ6e9DyFF/503efBDUzNAcUv56JcDnY
ecbe8nKWTBB7jXVkUEVXGYzwbWBT9x6ICh8ZjEX9eyPkvvQGUZhIiAb+uJCjZBBx
1sZ2Kc/kVxNPsZ5eZXQ7tEXGB1E+0synS7MED59Y0l25gdCVTf4OfLYcCzGiGUc5
pzqv/SCQLIkkDphjXhsGOtierPLBC6bsKuYYDI8+Dr3uUEAWO9U0EIX0nQym7PdV
a4p7zo5NgdYAZknVQms1r4QGgGLjwpYKb9QlpjD1bsO4oGTn/73src0unri9wQVF
iJ0tLYqAxkeU038kI0v9hue68/TSHy00Yn0CjfJi83ywfo8MTqQBqfCjmEcwANRL
7vJ/Zdz1jGFvjYnILgMlN2KX5U4xHuOLbE5vm/jwRDISqraQ9ZBz/+ALY74jn7FZ
B1Nv9oS6auNVWgiNEH/Ma/ZFTLn0/NMb0e9ET2XsO9IANEl5MoTY2ISCpdg55vt7
PyFbAce65wN3y46slAMLnAKteMUxUduQU0KvnddeLA4aWStQoP9QC5qpxH09nTzv
VEG/ugw7B7nFrlfK09LXh6IpBFfVjM9VbecQbSAFXpDqS/RF88120CVvIBWdo/Ob
Rd8Ydf1XJGdHxstkYZvq7H2Spu5/FqAj+025I52UxUHiTryAZTAjH+cRpQSKVbik
VF2/QLSULzYwjCkyMfpRCmJGn8NNVTCIjI9fiU/3s6VWcNoUYXqWYjbRaIhwM2XR
O/QzeC0TLb6j0ZqHJsMi000poIGZg1MZYC7mCJIWZWwMXWR94GkrIUZ2Ag///EWJ
g3FgTubByRe+CZvTc9Ip3crw5Ginr7y9uCREgwXWZYzRkbRUxpP2K59wfNsU1hP6
UaXqwW/O55x0rvtMX7HbdgAREhoq6E8xwKCU9A2fbiV9Ug4UTIGVWbO6PCwXCv/J
YjfGx79q3MtRB9R84QjYsMRLKbeTalEZh025fyNvUEc9Duh5ar4rHzd/Qn8eOskA
Xc6sQc17xobnz0ZykUE/XrX/1RO7ADFd4gkgKp4lqYmWr1Z8t7U1+9ZYOPoT7Ler
Z1MitlIJGfVZaImVdkVJToHFjpkdXyHcXMAuchm1YMyhoWA6ZHGXKATLIlnqXi2P
ABKy3bytSdRGK0uch1ael30+l673tEwVjFNRhNRlwB44RsCCR+/V1hX1DBMihRwx
AxrGtEnR7lXDyWAAC3/4yUTxMK52uB0+RNt7kPg2JcbK6MXBMEoFa599uBm9GxHm
TZP0YqeTR13YrgDmtmGOrXTWHUlINSDR+4KYcZNLMS3+RLe4WI3165SCfOm4c+q3
vGsMUgYWG3ToAsO58d/5RQiTjnl04ry4zpUbpXP9BEUlNmGo3lmZRZbbWXCMLZ1Q
aQk1qBinTl6FssSPtigSuGboCuK1XXUMybnu/oVzv77mArdvqrPNsOozOY/hM+cA
PZxl5T9jyLAk2n5TmN9KsJfwSBGrcuhnOAIih47wK8TU2juczLL2L7lnVqygbguZ
biZVzFClc4z4DgvV0S9SjTl3tXYTNJca0vjkO+7q936R2CJJnUz1v6CLfnaSbAWL
/glXX7rin4CpP046Lnr3qTXlRvfmIQ6ji0NNnIpVlfBsH/YKb33E4x8bVZUz25cy
GcNz/2ulQBwvtlyyvnJl0NJxgmTujYJw15L43VPr67CoUAdKGOrwcE11od1Djyh4
GdeO9J64auZW8gadujj75gnbkALV7tjgIiWYZoxutJQYMZ1rRYa+oM1h6qjyqc+4
ZU5YqO1BbOFsOXiVolw2Z9G/zgz8JconS+g7r5SqcI44q+CRvHIDhkiNc71rOCMl
vIdyYiDMPdRa2Kbv+nLFVg1DancLg/RIUP8egO2+7GUqlu82r9A+LOmMUADRvpkl
14sd2A9RBCo+BcQLYlEc98//WUQJWFfO1f8BnSxziLFawVxkxaoq2+ZNo+PqxQ4I
LD6whS6uYwH7PD6Vyk74NIcyo2yXJSYxYUnEI/Mfs/8TDalAKt7fMLLU9VHfn6bM
Eb3upC0J9GlgYCFQ6UhC9Dgdunjub+4nYd0D3BcDVAByt48/Xngt6IPo6XgeiPCU
etnacWPngAqCzSz97qlMQP9GzbQ5QJhDMiQenuwQora/3xKUGzfnm4YLmcUNnlcr
Du2M094/26tgoZpIZbs8rh6z9m5sf0K0w4ahDaBKYrQZ1Ijr4rho2VDAFXEBnlkZ
Vqy6dzpEUWBMBhXe0lfg0bz0Wr38zkMhNryVx8ivOEogTpLQPGG/v9ACxIfd3cuV
yK8ydiZqmSCBlAuCRZ5+WWoPqiii9ZwxihMZFTWz3dxyjHDz4U+448DFmzOCzXag
3P6e9x9lS0baOGCc0w1Gtk6Y/FTRds5KDfukvRQGZF7unCrYJ+y7EUzubfzldq4n
jlbSViG1FLZfJer0bHQg31czvm4D17GMFY/o1PlZ1iE7AmL+ujGMGxI9SFF5yLug
COFxpmosnPVNewS1tZeSK1PY0bX7V/3MzGNYitLEgiy9oAAQjdp8tWd2bLL1sGEx
adf6/XnQ77oYn3N9uWFkb7yry6l02ogwD2w3bNpuKetao/fr9WLkTizDt1IyFf/v
LpBaL5Vn3ELZpQMAYxswDS4lSkoPH131o6rAFlBDiXSSJhi9zJFdtsIdynTp3TZy
+W9iDNODLAGZLDG4qa1EfAnD2QQ3U2jjU0OGq4oYeoP3QDeS4lgmTOngNM1Fj+f6
mishA024co3YYH48owQQIoHkEqdHOz1TtiMhEu+gVXrv63bozk+iPZLimdmcPmdo
eagB5KKwnFcpmT9igd2DsXddJCaoGO9gCM0e7f9bNe8RxWGqSln5yoezvr4xXKFj
OMrsSKb5bYvsG51ii38LHSqPYC7FGxSIM0Pn7/MS4p0CLOa5KJxayaCbUjF7Klk4
8rT/+IpxC7lQ302mMwY+CXFhdKzFZDRpUr+WC3oR7qlnL+7NbD+1hC554lCZ6Ovo
lITHsLfjpVArxoQ3xtfa/8zAxYQM6T7G5DLWnB/JsU3xONmTmGyivDI+MrcihucC
BykxCmZZEQ2XFBPvhUXN8iJeopOKjsZruxiCt5SQS/fqus3ZJgfaP6SFKybvY8ZP
RPi3kRVdEOEOoKSXfOzxVrujthATPU1q89b13LxI8QiU63W7TZuNHh8M4vUlmNfi
nqs5Id2N4715Llgjm1TwQAWIScABekSMzS1lUx5V3qfsfntNFM/S7EKIMj0msvY9
d+RVQZC6qI/BiMFK6vMJzjW3zvxXPzQwYnB8ObwyHxWvvtukNdE9iSVir9NPC/3D
4oRDFsZakxbe6FpjJNHox+ioNvhBPO/Fo/BKbKC9GFY2xb7Z6ZOIJYu9yR3Ds/03
C1NCq0F9+f6JUuRrih/BtnaQwLux0Xt4l+oho6Y7+ZzMucRCxyAbXHSHSh06W8AB
UuAjHcz1ZNd4yoMY9KmnRC517imxYeLGcin+jM9AYdYkjpAz62pNcjw3CRGN4GcG
XWFjSv5rd1OtAKefZklcs7nGsue9tBKL/GawnUKSKRmC3E8nLgCkROeeyXvdHdaq
8wBP6nm1qlRf3LcWWDoeTFS0hSh+8x8dKkLsK73Xx1UmdvePQcOZG+6IKi/b/LVA
J46w64EV3HEqq/zeFx7isOuiPobJZM6XzhcTD1BcOQ4LJnPYM9vxLzq88Is1+Y4u
oYeDMhHJZiYUicSe/S+G8ttHivHJA+NDXWYzd3TJIccsKu3tOZKgd0xiEOpI1n/M
h0RaScvRuuoFF5sdcjaLBWyBnEM1PbxC6ZS0VM2ZpsXbVqCvsOhiWSAEaVMJEfbq
N+XJEOviAjC6pjNlITJN6Gpgal1uQy04b3ubX7KUQgqdleLlITGnKB4UQeIpNNlk
DFAWKgC0stBz+iuF3IpA2SO69YufG4+0Oz9wQp1BfsgXdWVMfmo926OajOWYbTxb
ZZYXtXP15+goHVrRsjNyu2Ja8zARM3HieEF4ox5KlspGdfruqN3Q7CKuw0R8CC8e
YU5dMCKUqV9GL2DghGqOyem5hTpBkAwFoNflxYS/JEVGxqzBAOk7kFFD96mll6N8
x2aFaijyjYZOi11UpNz+b0qqrheInCzqwPBpxXup/PaFtjEpZ5SuUaMySpTpNydB
RQs/x1R6ksoNKLEIP9iaxWPqEyZNhqu0+VpxTFMNdYEst5r6lPqqI4yBexCEfEYO
EmZ5A3M/l6CDTHQ+MsPsaUIMdhCA+ZPaRa26aoiIxwnuksVbq0aPAzO1Ai/tNhJC
70jnz5oftowFJo0illfL9mnvrPM8hohMfTv2fCnzHVapuyXkrJQwy2hE4HrJSggz
wKlLuUs+FhtBP9cNE14hYAKh34BLWJsLe82LjMjM/y9NNJANKXFjmhdafERgKsmp
oiRakSMamlpMNFNjOz5zbOHXP+LtRbWu0aWN5NQ8pa+dm+tKleId+lPEPPdHj3iU
UO8gKViVDJ3rFSjD5JgyC9ym4v2XsFsKeb7+uK7rAOVtfuzYaKXoAojIhYZ67dZu
qDYJra8xHBvPw8Xcehq7xcvnu5h6JMXneRBNtkANdW5lZ4s56UB21g9DWvSfqHFS
AQvXvAFf4cFj0IFPAFXLIQi07OR+LNrk3yzTt8nh0Sl1m6ccAJlU8BqWpy5ASYu2
CT7+xNoPf2je7O98rSUdCIzd2arXLFi8fibkk7NHivJVDVOpetDmORRieTI5ZsCk
die0sl18v5CiIn95HSHwos+Zuq48rRid1MVCtoEiisfjGS3YfMQEQ5mMhP75DCoL
EED/vtvG+J4KLAPelLsyBvq7b6uhYtklkCCMeTZHyPqvU3PCisfyHEz6CYKchqVn
A42oqzgKIKufuErm8jW/oMUj/rWv+0yKLx3uXfU5T5iUo/WpgjmF9jZIi8FcpUfo
zLieR0H1XsGx3XtkqkGaQEK1Z4lAUVP+Bo4LBB1YOz9OVb44lY+dNjUaRH0Zv4nB
VEZHzJD9imtVErzhX2wAQEHcDnTwHlgLoJGVZG2YC+iq7io2TF4+KJi39BH724y2
RNDJ/ftKR7xksUnwyJah2qFe7ZY4V6ycT6QMy+H+0DRyBOG0y8POAIq7e48pmVlM
EpooAEzdo0qUeuQqW/XZQ703r58gJKbRZnzSeeQGRUaEeL5AL2EpV+HhYZ3/f0PO
9LOcBUFp4v6IgPTNMQejBb5F1G2yFoWH2cKpBZ4vr7PF5BcmmbSErpXuHVgirr6U
DvMwJa30ytHPbMPFzZ094lFqvlCyD5vF5bih3h3OGaTtn4HyKJTJI3j5np3AmnGS
s6mplU+k6V8dvNoT8SFp5tsI2XDu2pw+VLE2YNMIDg+c19MLNVpKGDmn3V8/vye/
kirSQHvOJ1zeXFiIbdCbD2jPItUrbDaVc58bgt5slBdGOBaoAi6pWMLlGTcZprQU
NdAbwwMu6ZBhcwES9nwcIRGV1SSrcraMcCEGmv6v8hiT3m3uOuJvSpkeJDzdjAca
Jbpm/sUdBk3ADznC4DvP7P6xDQ22Lu/3thjRwp2XlDA+36/7WqEA0lfOXRD3SXI5
w71BjmsNdAUSBisGKB1ECAhiacoGE0PWUoE0LPiM0v770k1xY2N1SZkeozOZQT1w
zhLuEbXH5tl0Pt5mgFB4T/9seAwo2ZOZJ3tbmTzw98zTNtwnyZC69EYWVpT+LFOw
cjuQDHr93o9psyrGUyP+W3u8eeP3TYTc+/weR1y8u8LIrOkbifDcqNQkhHhrSOh/
YRj9uECL8jb5vuRUVfVFFd9LxCf3nZiZ4rPPgn5VcpoxFcU3oLqrx688+gDzTpog
d6fL4z7LtDA9nZnhVmmUgjK+rococT1aQIkDCv6jfM0O+duZMdQMYfrYuK4Z5dhh
qU26ahJvY3lBL4KtZ/Wzm7VGTB/2MKbJNeMyDVik6XiJpOhCADM59Oqm18Bwru57
DACguglp/j4K+s8PLQ35KbfQGNmlmKLIQ1A8LrV2bqTmfM1dl9E2zvGnnEGMlOBh
weewImQKablIEm2Q2oOIkG/HlrWQmj8WeYRh5hAItM2AUD2dh35+uifExt2inu8e
YK3QpvnGu04fGXwVL3cF3t+4T0DBKMG8+0hwd96STfgrDuH88iTHKR6/uVpe2q44
OM529VtXp3PyHHqWUQtO+78Q37+JcYVL4IEMp8MbeHcKn1LGYLzaIN91Jdggtl3X
ZjAWYim3AvqjM1Kuxa8I6r3ZdLTT37VA2U4xINNOoFjfUAIZ3N60+fU8ESUZm1Bg
RAvsJuQTzP+x81qtS6abKK01Z208Gk7+n+CfB6HbhvtkU+qZJSfxrGXaIB1x4rYX
GZi00zLouCF3Mgn33s8hhFzY9ZvBL/Eykkcysg5wHccdZeB8Q6CyZsg8VZcYxLU/
7otOXZ1NH0GusPGT9JuzCMUiwztrvT2IdkIzJCeXJwAizLD/W/Q3L28KwYWdk2Jq
okBRGIqiGTIvzVogIp4bMPh1WqMlti5GPdZL4OanLEHuHQ0jC1KkB+645i1vR1A1
tWJHhcG33grLmVeL7boK6MT3vRERDQzqel4dpBxGQueIOrnR45S2iJbccMxeo1mc
g0Pufz95ZLNEKUcOfLA6Jm3jY7+8F04p5Zy4dncAsNJsD4gqxlFe+GeA2Inbk02v
Sq1O1+zsj180udsKyForVwKz/S7JDWw92iM5m04VzvoNMDpO+au0T4EPvCdAbUnm
DcHvGtspAO1f4EPAUhx5N9BRx3GMcmOmDDv74Vg+NoKjSxtOvgMaT3InU9ROYV+r
Nu0FTnE82RZGVpI5miY5t6K3zNx+t4ybiNdnZqr/7MVqnoiCtxof7K1zeMRUHRRY
5XInKoxJprm4lHDGNOi4wINOgrEOUHmKz9Fi3ahWHTvnAfO+7q8Wr5SoXzeNnLOY
oVYM0oKVhGGSJ/QseV4pPixOzYNZw4cuwHR9iv0OGEYTSUGdkdbN+4zVuSrpTqrG
5ZuXJJY/woVMH+q/jOzCrJjrK2P1zsZzYlk92OhRT+tpN87XM2KhWBpNpqQTBdwk
BI0ltKD2vTQ3SOJgJ1aqW22n+fAr4zHg3omvtlw+GfrzLngb7apwvP2c+xSH1pqz
biEdoVHCNU7l7nIOI7ZH90dtygqZD/+zWdfoKIJntCOZNT//W7C/pLh7VRHCVfau
/9Fo4Nvq/mZu7D1q0yNVH9qdUHunxUckTkybZKyZyVyyBShH7YPsLljclKQRQHkU
Es6A8RhiNQoJYo+Q6+eUZrNRwx4y/mAf55pkgyBiQtJI4pjMnrlaxWJGRras7UGP
4m6Zs3pjWj18a+NaEfvear0tTIQJpR+F/0DMMReaAjOQ2lCheADCSHWOWxlbWZ5m
3mKNUzp1wJ+Mq4K5PZWPDEVCshnCbUUjp4U5MSDHMnnGZqjK8YFviX4TV5XTimIC
s0fR0ca5XaHitFKbnVWUXMoaHOzDF/V4M+coktUkKX0qIEQxWVyCm0dYTQHUXTow
TrDFjaBacLkDE1c+VvJ5r6JkBMllACSlFvU+vbW2/QUHgBFEepcIJOAOSxYYhW3Q
06Xps22mAMyikvUZq3fImddAg8q0AHRWWPYG/m4lcPUbfhwE/n4EHO7yrZdHYv9T
AkVEOGg3TA5YeCuzL2fzTimBm7qj/ABa2R1NxECi7jp6S2FfJRopFDw9dgV+cY8k
BROwsgKZnOkOpJLSSxP+npCv81+RY8t7KPiRtFlW1vQtJ7G55mYj3pdU65wpv7p5
PYOjdljMXXSj7vSRVApfbdlk9v8rIVQvFOyY+KE3Jj6BOhg/6hnYNkh9Bk7FPShf
3IMRhUfsWKyFDb2wvNj+6GL1uUIDc+nyQDMBkwzfzl67TidarICEieiTlqiZSMOg
voTzCFW0lW2AH638JHCMD+u4mWd+J1IYq81uftdOjN2IVnTGIKIbZxvTPj6Qld63
qhUfArv+QRoA7AJQl7kUhMt3IHFJUPR7pkfsA/GuE5ES9ZauaeCaWdxUXGDZgKVY
8OWwuyxK+U5X8QKssrav6KS0i8mo65joW6lb6WO2yMlOOn1Rn8owx6wwU49YU03D
ErjHg9OjPJ/ipVCkhrg34S7bGVpx2KqEJpIYpa3EoVaS2uMvVCU8cSrUcEnTL0JB
yslAPDPwoFWpHKmNds4xPYvIq4nQ8bqvgYJU0G/l8ECE6akRyuL03eCsvjt/QfnF
aDiJ2kr7jCIET1wLmMfHRp+akvJwsFPVJrRIdKq0PBBnMZOUpJOfGb9GnSEVJNEG
+Zv45WPe7r4jrwb41jIrxNP3OcebHDX4xTlGXvYxJE9z5W89/EsCehqtqPG8lQMe
61qJXypK6sVkiAZExfrYjXWBxULtofmYCWQpN/xwfNCCow0qWGFtAL9j5cv2vksF
0e99gP3heDMYzuwZiZGf1uBpA6aZQMtZ+5mc9nCAXOFIvXk1tCiba46M8U70wb7+
RUvQ1sNyuZd6cipFvMZOa6PLKYzRNl+eve6TxIhZ2t6JBDTZ+WluG24coy4fH4RF
tUnMPM/PuK9N0rdNwbTL+4qykfLlLs9GoC6hlSwInYnX5NDP2ANbBMlOvNmyFQlh
MVeW4CjhwwjHx6enJblxMEGxiKixebu9Blcykq5gXJ/fj6YKQNGJPUVkwiIOsIs8
MNPfA11UAPKukQtXWFTXo/ZAjCj0GK1i1C03oEpcNNyJ6I0j0mXnBkPb0sp9g6Xo
F6k8ymBbq2fcC8BFsp587Q3NdNtUY9n0xJ/TBQSSf3TpfnlVPW+ygQNgLVM7nK7U
+SJDbWJEOhFT+BNvgWPQ+yxAD1AQXOZscRfxrcbH3zajif1GBfNAde4b5Sm9Ibnw
T3gOK9Z7FlJn5LuL9NDh3vqFWReK0j/BdAUARP/IfKOo7hhHr5hrURaZyb12oZMQ
YtpZaIItpMV9Bi0IA90nbhH2HaVTANrKNSBGeLZ4pyiAKvNIpgFdXFXQEjyBP7JK
CM6IAEuWGo2YqKJN6Tqtu/7QsO3eQHATiyQXoWdZiqRDhvDASiPVAamxJqzzLXue
WvJyIoam6JhcRF6AnfbNcLFJcgucdGqbTNyYheMj6gJf0VBI4MT2N4oxOC4Dc8WU
bDdKfmftdjEPB5pjOB8PJ67iIU8eBJCPmYTXnIaHHWt2qA/raDtv5V0Bw1rSVUKp
A77xF6IHAk8JKHxykGhtTDBnmO4GqA8XXy6RW1WT43qxPvi/DLnaz8/jKdYsF40f
zWMR0gUAhxKkyLPb6l6qBLZm9EtFp5QW0Ki2zkOJxdGp44XRYW2QxKt0j1bEiCRr
cETMEGBoETgNdvWU1SVx9H2TX+I3ObTSy+u8RBiQu+6b9b70z+BIRyGSMpVs9bOS
jWa4VVJUEKRakG+uRgwBUKdBZmxS/7UNXzygqMshOBHuUcrgeMBFX9RuNMO6ywpw
Ly2vFUC2cqGQPpunH8iWpLfke7YVEOohTbjDx9myh6y/0TsZY9oxm47RKioRLCeG
VHDuZBTthckJwkI9DJaq0MFPxrcx4g6bc5klC9Ff2pLbKqzOXfqS5ubUEZ8koGXK
r+K4FIU058J6RWAFRatc7GeJS5wMoXj7iXTTI/cYdpIUts1awd5EWugC4TPwKqDc
xWR1PqO9VgPGUXsYNnPygP+DO/1j0WKPrruAFQNPj6R3vd/xgWP+UYvCdLnRp91v
zn9FMAHkQkNRfp5YrJjrFCldElkh29UZ4U7Hzo262kSMmQBHVhijDuZQg61A1Ib+
6GuckgeLcDJ69XhmI+N3xEg8nneZIQ1qJ4dWK5l2rFREOoN4uLDCWNlh+pQjhu6N
ru3b29Fl53g/BJnWOSmXdR0Vyioo1qTaKV79NGAF/7oXdartoTqN4lAJ//LKiMfd
n6oXhmL0RrlP7I5pd8EQbZMnu11eFPHRSaHe+ed+/ICIktO7NM+mR6ntKUfkNEh2
EQv9anppet/Y+xtVfEpZdjCsSy2q7NamLzjLai+Sj6Ue7OZ1H0W2Dnv6Epsk7n2x
54ocrKXzOl5Mcv3ICJ6XWXD+U+PKkea38YNGbyPpCUFCt+r4fu6qBOLVPCwq1IRX
8Z0oDhGevI3YX6ZWu62cdZ5PQTDwXQ+G6owr9mVZ++vAgnTMwH0ScNsgG298n2Z4
Bci+P1JTSsHKCNmPQkvKrrboFiB34tGibGk8Rk6qCLh7WctCztvEaWT3nc6jeEeZ
0VqQ4uJAOLEdTvl4jVEs66SwuIHIAPZIFKpTsu7imSCEEH3QFz3TR42ZSdqvf9sK
useiMgFRxjN9tJ8TDsWJFTIy4ysagQqi+Dt+X82oOtzLL9WjrUwWlAg/PGi0OZe1
ejwFOx8ZgF9zByBevRn9kdWq+1RSbAid//mggISdmBoENoPXj/SEoWi49C+r+jeg
u++beqp7AScvv425Ih5rC7EFeVt7hm/4ZpJJPrmmGnBEk2TTFSgBXPBcIVMa7axT
8jWdzMbe3wcflUacQXCBLU/evNmAiEioFAWlLi6TWlbMr/smfNKpKtDwB+ciuSKM
yyCuDviC/CzxxeHWSwr9UGjTohIB9zjK1pzz0zyNFrjMFXGXgYWcj/36SN5JhB53
bmCsV0LG/kSK8cOouBu1PEeNBLrvyK9n9+3DVHsI1jJj5e63lqvR4I7/dtO8De6l
I8yNQ3x07EDYXeLSEAetlpuMtuZ+A5c7vaF6WVa5p7IyQAlEhVgnaVF9ruL2+XKd
AAXKUXKpbL6S750HYqMHy5/BujFV1o0nXhABIvH7+NwfM0xtpNdekEDwW7ou0HFG
+dgMdO3TU79/tPHh0rS6CgfOQBcNUwEVc7ML8JccVlhqfe56k3BDkvEq8bl3jlD8
JCdDtkq2A8gB1EarfOlsUza/KJuCqyzoWpvCA53yEQczomCYAyrOLbwrUHD+1mU3
widcsExdsEnj/wYlnw5CeY89MZz4EX1qJN5ZvoZ+7gNwjgZ3Soz5rNdDQHhW4mh+
90SyKQonoVHPOsOo4jt7FwYY7Byp8rQM4DSVj6QHrW0XuzsMcRgqhuJty0be/2xP
zBJEeq1s+5K7sM8czawFauUqS7Xru83a7f0Q4vzxpwSp9+8iBfnCTOrj/oCa4TE6
LmWHVrZXPHk/uQW2crJgevtn0LLERLkmigPpZhRxxbSafOL70GV2khVjF8fMN5IK
WhWeLTlfTjj8x67GcBHM6e2cXl8AjYRyFrGVWnxlJo25AO8JgUNKlP7NFelcwdwo
cE9NRTqLvt63W3J6Yh7xcvGkiFzcyse3mNZ6S4WjkRuLpeN7wYmiCcXA/+uqPYw0
oQvziwlsm6dVg+h03v1HFPYiDrw4uqVwre0iK1QZ2mop7ysQtXNQ2A0dPTH1lFJq
BW80E0p5hN2SZVTD/EeVReQn6TWxIbi9iSn/BG7yOlRF8En1UvCbVQdZ73k8d9h5
RnZmkxiWFvCuMcAlJb42i6V26k8SiaS9y0oaYPbaVy5lDB0q5PoNGeywMfAbQYXP
jBJlhqLA7r/08A9i9HM5mI9In1UlgbBWD5urf0DUcXQ1gOif9gmbvpH2U7ThSJIb
dEUBRusUiRc0IFPpf4y26hf2rlDkmnAH73tWjjgH5U0NlHTZEPonrbuKPOYaerX2
L6gaeprYRdEepsdoiFK13XLi7kC7oqV60C4mMu3rh3yjks16zAj0a6w26H4CwQhR
wApKbfqxo7nwm8t7Uk7g5vMhFIpUb4yV622IW5a10YKsS0IxXQsmrENtnCzudDZo
t9S7WhU7jTQ1ECuIwBg5AACdmOJNCYQH4vTMBzyZeDUCIy13u5sDBNrmXe/cvqSr
x8Rk9dCMNtIS/klkQ37rt6cfRnMVGb6Mpi27LaQv047ye04I3uL47hriumvYUltR
AX+2BtA2XHgtaWIHruZsrN+lu1EShMQc1EhbnBIZjLXlB+d6SGeyI7fuUuYFg/Fd
qQmm4DJoanByA+oUBPgWX2MRUPkdoul5FiH83tbEzP6seZSXmy83edENpJcbdOY5
UcTTHEPvw6PN8mVlgqAx1BketOfbCLLkxDivLtL5h4YtZ97aB0nOhj/5hZ3Ls48g
/KYji2Hn6gORZ6XfjIYNSmPhwS8E0s76BuBfdxYx/yWzZmCtqFKBP+ckQ5yig8D/
2M2Ho19Pfm/C+GB4/NXxkf3WHgr2iix8ph8//NfLjeNWBPF0SQ3Hquln0uyvMCZ6
5gxvPgyFWPqPnMe19sFmiJzEQifi6IJoE77Bj7p0H99yOJOIacWum8H3e8GRkfX0
i3ukuTjUMGGxI+xmOztjYX1oxlL5YJzEFq3RWIIQw3FCJS3L6N3ZJkCZ50aeogvo
n9u6Xz4kNYSuJ/641JHfJnZg6sRiGWwU19AQdt8fJtr/e4kBZhlDkf8D9qeNUkqZ
pqCYLj1ALHdI4LpCxcBebL0gouBz37tFMlA3y2OYwbCzWCb0dWbeQ6pbFQmLw+vF
IVzAeAg+1l0dtEGLkLy60Esa3jG9ij5lF4/iUejDvLcyP1dqx3i4dgFYoVmCJq2D
5xOTm8h2n2LQQMh83dJJP4BQpigBfk4FyVQk4ZMKMAV1ra1vIzgkLeqP2A4HgWHJ
xBUynjVk6kOTg9rrVpI6E6em5PjNXDzWxmlE0bpAHtHXk/LG5fV8Uzd5BtY5u7gy
YpP449kPs3UweDg3CdxhJpcAGaUJogmK1zXyLr/erNPp/LIsi8PpKlstmdX2bNrU
uv3VXcUJ1Dlo2iDtduOrE/1UnsmWJYKFdIPXX6pV7TCZ0pB+YAiD92hhfi7ZpVmo
k8aOYHgCMALqHLnrwH6keOrj8w1hwmCxEZLAiAuEeRKun2KxK40HfXkPd579UrWZ
ZwD6fvEZme3SnNBIC8E4zn1JJ3yUBv5kHcNlGcr1bkkBYEGJxxJIdB4IZdgnNSKZ
zJ1GrdEwCO7QgVFYGZiZM/I9EyEkhbWCasm7H454fgZsUwrExgq5VZ4HoNU5T46D
vQCpzRYqEPswdFgNwibSUTkspVK5/DnKbpAUl0MqYR42V+EDJh9IxW1SvXv3QkOl
1yB3OX5PqJRHckPETb2A99Q0zCxAiU2m7CvPsDKIBrpm8aI84gT/mblFOyU7tT/n
dX2sq0eyCQj2Tg+5XipOvewF2zshrTHxF8xA7E87bj+pAPkiIP59a/lzk3TG8SJp
SdAsuwxFtEZEt8kmSpsJm0ETFB790yRpsP5sMKrqGwdR6bpipKebrSAYVVFrAfYq
hfV476D683VrMj476Fegc3BKY2po7IUbSOF1ltZcTrbdsNWp5omNwb+Cs04VM24T
LhlIcIKJRYhu4oiMIsE58U4oBif0cU07LTq5lSQF1ClMakZ64aY47aOJehsyLdfY
mUXmkOfpDf++ySQoQoh7zWyJTQuRl4zeQJLZ1ClwFbFLuhnnsNW481Ygu9EUjxpH
EzR6PqdnOlOyKFX+8j2Z83k+9f8aFGWjMLbOXs0dbVR0xq1G3Z/oa4KaMjFhfLhR
0lWSJlOV2XmbpCA3nydortjLuSSHq+a6J0/xs6jmqi3dwQmjtG6j3n49Cx4UM8Mv
Ah8GOzLyGP4n92uAU1wTnO5QD2+6sCKRAm1ePojqkWsVZnrc7nXVzJX4zKyOAyUY
mfyNbyUh7WPm+Tk1IP+dU1/7miJPEmTC5ctKck00VqkaneL9TT4griAfycE685p8
3cOcHMdCuawEi/LkSQa+HkrziywheIiD+4qbYnI+S7R0DxWSTwpreU6yc40RpS59
46ZQHR85Mv25uDEav1emHU/ks4SBmxblSJCzmfCqzaOGo8rQ/TYil2movnavPdqc
unU1XyTRGvymEaQx49BBdt90ZTiOAJbERx+AGbz72ge3NJSVCn7wNqgO3rRF0RV/
+iKpVZLSqol8M5mXm3nwdamoXeKE427B9FXPZvs++CUgc7mX0UQ+YdKCvfSSPArT
EugSR161A92UgXIfRbyszOyfxNdYzGsqrYsLasTruPdPJfjVcbMpT8bu8dhhbflJ
zRMmwhRaqG4TDtkjbkfam18lIej783EjD5r2obi2M5nyG6LfE1iS9v9OMf+X9U+6
tCkjvyvr9J74Wl3I95Z5Axx9Q7/FMZQ3tLXnFq35slBOerNOcRp8kSmgSVPf0EcH
03FCAQIQZQSeoleSYReB5t0jcfDpz7n/42sFlN1WCb0BoQ+fv6wZUuFyyZJAzG5/
AvLRw8FQ3J291RL1HlPo0MwZrb0/+XjZcCmsOAPOuDHoWJ3b+lt86KxZ7QaC0kpp
p8JeiP4I3k3xCWDIjnN1vuQ0MR21LM4H5FhjtlwRx5I0Yq4qq/OSo1cjPuM3OOfj
BdNJ+19mo1P9Ykg/mPaOQBQUo3GMqmnLy3Zo+QT6/q8ronMPJd6HHe0e0EAHTAzM
HjKc031gaLbJRiKYD8Eqigxau75YFXTuFA1JvamnYO/NbNF8Iak3cBMF80LI1TqL
9Y0AnwLeKDCsdssJw3R3FYDzTxNNoh11YzQdFv5cVqsPS8lOUJ++8J47M97IjeS9
Wu0M9AfB9w5F/IR/1UtBS0XaY9FjS37FaP7ue1wY1Y6u30NCaMRkweZkdOen3/0U
XyewklLbi/C8Pa95ca4JJj2r0naniUAWz95lifnFB/xuvNaUsWZN4lq8rcJBw3c6
zL0ienxdO+jez4fXnfWBcYxi3Y8tTbg2ilyzaHSz9Rasur3VeThJ32gydzyGeyCf
Iv7n6XYrKi8ZB5FaulpenWbOEXjU3CLD9JLFvMBwIjBpppzWB+RoU5zEjEKRy4Ys
zNvZg8Ae4k3tFohH7qglX8ACxVtspcGzW9Iza+HWkEUCwjf2cWkjYcPvzYRmQjJB
pVVBjS6eCroPxnhdJFd/fD6bGw12BpUaws8LCId9+h1HBSQh/LvE8oD89PKR1hQn
Af6fEr3/J2iLrcVX8uS+txDBAe1T4SGb8AenVsqEnTw4SYEF05zEZGhfPMmM7eug
e1R06u9MlDjObEjfsN5/feLO1wvPxenZFUzx3tEP1NB/RAAu+Ewckn0PsjIoCJ33
6uvnfcaN4mahGIuQVzmFGgYbazu/uGSVX6sSOuJp368x5oefT1R0Dv7sk2SB0Ba0
eDcw0Oda3j2n4fNSvCnD4HzbOiLd3QheT6V4Avkhgm7lC2V1hZ2jNCze6+go02B4
Kmc5cv0pExi9sob3ZV7SdIdlt5w55iVvJS3rfeVve+TYNXILge4OK1C1Mns76+MS
uo748/JoLZiRw4CYM+xl/sSHR+2NvrZMZS4NKhXP4nVgnY2HFb+i1FEPGzf8YNca
eQZirdItt3PmMlIpSGS12JvYDHTiykdpCi1W+VlZ6ALJifq7tXIT0wDWsPtFTr93
z36PjC+qaVHdgwjDVblVaYyMiaVmiKiO+wlKwBLIF6CHuvN3UUvjRKteQsjVWmP9
N6O3ZA9nCeioiZRdGDdP4sipH0Lh4G6vieTKJxT9zcgYjnD53/q9WquS2lHd76SW
cq0+FxgUQnSarWimZ3K6h4PjwOD/e+carNYkIQNgcnW9HyZXorwt166pabpYYqQn
uK3ZS854O9nuYCyP5tmyN6t3vECB9FDSz8Xj8x5es9AN6aUzX3DckZwqoSzwhMxQ
9CPmZCiO7YFtkPojQwPkuUVMYbCZ9bMQ/r3hk8XRddau2cs4wr/Mjtsa3KxBrwzj
o/5qXZzm1ysSxPEA0TzBNHAT1+Hu0X4xZf7auRPM3+Sq6PqoIH6OC7dE2zEokLvY
sHe8pUJ9cOk8FaS4XQehwEPanRfKBvsg6ry8kXf/36FNjHUcK3qsJ/5wlSJ8KdLX
kkquW3wZDDQ2598aKIK1BZXipnDC9vYkr/oESGpmAchDQCSoa7WxZyPo257GUYlj
Sb57aISMaDHHWIDcu8NTVbdufLOOyv5ZMZ3Fg0Q5cifdquO/JTQTuy44Mu6SmrCe
n0QGIoOxEUkascfbIKERgC7OzoYvkqTC9eHI5vy42muLICL83OhBBtjpXJErdZn8
hx2U0WMxngRny7/TtNoSiuEzsn/V9Ath2yM0Y7lWMEtkh4jwMzlw3nEWPg0dM4+o
ILi6i/JOHKrKPFgPKugaBT8w2ufbtLyg3BSvDSk2I63YSCg7qozwBid9VmCWAdKn
GHG/9UOavY5ar8gbF7dDIMTZVV9lJBovYgjrEHUQlqOnpDLhhxoEHrrOPpPVwrCj
s5qFyQ+UAPUaou8ZlNDFB9bQeUEcqi6uVFmKgzlHzDaRp3qfaEfKdrVaAmdflqK8
IUg2CvvbjF/XukHKrNl0J+anjFLvLJXClb3PTstUvbRAcBKRU/0E3c8hQZq46/EU
nhD2tKzpNcECUBeE3bY5CSv/WPekgcL+ZyLiHIYsq7QwWXbaWInhqOta8Fy3rKCe
KKlfgyD8U/fMXSDcEppJ5gnTpqg316Li+QdXkUlgZ0hb2ttxZbL/BIdC9a0n8Wt1
X0piBMQwc+NatusYn09nDjMcWRx4UE5FOPgVJLngv2ZFEHhOHxN45IPszfuijlEA
0bqtfayPLlltqMHD/UxJ6AjToa/p8iywH8L6Qkg7atBFlVCxBB8wtg7ql5M8HzKv
/Kru6QdIolrW9V+gI+WfxEAh8o0BQVSK3M4UhpvF6se8PDOn327XfQtFDkycszCl
DTXSX94UcMI6GjOED797f4FHV43ADU6ZDzgBCQUvi8gvCZm94pKxhiRuwek/bvXM
hajSslZtEpP1Ln1dhq7lxbwU/JjtM6KHHaLn3D7bAY6HTXgHjZCj/PWPenMNoTOn
3Rl9HZgsiZQBTUYAMCDw06gJJa4AmkzHlyYNd4ySyxbRpJM9x+aacqT2GfLC/xfz
DWxIbY0Hk5ENT4yE8+yGDcLiMv17/S0YMc5KxpDf5ZXf3cMuN/7AaQ4ZuVakpBL8
SoizowcFjETB7QaBDk3P/Ud7iyzm2/VHxnwgOIcMkGTao0LwIawHH7ipM3G6WPdp
5sK49Z/McvSyiitswAq/dCW0AxqV8xCfcAhUsGcq6M9YDKMv/J5sv/OtnIR7hY2D
jFClMjLQF2KlbiwyyLCWc19Hc1iw0tngkdEtrfW9QRAcfgzzWmvh7cyzWX1L62dA
c2VSC6rgArN8MFhHO42wG66SpI5Y0phiPpYXL1tyNALya45xW92ej8m0c2BmnL4Q
1T+jzuyeiWYoBWLlJP7fgphY7D+UCgPcAe3sS9fcob4Lq7YrtxUCPIB/i5NnMWTB
CppdBX0U1iXtpaYzkho6lQhyizKyLyzSojyJu1e1L1KqVdT2m0Jn82v9hM4+ztI8
i1X5l+Ia+nG/bm5WQYUJrzLfn+WKFkGKJCR6FLa948IgGI2bEx45r/6NoE0YbFF/
GYzwwLNxQW0PUOp8vE+sPEMHl5gFL8UTrdD0Z0nrkuVFS957RrIM5Z3h67rLPVOU
Bn8ZzFdrfa6sWZx2X1h14CAATPANbXC76zmvspLl/6TZ+L4jsrGXi2Leu954qP1c
isk8HHMCqrM2GUV2QQeQTmtKUns7SQdw2QqemR1a4CoHPmvGaJAEgPTKVA69+tri
3FwpODOX8vdH9I9F6uqJwM4g63lmOTafEr3VQt7y/7vHBALxhwHcI8/RcRE0cA6L
j3D/BdAnlonZyxpiVZhvFJYqWaVtCfsG0vAT0wtUa3WJ+hqEEcctIUTKObC2DO2B
AIGPdMwORyMdwDf1ICqJCJnD8CSpQ4HU1h++MxkGK+gsfLRQ1K79vnoQqHZJ4QD/
tQmXWiO9t6Oyw7ayzIUHYkbiu88G6Ws/DVmAGsWS8clenLSyo/UPAwAhXDsd+wx6
EZ8TLy4SuSW+mm3Fq6dDjHBuJ7KALPO+SSSwzFGC/uqE/Mnt/dTfxtzIIwXpRByN
y6XEBX+YjReEuf0IMeIij+kfNeezMYpBqWsEMvxYuayUelc0uSygHQ6C4pKZXg4P
Tc1WjgYNOcyLueZn1vRo5CBZTyC3+6xcEQW8YTS9m9lPuht3piPuoBddexN35tZo
iiHfYlMUT/cyXctYpUUawR7mKvEZZKC1B9K4+3+T6TY3WehcN4kUn3XlFgB9xugq
heylVXFwWdchmDjGCeM7wrMfdCjgmLr0I6aM/1OPwbN6bWu2A5XGc/xvxmhWkgAB
4pmTjsWoSuJ9VpSkzPNrOJCcv+bdo+BzBd7XWfzUF4r7FcUkpukMa5yLDcy4YzhT
gJSnwCJRXAomdVMaF1p8v/g0IMyFijSsdDl73RofbtkcvP+iepK83OZqY3+qvXf0
lbj8BJlYEovdeTlkTnmjoL2+bkpOT2VKdGVNqZSnH2c5gG2DMdzFOhQVJAnU4Ryy
O1E8sjRNEOLp6A4ey+WOm2KYhe+vRGk7E+XlvrhhKc1o5G1dInyl4Ht78c99FcP+
lA3Mbv1SM4Vo6uLHmqfCcz7nj5SpiSTVU9+wRO96QuCmjI4+SKtTLqHxNLFaJ/9I
knLongKvkkjXZOuSGHo1Mct93zAK2ZC81gIzER6pXdugIZN/F9aSebK8E1/FfQI1
RvA7X0ze+TEUWVIAMVY2A0h7WddEMI74h1EsD1sKpYZ57fAn4ToAwwJgrb867ClU
suzIC4hEhFrjcZxK6HD1l7PO5glmzxYnaQ8mNJOOchaKuOjGs+UGvH4qBzBxwyzb
lHkFlOj1CW3w8uRxU3aCLYwVhHKKEel7CWlAQFhP5H7piF33pSudB5AwTiWhucK2
BKaqdlfCIS2iTettEBBEAqEyCAwDbCYlD5Je/1C+a/RcpYOqeeujpSwvKsXGj6pj
hw/HfkMoLaEL6KvRawWqMWd+UTF7o1IHIwL6lTiTenCBDZnj6sbmezm7pUDVCu1x
gFkyQbSz2RhVIQA6sZabibFcqHV8PK63gAbtJois766mYkhW+AShOMFjSlnrgJHJ
FazqzQPZNqBK+kWOKN+4wEBuufSnrDATPVjhZiMlsRGFSnvCZHXG5blm1pYggCal
xag456y5vreyYwJLvMFY10u4Ew6rIe9DDWa3g7BCUn0Bj8aqidMOUuPu8kOMU8eo
ix3igOO4F2o7lLyxopR+YaQDKWHDoI2u/aMpCyKvGIONW3eLm7LwQ3XzTD2JwCFh
q1THq6rdIx0Q8+ioI/cQOEVR1maRY0J6ILo+pjSXZwXsLkSYWCbLuf0mzoKgiU0u
u7Yr58ZN8zCrWf4bqBBqs9Llexx+qvSsubW5NS13xLVMZIpal9A6wH8waF/d0kt9
dtg/EFFbilBNrEofKh3ckzA05cmw3xIn1dHj9M1tyPRDwv9y4QtS7/03DN7CVoS2
3zMWK3rk8IU7ZJmXJYJvv+txjZz6JfJsSyObGJwU1jlao2iqOtK8tka4T05Lx4ee
eaWh0IDkRCABz8GJaCfZsDJrFp67KHas/BYp39K0XNpv21VZ4K25HmK2cMiWbboB
IRYdXOdNdnDf8MpWN8L5uOazmrfPi+0HH5IKzoty4LagN6o7JCXAoM6XBZeIa+Xg
9qnyndkv5vzLVIrfilvryzaQee/XLzKdiSuT86h8F1xXo4TpkQKJlOsLU5yyA0IH
hPwkZTh5ZOYIRdz2dRhwSAPrCHRNz/U/r+UojtBAq6zUAEX9NoPznSwHtp0yQv59
5xlDY/4SN4wjjkQq2tIZCi0dm5wGSeFL2Kllzw6VHpqVqDzDYgQT0SlF1nP4v1Vn
RZmFw0gBvpIjnAHuWvybTWXNeYapukn1kla3M3RFtn2qD/eguEw7qJey7ArzJ0x8
eN8uXeqpGXGnj2R4HOiqEBv55oMUiM6ee01ByP2yeicchJAWETjbzsqmKDcevQat
N5uEW4KXidpGqH82Y7ixj8foaWxYHrAaj/RtAa6lN4o6TDGOGYowVx7DIEB872Y7
BUHS4GBqu9uW/C8QBNppCtk9N3N5AsRniGPUFJnV4ZRlg/nEPaPQebnYG4OQ8m0y
5f2H4USHxD1V4FCSNzOgj/+TT4f/dAnRH0bxJ37CMNrSt6NOWu0/N4Ydtlc+CkuE
Mp/GNOyeq3k6vpcf81UpvU7zBZPmOOSIp9BYh5Vu7SW2ahdv5sGAv4KkNx+Tb7B5
E+TL4TDtH4cdGiXbnenIxd/zXm61q66b0YyW0Lq7/NQGYk+BozvaYFWpfkIZGr+Y
BJj6VBxLSDRVAmYE90slJQItnt9UJ7QVT2/2lChEMA0DKfsyI0F6JXcVx8ZlupET
70mxgyHpTy5TSecl3bqsddeTV68i3ykKACQxbsAFkOqRyHQ6dIPj3EX2dNDcNuG8
eaLUCXxYWktmVttDm3MRKbc/3KAVzIunjQYxiGesM6rghqibL/AOSnK/ub+xk+Qd
OR4c0WiwrKypQtP8oYoHM8mM4gtlhp0D8kN9vN2DsW0PUG1vMlYjsHdvV5XXwbR9
Saa0GLJGMC4XgI8ZGdMObShSLgqsFML1kzqjU7iT82OAufp9VQRN9QJe6lV1V7wG
HnakKDx1nbqyuN/lD6g7hsiyAo2H9jHhOcV1k12MIdDNOnqIA6PhBwCtN5JWnXsU
JlQWzI/Dc63uNvsxthvDk8y/nmtKWsLFvM2BdHvxIiwHOZh7krnl4EPSCX7UatmA
SNMhS3v9AoHB+UtH7Oz43kvFk1TaVGsZUVtaK9yDBbyTQXy0z9OdCyv05aQh7l59
p93QDhD1LWDolVHI9+CwzSB3K+yd6v4GqWMO9XJv8jH48NHEVwp3go+rAMPCRQxA
r6WJ87o122WzZ1dm6o1KzTlW/d9UAIM8KZ6XtSHVM9msN5KSygHCuOPv/UuKGLVG
NcqV1MeIBEmztcVLTMZMU5g/v/3YpsbCuhBzR7XXku4DNPWKeWXSaqqXnOWqFU6Z
ENoxNwmez4MGZPfF6U6bVBMFExiSE9dhyIs6S/af5jpme3EXr7onoaY0KheZpr0M
EP6lmYxAKIvvDVn3sz36c8Ws96x+ezoGmPhfBK0om34RWSYLe6vETdaDcwqGq6cv
8h0cN8/cxFVH+mbEFUnXR6sr0/ge1j5Rrf4xSxul/FW2YwO3k/wfd8laWf2pWZTt
xxa6GZVCf/PMRB8akGiiiwXHaOntJbr8/3R90AuKIznowO2HAFB8xOIHqOvJQ+Oc
3jZUpFRUfJd3rdWB70MLWic7cylveZVQY635W4tu3ulvbeE89bKKmgwcTtvb0m1i
MFVmVxFZF60k9oND5RFerMwiT1gvOCn80BbWWOrjWfhypSfNylb9Z5rYWXNPQsvd
xdVfauWQXtefqawLLkPYz3sXLGzGLDcPCqU6NTzC5oignEox80aPHQqsVMrQAK0T
vdDc1WK+RCOqtKKMsU2SQMyis6FzukwbrZuD3iVv6NzgQCaknn3BfaZOM60IHndu
qGUJjNQO49InGZr9Zq6+xDljTDnywOrvRZqaS4mOn9A/VW0RCgCAfgmq2g9hqnb7
3nDdM9mEbvkhP1u0djvK9UmZ8gSZHMS5CRInzcevtdbHlqOEL54xHAD2yjLgf5LC
7P6OZFCy2n56lTcB0+rj6SXIigtc4HJtpbMOq9tO+WQJ7ViLt4YeoHnnoZs7DioE
7RCDQAVga8STVQlXybnDboC9j1vg0wUmgA+VH+ejki9ypqZJAK3nsjKRaZADqVpo
wmtaGqjiZHZHDu3xOEymqORyV2PoNZXw0LWpdsNhD+YAHqp/qqEBYVnwS6iSrRTv
Q4FB9Y6LHlByPj9N04wMqwc6YMti3ZEDFQ5Wqe7jz2l0fT0IrJOk+XGypV21WZg2
hllZ/5Sh76p4JV8Pc3J+x8YyJU23BTPRilznDbtNiZl8xD5kmapAZtgeMnyPYQnW
qlFIXPJ9/Ocw6FauProCxBIdvbqxSZyMN9dUmhW2qkdhBlza3v3V+1MZCGkGpYso
TZoMx7V5ejfxDiqwGMlHAf6Gr6+viY7n9r6fL0cAYDcOU/ynurd3NkHGlOG0Q+Vp
JWtol5oD0zfeCNEebFQBxKBOROw96TfUXRlIq4xSngPfTGYxVQYhe6toMPWe0tTY
+O0ULjiym+4AK0awRIB4ft+QJgAR6ltRUr0jwVxn4krEgpQZzrj+dzUIM1QCPC0n
PJ3bvoiaGBygHgdWTyiZxA4MJrWixquhN5XSpnvXXz7A3xbMKkJPYGrc9UPtPfq2
z+N5pSGO+svJ+JUlp9AA6SI7NAoW2JT8UZBSK2kxzx/6oONMd3rqA6e4dRdztanG
2TofYv41Ti2MlWTNIUNNP6wMCr1Tc+jqiAoJ3Pq3gy18v+AblGPrlva/QUgdNFUn
AghEUXKsG9KC2GRGxiAUrOzDDctMpi9W2NpGbK/9hxWRqpVetDJKG3tgktL+iuUw
8DvzAapOnAVA05Qdn8vfaLh5CKK6s//aSdwFYNfpBGDX9iitDESaA+WvpFJUWZvI
buWeU418utvh2FcvN8nKiD5ojSSpn3DXPaped8BUAteFYEiAFeOYwcsCtIqHBnZz
3ScDYXcnm0nBln7ULjyhWMio+HYnpHnaLyDFOsVGNE02vDm5/w7xUzclY/fAGlgS
6ge9hZAiHMcsJgftpDZXacsD9taDCjRqXMZQlGhQDFwYxHWcv7iAD+mxOXNoTZt4
p7kebFSq2xyx++7vWJOSz1E+1wf80SmFlwOkN1sV9RSNtYMOAioTF+D21+lKEhTq
2o6hXLfaUd6WcsSbI1NLRh+zEi0L/gM988OcU/xbI1lmdlLCcwb0ViySWXdFyLRi
GCpI9TIIWxLiwjgpGHI/k7T7mo9shRLhWZIEIv/uGJTjuAprT8ZreuPsPalL8/Gr
102xLRbQPNU5OzSuetfemCz3ojQm8+yI1zbkbYJXLSIXvEl5rcG1K6LUKAJ1Uekq
mxUDhnWi+Mqw7kNScJ1STGUGJG7xXajro4LPJllPqtPm8FzQUtDtq05B5jvcREDZ
qEcAJyeDzkU78U00GE/Cdq7t7XHutniHsDy3PLHg0rv4fRaaW8on7LBTvTiT61CS
Nay7FXcGJWtOfv9WJZlYPY95NnFhLNfe87dnoqnZ5AXLYkQe+/WZqE1SdVE05eZC
poat4eCIS8FQ74E7l+xE0SwWeEWzSZDDMRtq7FHgqtlgmJwmTVd6K7IqRX1jbify
mR4awoClt8tCZ/U+mgdsMWrwprIRTicZIsIDLjdlEHbTKCOwQUu9CGeHA//YctbW
0wgrAZ/dxnXpiLYv3ak+h3nAELd0vVdQhmAHpzhLOMxYMb+mfOMWKoc6QSNX5BbK
79itltUoWP44wMdtXPuVubruaZ9Q52SCi+zRHvBy2Q6Q2Z9U6sGJjNa79kuqeyor
mtTbZ9iFLOrI3palgGAVe3+Swa7x9voLUOQKuXCAp43afwGoa18/2ojGt3gcwObH
UOyk0lNMGm6wmtctVsvFw3mJAvjjwZSkwscnTbGRS36Uym92GdwPOVLLQCJJ8EfR
8se34IpKTmF5SsrjvOi127YiFeoQkmgXWBaA23wXBQa8uad+xVecLltac9CQ+75G
EzFXw7h6yCn16nosBs0bvTqsps9F23aXFXLiALqI+WHB3AxKHNUWuPrc/j9kYiFP
3x4yM9T4He16ewA+X3zvlpkXnPtg21um1BLt61PZ3CcpqRlxOq3Akph9bErergm0
oAwmEG/EQ3GDXsrCBMWvRrxFMRW8TG2VO1wjlH+Dar5+zlsf3QW2bO0tW11RRGI4
XX+mPLCo3s2Xp6jTppHbcbAq3YZjHhjZvcHApiU3pRUZLL5tzzHjuRB0gNH219qK
NlhSzgvkFteIY1ak9HErpAxhQcE5EDgr7tkP/Gfd40vvWbQP6Ds3jLLjWArWrDxX
xs2ZHQ5fOrRV3B8xoDVDIMTjvCS9Mm/JzxSMKrZ4/EITGD/EVvSxKF7fC3D0hs4H
LDRcDucHghbnr29qPetWzKkx/nQcqlQ4CeZ5bkMOR2jt0mPWwLlH940+jGdPh0u2
4j+s8irqfSZzP+cUrlK8QA0RHcr5ONhhQo4nStNKkefR4P+icgZrsy5SOAtnMmpf
RdNFRSU1r3Hu8I2tqtyvuUBbJ5K1yFt1cfWmtwza9tDyv5R6iplOuwjXD6trp1Bx
u7JDjqcm/v4UR0V3DztqeOVGoCwIU/jOHg/1Kew2bgd0FJfdZeoFoGVD0V+CNpjC
PJVniwz8zbm6rISgUKqumgeE8v+0gIkgXQkXMrPNGCyO7MYXkD2yBj1bMmTMsMD7
v/ikbG9HkL1MV1p2seU2gqKO6jYqvDFDHmUEf1YDrt9/IUhw37j1XBOhFe0k42NW
k+Zl0SJHM0HDKr1wk/v/m1quqER0vFcpmu+FSx1parQPxrmFixr5b0U+n+ddAv51
tCWYSoJ/YZE5vuNm643iyY6S64T7+0u4YKMwqNPrLUKfGuTZRe5vSNSDjNcFFSWz
SSPU/pJ0Rp2Fvr2kTYbHZxgwclSD5nXcHVn1XJXaYT6hfyXJwU3wyRe4V1LKOqTQ
iQYvLnH03vJKTHKb1c2lSIvlRdA7zkhu7lnOhykPPcBTQFHTVJXJ10a3904hPaSK
rHxdUVK+ijUjoxpvFDqK5BqtF4bfqc2yFgHEHNeUr7hXImToUfomhVHSWHn99tbv
t+X9PsY1wq6lXR7qCnXWyNTxi4PhFwgyx/H0Pz8rZ7YG/1VtwiPqFtgt5GH9qxfZ
ar6k1DYGp3/v879WBL9itARBgs2jkqxSLGWewV9WLsEzYwWu0P8mcQ8w5YxVBgwg
F7jMl6ebD66aLGzlXIS68GDF7J8XfQAUhjGv7ECBxG1R1b7/zsT4polTpwh4nX1K
XI/uiIkRbD3gqvuT6Uvczsv223xg37636LByTdRK05uEvREMFqMDb4OwcradwU2A
0PwKz2Ag/JypSYmguGayf8fuz1b+SSGGamTTtZCwckp+1mmIaCs9hIOtHggZ/K0T
cbA6r39BvGKjzaaiZ9OQJepabrvxk35nGhLcL6xIwuybsYxe0PZxdZ5ojovLdc6v
FfoOsuVhvSp/ETsdzPY3rXXiacpHnlqZWG//bkQ3xmYpA4fpQir8JtjAxbYaeNQB
R0KCqqGWnaKT1WGRX1BU1Eq9xsKCm9chpQyAwCa9H9zrq/0V+2E3U3DQVVR1hauC
8vn25zTxjFB+EQ+TuHnW42zwR14u8NC84lCmpqULPhs+rgneMbqxPL6ziNzYCJsx
DiS+bTz3jrlDAriwXCs3/S5BCXTNMypQtGq5IXkxD0z7Sfa/vZ4fbWMk3+RHGkRw
GY3ce5CPlXrrCzeA3jgvJbiol7yXhtrn4SUHrhM1IpjQvngBBA4UKSaeyeDcJnR/
qFLnTVRi0cZRkjHcD3l7DT0UjgqGiyZcw3o928K2RDrxDd9l4DQs2aK7aIrZLTaO
zKg2120vRA5Zrz8ol/vQgc3kKkx1Y2Z9j48KRfBK2RXBw3PcojKinFG4fS11Ml3p
Nau2S1phLPm313rV7ITY7tZ+VyLCTutb21Ow0MH7U8duR3e0k4CL5ORpScgfvxjC
qsUXrsF/w5ia3VZp0jm5sH4lzY1z7095mYE1QgXhi5l445Y5AZPwyu9Qmv4BWfG7
HYT7aB9JvoeoaAtZDjZIMDMi0x5sbwP+q3NDp26SQy6aJLxoZC260tDKoE5E145S
eVFFgfMY5GKSF4NRwr6qTHZq/xsEhVDG7n/xjDkIzCXFKrjTStnWunYOiZAzdblY
IkHXE2Aw2p0uuHyJU7lxkzXMjZs7LGH5ZE96J7A2qU6a58yIiUVqOnuJl/ZB247O
ISDEipyWMCI/Q/qd7XaKv3B6LdkSA9190bmJkFKh+IIRnvyGxu8OZi5j9kZh8XgL
FZk9jMrEgGwWynXqGaUDScB8zlKmcmmdyYKrdWOsBXm6g04XuIUhfcGOf13EWUsl
XTPq0+7vCqH+FT+hV4lgYSFpHkW+4rCKOPbrjL9N2ejhqXtZND1m4Zbc/7dQXTZ8
IPvOcFFMjy2UduUGWBWaPBfbDRrdWC4CBe46D4O0BPhjcBKHLZ123VdVrfDqhfqn
pLRd1LUi6iCCSD5Jr+0yYQaTysuRZ8+olfltXw7l9GizsRW9ZZnsRNNFFg7rfYoC
GWTdJAIEofHNLPNS/3KZRCFnxt2Fy8LVbTz3zpd+GZ2SAlUjPJ0oTmpivPYrRuUl
4ARuyGmariPfUpbdQugeVWHeenFqvXuDpx748DBeVrhfOGFpwxaSOw5qnUOIb5m+
jFOtXRTCRpD3ItCalA/dECyOJ4Pp6TjP3Tp7hJcS8wPtB+JaRNBG7g/tpMEFHbKB
jQUHOdoFT2FnvW+pMnorPpd3pFDhGJv5QbdHz2B4aK1kXVUGNBUXSSHb/Vw7OeL0
30BC46oAbu+hEhppkrL0I3cWpDT1o7tzNGRJEGH4M/RwGK+3lb1ruq/+2rcSum5K
hiWnhN2qTNfazzZ2cpYQDgroOLcYtC7zTv2seJCdDlW/SnE5gJa2k/9oPxY3qXD4
kFQkQOXrk3a+2jPLE+loIXikOlAtJgEq+h1Q9VMGyDSyOZjRUDQlSWoFrnn+0Ngy
dcWlNO+XaOBKdKAtDZhQfXp2j5JpsBhwCSuoChYlBdvxVQdzii5FlpLLp1NYyOeT
7bPCEKKwoffSyO1WO8F4liX1pB09qcnHTyMSNgxRSGa49pCSosL8B0lD/RdR/dLS
Lz+bLT07K0DclKhIlU/BsBMtBZKZQ6G7GmjTUwYzNa55GXbjtqnE51rBvX22jV2f
ZD9QrwWMefcQBeCqX5VJlKS3wK7PsW5TcDtM04j5R2YiRffcnuj/ApraNedsBK8e
DWR7PxZ59BiVmp4Cgjxyjn11In0/5VqAVLKJKtn/GHQ6F/LZka+FjcuNyiCo/TgI
q5N4ro6s7qLqRs2E4kupzF5Qp4SQpWbwWnaBxFlYuLvrGlC0MStHX4bVdbUVC20q
QId2Ng1ei1srefUwnFuaNm1Zv3IVACYYlmnedsWMSiG19p04ETnIGuNlj1sACQu1
WuMdHGCqs9axgXFxv46Pj9+JRm79pSSTKC7boFz/woVSFwUjQwVX3iU6+D8QrxBb
hDlOLBUhbkb0Y1SxI4KhIdvR5og3gdC6EKp59n2YOZcZCJi3ROWXtbsXtPTqI9I1
rWDlCgdxV39q3QWxqEzXQgLDmMyBww5JTpK2ZmfTUHu+V1ApzAP8qY7UUJOs66OM
WgSnq16xvW+ZUaEFzSWgPG+jl4TZhX5SRbKHvIZVJz9JXKLapHwvZ+5LTX/X7Q4G
uUoDs4w7+INMn9SsEoIUdbigHOcZb9ZeuNoSnSjIudGfInekKErtbbfTE/VJOkSy
GwCaMSPz9vVflfvcdABcfeA/tBPpC+Ow7+pDOiBHsVPTyXM7pJiaQzNBkCQ7cT6y
QkkMwAop0UD3344inGRmC09orCnR5RIqVdGrl3xc/bO+HWRNrFsqHxl0V86ucC6Q
xlKqnXIocVQkVkVK29kyIFVLJ9fbY8i4AmkWSIRPreu6JtJB8VgfcGBFr4e3r/U1
yv+wbmlCtKoBMqg/dJ8u4TDcaIPJmIaV/yUwj58rhURRVMWOgToUf97Vu5l60hgj
g6HDMuAKCRJMMXnEUz0hy+GC3cesu5EJMr6dktf+bOdfLPKY9QU5F2qYIT+zMltd
WciK5sepeaez+I7XBqYxM/9RzHLluZPM+nR8ZJ+0gxwHfweFmNtTZ6pzIqxyknhd
XQBP9RpnN0dbi4Wx9/XlXFZOdQW5zK4rttzpHZsXLSLNdohiuNyntlgxRaEHFWLg
A+7PkpcBaD2UZq/qSdpb93UFRv5FC+qDoqJt+jy7OglA2SAbDL7lC2Dtyli0QMA9
pmp9ZFxK0Y/DPr2GGmrgg4NaVgZMyFMmmWJ63iwbulCK4IC9Ts3ihc8uO91JFi5L
hFx5UQaCPQTj63KJmvSWIUxKBDODJCcKTPifBEJQ8MEY4q5xgRlyqbFwOT1P+IDC
LeVN6pDANHvzxsAEqVvLWEEU++lqeF2eiY5aWfxonXaRx0ofcGUVFlfNXtNJgk/G
W5s1cuK3e9DFvzWgJ9oiFtMSWB7v3hYIHe01OBqINwYF8shpVt7GcwTBvda2HW0w
SPs+Nl42Yoi3XFrLoPBBJ5fCV35sMXrxTinS2R6N7gHKCaJxZ9j6UXirk/0Wrogb
K1XYfHo8qe8VqTioO7cMx8VsP+dS9KfRv9ZiWGvqzKd38TJuqT0b7BAM3Cizkqfp
K3JUDWZV0WvrEMJ1+dem4QIILTPPeslEiqaas/FMMRyOsZ8CeRdumfi9MN65rHEx
oV5NfhYSAp3j6uc1Cds6TFuBSh5b7khT0PL72XkQYAgROQUasCbLIlz2jrGzIvfW
mew1GclRDTq012Hbu0t5wc07GUpjroVfgQ+QHpCVpljlD0tcMDbQcQ5P6RPHOJfE
JDbFnaC0RffmUC38j1DU5nyqWKofvT914Lq57EVpHQNWpk1lhNr5jADop8cDmt8c
kRYy/jFfwbsObekJmSyM/dX7Mm1Umq//QQtViI1RAEeIEJcu/DY1BXqMStve+BlW
pNLPA+5uqVwRcG7EPuvX3KNKZTrKLxqjgQaepKFFNJZlRlmCKqRamQhLh3ha8e9l
dJ6UBs79kXYTDeEFFmDFk5qH7TEjr7Mje1YcP+bIzo7P8Ebvu6RcCwqRWXptT8ka
sHsy5Su/d0vFXq5C5HfAj6059EtP4Nfty+yTYaIHEd/6ZHiMsr8jg6uVDld/av1J
ThqzGrSjQmVZzHlKeooNihAhJTuGoUqO8xIlZvSUK2Cc0UTlJ633Vw9gf+LNufoK
+UlOQnQrlpd+k2Z+lEtfsdilTxTjfuJzF7w4pntAP+BYibaliuWe7hb1DUWaviMh
pu2wQPL2a7VHszZcptNOgGSwMR7zoa/FYn/BcUyz4h2A6vt1lVC3U0Rv9DHo5OD4
1pjhFCRPpWhaUXm8R0E+jCMN9ZNQ8e1FiLJoKIxvC6F9+YgtpzaGoxDPWjOZvG5e
UxojyOQgjbW8VvoARm7dvzQknYR1T+8RnPQopIBlKqht4PBJbP0944ew80Ow6brT
OvXcFJV8G8TITCjI3N8GKHPj47v4ZBoDeaeQDC7KNXvMZQnjp5+ZMWqabgHq3OBK
JJaqrNLbCzIVPZEYb7c1WbDHR/MnleIySJvOyt2aX1p7p44xT13B0NPnDZYqvhWs
+PCFyDCp+QDW+7qKbInWeQZkF5CPP+vW7QpQ21DUrldfERceMc+zFLKHjyi59Wo0
DkOuEeBizRrQ8WicGgDDgJ4HzsK8vSceRdsb1mxlcl1ITAGXX1vPer+4rxZ7RcMo
h/nxCDUMSwkKEaXmYE0Hn8i5W2FUETqmlwC2wQVxOOtLjTEUkWGbZNP298YvykRl
wx5609dJRv2aCI5UgXHTq0fH7ThaidhjrreTeRzEtyabG2IJIkol9T43brU032Yn
kpiOMypnl7fdel7ToWmpDDoD/R+UrTvZXWZxAqdx0mSjuxtH2p/Jy0Og3HVdgaKo
axKZKeZTwMfxdJ8uSGyg11rBNcNeeMQOzDAJ24tvaLiGiMB9U4QshRXkdxuBNekP
8sw9u/qsUZ74C7bGwUfVjK9kZEWBV+bvBMQBXnv9qWiFu/38RRhsN7OL/9Q+IGde
5QoAhjJhtfGr511XLJctXrk4xpVGtxZN/l+8Qb66h5vOjL/P7TqpRbwRCaw6OiZO
RdCDpzMwgoxlsxqevl/SLQvRpByx37NRAF5eBkbfA61pcWlPeOUJH1OfnlZ3yBds
rwt1iojPtWnKIimg7boHJRPZLm0ijdzYIN/trcRns4MoiM71ftKJcGWHXpNNMosM
iDHkGX7D4TeenRC7TyXj1LRGLB2wPP4aKTJ0ODOJ/SI/OX3hX3qCU9SV5bkDHQFL
b+4X0H1551bz/fqi6MK8fnLq/0Pr2716h0dqfgU5JFV1SC15M1EHY1sLjMjfBX9L
q66EuqnmoQ+2AlIkNZkjaDgIbyh3zQpDUJKLxLXzG9icWEdesnRCIyuf6Y21o2DJ
RheY0yxGiFP1cr8VGNfZj+Ujfier+PnaLXiXxwyAiOGrTsAYVUTvLRgFSt4UX43G
FgoWawiF0tHZjSJsg9ImXcn6NMwwP1RFjQ9+sDEBjzsWxK6PkTLeGAjYcM0fd4aN
NsTvU2sBNEPfuAmt7lsB8o06C0VpWN+MqG5f/QMG8TojGQFrI3/Fs/h6sL6sSCkN
aGv0NATUB/uPu772x6vcMR5OOmBtmoQ9Qpz0b2bWDrq4nNOosCQU5cHOwuq+K+xb
4D1bDkniryHYfqYk6hIVWncUIJBq/gcjyO0hZi86pLRHRu0FKl9u6CWrDGKYmLLT
3+BKrx41c/XxXHoR4xi+9MzvLon01uYAvPA5D1zfCGtpJRn/mfhknSDAjJpBYqAA
kD2G/1cvZlrMZDzcAlevegkDqEnMfKFTn6TbRzTFJFOb5FC2FP0jdraFFpEa1iB8
vmSQNXfwGcMs3NFlbFjv42tFJuOLgyFKbw8NEP3mrbZL5VjPrHv5M40RepIoc2No
K9axIWB/LsTBOS4/Er6A8L65vctMapu0G3e/ExWgXcJvGdBn8WbiogP0IdatuBj5
T8HP0eXyOSK+ft1OuvP0V9/VoxU0oSbqmD10eqGVLZhVivpsw4SF2SWQDr0e/sV2
JRYxCmNM9IDmUuulaKU6UtLoqzIuoFU/HIUt+0ArCfT2UvgG9kRSMN8LyF5WMGcF
ErM11/3uwlne2WLh5S3h5NVuzDMPpQ4aLJf85WvZOKw0AEJYP3IYPgM/qWj4iRMw
dRDoa5zQLwPg/Ig1jUuynPRPPStrw0P7CkcbdJAwvYQTrP+Pb+38tlNGdImmiK45
ZlKKGK1OVB/S1vScSjq71ZzG2kao5l8U5uiQNyBmV3fJR0oBwjz9DcJanOBLDUK0
F0yGcXWFeqXewgSQCxB4+VCOt/n45U8/LhYv1TLia9+gfgU3gKDz2ZKjUfleg3np
4CIYwCgOxw7Qxra+VKpoIkA52qzz6BRGIGItZDhUhryr3K2JL/gWNCsua1HA/IEW
8MxXSrXqi+WW6BfSWhHSXEdDKPnd/r4krCIylElNF04GnAq6tESUet3EueUg5apJ
geznAMhECGQnT2Q5x92JRvjGi8NdrsCJ8xTU7fAjigOVtLuDzVjp0LzeBb2JNUAA
GhMvFnp1Gg2NhkRjJjBy6DnldJL5SNHZkYLZM7tmkFsMAp41ERAckl7ZAatJrB4v
DqvZqJTedVHmY7o4iUeptBRQyfyOs/O0J71mDPJGwURh6ZMngnJetgg2B9pAo+Sp
EJcNpFPOM2CZrMUqCF+dynqTWIXeeBQsPjEMA+YA0sAdkho+nQEb0FUXZ3VQowMS
FptXKGk45UzEoqKaZnKgqmtFSsb6mur1n1RFABe52davK9gtToFKrJ/RiTUQQ+cs
hVe6o4sMZHO4BD3dh/GIEJMHtVlFT0qgg7rHHplhJKtjbyhBFQuDq6LtZWDzT8VC
56JqAVndXIVbq4HWqye61eK19QUgp7QniGBeu7hk8tNWX1A9nZc+t/Avp/GIxi7S
UK5meL2bqcaOm4V3dN080d948ryvToUF6cABNj8ycjAyYfQLh5ZryArPaX4uxZi4
IAdxGNo/VB/A8g7rYrenoSGn2/ZV2S7J9Z4f+z/YlJCWmHyc1R8C13fEzCpDYUXe
s1gE9Ssh69yl3yu+f+ow4hcgi9CBg9AA748S/xpmTjARhgTLEcwVuvllzrIXUXNm
cyLskHc3p9bq83cudX1H65GmNkwrR9h0lHLISy6v9QcCLq4G7HfSKqe+U1d/ei4J
DoG5/FWJUsIx80fnp3RIzqArW1P7Q46hZSaiM1xxZryZz1kJHUAyrdsGNsZguYc3
zcb4GuNnzZUVRoDYpRkSaxaof3lr4FH+Ahn6FFpGZG3RYQGJvb+Tfoe+1+mUk9QG
l/X46dpNo8POo/w767yiM3Es/+GZz6/z4+y8btvEy2k9r1tQFRZYV9ZIpBKzxjlx
htFixTr3H+bh48BfnStgoYowqOK4EN4mcTeEOjsC4MWc6MhldVJ7bI4SxifztMw1
0xhPc7lLYCPpiSMfGhxgrLsOFmNScx1A8zZyTuCRK59UxtBjX84ebCry1nrlj4j2
YjbjAu9jAoFRe+XGnR2aTKksQmRFcrLk48PTeh+lj/BKb2Fe9Max5CCtCvuJC+6I
4Mews1Or4AlJCLhw6sueA66Il/5AbKsYrldSPOhiJfq+SqR3HUW8sEW9B6NAICmK
URCRMJ8LOtzqdcSQgJJgqcB3Kpyufxz904rqhXTp8gufbOzkNSKv0H48av/uUGhH
jctIfDdiDlZFRp5wkpf1YUM5j534Qm1IQoV1CA/NcW+BFlt55E/ojAcu4ApoMnqx
MgHzTthuzyOeb8Jn2fss6ogrETRXd9NDXoVUZ50X9620effd3vaE8UhShuTSf5s9
UHMU4QZNiyFVvL3kqVL/JBqBQA5Xai3mBcc4mSK2+L6YhbdeTLQzyVSlM0IOiZfI
xCSs/fRs04H5zUrlDzFJIItKpyDGyBkfocGxJEBU1Rc4ThQ8ZsXn9bSUK5DklDmJ
nbvN35FKEdCv/UYyQWWw+JMXu4QCDaHKRLIZfn4iyHbkPO7umDcvcQDeDAbLXwN1
IZIzMdZztqF1XH1NO03Y74aMTrNl9AWqXKhNFKzUPD5jHJ943a3YDNbONOh5+wji
ppWFDmDUuDoJNtpi1k79LiEDlEBAELxLXy8OmuPSk83kLXRW1JtETipFCAWCJB+j
t3vfAC4DAE7b2rEiHjdPtYKUfYWSWp/2NGAwgp1PkNyg12wsp7PjpQKbrhMj1StW
g6Cjhc9a9HSUHwbFrtCp9T0w86VnGBWaXFIHWYwmhUZhd13JKHOr51Q5CnS3SaO0
V/8UpNPRaMVPPYpOhITawjahOZ0Hduze67xEob0pTuqxplBXCF5dObr0pia4CveH
pzP/q76i3YjgV5GNf+BJn6wXyaimWZeMcMOEoso39lFTDrkmp+to8S4G+xnEC7TH
xqfeq/200MTUuRr9iBsVOQanNCyfgSdPUQu2qV24viA8oHRDc+EgDUmaU0RmP/y+
KVFtzGzlyXX/hLe9rAx7Rn3dNJuAMBWaqyGWkR3zJgw8Zdyj93IjSU3bugrjfWND
WQMrYvxE6W+CZwbZ457J6nYx8NZNFdHgeTkkR1+dbuJbmhxUzpg0qSsL282XZs2N
o+n2oMs7m6l86pNBHz+Sbs28+b10ZteezsYPC1o3D2ojzS6/JZnW1xeGct86w+6D
IJ83WPNMj58Fjf+Deqf+fKhxO1SYfgZBBIJ5cOTYsDVCWtV+JMOI1yAfiwYQgFHt
POBYnQGyzfttNPPvHnfldya3DWFzNlMnazSJhlCOdWeFFy1lMz1NRJEtzvQ5YQmM
IKPUNg97gnX2ZoI6dbMvrSTxIeDjxXdrF4dy4AAmjTH0LSo+b3UISd3LJVXhf6qd
KzJh1040xGL/jqJm3QokjAV0SFojUrNjnKK8ZaQdMTdvg2DoikOiHU9e5yBoujA+
IPYgOMBnQyLk64zainSSDhESvcYAEHMFZgjooMKlw5NSWkOf/WybNm/Nq7CsZYg3
igf2S84bmLAJvYggTKwovqriaBHt6f+NlDYIIWhujNtsMT2argF3H8Bi9Omn5Y4D
hrEIzQwIy2YjRvLMEamJ4BjvY/CcmUHlEWFUFHNb5X3FbeuJmj5gyhN0zYocgY6+
ZFyoCjEY9IfECccyyGsQOzXXYwGHzSFXR7au3dqDP2VaY3qKyyjDmDlobDcgaoEx
PHhGdsamzrjw5lv/9/Sapih0KdlIOSlh18f7YZSCwPxzhEbkuhkxBAvIMaodpOxJ
v1BPjcCpQTp4s/oHRh+E8PiBzGdNGdgKW9RceIWfp0PtCQD5CzcOusSf8Y4wZnR4
RVEniIGn9yIeuf/MKwttjxkt0cRBYte0uLIsMqTesPqg81uzfr0EERJZfsMzN8Fq
wqyivHr41Gbj02Jc6ehZkyEY4T5ObWGNkOP9UFMOhPTnYZSWc0SzmfGhRXdbD26Y
w3OS8O+B/4WuXne+vnJ+B7Ya86FLvpueyjvKSEuDN2TOiJNbN834PNKZdLWCbQuP
X57tfh+BfT14GN5MMRryaXszaeol3/gMrZ3fXhasYfYTP/HuMZQy4kj17VIZgYSn
vYqBsVJrbZRBhfbNoV4nP/uB3BmIe/GuHoCgchfIgzNaR/fBkAe9GY5EJ9Kcu7Iv
2PvY+dl8B/oVhQD3pNGhUAPN3BoZqhSvkYu5CsSNfJKuawtFrkfzSoYLnQQeyYxQ
A9h8DJgFexYcjBCU8aHShwIo/L6hTmhTYg0puiRBzifYZJ9qF2FKz/nIrqiJmvyg
W1nUzxC+/N/bTQSsyXuIDYhmudSggClPAnJMjOTyK0wifVRJO/dmUlYQTIHsBMJV
efDGF9sKBd3ygRf62wxiuqpea0ACHZzNmp04JttlTpKLP9IC4eYnEIQt0RfZUOWy
uksyrYvjCIHKPvHFMafEjcWzgOkm/j80fXm3vxYrjig0CbFJVjGfFuzyVP9NKFxv
M7tahlqq+Eip8gaMQvVuefU41CDrvU1JobAZgcBDiYU5u13joqjDlXPhhGl1bq+4
L+LGnlBZTGZmy85We40xY7fKk1JuNKJzvMDdnTCMfem9l6oRJDoLlbF8KgxBAsSj
otsPvPhvZdRlmbRjvutkQhc2dAvpu9TDM2nvwrUh9CPCR+cc2oNnyOc43W6Mr3B4
LWh80k3IE+KxXnkSFP9msSz6yArgbykJaR3bd3kSjHfUd+AkX+7eGOFUx4hbCQru
xMH7aUqQpm1JUoyLb3z0dK1Vj0bkhaP6fE8WXRhopJ6ioR5SeRZmVO4OWeO3SsAN
VPO//HDrcxUBwnSer/TkTFt3UnHH3eQ+rxRmeVjFY6/ofom4F4Mz36lvCNA6qfGv
+swl9socrpEnAR5no0w/sD/dkoBMU/Uep5Zg0WUH6lLEwRxD4r7abfGHBhdpPQ8z
gREDKs8EP+U/NVgz7qD+JKbuTyrOggPI4TivHXG3CwE/2x/yoTbmEWsoGBnyDDTR
Vh4d/jbxxoL0djFnaGVVxQPwW73CtAYfbg5adgDNmZ33P8SANgfUdhrcnCkgQ2yu
RUwuMPA2/Bm3sQoWilUfpSY8NHVPmY6mLffNOZtE31gBa8z/oYV6qMfn1/vJ34kR
E4vhyPft6zWfQC0KPuksJOZIzLauWicZrBqEMrYorcGC2lo+2JlG2QT7k/e7EdJJ
QsHavNveBNsJdNcjSP/FmZXUgQaiTqHSzrpFrmwV1c9ed3a/xKkrqXkz8DjJHmA3
tOvygrSl8kz8r97d/ojVMACh7OCSEag9cmABxeEanJoFOnXrKkxTMATEtAjxzr7l
wNd88XAM+EJqID2cfmRmfSLmLPyi6TwuDFz4LAK0ek0DRuh9DrwpktZ8KinRKok1
WqZCSc7sXu6Yg5/zReUAbNMnOOphq/zhhq0K4fMBGRgf/xhOHCJ7RfCUkX6s06yQ
wSN+7efRtZl1o22KkekzRLVzRlAfPPSNnFiKohX7aOdilokYYWBr+FmmN2EbrXQB
0rPi/vD8ptGXPzZ1eb2nzEKRhCXXYR9gDG2bKmky2zEsSZiT8VZhZNaL0qilOp9e
Cx19qH/fM7wp/G4r5zY45gm1VKV5plJSfAhMKYevlGE2F2z9siKnjgLVqVQrtwN+
bynvHs+4SoyGIUGxW0+hOpnQPMMck/2xNovO6C2eMw0ezLfFIWKhj8y1BJD/lMG7
OfuT3E4HFjl1V2roIirlnkKzZPwsM8K5yUL7zyQFQxxQluUhw6ZnSV7MmEF5FUCM
lDbXoUr95UwjIE93wZwqnKgHvNJPxsYpHH/2dN0JIiinmp9IuWq1oWecpeusU1yj
ZWTIx/+tsy5ilDhsJDar3xn8+hudSHqFbrLrfd84NrAXIkEwVtS2cuTfNDHXQkvX
4YGah5PFnNTjXy5YXDUlXahDKuQmYQDBIDJkROPRTMSp2Rxe0q7ySeqAWLANzswm
j4X82NZxkvOsIQqY8DqNOhVFgYoD0s5pbZsLv9tfRi3knor3vAhs3JvBG2lE46hB
dop7zrkXQQa7YNsw7t2IgdJKWIeHS177ombC3mot5BIGPNGlxpouSrTh2FkuaLwx
mYwb004SKXRax+bKoWXRhW1IP4gD0H1Mldgx7nO4hZfTRzHOZ+Rzr8hinu8ymYXV
BsbSYqaItq1EHfg1yzeMTSG9/b9m2yVCSHzIGa5uJqSc+3037CHCdVP5b+SlzyN7
B2gFp84MHonNioGdwPE/b7CjYbmdARyQioYIDVjMY18t6929Tls+mv6aiyLK2H40
nSDu0eoB+Bd2rl0Vm1f5vipi0KPcsOlsncEDP65ZF0QLSuvNPQXIzv0pr/a7RR5A
HAdjnPOG+TrrtOtgLDmiFORfMjl6j7cY0304sFcxVhL0WLTsBSV+V8Kzte7grQT4
7h2XfCOniYA0cSGpUe2BBjA8T3l9ZkbzIZOQie7KxkDbLxvmIIQ+iCt7m3aNapVV
G+VW6wuUM9ajzMTvoO7lX9l9mF7BCp5nnSpIxOlSKVGg64EjMHoLluktoi2t2Nwl
RfHiw7VlzXtcHS/S8IR+UKHdyEccDTKKjYY00yoDUEU/BkK7kPy/8PCpWJmqFB3D
qT279gd9fZQZVE6Q0+8a/zwlCnZtmHYCtfZVC17nJ+9oFj+hWadd9irQDLR6KbLi
n0oczF6+FDICZ0H0lHdM4T9MDje3pQWSUOZ/PbzEziRE3wG1GW1djN9+RXsyX4TA
oPSIdicJaMDRMpVj2O4m9yuy5RDkNEsbfP2r4CcR3G0/XcIYXNeYN/0crK1RXAwr
uo+tjTF5q4vC1du+AqS+biygzduKs2PNWIXjxTuxMLl9zsb6k43GtzNaDI9/Ycea
JB2n2TGAB79KddEp9HEa2JSmTiMfJe/PUKN+jBkz2QAGtJzSN7H2S6n85hUdUvpe
PN5Bv1NwsY5lY7tdnsksf2BXQP5EeThwQkKb1nraeU7uHLEjKj2EgJh2afVZpn3C
fDsPdQgeDmQQf24olbmm8Iw+EuGo93HZrxbGznpKe8MTbl1jV3Ey0ayiBdEOOrDh
l8sdkD/yBYOg7IE/BHjcdT0Z4OQjb1KzU7L+/JGMbECfmLHMJqSg2Tf/1wUO7D35
9ldLiKN15NmgzNXIvUiqGlDjzMBt2FNugTEW/3TgrX6YOW97UK7ZOheLN4VJzSZa
ovAUUTVxIaTAjU8xJZ3IHvxGotxU3r2s0IjofuJZ19SZl8aUCx3gstg+4tGNiD7S
Ch5HHKJmYdJfWlFahyr5ZkrS9Vud04/rVg4H/S/MM+wg6mqBugVkhnCFuhvzqKni
/CB6KqTJ67Jh56bcN2BS3UvwwPz0McQtNEmj4b8KCDMw0B98BK8dNo6qLlphR33m
MmiTJuCNEmlkgf18RnhUnYlxJvdPaWtYaOJgyTN4j5h/lndNhgKS1s6BOL2br+ip
muY7mh3oZk/ULNYFSaIWKc6WS98sNKpuloe3d5XbcAhXUypPS4AcYc9qo8aPBPW5
xUdHCh3gxX+ClAab7dKYXsXf9DSpcJPQAjOLgtE7L/G1RANF69UoD6h+n3N5D8ac
QrbC8IP/XWZUfO0VeUP25vwq3//dLQhi3kYJdw3p70shO4fyg7Dd1wXW/AXSkn+o
5fZxhGbDzv+93MndCdTo+7ARwYbwQEOR8bwEY+IwWxA5QICAnTRpX4mkOMNQ+07C
5j/H0M5FdS0bRCjrXZCMPqWy/FawDl6BMKWBL6rtHxMj2pDx2yb7XNZGq00VXTk5
aFAqzGNK+AfolZ4+6QksH3e+1BONpYNNV3uKq/kODVWv0i/2W53JUFNRJdIxOf4o
L88eVFfRSlkZWAbm/F3OVEh0Xau0L55D28PQ8Q8WZSQRoxHKOl61FIePuvxl3Lo1
QgEL4tjdNR4RfG/T+f1dlDUILA83pxsNXnrmiM/yCtX4ixMtWJYMVMZnqeHZ/eKZ
tIPnIjJKHa6UzCL1XZu6X32fJ5Vcl+HawMiNqAJigkcqXfVKgAWPIrSYkDy1Cxd1
kfdrfMGGsgQaATPJj2XwILesm3Am1UzKBkgDULlHQ0Z1wuWj3WPDVNBJiFdsS5F/
19lnYsJOnGknfGiENGeQTu3jT0Z+WJ5N/viiLATsUPR1Qd4ln7PeU7KcZrPY/jdz
RWEhWyOyED7Bo1p7QP3iaujVefx+gbtrJ1UohVcrEM2Jg9mNiXHrDeO23hJUBq8e
7XIX/GWk23IW7soazrWklYKk7KxLlhDeFDqd9m0etzgsLa5pcGIDKgS+/lgRnwTG
Adu7qous6i0sP+I3Jl7bobzS+s3wxVccouLeB6pcKJuPT+e/+vGb7EjhRyjoeEwa
TUwHefppTaCLDHFN6eORebbOlP/pDcK9pEZ+a5iZ+zBTF1uAs+jbacfy/XM7/nct
4d9RadrkrFVfXDepXAofQOMdUnA751bf+A+eRQ4tF6bURhHXnzCJaJ2egx4AxLrZ
l5OJLUqid963kJs3bDyK/xnYkFopb0YFrQqN6Yh3IAYOBmbUQY1+yvFQou9LOXpO
McWBxXfvyLA02kUSwv2aIzIconPIEQHX+ELx4kPPmsy5sp2S8NPxV/EnuIUCegGD
imDeE+l52VqXnnsdCk4hUN01pgXLd+xmqDiplKLUnjf62LhXZR4Yos+XwXhqqTi5
S7nijTdPePBfO6L5+rPKvPAAOYzghPH/J6b+PzTw1mA56h7pyWyZ7fNtByHSDpgO
6RAsO+kZvNkRElOvxSCtbtVNg5BAWvlHza1op6Gn5F2C9oW/E90EMZrIs2gLwAOe
vriFhM3C31XHBiexxeJcWmsrpjir07GBsAkst98/K2CD3HedKcfOPh9ZE15wNe/s
6048+jgal+HB0rGSh1YpDYTvmTUxpsIIbWQK7sdsAQgNUawB3HSwRwz6mK2aW4Jm
Oe9sLWKiAcA5+f+3BwIv3seZL2aPaNiOl2+IB5xlZyBmsF8EqRELHAOFWBCgUEGR
ATcZ0+AS5BxyrQza92c6wx/SpaRVCTMLb96/NOoX+kXEMeq+uYKLufRWiugGG6n0
+vZ7OjIJNvnNacoKAPgVTPI1ubyAYJ1IUZQQZLW/0wqqfd+rDYSpWxI7wZOf43MW
6qdWFhT++DTfX7dyuRPhOFhkncoFyGcbG4oBY9XiTV4rG5r+PkPXH9D/TWtRIcYB
vQ2q+InaZfJWJO8Efd2Y635pKW5D/yor1XtHQlIYUTB8b0xDPlNjuKQSv61p7E0S
2Q1vlakJV2YWNoCgjPpmTTc6+ZN1U8rR/7eV4HwpdlEL/F8uW+U8NTwVuKiMKSSv
zqIwj3d2AGozuxHIpigK9dEXPeC3dzyk/y9My0Q5U7LeOY7gi/l7SMKmya/CXJAn
vlF9pJV/+qCGYzItOavv5akOrhc1tw1IOOSCiw7le826BbkVdewgvTGHYppY4dwi
mLfzxP4NpJDRbKB1nNKiPRLfleoiZcmd/zsLajuWsruyAJ4oyDQbdOsa0+yb04m1
vicqNgEB1ZAF1tTex1bxm1r/SSAE5fow/VjN6MpCoCILq2B3jA9F04U9ijc3EXHj
8CEhqwtVqf9usKJufo2Yx1cUWWT8WS5CNL4VPvv0HLJPqS16U5/fgOvk0tgNIY+G
u+WcLf2QVXVvPPuuwM9BRyM3ascoD7vcuztmfmfO6bg25lVy4v2FpcTkNRoQ1X8l
IzG50phxY/sSp0siV3iOP78oxE2XfvPq9oX1J0S3HP5WwimZzqku/Dg6MmINtCCW
wdZaP2eB3aO8iamg4LwWQsVunBRBGMVM+ETzTBpIEoYPNzgnO8cTOKnRiC1B825Q
Csmn7MpB2kgAeveAZVOhblTEIiDvyPrcSxEF4U40pJ2x/ZjWnrkn3v79LIiGqAn2
ZswWk7Cv60MFPle8OE5kihJ3mTP7dY6mdQ61wdN9qYgW0DsfqDJPEqkyktz071Yz
18+690u1fbYzDU2O7tzbs3BIvqMz60eCTdGU1m4Fdq2RoHdMTdhY/zmDtWqJh+t8
GqD7Ci2smieC6e6XCh4HMeb7sDlXJzqf1Hd3aY6IL16cz2aBrVMdNeNfxngBmSD5
GAPcyicuagE6+Rzqdx/L53sPM2xODXlWbrnIOz3EHSbbBTjqcxzUdrYk+AvlUPV+
M3G1cYUEI2w/gqxwx5PpnjqFW53gZHteBuSTVzftel5kbYnMs4bH4B2/Vtsyt01N
PEg/vZwmyTYsZ2nmlOqCRUqJ9+WNe7W8K4aYcbP2NBHAb+R0xlVeHpJpxZoo60qJ
waavWyr+FRujegYngl16XXnYq+I55nLk2smNLEhLx9k+uiqWOtQZDpjCv6h2q/gf
4RakMWFUybyO2Y6oiWJgoYVKUBe4vN7R36RCHW6TybsieirenqLYJPZ9L4LVq2BE
+Orc6PmHz76oTFBF3wN1AWEGPiT/kfRnXfW9rrhvOMjflv18/X4ZSblFbalBv1oA
Kho3sNUvB0rVABXq8R9UYYpZkZPwqdaTHkUxP6PwyKgo03LpJ+f3MZwlOjcZqRQx
xgdC6PNYlqN3DDMNkqGkTjQkiRltcG8QLDiEADjwF+Z4Hy4mxNeMkv/t1PKL83Ss
5BPbwa3JjWu4TXrpBQUHcE+2qdQpzB0MgyLULw9o7Z0aUso4AZ9/sX993i3zU/RF
PVdgG5EvemO4EmFcSsdbz+09z9EvNFUwBg6cmLN2jMaSWsMjPwlBclCRZ85T5Q+C
fIeO4Cjj0YssnLGlyvXvT88hfFcw0AIzjt3k+ZZXtH+ZWZ9Uj2ZUEwH8gqLsvKb1
rc/ExHF1k0C0Of6ddxFFn8bnkbPnAKh2uUU5RbVfqcfKAAbzIRkXR/C4yheUpmGs
Y0BjVFzyH7VO8MpycibBsMPOYFbvpulWAqkDPqFPSQ6oniqX1pWShN2gMXWWjNFQ
pA57yXGcffyYiJ1PNK+m+W0nuvnoJYeoBN6Vwn99M0o3o6mBJYyQKw+LFyw7uYtq
je1klq6B2MYKlSonM4E2j6Mx4nTA9KD3T8J0g16+t0SaI5d91+oTIKJaoyhIDYOa
SUoqbc98JYyHqCv3NJaY8UDptwnxFv9LcDfrUbpLalXTotthmBgPYaZMgjKYSMd3
iJeQWeCqKd7FaBg9Pqm380E5uEKnxkYY4XRHy4ZWlI12XDdzlD7u3fj/od117rTP
ZA9Dyn1qB2ptdsIJQAVFmipHBypFEVb7SPfsZOiGiIjRzzZoZS/zxypuolkbd3yx
QDx8dtzzdnaI+D6u/aFJwF8eyDRy6Nnj5xi1zR+rXS0EcEhCVQVs5xQMIL51GSQ4
aftK5dvjf2owB2yMRsFQD364otZ2kzxG/vDGKFgIJbmZLwL+gsFKtmeEhaefcSeK
xVLRfBc2WRxk+FClR3guXmlt57K4tTWBwWbL8WuwwU0r1I2Dt1IlDSUA4B5IHP1n
FVDpDDSDfJrs8MtvCy9vcEH9+UZLXLcV2HfO7H3KlwFBnQBjk+Gs+dyTRNj3uMKT
2+LtmS+CR623d9Uky4QNZIqznUQ+3npN/f1xQR+XyYunSfPRSdR592LyoUtCjm//
7aVmkoNmzd77P4OzYLRUiaPjLsrooV1/0H3BRVBFUKXXanBwh7HpiPiZ4N9BlDZX
lwKHc/pcEY6D7tJC4XQ2hrk1DZlsSx0hRlytvbaGD/GIKnlWSPKjfYsDC+8s4c8q
J2LJLfKqNRlScTF+U+YhV8zB6RJdsKCNvDCHt5Dc/S/RC/k7FoauGKGgb0x88HAL
6hBCUkBvqg2nGVsqL+jX3dk7qj1tGYmXAxyli+5iVeUgKpS9cRRaQK/uaoxv7yIg
dDuztnjhKPJdkuYBiKw+WGO2DH/g6Q7oKhcwbR5LG+cUgRUqqjJzsp7FmxJuulVY
UcaawmqSsp0ljcaQJw8W5LHRfAeA7rrQysZQMkN4w9NZdoybIYEpJqUozzl5A5ZO
f3lGoHKdL9+9bVihau4hVzkT0jzBmXFuyQdvuKu4q/Mv91g//GAqQ/4nL6G3H241
11suheaGVA4/Euq/zn76cKLc6QcNBQQ1c+oA3bKeJ7mJ5B2jlSWlPRs4hGJ8TJCT
kkW28Nm6AmBtYtX2KartCQO+EM4RWqwV1F9MxU5orKP3lBxOjOSaSHAjHgnvNYY5
UoxWBP/Kk9Hzpjylw80DCjBN/WYMv3HjtHPog1yCqS3zfVIFCmQ/dRx6hDjSBUDW
k1poMjn1RQ2ZUKWd+/DJ2Ip8vIVb4wtBqg0Re01zMYQ3af/CV/PG4Q92hjNYtdoq
tri/b+mBB3gMjMaLs3s9BKjrdLyxww1RIuKHVSPHgy7uW6ZYo6jy1A+ei90bHlz8
1Am2f42DrZFEg4/TfQkkA+t9uaKLngQtwpOBH3v5zxDWGXlw3aMDUj/YfnsshRPB
sY+N5/p060wRuz6n1jMAdK2ZCbHNEx1yMa7gZVSV+H2SY1qaw7Kj1IsRzwZq6Mj1
6icHa5Sx6EyJZtRiEnUBYs+4QMC0/ojIcKPOFsGVfqoj0CBiDAPlspFnREoZkiva
31DPxi7BhmZsV0G1PoSutZT21hX5WN0cSjN67LdqMK/j8OvWC1nKxBYJQ5tzWLI/
PtN818oSA6dqsf3RAgZ8KnCIErGOYtvqeP+YHx1HUMW2ug1wefikFGO9g33wUan/
fli3gq2FT9nOMdPhEvKu5fS8pLFoZTHystJG/M4/fjnodjcg2gAHb0UUiz9kS5+o
K0NbEoWATlxHqQn+mzvdpSDPSqOCXYvK6YReUp1G/FCgzxIabS3aeCUDiRDfzTk+
pZh1qsksh1CttWgbFm+C229kvNJjwP6oiGiwMQ5CyVsjA7Ircym2EwZ4hZzjuH59
0/q+2eFDr5hloaenVhhCUr8pvgXEliddE9kV72mV/9qPb2AbtvUWaD+FJMCYUBTd
lkgusdDeW31dac+0bYLtfJ5Fh+RT2OPB8iAJ9l55+w9eZ88hoUpIxvF0+YICdXGO
v+5LJmujTf6ygSPvCddA+Agw6Kc7nomFEcyQByPF7JpJ6oLo5MFkY0qwlsJBXCKI
sNtDAd2eoXeeHcOgu22VkSCspPIPYrUxJOW/Nk1HVpYv812MErNIdqjI+XlC6hTO
MJ/PdxI726NgXMXu4iU7JtwJPg+FNMnBJwhCmMeRWEHsrISMhRM2nd4fPsLb2n4R
rTeqDElPkGlDFn9rRGAjdh8X/LD04mtzDX3s3h6y7zuHHiCZrMmIxAdkzZykM7xy
xZBkwtOEpc3GRgFlU9C/8s0q8AYXtdHFBXMwiti1e+BoqAVEo+w4euyub7eqqjnP
48dlrxz2w6zFozH5qUdYtf07lDGBjKxPGsTvmfa/fyzrWVExqzm1KGNm91DYwlzW
26qgBHcGWjbSN8vWQESFSF14AR4x4RJjDeaO/FBrw5FUi6Zpt/PynLx9M/Eg/iA7
s6wzaBZ0LnkBjuMxxCAggqnE17uZJDSYoco4S+lJvS4+b047mWo+YnTIdPF9HKLy
gDGCiRhlMTXnApHxFBBl6R3tMTzmzVyDFa+X9Lp+rkfd2qMugLfxwZCAzrsMoYXR
gBBO/Ghn/qaOHIn+kaU2qtm1RG8G7w33bKgHducYc2TckMmA3YD6KuagQS1B5xH7
Hv6ZwgghCVw0NkrnFvUnhkjV5xAVjZ+fZz/46+Jmpeyb89H+1PZkSF8UjdpA8dFD
P+B6br0qknpJrHJgE3U6xo6QnP7/d3odDTD8AFS85nabwAJrp0W0/H5btOA+zRVg
i/AsTKeeunUS/MCQpwOx04FCD9JXKzVQFfU3s0IejoHYByywKjgtW0DUGeAtPdDf
rQJRJ2pBwjiN6q7M/joz16LFj4eZeqM6pbbQmwPIULZjs5lmCaigvyl8jKa6oIsS
XXU6tDGI4bUnybuS8Stcq4eDHuBabhPOdkGeVsKM2vcS4CJxYBiI4oC4miDPceHZ
Ieg90rEzLuH9w3B/QjVWuMMQGG3uwi6acWqx+fRvlwRKDPzMT6rNEI2jZzhemIPi
Sw/cpbEf3BZKRNWzKYQT3+0hFW6f4420Jfkhxq/fqNO1hVTb9tHo3vQnxiz7yJnL
fDFc0+bLRqnxgBlBqxYIrfuscwcHtuCRinU+hNTH/2Sx0iefW0RUBdD2hXpc43mo
l85u6Kd0RMRb1o9DlnmjkTGZrqeWU6HHGshBWdRAb3cobksOY3krxPz49YTVzLkw
9d7KmN96BzMYa6JnTSffBme1OptBhD/drLLVRVaJi3IZIf/QE2UnuW7Wu64LuxMO
twhEOGGp1MhPfTmpK2St0Fxkrn6JJd1fRtVuW1UvejdpEnlSVGvucy2VSuy5TYV0
ONzrj2HNp6YAXkxuShYO0RtzBz9pKct+c7wyS2JVykx92+Pg7PLbxC7oXCLOMvJY
KhGdnqyDOGV1zIx/wCNdsLxqyQSj3jo5dIoxW+Xgu61jrTcBf45Hgoy3unzTI9wS
ufjtUALo/Z4RSKMkWORqoxgzYsUJmU2UBFLOE1NVCLFVrn8+ZmaXdrcz9KtMJ93w
fe1ytAOyO8f39jAW9bXZc+7+C7ZqWPQo+VuQ0Xoa60eH/VnmXNJKj3SS8ksd0paA
N1QUTJ7awlZYniTk+ISu7LFbrpdhXjzSN/F0VISk1wHnmxZ0wIg91HwGHty2BQnX
fAErdfwzlui39fwddV3pY30Mzo7/QrjFo8gE5s3/VDB74+RBMa3DUTLgZua1ONup
ddM9LuLnHZWD2RW0HnZBj/UEgGA2q5iEtHO3/ckul+TNY9nEW56dJbiiuDxqDuWO
8MxAVOk7z6oNBEoMdwSVnmeIHhky506chpWvCZImshv40A88XKAl6jUaQZ4liXOj
tMILGfSCc3YULgQG7+bnuU1Wi+yYgqTiGI8YbLnT1pvHGRFoMlkqzaJk9OmyjcsJ
vk1NF8BA2GpcyrOsxtINMTuBjWDmmSGQk4cPa8OH/dhUeHPVHSucaAmeDn6nMkMl
4zojhO2bV0dDY72RlnOA1ncfW0tdEMsNNM0vgflHtETdbcWPFbimKKCf5RKR4YPE
YwDBVZqn6UsSqLOJzVXZkZCC/5/y4eJVC/0cKeUbWmYtimk0Xl78P8O1A4B9HjdP
1JzlGNCfjmWKQLwfVr9dlEmfvF/6pBWLNwYvxqiUKqYtQgiaXNOgfc1wX9sCZFjB
YDZmlg0gFt5TxbI+FCVA6sveGAPpE6qimYf+xyONA1COICwQCigxZymd6yCpe45R
wRIzno4QSM5OD+6MTKKfGEZt+6HkkV7X+Bd1kbsJALCOFRbZQuTo24ARFPUlFzFs
QTRujQPdcjrag+CLl0Lw4yiV5zNfcbQZQjVBp9hpnvCKRqfibCgxk+vmNzQrcxMq
yrlhpcrJSV0hl3lv2v1qntQgXIiGe2mQNbumieoC3cNZO2Z1ZZEMrQODgtec/u7g
y89f9YERWwvIA37qERTPqoemzWghUublraEN9LjUD4M6yp+kbOuBqr064GEsj1TS
qRwfwt7/9WHhSG5TsEOWLEoTKLb72rUAWtWhvsT4EfeZTNjYNzTccONyZwkfZE94
BS/IHnDkXCrYA0yAZbbbgmQ1jCauU77IkBcaYPNGnuoMWmeEHwZ1qIBORC3ykQF4
9uG5xUbX1FH7NUS5ACASky74XflPs5zTMRi2h6GN2/lDZcu59uUJgfmNCR6ZRgug
m3DGBTdSV2FmM3VGmyPpCji6lk2g5W+6EypqcUL7tS7fLIIJg7bALkNBtGsrbnFE
yJeW/RJmrScD+YEGP6uFA1Pmu9xi5PC+7/LDGtsk89Te1KdKll4kozIYqLFBTvjU
r09CRv0tmU7XUg47UOxE+vxQPMPCH16GjMnKd7/Hu4t4Ka6OUNarNNbzCphyVqIt
Fz2HyizvO5eMyfeV/pHi5qvxYKC/ZWVOLSa0eA+9ppFVydB3g2VE7CFTexgHq+Ag
wHvetO95qW5y1iXBPbewTpYV6UkevIzZTEen1urGOdj36wEQIySQXtUwYoIKGw7n
O/rfRBzaX13VS9s6sh2lcu12mduZUqaf8BhAD5/4rbfH3nyq/sC2d/gNB3XJjRrJ
TO8/wrKur3HLQs2J1/Cn8FZAHxkNLhoFL50gQRLmMBE3mzcuYYUHDq6/RkwiOsKD
ZqCttVr1iIsBUAl23upcYDcgCoE1XDIO3fCnl9vPBsz5URaXvDTP+hALvu+jV7UR
T0r+7gecE4n+DFN9q1kdXWQpXe/uOKBhr/xVviqkCpxgwC0RV19VOcnBV7rwrS7M
dMW3PoCoqqCPHSHbt1eh3R7Zrqlcq7Z4Kt3C01NWklhO3NMLKN6eKoMk0SQDvHLG
BEnPOFNa3ZUjueKTYf7cZF/egc2cW/asbrn8LkcIDtj7b4ZS9Sbf33PvrID8bTq6
e1XNWyjAAPJd4soRVOscTQPv3OQyU5B4gmNPA813gmmb1hollUNw2cC09x5niwNP
6ySddFWDvWnQ54JmKikNNg7CrjhW3VRWczxlhbNjeCyoNZpwNKyAzB06cHdj04lJ
yLbCRBpjAKtqeKgLSXHKhhstKWKPT9ExtGSmTqFLS9k8QpLz5WAJqM1Fqk4w6a7T
qqWCu5o62w5HQQgMZwutnxnzAgBpnj0YymfRQ9hYsOKLcctIB7OgBlKjKdj1F8q3
QiFwCNvJWUlk8j86Ox3/m17p7/SKm6UGNvu2orqqXpGPBLlsbCAMWUkzHtd6bbZ4
bzTRDv9diD0vM2zxrwgy1djdUBWLgAwxDqk3j3yah/HcUa+GM73XIQTbr9LRu6WU
vZZGhl8qqE5BqLRbLVKAfydtGDqYIxLz4rV7rxMzymXFpYPWvo+M/TaNGIkWW9c4
wSj67Ej/wXTrQ3WtDviYwdXi+xYuHVb9vBLgw7JuKroF59Cu8SqucxtFHp9EitE+
UN0Qaz7Wb3hN0wvsO2iCXr7VfKnts5OOgeW5D2s1WEsyjrEa8zglsMFDEwkotb33
XX+kXwbc3Jt6UQrglf7WSjKaeuAHsWC+VhuJCVmCpcPyAfv1OHM6K/EZeyObSgU5
UrJbnmi+1zgOJPvijRfN71Nom/Yr5WisyoZOvKpT31bQM9ph5Oi2mN4AJ04w9hLg
J/eKsZQCxcYGbE+PH0jc3i1RP8FZxsWbShhiBSeXmbmrCU6MY0XYp9+QHVBKvUFE
LysfGA8zNSCfHl5d5GJsgpyj/Kc2LFR4RMKmJcRjuav3BZXRNMttcENA94LEqA/E
k6JcPP8Y1Y/2pWg2F4Bzukcyio/CvnzktHnRZ+suXkftI7nxYRDN+emE/xPHlN4N
nadRrepOyZ2CoijrNVBLVyMv373pG73j16NTi1SZtcX4tz7u4yVBLYdtt4dcY1O0
f4Pk6+z/e62rB8mdHDBFwtH+RenSjnj8TjHFu94F7cWZbsmFlT5MB7k3XeoZC3Ut
1dipjm3Ca0KYJXS13wV6mshgGyVWmW56sN5V7kRQ8BqUnVGDTIkEOjjCglquPd+D
F3J0g2wFcN/OHWsaI+knLIXuRyiOoAhMHy8lyDPq6+mLueq4vvvJjj/ddbzVVOHp
3StdvhGUONGlgDsWPD9ZEpROocNUfCg1/LmlEpx0QO91F5k7UhYKG2Fkm2nE+/MV
QrvxExeG3f8St9n5CejuDqhR9E23SjMt7Jgs4Dd5azXYZFa/saMIUt0mVFYRPWZE
h9iW3FCWpY3mGt7uRW96HKMIjwUOBjWpLh6UNbHCjwLuEkLBxDac+5qMvfC5x9dm
Fb12OAf5gB+Cqwa+f8v70S0y7syZk1lNG8IyXPiIV7hGDP2rQK+78HGt5y/mN7hD
AuTj6jLOZ0Lj03zQLk7z2YwIOWjriXUm2tASJnGIlf0hJbVcUlvTzYba1I/FHK5/
jocVofdS+Z9vDi8feM/Rnr0eXRDjilBRblm6ALiqsM3VSAHNwXSR3lpptjYbzbO+
p8n0QrR5/bZUktI+6TTkHDWwX2Qyii+FqMUTygkAK6TtyMM9JpQD4mD9UJnAf8ui
3iQzc52LeGhjPH9lMLgdsVBGkDQ6nn9eOThYSwfVJOMSsszxLrGWaE2U27Fy7oM1
8uGCKnB/0cre+avTnfHVJ7wlEdEphTZNKMJAEMfZ5eQkGi0ZKoV5aqPi73L1sa+d
jqgQw70IbvIrs7R1jDn0iJRFjyi+ILFnMpBJJcvtw+yC65qw7nBsss9xNzsfreXv
Jf74ciwg9x6zXnzW/MNCGe/29F3IwkcT6C6bp7bKz6ng8AcsRWmEqlluATQ6e1pg
kZxjgSaakzB8WlLhU/FIGQsk6fCCiCZ+oqpjDJQHg0nwfq8ohIHqC+gHfpff4scn
PzXuRDuvn0JnX11PtM5b5NnuabChbe6E6nJW1PWHp5tCNLEEUWGXrJG2Ibv3ft7Q
b7HcJDsE2kmVhhiDHmQl2aQPF51EI+6G0NP2xtttX9xGNWTLb/otCrwtFXS1enis
3it1UYSiOPAoGXSWMelHO78+xFA4AS3zLLDRGcVM5lIWvTdRU+rSCXkgWiQI3hjP
x2ewd7drD4pP9vQvuQo4/VXcDtAY/MQHF9mZIWupVuCQukq5YSdIdeTXcDbpL178
3w7wNF0khY3uI6ta6mSPINhxkna/u1zLtd6LKB9pYkF5D1/YF7bkQ9NvS/haISsc
cl7jsTcLtSNVxh27BIJtaq9Wiw0q9bUHA9OuDZvFe4xxF5FX95Eep2Mze+YPMOzt
YA1kvNB0wH7z2OrIMGlhoZqtVb+7YUyBHNfns2ABBRQ5NqmAsrvrniik8buRTs++
on83I7Ds8EjnWQz+trdcCbfZvbsc7I7EPd1m3HupLURgdnxOBMNr/Wa3DDwXBCLg
DTVGuaUxA1aB/g8y/IEuc1gUBsEI+5Xpg805iBhjnlRDE8QQHRyMoFWl+NrW8BnK
0G4Mpjc2uwTbFHVucTUCeurza8n24zBML9rC64Wm/02wnAC3llLhsRs9+zudXUc9
VO1jPKk0TuSI/nTMuCYeHf1+LkM6SO7zC8+9prlO30rQ6rW7NFkSWo6QsGvBJFGW
uID53lMFi0y60tX3UF31zwXg+r9CFwoRjkqQ8Rj/dU4DVqi/daRm0VFbprSDjjQx
UW23iaik++ToH3GFN91dhBvxI4C6Av8zN2KSwDE5UJsyl0rs8bD+tlwkTHtM1sg4
nvOC0q3HJasFVpLHFJpDNpt0gg7hQtTWRrxTcttJp9op3Hgxos93nfciNbdvoFVZ
n8FIviH96iJrQFNupwUMKYXRPo+/XGUCF5j5L6TTICUev4Z4G7wVbPinZmhL4VPy
FiYUkCGffX5UaNkXYFbhAZJD34UAnE1CmXl8TZXks0YuGijWbRce8Y3YTiaB0diC
32G9Fpb4WpdltbKQrPdSW+eOxW6BbL2dhXCvg7H9Cl9+EeSWUaICwQLo0dWJWGgp
ExTFEcDwE5WA48dm4kAeKf+gnlmauQ8a9mWkKtw2htj5FbHHCq+50d67UxRC428V
CFwgbnA0BREWNROAZr1yeZwPqy3ELItmVYI5oDtmUYAV2gjopgaKK0zv1VEO5WW7
heOQTjUeOuRIU7WatIiw4lXaTDytkwDxfHXjU2qAEZvavn/jSBDkERAcw6rOmymO
lkG538TDVWbXYoeSiw8JPgghDvzlagwEMstSyHaXf+iIofdro6Fdxwt/S/8RZND2
kkaUNaTIHtsWmaaX6x/1MDYf4i3JCUwbHIO22VEyCWeYx2BdbTNxBLWAZnSnsDXC
+5vee0+38gbDQJfvfKs5DtPM7qhBx0Fvp06WENc3Ju6MtLd5M9jwFMnpR0SvYPnf
oQehYpPZheCnZTVudkbrPX9p6foE6+Nt1+Z5PTk5wq9x1bDNXy5rjizyBRtSaH0g
7IdTfZ3dO04YcJABzA3mZqK7zGRqQvi1tgtggDNSs7JoY09j7/BQGrasy1WL+6Is
vFNq5cP0/F0ZRTqhJcGvgqDIbY4NxQ7ECUrUfcwlGwrGIK6mhDXvTrEXJlznF3vL
Qs5XTCeAq83u5bcglnMCpSj4/HJ0laOds123Pt4hZq5d3GkN/yrFnBdu7k8j7AnB
U7Y8RdxcPTjhthxRx2AditC/jIwIJvCA2cSHGN4bJjwtyW/qIbBX+V04bgLDpNTh
uYqPbHyalF/TtmENe7BFYbMygTDJxFzlRyJTbkB+8lyaIxZ3Bn7uZInTvMMobrCV
flBuaUXt2XiSt0H2InfkcuYrWjwHDVtIGHwc41ANj+ILJGJUqkAlWxZtA5rJQozh
i69AxwP/9xu5PHZAz8aCmCbz68dVQVjza5KoTMAzqpSaATV9XPq68gPmX/rqfsFE
hFJWYBoYPOXjxj920nfNa+Rlgz79ONpHyfUaxBkY855+CWcBZTHPjX8PqBiGFnDa
plAzezYDWj6igPkuULA78aGA1Dm+g8+PPwbDB4GGy7giZwzkFi8pWQSL2BZ5ZiCY
XaDgz/0vmtxpXmNC6AjsHza4xDtOD2HvDZyOrucmm/HLmqDtmRSfhQqcrK1G1FE8
VJMLoUP1f1+w/9Yy9YrMIXOaFLXhQyUJjMLAo2hcLqRQk9xb3rrbYBGxA8x4EqXl
9BBVvSTvaGlC3AdgnqTcvJ6tiHeQ1EACn/WIb5KeiQrMPpPV1RR3K0P0hPhk1XE7
HHRHMtewHdZX4vhzX/PEE+1qfziE54eprOFKRgdwi9hSLM77n36KxHjg8aEKig/M
xWnC58FtKnjvXg0JE9QI/OL6M7zqUbrKhYBWxEqM4CSZOxN8EdktE8jdTKstqcoK
x/iQfWsYgDOHqF6eFkOWg2KMbLKkrUBvjmOY0awbNz9iIS2uTOMvw5cX3144FpW0
LnlF30l+bLOlDWZXZVJTOJu4o4EHITR8R1510hSY7ZHTRv3FvseqfdSw5YTRPnMA
MCz2wWX9nupRi1IB45JPE9I/3xG3VzE/hCqCpuyjdFaf395UYFtTybNpEemtErWs
f8L+3CxtG/Y/HO+eAXBY8xT5KgyrpM79NBkrP6IteNl5XR5hoeffa03mTqWXUrI6
e2Jp1SHqwWAaJ0Idx/NkvLkRmkgAu6FwrW5W3kCDW7/81cbgIvRYkwZsT8RNZfE9
Jb+VXZEPVg2hyMzDZ14de56DpvRf/6lU/3LHQDmeQCgjf1c0hysayplqdBvE5W1z
1xjOG9kwxvWR1N5w5/YGfmglHArKXIcoaot2W+S4UhrLgQHVxUPiMUuUaU4aI/2V
MlyuvpZlZBjyCAk/U3AeQ1q3gjBPh6fbNZQjpwoJOl0sf+MUK2gZtzvp44xtsc89
1VMl2TEmzLNSIi/2rLdqPFTv+Q/BUF5tCfibLqHvOJPC2WHoPfdtu7O1RkHqb87Q
oDH9o7N247vPqBWMGeUmN09ED/zbMsPoVj2/aPtmNaS+/7rg22qmVPLjLb8nkAU4
a462N9CrQWZ21HUq/v7MoBVg4TGr46w6daT6X6C99FKeNML4rRf6R5vqv+AvLr6j
RcdDpXgqztjPVmbxVaSDNA32m4UnddI0nULjhlBqXGHkyRxzRWhhIgBhRUSHLkBm
CCYkMLWGHQh3Z0MsRMGVO7R0PAT3PVTcRq/qcHUyQRaZ8wyykGKQDFG9rCyq1VVi
1rjcoBs9GGwsHylzFTLDoX6eqV3h+teTC2gEVcMDDHycMHetQLZop2s9V69bLGU9
XT73x42gkbuA4hiBDnIf4/0yIMaCpnGlUnI6QajJ8dEwoEImDLL44RZacJnqhKrw
B2L01dTuhISUqSyh4pTyfTn5GVj3xmOJv8/MyDB7MUcGOx3VE5NwitBT/3ou/hB7
2ddOBQoa7uUEd5/jM/0eec/qwFPGb6d+TFSOTFw15GFRCsQn7ApopxA+V16d/bnY
fxt2YB7gigM+8lKQWZi5r8PPULwd+gZqoCjNnuSJ53wuE9/1lcFbRUAdmetiqX3v
YSWhssE8AwjUiWIb9mcqW7aYpDob7RKFFW2464gLdgwnBkIloFzh+sWVpkrXJRJo
+ca/trlKEFlcE6EtlyujXmvkNNKCUhXI2uvUMPGoXn9fHV3tR3LDF1o2zfkSA87G
9rX6vZFIp1l1W6uAFM4OJ605XQG091/pxxJr12jn1D+Vh9noH1CdkCqi9deYMvL4
CK2zMOb/3kERiDditvnCL9DUHyO0vz3T1lUJHv/4plwVZZfjXRBVb0/pYLMs+Su1
Rl8OBQOSA7DQRQ3U1x2f2DPscky8BicIIiuSW9ayeE3Jct+eUABT6raGc73eihWV
/P6ystJuxPptn8uZDNO5VPTk8mBnbDQVISaLhtWUVlEaeMusNm/T6NyHx6OdnizW
64DIJoMpSEFAJXy/NYquVtETv5+JAgSU1hYEbrRgShpLJygM0fJ+kQHE2oGfcsY7
LtO/U24Sj2DuqU461z4nvDuj7ADsfN2CD14zGfcXKqNCCQhS5dxemag3JMfAxIgo
ru9Jh9i0TC6Dv2GmNh+Q6thCI9A5arRU+Ms5iiV39UvyP2aCQLLd8Mz3/gB/AsIr
oa/Kj+4C/hJ+3s6n4+KUyruL1EfSbiF5CTyrYQO6Hhzu39pLYnSz+5Oihr2JUgZN
63TmV/OekmRRAFYMFgysSUlXoYf1gvqf3Og/NjzAuECaA+YcQfuig5nRt2Wm3l9I
yfGMPGvxRe+rKV8J7a0gP7WW1TlqMcXpq7qcO0oXIgC0O642wWxyxFxRFhpBFRkE
M6bCSMofaJLmXzFYWAtp5l6keLXcdTEF5DnDW5YtxCGpDyAk/wgsv6GfUJhZb93C
d9w2ZNttAWiA6/TGU7g5Akz3rOY6ckiKge5/g3469TnNuJ4jEmL/njA8MLsaPDKA
Oh4YVVdinexEq3ted5nrInc6TtxG47a8me+1/y+OVc26d4ezwcFrzkwC76JtzlBP
3Jg+PmCGYU0tFnXxquEmUaDYu92USiFYbsjK76llyL5ZVjp7ag4A6yCd8jQ86zwI
sy3R6Rw9cNRhJkXPeDEiM95hp2V1FYck6K2AW0MAzj1vRSqWcszmRuag7QKZMB9F
9UTSBN3bE4tuB4JfFI+hwl3MeR+byd6WoOwg8Qo9xErFbQmFASIU7cd7JFHl66Pq
ldtXa8oSs/iJdrb7iBwZNLIqUWBFll5+G6rdjdX6gADHJFpCRgqQk140vp1itDaT
na/TQmb9rji7emm93kUotjNy4lh9mfhUGmqGjczU6cS8CnlxlQdjj1boNEnlZIT4
28ODTZyikMoAiG9y8QCBAqEN5/qiF4McXDy6rBICWcvZrpxNIDFZibHuqVMAQ7TQ
LI9c3ItVSbBKQ10bQNeZtd1i34utDrRRtHfWcw/ZC0eZSjH1VSVIMTekRrDWeEQj
za9uBXT3oN0I9KSogkfZjeXHeEPo6k8xPaZ+e+hu3wolhF2qzwbxNiTtBQSDcJw8
Dc17v42DPkoBIxYM3OG93GKHWYUDWq0RHK4C3t02+2e60PMBe+i9cG3nkBosDL/p
u5B91D89QbzKU9vxFQ38GDxXxoEEdTqwfQx5JVof0uKNRCaDY8vs+cIBl2u8FxWf
gMgY5z20vwKep1SqXLk1/7b1xYo27DlCxOxtKsCOJpBds30rp5nkSD/XbCEmxOsA
gV3AjVFkGvsU9nSpjVyV64qZ6aTIMnOtreNlFIcxSxGsaMlve6fZBkhU7iObEkNQ
8A73efhtaJDIHf1HLtOJlU/0e8pM7p5QsVtGCeMMDO82vYcqf8kzlv9u+Ba3NgCc
eRUkJqbOZhnBuhd98xT/OBglZW4qvbWXw/fdMQIkPl54gBCdtjZyapfnZeZes+uG
Uwz/alUREkSsImaKRGb/mRX/F9KYGiI1iQMn4eB/PGLAaoBDWpSt1/Ioxwqa3KG1
4bXBsTqxMer5UuHapVX7rAApx6dEPrbat3yfXEN/adMpVmwoAUeC5ZZEiuLiXYfL
czXiUzqmvoS0RV3zstBu0WQSYewodZbBzqyM/wti8bmvj5sSOlDyLyVO7bShd4gz
ZOxUW2WHJU4A5s+72IqzXZ0LEcLuq39oB9FsdXLFMmQxEN8LYZbUC7Hewg9IdYya
IEr4uIVf2Tr1f2bAkyY7jgeO38/00nS3vIr1IgjDV0LNOJ4cLGytWj90SJbjhVWq
0N8KAkXrPNuy+PdYA+kyxfyRbbw/My9WLDILa/rEp+oXhBuQiESCotaQmQEJwyxj
jvDaROioKOG2+6rfIguXCvWsmU0fmD/14jC0Uo0ZaQHQ7GyJq8DoYo/6VR+cU/xp
ZwzzgkYQYB5qAX/AnMjQzhUqLnz6e6VQT5Tvco8FP/cDKiE3cLj7Y67aUjW3qA8L
9rUtWgH3FKJJCyha+pcZtVf9FoNU4CqeVeyfOSbAhCBWQB0Bl13uguGIKTuo6dhN
zWoUxrpg/yMEGQErSsIU+WiSeh1tu3sBoa6cAXYR9Pu82Y09EBnHdn4dGf5dvMqF
snsJHXZZ3hOfsi6n6WNu82agZL7XbXyvwqmIGiAaJnqIVpb4SzdJkTXx7svyLK7U
rU8RdBqtINgmGQAzTFOajUvnc9QXb4dskhHqMWuKqL/0Wf4XE62jnjo6FHxFq0jn
5W+2Qy4An6dTzPvZ8nua/bbyuXaGKQLO066WNnsu3H58EiKpQvXiTSrt4v616V+S
PqcP++UWtcJmJ5uNEgAvIk2ZGwDVzl6Wg2ZZMunDYx2fgkAR9JU0ZeJzkNLob0L9
HFzNrvMg4ZiKxrpOlg2kn8fvILP3h4xH+n6scF+gUmYi+ngnYITI7M27WdKLKoEA
PJNS9lVGcs9RTEYGnd7C+qAWhlWzeT9n6oiLO/DdzTydqv3hgBhxzut7zY+Ir+9U
HZaGEjLnDvSBJ6spQJoRIBintDF/ZsiCw+VBYjWllwzmqGcbm1cNXEr/7JwU4nMT
agDXTZiU0uoE2vkDuNRPlKBI6u+QqUpW4tcwOnlMn8e8UxRgNMmJ4WCE/VNLecbb
y59+r2CN9g4h0hZ/i7ZQs71VlpScoVa2/etqm/JyxlK1EW56u2C3KVFquSMZtldk
PWyDnAOp1CbtbbTo2qrScHlPNDWAwLh/jmnTUtLmueqq3K87dr10NiWvSV38gWTu
DwNy0XrUd2r7fYzSGwRXVVuhh+C74S9Gyy9HBoK6ftJXzKp8s1vKAhICA5AI//rK
6F0Br7J4+BfxsAhYHNoH2kl0WKrgySAjFoUAGoKI5B4bpo7dyJ7xV4Qapc23IKID
zLoelnhZPmBWtruaTRWrAfz6Tw4/Hp1jQ0vBsM7mBqMxrQX7moNPFyj+EE+/ZetQ
WoSpWKXGm2GEOgU8bRMXTXIN0dXqHte0nAMiTAZ9htizD5KkSEueViRpO9w96XRs
E5JBJsgT8XCMxZFmwkn+LbfQKx3KHI9AKLN0ncSueIxFc0lVAEZ0m25y+52EDc1J
P+RKebUvynSj5H+cwmPt3Jt4p/6ZEJGKu9z087KS+vzk7MKSgwty+SLL12HX11nr
5nQtw0u6/edAvhx8GoaBDZKCZVgFH3yX5in6OHb4U/V9LUIZUyK8fDrjW2iboMgv
gSsxcTWd6PQ+EuwSAXj6UjiAq1nliDHoT81hG0CfsCn2Hu6M4xpQ7ezy9e8WUijY
htHf0f/RVsq9SEq1aoRpf1lR8ZfQubjFqszOTQhQF3C+FIld/0sHSBs+Wgs1rvdD
syJGRKk11Wyis2jex/MdM+yhGoOpPNEinKzTsE4K6NEei0vknCUTCOyc/nzvbaYA
tsV4YYQFSUDmLIX5txbT1pcezQynAUKWyLzT8UXyebfjzamV3XgUGL9rkBBYrsuv
Kml2EfIVOozme8nyq8qM4gLfPBB1F/qH3opm6u2bQjB/8uw0rLGtphVYgQe3gBNQ
ijp7O7vtcyQuaInthibidUeke/O1sI+h8/ItOmaZKW6Yp07KBOZuJYhU58pwre1r
7mOsy5QSZWER5MVSdju5vxUKOrmDcONRUHWzCuskZ2Qn9y5u/AJDeQjZSK50A6hD
V6k/R1AE5lFqoVZlZMVU8C29ST/QXxiUXpcqV4YRZW7XFDr7L1oD/XsTKfCF9i35
ZFna4SNwMtGso+nHGSfp8S9MqaajB3qh1OR78OkIlg1aevz/vdcrmsJn+BBGhm6c
FAkKyUsPZiY6LrlZOa40bdf38nHZG+iHgbXz2BHnNSa2H7JMyUw8xd5sUoEm4hMx
I7JjeFg2APLs8fnw5Rfo4u9flQKwlxFCy93BBv3McyieUUrBRMPhw4EcV4Ymt/D3
ePCz2r27oXu+yswsq9BS1gdxe2W5k2BLbhqrv/1EdDSW1R6kmuq6nubhMLXI/0zJ
UcGxWSQ17e2VhOQm0mUCg7sh0GOMrd0CHZQyrii87lwEpBQkrFUQgio3jxdWsiRR
KyKZ2baeK6siGRSYtMIJOZwjdbeOoS9bitj5jMT8rzoZddKXIQ/lMJ7dJ/xrAWYb
J/v1FzTYdehtlHD/b+X5A+T2nniBg49pcxJ+7HrOJYM7bnWnEYFEUGpV41zFW9+K
fjJQJW5ZBwyyhMdhL8MRA37rOjkHhaJyuitgY+pkWK86AAn7upfKtD7PJ2gjRHrS
7whBtA5Ew4Lc2qys3JPW175UhHAOsJxD8WOxoFiZb/4offFMp+CYxNt+Ufyte7Jj
L7Yr1c9EwqT3iWpXVbC4WzWfSrg6GhCD11nqxOJJecKDcumqlBKWEfJ9k/OeIeur
Hgg1lECEIzTlw57tKTahlANYCCtWdf9UAxwkm0jRxqySuQ+WtMDZMcJCdutL9/IS
rQqB3olEYTVKMcbV6IbBVOgfHNEvwuPID/Dq50llJ/L3YvmjWNY55fgLkuMNcRvN
OsopTFTh4+bAfj1NQjU63MZocjNwplmx5LTUe+SibhfSA8WLfeJsk0l7v0NIRRGb
L+z+PNLm/GBUmGt5X/1f84iD1jNtyLrkvo1DdB/Bp2hltUiDXVBn8ToniBGuJaKc
Y5t9mA6Y+v/B2HlNpP88krxK3XI/33jXN7hH+wMeHT6g8nzqeYKIdmYnE0N9y3Mo
bEOhTawGLGfnfNTl+g+LRVQ0SROjhCC89xC82rcgWAnjaG1m0NJvuL1ulX6GJF2y
r3ozGLBNbBj+tVx+FB1lJxUSFTFnKIuRi0R6AkcybuEW7BPH3OLnxdE1xHXn2CRf
tJpIH1GbtiVh+EhUNAn1n4IxwfPovb1o2NWGRj1X+CzOa66UljdGG+xAiQox1FVm
wSDo/T7mh0Etm+ThJquZyaPavjesJHmSEb95zult2E0L8Bg2WVIplTTKT+W7DM4u
/TRmeNMCYQ5tNE+yuu0q76nzVsX/PBB0S4xHa5JUGy5r15lA2POzmYr73ZAE+IXW
CgV7DuH87oxHCyqMC70FbrctUit4hLRD5CazLw0DIqmdcgr13SvO5UJFW92NfYpS
DNUiI5GN6dckSmuyn/RZgLtjErHOlKYOyP/LwRnmuMO/owXkSwCPRnSgH15tGifM
YsaEJe1j1fwwnoSfiGdJKNK1jwttokcdlYm92JcAa+mjXORRZZiLN0mbdVyWSQEI
JZXFNqSHfGsjlDwL6P7b9FD3sZrD+zOR/yHJey+/OxqDUPIkITHzPYtg3ElxxaOq
LnjupWQ/JnIQdq11sY6vyHAsm+Qiau7xhtaMbE52/Kuhcbjbd43vi1Ojt1Ic6s/j
wZpO1zUDdxLQoc4VOJNZ0Ln6cGFhc9o5Ve4yyCKF//5Jzl8zSeTkVg0eE9NrtEaJ
yS/EdZbh9PZy9hKGWPGOhnySny3uNGD74rOTUsR/RywbS2MHA1zvP7kdf7OMlraB
SDIBnf0mNFPsHOyoyq1GR4jYRhgsqAb9h1EYLPK/4giMVVtRBQb98hZfHKv+vxyP
5KqwEOZrTtqgQ2Qtrt+42SvAJqGVPY9j7/LfVG65202ZsTaeVUji74YP5ORbyXd2
f3HBYClfbRTKpHgsyI3Xi+NF1HOm89RAhDFC1vSh+fFrOVGa0eXbc89u0xIsiaA0
4fny0NWbNRrsz1oQ58O0lp5OSxsaEeRpb4Bn7IgLK9iwlZ0/BKvy+octkXFMsqN8
EfsI5123T52XFLwVD1zuZx16jqII3DEEBf3QGtV1EWrTsmdLenQkWPrh7Q+KUxlg
vuEuSla519aAYSFmy8ZeLMheZUobFVPrtMIpPLsyGW6OVtCdxEIJUSoDhyd01+qH
M502edyZRSIfd9z9X2xZyY8tIj/u0M7UGRY5bDrcit+tz7oijjsSEhiLTdoB+NUA
QW1oT5OjTvQ13SHeXVVywD647IeKoirW+yJhVr5ozkSbgZ95dvXJvibWBD/3U+Oa
9QOglQjUdYhG21gDZG974bv3B1KigYcMkXfzhNUsBDTJ1uBwXEs6WpobQRWOBuuQ
PwYHBrpEOMMD1G9Ncry4n4N/Ue0iaAj6VtORb6wSnEHjJUftsKBK1+pgHZdk84rf
IDfghvpf/flBWce8rdpB82sLCzCHfnUCqnqFKJZX8Z+6IV250QDw8ruinzsSyGfY
vsj8RjK0Wf4vn8rGF7Pem/ffEJv1gct16OuuqpGJTrZU3kjdL73LGhfKq6qUjgic
xETTGKvpfteNntWo4tVJebMRgmUVKB5oAyYy870ZjzNQ22Jz0msAhnKNnhnpoo0t
I/rEl6NMS8fBzuviWFpbHJFRTiibLSCR7HS+9I71wvnc7T93PrNy/GlXwQRl3Kuk
x/u9w2ifXjBc+/tb2FduKSoi5292tYy/pMc6+/bUlLiKgHtRNUKQ5qbmK0JSO/3T
t7Q3r+gBe5uFLie9/kUUr9sLxBzmz+EVRFP87DrPQH3gaaQt0SBcxT4mAppxH3VZ
eFnh7NAsbOBnfQ/JP2+J0KsOqZeuZBZIij+Rlo7MXxiqvAEJ4zF2npSKYqrmcJCZ
whYEl25U5+qQ74QnOlycCqF0drjSMc7etCHe/Gn2wjb6KhIaVmvga2JnNXXdVQd3
na9F16pYTKxKYikMPfu1N7yIoCXeiXxBds44VCjX2/LIiiEIFUmBqlQ09XxR0WmN
LiYGrex4Yg/b93bDC+IYDSYJRcE4l57Aw4uQAE+XRukYIbu4Snt0qNmLEcesODBn
2m+CxOHCYgPNRbSu7ItrqgPAgksfCD5AZuaJUmved4IeX1+cVFr8zJ35aeQeEeMn
7IeRAWxey+sFnSMsH+cb4q3jnObqFR5p+wggHmOrWZkWVlQlBkcD5bZv3SwRKtRY
e1bMBedDII/OiIiTotJD/k+Q3WIsqcOMeqsTUcCmmc5zwLLzL1v1k7SufDFM4nNo
GFGvO/Ts/fhvOV9ONHBH3dqlIo3vXrzlFTFnRV5HOhBvlJ/cqB3eCUg4HIZBw4m0
8jtJvrIBy0ZFZBHmcCyeNAdoqtp8PhjCwwpgzRMaStZd6/j6FDjtltysfyNoa+ol
W6D63PlI8kYdbDSr4aw3sQtuX65OoHq1qH7qJc2HurR+rQZp80plOFu+pIb1epyB
nKwNV9SnuLM5VCtVDRMJBx9B1tMDbADdyPbxABNbXzVcID4c0WWhMXpl8S0PL/Rk
qiQpxWLgs9t6KJU6gcNoUNHpJ3qrHxMvCyOQEkVx7FJe7iQIY+1lb7Hl+ZRM7ifS
ohM5rLGzkktyxVoxoGhEEiq069tndrdtYHW93nNkCaRHrdbxQMHYuIxf7F/yDtxl
sm+449lpLFcmIpsPfOv+wM/MWeNOhbrfd8R3sLqfYiJB/XgnfIswTO/Cg/btLNiW
/6FyKL/AecADbYsWD8ZRjnmWYsUX3XXWGlXLvrRHvtPugMZbu6wqxpJ8b9A+TxZa
7RcNtB/I3POBID2l2v3rylWxb/oTUe9DiZdFWs7/02BaDKcjaa31VFO9sqS+naMi
9opw2Ndm+7pGF1y0exIvZzSE52+fADfmwTEA8yvoj/N1GpmWg7w3qH7XL0T4ZQrw
zXsd0EuGMYpQ2yiHMgH1Lt6LLMIjUONc/ZGMurhrVHbBJ0X5bArxHtchYEgPe/Ss
2dTLljqZlOm8nre99pB/X39+CF8CWg1VYus6azJcXeydYKtrMzUE4SIVjs9SPUe7
QzLQkApHwttSd+svrOqWBz81e1HxDXirOlWEVjpbM/y6Jav6CYh93CX4t5LqjJAl
ZKeEXPW1A4is0UhDKAnL/AUOCAjcz/5Uhtekykfsk7Ilr36ncEaRzeVeqqTE8eEZ
FNGARuHJtLiM9xGyW3hjG9YE1A8y6rsb2Zc9bLKGdFghbH1WwYKbuSYB66jMD1pR
YAncIinzq6yQRoJion648SPBEozcuSlJbV5lkRNs+3t4SGW+tsaD/9Yri1e4JA3r
uUQb1cgx6DQfIn3ztPaJX2UjXbev64hVz6tAfgwMaCEGIu2mHby5XyKHI1gFQDpp
ExZZVPedNcJyj853oR7GKuJGlPFUgewUBEjkTVjrDq+PZIvTPlR/kUM0aSOGmRMJ
VjbCIbzTw3DBbih/U323KUzr/jwfsTpSUjJBE8BECrwffyY/ynXZ0MgXT999c8hJ
GtXkcXb6LZ9kB1YAvhN4ixXc+joGVpO0QrfHd2vR601bHRdwKEuQg6fHzZr7WNO6
rgZbuSu8uLWtPAT+yvMA+dXgIRl0bSIPhgfXKEH0BKgNAGvtbpWDPXkDQOHe89VD
4NKulu4Rl86pON5jFAzH6XEFjQfBjO5LMY3+AcNvQtF//p7BdtrKOAGBRxQ+tNqC
JGEwDo3/2XgkAFDDMijNF8AMrnKJWQ+B/SBn9azq+oyqSjRUn/bsuO/XmHZ8+7Fd
zIQVuoh3uo1jCt94yPq1nm70h1CuZyZ4ATaUjXww0s7blsUapAMCBJhg0XjYAkf+
fg/PVd9ctrQqXBNtHay2TuiCHL7Vc7QXIOv/KZ8EpqGdBtkcj4WnoQ68j/1YkLDb
jGT3y3XpQoymmt/W34OgxMlgen+1ffV6tuqGjxeHyjYC0yZe4c7nfo0nv+EUipAy
QttrOCoR+L22uJuKCHIoGYt8KydnLfTcZaes4WjN96/SrsCenE+VQeLlfdm+84/s
7022F+ygS4kRbenOMYXWesm9lqjKwanuFs+RSUMj6FmGURYO6QtezfzQYqFfEEeg
+/16G9bwo09lJzSyn1h/W+cWlme3kWRZOFkJ7MqVSE402ITm7RD2OUfiB6/WY6Xz
DpPJ4o5AC1qcfjzLtCLFXrBtiiSp3JfznNOzvktYA0bzAlfQbaxuoQMAX3fI4Diz
v2eNydl0FMC7Fh3GnmhCowUBcn054WDoghd+GbLYPbodhj2wkw/05TDypMlDiCII
3A8xYcu2+0rEIgQvbwE+mzeLQDNeK36z+dPFqxjPrrPNGRjPoRRzYJYSZjRB7b6B
US8o+2FjVN+Ylrugd+JWeBnHubWf+v3oaCiG34xOu2qsci3clnofJeBY3okPy2P3
UOqNRlv9TNyU/OFXDyEeiOJO976RwaSMvUpYts0mUggohC2TpKp/1EczXCpA6zyq
8B+9rKXlNqEGz3Dhnj2eqWscrBWP4nxJbXhri3u9vFQIQlPCDX8HVKOPvuVdxU66
ScdXasgsi50Y1d1sp7btwTITuofgYVjgPRewy92caTSN9wBxNtNfoh49IgjHjq6+
G2TSB6ETTDT5IxmRKa8DolS8++IS+HI5iRNYGxQnbH4gLsDM5vTHhQoXmWpMKBY4
CCjqu7oDxF2vZenvPYavcZ/Pjn3/C7FTp/kfLPK4MmB8AbzyjtIPWPuhk1pDxNyz
SVFrZ8kt4h3sVFJF3iSgQDO8h2XC/ch3nsjVJ4buaUAg/ah/87rq4j/jPMg8/kQB
b1Mlu/6eLJnsD8bovr6+Rzs+IxCECU24xGlVJHZoso7BSH8tOn6jWIsBkfWfHfRF
rYFHxvSWDoOZ3VKaORbwMguUoy5ILrA0vujNr4mgwvr3/HeEFb2T8iColy4OHXRh
19U4a0xgCs5ceagL2Q/sdZsyCJ6BFGc6uf7y/0EVjcKofRfJXE6I1CVEBRdgk/Jv
d/dJ64hv5+7jRArgHdCbadIJKcvatk13A3tXa8cbD9GMl+uvksz/p28Uebwq49LE
pSB1qPTj0n1GXMbiQnC9m+tJheKxMVm1+4+vwub+6sqzAQ88ZYcKagmXC3WBpeqE
rCmxG66o6oXbg4rt1GK+a6zI7YcnNAmq+jfXigvb1UaTz1bJ2tawP87UwpkjvcKv
Gw7MCQfPt3AF1nIsg2bpBGlrsNEzDe2RF9qT9iwAho+p9uoJuaZsq/ZAPJPQLrnt
QVe9lVdBEMkYppVvqi8ii6YBr9tnYpPx5YytoqyF6k4SPznbm2JSvSEUdqUzd0Lp
tIQ2VhED+AZFfE35PKaDrqSQAYPKSZp0tsL/qb9A65MWkP7HQGYfv0kmsrUzS+RK
UprSwdEs/FguBJASUzAGbEfiioP9BU+8Dh6rCPdiTwuRY6MQ23NAe/DqLwfsJpHX
7hZO/P65Z/V6+GRqawfhmPPnLFv/Dp5KWdR5qLYe5Dl/z6yiJcEWKQoowMlUDrme
nL6+tsyXKk7rvE4Dg819V6zLayfmpm4tf84p3pyMHqlVIlr93mPGNvffHfsdsTlP
DhZZdmzEXa4+Sg8y8fQZEZJD9LkmAhpj3YWf/FozFNqdv79EI/8x9oYEQg4DUJK2
orcQKG770/ms7aKShLcmWPu5Lr2faxZvFVztvkZrV9RhQysQ6xUa7vFu/L7NcWh7
1kZHofOnML2Rtx2t87BJ88cSxYgV68dg/UZe8/cQ2/QDabhUjKAhwNROP6Yp7Her
MOkPNmgimu0L55yPXKPEPk5QGiLeYQXy9LFtT5TAxkdQfm0b5xX4d2UyZ9RgkNX2
EKMvGecti6qKYy0to9fYStJ9o5xY/vxcDUaU5LDKQHC4O2tkq5wVJZEj5GZy0AsL
ntyMmzAP8UqxS5X9IIHIvg1iurcp6EvIoEWsNzuWjLvH2S8S+s50QlqjfXsLTOIb
bK882PVjWRmMhIJelg2O8GUhgZv8BwpAeUHUc2ZqMsUDHy9ggYZ3J51cr+7/RPgU
tGmj+vWYCwCBPJApn9kRVCKRWvSXFhAxKUgPnHLl1xnVJIKPvPkPygsCVx0sxoDE
8PjWz2Xx161NRp1cPw7uQ1ZLD/8LMR48eI5PG6WOUvo+VlQJIj6OW3ZfAU31GSl6
fybrOBDJz8H4iQAShizlHUZacdfvIx427PadXXUS2UkyuQAeOA8xd0IPelTWqQW7
IN+jdgYZyN20stcMtJNKFsRjyS0/0oKEkfm2MghndW8eBRreR1UWNj3rQOfkW1Pd
V34AdeSpGh2c9aEs7uBWqRGAHj6RVHxcV0L9qRqC7zzRpmIT/2gLqrGgc7RWHwZZ
uHdP8WyHY3AZe2ZyLYOEPKza15hSZ1YFnb1f3YXVJ9E+B/vW3384td7lCmq4xprK
isei9I1vgdDeXaQMJHLK8NSwtxy59g4uDNadZSRGeC0d5FgceFRGLFKcOFCsj5h0
oAYSIM1zGyteFiCl3MWQ+FWuU8nHjS/x2kuv3vQpM1mtEa+h05GQAgdYIJSHnkWp
isMhaTnZzaOKWcLfsi7NF2nLrdr8445lbONHQ0RrCjHRls44Y//x1IQtQ0/SOUYz
VD5oqoNPEILnkn9MH/rT1MNsuQV9lR0bkI//aDS3Dquk644/noTuzpkaoxRJfEhr
lAwmko7d8m6gi0Q9n95VLCapwu9tu1v1RZoBv1Cx7iBUVwTuATQdTHM7ywj4sYS3
NBwdd9qJ9+o+fHN1kM+uyMZRJTH6qeUoa5XpVav5bv01eFbLba/cd8OOatjmHoPe
QZ7FSK9sMxm5XaPX+38bp2wRzKMVdPfqtQzpZuXHEZeiqKb2PW53CY62gJPv6J2C
/cjmKUkOhftqehs3I9PnkQ4XqWS0pyPNvRjOCyVcnC7P3zcKXGHc+r5QTVJnnz2F
mRTq1kV3xNlhXsc8JKqL88d24zUaLYJo08QJnH5a43xFBNMgK2Wp2vfn0bQfUbds
6jtTfxmEDBGZpQ2Z9oW/GRnm28sHMUPkigNA6PPLSAuaqRnQ+2A4cPrOvH8bruDl
KyTHlM3taMILm3XtneMicx0oJ6qzHfFiTRbPSkeOd4/Okc378UQBcT07Ma4TkXn5
ZXVOD2YivH1pFGANYfL7Zk5DslExFHNG4ZBjCF6MqrzGuYsiWNZS6hq9nwcqfxeZ
0FF80fzuipF5NbETzvxkMn3Eqbwoh1a70YRfg8jfR2Xh5ZV9rBGlyUP4sET///oT
KLcT2+3QdRiU0re4alQIiN2XGIN8uWbqebLo4fQpZyAK+17g8ittMY9O6uOolGUb
CTDxR3Ov7ZwwiMIdsJZYcjvev0UK1RKe33A/HluoQW6Ncv5CmaBw0fpAfRyM1+nE
y5pzvLrvcuviLMK5UP6RMLu0+j3yHitXvG+76d83UCsRH85RIxXYkAUe8dEyIpEx
QgmoSDxj7U638quDZyRfjU/tOHTiba5+QspHxy7ulgq87M3iWLKNQ6pLg6dI9BTn
EFnaQX4O/WNPuLg+LFNicIrMvaFOFeQT2TLNZ/Xmbh7M0JMNhQWQLt49hOgZki6m
Xu0GJgNKjpjyaZp1qxhqmoq4/X7FZ8hJhrIyxfxOQ6EpOv3wOtLZgP9wE4qXVF9+
Mdee/hIcBwpPWFovPZEFwmUmgGO95JWqrrsahCgYmS97VQD+VU+DAJ+yfgntvCnz
P9BWvpHbwpbr+Jq5jRKZi4t+qCscf4CRXcnTAKrx4eDtbjhJ6VGesbdG1R2BGFq6
bgC4sSXGL1vyw8xJ2wxTxed4TBefdkF9uzZSDwQoWvLu/g0vp9UNG/HY4L6kADAF
OfTEqqJS5HpbgaVmllQAFx2QiISKZbjNobuqCMWCef3uBjtei2bZeood1UgFYcNE
PpyrJNr+wkWD+rg2epSD0khUv5ZxoHLTK0tadR85tSaRQn7aU1A/Z1BDB9A43lYI
TMdIv7Qd+wdKIT/5sEEudoss0WIfEdy35IHsASaaNkGZq4dHYCOneNm2HA8v3CwO
TdSapF8AUfLWu5+fIYF8ALNjuX2v86x3vBmx2k0azO60Bsxn70SGS7tUAmo2e2GY
VfZqxvsSNy85r5vztgXHGV592rQ6cNiPJELnPDBptNA/pDj4xvYYIUTCbrYXav8H
0Y9j0vu14U+haSA9sV6Mq2cF9NSx+JvMxFyURswUQuMzMGTxT0N5lxf+hsfNHTMT
gEhg96kqQFcbJe7YdbU03S3iLRBpAMEsMyEQPlZL7u/p8JR04nqDEwYpunXFUK3d
ddT5IyvSfU0Orb7vZ4vdgNQmLASI7C1uF7WYKO/pVLasrixRBUPtcUOk15aNhZKH
YuRyDOUR0u+5g9gy85/OTB67IMNdfFFt0i01tAGCut/HHYcwkatSp9DExb6Giais
L5wZ1VmqzpzCmswiKTR2PGS0mOrCea44Kr5FrgrhoO1bgwzS9+W246Jaaq5sYImk
KCbJhJI6weF9WSDuQqta3/NZvBHf/+KIj65yoliM3q2/R+PBWDcI2gEIPl8Nwy7w
4XGnjDshsBQNIbgJN5mWfr4YwbJczGlRr1wvf5yqCdPTz09+5z9IfO6JB9ZvoNgC
ex4kSJzxjVlaRXN+3qfjBA0WSY2XSTKqkX35su8L57fizdoMIuesKXjStqgR54t6
uo/Klp2kYFpfTcVBjiPCgSviE4x3Pbu7iGajRjRESxzuOlGoo4SRihSNJn0xj8jl
J9eNL1ppY+CrOiH4qrKvIiNkeapjOQvkgRjD+ifm7DX13OfK9Mgb5ibdrc94BH1f
H2DBjlcgsFPFpz4RvM8mFtE8xpXbyrgR7kvaHON6+1P0QzkffJTCb0aJj0zzS+Sw
+KMptJnJeRDQEtxojeVG9LTmSu1+5wDgUKC9ExxzJby+s/pIsEB1thmKyIpmZHSg
bbRj7DuORLvcEgz0hp5+u13/kVy8jYUVom75w98yBR10kfresnQPfUKC8AoGHkSR
CK1XLEOEgFsGY+WIPJqdgkTXr4EmntqcnYtoAwvqe+95Ar+TasgTD4U4iWyAfQMI
owoDYgmiut/z1XZqoBUhyYK4pv+nbanSG1BfYIRew49tB70XO1XVtRVu0Z4U3zhS
SSGTHRMtBPIC8TeFjSCdlTUmuoJFu8RuBM29q0/zkIZpuPSnd2l/NmFDDobd5CrJ
VXp2efD4y3FTzVC2vQayfolONyFdMK3fNIZPBImslte38EdyCMMdF014/F2fiFx7
gwEmB760SuRKpOfmVbOZW011p21mEvTpAInltxao8wmLi3apNrtzXsSurGaC5+HH
ZrjNpGJT61pKckmwFs2kffv8OyJa1yLalO5tTQAtFTk4s9qB0/mBEzdU3M1fA/ha
QwIESnbOiPX6U9xuV1aLDkRP6vUANN081gEpE5O7+Tm95BkeLkuD6VeB7FynnzKG
QeMQTfQJD8Vio7GJsQIzf0Qwx8afDc7FKflbSDyMfWOzOymDShfG+Wudc/CeZJSE
t9QYjc1ac6e+21JKcXpyMTT10GBGldAdDuuwzVIXw3SLHoy7JfaSVeXKvB5bC6PI
1fePODdmnktOjx3grI1NjyZ5Wk0B9ND4YTfuS1v0iIG9JxJgJQiFijao4YJpIJeO
ZvhnDAZgiaI+lcKUwCaHhLs02bFCw+Fec+hJNV3XGVcqYeLbpzSknUb/DX/WYPEx
HuXuBEaKMEYFc+NBbTt750yglGlgN4aTeagJLRlVldJ9nc7E1Ry7Rj6QU8EIGXfS
SZjW98wO0khqCI7zeNSN+CpXFRCpephFgjbhhneE034bIPcPt7/fWRx8fp/SIUzf
Wd4R/p3S0BthS19m7+DjqUtosMd4BHhMTdry/HKxYZYSnOwmuFIAGjmBb+h83Rhl
wcuvm36L+0efqbprwxCypoFJPhLR7x/4b7GxylFzfAWgtuTJmsSg2BBNFRDZp3Qf
dHAabIkSoQ4fIdTm/gSTCJ4Y0fuzL6KS0iAukESMtmDnzGxLKtrl8d1sTx5xLN3X
K3b/QyiXJon/kWbtFlwxVxy5m8XLfgw4fC498r/x2MQ2WQiMJes5co54RyicLzPa
eMXKIZoxLJqHHbp+t4TE0ZWWtShFc4RxbHnRhCOo7a97mO6Kw1sBMLb5V0N35ChR
hZp14p2ST7UluL2iESEB2xlY64vmONuw51HOf3vi6cPD3/I2vcIh8PfpAEsfWsnS
9zn4wqIJW8qJQRCH6frx2Ozw9Bbo/9NNTv/8/1mJsUiHr77uknL63LjqgLc0dl8O
M/OlzNzsH0UsorK8c5QHx53x+cSj+5kb2BnH2v77SXbYWTCrEdbmoEJZabMmmcso
vDxA5GKfu9OlQ5uBOVQLapW88VqmvTc8dMmQby/Yro20wWGZh1nAGfG/pWjcifNO
Z7X2CY1xeibNgiB4xjAXlu5sO6b9OgcUEvsNdhs9CLkTvdjraOfguvGYzK8/vB67
GdJotA5QqciMTMGA3O589pzg8y9da97RrSaYh3q50+W8o2sNRxbvwoVT7RGOip5/
BGz9ysr9kSwf2HzeUoJtxXpPZMRXwKST+0XezrkaLYKWtkqbioe+d4xwlJNlj1/o
9myr4NJK9Dte4ngQRvi4yXLOZ7jW1B6qQ4n5odd2WuF6WKVJnz4MPPZDIF5GRlBM
zvQTr8q+UyvSHCZ/k7ccDASOiRBxOPhTaUtYTDLlAsERBLQJVipRMRYnu4SRc1Ud
w2gFBATwh9Z2KpGKKe3CYRPc/UrN6U7gZpl+2K+Rbnl4BWXaDgYcJ+eqJVJOoqJw
OHIUK+1NfB36eI8bGm7T4eK+fOoI5z0p53XSmKpdl6te3uMqJS6vY4U4JTWwWfPY
CGamlz0JtSqo9imoCKqVw1xwfel9s5g/Sp+rJ4HjlqJcpViwYVeFL7jfdAnYRDo7
b6sOzlH+xTmqFcrJhBNe0heyj2nzoX13oDxHLLG9rdU9AMg70S0nHyKXEdgG3zFF
gFLM3nDjf4TA8CC3GnFu74kYUUzgZCEM+Y66jH9DYS3kdI8InuArlX5GxZVvF7eT
jOH2oc3JIQPbwmCQgutnI3MsFA9JkXxMtf3K5Jgl8Y2RxGwz1ENhE7BN5W2sLvc9
mbcz5c9RpjMCN9RRTdwH8OBI7kbse+sU8lmcBR8Rarp5BCtrCkCnY8LJ9/92fbzo
sEAakfSk7dAUQ55/sVzeDSDis/o1GecI1f0+PwAzjzNyEezigtfHLls6mTLa0LPc
lZyDEDFuDx1vNUU20tXxhd8LYcML7unqqJNxee8XdNEMPw/NBLQ5NCgej38I19Td
6+ifgx69LB76awMiEh5NdmmIiCzFMdJVwJMqwVuuv+s0MzXX1OYunToO4orPYnfJ
iy7knGFzwOCa5LpQf2TtVzrb9LMoMnpNEQhLYu7jmKGeA6+cH2CkI3OKNWsTiL3o
iTfrnkvYsXkVKzoEzOTthJtb3duwopzHW4tYI3uqr8tCSVW4HUgx0W926PP9LEah
rWMki5vKE7axd2JqexdKuEWXyDG/RDf39jg9a3Qiit1kG/e6c8FidVi9eZbywA00
7N7crc3fjOUtD89KKbIiQwnBIhSDFGdis8z1q+gBHoa/TV+FPc/RS8jcnZFLFHYc
VPMG6SjBYvMGQxp3jhBbu82ZBOv34zCE2Fb+nc5FIERzENSA8wXALoJWfvgy+1id
/A00Sa6IJ4B/CmvFiv9BY5xecSXy3E8M9oDLXUYPsjJXkrxCRQnEUDcdGKas9QRK
OcuCpPYXwgNZsFMkDPqDnT+TP4nVlbVQDjWtew9u9AtHTHt/MG4VJI39UHuTfKdD
tOY4ja055MzAIJ9inkUrinf9wvCn9SZMCleqAUOIi203O9+IMrvvEDNRB7MFKS2W
4pnl8n79S3WNh0v41SnFu5NcmI24d+r4a8rRPC8V/0S/UKye30skBv41eLx7AmBj
mvPJAXVU7/afgvsHAqCah/3NVXUwBZc1z/vJgh8KLZQX0rMwT3evJH8bZzi4Xc+o
Xshg7QyOvDavcq39ibp0sc9ctTLpQo7T6wC2ipheM8aX/E8cHGrd5yF80visiyh0
d7OOo2g+lp44cdhO92rFLemkNLLmhPMbtzOXBjxrkBu0faO4+3AVXEXRBRIkYz+I
ibNHQjOEMqzFsxmdeTT/keqNc4Kp5NWrqKCa4tJNRxiQlYkql/R7RaTuptXSP5qA
FflTZ9u/DUdBFgXjkzMtmR/VFt4ce004Vd0+m8nbmo5MzK9Lqp6Z9QpKLf/JWKfj
QSUFpXlF9RxL78gq2/bQPEaWiIs85vaNPh+KoWww+7NR0YFLT2gjZdzGD/rcAHwG
tDIwFr/VhZHQ+rMfjmBGoVDXurMXEOXfbtBKkNqIz+MtJhI/PRYCFVqpPx6WPGuz
1jlwXBkBNCwc0mTBcM7qx8FY+eZm+CIMYGA6TSFULw8GwB9hCekqjI1MoRa3tGf8
PHdlAh8dPVyQnVph6CsAvZn+x10A45aU3BEY3H+8mv5pr8LX9asjTMVx4TV37581
Z4UsipXmbtGHRb+/c16kRY0Fjdvo3iEyTZbCBuw1eJFtqQjL+OQnDc2TiPQLZeLu
lyrTRYjEtcNfEhNwcCILZbhj3sHeb/UmhEqPC+3tr7gPD9tg5PFjM8pgtnhIg9uz
7TUQHbuA+MJtQN8DhP37AMUK/NSBuBv8QZGdsJrMxQGlxejgtL7y2M6YrkcMLrhZ
5R1jih0zUQiRpa3l0BXQp54wCyxMRReu3OJsef0TC+Yu8XP+RR1UIFSMLDdoyWUu
QLE0ID1+zfkANXH59EFQQjMeG0HZCmIu77pwt8qr+I6IZgVwRXBZQLvd2Fhomn97
TpMJ3v52r9tPj040tBoCCet9CpyBrjTZCXQWNvGRg1HD2TAmO3ZPpCKba7nr/zFZ
n9bSXWKpxVbML4vTp/IyeG4PCNenrOcLWahoSLHVAEh6OC+DoQLHkjbMdjJ65JfB
nDYAUaw4kz90jZe+ysSCVMn9fr10Xeveo228XDTIEw3KalmDXKHrtCPFGMFDUwyu
7e1uoF3XYjsoapmS4D55NkXU0y2UzeOKIWsO3uBC6N9XT2ICj7E+dTrfrz42IRtZ
emNxMZfEPfTAuclEY227eWjetsZRjJ6IwcTP6wW8kQLOFipzZz2IEaTXqeXyrJ78
DczTv1ZW51WUtAJ/3sqEEEsM6MVvZGiaXqFXJVYG0yssHhN3CDTZRnxvFlIkA1+Y
RtKxDZMlVgC4Bq8GCn7urIT6SqYJi55RO81ff1JWe+ulfbjRRNX4zmPtzcJ/jbsc
jz5jH9LEhaBlcJDSKWdURn9arFM60mvLmELgy52ng2NmnebiU159576ThGxjiQsJ
+TAZkE984yiEwMWX8OD8XPFsExgqDCdHic04DG2wG6xk4qxRNPjjDbjwsutKEny5
kPIVl0sqSkhKaG5/uoKNq3SaKrMQ0zfBJscCVlDttKJWNRqzzLoK2qk6aZOhDPJy
z1jWhjx0wQ93FZKsJP0ddY4h74XhrcxIuDb8IQvQ/hgEy00dq+JZzifVfTCyFThn
xrK5lyrMsXFxOWNTUXbjANdHTdCusgDuIq4cF+dOm9QqzAHYaR+22eOMX+4JB+KZ
9Oar5OZnWQbBVdTKb3LLpkDDSriRuKZf3mldcwRxiZdYGPm/NmXdFHlEkihDDJTW
IS9wI9k6hhZ3BiIlhnUWTyMCeTyZ3qVcOCLUawSNXdklf+t/QOPIqddf8Exjt/lh
2znsH77/fMr1lsGcM/rD8waRhUYJ5sbTb8mbbaRtlMUG9n+8yi8V1IVnALTAaq/5
vUGm4QI5+EcOboqdkra1KjEloopxE694Pp91QHRZjDBZTr7/XBEPvi0N7HC036QZ
wojvsh7HaU/aJ+GxSOJokuzKscr8AM1aONaoTJDX6Pd404aY5JwPqPWvWEhZoIap
nd0QMrQ8Z62o5nncSvfludB9zdQoffeZigL8djuRHS0P/Kp08rz0kPDpk+3MPnPh
DF5tMgjr0K3HZMW42BhL/zGe8Ml8vwC4D1Rq6XWaTpYnhYUYbLZsFjPM9l8d28/P
p6YBKTkl43PDxk+0aMbtGBFuUFfgu0QhttSL9OExy3xCiB/k6+S8r0Plnf9hs3Rp
Bva7u70FT7tMwr3J1SkZfUjbihb6G08xeu4OWgi95IB6u6P/7huhfwQEJRkA3zyg
U2irZvzYicZCzaHAoizGEShBEB0nnQQdtcyAgZu1aapxpFVu9OE9YpIlsmcgGz6R
5wpcrDMLms5aGk7WrPUG1mPNFAEmKov8/EufU4lBh2Ppn15DXKiWBWUM/5kDIPIf
n+w+4JqNivsHBD/OkoQ4h47Oe23KDcvF/bWochgSjGNO3C2OeGaNuk6ySYuxAhUK
QaAeemRPqufgBxkilRj60cCCwIExXAEJfWEUJSq29sPhFxy1V4imzA5IPg99oRZC
FxPt92NkEz60mZsRo4PF8RrsBlYMkwMMn2gc0LpyKhuOUGOzz9ZPHtQu12dgiaCy
k/0L9ebO3wZkbc89Xd4K6mFwt3eWXvRkFjwdFu1HfaPvaLsc6Q2a0OiB64+dkxDm
PH+mTF2ZQj9kZin2BM3bdNJYVM+WfZaEKcPRtLGA1kYhbEg63CrKhLUPoJ1vjLGb
QdlDsb5CyPI59cFfheHZ73lDBEdjbP32mprtaZj5xXoWBTwcQXlzaVWABrOSy/kp
yCdvUNYNFBL/78bNbFeFT1Q4pX6P2s1YK9dKIV0wG75h1UtJpk7Ko0WjCMIwqPuk
/pxrwlm1It8ZNF4JrPh9sAJwgUnxPifWrJG0t6rZDBfOEc+X9rWwZy7UROEIHzsw
IuMijvPg8EjFApxGXNIhrydli+YKsC/UBUOh5IhzoS0zBxhH6csPFaNpQ3IrR6Wd
6rMkqqj1/lxGxw8TGOShHguhLWtIM5MN96lz6ujT5NegeJwVPqbArbQvq3h9Wmat
4Fr8il9nmR9dRp/IV1xOJM2nTE5VTjwisH1nZdg7QtW7V8n2QVVMYVpJ6e26Bp0l
Npl0780ah6MeFxQQ/UqRutLVJzEszKTjRH4NQhdeUwwv7ihfJIAjuNpn5jaDNzj5
jItKPtNMFK1tpzLyWkQBfw+YPYaha1NmffGXlcqctHRdPUiRijtMxyafxyPQMkWQ
4X5CFUfEKyRK7pJmje533dP9eKraV9yJX64uAXHooZtFR3ngvCJaObVW9YnaP9/S
zjOr1Ebi8ed5b6cBk7Gk+sBtnQOkvTXsAUWZtYmzysVFCws6qR//gzXYEeMbMxkM
By7qrxHRF+zfIpAqzlzkPTzVMKH2sjUj0/qSCzhK7q0YDKjCmHuiuvQM3HKMcOYE
6kpzRcXsGs7OIwPnfjG84NVsGFB2Eg18KysQEzSoCHF9uli4apXEJcBUDxiSCKFb
/R0hlL2KGHtb4YgJhDh1mghyqzfuff8dyWDPj8Xv4GawX4J/b/mAcLm2VpN+xzFd
pLO9wE83D7fiHXD8jn7kXS+M6JoUTnrdKVODhoWoyu1Gh1GwDtNf4J2a2zXsxFaN
pFkZ5pdLVtfShTONBhKbEgVe+hhLBYsWeEAcS9PlWdMP0Q7WbZ5THxFn6AoKsahv
ILqD/4HgNSWPFKUTRaXbH2s2psuYhhDAC+AQ3HGV7C0aWndqkeFaCV7hnp0LTdvs
uVkjMyTB02lRoH7BjdCZdkyBjI0v/A2UPF1y8HkQq2f/t/6D1pV+GYcgGiamLXZB
MqH4ea1QX+ggWkcOOKicFkSyoTTeRsd+lU5mkfu3kmiQyTtCmFG+oUEktloN50t8
SDk1bWvtvp2PSNIzK998pwP291abXiEEuLDLdHgnHbw6JnMyAgeBshlIk4gP1pCr
xGA/4UXcE6PXF25vsRBYz2YN/CNdlP0aqWEp6R1kmKeFl2naGdwsqMOdGLFfuwp2
4yCOywq8rRwTzY4vq1K0522sS0JRlA+RSUSgIQtflWjHfgvGaIaUF820+33RxKfR
MxXPXpiNdKG0gzcKZsz2pUy9iVGL4T/a3njBJrJUD/K5wra4TIVoykMTpfAk2ZKV
i38Fv6WWK0G/qV2FKvZgm2bRzrVCvPfozz2OyDAgS8LPxCMAE4ikLfHLjbTj/Ilt
D8FHLNC0GUqwyLFoKEmMzYfAPNWOq2SYydq9clZsYWCJ3+H2mvIHT5nRsUNFYWUK
iyhmFffsmm4tn6/zm9cuh4SAz/dvwmQ3DAv44nleZfIUtpEGgBZbwYd0p4GhW8qj
s5wD0SqEvSpVauGocXCLmMYKz/5v4ajp8CtNxEO/5edg6yuFgbwfEcKkNxtoNPX8
ca6DIWkI0ckbMeUQnnr+zBttHieTMRM6abxgiCVd19aiiRS8K7RHVeywgiA1uuY5
nVmRsHNXCK70IMPHjrBiztooI8fK/dh/8NoKLHatfilWHS1RjVzxlskobcaPuBe7
SRUbajsfCTgV7H6WXDgjwE0CFfU9jVfrRxxrMvowb9ld0E5+d5MSgoNMyJhQ6Adc
OE/vBp0wWGMyn1Y5OOb/+rsT3nt0a3yH1WP401GH/4OvuejcBpyDIONRsMylska1
Gbg+hteB1v2Z7IQ63AyBoSYvXq9Q9LA827w3uOgUDAlBHwmz1BawVH6nYr5qts1L
Ut53xpEq9n1/96igA1vSyoCwvBCEdQUfINK4RMbHMISqLvnfHvcEzC/xhAEZzqeq
F+K6bL39dGDcuSCvy8rsPR9GHUvWLXODD0ecZF0SXVwcZv8667w0w1r8zTBX7cXc
+rLYvDRj9vAu1ho9zwPGbN+QIC0DzJTtCrp+TV1+HhP9wUx3NmmolYYhn6WWFS/V
5JYif2hSbEhNex0w+4AZbXnmq4hnae8OH2V9X3an04SsywJ1YeSqwZQse/VaCqRk
mzzV+qMw0YIh4ZjSPZ1QN0JkejThml2PW3UkPQHkRGBy6Od3YoUSxa77yEIg0K3I
XpXcw0C3hVKvN8gBs/8iKssjqS+Wd+wCW+6gT0GwtFixHsbKSPBcQzi5B/IH5uoq
zLYSoXLPUb7bRXfsXLtGpqQY8zudMdzAnFQl+Ln36IMW9YsnMmGFIJvBt32tQi6S
vmh+Zzhoa48HxYczG3twHtMv43iF7Yfb4XRh4cb0zyOoyfw/qSJcq88HJG6Qmbwo
pSWmcrk81Z93foytfiYSAiKDNnVloE+0wnzkk20LYEnp7ftbeEakmaU6Fu7C9+Ml
Wnb8rFsSFJQjoL/rJUyIak8StqAASLhbnCG5quar4jMnxS1IcYN0FMMQzVJrx6Xm
PLt7oy8pKETKyk09HxaP4aLAvbl+hRjTxYj8Dzk/VUjOf6oakOzpw8XDtHiwzpgk
iAuLg+ffmn7raPO9ALmK5ROgnMWMtjQ/OUxVra0hkS0jTJ6XLGgAGgDqtn4+4qEt
JjqKEIJzbSYSs4WWvH/UFEmPyrh2Se7ZoC93QgY99veFnbd/xgX5OojxBu7PRUS9
FSAns8iWnHfq+b/+U0uDTYqjdsin3KqzsSu2RJiuTavC6iRyD1nGcnE7X+Qpg+OB
RW1bsfo4b5eCoMPiDKN0bQK3668fyq1I+RrfkskVwm0MCgzbDjnb23fsEoQD7i8p
wSa4EcCEdo4F6JkS+mVGFbtMdDR1rkXjndZ7sfuvO/zmHRHZ7ot6HIuuA4ip7iTA
kDJ4+XoQFo+PeDOyZZSAmlu6tOhT9pjrNtKXM+yqNA1Oqq0uZijnBg10nnacGttW
BIfU3jhuU2ys6e/ati6GFC48/MNPEYTq+15TXdbOE2/t56ueWL2fRMRqfB5WMc7r
hzk57QsicK3yyQP7Nmn5n1AZu/ggm/yMtZsUjXnoZZpYRZT4BN86ONj4iA2XFb1P
+um8KTYmgxsyARDDKFgoly1XiW21EkTu+1d6VzrK2mS2K78P+Y/XAqnHBehH4+1d
VeahvGirRk2narkn1oqUFGexMMnDsgflZKSW2yXYx/r9M9g6m44JG6tc9uRNIXh5
cmaHdyUtPNlze/FxoM3laaWtDqb1dW2dSwmgWqouMEbItdhyeOVeSZGySOZZmiAF
3XbrHvS5I2KP/K+++D178qbJo7SIitcRq1pPFe8wwOFRYKwKJgBleo1x/rbbR+Qb
oVNWbovqIsaVpBcX44mWVNHCeev0rqxxPZYzwZehfR2rFBgAPXV7F1Xv7CMdXEGK
+vRWq0MH9DY7wumucqaVtYb2Q7qyctjevOMdz85hUrvIDrqgMfhCYEKMw5hj7w96
c2BWrNwqVvJAyRyRuqNyv8uj/XsEe7N0ehCZDM8f2HQCEbC+haSDOhbEva8d1KCv
Tdx8z7cRgEC8u16SOni+2rrmN2Iyc3eoXy2xzf1dXDSPVqqzDzD983JM7U/YSqPo
9XxpjYLPGXAcvWg/YzThxJlpVj6JVyABLALnS5QndYIzUF82xOD6RWm3ph98PMJd
IzT4UtsJSeLyN6rE6VW5foYI5vrGso3A1wqVAFDTnM8x8+22OQCZLy6CZQC5EH5W
K2/JG4gLXDuoBfEzEm5YaPWYYdm2Dl7P+aG4Kpc3YxtZ1QZC+JZ17jUSMSmMBoWx
NlbsN0K83bGc/8N9xGEIWebCpRMlgQ3Jqc6luUCHp98poJTJ0x23ZZ3KJX2ZHL88
Wq8NxjIOveZye2a+M4hgEDWSl9FxVNjszs7Z9AFWy6sj8kjSQa9f1nMAM9J7hu5g
rd5SiyaKGSrVhY83bCDY/1SU0J3w1m09SmqF4tKEA1F1mZt2qLdrem2aF/XfF+m7
7n3hVCoOVCrb+hw9BAOrxOkupA8N5f+z8wDEYL9JiPNT/ScAZfzDstGMiG+VOjBq
kn5ryFZajcDzZqdQeljs/glGIEPWwUQRO7ZsiGDN/SGk8rRoIKCIpivsLa6JII/2
6VSRHAC6gmapEdfwCSy2cF3zmq7jNQ8CB1EMw99Z5ze2Cfgw+h8XP7PohejPG01h
5P3Y7ThBzPEJNpGEFmBK3mQq/l8cKH5VWYjWrDwUTcSwLvMyBo6nOgG84Lx3y2SJ
XBkDsl9k99LBPDNyZERKmHN+f/20ZL8orGN+xeudDv5di/otAbKBd52MVpdhY/cw
WVIPWYCsjJbzknwSoZ8jnp6Gpkp5+Po8y4YvC+o/UG33u54kN2jMmRl5CQ0jrBTj
UINJIIfC9rbtHFnxs18+yjiimZUH1H3BwLjDoQNRn2W5pI9bJ10L/eQX1QZV6d8C
bta7+uFkUmr/Gk2aquh5RlvKk/CQE+9GxBswvhhfVle2HP6VEIGdkz5qqaW1Iv22
IthRnrYCmJxmCw8Ajp6tND0W4eucia33kh0boqBcl30ITwwdqdL8cqhTOV/0894/
825ax2m2ISMf2DBHqvT9pd2e7o0OJlzroa82TvWHOJ+HsHT/95FetQy3mzVMsrzZ
FbsK7xyYFDvUZu58tumvi0BmMKvjW4+ngv1xN1nOgCP7QjOsEQQr07arsm1l0tju
Wb45i+EokExmVXXbhEjtg6rZyPZJweSfQsRlYO594cLZNIfFH+00aNPzcY6eD9BQ
aUbyPrFbs/x6DEs35jri7+tg2ShnIcEJP2GItbLs85jyd7fs8Q4zcHNMuYf75zAa
3B0oJBNnfGCCbB4Mb73tY+2VEWuyePCYqwK3DEwcUEcsgXEOkHpZ7Fch06KS9On5
38fLxwJXILNOZPlvmniaSLFIXV1FOT5oGRGpgYJ6xONiKbiADKNHAqR+12Gmj+IJ
QnyDXzx7xxO8TG2m1SxtMYnHx2ZtKH8DVdEe+swe5A43RpkbBxIC8w3Pot9g+rjh
/K8g+ZhE4COKMu6sJMwN65J7eekZLTYucuM/LSKpGjV0O3ZFLK8r9mNmKwojqbQD
xSSoOHzxZXVFIOQlS+UFpguk8/XtdR7NmAckAa4DF5ozFv6TYZUksxYl2LuUPij7
nlHiDfgt8bBESmwHSq+O4mxBXYxesa6ksATAYd8Hcgl5omdgbWrmYSACvb5hNx/n
MwMwln1iG4oaJwpm/FAIJG9akyRVfxpPFdgMbNOBi5y1Xqm0qNayNHM/OW4IOGGk
yFvcKH0JUT9GAsSLnY6N+5x6UMVjrODssnK8yeLw5vGKj5wlFulIU/Z7nvIt9yk4
/3N1oYfCq8o0D12MSgVAXTqLqCcu7Erj2geAskrXm9bc5t3NFBbH1dLBpw+2JyXr
rt2AU/LWLsqzXoYawePyoOayipheHtNKG6WL17K9XIn+LpYoOnRiFqCCTA3kYFbz
6gKbeS06PPE/2YO0lq0Wg8E24A+4oiSOgbQ342QX9xLyYFZ93kBlrbljzq2ydnLM
K0D3c6Wbhm78W5tnFor4l7rHzIhTP6+c4lebt7e/K4wm1G4KgZzofBl6Lsjg1EvN
xDGCEs0KDT+/MoI8swuCL1pC9jVYEptKa52PnGg9osz8IzjIVD2JSL8i4Ymqfidu
4AcIufODZrUcynlOmnfhNV5li7KoI0biu0EJcfvxMH77rg4x+s60T00Ry8XUymqj
V8oRNI4Y3RLTg+XYHGvbvU5ltVYxVJ9qQtscWwmyHKltKqFWaLT5MtF5ZM85Lux0
ax+xsL0AJCBZ3UvVuAJ9gHCS+DSMENfr3juBAd5r5aLou79rkwcz2/L/rGrCk44t
vnQtq5nMWje3dDXoZ/7Vsbpbdm7wo0x3eA717vjjOyg2Mrd/K23CdOerg3MJFZdS
uMFLHCK+Ebpk79xh1wroHhT4FWr/hZW+05sXqddF1wX42gDuNVFqUPVQYAn4GHWE
W/ySI4FlQgQR00fuWO2gZKSJMB5hLEfC+Xlj/LqWtNk+XFjTnvHdKccihxgPpvEV
ocy+7a1PZF85jDI59sSbSO+Hr1dE5Cs8mOnIF5D+2xV4cmZmQiqmGVBkDEMUCFz9
jiD4dE9GZsIr0Vbu6+vf7Vbf6ccEFGJZoj2HCAu2Wa+UhVu2Jja5BNAP9p6NIfAk
MC2dYeD+A32r93BcQxCpUokjOLnMTzvWE10/ZiQ8QXKjrpZRFvImRhhxNSECv2Wv
t9qUrPmdm961xBvgg0CFyqf3WU8RqHHQKQkgSrQJiK/n3ZXcHZThqGXrRkFj69pi
0Ez6TaSh0MsTQQjveFL+ebfjyACxbHiYd9dMISHSEK3Tbo7GXbMlJwD3nEtW8vA2
eTKABfQyNZVVFHsJRpqaoPjs0fYMwXUcEbOwnQEYpv/HyVG77H4d+Gs7L47vDUjA
DicDaO/Hu4QPEaeqHZJ3Xg35e6ixDJZIbCMVCFa7ygj1ESxu5hWwkSWmYwRHOKFW
shCxPKSWMVjCV22u43tfgcmnNNhWgn9iix742RwrKBAm+JbWl/773PaFb/ytTCPs
6njCpOmPV4mhoNOwbDUdSGdymqeUfd8fxQErY8sWz8he/t356ckpNtasXFuzrxdH
4DZWVNW/8EUBZgihIOAnS3YBree9yzdtea48hM8sXsBoIrkAM6qSuVzTFiUyIqbA
M9Bx5eP69dflN0rq+ugCw1DDnyfQ/KNChg2u0+R6KbWyTPxLSd1f+Fp6VcqVONjV
4S602x8CDTJ0DdfnZ1aRKTQoouWhq8bIfGV8m5kgSvK1jSBBHEN3+1Y3YycCtX9N
NZK/KeNKZ67kNFBlBya4rmpVe+acvcRzxWgptWgNiixrHV2Hxs7GTL9QTwc7eP+K
st56oasDWLGCtTUQVA4PMfFbJqfFmUJVpfGAD8WIbnQ4kK6/HHk3yu/m9pKA/2Ss
TYLsq822LKOYDHQAl1A1rTwA3jGl1ZzzBs5JDiBVl/2Uv9fVWUf5b2MV43dmxDWo
QCT8lZP1FYqbjULkjh0p5Tza0gN6UQXSk2Ra5VRQWr/0OAMggwDa2sKwgDCRhuTe
/fC6AwDLgzTq0xPwhB6IMMRSqzjTHTK0c0lhuGamuOI6vZegENme3iEXqtXvBYcc
fhqf+821dHjT7gPshO9lGMiS+ENl96TilEaLG1nsYF4eJXZ0AZ8RzeWyBP8paIiY
4cjmt4YTYeedStnoAAO5u4S8iXeX0X9rLbbNIoD57HIfkm23sJh3wJl7l77Y2zqn
U79SP0pnXXQqLtUOvDUXcltyZ6ZeaKUIQ1g0CxNiLszmWpw34DScM94ZGNkGK/7j
UL/9bFVGfIvYQDH4Mo3dfYXvHl+VZe/QjJrsQTYJ2+0umw0alqAXRzD2a+p8moqI
csBhjJYLWLJT7ld2Re/U+fM5hY4KXlQkKRX5wU8HqilPlY1ACwovvAGSYW9A9u0u
dTCWWPLlcQz0Pu5o04vkr03ay8mmU2CYOxg2lsVfptn8Q4uQfs2yuHRW0dl4YhAB
tYAravVivPsuCK0rQ4Ugql6D56ylIpfdF+Ym/5uqXtuz64iwyta3ihHL2uvgI+Qs
6i6CFvDYUw+LUuSN+3TY7Lf4v+oRMd3K0LPx11V5C1h0j7BYOayq/imOUOP6LMyW
+QA3APP6z8kCKUctypc2ZvYY57UUjNRCEas7Be1TLeXqlQANhdr8D3i3/8LaeqeW
obHKsT/JJvRPey/X7ryXLjzmFKS3jrNXhDLuyhrMfGrgMkpCYoePGvQuSKOMGw27
XwvHRPympzOga7ci+tY3OXR7R/Rbwn6Cy1KQPNS8m5nFHcg54xQfKMhMZ1602AW+
gZTSjPyai7rvPv6BvPVzN4/Aw2WOyZJf3Osa2zsu3Z3V/tOs6zKpiYu9T5U1Lt6c
AvHXLysT9SjCf7Ge3jpqoWvI6AXCblEpHVMm2xX/D711GgCIAXMGHL5xHYMWPEmo
/8mve+pMqlQkEM+FR+TzBQgSJJ1knivPndEDV9I10TBV8lEylT/gcHM148ket0wV
kJkUj95LvGlQc8T8HrXQhXILPIfDxQ0OMFZIimpV1mnq5uMA9GhUTfbQfbII+zEo
GFqYKB4aIBOhPiG54rg1ovdnERD4eNhrH3SMvcwR/dOmbPAFXOpLQXezeaTsqrXU
ilwhEG5rDsQf53sLZ9fQNUZ6eYpBmfKAsUlWp+uAaDY6T+adpxCa+rAt1MxAOTwD
loFLOL/HL/94KxE/07LGZXMVXVALDdeFPapdRL1UNX+qdwtf8n2m/jnq2r8yLXrM
QBcTMsyJnRsmRP/Fppui1flvGJVqMyTcgRyp7yGZ7rZSpDpqe/GJsts2xjs7jJw4
unSIgCdAZWjZL166i+ikKLJfAf4uSmdvU1OKQYp/29oJ1ywhkcymm19qk/9pkaLL
um+itsSsQ2McwSQghtWnsi2UX4qImqYosPJeHiOMQZVki99FSTafuflR5MpNwDHk
Ft7rLOWUF5Gk67CnBU0yygPQdYyEn+gOM8MisDRclrdIp9aAb9w0eVQpAMZYPATW
5WCNZcg5pgTyW/cDSfIhW2+AHVrTe5R0/EICWQaVzz7OYtNc1mT+9Y7EaNGwyL7H
UAcgEJD3NxopnTvmjCipNeyDsL/cK9MbtAcdEnRH6ygQE6bcwVe9OevK1nzBU3oR
IU0OyFbJAUTJubA4hAyr0DBy3OcWiAL47TWeStaPY25zuGwRUohj9yO793iEjkav
H+1mv+GmSXZZBUAmZS0Sv4j0tK1jrk1Xx7js86MDmX78KAJXbObVdkvFO/JZPdyS
hwv6wLzp6//O1uvwy0brnMYQpzL4mhwOueMStkdlVGWJLH96rY+A1Xo/mbKyYwkY
Hhe5pUDayEKASFRFDYBTe7O3/4+pMQGPFgI37PlmgFYJovljTMmbeG/vjMJfb7/G
+GYxYKW/LLl3EaWWBnv29olD8XfIRknboeCdP/L8QL70ULEYWm55mIkqGQCugSEV
NsRxsPQEZ9ooaEiGIi/DwA+lD3VuUsvxcRIKf740K4gf2XMUcVWsHYL1N7S2F+ZB
FBBfIdCHVkM/u2OTWa1IxATn/RybO+Ak+WsORvdRxSZX/JJ/Pz9YOuJq5Qvs4k9Y
GmhYfa0uDdYFyPDO7Y5qoevjMe2qhrka1kDoA4Z9G8ukWfh+fZZ7bshSo0Cnw5h/
r1BqrcOqIbTm0+FGOywiPsSdKT7ty07iLP6RB7PUjSPAZxb5aLzUVK1RMN7NkUDp
pzTITWvL1+mPkJ/cD70Nc6L/iOYgm3XYZsovkyUDWqLJ/jrOEJkUWlSKtZNSX2/5
AAWlEfmELTwsqgmrjiEDmwV4VcrXIWCW8kCovVuapOwMH80/A4nbh9LXcf6nbc9x
xSNAQDW1RWgExB23q4xKA/jQGd3CVInJ+aw/pYk/ApjJ7BLII3neEo/uNhcgP64a
s7AqLuaugkHbnj3IcUnfygMI+0iY44wLSJ0OP5aLDl3bZthbOkUF2U4pvyjSgxSt
hf1vi9XGcqSP9UJ3HR/YjZOz5Woc26rRaQuMy/8F3FsrWJ4G2GtvdJqIktIC5COl
Sdhj0t3sn03hYbPe1BYnHN7Mt5w5qJ7Aqqd3Xwv0sFUjfAdxrtunRKKR8H0TYM27
p8CUtKTZvBg7IWhbO4ZTQS8hVBmA/3Atqni2ptpexNMpyR7R/O+Lu8XhAWJHS3WS
PjMlPK+pTgM1+LcVtwxAJcmwnLOI2Yfd0OB39cRizrWVbagGT8w9Sk0muEzddTVd
9D2/qRBpvj6qqOcjl6LErtXxIgZ3167uCvPU/BfxdmrePMHalDS09V1ML20DAzaW
nt7hA+L8VqyEInfddLlBMsERCX4J2Y5Gm76oAfK2XD6aPJC1qj0yByWKd+dFjTW8
41tD+e/IqmuQpPli5VNc1TBsEXtQ68L7IF+M0gN0KYpe19/rhnx/AY0edUzZPXK5
QjtqTwG01Ndmh8mVcV5wYGI8nJBCaSMrD74Ul5rsAeXDJPfNN5sdsKPNrno0RJIV
WKQS/34xI8amRVZXVw3Ik/GxgxXj0qpfzJ0x+aPo/aC50n77KVfUy3eRbMzZPyEX
1xX3tIY6u3uT84LthjiwzXo+Ff4eZzFKCjURRyYgq3eMKrNQQ4Go1dNBuGEWNl7t
7zL+oZK8IHGliAFFRJhBIw0Eqm9VNc57+O6BW66eRlUtXBdSDZbys9R+tM87EDqV
lWdmESccIsk7O9iUOwi/q5mHlKC49RQRU1Lq61SL42diZNarM6RVpYmmJXdMNmFx
bOQrC5eCePJm0WqKCfdIRB6HgiuTOM0J3tRIxudLyz/brHtHMUwaCaZ1SVDsAp9E
Ug4VTP5qTil/GoOVzxywMss6yXvfaN5HZuEqMVBeCmEKk5UikGdNsLnGl1Bs3bkG
XmLqARCX8kHr+8eOdZp5seqKXyxtacrLjKwz5RODESmdrRvFxfkaSWj7io2W7Gbq
W8Q7UeSy7u9FPdCwPFOTutvZoRAO3saFfkPMtOMgjBhi7y8wpo+LSbfOhhJxoUUu
K1AkFg+Rlsc+g+DZtqHxoL0VRN51GQyyEgqUvSuTu5cO5HpmgKdH1dYx9MrjsCrO
47c0BxGcSIliS+kzfZARdUbWPsHSqc29Av89TYu5ujCm2qVW7J1gzlPY68vm23Vf
U+Jy0eIS8KkboO4g32ot3/kSh3bkqhcckaSgUMJa28JGBbe1kak6GRSHnTfw40MF
cbB35Z1CUruKkkWcNQNrMk5vThQ6ter5JiEYr4E9UL49E+XmbcG3EaPtaUoyJjtf
fnGHVxi2b5vQoW/+wvKpfDX2lq8JFbcMwR14uBT6MzyrPBofA6nVdPnrhD75yPM9
FBrWeCsDc7kvJ7qQFsLZCaBOzytjF1V5LJblYo1efbGcEwSx4FlT7LMDSNzfQALL
207REyW0esdhYErO3ozagi5MGBlPjG9DxI1LLMxBi1YH+3I16Tz6Fmvl1XmLneMw
no4wdy8NwdcpzfJU6pJAwR29QySxFTJmsIjRYpBIwYHFOe3kgoX+klK1WJAnEVqt
y7NlpPut1FBsMnGr89B/b5xCugUJf8/VScyXzQpKZaWeaS2D7yAdoITFCFaV9jNC
ihiRV8TMktCiaS6cbgsvvwIA6xC3XcuIW0QzprizCn78dfOjcSSioKVS841del3I
k4WtT3OGg/pf5rkFnhNwz1Grx7t0bYZPbfeMRqZglObwCf3YGpb06que0xEHV/Sz
e5CCLhsvC3LEMSVa05SnBX1xWxXJ/MnXlZz8R/1YbKDNMXKXdCXK6jpgRwV2cMOf
Fbgv7Isq0MdiHxmI120nbuPXfSmnKhWAwJ8o4bb02sOvs+m5Z52G0F6cgepxpR0u
40fGpHFjVngfntu85+aVjpqAMNlVVNJ5oyJf2ybhfNoT7iOXrxYnNXukfvmBh1Le
ZC/IiOdnk73yQmqg6mMvX20BkUXpx4DzYcWL5f+JJBempZPm2NbXTOTAzkpowJ3c
ujK+rmIt0R2uOiVGpxysJAMigA5n7nKz35tLhFaJk22eTC5p930jkZlBZXLg5yUA
KMZ/+tltdC5psKNw8fu1UwU8+mV77ce5xLvqfHwqQFvkBneLa0eAMTWmOPA/LOgr
qJXsEfM0ezSOzpe1bXy7jykk980v5+Rdc7d9FLMHtwpv8ChI3/fp+AxgeHZ8QymU
sCLPi+qPV8n2Gn9z1bM3TwMSVUz0CmihOeu+UnlRaR6Ocq/pZKPAk5ie3YnYgul4
QdevWjVKWxjD5xV0YC10IMuVO02c4zBo3eIbeyFrqjnqH3h+hiDeMXmep/Ys8VCN
IPQlofrp6VtculkJDuFG4Sgr1h95SWptVvs6FdA8LgmBpeJzUHY//hYMEIoITZc8
aohFd0k1ShgVZMG1ST5/dFg4aeGB2PA/pAvESoG+HwT2v8S3vkDuycdqAAgmKM37
sMRHQydQMEHtCqFAbUnYlEyZ/jID0K/qm+EP1sBwXDjxq5CeVd558Zt3IDIVBUdP
7r9PiDcDun672cC1Yf7mQ8UMws6Rytg8tDa0WEj2fW0Ga3ELUHRcRJuns30KYB4m
cq2WFFNwC+4HBB727NwN2NjZg+AWNACE9ofao9GQMZF2VIHYU+IqUXxe/gmFhqSi
h5EzUbkyKwRFYFkCKzqSQTnTy+hKTEW7HpsNE5LvbkhGT97EJaTTwcnluxKoL4YR
otuGO6UGnPfixpDjhTqFkhvKkIMRBsJ347ehE/63gaOsr7Q3qBv31VdolUzjnq1R
vbdSN5Vol48GBsYprZmtKCXNyIhrHKqu6twwKSxPX9n/fq8CzOpYDahgpsS4aSAk
jjMMNU5EbKmuDS1o/NYCcqQmcNbuDs7JvfagubZSjRs0+mar9xscCOWX+DysxWqe
/wWOyidgd9ay9cfZyxiaXL8IKSTMTIC47e9NW1lpPZzxi7uzmc8kRlQfbJDc4vma
wEoLvDBHbn3gzFo45ALZ+lak6pExDHsoBipojMZysfVT9eow85HaWshFEhGjK3NW
6qF2Do9oktS/boUsDR5XA9ZGyoDlp8bo3+g5mlv4vzvCmTEj4vMY9SGwHhOeUiZw
AUR75I4Qv/aB4tX7A4TuBxPf2MSwTt9v5F93bXtz1z2eviNU2l+sRTNl7knaZf6o
CgWcWoVTskTp9XS3RmLPVmL+pRZeqFRgU5migrjabwJB9d/mt3fNNWOchS67KuOc
I6kMFxGQsChtANj9+3FFdCadqwwWLHWBZ8jdo3p6k2M98w8JW/7kT1qjQGsiDtF7
u2raTC11eksHyU7z3JiLlqX9LrRKkhKeFvmTNWaPdpsL3D/OWv7pfKDS4cAZedW8
WFPDMcvKX1Zbo2SakUyk+DwNA97mUy86/+VOZNoh3c44Awb72eKqfs4aPtFFak/G
LEcvxt/dKEMzzrW83LLiifBl3UEqY2ddXff8dgLjObn48nekQIcdSaD8aIwTUB3v
tVO/mU76Dfd9wqJ70U8YnKU7zdg/tHXYM5JX5/XUQay8ymeIAtNgESXzeIdAuf7E
uJb7MUnGkMFjnQGjneGJNXpoq3wfKIS0H8E8vmHCzqeonu5svacbG2hnUP2E/Yk2
gKRzb+NShBla8boXKwhSXmNB8Lxjntu5YsjLXYa5WUbaFrLaLtG3vSmQaEmBCXcs
uZ6w29OOnggrz58NYf7BGAfiK7xFNRKazQQ3tGhhWS/pH/OiOKiFtBZj1m5jPRVq
YSkqz9+vUei3LGLFKoWQ+2radxU2rJo0IEsGo2QpzlL0eZagsFxbe/LaMVNeVe1P
lg5a5we6n5lV1ZHB9bq3RO/lMM0xOqajRzo1FgLkX9N+VeiFKpFxYLT5lCQtCsAD
ad45V6v9bs8j0KGzWkTVfOkFjm+GCSWQ6xAqjmlRAdkTWDeg0/+VzLgbzEW9+Xt1
OdBVzZXsa9UIvi+2eyL+V4t58ijMiJ2Ap0JtDvAmjGAKqYSZ95KoUU+H2oqsa0wx
8LQ2eybOpnvTPE+nNsDk6d1y1do3mQxhvRW+KDUgxjkoIVfi4/huTnMKxyTSfbi0
Vtw6ALP51OslgsgzydWHsvg4Umlisf2O/hXogCPulkRnpzeEdveAkabVnF1sHOmj
xEYqsaC8yNPx7jWc8f6ZtrNPfllVq0CPS6LVY7HmeWg+8UJg+bIvbI69FJmkNrFo
COm8RJmrcfS16h5sZzkIv3UOKcxC7Bz9kyukH/diUy96hvIJazhfLwJuhg2vYKQC
iASGTvTy0dH0y8AoqoqJjrOvYft0jTEzTRCQSupSPy7rdcTZRtfQq3CJqx5OHGCm
dT7M4JMyfGP6eG26ofxC6lY3KX7iWcAqcDXkBm+/S8oNLuFsZC9pExHroju/0EXJ
e8BDeFp4tK4CFARWKvYue8iCEfRoj7CNbrQfceMRfeCMc/037NJ1QOKT5SVpVOQJ
4cKDVR7OMvWCxIFB6Se7JdbaMEP14QNZ1m5dzGBFwQW5ud5vwSGKjITbzzIYLiA1
Fd4DSS2iTIe+zJxPRbAWsNS4KAP5M9U7zelQJpqAA1cDw2CmBAD6lm2UG1+0CjRb
YSXlishdG7d2Ic8w4O3E1d4kIWKPg2xjNQmwGXitqfCknjdgJL/nFoqv8Ta/JBTZ
4bTVCyV879bHigds0r7Usjig3RjiTbBvbjMIt0u7gboS7lvlGWZSc4g68vhUKRp6
f8C8/HcWSqE9zKSBv0wiV8lWCAYL+U/qw75AlQ3agPF+qOg0FBMSLA8AfHWuYDbp
OCk4zo/m2a8i+Fl+l7PZshJdN9xcfhJz/Meq1/5De9dO9ZkD8kUg4tPIgSeV69cd
owRQghPA2b26iq92YwK7RWqgRCpan6fxm14lL0RjCNh+Z2Os/Imi45TC577UZpUl
lAUrY5b+xfBrnnWuJr6Z3BbxJVqDJooSC+YYkEmk3jnUezFBOYdDO4fYY+hPNS3R
EDl90wr+6qGPfW8zPvDFRX+JuXOsW1uxk6nSYZuWukwr8/7eVlEUrJS2a1FUeMCx
Zc59XSw2KYMco+VT2ZeFNjSjpHDgtjy+f4IdMak9653dsOsr+r/UHFAvAJGJf2ps
qYUwX0PoHFk8KaqmHrh31PEpYOukctIJ1OGBMXSDjRWqcA5ZAnFldQlxdnHVZGMW
qAsiczT8nDwz+vf7PIbZ9tzmc4F8+0Ey8q+tU2Y99qC/wSkjbAcdYasjE1jSegUE
SfsVFrVFMLsqt5wQTptTlLyYvsFB5MucjEW4iWyWB581K9PfZy3iX+9iL2mrirSJ
w4CkHUtM72ksSZqpiU6Y0EOOiyL8CfIZ/IERGMkTwHBSiNOzJ78oFVlj7e8p9Vr2
925W6aXPKO/2+cDDRb0Bj1MQOiFyhzPkbpsiw1UtoSW/K1HwrPd83BNJjEnIS0WJ
ofx2CRi8BbgUNDDMIjPyGAeVZ8CkzoTYL19CobwRXiIMY4i+UW9jh/pHUMMEEgsG
+2/hjry6191MC/2h0ZF9kNKn9vSTG60T+YvfkKh527LXSXJ2+9qDuhzIiCFG/8o5
d5Tq/1TNMQWLjVjsCppNWfOaVY0HGrXKcB8MZXewSvEZZsVWMcoftuw4dU+LCPGA
C/IBj/R3yK3ThE0XVwxVHEMSSj09XxVgBMiGr4X+l9VBNqo/tm75oTcTT9CSvL0s
fuFyre+pcs/7i6/ahgVyPNtb2loIOiRhn5FaBMy7t97cfxIlwWG9VFrD9HeOGwo7
jGadssEc6f99Q2ldN0NOay74iq49GtwGD+0K99BeI3ZiI1BStAFvwjAMkJgHnxl0
Gc1eo82BJQl6aia7ARB8tznHCznkMrYDdytau5w39W09F0D0lRnl0rHqoap9MIZX
klEzkBKz0/twpHuY7nVORqi93MBO/Nl0GfZAhf42PMpJAwpBxg+TpEamXqBztcyL
JFEPlC94DrNhsPLM4GpGuu+iyFiaUI99wzomp5czeAsMG9/hzMQCrI2iwIYKXCYJ
zrdMgpDCKMSEedKgQUdAk4UVbcxEdzCp5I4Jr4McOrjxRHeuyqW6L3TRIs3Ka6bt
WAKkuwZFqHBEBxZrgDhXBX4fh2SXtKW7XNpbBd1Q3ObA9ZzVu7MacPZBm8v4XIoy
80xtBb2vtqdxvnlxkHBAbtBBXEIeRuXYbffKylMxomLeGyVRwoH6aN2Ji5bbf7zr
h44dP4Gmg5HNUXstfNqhLPoQIiyhuurdH9QGrdkN5Q3+O+hxKslnit3emeEmmSIf
jcPPTxknIUQ9LqCIiLNd2DxZ8IBjo6XyLkdLzEL/NS7U6rmrWen2j4EI1kgTMjVx
GcZKbAIDsH5XqSON+3evLy0XxKFngEpy863HMer/Bwzqy7xalUyGR3LUsAvbARv4
JFi0PXjopcRQykffe0y+v0hTvaLIWBjs9rLgQE7KR29OtfhyNvpv75gmba5qmrnh
dICLtAN4513ACyHfFg77e/2JdyKEimqz3aS/VchJ7gGUpzBvo9UHC7xGq7S98MZm
UKYuXvpe3p6Z6c5Z5ejLg3P3AYDgXwNcPhxXz2CLnJ91Vx8Hze/kp+juSORXTWMv
FpI/7CjylDWEA0ELz0bTmeMr/pq5yPN20OWkdvHTtbNb1c6RorEzpDvrFfkEFhG2
1ega6W4ORopjy6t8eqZyQMfts9FVoYYrTQ7AlelNOUO5XeC5T+gDGMIt9MNcsBnq
M0weTsDlTjp6ex2Q697JHS9/zf7CNtRmrx9SngZKW/W687/29gqxSoqIJKhIY9wS
tDUOQR7IqNxspr5KLTMsjn3E4aXLEbEvvdQBGk5f1PThpWuMNqfO9lweWp7vJqXq
wkgjB5ewpCu3ggiC+uY/HGWjz3uGznUBDgFMVyElooZH37ko8xp+tmTsw/3Wumkx
1O01feMJFqfZuLVbmTpfciGTCBVYimAySg6LYh6XVL2JgLbTxDG29zO95wcS9W6C
ZniFHzeQjkACD/tXn3iJfBoQWvKF1Ho6PtZSDdorPOK8/NFISBTdu5Fn03pSsnJ4
DU5AI33P3SiATSK9Cb4EyOKNX5DCSpQEUoSOrLE3H0cinK1nC/OGQIRSM5Tphs7R
ET5X5KS67kYvAxYfZaHG9aLIT6ySKBQOJWpy59jh4hrMBciRumG/QGFJinupJmsa
jrJE0YP166cLo9rUTMdIPJm3zwa1uOyUjAF1H0DaLce2O9G+LRaFz5g8epozP3gH
YkI3OEo/QnDOyOIQZqTs09vBzVgXgEJMVAuUpr0xxPEny6/BkjpM69QicNML2kE2
iMs76HpfQW1jiw8cn+qnGVIWSisWNGzpvLMBWdrtFut7RZio0t6bJEo9QchNeO5Z
aUGIBLK44vHoIfCJWzeyV+X5eoCkxH6P8Aa1g1EyZxDz4lPnrrMym/GfxoczpR+M
/ZrTaioC9fxBQ7m5S4tx0wpGmjT8/iIxX4aJd9bJjkIYY/2apBWROBG+iYnsMBri
FWZEANboc/ovSh6OxfhMLmZ1FTU+ABAnuMtZc8E0mGRdqoNt1AuXQOzOv+/N8H9u
fhYy8gSF4DMPlq2QxNxAVib9Ky2SaaYQVonwIVkgCKdwBEdh6+3RcJpXvsyHTcOv
RjwB67+Vv0D4927Ciw5B1347CW1mg99RVRTWnBWSnAEErorIXx4vjsH/vl047Di7
Y4oGu6xlyDjJ3dbbMCZchaNyWJQr5SWMBirtWC4rUXyL68c2iGSVJLwVScHIs8CO
jBzzkcSVeQ40nNWC9CcX9IJ2QJ3gBgABYfLPFwjhvL7EyxmPmY70beKZt134h7ja
4U1UPYblxg/mpJ4MTQQ8cJbzQlLklg0EK+w1ySrbgBS5vsTbMArzYEJ5LjAeXE/T
TMi76VBs9b+fDNlJnImaDvg8jX1VB2ngDHT8nUQA5bH2ruDHzN4VnQ4XRbKc/3Jp
KuHr4L3mW9Z5deB7/Y1yKxBpoOXjFMJJ01rZ58SKrEbqM6mZEr3pJo6ekgjrZVpd
McJjV8VzlWT6Zu5feVdAoDRbzeHK0DPi0CmXxP+fxvFJjMpzKYD2ihII/joaiY6y
BoU1XQUaf99+1U3hIiLYgcvlSvuklquQZtJvPhRpHblG2F0GmNruEVR3mSx9YmGO
R8K/+/V5WmF8MLbkLSMk12Yo+/EM8LA3vFW6Hy3oHV9duihvzi4dH3w8Jbihxs4i
tsGU8FmkGj+VCbfDMC28ELrmoN+1H4fEwvxBcw+YMb/bd5yFIa1LMftguCgp9sjG
sNmru9E1Lnh3Fltt8SCbGfGkc6VGKozNx0mphSDvEIMWpBVAhSW+/AZSY1fal4zH
ImuwQMAwC7j4nEnTsvJaHmJyOPobmgQJuKl+yyTnOtBdK4rfSBconfiFirHAW32A
kqrtZaLvk9CpnC8ZCYYQu3PazfGfxGqabzxhfAqDXmWhPiqP6bhsXGX05rhvOKjd
7sdMT/rHcbtdi/GRlygtfXsPK5+B6CGY34is2HfZ2JM/XmrYeY4k0orfEY2RnnrT
ozXILDGGWIViTZ1uGA/9mXSYRmDT3jWOWlTLhT02UzyA23McRXgECQ0LzdPi2hPj
HOwilDmqhqCXr59lvAhBAXuTlm6GXT5XHX77H1g4UHvIMEHbpcvD/GvxUVMh4a9O
X7406IH+tpB/jUhcUnCsJvBSlXiZ+XfSJvUaUL7zqOzeNCUvOEPF8HFHxvzq+i0d
yf1Y6bjmFbpxXtyXr903EWO+cUvXTRVOgz7QXdWDepsKfrjRefcvvWiSlDH3G587
jEd32c/XmtEW2Fhki6GHn4n3orvYCWTJBqB8ImKvUoFREbFijTlSp+oQ/TsmyocN
zNXvUKDqXw31cJY2z7fNIvZHsEwfw8sJYkihfHc7emfw5nspiuN3DbgiTeiAxxWm
JlQPwkuRLd/1Mg6ElCSqhL+hw44N0k+fjiPVGKetiZbp+ghJVZMwjVCIFFUuZjFZ
M12LIBot/rJQqzSOVYNLwTtU3d8zOj32xRn98xNWA03jDHggMa5ArNmj/ZuCcS3H
Kn3cqFXosBHdLJgmYmeJ9VnGXnrycTbuyyu2fDpaaG12mz6KDPgW1+tCOndAN9Y/
kl9RLA6OSjRkVxx2Jmnu9VJnzajXZqsL67ouqwgNVZzbJJUuGGd6th/6umCQPPS+
mELIQcTNxuW5+XqnDNE1HDGlIG6CYPhaZwWgmXPZZeInLNqsQgfHIRyGmPLjv+Lr
KEAmqwyqOaMKc3G0xe510DPCy91uS8+dzL5WmBKdE4op6jGDC8G3TtVcudIYQF9y
OtAu7Lvv4zPHCruP2bnQQwnAUVmuF6E0AMMettQQ/RQDKtWO5e/0BoM8odvjzwMZ
Yu3Az9sBMSsPpylA/ZgccaWiMV6lf1t4WyNp+LCkggnjjlCGrEDrXy2Q4Id7xdcT
YGNICXfI7IHpsnU1R6OZk43TaTdGeLoh6tF+j1bxeOeISNbVpuG0pvimotLMJVHy
Q+2snEznUmyQJWs1ax3WCdByTRyo7lsXAcyuDeFyu4I9q63SaDVomjTHY+KJzGeY
cC2wun6YICj6QTCgViZ22WIuM6VheCtM2+acYNOEbVKnYuqEIduMFy4GmGWHAjst
X+ey1Lb4MH5oDKIlrmHVIq1hcps6l9t/M+0vgjVN/Wg4OO4YlSTwRRQtNv0kN0+B
GC9d3F9DNkF0VZoFDgXxBrDn6oqVkXWbNID28cZyr0hRCJeokvvTE4f8Rfk6o7vh
OBr+oryCVYX+0KXGMRGM9OZjMxdGyAVFPRYctVcROCwnuso4G8J+8ogIV+V3hAKU
Pyk17rYiGuMhsj/vjTvvUadSqRpqNvPNz12ajAcMKd0yZakT/eDL7et2Ussf/BfY
Vqe1PvysPhGHMI/N2fuDoovySsJlXlJ9XT85FtfkabaMdDj5zI9fGPMzPMKmc1i3
Mca/wRJJhL7uY74UKM8DW+H2AZjPTuDuoy11MCpVsNFx8cenMfNPOda/SqYTgWD4
pf4FqvDVo5Yrh/bidnJm+q8ei5HC0S4EY9cxc+wPfdjNWdakx8gyC51CgvJaOax/
3q7Ob8JYlsBpGiD7n/LkYVFoQ8n0b1TYhT+mfKxOD5kbmbiMidG7VmOUwPcYBKdX
YhA5epHU9DMHL3YEToJUCh06zpTJE/vQgmPmIY/bb8dpavdRX5DHXavoV3c37Mnb
1ngPyGSmcN6UnuMGSOvaX7XqN9tMiFUzKAoA4hbusVnZw7dgWfOGM3sa7n5ides+
9GCLmWMX63Bv24y2lIHZ3efyim+JQvUNHSXwSNzOM41HHymdoD7e9CFOoV+L4SR/
H/pdZfRxgOSACthl+B7Rrni8MY63g20s7WWxTofsXqY5EkcOeS/3BwNjJCvFttN/
UJmHAjhDVCcezSANfiur1I6NS2WVw6ZyLrAzR6+NTjw8HsYdq6D5mbtTDcrDi+Xw
PE494kxoyzSz6ajqtSWnSMmylkeMqXpOU9P6Gm66mdAxRFPcA0nYFZl3lQrvFbG4
FkO91n59J0KehxkgE8EU2uGlmvjAURgF8qnZWMljE0BL6u1eEPQur8yjQ8pRM6JE
MxujqK9YLt77KCO3i5logi1Hui11BKFY6ZdZx2V4tcNLi4RzSw4pfmLQzZwPQioi
hpVjewr9ge0w6fzI6xWKofu0dtBSAepJtf+iwkvyOEdYefSXcXb3SyMpuPwNU4se
S5WcN2eThKSYq+ECl9ueZbHuFA0YpSIVvDiZEU7heTn2wnsXW7f1/tcLBpR4k2VE
RQQwAx+fHTD3H7D3HI5C/uDlhOU86+Zr6+/y0aADS5DI3s2XRC5BQH0WXaf6GTtZ
eV4LGGjzpMMRr+YJ53kRGjg19rTHbC99h7WrCdrlmuTUoZwTJpEbheMNxXH+EZ90
Ac22bJDdSyolODEuP7OOJo5XiX5p1hGsYIlbHjA8/SN0qjOn4llUbHu4yshGS4IF
0dCKPuBIqglrnUMCvXNUAQdqcoDkNqxLvyGZXr1/cytfQKfQTHTLbHZPxJYKKq/B
0+WW+2nwuRSun6tY+Bf9hRCQJX1U+NERAs8Mq+ZgEMaRjrOFnTLtJw4LynlA08yD
bJ1GgR4V5cDE8PrRNi7f0DUS2InLFnAu3QpVZMMOuSEt8XSK1V5B0/C8sSGypp8R
3XJakjed0/Ktv2tVGxybFZciXxqxwDdIBIgxoO54HfO1TblUOeT85dlLDnfGH8V4
yZo56/lO2grY+OZKUB3eN/qiVCQ2FfMsNNLV7xmThV7jkA0UJZoq5+Lp4xZhVRrm
iLs8NW8YBmnUo9PEDTh4Qvp2m2lcifgpEkJJskSnZql0LgCu/1/GlErZUl/kkuhl
Ho7SiDAvlm/iBqJp1lcCTuK4crLB60h1dffb18iqPWyN2vlDmy/29wZqkv8f796O
B3Ebg//WlHrmQtcvqmqZhUwFZQI0whoaXrxHmlP9Odi4pNB4wiPMBJLX714ZavUo
PnQE1GKAwfYQNhpXuDomHpG0aqhS7O/WA9ej2wvimoWzkI2mfQq20wyufcim+QOq
uRjIgETpuxKFuAr4sGvXODOLRocT3mFRwU5e7qCl/HG77+JQukGQ4MGW0UArX5UD
HXai9yOuvIPw/jhClt+3R86+4OiBFVDUErootk1DM04ZhDmIBXjXC6qbpCm8Cu+Y
P5LGjyF0IVdCYYr4bkJn3eWH+ArS7pobQmmlwz1UdzLBJyboiCx7FLy3/1HPAGSB
Uzk1nJ72fVyPFT87KyFik8VeQAagfWkwb+mEQBif2UiHMHdE39K8CKiHjaqW3AOX
YnvJ7MNh+j7hT2Ji6hQxzI67cZeR7KD+Q+YOdwT3QC2tDOAKIWuzqol4LiJvO8e/
WcFx5zS3VygfBSCZEPlAQqoCEFRrfFFXWTY6+2lmq5pWbALsAsrxbpK0YK8aCIbR
yh0hoS3B7UeU6D6XRv7EKduuX0Rd2N4wgsYvnAuV92kOKLDdFxLxBiswqe5RFeyM
DuQkN1yDgOLtg1/4GIeBqXDNRw6IYYIekWCT3GdAvtSt4wzN8hZiDR2MOl7ckoxY
6onY81QArtX8rHlZ5JW3jVyHHB0IR1JzfssL8xvq1feu2r8byqNlOZq8PlXmwn1D
0ZEU69kslFwtcRqWwVxrngV592V3T6n9F1x+VW/InUIf3MmWX7lp7zoI2JvRCYB9
VDZFsrf4UcBUj0EhKwwe5Zac/01/fOyTiqnA1Crt8f2Wd1rlgmcguo2LuHOtGOJl
Yh8dTO+W3tPGn/uDEhFeGqNhwUCJ/UTj0J4ERP3BHwKMmBkLITJKkmY1w9KoL8aU
MDL9h9YsNq8nYMZFMuqd9e7d6PG+8Tr7FpP37bL2EoZRjZTpujheqFQU1+eKZtSj
5mcz705RUoiJi/4i3t8eq5Xg7C9KsflFGTxpHNdufWvx3A/Akdh56PPxGvHGhjqk
qQoUUTUzhn0rBMNb0XXQCrFDNSAMgxjra2lZ7tBcA/bXVi2tEqoh7ZLqT+OczHH9
5c+VvXB8tFkhRf1ltqnsKJ7DO3WpHuxGgaP5GrSLfv3BEJa9ZgqvAu94b1DuTjbb
7/7+kdRfsbKkUsVj9DVhAoZ5h8uTIo3YMKrB+6F7prH59Pr6UeOdJiYAd0gzu5eW
iWPRqXTranXTRUdcM2JwqW24nuI/qTO6C227/hx0RURgTlyVx5PbkdLF24MJvjNy
3RKXkzVRbYZ/4qNiL1eld2+0/VhzZ36iyGJUxrgQYFHEqCY8mnArvv2aXugk4aD+
soVdlCw2HkgJ5ymmxQp79bJS0sbaylSx+LP8JnfKYQuFWYuRfJabFdx8NaWq3kMn
l83tCKaqA93tojm30wnKYSMJu4EudvP7Td8DCoTaakh8Rm6jTWHRZxca7MCvqrNB
hNZ74DPCeicuc4N8bzp7XbGmvB1iVQh0FjwNQIQ4nw9H5Fep2o+CINSWT3lK+ozB
6VPHliZA8dagSwXKFBKi6A2PZdgVx2pLntyhHalQ89fypyoxnze58r4Hpr/u5Ult
QnLo/2j8U7DFH4Ku0pQTT+W0HxUMRCg/j3ZJo+l4ZvMhipEwZUecyZ2iDetY58qG
C5IXZ+UM7svnF4tueG2vTO5faIiXbiBrNLE7aH8uV88r/dfkKVqplRTu/MvkpdkU
5xISFff3SVKtRQxlIaMNcCoz4NxkxwTLUS0iygZeXmNBHD5tX1q/jjBbVo6lh8Fs
E+NIprc55QeRJ+Fg2gwU3gykVeoPWekOABOHJEVadD1Wbz26Gw+AlXZUt68+6d1B
Y4wAxiqCY0WelWyS7oDS/BAS4E6RTNZm/RnUHwHUIoHdM1PzQWKTdKwed2k3suW1
tGpWi8SKqDoojMTYxZ4E/y8BsCwQr3Gx9zJ3psjx+TvnhPk9927CqdpHEYW/xjf9
sSgYC+w1l/pkp8HP4MSk5u+Sm4NvPRUSYLjmc+DjOz8erm0N/nLPn/WC2Jsv5veE
/exrOlWJk/tTriTusKiuxzOkFsp1eRh9tOASjdjTOZDbq7GiFNNfpDgJjaY7olfV
qiGPHCaihnPVnhn5H8sol5BWNIK1tD1UioSD0D8h0UHrlR5zQN08x8ry0gVtQrlh
OJLQi/Df0WF5Jg1UULYEegkaFCRqqqoo7gCYhQ7Muw0mtMFWgy3VVRs/WMNpKJb+
ii2R8MSw+lM0kLT4U3krpMDRkP+ykDxm8bYGqiJcMdtODdYdfIKwuQF6WHqj9b6r
0V9cDAf6zen6h8wNNOm+rYfvlr93MMrIM/2jA4in8oLMCkdQiGPopBKpo1J7PsbM
F0tnMZ3guGIO0O+2sSXm/Vrs9WC5vNUYTquQBB+HYknaV3fQq1GeuPq45hAjFWCi
vtX6jYAGOCppKC+AqERFl9K02Sr293dNjg9zoWqz2/ttG577U/2XoAxFrZnnmylk
cLeET4ig3OR/tz5YTqCZ6bt8wsHHIn8Nzpvj/hEwqm59qHXDp8wZ4mOIxykVcuNi
W4b9kH4lhc/dqmWicBiUmXeE5ZArE2lWVCghPQXGxIPToAbyfT5ZZzpQ6KCNTAMC
3fHIbO19lQ7Iy3PM9xCBycqIONy9gfzR+NkNp2iOpQsIhWiH78qeEdRJgtD1b5ei
ShkfVbOpdTR1piBYimWdj2bQRfyqmHkoxfFK264n4kzl6Owh8HPH1x1qRD3rybA6
y1cUsPp+D47DTxOLSQSyoCcdpQ2J6c4iXmtVeCyWWiKDe1WGa3HNx7GvOLgZSJh9
vLMimpYUL3uGk4d9F70Y2F55mHiwNYRnNcmDG8hno4RZCx/uGRJTswVSqUMiEn+t
sRndK9Bovoot0AXPhg6CoWdvsyIty7LYSfPur0Qi0/pX7tCInpTZsdMGEkdPlYIH
8JgZ9VSWvOxQ19xc4wsQiaI/V6FGsSHMoVCmZNrbjxH3YZOxnbrxLkBXK8uJIE7I
xXlZMEg7frciDjbYq9HTLw702K/Ni26MA97uGGHDQSuFOXZZzEP0bvlEqAfDjF+w
4gjGMUOGP0DRKf4xjtV48LtnSHlPIXanVRBy/qvmL5wpO+QaHpKv6atps6PWcaDs
HWbdjaO0Ww52n/P4kwkr80vD+l2TDy1K1T4wlD1chPQbpHMgAHYnLQiYyUN7iHhJ
M5YbAvXWw7lTkTEVe0htDvryfAfIjFtl5RmTIeu3VliO90T2zhq81O10VAk1CjnE
M3xp3d9qS03bGT8pFPFBmLm8JMF0p0VNY8b6OmobFEtoEiLbs8t87pjsw6TtCHV3
0iJp4TtDLDOTJbcaPPK+GjhQUd//U9NDp9FRnzFxbKTuuM93slZLkMxRTcPaYLc0
DJB4EGuaOtAckydDD2OH/Ixu/eRx2fpPMzYel6+IiETGoik233y9YlVSFroS5N6J
dBJnnhWlEAAYuwF23YyGv9MtoFk2g5ZD8Hwr8HVWJAG8jHKooxZ8S0BnxI3PJ3uI
iKcsPKwm2DZopEJiHaWkwnOTM50kNqPO3YusH4aMGTvVi/NZvQB++E9RfuANL2lB
hyn9Fq9f0VAeFRY8GwypucSrn5jVRz4DwVDyocBHAdzmpLr6SZyltcu2M4GFbtyI
NFt602KYQKdTBVDQ8HP4TjSACu3sj00DlaStS2P0V61r6NlkPpudK2aVrz8fvgDw
UAwOeoFmV4/F87uPBerEsq/qRyOTUAegPl2roaaYg8s5QpHULTsloWiuyCy05PxQ
cmMADpV6onZ+0W3UwU/8rc2n5uT7Hzc+TwJikmUn7MpLBFkGZ2a2QMz91ioEH0XO
8oFnxk+kE7sPdCGniPBdLsssyZsWVK12WgM+6YdMacDd3zIppFHdcjZxArFV9tpl
0VwHlrvawshAjqmTXpTlKFJ5LvFxRyTs69g6lvm0w995GGC1dTwaI+n5EEzmr3Gw
XMIL8Ir/VjBPqMNnz4aOzNtyIkUtBXgFznJszCqKYGHrUKrF/9U0ELm274SMT9vS
onJ/vFDxxXMw3XaqJ5ycSFkvTZZub+TkPg0peD+Oqz1NVkA7/zndmSuueBaNFiOP
elwDVNE2eSWkJWG5p6dae4RZvBggjSW9BgaOp2fYB/b81CU4mNTLA49ukSRJGOuJ
+Jm/1RVLo44t++oVebb2i2A6yxyUe3xANJqIteQCchiCujEg5W/5dulcmUbZtsJk
6o8RnTzMryzje0lexXGQvNwvMfSvST1NpPR44wAoHhpFEk9BE7BeZEtXYFj/k/s6
rUxxVjz91rgyY8V1u0Kmw5mnBxr9vRJm7tdtsilzCpc0ZeDJDKD87B6P7ekNuUyR
G+38Lrm/qUv/qkLlRCk8vWcoNEE1iRVg4lxTKWPVU+ogpjpVJNfH1m/xfQd0aVUH
GS8EqP2RU1tAymOUJRdzKAt6VNDGCE47gx1mEUXJGKUyv7xAA5f7wQA0hk4T5Nwx
Ch/hrR66X1ID77QoGU4aeTjO1VcpWws26suqnSD3+qOOlHPKMmq27DxjpisirWtV
ZZBID/Bv3rZuKu1rHs6H0/sq7rzoWXeAyiVFraWPanLI5sHti0ihKxnVSS1VyDz5
pnh6VuC4ydT81hi7XSr7kZ/BSUBg2Uh2SVrmJNKLdnZJ97Ljql9jzjPhWjdH7bL3
ZCe+8bmm5nIDPadRZH409DPRNWT2Hw2UzJC15EQGNXdnvHglGJ7gCNxWM83vsFWd
V1CcDvXX+Mo8V+iZPuYRDbeTAtbbhv6ZWWrkNXncuUi+88SwjgUkF+HdC/MLOGX/
zYuus3ots4d3qTtoCqk5/J1vuVQZGvrAqFAZHWSjReV5Fm3xMaGX/IVo3rMCRCWl
UQJpTCLPLimrcz3GXcy7Sq+CwMM4Qt5jKp6dvHTQxbwo0fHNBHQ5m0K3qeGpQkPf
uKD3mIAJAAhwP8JBs6DyinuO/Rx89ChzGn6F6bNqNcM9KTxuCxPI2uTEXQLd5gtl
ih1IonfCCD7jVWc22ke+MDv8rPC60qztdMdo7vQt3QrmWu2IxiDqE3i8rrV8Zed+
ovBS+4ECGecW52WbABy58XCti+Xus39CN4NvR0Kpdk/LGRDFEYi+P7RrptMPVHWL
bOPjmjnUCh+p4xgMikIanV5Z6dtRM5kDbyVaa2DZlW2yl7IA0jM5J8uWZfUT+nq3
88n//CzFdV3MRTQBDKTSjLlblY92AMW16OPag+7DQRYWOzmj714Wmps9niVcEWnb
M9aVHQJUHb4xEfTIK525eqB+At0oWc9GvA5V5yGY2xwagh83vIUCQNexD9LhRyTL
NiHkF6OrcRJ74VdngR1WK7MMhtf+TCgewYmJe2QRTc2Ef6tWuKj0Z2HFnlAsRMpR
GuuZzWrCxYU9UtNEVFQ3qEkXt1UEcfmV6IaQY9oXxOJ0DJRZK8XJlcCgbR/yT32n
TDzujtznZWcnaQtIvQED9T4hmiUDDkXn3rwezJGaFnJqCBu7nGy81pLR8JtdDkvA
6WscFjPMSdpNi3YLZwgPSOP6IjebCv+3SKIr2sycwCG5nKXYOgGmC8y/JqDqTcnH
qcirI06nfNIbCiEBHYl/EJEgIfUFP70dC3TsezQkdvC9QUl3zeArY8FfoaFIkaD+
hWnM43AhfK59W7aMWO2g+0KHZ33wweIGgWJgBlS4lfEM3HUofTuv0h+lUFCUgCAV
2kysdhq7NE/npYUcJxN+FebwblNXmdSWt/jwEmH36F7sONh4rTCsKyNOJBii+iLB
3yDz38RPDbI9lDUceMPked7WirXtLQMjBwN/Ic7DdeKytTDFELHYzOjSSeiUILMh
pxD+wbIdW6m8xbGFFGKJwwDQjgLTBXvVoi+/gIjWmfl1wBy0s9BJ5/YlqecPmwyQ
SJOoPw3dDfgbiuiylX9X2FuC08hpetxy7K10mcGZngk3w5c8FwYmWfs8slkUWN5C
zQtYx4s4AhYVOBf9dV+GI5yLM0NgNzHKFdbgCBXyVnhfMFtImP+53Wav7lTb6u0N
tzhMIIm0Jx30uDsBC7FSn0mPetXGpAFIa2F6qkGWvhPSCDNauMMC8E9PdfmL94g0
qc1sluo6nOymIiBszQ5Ibb+Qo0ek5gwv0k9bdWNgXfXrwq4GJ+YrB7JGHWr7zMPr
FRp8UOIN2eZ05lNy0SwMh4lGcyjO1b2KOAWWWGwhHWewyNZa8q1hU5zkcSHpIuj3
KRLdowJx3DUVq0EURPBsosOaiqQaGridrbZNzProUhvk0D3GnKZbyokE3aeQ8WC7
lnU/HHmW/RuIfv+dFyfB7W4HlUJr46n4Nlzcd4U9nwKzH9Sq7/Zeo6DLjCixKHVQ
Q9tvBmTtwDfMntu91RZqR1uTcbAXp4cZvDQG/u6UYmc/wyl3sWe2odjGoUhRhVOw
FF/rL2IfXPCNp+asU3bwCyBs+SNL1PoELysKvgcZSkiexA0rH1bakYg+nNVJ8CI0
yS5qF4qG8zLOXDJfH8VpKwYMoxDL87/jArTaxuOSpwdQnrsGhi6SuEGYa78KFy9g
oYDVl25ZABQdC4+YEyWi40O/BsGvKLHXx/0J3uFAfqVQnZWRawBYJ2jrPafmwiSa
roqnu5Iy/BVeznglA/uEoEeBbPxcZ1GjGuvd1xhKQmXrkH2k5Dxde+88XF+YMykk
FxIjxdkUJfE4NLL4pVnPOLGacmoXhvrVn6oc2rDKOi7Xhv87fLXBp1onFIaWnuIQ
/+qFwX6V5LwYlMlUqNu+kJQuUenrJuYRYQYpfvTp+FCicnF7jenP/wX0K3Blek9i
F/4nUR/Ok3GLNe+4tXi3BLNtOBXFsS/WCfHCFie1boyKIgLnQDRd+mxBwAE5KYVA
cFfOuV21h5XaVMLUqo52GD9QzElfWO2qpUulIsPftOFrC9oKmrKf5Fb0YwOpviLC
tRG/fDgwdex76gjaaw1xNMd6xODTvx3Mblk1fJl3joh/ZjVe4LQEHNCLp/EhiU24
vswSg7URuilvA/iIbFz+JYOvwGDLyXX4kmBGXM4vtsS4+WVuAQkkywYDK2JBqbMu
3gmrswUYpBia+2/Jhz+9mXemR/1+waaDC22joaZ4yVYnvwRavOQ+pT4tvuM9KJAK
FTEbVxyUoDGlNwwaqZCJoUx98CTeQpz0FauD4wEcDAqPZQfbfkMuxzdScKF1MO+v
9KWb2A7yACFTyvENMCkjOs7yla0dzl56QGA+nWK/AnwIRBVJOlJBl9xly0oB4t1o
NizGP3SwWWewp7LKYUV2UnhxADRXSZttRF+fGWLg2exTAWVbaTDiEMbNBZXGmG/u
Cgkb4oevoT7pYLNzz4DNaGs2Qhdu5ZXp/iKdiA9wDIvo0mMESDFeLUxxr28GZPss
PNeY+R2JrI3+jzGwK4rMxksEKFtMVbaTm12sLmfKMuhalyum4UzXijU3Hx9mw9YM
MKNPOwbgXQTz/bRn3Lm4Xj88KCWHpHOk9xp7Pr8c3HzqgvZkmJoovWIvgodH8b38
7L1S400wwHZMO8llRCUMVQhB4keyhZ4TcY9xyq5lsi9+hogFFm2Z1FPgzZegGE+a
TEv4KMCOk6Vpl2FYm9kSqEz7hlZYkMkC8BffRqpHt9d2ZLcILSYeG/yLDI5vN5o4
Zt0RYjcHaWvfg4tHLrz9b7FkqrqW+zQBAPrjky/UIP+6xwi4UZz6lGWNePv5NRDD
lp4vm986sPMiF4quMU/FDMNtOgCYnlgg0Pn5gYS8B+WGMSf9OBRUnQKu5RghZMpz
qEVM74IB+3oDZC785n7irddZyIKM5uMluO2D2q2sqMu8LhdwO3EghssO7kW40n9m
u+jIcb1VLUsvDtviCAjZ98Gi2+eX3c5LKyIYVQFqfM0uSeIeAcnT2E2iQ8k8JdQY
kQSfWvUcEfMxfJqsyPiPhE12Az4IdyVop7e4ivXge0t0v7INaoqYJtd0MUrnp9Bc
rEYqCq6/Ir3F5IwGNvNnkjaIL+Ox40r8CnNjv/4/8jJcmevR9E45YiGwiBFGcSRF
SKQaYsSlU4ui1/eVnmNDfWkzKRigq+1xCI2N48cSKWIZdBqnkqVGYSPKsV/3dfam
mI2VLENkY3LuQ+4sr3AJRXraB3Iu7aG+ZrZuJR1xZcIatX7MUEJoGUYg88CLeUQX
V+PN6254dhtB4rfj2C6Q3oMP0eRzDfIinwBmqY/lhltnmvxhXG6FocUljbH6JdMn
AlyEnNtTcZTkIy43EjScGACBpOkO/i5hpZbvyZ0pce4sRXboyXsHOnW0U2K9OMXG
nRd1Lt2wD+EYW2qWmbEdOg9oU5ouUryub1dnG2RaX8/al3deCmlUGGOlH9YZrXCM
w9maTt/hA470Vwpe73wz8rKvUGvQtNf47qear6W861JayGgfjucnB7CIEvfy9Vkr
jZ8XMAY04mhJHjhvA5UMCLIyguYphTdzyNBaoMWUv6HxwY16H9Zspgsajexo34/R
g7FDI2Ges7/TbiB4APjBsfhchgYVuaxZWzyRdkOQYAPnpr2nR+AZT8iC9+o4ASh+
8JogeKmA+YRRGn7S9efnjmTIfOPzfkoSGGwnyFEAi6Baf+DfUanuGae1UdCrFOXu
u6wKWAXLLzcDl6efeNrlkg2I0lzSTiJ4bB2QALc2PwdLyUWbkY8BFOpzZBwcWr2j
axBZqyYH58nH3mhTQ2RYYD0m6Ja5vDobUasP/sjOpBcvNGqdKX5vFlGt1iXZhylL
yU8PsdwNjNddGg6CquBbvGTrEEEPT083rQ/9sbRgjecBaP6UCgmhtjQ7YVNdXvWB
olN+U5wLmaEsmjWfd3HSNPD2XXmmS3u2ykMCdTmc45bffAu3zuYMhCc9Nc9fDq+6
sUDoR5RYRVEkiS43Ke5eUEcMGEX65OmafrGw8xdP5m24VnNXKOOMe9cu8HuxK7GZ
Rt/6Zm+16bX9V9a31+RbvY3lNFU5s7NSr+nlWPg9wUD3f/HK3T7qRx7yu7y85i5B
eyjnyqveVUR1/Gl74JAQKywFqVNdVfzGa2FM5CmM82ZHYI58046y7y9qWRbvRmBC
daduoA5+Rl6vbR35lF7a3vG0AA7GQN1wIu3YouV9AnZ3P64gCfZAWna/qVDx1w++
4zin2E6KBjdhSu9d1IDRoFox2c9bARTvTA8NQydXy5yyNNiKoD0BA1+AAGXBFZmj
DuCmWekmAt+09HRlmM4cImu2T3RR2pfOi0uUC8ncE/S3KjOC8R0cGyA7gVLOd4Hj
WodO4UeABBON0vNGk6N7vnHmVATVU3rgy2WHoPaS1lEmbcxvQGe81Yvv6F5ZDR9J
Ud92CAXzuYQ6aWqH3PeGKXbGEajojv1PaFxnu5dHufmDUKVAVhl2shmb6ZbExEAA
f5JKaUQTu3fLqdAV1gN8NebEXRrBlY9Ulj8J26m+sJlCo8hCzrXnz+UloTwrR6W/
La7tR8gxxKO3OdqmKJY+pfjWW1hbWExh8lObiZBKtaXkXHZ1HXeBc98L84mcGvnY
X8UxUOW4Rjg72Z62G2Y/fRABOYKdEp9TY+K6JnzwgWbwlwFxFYinXvb29FvhnXqt
1sLEBeQyI4y+qjvUiokH353TYtNKJedXxc1VTpSOF0nqQQ1Tr4FOUABBLcvob3UZ
OgDqLJiax/OrrMOn1z50Q+r/+kWhTUI1p6D0zYIqAws4LYB2ftRyBBRH9vd5ByTQ
ILumUfMkSXGI4sSO137yrz/s5H9pW6qEdCkK/QUZF2/xPb3YFXLToKlGtY/N0rXL
v5OvE21mmkRrVkRH5Ts1qyROMMyJUrHOsOBgeFYZPM4w3Cg3HW5Yj7h8I3E5CAiw
qm1hMW9Vbrcdz0KaNkXYMSpGb1taLm6sriC1YxcFBUF+1yuS93mjPRnpkI1WC0Fd
qRFn3nUxjY2c/PdlnthjXgtrf5k1QWhCXYMFgtP4rGvDEnZwnMPfEHsphzISNOTZ
LHI4gKJqhG0T7Ul1DWe3JVNQJ9Qg0o2afAE9ppCRaSJyugxcsm8eQkGD/CReVZEj
gTmT/q+xPE7ubEXFYtj/hX6JE10dIbVGc9BUMX3hSPf3YjUu6usWBOfhBX+duz76
YxjX65GUq7adGqhEgRDHc99ZbdtZtjYP0Hv2Rq6N7J9X4YBsGsSi+vHP2yGqUNDk
pD6KaCVH2VL4PNrCYL582nf1sRtLRTHmS5ClmMj89/wys/dDnpX1BkWT8B44nZIg
GT/uk6RfTf5vd3OAIXTqR9xiuYH5ImLlnl1kbkNHpExqPGrzO6CY5/coPuXEBYFW
/C/UZ6vrnc/c5CYRWCLVtXlk/VQd1XrDyN+ogLtcZJcKxgb0AufqVn/23F7GJI0Z
GamQ8fT2iJ1Ms0kzbXunhd3pG2e7ZAQqroVz6hbv0NOCK80i3kBftHQwNevTVyHK
fF4yxAJAQaPFBUloDhCckXw0ADiypfPw8yNgV0nWae0uDt3X8+a/U5xcZE5dxfFf
BOzbfpZfNFQGhIvjcVqs2VAuWPEL/dnzAVhxjzB78Auq7dDDsel2NZ0EBdegcZwM
GV4qXExOYACJ1dw7cnfzh7wn0qTb3NxWNcNXrf5L+CRwB9lmNMnl+civ63yj8vxd
biFRJHtovYGMZzoBm+my6OoCCmCFe3BVmkJ/uPq+XPBaDA60N37LBmtfsBJieZtt
eJLpgckajYf1kDdb/dVztToiBFgAzamvrFGzc8B4AtHWR/j+Dj3/Ka264QKxKTPN
c3qRcbj23oxothJ1eBrF09kUownVXv0FLgq41z7QQa/3kbFK6hRY6Y+/Qg8NB7Ca
WCC0jIPRmZGm2C4PuII96PX7JuQvt6td5bSH4R7/SykHLsJx3kIgDsa7y6qcOMTZ
eo8umspZp49SHqQDoFdOXdeWaiyXAiHX1H2ewB9tU7/ZYVO/L7/p2/uuDxt/4kHE
Ae87kmnEiiTpaxLZa84fLdE+Ju2IJAwHH1YVdAe+qpyqVcd4gSFvll7eRT+O7tbZ
B5LXzbr6w4l+ZkV69eJc0WBI9zQsxTKXDQjkXvXbf+jTct7MeSEIw6CeKFqg0ucq
rVLppfVyfKqsckhCrSxk07+LkhcTTW4+RbwzIpWmS8hcQc9plTlUOtkjlopQe4YF
BP5w397ORoRytfyfHw1YooEbHtWn9nKE2fHkYkHh0VXIuab06lc1tPD1NhUrWVtk
TEuqNnfjZUKWgcIN1nrbw7JKaZSN+8Q9OljTmNzdBmLqD8po1m97mBY+FO2QU+kl
OkKo1yxD/M9icBbs7/XfzQWxAGfr+cE9voAxxLfNO8nrVDhbMZROjukkTB/4EPq/
XUvNbpWJx9Rf4ukgFUYwHPNSkrdOoYoSS1vNZ9h3hU5fLi0MKhJjJO4SRrMpVx4E
mnyw8B2MlKWCmqz/siVV0yhavWKySyjXheTQJ4mD4gEL5BwxgyGOqISla31JrNrL
PqFQb1MLKBuPBp7CElKmL4WXX62y+eommGz8oj0a+bPsfd3UUQMVe+mIBm0hgrVv
Kmv1SsK0mfLocale67+XBWSG8OCdQ0eK+ThcEKwRrM/mubOjNxsBWT8q4QLaSGLy
L2HuRWRbB+iFN/8wUDDnrJLcWYV4c3ki7w1KFLIAG+324KZJNcpEZiUHArAEzX1+
JHRLftoE+iRjnK8GWO15bsbIFvt6iVmXRby4uQKy/PTYZTGN+94H45PjTW9CBXvZ
hWOrSQP3jV9dwG4efx8CFo7Mrq31F+5mrLMfu9PlwTCqLbSFyJe9unNoaOqtEAwQ
SYzzj6Pggl+hLoUY9O9Fn9hEn8YW1uOYP+1Gm0LpKlw+kJDgpavbL/ByfX+LOPyl
AH+aPu7lkM+CxUobtqS7bVpVZSKsrUeoUN5NueSG06R+jJUPbD2nvO5IUpcW7Ybt
Pa/cDEGbAj9N9x54Lpwi1Q4Z4DWgh/zO6z5JoxVB5MXW9XopRhT5UHiob0S7Ajgd
OU9wYCPNzHMiws9DqdpeW8nkH6C2yx8mtRBCbhLOZ1sZ+Ae4QtWhgayJ3FJxmn6N
myMqszOpYs66YauHN/h4iWp3tcAcTSCEzlRA4YfcTcQOJhIzydfRibm4BR3BsRuN
qjpAu4sR0461M7dsegwKVjoVld4jMuG9H6dWtfTh61zvpvgOD2vYQAgsUwAGJL6b
RY6nWtciP4EM5615ofqKUuAeSLVvVqUuuhdysKPrAmuqV9woCtyKZaOIg7C6BgXe
U8fM0zxBk2wp+i4xA/xSnftq3PRp5kV7CHqnY/jJKFgXlkKZph+QQGksu6W3gdS6
KbgzbigFGg3Ya4coy443gbBt6ApnWLChbosUPIUNIK6RGSrUkFe190JcU9x/oyNO
FlgxEfpg3hUv6ZIH1CwSMw+2Ineav+aPJdhP+xmsRVY2+YvDvDYufLXqCs6w6LpZ
I8JYbqQQdPMT6j+co312Ft5t5KTDxn94h/TddCA7Zk8RjMgQBUEurxcwt53IMsaL
dlTgmdClvv/LfWwxCoETcXcj8raYo0ttnSPhTS8Bi+UIRqoMWELlc7d5m7giAWOZ
JJttNcznbLvnAiIoyKoGKFUEfVL7JbXOrokgNbOs3JC8p/im1l1Xe7h9EA6gvoOV
C/IYNf0mZzsPV2tzd2YcmZMZRS0Z7fzeh01ruf7FZiyqc6bKf0EZBgZxK0i4uS4W
lem9Tmk/q9qUhQr4/Nd1VSiGiJuZJ2aHcr8Web3EBO7+wF2SvhAzvxidj4Xncx8Q
Upme43zCxHioU8vh1JaGY0Mm9yzf3h45X6FKEKcbtFGFs+c7HIg+E7kWaR8d0qPu
BTqGWu1sghXJhN1/nOAEOKfF6NF8pEoWJRI+uZyThZR6rTaRKsQDbLAa9926WnF1
t6QYqq/L+fjGqXyeqnREkT2tGbPU6yOixthrVKVgWRTms5Np0rQGflxuW5fmVzrH
0FQiGsOW1EuX1n/8So0MfAf/casijNxLA6FHYF98Hy+3YVqQRdQ7oUxyocaYgx3o
jpORrxelffY3KsUQEJfmakrPNI7EfDwGvHiNT712MYHPuTCNPSMBrPdV9qzOWjpb
mWY3r6AdXEXgBFccGLdrEPTEStf1UltqhPt4bRmBQu3K8nUuVF7Aj5ICTB57fGgd
5n2GsJWaKi3hnXcn+pYi6t8Ul0KmnaXPuvAWWmuDzW+Y/YeHaQ5NWz7bSLPFlh8l
uctoJuozGpLLOLkbHP1E9qYxWDieCNLVG8bukuEkMJJn0wjqvQvIy3w0MIrqDVWI
bjkiRbYuMNe/t1iqjfX0b+L5x+CUlDxAuzfuSbYmrtPkj07Z6uYWkfwahVB/SIvK
FMblioaNM4atDFPw9PDJ+9fivFZ1ihafSwJe6uBnBiQVRqjRctWqse1RFPNNWio5
Ks/DCFxPPY4fNAYdcV7O4D07vado0mgmCHmI4eX7uV1PAYbmtCNrsezxh37OZ8YZ
J5M+GpimD+NnNtde6975S3Q/cQBrsulTY950pS59uMB/6vVProCbNMgf9bVn3+oG
kklocar1I8AHKD5JyrlI4LmyB5hxrYl3HhbAwT5B/s3494PZcpSLDVLf+Hs4F8iZ
j6xry1EMzke6x3rHmUxJiKFkp9fChYh/i2WUBMv4EehOGOOTSfIBJPMapt/L5c6N
0BVvgFtxHzLcnltyuLWoyzoCJ8USwJ0tbF6i9ab1vEVGBAwVxsyDDh550u/FmPmD
RF1nuLgyWrAvacj8pua3ezidoWc3MpPURnAZT4dlaay6rGrZ3qlLbt7GFwe/rHx8
vKkBYqKg5bnvXobxsU0f/Hf7KYeLKA/30mWvt+mqVPENza/c0ffGUY0j/OyhZCtr
pRx7AbepVoHgFFEvetqIex+Xii+aFxCqd/SOSxsDCFUdsQ+7YpB3LLS3yMYjk2CJ
Y+BhUhS30A63en7a59eKU31rkvCO0vEPEtldpQVHhXyWtBM9eOqZrmFQCUoiuqUe
z0cv6wbRu/HTmXaJQid0R2FiWocP0ta2wrbBEbaioRtmoXXoZCMbLAkoTKcvNbY9
zwNf2jo6fKPHOLkujyOXJ08Ht35xTyPugJC5xNgMwPab8fNv0Dhh6WqtCSyUxbqX
ReVNOnsuIHQOWgNCXGas0B36eAuMY+FqRON+1wnVKK9sJYZfO6e0Fxf5nP6aX4iR
z2zrGT10O/dTcK1Lf7ZuhXbzn6Jv7jEeXExOo5S2+ARrUWGH4UIqSKaAbehs+Dv3
qiWCzqIIaFsNeH/hqDf5ATLSMA+vN+T59S9fl5Xd6IUxCZrAYXM4D7R5GLIOcW/i
Yk6F/lXmwMxWCFxdQqxQDrzDA0hk3p9Zqdhv9t4cjwuWlF7t6wjWM0IVbYt7/GdK
xfVzQw9VD1EWvsO6HWCBP7qDFt9qSLZzDDp6hS0WdkOqhMS9QOfc6UKsCYq9pNYb
Bav59vj2GAZ5FEO4oQNnUy+p6hmWNjRo7GJzVa0D9SDWWIXzw3/a7wmkZAajPBV0
BKnf4HLsu5zcDj+gsebADf02fBob68T85b6XBmVwtvvZO66vABtNHh98j+t0Hcos
FqxhelcNf9S0M0+ofs6v6fAbFUeNYhIBls0OFJ8to6jX8H0bEKDFRRwrTu7jG7Cg
MDlxq76jLGJ5wiBqIDTiAJri9tgvURBoI+n2kKGhg3gocil+7hwD5Nzv2onXhliG
965tmm1+PCQ5eKn8UfIlgROTu52QOcHjjKPOH4Prs0GZ2JpXgFgLOiurxjdbnWGd
4HaDlJC5EeDaieg3SAVUbvCQGlaxIvF9iRxojgg9FnGjmLqVoW76DmP1O1y4dQ6f
vgpAAxGI5RpgCvOqp+k/bteGTmm01XomMSSqrk0Q+Y/2foJ7v3ShxpL17tG6jMZA
lCPpzgu7Jn+C3rKp1a/MQJmIgasVBvzNH4yQ1WmPeg84aIajQ6S9gNfL3/kBbJo4
TJUmIc6p3LXVfSWIBi3zdqbNylQxSGY0LNwoQ3DjvennXRYsWLlRZTNAaigh8pwC
wNs3Uqkuq32a7GSjLO9SE6pRjXUJmkd/3AODExhDFhqakkUuAVyuUh4eDtrKAsdD
RhhrjhLTlCsUihHG06Z+vqkcQ80hPOwWJLKbxGocQgX/jYv4QHb7moUAnRr/gqKd
aEyQgBHY+ovKtuCCVIdvbzEgPINy+FoW84JU/buaLpyWknN6E8hqFleVAqArl0v/
baDaUY2b/3Eitp/yxm7PzsUgUPD2l0utAMJm9zHvUdndsWeXaaD/9Az97sQix8L0
801rClUptPBEvhraYvtbKJDwxXOeG2qHKdcB/hW1Le2Kurba+yWmluQudP/HVC4u
N9+b/6XbMevWbdUloavuHytD7hqI0V9MBjwZoWTt2nVXj/33ethUIKAyZ6M+QVP+
bBfxTa8T3YF8WuBThYo2Fhu/b1qOM3g36VboqW/IAthkxsb7JvJwXlNR3qNmfAl/
DcT1QtaDfF3EOUrmtrE+XbEcQgg2wkivuafidupT0H+mDWqQ8JOL4Rt/4WgEnSvP
MIIBlCNhnQtEtkKb4GXpFPJ/uWkP9StnVlf8bAjVF3+fI5qRRhVhm5ZMmKr3gqwt
BYlSASxaI9Zou4bceTEUKpECoRYOHgJkv40xjt5g+aYegTws9+Z6JSjZtmTVtl77
DC7CREru9tb+awhi2dEvXeur36szjyfcLiz6H0cxfmml2zyo7rqG2+Geaxssgbel
HorkPASSiFT7I+NCZpjAFnWJbco3dqsYv6fjwZDZX8B04N4vRM/+VLxguM/+WQD4
PS7cl+Uoph98aIJFWzUI4wYHmYrpwhLQN9gUlgRmCllhtWTuw9U+uumF4AeLBScb
L9jgdW61JLUBWazsXNZEvzR1+LxDZQeHXrQZICc1Gj8m46UgprgQ9iSyCN2kanyd
B03fG24yTr4NSb+UdRF+gxA0ukDHkPsdnAYvOAfsEIN/zy+1muBysSxP5Iry+G9Z
SE+SkbE+6vbokXrIscBYVvlKPVoCwemrgWkJvqXiAr1CbZZj3IYZ21rc2z4xRs9W
fTt6A1sDcN5cDyID89b3TcMWGFgVkNSOgOhCPLo0+9Rls+IaCbmrQKhqV0uhum9o
aNKGMVauXZUHElm06QxWwM4e1RUy7+jjcX9xHwD2I3tgXvrGAQ8gMHwngD8Ba3Qs
xk8miDURcNmU9lPOhtvXtSJxQPOp+JIQhNqEpP25dwbiJQGTGpsPehHe/OPPxpRK
OhO9yghZfuwoPsNVPQI5moMdDz4ERuiOzRrwBdnllz4kXxjoZdJNEF2NiIoW1Jny
vT1gCXaPggKSG9wsRjzUhlSoLW6wgRxuAehf7XIYtZngxnOzAa4MprIaCdlf+vTQ
NADtKpkl6KkUzPy6w/9HBKpqSLwp1DvqWWRDss/wRfTyHe4sdhmb6EHbDLHcQJgN
HWzzNYGgbppFrO3Se/HzBd2LjJ5++d1cn0oAi55XHefmjKI1j3mm1OaoHCmWjWNV
URv/4cmVjOy4LtRacOvl+opLvPXAwWi+Mk7AVqi8WSSnlATS8g+ZIXK2/zD/WJVa
dQt85pAWiL+mIWorLrgMIguLDQf6WacI6kqkhDxC98akmE8TSWgr9wCPqTm918Jr
m700MsK/eTe+5JKVOdIY7lGEiW4/KlatyoLE0LPVm7N8msi9IrSGt7iz+TSsvIyw
P5Rlc0gIa/OmQ1GHmbM3N1cy47GpPWE5OD5TxRVy1T61e1JvKxBbkLBY+MCShOvt
d/rq+nPZLaEWYYUSGQjhtFuNClRzyqz+BMYttEyMuAXB44hUd0lA5ybuPquCYj9o
lEVG7G5L0cKv1KDFBFxh/U4euqs/Rf/Tct+letmV6Gx/GuAhz04DoJ90bOMOParw
QCtaxzcXnEk5KsHs4qIObDmCG/u+XQ1nmLt030AQIwvNDpqGUmeFKlZyriwa+Xb1
nUvyScUdP/CaD2TundMlu76/u48ZOEr7EnPJ+MAcuMTqRwy6i0iDo84aWDXft8Jv
v5wA5pLNle9+QvsbcAHE5nAw0SUfPU8oLW21HtSYeJu90u0a55zWkTxe+ejVUsLg
S6Do2OZOlTeUH1yWIJDjAR2GVO5z58EPA72Bx4LpiW8bveBf1l/lBVEWIpotwpXd
3DV+Rz0LxsgquBxmMfAZHNc9LUo6psshaZTZ26tdIQDjBYBbU/AM4tu/vjF00vVu
op1hcD2mNwPhhASt7U1wdIPKt2zv6ugVlIIM+AM9AGEUwSAijrH9EpQ9QNOw3PJX
nZcU5cMCKfjB1mcnBA7R6OTb+ijIy3diJWxTUHI86xbUkFQH0SXZcmGf8qgp/RzU
dP9QxiGuPx/zIxu8xC1WaMnORz4UPTitCdzqytfSEJWpt7X4Pugw50O0TQHVsb2r
Zsah3kyWHJG4DyNeu9rLrIGbyM5YXZLvdc6Iz+mOjJZGDBCXjDG58/+QTVqykGx/
17+JVRCdkYUYB9Y4f5GCtQFz9f5YM+/colcEfg/sIvjf+SdI7cDItmYXB/28rTfX
2RfxUdmisKy8Mf+Tunp+U7furg9a2sOxSruH3RreySHc6qyMu3bWW+rnxjMYtX3C
Rg3QREIo6eZVv6V7REtrlsPV0c/9bpt4fq5De2QSv7MnHp11+kWwSl5SM40F5X9h
GEFL7RnakF16H5yTvQlZvJ5Qaod35cm7Ogj3b1K5e8Q6yeiyzAnfOIeDkaf2i5Q7
IXRRCOvOCXXb+W2u3chjyCwxJhwcQ5Tvuv40gmYFHM6MMLu3NEOXL9RiNYOUvJPE
bDdtddcuDzIWQAh1an1Twci23uBaNOYKdQV76JS2o8A+48cMgCO/iCy4HgqcENOb
DL1w+aBxGQ9F7FKQfAC8c5oSYiSTDVHyHA8bmmWO04OpuDtPRQBsPHmV7cNdFkUz
LFRk4kTSO559IqaH8mAcu3cHt/lH43s/gXcd86Ugt+qz38xLi7pcWWzcrDFxrKXh
W4mZv/fwRGkhkg1OtMzmIvpfLv82T6zRXHp31rlew2O5eKzsay9gSwIxZYk2J7t8
BQ95+yG3fZ1F0/XGPZFe3Aw1nAAnywIuet3uJz6hDItS6lUtTTT2T4kTur+yooRf
AbXEHE77wrkLnVlDqDOrSNQR4iw2MUk8Z33cfU+kyoE9YU5QuJElAsP80RI67qOl
oCChJv+FtWDXwR9mzfVCyYg4Q98ep/1MO1NfJus29lqA2x4YQQDYdmGG78jK8a6V
RNDxGNxEhjBXTcZgnKjXgvajrOInTp9k56S1WWUHMRO666DuS9BY4BEs3Z4xn4/J
gT1xg5QSJqtVRZrIDV5XYD4hIpo886LrLyC6bjg6wEptuyd7DAOgCoUMe99EPaaT
H4ffw+WU/z2E9xNi7MnSQE7xLhP9B55/7+2YtVw/92629yLLtISx0NVPm0GwQ81x
U4jRpchQ8ZqnPCDQst72N5cOPanXTTYleug5pQILq60/DRkG0fKjNn4hDi8QTH0J
Gmbz2RoW3QSatYJNuIvhh8ZuG6b2YBS0pHgRjuetlR/hwUfN/PS6NUqCzZrKfai7
Vla8MhG+os5+lejo7d1AlzuDUfg4YNk8AF8+uXFewQ4Q9IMLLwVfeZ9p52NMPTPu
LE8QkXBXk/it36fjlzpvPAo8pJcR8QYUwQqoq3t2xlp3YTv1xM6ffdzzyVR8iaiz
nXUGluSlNA0c1Sa2ooVI4x9bMnzs/bG1Mew4Tapn6UdhLDQrER0i4yKTmKQxyzvT
DT7Gdmou0xWRqVIZ9Z1mLmZFcd66EtYuGUtHOOJhAqSOWBaPczVOOQRzbBySHAM2
YAZb/1I6HsdRhocN1smfumH7+drbBD1ciOWI6g+k9NM0/b3rq6jKDYVxwfJQnTdm
Ts7+NmEsKPT8xRqgOQAGYD3MIbCHP0Lmfbt410XoVa1SvSbSTcfuyeQCZsdQuM6F
TfzNg6ZGzoBMp8u5/1ZFgBEKvX6xVDrpS691H0wJK/xTElsUGO0fJt2jk9cLSjDE
s8Lv8bozwkcUrob/PjaKlXZdt9ZDqWy8J4CnswrDzBq6Tujo8NjMwAA7BGFpv8b5
AGAYMbRWL8ne4haRnSLTYE4sGdeuxhpGQwIDrhhQm6zGOTIpnI0tbi2zBMvzjh/q
xpNvggantal4ojCKBPOhXOPqJ1LwXQyJaKNlUocSEP3K84TLWuGP4kox29pVWo7F
S99Kv89kt9zwcAFjZpkR0rNlOdEJI0iNeqFI515wme/6x3q7Yi1u837SYHK1Npmp
q86vUJOT1tKiaY1wTdop6ILlGkjlwLdRxo05yJ0CK76XjbB7hzYX58vJo41JtZNW
Le3g6auT1gizf5nLclfohY1KjP1ESoHO+zXbfYDXeb+3DL5NxY8oVc4BR5IrgDry
c4t/r1jBML1B0gGf4QeChqkEhYMnHOUmxohCFtX1GIxJh+nEKGagnH00/lZgKnNM
SP0stEvBc2SP5vcJIMLUsGZbEFgvDy1cSVJ8K9tpnOWxpOTJq2cAZDXk6aI8IPFJ
ZLm0TtRkuerhi4LRtZNZ93i9krTvbIeTF6biYIDHhy1a6X8jWmHz0zl5Hy6EdeiA
Xos3WAK3lfT7G+XGD6tvG3Zw1Xaqpt0JxC7WMy9B9C8HWetxUzuxIvTCXhB6WKLY
yQjeiULYuV42npcIIZWhmAWtz612mdGiuh0uLgVk9Y7QfO/ztuVjl+zI4nkWKCFN
iJwlqiBG8nwIYN5GHyORX9OyVIR/tlUwUdGXxfIM43mNuSvefhhO8VRc0Tve43ua
hzoXUDFp8TFgdHfNDlhltmADETaYfaBt0azxgbVaJJI/5Vz7be8FqN1Z8TxeW2Sx
R+dTyYk2fWIkRqbVp5bhAv+7sMSnn+9+7RnYVXyuoxDmfk77pxwV/FxGCXmJRJ4L
4k8xrmO0cQWPLctbYRQn53t0gEpkBMtde0K8zkWHxhZ+sbcTN26IA75rJmmjkW25
e6JlPqFlgthkqXbC+1xAOOAUujEMqxSyJjIoY2dCPPfdrKPtAPwtANZjOm4pKVl6
nZwWV9qH9QO4SlW+dNkgIoR/5goHsV6QPO8qO+1es9EcWPJ8ggPqZkzuP+CseKgA
oFuqwnfDyCY4I8ISWTlCYJyeWpGFO6RqosBV/eCToe5zj9XIM+/8RF5JeVTojfeH
qL2otBCEC3M6Opd2XZTJnEGlx/HdJIpjT2+nxp2z682GDRTF/tFvG8RA4ff36JKf
eDE6NuEBKFlVK0jZjvvJAwOrLELQKNQBHVGmBUARVtdoER4GOeT9JVE6P6Mwx4sW
IWrWuQCjjQ94LRi1JZLabBJy6tTjCO12kw3dG9HB3J7P2dptrGuHUugHl/l1QkNI
6nIIH8i157veEPER3nFT5ZKbD6FufyWnGUl8lj+o5zFJZrWH0IlX1i79AFFtrc+i
8ohljen959gBX1cSMut76ph76L8mJp0g6cENrnZ9K8yGgQ8ULFtrl/xZZ8XkAkNh
Qy9SrYDnkPOBOcffx/RNVqVU9kPG4ebd02yQ8TV/piAMk/fd868OG2npqKpSmj4j
cVS9JMUL9HKLkJID7Hoe9j7UeFZsbmD98t/sAKKuz9maMFiaqUBP43NmxQoIxNDU
9pNXky6A832HDc5Vv3/4jy9DbP5gCjr6cfh7zN3N8hoBFNgsoBU9FAi/uGFX9j+A
ynHcpWo6BIGF5llLimWuh6t5sAlRJbbXmOi6Tgxqf18CmcDir3mtDIvVdsxk7eVM
wR1SOwvY+m0Z/oMzoo2Dco62GeumjUBGBURA87v31b4vgJKd3orVYxxuE42rTR2f
XvLZx80lRQeOPZeX6lttr2GF2Vft0uNp6M3KQ4QDVduRk8MdFrb8oX4p6A1DvLQW
ZB6XnKknVEQ3SX+WrN+X0vE9iyhvEI6BdpJZdjYhbSadBfPZO8MMCEGEDfsLle+d
DPmIgexdUFW0jApg7AsEEIe2nyyKwNw+gxmxfik+j0gYk59f3JPARwMuy0aOX7zu
ugSCryPsOCusg9MXZZIM3gaXQs56Miw4M1wKDC8OY+sJgHqu4WJonpRScOfYNpQK
+ibx0guqhriLYPWgEvWvhRYUdKrD7KIkSe8U4CjRPev59nzCJmeFZnolAep7GXbu
uM/lCm52czbi6H/aQg/nmrJciMEKZHsQr+BX9X7oEOKOzfOoMkFppP24MdENYHzR
0xMiKGNTLcsP8bfLFHX1ZdXcVMlkpJWgT0djjt9w5FZHYn7toAyg8TVDZRQuzi3J
q/bDGTUFM4aoh67DJfmq3A56OWfUECiweTaRGDmHPevOwYkvZ3hOafl0W8W+xE96
8lIG1nQCUe0W/xuKoLIfjDAJblNIlzED6KiWXWLDO2cl2x/pdYF3hr+Dz/8vY2/5
1o3l5fJSaEQhYLUeYZtJj+rz0Xzl/sZDKjayVVxdTxt3hzcz3/ZkpJoobQJkH9NX
ajPmeLZjcZ3dh625vOMuYlhubt7psEc+rz1eFBGh1zPNFKrtt33D0N7jmxRiZlPd
SVUf2+orA9RGO0otSER7xqTgir6a/nJVBihGz422Y7gCdZitluTpAfOdTKGaixGZ
4rHh4kSLHxzLir9GfuskxeZNzekDoVMnpU4z8PIKJ3gyYFfpniva3+NmLGFKWmBK
7B53bs8Nh0XuflDo9rG5MgqWTD0N5A6jFaac0ShOUf0W3wTCCwf46KJ9IQrDpxGW
O1Wg16LvvZO3/7sYFXvPwdyyQQySzAwxWA93zALIyCQLKZxMA/iZqKisGj6RnUff
IMTksqBxka2+QBy1YsUQCFd6lY+av1BnHyW6vax7z9N8ks3U4LeUoi0Pb9sv4VGB
awUMTWjYff62XcGMgW5SGCRVX9Ea0k0Gfik2+zX7dmFLcWsmQiYXEgLDhIYr0sEa
6eFAAmHvT4nqSsO5dcTHz/srWgeviyMqTI4idSfaQ50pTh5USybnVE0dSTD1Ce8S
wSKWYkg6JVtpCoPrTE4yj+drodiuocy6X8Sv84n0Pp9Gvjy95T0lkzGdcF3c6cMg
+bOYcKUuNAKNecjlrZJRMeBeRjbNiVHUu45lQNtRVN5EhMhHtdaFKNeBxJVHViJ2
ar4V2Nek92xf34luAPocyFfwQMQzyvCC9MGSsDK9mYWNLtIWfvFr8r/4WseZDoP5
phLyL+8S7RHBTigOBxdGqvlLhSzxTDVrx+hUT6PWGFN08Ws6yIR6YkPcmYC+Yxng
2uL9QCCLhJBulgoPSBEhiEqQRuOPmoAjJ4iCXtluWneeOtaBRUVGnJiNAR1OaM8s
qhWvmaMrpqDThjOJ47JRKX5B+lumQVkxrhG42ZZIrceDKZGy0I9NU94LrTK0d62e
5dkIx8+aieSkKtutPLkc5aWVoVjZKZASuSz/PQUetucjj22L0gJBCD3hGL8pLrqN
DVtcp0o0A+Q90KD72+jZVJjzALc4nvNFpmwumKMMYUxjXCQasshm4EDb9GAPGltE
15k++6x2vwppMF+94VtFu0sNvpDpUjglw+SxZkY/1DKqeiKWClatahx/KxcDdDv5
0w5ekmlmbk8koTdQ8GTrVvi9eFr8gb2UlH/DFFoo6h2n/ytbWtqG59Bd/s3O7RfK
4zm3gJ09t2lur1iVN91Qax+jN52gOMgA3F8YP1YOVUNxFwcBMPToPYMEi9SklPFC
vQKjWvsuBmHUdWjhR1nTNDa7qW0nxGo7ghMhfsORnVMxJ3VoyTIt6FnjiG5oZB9c
2FW8B8sd81b33J5wnZCd/h2BoNh0+aCCOJ3tGn7ypqd0WjhKiyN1UN1DvPbhj0rc
kR3A6XVDsolDvlxBLIrVuZ6jpi6z6We3oHNW/ageeQOzLwXbRTWgISKACQ33XR05
excDPBwIl5c5O5cicUb/EqhA4ehqzwxDnczF6zj1oCdM8+hh5W7hZtUW6KKJ/CHi
SSQCmPjnFU49Q6hDunCC+zib10RQgGhkTuBKvdhct8ckwwNWP+LoVU/g7IW0JHB0
w9d7ym1j2usbJyS1M9Dp2HeTfsbmJSlzpryq5QfHcL+Mm/9Fd7e3LVzICAEzJKBk
z4o5tq+iBIGgrLD6Cfhd2lsOa5Iv82vvjfnxg7ulWKwPYc/cZaGGy6q2i94UKC6v
Ca43Hah3kIqqPmc8X90YTAlAcwUmdXjbA/dJ8oTmmJ3gmK/8TTdoIs+MnRQD3V6J
jXyMUgm4vmf6LwNcpJRZ/nrP6Xoxf8W+yp0qnYJqepp8HiZSCVj3AsoM8yEv4zY3
gsz6+MPFlax+MmuDQH/MUu3iysDsuFcSlcWW+I0R9XbDiQDGseDBbWZqp/PNpaRv
EwCzPbWyjqW9TCC4La+Ps6dd0ZKxphXV3dk+vQz4VTcGt/3wnU0ip02UDyqvQhiZ
/SYONnf3wmch6aMh8+mXdYC1GjkmH/CxP0kxqHTXt148/BYu13TF3PAIXylrFJ5z
ewEbfk3b4QwRFxymZ/l0NiiMaUHcZXi7JenOtsqJJ1CvzRGY6qMf3lOgD6uqdNbD
TA8dQtxC2HrSa3/4FTUVQlyuNCGkoHSe0m4hdEAHq77mz3UqpuYOKvZ+IU+bgdhD
XhCDchAghmFhWy89VEzb3Ni3+XHoZnbjzMbyPqnHjtWJ35CA7xex7UBiKvYriueN
zLuiG32GtPejvs8ikAAJ7XkcTSzQVxMyPpNuapm6jY0/MPt2V6PAvQxc5G41ohxc
GztITR+0MCl7H5ZsqQPzBs8r5ox4nvnUUOwRjktJh+1PMSBPfKhex+Vh1O3ZqeKU
Xvn1IBGI6tkwUQ0dosIuHZLs+S9L3qqypXXQZrZ6vwnLzkUMnomrxSezcnUU/3Mj
pExhNr54KJSLLI/MzmN47/FkbhvVfOsgA4fblSoU+yLIVIcYLNTP2vVboWyAyqA8
5T+q0h98St1jSMR9Kf6c8RYnJ0hp3Fb1tFCPrkPeOSuvA+8yRWB/uyNdZ0/ePFSa
RRhJo7OWjno9iGAPYbOWYqri6h6N48Ox1rD+LdlkzR/BmNsZjhDOGnO19SRSOuMe
HC1U5TQIo8dQ76ZjDOfsEAFg2+pqOdhzM77naDks/xbj6JDTrSowEhgP9JHj0c4k
D/k9bd1sE3+tSCe+cDzKXLJxiZO3FkZyDLYNnOdEgOgNTJFFAFhowYcc4IAZB1I5
s7zWyQk2WzKAlA3foovOA/+X3ijEQpwtbJFcJVpxCAwK2SOY22j0PinzZZ2qOrUz
YvB8DDipubRcWgIFUEEQkNIp0SzuYr6pFI3h/QFkwqYTxbfY77Xud7Xc/+7mnk6A
PwDqdrPlhlJgsoNyCTiusTestWDF7hBu5IiKONi2n3jdevi7Yh8s7OJw0bLYezjx
VoMwyl68AWmIciHSLgExQcKHYR1vog4bYusT0QQwjbYmFRpNWqGRIKP/S5Tt+TiN
gUO5LQoFCeB/qIUBvNpLi4x101+AEM3Iv+vyravldaRhc0t2qP7R4lV0lRSh6Mr7
VOmAxuyB4JrDYxw7z42ZG91vDBSFuwsru7M5uPByF1Y5rvaf3ab043mfa2OBkKT+
2+C6dFLmvu0Kn66wGEnnjbDl4ws1DV2zb1eL9qzGV3E1/DUngb5AO3oYJVO2DrQ4
VvNAVLE3UymkY0g6ErkTD+eCr9nV62IGh9vIRX+EQrMIT9hlFDAlb71BfvXzN/1W
G0vHhYFe1mrCS/vOAaJZnWtvHcAH3TDpyvXdTF9M56aSi36PkbLm6I5xu/eO6fO4
MH77YM7CxaGw/mmZPHBmD9MhYXCLZd7bs4fHRB7oFLrJR40bBsz1qxoiBO9pqtoz
74bzg3tn8lOqW/Th3it/QEosCa1plNTKamYmwxZFdC9INJsXnwzwy4MvwCeryQms
f1Qvz0gwe0BdNPX1qXRPE114MAyaGK0bgIkb1VSczzgLOuNnTCNAAAb+wo2CqacK
Ums/y6lB6FS3z/K+vtRKdkK0Hi/DdV7ATstFrwiIyJfc9orn/nk20s/WWbIzobGj
QAhdUDzPn/rHzPIO4FsbkLBvZytbi7bveJ4uJsHNbb4lJuPhNrjSGjiRVzojCQUZ
nbIE4OIufABgPrBts3pSbqHMOyWWjBE2wxjUrqlZ97VZM9CMiZOmQHDIZLrDUgY9
atNlAeWIW6KC46/goLSv/KUxhIPEhf8IDsVHjphfRkTJG2YvWc/1fa2hcr7I95Sz
RgJktdfstGCKPhmN3bMvhOBCR3fqxV/Om9j8zSI6uacJ8WUc/Gfxtu5dIe142ZLq
g1ntPqwxrPQlQKbblY7Q0/x3GVrf0G4nDuVI0hOitThkFdvTMvA3R5TEKFLQ9Y1K
PUHuOqLhZNWbWxy12x/wcKGUUt+ZcEZdNnkhdw4p/T6o/18oYVW9Yt7oQiurBAXI
NWF+efvWWbvNM8b3DU8KrUsUhRw0m3HYuMpJAZZfg8UynJp7V/wjZ6fAVvQIKb0s
RBrDeyixZz3uSHZf0KFgpT/RAtBEoYJDuqPXEU/CfeXIj2ZnUgasNMDRKHYLgK/X
PIbTDOXxyifBarGwBc/DeJDDDmHIEej1KAFeitFUUy03CfULAdOXxymF374J2sR1
IQT3kf5vnuF5DNPOAzgTXmbol08Oqb6hfRZ6lBwJqbqVBJU7ZaVX650mI9ecArHz
bH/FQ2PxU8UTaESPdlwek1w2YiZ2noVOHUikzF/7Wmdv69OsI8Kj6YJdxfseIBpi
B4MVMAJdATuHGd75XBpM7tb9BpAsne0foMYYC+kPEkm+tcBWvDyVEcjnEMK6cEex
h38c+QHjTP5k6vKymU/aLnlqIDE051WQI0BJCueRcW4leUvPAKIC/XA3Rln32pX1
a8PBghqkRFmVwSx7Q8U8GYXtu21Vdl39ckEYNzB8oezgY5bOPmrFzU1id064l8ZU
9y+SPfwJMzvOLNmqdMVpCK4ub4rTtbewBH8ZC4Ro2SpsJbHHi6DbBaMfF43b3VGM
LckJl5bn9j1WRisQFkKgKi8VSvewSVpM8j47N+pPuUcnXI19Vnt4Kg532Jf8fQR/
C2OKdbgXW4defzSGkk8YBCR3zJxQjxFmDM1GNSGZm0TsgANLgp5wfZPKz2bHaPxY
Xf/b4kIcNEyzXaENCs1XWXhlAXkKZD0aHiT+7sTj3r9hy4xKgtArTLxy6E6G+x+9
j+CYVn8NSwd9QX8gwSLde0/7Dz1MBPwfbe/f+/vvj/R/1A1Paf/nbigLXhxTF7rN
p74Y32UmiHXDSl03QhRZn9Fm0OUNs8n0VZOBmXgEa+25gRZso3jfXjrDGhOE95Ug
AON6ZMYenGuwsUCLMvPVSgeYMx9ntSjx/tmxoWINFtApgrQ5fth2YWn4jtBqwpSd
yarna2RXoNCfHeVRQe71zf/1Ebo0RwZruabbFQV2b1RQ1GRCGgqn43G0TrtgFn74
0KMP8oz7HcjkLLAxENlJ3bopnYDOCTEpu3YgiIaoiUr9N/eBekHwRnSSWfQpxCCt
p5i/U+CRcunexFmSkgsPjiJE7GPYmdeii0oj7xDVEf1YULfmwYKyuZm3NhHuMmlC
u1WycK0mH6aeU3cRWVy8ELgEdqW7LrE+vTI/jNLX7qorDSELT0J33NMyEoLBNmeA
erdRWzRBN/VFVufSYSLiqnARO5os+yfv3XH7QJD9VGQ8uzTyAUil8N2T56ocRaou
gVgp0FIyTmmxlX3pfB4IE04EIl1RYMVLjkMAovORZ4H08t1ZjV/7qTP5+X/Bgxio
p5ZX6ExSA8w0H0oR0x3MlB9xAwWjr5xxFTfToqqeGp4y6tlnyqYkUK7xK785R/FG
zt0mdpBv8lVyWRJtZnQErYEEIn28qMnjFutOCn3O7qNeEw92Cs6W7KGfBuvkX8nT
OhpEO+iuNM9DFUX401THinYAocBGfUm2k0ETk1QSOvMjr60RUFmi7hvBiK8gDZPe
acSNJh72hCRkz3awstRURR4MCQqR/O59lmojw/KRgVHYJ1wPfy4CxE593W59jbiq
2SLKuCKULd61pUfxv+sRUiozHv/hZIqueTSlyNWdaaw6+T+7o9lkdct4UtIvkiMy
A9HuAmxnUW79ij3Yp+T40Ao9Q6+/cSTSWwhpoqCJj3kmpOv6DLd/knVYnGyegF/6
x3AXWCein7lcvoutTZhyDWpJlgCftz+gx7C3QvNy82yCUVvrLZ+fJ+HedjPXLMWa
DuFfgo9Z9dyNNsaIuihktF7NiexvZbhg/MZVx/kQclqVL3UT5RzPNZbGq7RNm4Vy
fWg51rsNV7Hvg60WbzGKLEaFSFBOjAJcMp15td/YXzGVPQZQSLTUbQDBabGTa0YI
xc7tuexdEPVGShNN9VVS7A5Fb/PBosKMwwtd7AscdoWJ5t+PgWqpiMPo7kzz/jbT
cn+LSKNbh+lSY2mh3bWzrjvGKnr59acEmQxR3B1we3CUBwUdPUYgJs315GbnpOx8
2xPD5GoZgFdjBxw2tfbLuN8DdwDuxdGkD4XfKnAcwfbn955MylkDN4AwG4cJ+5Ef
Ge/SsWNf8npGIrBXaF3FA8vEYUiYx4xflLi0AXEOopvdTfu6woAGhKqRabj/8JBE
sFF8dOBLfv8nAXrEcOjCosx/ybmwOxO2HcfhzgTIubwsAHCXwXYAGLMMbVe1Kje+
zSONcV4SQ78Ce+oTMkpXrjoUl3mAF8WYcNBlhsAJ9v+vnoJ1myk73pBuef6goUE3
jY0gMpDUpiawaLZQUsO/dFJ2Mp4B3SLjRfoR8dL8EzDAjnYgz8uF+3MyFOsZWHWf
FtGzOf9b1e8Ze49L3dlPZ1tfXUudyrRbcimBweK/F9rPIcjfbNEWVC5j1sEIy1ot
1mTRkXeM2EWZix4ORgwqf2kLp4tdFhn2afa37CWRH6wXPTWZVAjX8RGpS+67gjSv
ygfbbVYrjmBEwX8CSMBbM1+eBgUCQtUj7P2VAmCAldQSbfrE3ZQrnetdzscyepUk
3x8TZzA7lZ1R0Pu3Kf7+4VxWgC3Va81jLOIGW1X8zTYsI3pZJmuJ/ha1OK2lsZHP
F62bjk4PNk3o3XLouvkt1F5Ng38V15/aJ7gBDe/t4vXjC0GpXzrjt56bu8DuAdlv
4ty1UfuqfZvS9EZWNrikUiDGBGTfqFQpo0wRo0ZufsbOVoaovuV6GnXuuGoKFhca
dC8Ypng6vfD5LrDwwTdxgJHqtTcx5REFLwZSuaDZ1NVplEvEkpYu1HYq9Pp/5T+L
6PmvgyCoho7D6vRK5eoH1AnkFGiFTchjz/Yl2apStKWlpUNIjNaT/utbV92dANub
7jLtJ8syYt6nKpJ/iP12UUHkBEG/Fl0169N7i8Tk3odW3+7SmPAOu3J6l5HciQEG
0UT+74Kq4HjxqzVNx1OPEJ9YtajpD4NG4M6u4v8/5HwUtK/QtFuJvT6l3WbUTmIM
coR63eGxN2ev3kR+5QgykbUqCMfScKCRckv5clSoh9Xjl0A0+mrcr5nvkAN7+hDd
ScYdL7BdTw0hJKW16Ktr5WmD3oixBSK4IZffVgv678pPVwRwDkkvlxHAgGfCeVaM
k1nSou1iAD/yS20LCuxLB+QCU5rSAblDWNa61v3ssZ7uVyoB+oO8R/nXFXi115YF
AKS2646oyl+JdpxtP7NfGYNLFmfYvkSVRCdBt6V3MECxlJoYw+uniHsWKy5dFJGZ
/+GVCGhSOfikOzKCKbJ9j1vjG4vFgnfNxBd9v+s9qV0qJZTdazan/MTVdN+6pVZc
9zqqlFnEKEnEQU3SQs8Id04eXiHlmXrqvISGaQx5h1boQ3Z5wpqOuc9p9HyiAqVu
wMi7gGXZQFhoeuf8hz10IB9sdROb3SWLBvRP+2POA/FX54qmOIiaAy+Ngrh/kbGT
PstzPCEfTnKhpifQunYR8TaB4jsanZcfZ0+IUtZ2Cef/CtREXng4iiBav67rhPcG
jJbw/ZzOrtBC3St27meXE+lpQaf3vRFiWNAIwhakhu4vG4XnAaUSarzuRDiV7y8E
GtWQdc6ksuVF5fSbrIGZV9SFSVWoEre/0TfANcJVl/f/JDjOlkV6EEQV49/moP9p
D/2EeCG5DewtDjEHgjkBEJ0GjPQl5U0Rv1qEnQIwezolku794UcxLZSXeJci+tA0
Xr9FOzYKIib05d+orxiZgC6v4lCeAZscIBjvLl0X97m/da3efCWUr8XAGoX8+Hcn
zwjOBMExY2Y7HFSVpFXGV2cjBL5DX3CyR4Ckl04InzbOSSDsA96uanDGwCAEXLKf
e6rMOzDi3R7scmBkPuAStyVEDZWsVBd/UY2Mb+TX+U1zpjx9Rckmp6VpeX623pEy
URMGKOs9yWNOZn2N4K7nM9vYSZWQqb7Y4jEZZS4VDu3iWTGnHcHrt+XGbM3Lv+kV
d4p040/vLtCyG4eql84zhKG7hnnb/Nhe4zRmEQeOT9gRdi0O75/QC81FF8pc8CcT
9lOdjwa2b7cY+wpLFGBEFok6YSXUCjQjw8ZWDmRcfKeYpvMu8kG7RuxOyDvDOQJy
5+Xj8C32N2+bU7ZTGaghN1w+8Zx//tDwPa2KwujI5mfd8fiYnN0d0u0NDFxIv8tM
ea2nOzUJ0AOyGR2EcXKei1FiNExZAkRQisNGTYx7eypjuCzOvYwvT4Cew6Wkj9M/
nuGJnmkop9PIin6QVZkoInS7U/cgzLU9gbDjHx/AOkYb9UEBv3BzVGUVsQCh3V1j
ww+sXDDiP7tbFK6qLiAg7n+Q9t8lMB+wxAoj1tLMi1FPsZYpmwZHcZ7efmDKUsVO
wX3op9J4C6NVGzpWYFCcj1nwXBb+41LC4G0NOIEeq4B6+6uvFLcum1am2HDh8+Kf
uqNz06trZLQwu4cOml1TxaVdd9EuYDrJw2WKPCANokAOVg3t7ipkLiwv+la3y59+
NSi9GTN/EAxre6KwDRBuW6bdcZZ0+qrtx3FIwd6NhB2GHzKlZJVpzTKg1e+NRc+K
KjKhsrfmykAUdnSyHyHFTw7xRFEHYyeNHI/yosz4RfDqHHJN/Uosb8qQXxWT+wjL
zL4KXei+qg9SX/yky/WN4MAZbi7aNI9y9nbpYiXvHuHPDTEDsYPdjFSiu7PTNqsK
lhrDlfqZJGj4iX9v0d488P4VjbMb872TeA2IYSJcOc/LTXqjnLscojZ6RZ2Ec1h3
HPJgqRevqt+oNqN4JOYO6OfSACXjIK+QgYklgY5pwJPJNNi2fNtvy8LAtVGGoMjH
1bDwlxyDY2ufRf/xpdE+myCIlZBnAooiGEuqggWsUGx1dqlLNJ4pjvd9FoHrUe9z
gP5ze5LCAURz0pCxLs3Mbsrq9ei6AbPCUHHgNAiHWZegVn8rndf9s0/E9nsgZFvE
tyv8hn+YEDj71+3A0sRoSexsPQXbkO5bZ/V/G1cnLVPgy8+j9Oh7iGgVQpdZx7S5
Wu5k8m0Y6IiHikEmx/7J3s5tKdO7SZz+Vw1m0ORmdQCRm1AV4GnxdCqzOMg7zei5
fz1lYIIl+K0C5fUl4STGhIToezehnRY4GBWtWAjExaaB5M2cpURQMBw3VyYmH+Sk
Dkx66hnyHXsteaBo07dyLjoA2K8Ts6DeNc/hpdFaHCjNRUkK5GcEsRHTVYkhhQVq
bX6LxCXIVNDoatyShaXjrZPVBxqgRYIaVfY/BGQt+TnYcB7j0ajJCSllR7e/Rm4T
ZVfP2eTbtDacj7Gyp69R4znAPdT+eBs7XysfJUVXJOq6edg/IXMTh+oRf5D5dhIG
d2e9dsyBL/Un40N1Yp/oYsJWrNFfAy7gfAhlZcPUboLk5f6EuTLIVODLaejBKLfq
8/PI+tHhcDaeJKJrkX0gDhY/ZYuOJ9R7uZ8JIaXx/sOsnn8INWFEjBQ41drhlNwJ
+p75iEDltJwNFaeD1MUMJr8grmLJboynqBH2Su79KglqGyKFCmp3NatMD1Unp3k2
/Jv9PB+ETw/dMmwBBSVxpr76IomCBKK/9jH9xh0Hfqphg/fW/d0OIZl9MqAHDBvf
L7XBQs1PcilwlzCmRjPZRPbS6gfCwo5rJGbdJYOQvkwLMzStxsLAGlcNPQEKItbI
v64NJPXoKLv0fFvDW5t8gGzBHTX8fH3oyhLpjKx8tIxDRbUQHIvUEHq8+hldNaJl
/QO13Z3tgN5cgNBwBybXw0+sH1hiY+l3jooKeasP1AbjO0tDnjJea5qKayoMpg7W
zatI6UFxd2CfvKuh54x5ppFIS/jcko57hB2kRqVr3TK6InVNzhLVi2VYbRSRkGZg
y8sujP5f2Aqiz6aMoHYe1U0gEaJFBV60oIQ1y4KNJKmXoGWmnVApiWgtrC75lr8/
gbZh97OXSuHuIdDj7l4xX44lMz9mf8iUB6KvMmGc23wkB7psKwz5Z30xk+Rnnnve
RS8f9z4k4ECtmZq+3OKPAU1WkAOTt5ntWhDNfMPvwV+Aa/o1dMUMgcSr0DDcUAXy
4oVEYLppPczQY5nn29V6XEDjraxu+F0xhWWDi1ZrcVOLBJydtCNw8AG75QASJOhx
BFaDYv/LPEsO6G5fj9mwM9Ffk4z58oPS/4Z1gReIW2fXdOdXkVj3PuKTy7x+rwZT
ptsaUSk0UIZVscg9N2J1mlc7MW5k5UH3FPs2ftO/OnYIs5qFr46SHaTXsBw/7IKo
ig62ZBql9UQKJCriYHzrSCI+6i0YiRyEjHvH8JATqgjM2hIZMxoivdbyN0V50N8i
BnO6XCG6oI5oH+o0YqE9fWQ9gz5KjccK+GotAz+hbFneOvu2ztpUJEXtwWjue4o+
ZVsieKUxSWRPacaHzgHfadqaAjAyhVEftC2C45EZu5P8EE2LpUXjWx9T8bnze1Uv
lbFca3LfCxPgzIMYaT0HSqfAKjDW4BFwfNDqttK6Sla8zuMZS+w8ECTvXsFjurP6
16uzP3T0sYD8sBL6UwbQXjhV9vrvJU5OQ8RJv67NhFz0m9fk9S61/7HaWxS9e3xC
PLEN5hWUubZqUJ2aiKVSVyejCVwhClOpyPVVpPORplg7gz3OtFV5nvXhnRzW8H+S
XJkAy0EErJ9R948+ZgvNu1Ol+uTISEuhkTJBIXcf057tZSFVs43PdpCxo0kSZ3a3
LAJEIcSMb5NYOr63vX9X9bbCFMxtp8cXNJwWpzPkNq253XJxdMpI0txnBLJsEkTh
DqrUdfPQYHsdcEt6C8SMZW6H7RxEEbLdMKe9r1NY4Mm9489AqBweOC/Hyv0l9Ggh
kfBSKXNuz1p2Z2Nw+7VjcbBs7n/smvbBRO6BQZpSgXCFQZdvNSfpOyNO8stUKHbT
ICN9NwfmnFRjRgJHJ3QNG3zdmT/TTZ6YpvMzkBVQhGjgMORVjGnbAen28pvUpFyH
fdI3lgdUMyKK41WgH8tBxJ0ffqQDEMZgom5vHfpMPySP5329ZvWnaaZtTycQo5PH
fO+dsx2IzdBu+PQLwsqxYu0yEgX/dtJUQx1I6WhYXb4P14yC29BQUc71MF/+d93M
7wIIKEZ7OSCxXs1rbnKyd6zmIa839Yb1q1ljnoJL2lH6ze1vFMdt9jjWFMvJyx5f
9Md/P11zDuaNdZxIu/PH3+eOSDFyipOl99PvUaPhOvd6A2KEbzF+OHSziZMuSP5M
MeeziyVATtLAbiz69VS6j7tnGxL097qzWwwXevtMv6O/gRxfow/jpIEcjoRTXETW
oHOXiPKf8GoE09RXK2xyPAFcE7J1q4eJp36i8k5jlTGjsW8AIuAVSrmAczGjQzL0
HZxtx+SvGglVxSMJSup5AvRupQ0EO+94apDpCxdiR9+gdAjEcelzkBjVpdpsU7D6
mTSp7qukDBB53IAHPxURszcKsZfYhZbQ2yNH6d/g2TtJ3tHeqwIWhb2gnlTX3JES
aYekTQUFOb/GuOUB4qkvjGQxd9jflg/VInF969S/miji0WViZfBJQCwY44XEpIOv
+S+rGshpeeEq43mImqin3qmPk63pN1or+V5PJ4dQUmelt/r0F4s6PALatqAHCfZJ
C2nYy8/p9jQx2SG1SFk8H4ULmdXW5+Y66d6956zLFpoBeEIRY/lkM73kiyTCyIOH
Qmxi8EEQ+66Bri9ru9FRJfLsusf5IC2fFe8ftrqHFdXb5AQjj9MqvyeiVgULLC8L
XidH86L09T1ar/uIfOSK7/FoGQ36iGfH7p8YV8WHetQM3LUl3o6h/MGnubDxeTzF
Y8k2zz3hMJC8ZudBJ+s4X9XK1k/TRftUHFi+Inp5opYUwEX5UPQ+PBpQ+ckK8iUC
zK8PYlWw10h07wHmpmvPEmUnFToQyFurIkOx71rCYz3NYxRsBSDFJmrBMlNFblNj
3XBkbQm4YziiSXohh+oboeXsy65vwI2zgYIKKhOvOZwHvmnRSML05X7UkQqLAuNa
YwmgzkqaKIJenqWZukEGMzDUGFq7XbcH1+ns+CUhC1CIibYgrgF+youSLJvkea4J
g8RPYuJZNwcfRQdaenjqG+YaLg479QerV4tMxSV4gjf61aXlGUiFjnQEh1An66aG
merIJr487rW4vhMgZuP5OyGRVljS8viv172ORaTNW2rtmyraY9INUDbZSDympYLW
GyRQYTB4C8vmyxcPPAFRAOjh41zwALrLgl1zCndC1XW6fkJGi89FZ2u/o0+F9sqw
/OzA1jCrwA8PefBAP2FhV9Um/fEZA2QLvaojuiR1FyNIF+nUZF8qs8qE5YTl7KSq
irwjEbPpOhGr3BGV8RfMqhdV2U5Ata7UX+D5DLhq7mTOgj8PrU1Gt8kLtkr5LNR4
obnNAYt3GERhCftc9Zb0c5SiaM9oGC2mymlkc7cQajRKSQFGlynqlovWhF9+OZyP
DUf/5+x/Tmjc4Nvu6j7uwzKvOOF64TXgFrnOS/TfYsGAZUHefl/SGi/5jXaxCVpD
qxBX6QGjr20D6++Y/wi2nJKbbFSIpxwDuoV/K88wxxiXXCD0srmcuqK+OKPHXUeZ
T6SSD6lmQhfewESQT1ji8Dic94tP5L9K+XMwYeXm27cocS5g5/zPE1Xbh33ACQ7x
AZnZN9UXgv9sdACI3trenOxgRu8yOkAY0kXBpJP5lPZ8+VO42Yk3qr4vw6+ttIoA
HIMA0j0G+3y5zgZmGfwmf2O0Kwem5L1sViN3hNwPfN0GbcH+bHOaWV2xws5nMiwa
tMgyfHR8yomef3uOI5FrKDJM7cyLQYmCjX4gQsEuA5M+6j+4n5UvFjXQAb0/BQ1E
JRVWt2S/8JZRbTZBSdb2n8/ECVzKml1QTQRivUYjyOdUomcCWFFED7IJ2Azr2b82
dGENYmc3wQZ4zAbhxzhwAyp/cOoDMj0LGDOhYt552ukpR4YxID2hxmxnjax0+2PD
Uv7W2VtkU1eX0pk6BMnoCa1UD7lJU2JsY5RQe0Dh2DdJJ6Q/WI5Gryh/6MT9pdYr
WZhYb3U1pIzO9KiOITFjkN3wFTWzXsseLWjatvqKE/BOwrU14D0eI1ydrnGxItBs
5PxOpC+eZs9ttbRWW4h9cNfkzb7UVUw6eS+bDtTJ/ipv4z+n8npW0btOmFqxKaTJ
o78MQUSZvPs1JKY7FwtlY0ze7VVhHDojRq40SCZifWAI9v4FlhUBQjcfJmIc1HSJ
Tdjuk8k7sm4+e7FoLRz0Lk0vw0pTv+I0QU2Ub4537vWUu9n5pEHjSFub+cJtDG9n
ekgmnCzaSYTflPc1nXbjJLRztlLj2mBcftUqyeF/zMal+eUkXr/ou2cHSvrPuxeO
d/dimk0lqpLwaxg73bt2VYgRvgPIPXpNOhUmPixCaumYrQarnU2XeYigy0RIBTXs
+xOKCsVA1wX71evcWYSTPHgJB4FSMf47eJ4TK/axXGEYfjwGiE1/tEsOT5/cPSEg
jv1FiiPOcNMB6tdKsompZ8Du5p8g6NoreZMLtOF+D0Rmt9WqvSqx98HuTcKDT0mH
8MzkjBq0+rx04dH6aQNRZmgTkev+BqlfD9MxOXpjeDNZjFJUGF6vMWiNc/+T4Fno
EKOXq51ZbHHq4cGsFKaB6dhkJi+Jx72LvWYaqQgsU8YXNQ20MdYuV6EtoxG3OcUq
YyZENBr/pFM715QgDULxQ2ETnmYEsXDJkxP0Sr8aaCLPpzU2bZF0sUqbDq8d701f
E36NUZyESCgHepJ1lbnW/QileKdQ1WOnltzsQm8T9SXZn1Tu9cyTE4GJgSBkQ70E
HxFFjZ6w4ggGvdCcgsk2xj66C4Bwvp5JobmL42tT6Neg0EV6Poh2pwwYet4HBGpx
qri9G/51EOg6hsIozioa5wlMwSeaa1VyTT0f3rGd34xllOM6idd9+jq/GvU0jRaV
thqbjT+Ll/Wz/z8ahvrewC85qUcQZziMGM3WRNoeyHSapK+g4ZxmiAAPt4q5tWcR
9Ba+66yVfBwq2wbCmvGwq227UYKu/nhqfA38ToZ7vvk3cnogJBVb+0UAf8aira8D
H9L6kydr+ez6da0De9I3WN+m/CMBGg1x2ZUQh+0jJEDI0P8+yVhHPp/dAjc1e0uj
Nk0oeiKVcDs01H2h6poUaI2O2Lo6njBLf3yScgUO0zCyDP+fpWLkLxf3mUHrsHvN
HtQzYIwysm8uCFSZqjRArIwCap4OgqI9jH/lFgpomRHQQHj0cnIFnEXW9CaxuR21
aQrEAo560m7J5W5zwICVeacH+zHTNitGUovfUwBVrov4wVGI+qdSH6RxoT3LUYlk
MMd8kFhqBaulrtjw2e+P9VVWBHkSw8qPs0jXT0ExgbPDiG6n+1Pa5ax0tUb8y/XC
BpSElopsJlD3557vgb6V9zZ0NLlkmD7bI/d0TckQLezrg37X5qYAGElHZT0EG6o/
SkyBkk9Yu3XRAaurbKvr2p0H/c0VBBUnzKZqaEj7nwucwqtEDomo1qe/9tvZD94K
pOB2MSrlS/yz3GID38haN0/aFyO5BKAMNuxnhtgVAzIGUC80SVB/LC1HBzgxNQh3
KU09Ar3QuIxUi4+ZYWrvWV03PGI1CIitlLH3oq1j19eB4RUHRt1S5F1xbNRXEjbj
cIAMrn4PzqVtJRXC+HGZ/bt1RiTxvMl9h45nyp874GmRe91MyFV8PzKJ3D9dQlxA
iIB/fbJ9lUMy3bQbexwuL0ra8EltIcS4O79abEaAHGBkIl/tn0I5aeNdibCRuyr3
w4yujhLtgyJFLWISvUDz9fY4FZHydtZbg4zudsKC1IlmPCXIUrEZ6id4XtNnL5OP
G1EcjPINkSHIUkOBss2d/FS6DVz+WU7YXbP1S7xDPB+yn8ATOByruzwa5iBOsMEr
eUXYgwMhjZ8marz9hCySxGPaDcAe7sLcvRsABa0TUeZKutKpnvc1Ao/hK8RfiLwU
4LOF/gLTuGAdD4GIZZ3Krr+bH6k+iB3VZDsPOoAQcBqonUjdaRXek88gSw0DQ7Pe
Qf1pEj1aanHkbv5tc7X1miQ83gOlQK3Fo+oHGrqDlEzG/C/3QUESrCY45AwWvrdz
A0Rxf00ZMk1QQ6ZEHBYK3D5hZdU03Uz7EeRG/McHLwwgy8o8/digES+z6oM/HZEf
Wc8aslVRckdU4wKNSvMo/efto7FCsQUp8ZEFgreQLAdkq4y7Cdo1G5AAnmbjctFj
FjEORhjKrjdjCX5UCSjI3nRCpqHSDTgWQ4qIdMNhWOapPmmz9b/O1+3yNomWY/mQ
15SMZugVhpnXwsiaftE+tJr9Z6b1dDKhWGVJNzTzNjCpn23gcwOvhzw9GuWkDSQn
5LStUp+mvwzuUUFLIUBTfotHP2NxA2diUuIH365gewL17vVBw05y+vZClWlctvXy
T0pnkOCkpS+OOcmZteYFSUlhB8GQGpdhiZjPC7mHZIgENcgGqiC5RIkAiYRLm8My
NCOAFX6lLH+S/gP3pk4yjvU0UGI/QNdSG7qimQlrunE+4k+d3A1MNDwsLKfcL2cH
0c99giPxb5bdsPqjt0x7TSyMMDOnsQ+NpjLMO33W1Vyy/SFEFhjhHDBSIz+tPBeh
4PqGJUWhscigBZXALx80/3hEkdE8PJY57XTVf/op5Q4RknPFSnyyUDpVqnHhB8ci
mdjOct9htFjgUEAQ1xf/r5DkShToJ80abPux5mN3tE4bcO9/f8N4vSFXTD5UP/Xv
eDkPi/W0aoC/9xJN+7WWeRxyxBqhErER2yIA3iLNIxa4BRvg5rTDY6rh/8K2OaJw
xRBG5MGYpc+YRokc0YnHNfSkqfFS0lUxnLGJZBU1aZNtRzezO2wbAjR5ct0inqkH
MBktjJB2Fau2LWNn9lisyEBCfXTSAoYnko99gt4ZwUuDrTP7DdNjFfiGzaosTObz
friitbcEg11vH1H9w1SwBTMx10e8Rd8XAqO/prT7UUbxekUxkTSyda5Ho1Mq1ysC
a0E2A144m/p7w1ago8EaRbQakUcBXK6aNNbZJKV9b6AZBrR2bSB+EQC4LCPvuSDD
HSfSatdrWx85nZALfY4NtnrJSYHplwAi5RZF0rNRuq53oGstlEI1VTX8d4VjeJPe
dTA6pBH1ZSzY337OoM9vGkvVqiUaBhtEFhlPJIUS8fQgswBFMMfxbcNM5YdCuzNf
i3VUQCrEIdO2HSKm7t/0fCA6JUJ7XjT2eV3oTugHZA5+VDzplXAGQ8+ne1T2wQHT
X+Q2uzP//L9qhoO8dzIu4i0JumYNJYKzctVomTB2rZf2c4lzsV8feIwcTIMdmYk7
ehJGJlHVRufKCTH7uOY3z+V22vj/0Mo4vn4AymLfV1ldijfcJfnIqdrPoYVT4/Rj
4IqZuiAy+2lAjk8BSCK7kDcyKvVBI2/P3yJBz8Nh3KXQjnUwgxbgjrIji7u/Ww61
WBQ2NLhuZKBsHWxuiqsrf7vMgda04chP7H2EgHFMNAotui4j6tcp19P5ciNgGr3+
9NZnhgo9X0KEswRu883kUhdSQEpBrYCtqeqFR7+Fdb/UI0Arcc5TUxv70PaO9glx
UDAr29EEMoq+oLWxkTCzvug+XD8KjEy/FvmNFjjoTbXbc6tLiqoF3d+nLDS+nf3u
W4/8x9hWjb5kwE9fY1XASm+LWqzIpuLA+hNPeHOu/PMwOf9RkAFYbuKBmZH+Zy+5
NjJoX+8F90PdK5lmMmesuWNzCeuZ1wo3SemIs/hQDxyBYFLZMBFF1i30hShmBHbE
N/fdyErVy65iyz6OstUZVlWtyZkT0gIKpD3EPkusILcKBeHuFI6b4/dn/1NIwSfW
lYzlLBmki7h79j1n6HU3fW2owz38yFEJCqhXMrgs2d/oCJut0eL+1ZY/OMAZd0Fi
siMK+RG7PgWEnLeY3GJrp9jDZwgkfZYKcBWm1S2ZQxPNI+zM8RA+aKADGr73ODKx
BJhTVExNhCe/JrzW5AYgBSLzP+bExVEwjiLM9oLmXLUL2MIvlJczl//UcFO1pciq
ZrV2IlUhYnHorPgt5wDvu6idIct2CSUvzVo2UO8tF1EhE2rGHlTYnFwmdf4wqe+Q
cudosTkuFnv6i0pq+6gDPPrGUlzujgalt5DGydi6z7xW7AfpzTh/gupq4gm50qD/
jGXz9BOHf52Vf59UjAKZfXC4qsNEsBOXkEw1RW2aceBv+zUC4oyTM17i9mfsozqw
l8Xs1jtG50RlK7YZsbjq+zlbQFjqbIt3Gbi+gh3BK5AQaKVG8VWDnS53jVShiavQ
mHZhXfVsyn3c8Cwu/AyIlOhSlrefLoaWjfI+NHBimSKfKMgT8SqLB5AIF2gTad4a
Q5M5P5f5Nx6sOcvsWD0Z4lAjFpuSIE5n8Zp+m5I9CNjNhcSpyOohIwrZIS7XHmcl
6VrhysreWI1wlIXBqKH2TePl2SF2P9ms4Ue/EeIqLXeNewm12VZ/1ETKBw8jWyRC
PmjwPZCsHLzpYUax3pmdQRmI+fAnx9zH/l0XNcgJqtcXOgFpnCg3/0/NrIxNkw6x
Vfql3vg1IhiN94rHm8sHrg+xm4AAXBgnUYULjllwIs1FKupTGM9LF905TZBcLBh5
BUMDAYyABfVlxbhv69btOam+FDcX8JEsjZLExyUT0Fk7943/TO5RmBu1+/IUFllX
JQZPyWUw2RC1Njq6Y2XkGY8Hpd7kBA5y1PNkabpSmRXy/pMrHN7JwOBAaDS/mAr0
XtnSlvFNI9Pyee1wy7XhzhmN1rtTRqaUAkkgbhlnS8ivbf3+vP1DIuOvaVM++N2g
ZvIopZMF97vegp5oXKyjtlPK5WrfN4nEfs9a+erNK/CsiZli9KhW4c6nj5YCahYw
Ahg/xDiVQaVluTlen7LxvslDnbeiYXyl7nPcpvJVe2JtSxQqzd21RKdlLdjQYXpW
w56TQ8BZJdT64UYgx8HyilW5mXe0mVJ6AuKtGUy9NrnwkwbpnkEpuVn5Kt4BkFXu
aZIukgofSq126zELcFGHm+KChLqLO9UbAbWTAjc2JUachOhWOfedq/WiShO8n4Eh
zv3sWhDEe7/yzYv3DJdyHh8Hh/iAQKoSxqPaXtxcURyZdCM56NUHPlFK5UGiH872
3Js0C+PNtf0f75vwTESO1qrad1bYH4yV4WpTZo8slK69cgM12az9M3Z2J3ymLc1u
kn5In8pb7Pg0n/2Kz0uG9XTfwIn6opCsVpacHxPcrqj/XXvMcIKVpJgcCVpcI/cO
/830q8iwCb9aIxzlqBvJolD41V2X4sK0oMN/oV4nLrCAkA5c2c5BJHtek+mZygE1
ABIvAOTecZcWsOlJl0c4Dcso9ZeU4pTz350ESyZUetpoaoPWPAOuxy6UxKyqFAQN
Q/v0JOByLlxlQNhU0N8tsTerU+nWEGXxbC3IQSI3XgRorFSP+OiFWwr3trLamvrv
bJiBbPO5ym7GzfCYMPC3d/5H9nGBJOmEJ2kQJO9trsSdtALWetKUdrM9iHSI5Q3z
EWUWz5QVrrksIB5PTAb97EYGXlzThqfnlrZSqY3FLXvcCeNvdx33vqk+HmL+rdbU
YCiVKjMfwlZ640xkwyQW1HqS6HsLTxPTPk1+WA2i4FDkxXLux5aIvXhXY4bZnoZV
CjgcW4R8AWPWPNbpm/HAERArTuDzI6VhkK4iPUS7EDDyKw+syvl/uqxdjQ2rVC+q
8BUqd5x2YCxPT3JS5Tc7BdJdaIa7yPx5R/2aN+7liEVvzqFbn5HlN3eftcXoEq4o
fDbkAV/0s74m+sir+VSGhuYbqZf/9Zsn9najPFOjuPX1gU8O7O63dz5362BC5CZS
7g2K5gzqkKfb7PRoXjrTY454WMHuPOOVdBH0NXNP/cUZt0S/tOcCctTk6vzoCzXl
q1nxM/CWAtkavbtiwc3xnkcpJBDPKp5oHcH0az71qfiARovHPx66wfRxRO/U9T8C
weRKecyy/WLKKgEdfosYIZkWWJmEVvkcNuwrZQY90Ttw5zzFbuH5/O4Ti/WGJ4AK
kVehjwmxIgHwff6EJrpdoiMs3h+pm939zWbgJ+pPKJOqbs0O6tfSxYh1LUQIWdkR
8+S/8it9XP/1DxDeDpEX7IKO2zWdZ7uwaRnog5rPj8EX3cpW4saULd9r7PWajbrO
K+EXJulrRwZ3h6upOwaFMFcx8WiY1PTiCbGnLp6byHXQWDjRucyMgRmORz9nsyg1
uWs/rWx8F1aZoJINn6bWh/w7TftIz8vtbP7h2xY4u/vAKfnNhHOIa3g67w4hqo5j
sbe1wIujJGrR3SNjvnZglu8VOMc7dpt8MHJvi2b9IOELdAQ+irbgVAYU2W8PlzuN
Ys8j1BOBaiY0lXqc/s7+ZztjRyEDpSw+pit1N9Zso8yDIIaaQvFw9P+fDC+vBD0y
Fi5mIAlBRxJYQfYspM3L+rhmfga3Gl0s0pGw8I3Lw4LTldZXh7aCTHXqoGDKJz+C
xIQog4qZmaTipGy9NB4txUT90/3DryORLTrAF7n7tNRZeTT73zU4ALOmESdP4wKS
3FckXHT2LEkJEIEXfiX7o8TjgZyRahGt8d7MK31GUD2m25b3Bsw40r78kJtoR9Wp
mTFc4pmfIJBPqG+IMvw4pOMzYR82BhD8z87BZ8Z9dS6OG4fcbt1M98GG4yn7szWH
UwSFXpdIYntkTV7rMFn+CxKHWXXBhsHB1NwqRwCKPfgOIPEWYWP1tbtyDw9fKhFm
u+L3ojZZygeQfCGVW8dzAryMjZOPHVd8Aeg8tziZ9B5xjHveVhs6CveeW+2I1Hxd
qLU0dyi7chtcM+WcWm7fVndLATu962VXIQegwkr3M4RSyMAWRm7iKG3+rQgnGnD3
7QyTXrF2GF7vD/8OgvoNgkqnfaTf/jlrQiAwurBsMSyqhuMKz8nAu6YPNFaHu4zz
wBTkiEOBrsTLpmcfWlEQ4q3JL345oJ0i3D8IkvDCe5gWQ5XpdymKMwXuKVRBm5Ln
X8H1WurZi7kbdama8f2YfaLwoxGz2VLPtqnGhrKBZ9dAf/cDizYU6VOTGZCniZ2x
c722jVqrS+8IkUMrYQo0ZLw+8Ok5gTH+PSRvHHKZIHyyCXSTRjgLezy3ctDe+Z6v
4vtBrz0vij5B6moXmlxwD7PfWMd3sNAe3YRTz2plFgFnRZpLJlEnkXJOmPu3Wq+j
1XAj0DriRWkAh2rZ5I6qxrS+eoffHyhinB1z7DkVfuIe5bnnzTA4gtiqnRlSNBKO
JbmdNyUTvEwcYrOhDvKCBOo8x+5mubt5eTw0lI99hqwtSFsKBSWdD8dt3lukolN9
uJchhjvXiuMnrRw9b1tFh7yz2yBctr8qbdYP7L8K4pidlvIO7Hozv2BZOr2vn2Gs
aSenAGrIs2jfpRR9tHFSBOZ3wJvAInQqQfKL821Fect5z4brMLqHOfGa7y7vq8BR
1j8oTpH9pU73j6duQg998+ny9qByWYW4Kkl2fu0wfHrgRPXZ0WxI5/lI2yPWoIxG
STswg5Spwz8cgK36ODXZfG2iOa6KMl51ECnk426u3ztHjmyqa6JLkoM23KfyTTgo
OuTJqbhkSVDcrIK4z8Ucy1vXOlZTj31NYYD05Z58GPR3BN2khbWtBUxtEPpyMjzn
4ic3ag1F18qGqVcO/FplVV5Fg51fxWLmvdzpr5eZDdadS+h/D3OvDQmyWu59VNQx
QUWwXvynPQNlTGiBkAFmE3V3oviCwgQg2IrWTom9S3er2b/YNdAeJgPGjgAHwJtT
RqDUyOfDfl1ytNOSDiDxtGS01seM36Tx1St5oMqqVlqXHSVc7CN+HqJDacGvi2LB
Gzh27CRlB37zchZIoDO5EP7Ikr/123uE7Rt0MRl7X32kn57DIUK85p8ywP+BT75Z
Ho5tT5UVsGdlkEIW6qRaSGVijoaNwaV+m9j/oYiI57IPgjVgBhEd2E2P2Vdfequi
nk8FAuqFWgjlXeMiJBTYC8QK6BAA4c93cv3HnxNNyfbc4HQGkOeNRGh1p39rHGio
3Ee4twd1wknb4+MGQzYQHHZiuKYK2dMFZJwGYbbaS0XOlbD2lRLrzjNU19C95IZf
FsRBaRbyKfpxT8z3tRIAHOS6VyeAreBn6c/utQJTD5orx/35U0eIDPkNoPWnXsee
9NhzyAuEqI4aCtxnJIj/L/kQ1V9NM0dlSBIaAXUFYVuwWU2yhhKk6UYCvIPfFRNX
BmiI91fC1udQ8UScgWUqVWFejzaVBYCB5uwQIMOsQIm5FJR63xNMAW7lg1HAkd8x
l+vkq1uRXnahFPxXjsA9JixfMI1QBoo8WH9MtxvUGzHeqtdNsqb6LSzKaNCFO+Ev
lPvLZ+I6mzogzPmLeM0yax3cw6Gkfj1INS/9lA56O0Pd3qyYUo1JGjMpyLRSDtAZ
eV1PCNqspC9d8rUvLBjfT9cgrX7udz1a3OAECegmTjKPDBIlFrVdrTZUvZIIJtMt
oRfJSAUxIovRuuHXF8+QHHFPmD41krAXfF/24b4WEf54xN4/zI/sx5DQbwEE2V2M
Z9X8n/hXTZYrKqDxbpTW3NBp26rvz9h5Dd5/gQ60eInBVzWnhdJtHR90ynD7EEeU
P004y8C4cGTcqPiFC5UXWE3iVqg12bYmenR9ijNKtsbE8YMrgkqD6E3vO7tR/0D9
qVubKnoFmSFQUBPLFtR7jQ4OHTIZ91fkk4IN6nRaGNbxcWyFo8GImr1SOqIvZDJp
temlDAsGPujp9d/JaTA5vB1Cosxo7qFtkNEfX8gtp77j5bdg8hoGEO3JS8EKBnQV
ndt7+DHTg+/k/8SEUL7JduNozvQP6ciYTYab0OGv4UsCuZ9Uc/QpyxkqUO61a6b5
CpV1xqffG1qUPObRsTc3iQ3A+mMvhQ4HkkPyr9YayNh+QtKYZjM2VsQAqE4oR7s1
Finpw0OywesyjnhefZuQBxd2XJ+Yq/A1BeIKdp4UOielRQkRC15g6OvysUcCeGTL
jNpmN1cDIBT0W5YPn4/Wu1J8eAFIoKvdS4cKZwmtkNR/ALNKUVLHHiz/g2dTPMgs
kUuCyWgviyRjbTULIOZja+oF+Cv+jNSQrKGm+2pE/LsWEgiNo2z1bo/vefmmLiQD
f39XDWVJWWHz/uCG+LL/wEdzJLZp/EwESfaFH4g6yyfL9AxmVvFn97PiZNr6sqQ8
2jKG0J2O0k+KWcaKrhj6A5DWRYuOdXoPf6l8adTru0ln4f8uM9FkEsd9QLWt+eYR
h3yAsDE4r1f2FMx9YcZF6PyMXYYEK+6TwzkqS+M/CRkZftti9AXoNQeWUc783QnO
+ZjNNYtVb7BebRnHrGFh8vtlprIu2z4PSm1+l5C8+W7iQaAawr4wIHH7c9wYeFeh
R2D1zMFdXSJL2lOVzTHykUIDHHh4YbOs6dg5tuqSrhJCbd7tBxVSS/dHDP1bK38s
a45ZlmwPPmrZde2gAOEzIKzITEdUusi8UV1+IfYawJ3vJiLHHA/bz5uU2ENYvUSA
0KEvdBTN8L41ic/TLIlfsgq4clOLHO297bMDOWut6B7y42HS75KMx4TYE9AluYw6
AUA4T2ON4MG5ddGIsbwamatsj+exh2GMyyaUH8loSPoc7DHlFFZIz/G/27XxFQ1a
WnY/nbLAoO0c5udst7LmzoF1f2iSUc3nwdfMiIi3GrqV7IzajSXP7YYW8IIw7zfL
OvQTHmVJokSvdWkCCWmYXXFxPmjyMCb21H9xPTAEkGbJf7wisd2L2IDueMxe5RAz
pG6eGQpc0DfWBJrM6dOMLeFAT12SILqNbVJv6xB3f9uiTXxr41cBuWpsXmoIVdUT
g9Mek8Ie1avKllka5L6Kqd/trLeJBgo2gfoBgkRw4ZImTDgeLpl0sAZoswhitLF5
BzGqrZi/yQHl0ZJu3E7xdvF6oQ3sTH+3L9B6k5QIGjm0Xbvyg0m8YhAOMKfLKDK+
t9Xoe4BGXVR51x8M5SB1SAwb7RoE2v5xM5Xd6JWeK6vB2sfdSMXNX2ebOCsQdeSE
hmPPbfbGpkIMuMXzRTxbiHLA13qsW7i+sidsu7s+fVc7B0tG3SgqGxFGNVbs4ufN
GhsAdZa293eFmXmpgOMnAYsoVMlX/7Xyioea9uPO5GOYXzrgZQ7kWpxn9RC9v98q
LQYTrRdmOROZ6TctgkZIofaHflvbLagDqbriOjCMcXQoD3CXVkNjUjPNtreGI8PV
bMOSyw0/AunKfi8hui+d/a4gIrB3jk1h5lylKl1e5opiRRfgssMNBpRcykWH76Lp
oQRgUP0SYAO39s2AFKJFakM4DsXEh6O9Txk/9grs5wutD3BMg0NMH7HgpaJRdvP9
GhWpERdVWZ9ZRAjhJwJLGfNz2v9da01IvKkuCp+e0ISyXTmIV1uKZae2AuYMQfII
I3AI5AjknSYWKBEFE64SQ3Q+wAqt3HN3PUgIWmD5qYZeFlCdEaih41jnKX5MbA1k
NJYK9kwXTULDnBAV41Pr+KueutXa2YXwFEWACxMOvNWX0oQ8VPBYRedcv9pPWap5
b8yNc3sjrtctYngFIGQgEN/LhcopnnN5qBXi1WjMM7KsC8WvV2QwsX69Rck6U9m8
FG1hW3IrkthNceoF7Ybcon+Xz/1aJ5xtMo2XXEqtl+7Glu5b5iHd1BdQg1SmI7S0
E7C3207KGaoXCl1yP/u60VWD6SyKjhruYRe7wtr+PovTt7Gu673GjsaHLN86K9XN
dYluGH383pBY+Ouyske/fGiajtotkHLGSSc9loDjOofYSp6P6GBrEBrrdWMSDOyB
DjkXWV3Xirm/S0uaS8jYanRq4dAmX49WMvHilV/T8UkEZT1tSEsL+x1oJFusKcKa
hn4UBIKxiLkdt+Ush0bMN5Lfw51GLj67sdpfZNTcHzG8C8/AWoJ/tmVJulymcadk
qmaaJORuvkaMlB2vbBl332SK8YswIP8rj9aCcPegBp9kx8ntzWPMXU5VW4lh62bO
agPxTYEiyVY7HsW2IvrySU9g3ULTc5sXfkOmXBHCYYhjTR8pI62w4CACcOAOQdol
W19AGDlsZc9KgDWDBI0JIXm0ibaYpRceBcyqi0m75AASHWSfxCS3Xiv+0buoXbgL
YYRjn6Knngc/MxCkLo5PUXJHbkmDhyrrPmkXoMk3TeaMk3i1Fu7eaJVJtXvNnpcl
8DjqewISds2H7Q10BTBIXQZ9zLbwRg9v6JC+jbNe87aEpS8rxFV4sxVqIcCTO480
iriyAheoKVZYiFUWPHvkQsEFVhTLISlifpmPTA1qygvKlKbTjYHfkMalL67h7Oxj
fm462z7RmLtXjzqLlS9NNKDvcyAsPXZy2fuk1aWJJe56H7Xof1rgdJRQlYTL1rJc
HbNLDJdoLvOqYQCIC5tmbnK19ZOjKhZFhgaZp06lbuJqpfpKSVbuWd7ELAC0XOjp
nBoqYpe9nLkUHH9cqgaTIZf3AKSrP4+xKqTAQzMQwU3vOpFkOrjDj9p1wkroyJZY
iUQIEqfiU7vgXM8A4olvIOxhpufOhYu4A72jFXklJCCoK/ghn+yI3IpoF3cOzZ5P
nmWx/5RID/A5EcH5CT1A+Vkkp1AmW6nh4E+LksnDXiW/xO0Gm22absCQGoHYDxw/
xpXw+jYXu1cPzQHWlxpQhS/Xvx6djir55/erC30+cOb+0YK4rHkjedbxP3b3yJLa
2+ozxgK6QgHm7j+tNE1ssbXtwxmK4LgRnUPDiStLg31sKgw+MeS8OQzdpHCSn6nh
sPbgLKCRjNKGaXlYKCx15zIxIDWpp+BwCaUi+5B91/SvMF/5b1ZTm+b5FtgFFTgf
Wm/+425Nx4cSscF/OKIgc0gqNo5AJjnSSMMrkO2uh1AYjgzlqHEeB1xi9joRW64v
wonGj0qEK7S7YcFgeA7TqgIijK06jM8f5waAZbJGdEkXoNq+X+ZwNYJIYrshrBmF
m3k/ddHnvcMhWYgSkAMP5x8PFnl5O6s9FbpmZaNV2aJmRdeo9a/pq2ZIzIM/s3Y8
itvw1YOlDHMo8SiIiO5hOkmiNmRk6/iXvhslNKtkcZu01Xb2QIMEPOFJddODRUvE
VbWYlZixPON6GhwVX4TkXtUL9ICHqDVQxseLk7r/5hp0XXr67P16TC8dd0yqTx9c
NFP65XRkySR5xn9+NaaQjYmbAuhC6T0rJCPIF2Lk8geIG7ev8eFzmU5NnEIx0kWO
vwBEIxf2LN+uP66DFfQYC/AQ//kxQxjItfM/i8DP9b+1kLn3y+5EryGRKExyLxxm
uR9GK9tEAWE9mYrjJGtra0mSEUucwtm1MFkTaPqSfmffJrzK23iJg/QienneTObD
LRDBPwIP4PvkTxALSe12U8OXL1F3sMeoyuOceF1nnHOxqA6sbEmO60u2JOr13A+f
JGkc3sWXr/lZwEBcrz+nWuRSmZWA1NT4jt06ooY2Su3jGGgRbVBa4EIrb4zoaFJA
EA+25OeSQaT8HOVc5ciPR1imw9FXfX8MpXCndPMnhUBdgdI6vjh3aGxRw5aeXF1f
5LG6jK/kh79gc7y6vgCb3aDuNUAVeha3e36ELmbDpJME4IcHK59piXcrtmPTm3ar
N6BG1NdhFHINslUek9ZxQOeP6ZINQGiNmyh7INBv6u5MohLySmIpLsaq1Lv0kYC9
wIoeWhXODyToPMYkoylQQ2n9XpodpotJqF0oVOPdpqK51aXdJoubWU12rpN78Ype
l8HJUuY4OtlNokQ6cJbWW6kR1v4oss5/ROFegkzLmJ/JCju1D5wFMVLaeAc5cDiI
6ZQsiBKOjYEv9hrlPYeIWaYx2IgDC3VGV3rjhlaITNPjHwlUk5QZjMlJ9CAZ9dNY
CR+OkZVsQjj25KSyi1YAYOoEN9DgUmsw14SqCqgxzPiP4zN3xwqVS7pWBMgCI1Fd
5YxIgayEg/zRrCAnxd29azjYp6wFO+0AJvdCwmDH4U0AzKLtDVKd9sfo1ccRDAyO
qX7ldp+VQRYK/NXDaa6fN6cuOiv1qg9cj8MPNt6sWvKOLNtUYscacjtSfVD9hfta
cToYcN1cU0I0oSdRO7jyS0JZ3Z6btt2x/EV/swcEUKbJ58OHn/C5ELUzI2lwminP
ZotWxPwZAMYDqnHzRm9Ilvgdxmf4Oejpc3q+fk060UWMKeP2Xm+otBwbiDlF3K0/
t4wY9tMWzZfyJvZk0kcpc2PybBUzQTYQe9QWiXJ7KFiBtvaKKYuG1Lve5yaxYrcE
3UdIvAx2A/lW9MgRC0CxAdYY0mDIq8V9E0ma93YfRcg6QbrnuT1BCzLCplu/EyWj
/JazkRQQhzt4rAhYGQnBwRj0uQEuccE7Ip2YtpNiCvRR3RvsBfpnE/WmWZpOy/uV
o/9Bz8nN1zQ/Qb0I37JE6tmuLPpaFkXek8gIcCDD/1D3Npun2+6IkibPKVM0LUhI
rT0xdkBtP9Cxc/JOiu90B2vm0fD11uaLBKLLW4lV5D9HtciFdnd0yV4JxbpVcDUG
T79YyWyhr/hZ6CdVkjLSweJHkcpBcNdXyIto0op4pHuiA89dMPuMFN5qga3FURbR
o2dvKLrfCNo594/6qANM42Av32yET5YQP2Qsk+oFMMX2gnsQgwz2Uy7zsgRXSlD3
p4gt5qF2azzvqOUWLFjXoPw7WAHgBFL7PI5gBOPVD90jhWvpvuwn7AH1IzNjFC0w
ezwwC9F68BVaD/Y3sOfmOU7Y7Si12oGwYUTwdtlWbZoEscff/83e8qbc1Ygf06bT
6cddc0AviSvZM53USN37HXkqkoAWdMzN/KeddfFm8kXvfBwsmE+3XEYhQv8ZtQM5
IPDnYWOxwmgzFa+eXmR0pdAefXqgC/iLXf+DBwQAeJQaB/PCLg4XY2LXp/CYQ/lC
XO6x9Gt1eeJBthjsDiBjq4ODexo1k/mbXCy8oyxm0urwktTLb2sTxYLa+dY6mXZE
4NFS6z/PR9grpGzDhPNwc6ZEy+bV+JSnz0HCdEH0X/G2MWEM5iYoVyTnMv2xJ2qa
PZPtvQAgg5NTZtisDJ1x4aeR2F/Wf/vtEek52fadfjFZnxyQ7qxMI84FgFXuoAFK
1PxSpzfjLXWNXnFVvfsNfpWrsT+LlCRuDXC80Fk0ZFiMVKN21m67I9X3KBNxIWPE
FPeXz9dyPpAyH4m3KrE2zywFlq7wCrvQAnnAKp8lNniBlSz7MbQr5bP+J9h6VBNP
b1F5kRWgo2B16+daPXkCP2OISisf2GePBRoeu1zm79nDMxket9o4vtCMTkg29y0z
2BwEF/n9IyYwtcMJupc9kfDWtWwHwrCCWhbLNi7diw0J2RIOo7gzMR2x9ceK3HlR
5hYkG4m1qZi6P0Ufbxae9iLIEvwP/wvNC9N3JOGfP4XmrDbeZxsZ0T84NBUI/Vwb
/Ma4Myx+mzhZJSTA4PdYmC3kc67nEUmOnRz9pRz1Au7PV8nQUdM//Z857EGdFyd+
LhJdW+FrWsfpKG2VHLcdAYAoD/pq855T9CncAtDywxGDly1/rctnxNWm+oxxRJIH
j/X2sj4empPMmnP70I9L3tTLS7t6waLaYUziejGGskEG+/lX71ZtyHnzaD1BArHt
VEgHAFkpx2iahuNhfM6UUQUNz/+KJKTTwS1udzEcGcuNo9CiPj7AbXynJir4dCZS
fjirhuVFPmYnAh5AOk+PxAzLFrouL9aizjd32JjICNPGuBPjfAlqW8euqayC+rCh
BOdQbl/d9escN59j/XaKl6FA4NkD4VHNwHPXgO9TSnxTfkLPdGMJ09TConm+ha8n
zdzhCN2oOE8IXSZbRPfBwQzIYS95M9wOdUfuht7OkdAYL1hEXZrVLtAkp2hhZ9hF
xs93P5V1amPUEQdX7m36CVXOMnaiXz+rdptcXfTUDyI1+MXL+Tem9+u1ZQ7CekP2
fH/J39+V2BNTmbRMnDHRfNyWguFJ0TW/bJbO15DAnfKD7YAc2Ct7JhV4J92eLJW2
mwNUCqcs48EQxGGlLbTl8YarCcHaCegRCPTs1YHrBctYzxFhHccndPt4ROy+wAYH
KLgXxBzMMIX/eg+fmo7Wb5/wwU8QGwtJzMPg9g00Y2zKk7nUAK9a6rYaBisTeAz2
4pKsbqMv2CeVtNz9n/NP52/HmydiwKbJZCiLKgQjwZzmLLC/kUw0Bdj10+XhBGV2
rlu7CU1J9C/vDU31p+kHttRMxNLArVifPPBp0kh+aagrKrFIAci4NeNa6C0zzTsp
hwExPjzMbB56dOvzHGYOoxG4rMPl/HEsxx/Mz8Ib/Ya0quAi2fVPzAXmU0ZOsFhJ
P5vM+6E2uHnkFxA6QfbtQmrThgWhTrsSVz2MiUxLTPuMc6o2uYEKwSxBdGgYtZkC
8fEsa0KBAQCChpidKE4KcV0o2qoDNok24ZVbMNQUnFoAz3wYU6eHDHyLoUjBqZjy
2WVnnHiNgx8cBeiYF6I9K5oWwuiCiQaxCNU/rTVhvynUP1dGjbGjshlfRc2yZagl
A7dcDFEBHWj8R+ToFa/5uHUZ7A9GngQvWAepjUGAuJtHXaTZWfMt/MFnnfRPtFrS
vbWZr+aIZYNeU5q2t6Zt+I/K1T1KZJoWmFHNYA374W7y6Bgyh8au/PKRkswzP337
YYTKZU8+slkzYtMtJD60fFJyhm3nI3FJwklrbfsKgCoydYGnOA5g8zUP1RxKG72H
QkwdMMdKkDay+MdAwtoYj+oodI9wd0GFIa0QSB9R+7IIxp2wud7c3GfFKxPzShQz
UuG4RBgvTWzA0LC5uWil7mCxWbihLUNtjL4kT+kmYwLlEsYpF34OlvSdSeqnOVSk
8sPhJENYP/2x6yEl5ifrKpMj0yhHmYz7v3rtRIfOAjOOjQxAhbYPLxJPtqLtwAH0
aCozfDBnh7oKw0GsEfFZ9vSlvdBat90bVFZEAH0aP7+WLDmg5fMMCVaV4YnOq6If
4mn8s02ceMzn8BowQ1hpsSQ7ujI/GgIotQiapcaUAOOsUhPaWtkfXeriD65CGL1u
NKBS/AnakqgYV+a2neBvLiybsvOt8v8qrV4kQZKxaUsDAxW4+15OI2zsdeMPidkw
GDK5xIljA2zNnRDgKwV/KM1vWfHB97gvEDBkDuPQ0/yqqJJ2huWr3KrIH6w8vEJC
cw5ZNTTSZVPwzCWZM16kDFytz4fMKkI+hQ41DQxShak/muqF7EWGfNXgbcELL6bj
RyR4JiplQQzUj7IKGz1zVlE+LrvLP0CHvdp7Sz6/O6N+6L6iD4qkSV5Gfip0ceVK
sxnllTMCLNsntbvUOx/1MUvsztVhwJV29eTTcOX6oFlrX209V40ZZKDkRPy/iR9A
YXOuRfDyJln/yK89xL/NEF3Z5gRd97Y6FD55WUND4rC+2XMFBSWR+rCPRpvL1SUT
e+yp5oGTUHoOUmlHPN28rfn/qa7FK48+zMNDYjpkb5NttDr2cD6tzINd1SDRfDZ9
uUae7pdzmlX9iXwUEsWmpWGvev8zxCsgx90aLdteZPCO27JT6MPFKIRrJ1mnAiPc
IfOd1FbqKfMqUUo8jPIyJ7imH/n+9d8EvH34LNz7p9ytswPdVSciKQoMvqKUOcGW
YLtAqY2DvjgVkuQopjaE6sAU6wSy3yDBmYDv8F1MF5JT3A+icZHZj2lTVCkVou4x
xGOdAUqun2W/1zioanKKLvUzkLSNZpJZs0ComUCS+mdBLf5CK7aaASK9C4RQ28uy
6Jm1WlxW2V92ProHLGmwM+4XNv90ZOZjpbPbbhcsaQrXP9icYi4hPOrDLAP8iXPa
iUispDBhLomzjVnBQ60xvDRz0zuCyX6qYmjUZr5GKCOLL7KfYWpDEuUobOvw29Xz
70tBXn2EPrsColNx8HvhAU2k6/BubuUxkr4VZLTtCJa3Q13pxRivej7Lf8EOg3RE
4foMSmWe8gqN9hRHotfhczOJXsQrw1h0gB0jxrJ8o/3/fOmD+RoMv3NRvzuoacwO
Dj0vTg+fakSkyQQqXCDFCOD5G6jTWQ4m/kr/LD5LmnVsEQF2nbcPQCz6cGA06fIo
DQKVs+T0BIyZzt4rYCZGfovVkgqom/GXg6fLBRDGEptLHhcvxLrkvzKLdBp9wMV6
abn6rJp1aSWOfQBusokAeVslogYLEswXCIrvaZr0jGecw6TmTQFa3KRKjLlshyuB
BwQZnt5C3CfJV1vIPyy6JmPAkh50qEn2UCdBD2HvCq+yNo6m4UWNSDXHWWFLxDYZ
8HiFufRPmWy9X7+czKP4CyIm0iGE+CulY6y6O4M8dGh078WArd6CKi8WF+DHdm+c
jRXSS3uAwn+tI/oCNF73Rb4KLZoTEThjvGGwx8XjXpZ/VNEQzQHQFhDOJlVdq8wx
Vi1jxhH6ulcTjRbEKWXaHv1U2N42ainWFb7nBat1RGkQ2RXAYAv9FH5/Byk/27+9
pQAxDGlKW/H4p4vRdpHU4257xMeJmOowc/hyJhla0QknF00ZHQGuRDcoouHiCuFK
NZizHsTnTYyaSwG92h7R1bAirTHW3QTjTGty7geElSwUURnjHQEMek6fhp0X6gKv
Mw0f6PM+BSF70wpH6g4WrLnbABgxdtF50w51sewU1uSauXz2LCMQ2wV8CrizR4je
N2gTH2GL30pOWYkwr0coXIvacasvO6KaYPVDQj2V+u5ZQeaO6oGtD5ZO6KvXZjqq
joD5vyqNNEE+xq+yRC3rWoiD5lrz+Lo71QzT0SlaegohuYWrWYXLwY3xzcEYLJbj
+G2tvXj8wyorseOlCSjZ9G/cBm9MdMy034nH1EFrQyk+7fCE71qSfUs2GVuM2jDc
1PcuD+MF/0uIvIvwv3bCLBLiKNmZVgEdCVviI9Fg3SQh5V5sfH2pjLOlePP0eF4u
zut/SWJnwXu59rQebSq3VzeMBHptnxcHEv2MMukMgyTNRRWIGJ/4+/J7pxk/r8LH
NqUn/My05UvMM3/CRUaKZtzRn/z/SAN6Kns4cnb2zDCrUAQfPW+pTCQ6RWHqDSto
j9BZ+Y6lE3+LQvGnub54AgvovSq6dKK2/9F8kNtnjZOW+yN4SSOyMOS3kINmehTT
kV5gGbdjdocJCtz7SYjhGAj25Escq+OCTXseK6WpokfK3KCAg72vlOzyzv4r5O1A
EXvibIy4ZLgwPgvFGTRTc20hG5NW+0Yfkz8R+rb1L2Krx+lvIp+FHeHn3Rt85a1L
ofHaUBDSpup2Dp/5x6p8wSPzNVTOH24+M3mG1of8OAuOaydKmWXBEpUPRLWFpWnT
2gf33xgbxEb4LW9yxcxgOsq04cU+o7GrloE2Ng3jsEVOA1lwoPQSasFMLNKzFpCO
FGXBXS2eDi5nroE2wcfzHy7J90ZzJ8LCZrZrfe93JCj/T499KC4JZMUBZ/l8Lh5/
BJECJfUt89uBXKdwdh9SRZGnl21t2fqf+ZYjcWY6fJrWldIOqw63c8JM7ZzZNlBX
tXCVGbb7JuM4vTLKHc/QXE76TdhyX44zbo86Be9O+DYmydDBbaJnQcGXFsGeYrwa
ZG0WN+qKQvZTA/+WWLr81XL+Xyy73ZbVZN0C26vkG3tcefgkgrP8x0WwyicUrhlE
4JNybbTNyzbtzHqxZDFD1pbeS6zcpobUB1fiH/anivREaqmRJStPIZ4OzJtB4pql
V99FnWlSmsFfVpLyagM1lSAle8nRwk90e7Hc/WabUniWWZrUrehV4mcl5gZF3J7s
u/1GK3QKvdpXEGulnacwszeepJ7KNW8CzzA3z0KTpzwGKdD/Ck6fItveWRvmxQPO
yWB05je89AwLgPPnZy7uqMcNIxmC8Ud9IY6C5Njw7vvOraBNkK9zn6BmcZ9muO5G
wp46bbuBvq6XCVn/hr5yDYp+gd0iNRbghNxQDU/PQLfL5sczwmsMg7GLyMXtmRpE
U13ctt5hnYVFy3g9sl/4euFcmEzkqTXfQwfsKFIEyjTonn44nGW8WZ1hCwgTDtq+
DVXitJuCdcLiJpZ2H5LJEuC+hvWOqLT5yfqQR/EOovo+hJ9EeUsDbQTX4MufT0dN
TZnVCD3rxXILIGEj1mnlETuO9C+7rRWPb3P0PrCyEeF/Sz8OLrvJMfWW/Ezg4A4H
5TG+I9r5bBn2kVZ4stGz9BjZhxYjxslnfFrK+7op2LFXLHTASWlg296SdgqWU9dL
hJufOtclx49bVtAcD6ohfSiSGwC96piI+bqWhUxhrXeZJQ24ZEb/Wwdu3ZGUiZ5q
o5MpTZ/f5J3b7eJE5L0NvKuMS/vAUaPwhzQM88eSfRt+3u7x3vYh2dxI/2J2Ulu4
UmgxA8jBLCzWVbqY6b+AEc20jHSY/hnaFNuxhwn47Ai4/M0vttjPriRRVlicp4I3
mlsVskvg092nL48okPf48oODdXg+pDs/dgE9PUZV22ANMJlEiVU477rwMd10W7X3
B94MAVpVXxBbHn9BI8p/IqnYiszUFPvzJBW8D6Yzkfsi48P4vW8q7CMIT9y/1kKS
Kp94sU/56WDk9JV75b+FEpkokmYjEDOsueiZjutcvXCBEixzn4ifU3xVAzm8F7Zh
TgoiDoBRcQZWwZUsaFB3fO8P2NZwz0ysMwd9vlspWBqYTrtZ1DyE6xRU1W8BSw3l
djPlDv0Fdk+sX2QOcRwS+blOG91yGNqfzU6Z1BVuPF9+jN4o+pD2Rlc+TN3gd5A8
d5EPUES4ClRE6Y3h38TN2OWKNpKUxn0I/Do/PRH4+F8SBN8o4Ty5NgjmEdw6y14Q
nRxmZ06mk/FMADx5limICAq/ICLbG9Ua/j4JguKJ0M9eUD6tbdHSQW9EkBFoFnd3
MLvRFYPos8MZm0nntb/yamB27aars7B15LcwZuZS2qZD29keV0WQ0zgKgLjWA4jL
UZ2KK6X5k6GLYXrzyb74nXAmbZOhuYVwXZuQwPO/PUGDdgNhk/x2lG7X7i/fS0vq
MS5U5BASgqvl8abaG2HJKaVHkQXf53LfWw36rtOWzLg8i9BIr3GIZc60ajCwC6Dd
fZbEfP5gu7ZB7lb2JUg1RFnOl49qSRBkGkOx3ewo2QibRR2lWFNqc2yIjq/L4TLb
YHsADM/GTEVgRksmP7JNLPvoRCCRd47s4Knc84mGBtGgIyIyWh7xWclYEK/WOSVC
wkyEJJvoOxI1lT672NCVg5nAxCF4BMyW7o7KvMYTqRyu6e0LjTIJiP5Q+BrxzB/2
u4rblsAuv6pzKh0xBzTF/Pa4QzAQ2rIZoYmulZ1YuDlPXvkRtvxYotePWkTzsXp6
T8r/2im4ofNo66TXbjdAkaZCXigNhNMjdueH0o/PxUzCV7LFLA5GDUi78jW1mWgU
ocnsLXy8YWSy0S1vrk/0me6rLOGZ/tmn1BpgZxG6Y6Fig5gGljQ+m4zL2wTkMFoY
nUf7PZgCryB+Geviit6codsPz3USOAW4CZlCwSy4zIFqxWZRIS902/eJOYSy9QUd
g2z3LossGlVdTkJyvFJY/8fl+FMQQ+OWBhrrBxQel6qcORN2DqUz6GVVx4EjdmKq
A7iDtezs1qGcfLSQxBtE1zsQLtYPqN9ULMTivkr7eRRVb9KrdRxNgQPpWzdovdrA
4zs1RQptlkrBJI4OUXKPqfKRpMznHGxQ3vwB7wIfXzkdeC1gpbWoduNk7YrE6JTr
kUjJ+vdlm70IQew3pTHRsGJiVFmxxDqGUS/riW/SXgluB8kY7FYIIbC9Y8MIWEQO
gWIahEAEHkGI6vdMoNPGC9YXrY6PKzr2+phI+jDXR7p/NOi3Di3vOv3c2XLIby5g
f69fabKlfA27WO2/xIztFistUlvwhY5TiDhpKqt5bsCtVJAVlnUHRMUn855kq66U
Lbo0drV3rPyi6n7L3yEes4qi7YTx0/YnpqZcW6ae+AAxtIYeJ14yiiyUzC6wI/H+
bmhYmpqXu/UQqu9FvNRzp/cxtVd89ukbp8ZhYuAikcGCXOYD8gTvQn0J/o93FsLe
bg6w3ljKzfFAbq7FlVwSMSCEsaCILJqmPBvAJSZoCVj9aMW22+ZD3KN1Hi2RlykP
W9KE4t+/rF+BPB7hGw0Y6mQGWrTGKucWwO4XPAyFPSp06gq9e6U9itw/d6J7zg8e
XLiO5aGorIzmU36uP8VaX15I4TE0MNHEzHD1/Ly0Et5A93PPwihUJX/AVsH+ZzLQ
A4mBkzh27PbRLaGNCUsYqkfWSTuH4+t41Gmyw8Jy+ZxU6n8mCLLlkVJNtKRUP+0j
0J16ZDT/cxosmyl8RM+HzNT9Lt9/GrnmYvq4pKvnQFqzLaIkQKingCRZt62YyXPu
OjASTZvW+pnPOMXCMlmqQ2SnxrcAijVVdHusY4A8sZ7ZmWxtUMtaTAK7N8D2CEh7
Wr2PcFwozl1xedJTe+riUbFhkmKzoC5G+CFLtKA7Y5cuq8KI0g/Wj1wfVHYB3dn7
qOMChTDueDmKwCRqJJU2KIB/U0zz6B24aGedgo/V151pOkuatwx3bes2XHWM2ZXb
SsMpuhEotKZAHAO6QgH5OqfZFSph9WnwSRVLKV2Ffuitstte+PQAHwE/3TpWGf76
AuNJkLI5MnVA+5rhXrI1jZn5kNWHC0cJXrg/30Of367n5X0o3CNqrxhb7BA8f/JR
/tvFqGTjXWptQovtveIBAnjC2VwrE5svaf3lHac0A2FPnS8E0aN0VXA9D9qH052e
dJQU0r1jQzyvxB6a38CoD3gg20wCJ5fksK+7DhyxdixlLN0FyeY+RR65Cs1EFnsn
Q3xEaUMrDnrJLg4odIobEniVWqNn7GN9dOm1If8njKO0+3F3KyA0DizGpFTTA96t
nsyCmLcPDPFxpoUGGyHmGTDU0gYBtY/8Ooorhe0l+QAOlUEC5mCUKU/qtosP0t23
PjmSC8VVxRyG/2JTCYCDSCvdSF2d89kQyh4jcqP5LMnzKwdLeAslBhqoV8KJ2JZV
iZ4cmUMAmjZFw9oxo9UaEIgmPtx23Hco90+xo3iqwEKQGRL3pX1BClWc0ISL/S96
dZYN5Ij4XqLsjM6j7+hKYinJ0+oNGgTr3Uw+mhKz7wOmHtFPFNXkZnZROQAaLHwB
rGZIdDPIYsjvC9Hoda8BBiIVKglqhqhicHhpr3zqKdvZdCxL/swqEj3s7A4Dsnfx
1uZ+vcwzc4REPPIli5XPfYB8094LqwNcuqBBvx0Gxdc9O2aqiZfRvOsGpE+Um4nZ
m0/x/hoK942HFv9hfd3KZju4rE16ps/VCLMwn203Jo1EwZrSLFkIyjnywqedsP1a
Rg4vumJcMxzuQ5s5WTy45shPTzCl2jpABy2YY+seco1VhlkOG7dDI/Lki5c9IjyY
HteMtNb5BmiNVkzKjRB+zw7qpgF/rZ6onaOiZDkeIl9vWSngQSzBQDxD9Cnc0YVu
ot4zZDTJnDdD2SXvqqoSVEeMrm6sF6hYGHMm4HUzFzesO7Rd1lL9ODffVsVAZigD
UCcfCyy+ZvS0jo/hODgn9wIUwc7A/+leFlGQeL5coBzMDUvNYQxv0Htu+n8+3nvi
M+QiZuNkVUjaTXn7ntkhPWSeDu5g3g8QJXFMgF2UpWmzC1GxSHykKorwb1kuGnrD
VLUDp7+lCE5nHWckh385C2SM/AvrhqUfR1CHmNpoN5cYhyJd/bzQnnlZfyHi79tZ
B9BXWuPClWlgeq8fKGrFVcS90wKrZ2gdS4gpa+qAcL/TZsmGtsl3HGIc1jsSn2nJ
MRJ7rkqOMIKfB9eod0ACQq7uqQYgS0bSHzyTQUoqU18ZR2hNlWmqAv5B62w7wDTl
tEAiN+IqQ0LuIxEMLwJGeVKh/8ykPjqVkb/ItdMoId8pbCaQbVwalTMMmdI+I9LX
4Q6g7iE9SpbWGJQ4m2KeTiVXaKcdPyDQTvHOSs6PRUCnWTknNVdGQ5pbvYk3HNgu
Icn8EvJWZV2Q9DzoBN2kDlFzp2tSbJPM1qV8WHnT3FegSA4wAxPW5fo4zbuVg1yw
oF+pnRrxUEP5TXTLI3ioRQ/FvZ4YT2QxLZBf6jyehAdHNST06mS9cmHPZ1EW8o1r
CCOJvCkeIysU8+V79Ca+Ry1+Uq6NeZ8sunDrzAoy9SWF+t+vVR4gn71culj6ylHX
P28EboIVZlJD6krMRF+YxNQe0y4LeP+To1Pi92qsK8T9xgjmAI3aAYpbad9YwBJD
iysy9zJ6LSTHjlArzWE8CbrMk3ETh3+c5vjcsS15IAEp4vyjfwlU11NNye5ywumh
siwkI4IdAd05kB0TJLuL9C5I9h6iLtLevrH18duut/xnYYRfShc/TICxZFbrBiPm
57cZU6UM0jk1YGXpdaKowhQi6iGuyBU4BfUhicKIY0DODcGYnQf8PK088lbCT3BY
i47yNCK04ET15ufy7TmH4ZpxkTvO2MQGoqCQBx1IAocRLUydzFvN8Y5Y4oVV9kZ6
lQSbHC44fOVO7et9C4ligBCVkcwWv5QKPYDQ3Wx3V69XG29QbwukOhMyumHrzgCA
9r+SbAh6IESmYjtYGh9Yxm+d/hIfwY2h5EhVHkSBREjxZEFbUtRdYmmTo37GUNcB
pB/0ZOFtuJfvPzXfCUDKETFZwwcUvSIghlNFZRJ8ShOEcLRUVuKMkztaRNBfQ6pE
gnQcpC1Ey/LZh5e99Fo8JS6zOUuNiezFEQRo7K/FlJ79kokWvadwl8iaKyS+ephx
s1OaMmvA3ZGm7G0XMBWF2RsFv9eprTxGd+pMKjE/lgNIYPBIIB8M0N03+Xjan+y3
pF8eaaealAqCx3oMQh0CxznNZLfmmYVP5eV8xoR16k8F+eP+joLoe+8Lh0k6Y14p
CjRi+NNddTfPtLDl5RT4ipNpsAEi4UJerSiqVrigDju8sQT1XRHAQ5EOqkuv2Zrk
OzTd/qoLw1lzQ8SHB4PKA/7gkX+5kQ2MV4MA8Z6qeYfUJNrMHm6JDXPLvY5vGA3A
AsoqsqJYJU4JnrJFctPmxc+0Ms0Nf6z9LlpApX3cTAiIb8ehAcCzea6AeH462/Ow
peFxe2dGs5ORyHoW1Wu+clArFcElPjMORJ5ON+/pUXTlUt5k2NYpyErFaenNmvI7
z0b7O5hYfNWyD/kon+7moHJkozOn0cPZG6nlix/G+EE5CETwGkZaDa6R5cZzrub6
9np91r89uBGZ/EdNLZjkTWsEm/0O6oB6n/2ndvpwndS+yq6zuBUjDQDVhx/L7lRJ
8OwxLiqtGwil+13m7r1MUn14uUvDQeSFvLjM/FULdqGdSJ8qKyrCRtdzZ16oIUyC
hBsOpiqhGZjSCbk197KSGYbQCQUhpGF0o2xN0cFKo/0n4SmsYjBRXWPa6bvkQHDJ
75j9a6BYUq5ZqKmLT4RFggPmgNVC09jCMSkht+sjJ9wzv6Aiby9YLXooMPFBqj1q
Rz0OtLVj+gpVD/YQP+T7IBpEuY4Ku8FoJtreCe5X2x6ZGYCQWQsOff6O/LZZQPpY
nxEFbSjatumBdYw2e1Dko+ClWVdk6JPVl4LhZVQ0lbSyrRsGJrmEh+o7rZ6P56T/
0ZU4FGZ9Ms5hBBkM4iODVCh5sFNpwLMcLfs3mPiux6FcvCbMEWym+APR2GyWdorG
KfFawYc08tTDMZRHqry27pq16X5qHyUlyjYCTj3KmzrD+kv1IoFDAfsxH8ccwHO7
BFJAe7VLp0MieWlV7FYxPx8QvcBUKauUhZ76B2HpytemlL0s/WLTKSB19DxvTKwC
ycbI1Udr1aZk7A7T79sWn68FU7NHH3UlT4MHpVfTKtXcaG0BnAfRYJeEgZEUnp5I
/qSJEQsubH/q4QZS+AlgikUhrzNgHU4QOpCw4zg7yhPEXIzi2IUNY6272klzeXes
PsHCpS6d2gI56PPmeEltCIwcj/Dr9ZMHTNxNvB2RNO235W+3p0ykoAM4qnnuot2M
ARFHxVbcL9RkGBUS76wmc6F8psI3D+PcgdcIngOHr9UArEjhvr9veCOfDEocRRSa
13NgJXsR6YqqeYG4mqXpDsmrLH+hN8iPAWvW1EmbIL8meosEiKMYNOO1EcWcXg1Y
rlkL1U4vl90biVVmaZwLjNHvxNgEl3cw8BkOKY0LzjG+2mXZtuqUUDOGZpHDz56W
FaB0DGHUGq02OW4MVlhTQsrcDK/uQWEQ994YhwfATp5McxoNQZNHmTwm0HSvo07a
pdOpegeG+8KJ/FO6l5K96EDAxMQ8cUbD6oJJdJCT1vSvfXeJ74ybxdujKGVfkcsl
qAAoC3HTxkZ4oWrJFA894IEqnpEs9sN2qJTUA8KMBmVyjahVfuWd6FjDfmkWTpJg
bPLwxJ03zQ5RvtRRR0rVtrfxld5PpkFk/c6oAmZV2FPatmLGilgfOK/8RxDcBKrG
rjLAMh2kHO/XxHqY0uFUb4zYbKuoSwkXYLvBgUtw6CW1BAGWvlS/2fg4wj16QmfL
zrFQGDnHx+nbsoU8aJEFnFlyQ1SZBvCEl8ESLfIyBaoEQBUwGrONfXP0I2/tyOQv
SfmOLRofCYugpU00fcvJd8X9fep8o5frKC0cLnGtzetoqTRs/0X/WhUPPj5Yuqnk
NUAYZteQW2sNgUPUQI24Xz2hHSLJ0ErqEhz1nUPYtaGHJPrYgeaAhQOcdAkD+yDR
YLJmdA4iA4v1fLtATnx5ihUJvM0X97JCEIX4WvSTiFQpqQwhQ8bwfWbzd19gCSg1
CIfb2ECsKrk5IjDlIH2bD2KogOqoIBRXznw3LOISxhVHtS/L45sTAOVnvgTaq7rY
6PhklHgACW48wlhkcLDZ0FcTFqga8PgejAEKXvFxpJsOYFYyv13CYLkbAMm3eBVI
yGlNC13wZBAfiqO2lwd7jQPfnxrKvraY+9xbDIVOdLBG7H7oFFAH+WxkkOSv86vt
mdkYZBi0+ca8GDgwKThoCNnrL5yryVmyOnl5aNfTQZRBCeQQRpqJVuZR17Vc1xgy
c0XYSIIVejrPpN0enrJVNHKGdHFaIo7/arJeOkFxmwzv419W9HhgToRUDTIJAprK
JBlHOJ6+x4xFaJs7Dgg6JrXGQgR3CaPycv08Ro+1lir6fBX/ctAQGRjQcDcXRNph
dVcxwMqHuW2L33HpiWsDS/jQK6zRv7WmM9rolKgTrtWY++fv4gCoC33xBj2YG+PB
rETOadbmoLe2exCTALo6KlQaUVfXw2zRSB+pUe+CNAKDaxygWLJ8GjZxmAGkbkDs
g/WNkgAo9kFRqgTQsWsWn0M/ei7XEj1kTzFF0T1/sGwLcciRkPFeE8W2LSA5sb4f
yDeaCcOk5tNH17bUsQn2a045Fza1wQWBDRL/cWLTmu/mor2AayGhveHVRgDymZI7
gaVKSBOLo08oBnnIhnLdAaKby4wHYYuBAgnUKaYZJ80Zh324rUG2Wzqgy6Z/lEZr
yWkdX4sHeEl6yjI5wfle0LAkzd+ac3N80KD8DxEgWnTFcOr5BIBy0uVCx1+z72c3
YWo6bK6nFUxRxB5SA57koO/iHHmD1rep/FeT/MCjsDrLQoLEWtxwbWXpAvmw/PkH
2VrG5HzWV5IIx+BJN4D9X9cj4yn4JEY6OYJZKvN5SiejR4+A9+yP21IGMVGFeS4C
9NA1WsaRrrbcS2DpV7hftpeterc0gaxzARwzKF7fIpqKZY9RigeKZDJbXCFPaFD6
Y5AVxmxxtzBI9aRvRWpv8rLbMRahLaVxwQflChnyCQP7jL/UtElNxKHTXoUpqwX+
DS3nJtH7SuvLPf0rDFq4Ho258ECp/Wc+nN+qvmZW6ngD/2I6CJw6dWLCpdiqiNW0
2lP9KwLf+yVacjR6QCUWLIhgYCJG5FicbTqi0u9sH+HRZ2Y9W5wkaM+jcA8ykP+b
oPMtRiJfsn1t78SqA/1xVt4a0JDdI2AAcGMGqvpke12dgl7x+PqU4QvWHlE3pqvJ
beFA4FVm9wbcnX9l60F1tWK4ZaFLC4KgKpkcrWWV9msCF2JfoNTGAXb7uWJmOMiC
sT0oiLFlCfneVchMw4PAwwpFnR+FW8kqNcFppQ2OPexnzap8zdhXixetU15lxFWT
OAYa5B6cdnMJa+wOOssSC1KzkPNQkb7/ffFzeA8elpTjyLfKLCbc7DW6MThCFv9G
+SiefLLr2pD/8kWdsaFSD6HOthwDO0IALZY2MG02JZj7GrcJKWwRodPvbzJ9OSFb
f9VpsbfAiDk3b7xRBYAmBWPlqx652nsfMO5TYJFLRO3xeFE1SFTq4SvsWZdwSd2S
MkhciziRj+fKEpI+Q/fpz1goo2oYqrCPD1PDRtcFf9S3NkMJKdiQjU1N3//W2sbY
bU+pA170yRg+cSBr5KmeGHfBYnlyvBmfLkCA8ii8rpevT+ooiyf7hb6KCUNMb2f8
Rd/bbuQREydARXJeYmYeD43qQcbAwh2/oyIo786hOS3ELDDtNsojQPM34WeyZpDC
HGs9DQh+t/MOl51ltyzTOSE1h8rcdhdx+ccEaOyJR6SF64Cl2QcMQtcDv03d4Cg5
130WI8njXSTMILf+qY+IB7kWPkkgmmS2z3RS7Q1eInAE7PVqBsn55GNipHz9e0iS
YJMNnlVr++8Z1AB8I21lRSOCaYsAy0LCbORyTgkO7TrweWx0etiT4Quj9XWB2bHb
e9yddR5Y3aa1KIovjPPwmiS4K1zcr0fFjJa98MFX4GjCC5e8EACWF9nFUOtBvJdO
T4YfqRi5XJNp3jMnU1aZ7jGh7EaPOloeU6TDz23/sLTLk3ui3oBEMkbZfYgdgVKa
UEygndON3Besdd5CMEszsRVcYGkPTLjbtr9Y6NOJazCi8lPGp8sD2mkeAw74Yk4z
6IMVdOcOrhPiZNRFud3DVVC0+JZIDRtgABEZxNz1+tytBAmNeXwpLV/UgPUpvxXd
3feZpw7HuOJJGzMbET7Mp9ZICxHxx1mbDJOACCQWrjSSQ9cyddH63J9BvqW6bCnT
RBzTsDJAKbEFEwpD697okpDdL4vUVMUziHi96VZHxDi11LfTSS5HInvAxEeFNMGt
nPGe6cuoSV/OAuejMCxmsnC9Zyc58bBiJ52/9TDomwkg41Kwl/NWZf+3eyEp00/D
SOT7ygazOAG4RyUAgNK+tNuo1kcR+BWPqQLF1nGZIB+fgReAUUs5Yk4il7k82p77
CXGKrQ2XbEA7JD9vBlPxzocvgCtr8Ysk0Iui0tfbFhOW4DLW5LAgRudabqzAa+mb
lNAxgJH0k4863XDLK9qtJggG6p/ACyuQOBfFrir0vXjrsJZjUiIB9m65tDg7UH90
c34TOpSmzcn0ogqjDoojUSbtFRrnaoeaC4YONmFMH01Y/kf55DmYpC8AYhEXiSRO
paAGIcbkbD6bfuw3YSZAgp0hD0Waxp3Z2KdRHQkVNUaxagvJLUbyFLwpGpbTvzU4
J+UaHDHlP0WTVWS4HvTcJ3LEQ3G06VpTCzF7sYmnTYHyvvyEeoxl2EXUr55t8S5d
kTj/PtExhuy985CSeWxP+NC6uO4FUAkCyqQcJ1GuOfLAQ+uhFBYrp9J3tOYseBlT
VFh9pYBpLW49SLZ1KjG6zUGA19UmBqIWxApdx4SZ5yF5UJ7GMcf93XQtLDyKdo6Y
HHVKQiDOoCNdFN9m/BdV8KcBzFHZ6orEUGTYgjE5lqbuL3/izaw0VgL46SttKCRc
0/UrP8buD6jk+9FOdf6Aagne5imVth3JzDN146UZb527iTaG1v5KCAQv+I9z3Gpi
u7QOd51Q/OHOMZ/Mx/YGkmv4g2Z2JLItTv/13QcmyCscY+lpjREmf4c3351NR13d
cEXvx9+fGfxVfBTBYd0xfza24rQOBRNC+bkx9U0shy1NpBBqsiCLOOXYtL83O+Am
A+u0e8X8zSUdOPDFzkbC7pEs6gslig84XfcvBjeRhn/15imKyyydchgueGi6qmYw
5cZMdH7Cyp2h3wy7opozQ4nGc6AgfhJXHvfTImkC7K1LLGr05VXpls65CyXJWUPV
LFDqQaTrB0vmPp07GrJ8aAJsx5cjc9j0y0PCeWeBqqASiQBf2kloO7DZcvuiBczT
OTIkMFqOLP2799fJM5lZJUhByx8uSLWMLkHWlLmqKqRkgdMSoIeazQrkg2EBq4f+
+fF7Yet0T8S8mBqoZtWEEPuYIuUomTryDE8hI/37S4gTH6ppMQ5ECermZwDvryaq
Q3f/KjafgbaKi+UfqZQvNtWIlOQweqq4sNvAwizMz2py6va6h2ReEAr4da0jWfm5
6yVp1lQFRFKnrqnN112Y4M7pKW5ETqfeaK1mj98ufwCtpI6lYv8gAqnvO6xtPdg3
5V5kzehV7Rd7Dt1XRD5rlitudQH+FYT+0hYeyDx8oo0pBa9x91m/uD04GIxO3Oix
nEof3d9tuMztpjBOaBrGg5kyHgL+U1OMMchpB2yRepgdYWkXlHSqTW4oitH98LeF
v34OiigSfNGmXcdatepfqGxqkQTWl1k0JGkKl6v3rQOjj3xY85AqkdGxlffAvhmz
pxBJldCCB0SPv/kl1FRh4khinW+XTyffb+B21LpnTh1JOsrGoryp/rhvvg82j0l+
QRFAAvU6YEhlCKSKfePqh6RQ1dUZfeiaa/Q2+BHAdMMW1K3A1PhtB/KOIN2AdN7A
RjdDrNRXw9bCQqyiMvSV431VnYwEa724W7e8zz1JA/h1jAHj/OnVXqO4lojfc+AA
oZREbeLcQsnrghjPDATeFnWeH1bQpKca7HAApTpdTnG4mKvjP5J/HTYslm9g/2RD
CJFvNUY+ITCumcBNzqMsB65bRg2rbrzehT/keEM+pQhfKiZFojuEVpPNdKiYobyP
1IBhL7mIHjjelIAGhHz/6MK5269xqMEMKYwzHZiRam1zrQ37SWl36hiiR66su4wQ
bMZrH0sdjaPWBaz+78w23JuILEb7iKIeX7b5wn3NdvtB74XREAJM7ob2AURX+8x3
WcKJxu0weREqbhSe4TbBpL14QSTHqsGeUQv8OQ8JL4x9buaJRW3016tmFsqQNQTN
IoKGZwhikgTqriBv2m0mVuQQOLijf0f4fgdaP6PIeu1T3zzSTOl/bGLsyGoGsLY8
hbFu/h/tbw20fEW2SVvSKKCIqc272rMfChbzLvRJobp7mpFZD4wjox+VarugHXPn
JXt+8Ygh1X7f+lisLC0BeznH6RPlI2X98rNFC/TehI1Jr+RyALFDzFf+pPsmReDP
qLIgieRACWQ/+gTVQPcdHrKfKYvBMOTxSDKINrCqWt8OrMA2I0ErEuQ0PcgDNpa3
AY856VA8PQRVQSS+Qtbc4O5whY6x+b9YFwypvRI62cuVexyCn2avDn49Y8rAmhI0
l2ZgAx2vaZxVdV+UgIghIvpTi/Gc1gQADsTVtSP1CIv6LVfXSODtpA2aalYAFKF4
2DzoUKIon7hgs0r4HLK1OM1H2fjo+pqhHRvruGo65v82vF+KuL7AwPB5nS4qyK+x
u8X4o+Y720oftIXk0WRJ8fgMAEu4A/gPp4R1WPGI0kBR0hBaMBFH9b+b94zDKcPS
9eiczZ6N+wnX2t249cpgNi9NLjXcVkfZtZtuN9fbasc8XNUvIiPJWIXGaYce8v8n
RPLhZxzfUlfjFq7r/2OI2TH6PPkfch6zzHUT+M05nQQn+w4/lum03uNV5AIQBZ7y
i+pNesCbRhUtqwh8jiN/K4oWCloWIAtRiLhNbb6G7YdiX+wH1cF6/lgekei6lZQ3
NL3gbQtY7WIn9DLoMkNppn0sWusg6bM8rudzjAzxtDU4LfvxXRum+dg9AgCXFYPL
dEo5upCjctrJTNc19gyuJdxnzrn+E/4UnFeC0uxIaABJtvrHnKjaWZ/c/ss2GWyM
5pAI5VVagW0BhDhaw91EBgk6j2eZCT19XRGB6HznWDJTmA7y34mKDXbKQWA/MLF3
6Fv6oQMlUVXQFf2ErPm3pDDISxSgViQ4Vu9z8VEci1uF3DGAx2XFWozbOTYbsrO4
rcSqDCF5p2gsXmHm6e6wtQr6tIRc3E8s91VNnZ2knjXeeEcrEYBLg5hARXufSu4r
JzuLOR479KZTxJiqoFjObvkRfUrwqBZLpfiPprmqbLw9wPL5UKwcP61dpbXVqhCW
MqXt+dnHAcc7Ed0nUB3f0smuEiAE8rphs9R6uZXPVPCkS5PyKNEuFaZ5BOxDyZxk
cGtf+5GJ8J3sI6W2KgY3ZCaAUfJvgT3PS6W89jPjSmZwGjw1eNk2Vubg8fkceY5n
BsoP8RkQ+n9KDMu54m3BLdTMcZIE6xwidnqNU4uvEiktRwnGDBXZTBunM3m895jQ
yLw8bcCbW1EovKSnEfQyl/6SdOYV/ixfFi037mo4If92aHzCwsZqPJiGC4V8igXA
TZSVxXsaifnZsdz0K9KGhDQD2l+U54/Bb3UjSrJUMlHM8/YgSJbJRSwshanRkxlm
jUaWLBgtS/WVHMZ5LAr9dXjw+cJ7tkBLOkbpxOXIcegK2NE0bf/bOLL5AEZT4YDe
3Cg3TwUe7psWmUDbP7q89mO6CTzzK9VlZHLdV432BBoG0jjoUwet3QZIptp3ze2A
HitQ1JftWE2l5ZsG+4Fcd7N+cSwNB7q402cuMKQ/TOrOQJ9vLL2lP6zWqh5I2ZTy
CItUbkCfqlq9C7+KzOUF32GVWgI/B3IZnb1b8BvEy8eakIltiBsMZYeJVIZWnFcR
cTPHTiROktCZ90LdORRq0L+CNbazyzI+wZGjD6OHGruN6hU+0z5o5KY5EfvFRRc7
EwuphFoleoFwfMZaWEpzZhkV8LMpxDQW3WavVWc7QsK5Fk1xbKywiT/tUuyxSwwe
Bc+IETNnuGAdpxGDScaqdsScetr8P+IaduEsyanndorL+tNHHNguNXMl8oWAU4NR
c/ClH1LPEbRWUQ2JDHpDYagiycUeoIM/cEkebFbdjEnCq+PgREYN41LSzJX1XjF8
9+4jOyJ6lVObD6ZjV/IZ4DgAj2/atsA4MjTFB4dyPZmGRKV+wdnfIXu4b54kdRdA
zotNjjZQ9B0WGkAg4sKVhvwKhukPI289IUgyAkdM5urS/W/AgoBbxDtYxfPXMCuO
P+oO/SHVU8fBI50Fsyokpc47QqltMSvKNEiEzaTIRTxhpXlOICiESjuB+KfC5KFf
DYfI6PcRj/wlnXqOQwLGAtssw2IgHA0FbSLinrLGG22ItlQwGKRbGgnBmLU+Xyt/
x/ejxtl5kWvbaG9sCzrjSgvYAho/DMOyWIPVmJWUfHY6VetitboFVpv1BWyd1zk8
OvhlASXKdOGMzquhHG0djewioiCKxSGjyWlSuc5azmEtFMHi9uT5+ovGmVOshz0Q
+hJgvJogw+V2S0RYY8nTvdvwGIBg6Lut8s+zjaY+G56FeQlZ+kXJgRtty4xUt8ZU
WmX66+YEChIY7PhEjWBcXyTGA+gsDZXtZaXBYyfBMEVM/U5Atx6TNOPvNcO1Kvma
qzOtTEJyjv47aeYRDIyDtK6GfL/N/ZzdKHVsok0aKPllREOS+DWfF9H2KckseqIw
70nIlNXqutko+4AHmBhC6QBe1IbVqYCf6JiYjd0QkKcWMLXbcnppHV9SZsYWgMOj
cARAox59Vt0b3KLJQZXhWzKmsWJHtnOkGbK2Kc7qlcUk5z7fqiCBj7Uf459b8pwt
W3BFpqqhWWondJLQcA+SnHtiK41V5bFMKuBOEjGC+QXQBuQxQrkFVVHQXI0RBV6/
G/eeWN+LwAxgpb2ea2pGNWhy9PJ86g0XsPGbwU9Ja/fSY87NqEXN40pCKOjvQkxK
jop49Qz/sVcr+udpi1ZDv+1/djlRhJzFRiHxVW3kegCFfyEzivo6JzPQUYXRh76q
qwb444ske6qY+yWjolxdE2/uFM49nRWtx1xONDLkTK7Y2rSV7PNCq523NoRn4jMp
boc5IWxWIYMIFENJLOX/wxsa/8NJPM49w4nDUzUqJYZyaQeXuAoN72M96oZ7i8RL
CY9Y17bHXvSLAxr/tPRb/c880XU9PlYH6KSQguZDHHEw4PVm0mvVYfOzyZTTkwZj
VMwrkaB7656/FY/Gc+rZAagZeJeQN4hXNaNd6ws4/GumBEfoEDcgVSwEiMuywGKc
lUrS3K/yphTKO0xmN8LrdwDYBePytQxm8eqbUm2erzHByAFGilp352lYpMhCf1k/
YojjqoycvbFIVe9qLG2rRgrc8SAdch1zOtMEHLX41wVNo8zVPkJ8rb4sIduelXL8
97HdUn+fggEk13tWkn6EeKrX7ALcDxNXz42V8cIOQvSqUxZfqm+znne1AyDA2yy+
31ENTztkh/KH+fFS0mX34+tp++sJtTS0QATXO9n1kRcDp4CipAUhoZHkFnVkRpzO
Ln6mKq5H01Ifo8GrvREgWjNlKBqK1nc8lUpw2LfiHs8yW2+zmTwUqiEobNKtucp5
4UsDuB/O6C1uEVVUeFDj/qy/IsOeU1lRVXEvKKQhXDeQCAXUecq4+U0PdCqtJMBo
Yvvca9y1R0TTMRv57Lof8SdRTmr7N0WwucEwIBmgBogRY/uF1lrgmTMr99lpIy5N
r+2ySYpDg9HXBfcIm/vr6WH/K5etg40MKB0c9eLVZoDanqfTPC+Awkqi1IiRcEBN
XQVH3ezv06XrMvM3kEhi4hQ14QrqHFQhDh0Zlr6+oadQmzJpnkQq35pw76hMJRuY
cv6f7kB4HWJII9v4QmGr9MnbPXWdoWQpYUwxjxf/zd9K2Rcs0EJuIstWH9Zx0Mly
SRt7Pj/MOTNiDAxgbSYlzI8DKNmfdPfOKQhETA7cUMmqaxW8OzrejPqmJHB8cXmb
qB3gAXy5r5tSapVz9ghiQegZLbYl/1CcV8hU7BmaY+oM9GakAhIMyTn5y4ifVKw9
vpzUQKyYYuFFGUNMSOaNBc0EbiTKwcpLxmjh1ai6lKZUNYpH8ioB421xaAzqH2GE
ru1KDSfQwtuhLUk7M1/e0Umsp2hW1t0kTeaksQm4f42HCJi56//Hn5MciLP3RlXI
4cg0xn/zvNe+L5DLhJvGLhWG4Zr6kgibXR8Tw97EmZfvvARfJPSy53YXWGSLCLN0
WIa0PZxJTtdPU3RRgK3+7syYqkU9F2S2fMecRvM6dqjBwQgTeMJR/l14pZAysPNg
SJAwil32EkxgbDt2Avt2qjyb+iV84y+yt4Qnrmo65l0UgiwfjdOw+MfaUfFd7pb9
QkWctJmzjOE+4GJqoA7zO5GraET1g7umdMQTok51MO2Qqy5FG7yfRKFyBNf31qXx
IkIaynQ0nc9Ndn70Q1y4cMbKNQasPiOpvnj55gEBe3PAXkItajr65lSIzBtY5MAF
Gcy+wPo+L7mna6Z4WLqF/KDZkwrh1r97bma/2oNAZHvP2xq6O1tKs1QuxNchg1A+
QJ6170MaBRJzJDOg0DEQm4lVQq3JRvQNRzxJS7IbJGqRAZhn4yH0nn77xQdyKj2Q
JYZFSSpOcygYcg238CgK01m0wFmVYkQcKF2se20zy8UtfgBFcMNaM1KugGvp2Afe
5jgAeD8zJtQvJ750igkuq2s78YlAlmF62uKM3/m/4kyA/fpz6SEKhJ9zyyvSQzbt
5eSg8Snl0J+R9w3LAKUhGivLOjYGRldMrQXhJDYBoROkYpjsJonAa2xDwT+tXl85
pX7sobiWNyuqjQrRaRXkUzTltLN+tWKl7je8fQWcQjhiqmgjPiZCYdJ2UZEA+C0i
epLZPFi+xnmmQUZgkM0AWcRjJ+B69Bu+PXNhsB0DhR1xtGatdfcvxUMC1i9TxRKp
z5l2+oNK7+/0Az62bCx9ftM/7V++K3/ZEiYEgPVEy5A/nx/RmV2xXCdJWLGrQA8k
N1fyhc4in1K6HL4BIsKwgdScwJqPtkVzMLlfRIOGrojfbKnVRv/xuJXehUxspV5h
u/5cq3iyJYyf5ICp60f1PxOhbtW0dOiAVnu1v8sf2EJfMPRMtptc5VV7d7aD1tqy
M4RIaCvP5cpI1SL571+5HgfroZFL4FRfLOxyH1wLxABVqWolISJd0vEirLmYMCpY
0nc5JUcSkem35djFbFYxTHHdUej84wwwANGYlcH6szERdcrZwdYlAGLGtBLat4c4
ijNezndwFoDaaLXPKelhpfbJX4WFdQ/GZuikdIudhjm72wMPIgzZ/GYTKmjpKobW
ndkCpOZx3uPxDg4Mp/ZlHdQJx5CbofmJFZRty2LnyCHtiT/E1oD86c2V+/3Of/HD
8UuIsayXRCMkfFKevXQ3E4/SpXHZvi9f+PvdbX5+bkQDI2iPO7c2f11fmicBpjGp
nlwM77DTtaW3MZ5lVGStakia80P+DDJvHB0FsmzgtkHiwEmE3Xjd6XOxnnGrVIZb
nndjl4cL7JfGz2u4Byk6AKKVjiOYUfU17YptWee/Il1KjytwwiYiioPPR6DVENTb
hAc2HkfRmqELF1cp+u2HzBoMAX2xcm3ad5e1wZIYvnSG1AQllABdL5GoknoybPCI
oDIk9bRtCrU+VXnpzBdjtmYgS8R6ZZyPYMZlwM5udNQqY6Lh50wQMpJA7GrPVMyR
pjnUF5hyCyaUR0xwkOxTvNMa65a29voLJxsrYhk0jL3DdsiLlX9BaTNYD48PW5o9
5P+VFqryWAW9fA8qC2GYGtvGKqd0MKnQU0pe+SJvKIsxDg/7VFEZmEltlyuA7NLz
Pu86uAK5FpfLiBNCrvjCZe5mwCDIS0fa6JgAGtQFBe6fMDXl1A6oD0aYBeVY6aKq
ARsgVZPDmT0a0YD3DXL6NDW3QYLgSRY7gKB8Pt/jY7UfvF2HJysiKOSWunFBtmg0
CBQHAZrb4tWgqvAsSwYAnGIBY+eHt6sLQuMuXw7t7Ehi+Y7XsdZXeNlvuXZ5Rq8+
x8tTdSRGOe2BcPuVQFaecABPwCG6BF9qPpm0OQdYQ9bYc5XeaphIlxHluj6HWdIc
/7boqRuPcVQE5hGuPiJSpuSiePFKNh1nreIgA/fN2TuJJb+EoHhjo7aBmviJiy28
KSNwkTJpt6Hy9EywUCF42A0Ce8uHjPSj3dzOwelEFFtJKs8BL6vietT4RJ0EUGOZ
Pnwx0oR2BdWkt0rXGgOD4kR5J36yUFowvhp/gXzrriq7CuMbjP2Rs6uHElToLJcZ
clkYGmjVXhju+xr+iMwkgWLPKfdJ890iMGKB0LhISmiwt6ar9C7cpM2d+tFtFv7T
mYCkYx8Q/m+KauIH++WLf5sa5czEkr6zdP/l2gzN+FiX/qOP6UQT9s40jSVC84bY
5c8ClG7t+8mkeaZELd8CCK2DKxQpw/3ImfRetdhkqXBIEMG9f5/OG/bcgQxILbK3
dv6Mhb9Le+vZ0iSsQfcRDMQyV/ft5fknIxY39S9YOXEkzHkaFsahF0JIBnYaSUX7
liv1DgtyXnAMes24WutgleFdXLyrrwS6iE8HT5m6jAAwTM8ZgxXIsJ7gRw3jpQhP
tc7fVLYsM4uwfGK3y6nXyHPXBfTeFFal/kXkODlE/8nI7FcQZKggAwHQoUTsKLBn
uHipmGNeQlqMdx5obOGdizJ0hZx5TN6B02Y9+VSjRXdYpVeirDZMbEDOaacOACgz
6sMtEaxh+MfXEEVrX8PGdwCwXyckcLJvHYhtUrVkyTQcQWgEqHT+focBkRmTKDsE
O2rOTwHi5o7N5ioiSz2ox1TUkazaRlbnoEZB05hRCfa4rnYZBl35Dk95dLGU8171
PAd3WFTQGQ/1HV3cTKd8x3gAEVs+lvT+jamWd1HZHqwb4i4Z08oRo7yolpIAAUfT
ebdRdl48lCqObZOjiBmG5RQ0MR8CUgd+YXI+Bcb0pn66qpXn8FO2wlVg9/fPPy4f
6N9+JRH6KvCLpX96G8KR2o7QyU4f5227eOeBKGLtLGL0/ejCffzDTZlanK0aCG+A
HrnnB+/zohaMHK8hrxCUX+Trw7CThqyp5S+HEef5SePlo8O4lWgs2C20PyyZctB+
YlyA/1qeBIn0Q0P2oHS5Ki4RjVNlJFugjr4sh6VIYQBChpgGJgOpA8p0NiOIZwsQ
vfURC3F02KciGAHGmx0HhlurAX4rwXKobCqm93+tMeD50YmBQcaLMIbWDPZYlOvf
53Wtsfy3/E/USN5Fd0JN8+MNgYIJuAXuY5/9/0k7pj1bBgWn6wbVFlDP2hNFrwf/
1jiLjGD0xj87eDdYawWp7nsI1qIMQdyB7yvY8XGHBcvzfvMTRaLn2dBXsC9+sEbT
PxAOToEupESmE1d3dl+fKQnPp1nyU6IreP676pvbqcLIqx4ESxlnvGc9dbpaD37j
oEk61w7GixaatHHfAwkIVfgL9Rz5Enjle2UH4RwE6vGUq6MIee1SmhiFZYyqeN/E
ahHofs3rqRTrw0O1zqR39D9NbFBgn6MprZYZHFAr0E6CpBQhFR5SjrG1xLWvYYhy
EQFUel4rDLyoP0TDPNLZzBDlpnrmR/tP1NJXAPloo7kwY6PoYbPZw8HeK7cQEbWI
oXAp/yHHvfyJ0SG8h2ANFMqw9Np47e6Zbm4bt8OLbGEEa94nKQ8gmRC4CxP+1G0b
wBPNX4o0i3qCUJkfqj7HjlpFe26rxV5tKTFJgzJcvCr4Cpj9vyTB6hFNaHvGDbFe
saYipAg8Dp51Kj/PnwRJZxTzLm3P1EQwOnbm6ia0AuS2O6wdwpRGQCe3oxfKIKBb
CbBUXuaIJPgxSZ9l4MM3Wbfxr1YrkMtTVo1r7t2keWGFv2FoPaJPYG4SrbYfA8vS
Upac1uSF1WWye6kh0FoBsLOC6Q+lWd37C9gmn/Yi5zb8wnPFO27GSGojHdyYMkmN
W/zoQd7pJzJyUys6wXJgZBGUjwaB4NSfl0rZQARf5Fx0r4BgCfX/Xb+9U1QAMJWq
1sfLGP3oYu74ABF55ywMOVZoG/Cxja65h4DnH4EQg3Qoj9spdjMSRObPLnvwJz9H
oPEmL1A1mY8LMpSTOzfRZMLtWq3vcpJagyvlP8xch+emdTOYX1vb7FbHzlCoEjP2
yFpLlBX6dZOW/XDs2lkIypkGZfbuXirt6aCEVlYeADZYx8Gqi/L3NuIn2j79nhHV
uqslRJ5iXqKzmnxsl6COhdu3UMP6ftKc3QP/jP8SpH9x92ABqXGYX7qEfJWKcC79
44w6KV5fz1gty6V24FO2xlF4jCvS5TZw+g0I4YQd5jlt+ktmuBoSebdANBqOGEJH
u9YXIZ36xxcyIzwlHH25jgcPHfHsN1SCBK36kXFJSt2v4fNEKOh+Ol5Bg9A6fjLs
5u61Ot1g0E2eQwDwef5v0eHYrfQq+gMJ/qDLmLfgMWHPZ6pPrcj1ECLp21UdlqtF
nNv+KJ51HhZnlhnZxLnVstnC39P39Lg6LDr13jz0kMLzp2bLrAJIt/Mbd3hVPMYN
TLZ0END6/95dDbQmohkxMXWRXbEQETXDAJgLRVoLFyRKwkXJIeIn58RLSFrNLgpr
7OKndYIUdx14cZRky7AQdY7E04B/rWUDlECKeyw159e5nFF+fvWDgrm9VRIWAjJh
zVQW1J0lZY1OSCTydS+SpuA8K2symks8NHo/EhJu43OkzdaRzlwqLeVJguSgVX+l
Y+O21N4lkc7VH6HaUGdUkjFNltb3zynlRPUvLL0idLGB+6cFFPQYb/rPD6FnhVNw
pCsDDG4IKkOwbvZFGAuC4cmI0MrnHN0F4l2A3FHZ5m1WVUHZdrW3pif5cX533Cdc
Xc2sIcCQ3Ew7aSBGgyobWkFoG1DvloHf1KiaR9zDfPohcPRFqNNa9WTBbzukahOb
WvL3JY+dZxMb17ryyIH8a3P0ph/dSGfFlaaLQpNCOlu+cAlCAJMEB+iV9hof8VCO
EoKA2MxKP5zqfUbVvT9PzWGIkppLyeU9Mr6Z0PG2f23PiVJh2O1DlADdv0u+ojBL
ByUZ8GVkdKvSlehs1FLHtk0Yi1bRysRD8APNuZWgXxwNEqf1QMSMVeiRhVl10LLG
aj/VTwnmK9BfYzQ/lJ+e5CzldFhTXynhTZ3s1BDMoUs8bU0YiCPsNC4HebNF9iSL
zoji+JRznAKTOi9GiBIQmfsmg0J7U9ct3JfF82S5ZKKamOucxj9tiK2anoEgjn7I
eDQ5pyyqZGUKM+m5rUQijK47lOwOrdNin8LcszLzcGhBBubisTal0YdmGclN247+
b8t2UohN34hhBYk8eO3nOWzyt65UEsG5sfunk8bIvYbtcALA/EjwSkc623rIIm7Z
rk5j2/j9zNXVgo4RTokpCpNmj87B0tWyWav5EYFkYWF59f5hJ/PmavrADtfqLFG6
S6+dhfdTxECr7/EnC8uRQzkgiKYwXxara9dj3Gdr+H+/2vcm+LcwkZJZuXrmfvBp
W9VU7t3FjnzRykIOHm/EV3hAB6AixplLRtsUMDu0mS1kj5WJVfNVJPXLUar3dsmM
2TpI5rNSWktxl0+fBCmQf0vTWxlN1FC0BHqTlzpFXdhMY0IWNCg7K83twLftfD50
QUI2Bui3GSczoaX9WhIMOpdFauUq3I+CtGlpMaaw6zcA/KjBMzjYQQffvfHjgpGs
pcch4+cdEZKYtywfsVWMuR5m0g6KsO7wss7PyKLedAXmMBh9rooWXM85WIbpsEuV
xRaWM1qTaZ94bMe/lTOyAI2JiXCuDkDQdVQaKWC1HiwjY1fS2mMxIghzT5y7TVmi
z6A9Qd0rD+ei7x//vAnAPnPgF08dSTmU/cJ+DXW+kOpCjfHQtAJoNkeSP+s9eUfX
1QYxGRWGxzxdcBY95HTt9ehl+q3rEMiFN4hpSsG2+CGNfT+MU9Zbl4j2RhWaA+P1
GLWxIidjmfA3qdxygJ/o5+NW1r23uutGXJTNXoaaWXhU2aUrK3KxV4W6UOdjc9N4
KpXWDwsZvHEMH+xKHdpfbsPb52BXah5LAWhGVYy9vLo0zd9IkwO7udXO+9YfmXpY
X3RzPJgFP0moC538vwNp9g9VAON3do0ixyRqopT8iuAa78rr2x7Nfh4076NNVcZV
CCxiTyBURhgnoeP/vnCQadc9vUecjjKucY7aNaKhCWVQfudj+ERBCRAymbUxxO/w
lLqigYZ2norrhrPYhByLXnkvzwVfCNGF2Eh1oP1icWmP/0qgR75JLehNE8k7PdhJ
G3aTbyjTAlRKY/L6iT5WHX2zaK8f4+4xjZud61e89IugsjwmnYAZuFH90ORXqXIJ
mFUs9zdmojkbDeOHE5ePI1s8tDSP3u72bTjfR43NyWR9EdxGfelwQK5AyOS+jkez
J8JkBNwXJ9Bb0iZiFGFGAy6LrxmVY4Jd1GJiIm7yYNW7l3mpsAks2oClkEUZVcNK
zhTMNlbHoVVEY8lv06BD7FVHcUAgWoc3sCgBMc/Pf3rI9MW9pjduDcSJ0pYEBQ7J
C+ayCdc6/8/OBnNfJBcn6kKQyAgbHYDNYf2jUbfKmMpiVYAlQ1yovjQAl5uRZ+xM
FketzNzNfeI0/UpRIGn/ZThsUm01U1dGZNdi8cdvM7XoVQ4rF6xBlLeQd7kgtyVW
CVoT1aAW/HnFTTQ2b34TuvuDFxIrgzPLQKbZgUdPjA6cxZh2DPk0uLL5gflUO8ed
CObwwwStv20zRiHemQr4CKGqQ1/Mug/qSBCeZ2NZH7imcRgLCQaxfLgXcNf18Y6t
MCFAmWA135OmYG/wfZ0BFGB3HL71/x2QFbIM6ZxM2zvihuMwhMFwkfWvXqoHglP9
2Ha7ptaTpqaetGgdLg60UEcqs3fKmor8PO7HsbvihSo3bJwZSAMsVrPPzUlugpQN
OZTrOvxrH5p06aSBapBwu/ep7v0dyzA7C2KB4FR7R6DJux5nNjkPNmuYBi9TBXdQ
fjmYXZdy9ovMHBLojvzQ72Cl4caK2iQhhf/uS6LS1ELs1xA2n6j/iyKAPL1Fbfdj
coKOdBgZtcaE7Mzsco5Y40p29C8eQQdMzyM20z3CQi/r0rhc0GUqOmnD58I9V/Ie
+EhuRg5hrd/MX9e2mEHIlzTInIsLA7XbSchhh1qVTU56N9aMWAAZ1jaixO6Gj41U
qO2ordAmey2MSeCxKLSVVha0vdRy9InJv709nebF1JepMch3VTt7nONiu7Hwdf1N
iz5DTVgm1xAR8jogQ9lME4NrxC1WTtWYzwcukUI+3SpzsWM3t9amU1oMEJ4Ljln4
GV9y+fSUysdtoB2phrlpFhXdzYB3I4e2McYMYEDhLpb4tUsE2G8DpoPsbIc5EcGj
JS+nmSXlNiu/Kslb2nzVXfyj29QebffAO1tWOh2aSexGV2EagINax1Mk7cM1XPy6
EH6FmnpFlBhTJuLPakDQm9Wkk8J9r0yNx7UOwuSL3aBtVfA4AUX7ZkcjbpdjtAP2
CIegSLGFafOHyu6AiISinKffup1V4Wi/Pi80vbywqhVLGjRhJsx40BMH3sJ+TXQQ
qDM7MOeapPuQ2l/Pd648hPgxmA/IKMHFaaiPdMF+Y95kPq04tOWcHala69DIr2iY
EH73VVv6uphttGuPkMT8wf0ctOzmIJOT6EpzXl+HMlB4n0MYRqpCWl8R+AoeaURZ
PfWJkLq67y3reVtDFlpWbBmFjxgR5nNxUdRNH/RcLLsphZnxzWCTNMBn2VI3+AX0
x2uoffJV13WIsPSsQCWFE+8tigqzHx7eO2nCtTNdF8PEG0q/3gPK6rdFzuoSlcf7
AkBJ3GJLZNf/TTHVkCnyG7gXQZuBo7BQySTzMmAhbjHI36foMPvBJ5J4j8Ns8d0x
my0XZWKbFmT4QCVw+JZgkDZELvjWn6FK+idib6Donztcy24zYvbPiflZhuE4iQb9
SBiXBcJOMsC9zHRXsE1nzXj2y4ZykPg0n32W7wbbLRdKf3fPkawyD1lXlRHQqS5M
u/u+YNl+bT18tw6ovFICXav9rFQJ8x3Ld4YdSxTcExkIpbKIhdoY8B4jrANzYKNX
YyxtRam99FCW/d7kGnxNta5erQSa3yzJXtDeP0xaBid6GtxRgrgZxsq5v+KoZTp7
8J0nXmouZaL+rRGe+aCKDaHK7XSIv5iDc+HyZOmfWq1RgjEVLvQAGPyc1j04a3et
OASTOP3fIRqO1H9nseEpsnjUGSWm41MrLYJD/pNSc862P6HsOnMX+RpJazssZGem
+wmpBtXnxJ5OXgqsNvVbBHcIjCvbSzlaaGdyFIVpqFa35FankXatuQ7l5vGxPqrA
zl6QyIYRNLhRa7TbTj84wwKyq6JpD5HxYVgkBX4+T3ITU+hAHQvSkbJvShIMoTIG
Asnve+/RpYYike9ld3Z9Llyhc4PiJmRs2u16EUifzab/iDXkLPqQ+FFZu7V0zYTC
fcSFN3zyplmX0E51kmCXIrXHhigdZ6uKYOPcrIfK1YxV5+P4y9idHguRXQs+j8Nv
j+k/WAYgOxuc+oKR9nWzahmGBTLp16Cfgx8MgokIdwR56Hz6Y3jTwtB9MnlIvtWE
PUimBhDPO5LPmZkpgXuevpBtb1F6BMeewMKt3J2zSEtLJM62rHq0qKg27Pm1DJtt
lTfZrT9w8K+/kUOe3j+WoQ845ziEeP1Fja4fFwQ3uSB/Jag8T6RKgLMA6Q8D3sl/
By7s543otJB8wbdEgqub/DVeGL6JF9s2vMaicYgyr5Q9NkmVIG4guGUXkztX0iHR
oHwm4o4mzuFNKdGlRvUOH//mR5Ro2mXxZ9zvdRE+lPcIqh4Wm+tlyUY0TQKEYc/5
W34OU2ee60YLlov241rk0+ThhlOiiprUstnTQFmA3cQe51sjVQb4VLjziAWEV0D3
x2rY+QIVt6cexcuBLt1cDl6ey9RgW7BFxNiaMieQJ1xyQfuh/9VX1ZzQHJaPt1xl
TKkkEjEU1ZBedNJsAlRWj4lkzQiLjx6dV5eK9OzKcnl7mQ/ODmso3zcUwrE/UAK8
4ZuTP8RKat+OsXqT57AqEvNn5iGGbZEatDMxDiH0oVrXGCltUiPMymSMSCfgxdYO
dx9M/6kO/rgqEFPU9LFJ5ArVKJud9j+m6P6kOkUXWY9CKjsVo0NCG0mc1FvseIwc
q8cuUlfSYmq0lcYvaqLoojsvD0PpvX08fi6WmfWp4Kk7WRRrj737A8OVuMwxYmnG
GcJQgGtq3CznsgwxMHVWFICf24OwnHor68iSSUOC9HhIctSeQpbftP3wGhvu031F
AXyGpb/+6xZVp/wETbfO778JDIuSTiIdXk8r7pnS5M8Q6p9ARvAmpxLHb3s1ic1z
dzcr5QrSU1BXOyG1EIgTXW1KKDRqFFTEzs5Yk3ZP3LByQGfRlYl0B9ECQ57RPGGS
HLqZ9j7XkDUgvasWvF5uer0X/WipTBinJDR3UAjrdpz47Y5iZXkIUeIImUXNfpeb
PS3EHZRm5YMwfOP9vSuUdRkSt44MKGwy+MgTGoEeO3JcpSlYQ2tUES52lelT691H
QVKMMSD1q3hV3RsI6XHtXTtcY6iK4AKF5/Z3lHRad03cpcfGbu3pEwJk1Nf27FjT
pnpEWLp/cpKtg513VKmTRfXSzU5SB/13VooBTwBjz75cfO9IxVfWapIRNLa7wWHX
QvGsprGOsUSxdjb5TPBSSvGJt3656lJ5ptjBVdfuWgJOlSysDgbhaTEjohhtyZNd
9dgEdN8pOy2isZvowJI75ILacEbC401txky13e1gOkxmL92QhV7XrbI6yXKRcoo1
oImBTbt8ps0oonsEwH+kRm90DVID46hOeGykPzBVbv/HJ79R/wGWBop7f1cHsGLg
6GGcTMtDa8glPpCbEN5aCjSUSkJxpQO8rvjRGDaXrdqfGrr7aZOkieLEknGsOEKa
OXCdNuIz8Nfw88+NSD4NjmfnBgvv9VWihqKltbObnC9w+HKiL8LhLu4Mon5tkko7
L5ZC0SOJgLRU4m3mvNoHKyWCBpXDdMmw+8Yl2c5rGXH8iF36/9muvzilwfuqTvZl
EYnSLLYwnjT4x5jtr8NuuU9uDAV908DED/mqXUeF5u5Chka8tJ5/qjYJgizf5TUY
RiLonDpEZ1/Fi9UQ4LylKAUizZSAAST4nZ17VrqDpwzghAV/bOgj37j2g/D3/9YC
zn8XGeNfCfpv5KJhn5qwG/62IBIX/zIh26UgIl0eT63nwDg2l254A9SAFUTPacei
yEMmZXm1b3TfiYUVz2VwaYy8KlEZLwl/zjRgAgCWdJbDYQswGHDyr80ycsiJhHEO
Go0PRAW6Mc0ZM0nd4j5q8N/X+rKY+vtte+5tkaBMorOYCs1B2/Gb1dHgmiBMdUY6
MprSvdSvq6QRZcWu2/bXdhcPNYBTgPoRLYhDj8YzBj6rANSD1h6PowiavGMezl58
/I5qbxDQQPtSvHs/S9EZ2Pix+KRGQ9d2HayGAd2DbsO2H0WOB8RNaJUxEQignhzf
q96ymskns+OUNQL5qZ1isuVQ0h2hIExOIGW8DWZZ8blJi1IKk7SrOIDM/EOLuFq/
cEFtVwtdbrWTe75Jlo4QGdlhp0MXH44jeVtUKiktqYHwRNoIMuS5GVJyGDXwNc5y
K+z7L/v02+wB31vVYHotnoO9tz6YrpqYpHZmG71zCb7QeeVu7UY5qwTDLrpy1sZ5
tENUWwcPO1HAtwFXi1I2/TUKY4N/8+jbHQ+MBgLxbPyOOKNGxNIZNWNhe3wEvNc/
QND9tsDwkU+CU6l0hMa/rdn2s5Df+XBN5G/RziiMqCxCl8az42VpGpGz5sbVQ/2j
lFerpRw+/OWlBh9aIwdvf454HFZA8Rl9EkDxmivLN3AS6SFn8S6lqgHvdoAOhSDb
sR+QSvdTesFAx5u/1lKednFqHl9T2noWgD810lITBbG0e4fB82s5umO16ETNppJS
GRTIOER8rru9/ONxrnCj+Xc+JTA20OSNxX++iK4GhribkO0D5TDIrf6vXNCrSXjq
g3HYyR8mJ/DTvj1sCTowHYpsNBYHrB6ySblB/7KhvAfQAE/kiOC1Fnx8KKze2pwf
PQeANaFMPoCybT0AWkmTnumpBAQ7Z46dGLi3OIf+0oWL5ISTS2+PA4GKYCWF+0NC
8RF6ZbIfiIQb4E7fN0qjWyFHLoSX2U7nULbkxg0a/EK5tKlR4XQ1hC2LU17CieL9
YWvbHjpi0lHR8MMI9ViJVvEFaEXEhLIFTH+uGHrwns0nfoxr7QIEPiClUMpbZWtU
Rj0/uySUFkpByu+ZlWbmYpBNv29RboAYTjXIwsujraQDSzrq/1s4Rr9XyNqvYtfl
hG9X9v813ZtnRkIXvNgCYc0JukUBSuSNT6Ff4S61HmDojBULmtT+xnuPhRnuIOhK
zp3lYAW9oumKgrcKhF5PMIqGqnrXLNG6R9QdVdao+NY8+zW6zW3g1pcIQkfV5Vv2
MbUvaaDEZahH7XvamUK0fTH2XHhwFBUffNvCuoGLKYiEhwwMCL+0nrIgUHMfhZAL
0DuDSJJh5k6PY6PMv0I2hwcCLK82ocTWwN7o/s8bXJlnPy2kdGc8dv5U5EC5ygRW
KZNzmxVksZzprL0qWNJFICZNUE0565c/Lf3teLwUOQb4tYawiqJsWvntfPR9oQmX
A7SnBLWm1qx6aIMRQOb8/TPJYcUAHJ8GXJ0pno9mEuq7IjPOvYNlh9+Hf9/c8iN4
jEyUhsrrImzyIXXnS8DkgUX1K6xC5rZLB1Yl0rfuC7KTwm21zSZM96ppgemp/r3D
R2bSBW2vbq/lHxzuDL75/A89lp3oQOGEfd6gEKIX7kqlXRxoiUJtk+lneb6QU88L
nGIZGqDJXaEDCXvSq54N+GndCv8qln2Gf2wT1OqoCqZBnSRqfyJNXSj1xlA9RumV
vY5uClG1thzbbdXWgRAbPFjHEhUGXcx31hKJ/A20JJqAnQGmuPBmngmZe5Nk6kv5
3JeN1EJJgtA+7SIhZL5WgIBRg7HN6+tzPrxTShNVoqiDC3eFr0uMaL0WfGGPAtEL
u5rYC92+LqzuAcV7iGHwFfkcIN+GPbzC1W+KOwEFZLF/gMveyCoaRZi6IYdqBsWu
G9atOCGle0S+OXzlemgQIKnVtFXJNLDd5TUaqhcRYl1Hcft3T6ZwZ/rpuS13DVMb
M2UMgUM0179cMeEZrcgEqgeIhTXsOkX1l89HYh1bJYGXFPkpbYjAVqcaZAsDQo+g
o9TKEEd/NAJJ4DWD7WNELmEaYw3/mgEt8EUpYuSouZ6SrrOY4Lni3gnnMWM2k5mH
P9f6y7QxEkB5NO6DUvDw1haEtKMyGVZC/tOJnqjJjS3KzxUXTpET9cksj/m8Abve
//Z8FoRe/uLmCCr345aXWiZJxbry4QyQen9Hx/lauHnLgHtTkZgCSoCJ59bHdW3W
lsI8fKgrS+EZFPOQLzKeKy1YR+GTDaqzqcU2ew6c/elnlszdEB9lNn4HYjngt3V6
jyQ2H8d/hupbw97KscuNINqsRC+iirP2y3xVhoPUlXFkF2HDDkrqKI+DcYrf+OdW
qdPyRk3+Md9towecF+VfmvyTXuRHkZQhD/y+xxnOyHUPh5aHz5FzTDLo4olUxCua
o12kYQUCgcYwl/tsRJbobHxdbsrRt4CtnJK1QoNjOh8XyHTdcmIUIaqxYaO08Jf+
mpMi6V0cbqMcriB9yPRDng8HSr8M3RV/0WSKB7zp4J/zDoJmR3gIeWWG32GcPSDw
HZmHo4DBXjCIc5gl3ayMaJFXavRgPMrDiACzkBBa8PeSZzEWUFgdOfZtJTNDKQHA
FooE9uFUDHzqtTZ58RpI2hkj+TgZYW4P5W0aoQb5is+MWqi9e8xHh/XNv5QgPubS
3YDNYdiARWvQ/tOrtsnDpbaC8X/8FbFBRHoZrER1qt9z4sYBgWcpu2UvDyMkTTG9
Pl1yjwoHSIJFInaAGc/vUF2V0CZmB0OyMFIErtrks0lkTf/mjIzc9Q6CMtU38gY4
GSsRPqCGi11ZYmhLIBGHiHN4YSWdrRZOqsVX5W2q+0FG35Ka50mFHQjaK+7XMrkZ
gqHSdfJbYX/z9e2VG9ZDDy3NZcN4IhP5DUNyJxNPjr9fHEaec1t9Vl1YrJvLphPj
gHxjKY7WP0kfJW/TQA8EWIXcUyf8Mia8BvZzWk7RrdOvpDpLHzdeVlJsKru+eWvs
jF1VKt10Xhlgg6kR6UB1i2p647pCEr0bA8h3+VwOOyA0ks5LUuj/Rz4Wci3ysSaf
XSEK5Id9epf+bEdPLjUHED5pHpvZBBowUvz1AumIw/WvmYZZDy1723/GGNQ3wJax
dqUdAfBlbCwm4vPzdnA8UPcp4hRFbkwye6CuVTEXltfKULpA0BdCtWcwpCtds5N8
Lf4mf7qMnxJRKnQ317vHhkMMRMdGBMcVs7S9z9BNVLabRZhad2Vv4FUyVOLXT7MB
VjSbW6lQEEngY4UUC71lk8g5KOSmJ0RxOuqEJdqEgA0fgAiLMD6AY+rnrcl9xOda
OgjEvuqHl7p1KRi1CG9f5CWirHYbC/5hnAzjdQnZg6YSbd5ydcainaxrwSw96+1f
4hl/6jGwtMekuHPpBJ+9sJkYtbC6RNNNF8wjCG05zgwUV7TfT/vO5ZyiF010Ez0U
VnXpk5nwlZyL1c/bX6TwJgIMjP5MRGBeuhDIok8Rj+ZBI/WsYQIpvv/hmS1D+Whg
5UFf0Bj71+jZm3Gd3iENZs4lrOaLHfOfhkuQAwIT9Ada+ZusfJL22n9UH1HPrccS
2Sja6/pyXphciab/cJPw5OhcWFYNdMcGRsre7URf5E2iuWmKvnbfZkUsev5niP0T
fkNwOAjo1TtTsrV3lJ3OSLnIAwHT06w/Pi5jBQsveulE5k3XvWDync5C5H95K0Ro
0e+mGD21QfKzLgZv+nKv5saEkLylVpjUmEA23OmKFcBQvByH4GzZbBYvBiVNjEUT
2Hw6vK13OX5z6mYnVnQcdRok0MDlBR1PzSIUpUrGjQgXBG9zyp5n0HDtGxRDQWYI
58nJ8enLfUMlnwdc+A1Fjc/JVVmDaPOhbHoUsUF5YBXbxVMOfZaZAeLCeQEGWXIV
npAg+2xsUTt0nWj61Y8YV/KRV/88OcEtkp/JoW7s0GJ2KqV54pqiKJ1ctx7oO9ix
92VT4lgEjXHIYqfj6yGOoqOdwG31i1mMv1Eex+WD4PxGoaTFqDsutntfEmrls6KC
YcQ8dsDijnAkd05o8UoEImQRPloaMICeR/9uw7Z234pbZ3CBnXBUiEd1G0maksMM
xYyr76PXRcl0HQqOzW8wzsXat8u82qHNCpCEtEJZlD74c40CDVfjUMFyG7uOMMj+
xjViMAyPXyWIVrqdiEvIAt3t87bxCH32ozHJ5IyA+GP3tSFbMKshR4wGDkYIrUn5
oxOWnhcAdJh+8fj37Ewx2noXceQI9AdHTW5ehAhrEoNZwi3/eH8GjfWDco6Ozh8f
MlvFILkvDXs3dOtJc61n1u3GZiU0W7QlMTxgHjeTtFP9JrRTFvd5z5hCGhpJMui8
zFC0ySB1lGMxkDLT2C1SqyV7jf7m4dHW5P3AFbiwnbRbQO26iNwaNgUYlAPsueNa
pI8XJH95KZlBWVuKy3iArMAxMbElODrtpqJQ3O2BlOIiHdgkvdV6VSx1DGgsIdG0
1OdWAZdeyH35RoS3ZZY+N/YQgkQdl2diZF9zasAwluYCHcPjgqAq8j0y7om3yo1Z
+b8Uu00JxFcvkV5JU1HfFH0RYAln5EGsWqbdkJ7XUKaKs63G3Q+kGZ6d11JCj3JN
rA59kfsIUsqP6Ftxi6DwkNeNYViiWHKLkkIfnWlLvw2TzhvlFethMcAPTt5MWHKV
D7J32VRGiSOdCe/R+ew/ycDU5Z1R5T/q3gjeDwcevvoOZoSj5D+/FAKJrcSJIj/J
54zTsRABej+FfDSrVk4/A2pXhOf1XZdsMCtqYwWhOYd7h/noaCgd1g0e2oaQfzfa
Aac0cydHsxCEdHs/yuB+7JRzeZU0PyFve5rdEPsa53ttihOEe6B54PqXbamigKYZ
5BG+US+W4S0DFbRJV0f2tBTzafwOrR4ifiZhpftWytCF/9XQ4TyXS4DL5hqz+Y4Q
0G8HLTwWmY3xTPaXixC0g57DYUxietGbZrfhOX5S/1OlYtxv6TdhdYvsVUWfEbvj
RllEdiWA/xjXoanOqxev5uCaT3TQqq4f5S8UHg07jfbOSMTmTRbrFsJ5fUrEuNFJ
E5hThMv5XGboYGz1gb54Whs9003oIzYrLQXZkAiZSc7QHi5JKnB+RMuF+EJMtCIH
rSlfl9N4pMQxcU8spHzqQ+pB3E9BFh4/XlMmd/9cTfj+3OArdkCTMn6L7gnvM4KA
7EyqMn8D2UZNYKMPUypI2IkqlnjfvfJkuKD9PDOFqkwuIx8Y2ONgZocxHASo6DfZ
xwTXYheQ8XCn1ncYc6xxB5A+Q3X1rVI2oYDAEuaFieAQBeYX4bfb3Px4EMTJj6SB
mknm66PZqRqDmYyT2NraB5U/9HgZA4isX5HO0Cf4Vx3oZFui/3U1AmY7tnRQ7/Ab
0HdUKTQbT8US/Gk8K/0BCwnXU8SBOt/PfNk5TNNGA8f02QI9wJlXHl8Y2txTC6KG
dSzeaoi4BGxc5xjBzZ1kMeiEkivDaOLkvhdd3ds1u6kbd15TLTVLjokGNFED+Nvj
iBxpiahB80bYyhnG7RzAZcERtbodHOSJu4rNChh/CrK7e4h6jacCEhsd3kRgSgH8
ZLUIVWtAQwUmD7o+ACcF3SUyR5bz7WmgmgepOkz8wGSe3Ikw6w/sBxn7zrF7ov60
5yYVuvnMG/pyg80pmBMzctLQocDRXXWzJZiTMQVWTh+cRAx2UvgTc+l753X2ektA
W4FnCMvQqcaKP+MdFlyj68XaWb+NaRwoL2LzSr2UJG9SsYUIgPX+B4MYX9ZjWPNV
aM3WmXPtQ01umJ3xsI+DVxbwFIk5FCOEIMclc2eILPXrXcLLkrFcEGi61IFtbzXs
59DBmsA5UOH0a/1E8ssXeXE5GKmFgtsezP/TuMAhDjcNDCHGtN3erRWcQ8j5F8wd
UIiE1o30dpLP1Lg24e8D3V0pxXgx4QONa6jaEU7X19VLW6evU1026W46IOq+4iXT
p7PXWzc2H3l1aKMGG9J9g8wkSypTI0zOJpgJdieIM2npY0of4TqsoyvcVBt1LUkk
fE+cZqpSxdICFXOBVIBNUdKh4N/6BVZsSN0h/5ZwZAJtjgD+7NjZm+gbn5ljYrV1
aqijYRVmAjDQ7vLm8+F1yY6NqN82ZXWeTSodHNxgfHin8VRZfKjXdS72rUtT4Py+
Y6ypKmG4VwlE8UKp9mSKb2aMNvI1XpQBSKO9yYHBohUmYmTHW964i780bUXW/t0t
M+eReJPTWnuJ9Z2qGYnyNdiIwnLJJcGIgVTh2EyQKwMUhMY5ZWBM0TvLe3h+698E
0EBw19WqnR3HqUKpUZLAsuitvVnlda3qExy9ORgMFY+elc+g+9+weGUi7e2J/CMK
/oUQPQMuIgKI+qSAgwVwjawztcHyK2M0ICEs68+6xOJzPhkomd5P90zKfTXWqSoI
43TWK6dvW+AF0JIy6ocAajeZi2bl4tcGmvJmPOXLfURUfzMA7AIpyIDM0tE1DXpq
OVoMPEeTaQFTikzhqXixq924pIw6LoR4HJILDfUsLoSBcjpHw6+ievTmNJt4gKjT
lRzGD0b8JxF/RAeL6Y+tu+uP4vNrIf9W2CC4Fi+yhgW/VERw+M4iiJYgjBWqYZCl
xZgorR6f8B1A6pHjQLBKtRQtWkC4CP7GrtJeczOaLPAaci5zYnXdbqdg3uPQc+CY
E7A7IeLMeseQSDColxiZvZHSfXaSHUPEjywNoVDgPuIpjOV2xqPZ9zzVoCOM2D+M
fYKN92f4UXWh7S6DOs+0Y3gy+OOn+shhqbKS3wi1d/6WdzRyqn70oh05dLe4X4Fm
6yYplHuJHmXwgAhoMSePJlWse7GUMTCZ0A9jab/XJrG8LhHXTIVpgu4alhXP4pdG
PKIcRtIk3ZpRJ5CeOJ2U3HeR7Kqtx0Op3MTkFKZwl0mAUc/rS51JCee3Wscdlcvk
MKSm6CniRd0huO5QyrELvizHhoP76J3WXsllOJPmMoqsDyEUhjsqDHqMmd52x48A
c2hbWdkRNP4UswN8vVh+pTlWPk0v0lRZjctGuybQqOHMMVlYKUsPHYdxo2gvQSjv
/2e8XogZ0bACltfBVBRAewzh3X/KCrfOfKwhdMokfV/DrINdTY+/7kvpc2XyRS45
KSN3zPgaYk00vJ/pYLiRXKXqEVWmE2Fx1qbUAEU98uTSxRZQbOK17NElIWjXgakw
GiVXkkP5jS7s920R43y0TYnGXFC8pTTCYBbkI8p6UyG+TFG3NG1bwGmLlDBtE3zb
Lg4FaWBxQLnM9xfyAnUFZOnFpTK6f1ZNGKcy9hHlnTB4wVkWcI+cEECjI1kUYFba
2o+46J1YZ+3EH3Ah7OofETayEyxFWIR4R+C8VQW5uXdlJCwdwNoqij8VXSaKJsAa
E/23wxQq/hBIW7vaVW1y8JoP2V08o+xFuNOSX+ck/0FuulTeaTfyoodygi99gPX0
8gwifNdq42uVWcRJ1kDwU/8m1FAlWqqimbFiDcJIhZXb9HjAT2eaRx28jCPiUD15
Yn1+haxjgV2/6RT6CcnP0Tx7EMjZzyK0no/414pnydPBZmn9I4ccZlCT9knyKd+t
u17zgoQjzozXDpMieWY8nPzp8wGmkIIfYBbRWH5SzWDVOwZPQOZQkL+nSZ5plVCu
Wd+ltYFssH7V2e527KGMKZ0oCrXG39Eemzm+Nl9dco7s4jgLOPHOoJo0Twm4FphL
nT+t5esWWUALjRIibJgPQpeJc2ylh5AFo2zFz0L/S+X3xejDDaVXofVJUyl+dXYv
lQehLytEDO46qcXMJsQ6EVkh/Cqj0Qb1XkIzdrzs8KRzXarwKltzoPAkhCUkUVIm
clyHUe9Hf/t2XHi3TCrmJDXf7xfpZ6DcfMEl359gYcTEPmyzTn/t0IDlaYOaeV3d
mN6Evx7YoSellqF8uOqD7rzqedOwVdtipeci12zcHrndPpdE+mzzp9s4t678ypCp
53hVrWIzT5rFknEvpNjkCeXjqts15RG6+IKD+2zejjsJzga1XiAeRF17GDI8k1ph
qaPDgifQ5aFawgaNQ3ryHH+26gheTkTCEGRIuuzXbMM9NQqBb/nN6xuYg9s8qEcA
2HzPR11XKa6MzfO9GySYqKV8cdXfSYi6cdpSx6/489JUBxHJrVcqobf63vaLLmN8
yCI8THbApooLscTTR+drRqgteot6Zql0ww86ro14o8QvvZwChiYISaWcymb1utW6
Hq1QgL+HOVPP3tkoleGNlow+EfJAsaAipD7psgHoMUL4ohU1wUzye4viM6g23FdG
RGgwS5na8A/Pm0iAXyOd+QzyOy041lezSgOh+noor11DFeVlLPHIwtIyV9P9XfU9
o76avRU+k7sgLN4yVEnXqQd0bRzJxqr3bDo+J7n54Ytpr5BL2o4hssSwueZPe2Ez
/VYn6JTYW6grF58UZTN4zZ3+swANX9WXIlr66zFXc9qwBt8FPH10aH9C56KsIZyv
WFB5PyLoALYYT2h29hb8l3mynwg+SaO4quiF81FIVxdRQ8ktlulT0EhZW/NVWicO
RbUDqS8SqcFj3k2thIPB3S2A4WEAucYgyA341lyW8l5xQilKMlsNR7TWxzmP9TEa
GK6hlOh0hnOZXKuzYxFXhwrrj1opXVdnCyPlSafBBDZS79hBB7IsPdZ7OO+YnUkM
FBUfX+kXiClqQa+FBlW/jHDxNzoBeXF1cFoBS3DeHnqQheM4XTvguWevkw5KCbXR
XN6I9KHPts1LFuVVwTuhOBtS40TP9sBMjZsPbdUx44UAKeJ5Pfwh+2u64eJI1fuk
jd2qNtzOcw7n4QMjKnMAU7vps7S94vPyTAAm2BEoGLo2pLAv8i+hgdO0oky3V+4f
Hh0Q5fudSUBVypouub+z7RLCnjAE1+uvWzy4SVEPUZ8V7+zrP38mBHQ+ioeKJ7i4
brjouhXTZCPWM4qHDwheU9yYAH3o8k9upP1RR9d3FGE+spz7OhJIkn/mFkJv4E0v
cnaygumxCINETMtPgtFI6pr/q0I/s08HPz1v5SDJ4JtKHMYO0SUzSXDTQYaR1LHi
rfBSbCQFLCTh5cEUzwHCtPQ3x373ICz+sY8YTka1Pk7mC9hBbLd2gGfkvJQpFK2y
nYQTUYlbVW41keRtv8AZucaOAWSpmfl6Y1fRulDHR5IqqAL6vbglIMIFv8MQf1BW
7hGM2CscSSjKtyvVgy88Yq2MfyE5AsSKsghZdjUJOY/QO8G+vK8f8caRtE60LXRX
acMi78T2cmua740ShxYKmPjH91KBcUQubKNTHZw6Uutx3hzMzFUFCP9iDKmyf7+m
kTDegcSR1kSKEbvsNFczp4f70fUJfER5WJ2wVjJCazYSLax2acxgiLm5mliVnhPt
XyS7kg04FmUJYgPlk2Wqxq/cpN7Uat8BYAPlwuootkAdH5v+X1BTp7rJXV43KgMf
B/smZYBD30Qb9QOemXmQ5GZ/zVDEbT3vqN80amh5fk2Vcn6OzZE+k6PiZXMc6q6p
nGb3gIXoxAvfE1TD1Xp7X5xdkeZhJwDNVgxxzmEMT2u4IHRFMsJvQOFbShrXaUHC
QnCrfX45bvFNz0eWl28eAnNZl/XPRvu1B8pXHa1dT2L08erG9NiToKcwLKk8efLj
s0Q3ScLuHOXs4muxneRMi9ZQuE8o8PSGtWC8piXFfCPE6B3UYyKvnb2XAIZetzyJ
7p6e/vHuR3cBBp9p2rcus5vIX9sw5B2ENPJVrIKNgLewYFKctkRrSMTkCHrdJolu
UmD5acYYN7QF/qVUzesZXCLEjhyDp1dbMoeKefBPF/4V5xD211zW6YycNqZgrrtw
BjAMKu/ZmrbDRjKrPpAtXMV7dse5wBxrKpBudjY6izYmk0c3vX7M9DsjJ6GpTOnA
zfXlnR5XuvDrBdhrUqtUwC+cnOoz4KDBwRt3VWkbBqWUzGVTIy4dtM1mPCUHrYFr
sl3JpY3+uhMDBRsTyPHfiDWl1zGGy9vpmBc5IbrLIPp0Gtl0tJKevJzb4gMWohaU
OVPHY1HOTLSzuoEDTjYIq8H2qenrGWb2G+Gn11UWdc/C/2VwFB7YtGyd+xZhWSNc
z4HW4DsXjZKOwdJmNegi/gxU7xtZFqKLlTFyEqZdHxrpQJoza6Yo1yPymDlY5qEg
MQ9+eJB8AGL2d0WwAW5JY4ek2+CSrtCqnmCjunZYc1i4ylvxGqmNP/uj2y8ihUSP
9DqACG87ze7B6ElUDuhzfGMbSZQjozeKL5c3c/jrceGTKQHot3muHQdJjIzCHN7F
bN839n2A8ki0JxIwFoHkMPSLLJxmeci2p2p2MBWagmg3c/ctvX+fsXbV5wRqa9T2
yDOssPFU0m3NYwCTVcIj4sx3vMt2ReIgtR5hW5kqkRnEDqQX1Gl2+R6YDiobtk5Q
RRVGxUZwyOhyrshE4jZvNYsoErfeQiEdELVFHaAYaVa7F3jkIldpLtTO5SlLv/4S
zez8ZlvARYBUlEt7abLgw393OW/QgCuJALay46+1Dw4sCj3sCA14bw0+cVuQE8K0
tDXeprSwoF2//gzZiZRm2TpEA6PhAfGzdrz1Orl7dMGj3rVcqsZRhB8f1x94lz1H
YjNuLSxELO53hqh5lsNbyn/QTc03zh2v7anwiluubw8tY+EyJbRJACTh959uiwRZ
k8oI/QU80Nw2C0Y6w6QavASJuxWSf+Ut7w0p7Fvcz3pj9W0YpnEMMTtey7mvJUmt
6MiGqklrgm9elL3SKJ/kUwaqOxJl0ereaDKnabSMhXOvyA8bpd2nzJvGjqF4V13b
77Kj0TIW25x3WTsIPPAR1YvCJqrTATXtAyceGYSW2tuHTDRXoF9Sn72psrEQsfa1
qtRRN7XeFppjpL/b+Rj6OIrDm/LjFxuPPt77TllpJfPnPHqV97l4RloC8R1dlQh+
BM1xMEhexqOtBrAIYZhmou/JiRPOw20NQNvBX2uWBlNCC4eMn3BRktqKolaeQU+B
xj2Mlt+V5TbEN1U/H7jdL7xoX7aQhqms/NFGW5iDyMLZ6kZ/hyZZgCK5Nu47Sexk
t5kk11MxqqBwIOjw/wBJBLrXcY44Dc0K+gQY211ZvxRQO2Jj3PDB1pwx4zkTsO7+
4Kj0XJ9O6NVDQyjqeGbOzwXxdTqG3qt3KcfyI75j8e2O69WjjJnoCyjVRofmQ6jl
NZwR/I9TfPsMjVCgs3sbImrNLiniXNCOHQLxl0yYU3IF4lbHsh0ofY+FAobIsNzr
crG7DLjsp6py1IRTOeePb3mgjiccM7x9F8CpFq3/uBGuI1SuQSwE+zXLgcStHQUR
xecG5bJ0t/rQFoOF7y4KngtOVUX1Zh4TSWY6gh0GoS9F0ZfJ5JoQC88IwN71JuYY
qdDXFuvF0bPjbJbXdJxLFqpvHCFH/vG3OWYoVT8JmffZoPbamC/nPCAc3VlHoWvT
MUE1QHpN/Th9usjuZiWE/DhK0WYD/RlD1Dvv0ACHJu3df/x/EXSeUhBBuVuspmsD
V/Dc+vGRL3fYbD34DDxOrcEkquzQ5ltCpnM8WikkOfZOMxOCiF/IzhX093X8f7ME
vGYA2bYzsaUyaY+16CBKmez7Uxkqva47DTAYLSZ+gvNjK+nGw6hKCEs4lXlcFfIk
PuwvgEFVjHNoqt4sHcfIfgaghUO7LuBQ4kQgyneovNxe+D2L5mzmVoo8WOOzJCPf
Wn8hfgk5xRpu7xmXwMMNnw10E4EHPMyVJCiqw3jFm8FxcrJ7QwuCXiFAj6DXDqwM
GcRs/qi1VZw0v4dRGorxPMoRUxeApMCtkw2u5NAXcUGA0fxen9YLkKI4k+yuw1tk
hmZhXo4Ks37WQWn1Mg2YhXcIzrc98RfETMi9UGxJlWYalN9jMA5XQfr+JyZSCLOJ
bin3z706PDrglX+ws/qIzMFTQ5N+4sQj1vQzXI5AZofRVxXF78ufeW9QDbHQailj
7XG1/d0Ysm/so/so/GkMfJxvvU+9+kZqaKWGumF0OQubk9PWZUudD8KHobhmJPhf
Pjyr8DgYYhEmy91yl6NHF4yttIH5V6wWGH8uvFUZaVqvqN3Qn2Zi6dn3sz0sE52+
vjztL6Pup6Qbn/vHe9zqJVNL2IH/h9GIuO93y9Eutujf9VKAdQ7TGO9rKrnObL3u
x607i+3HGlx0/+XbHyMH+krGyc9z421McORRMbUeTIFXlJMUIeRT18mGz+EodGmA
pXfw+wwAJHUVF8jBxddnKt4r6j5BI61xv7ycOGxaYyzSo8+KeVfrGjpUHflNxa+x
LKKDiqs9du03Q91Cz7lMunX3pvyK2CHPoatZMZ+UV2dzgmOYNw5W/r5REK/SlCqq
rfDVHFKNssG4dLGtr2/3abY8abKr3aBvEcu9xbCTPoBOSmzf/mPudPtg2NlBdj0W
swwo8Smo9pr0FNFheGKORKBH1bQMDtskvEGWYJ7LGNAsiS1EvMTtzfHQf+XZT4f8
Md5jf4hCvPPMoABrBVCzNRrJid/Gdp9wSR7ilnfvzO23ot4Do9+kNlpqDq6ixy/5
RR16UAWz9oyJcr4CyTXTFAGOMspUqd3LiIGN/Y9hBjtXuAK0l7/iApA19NwHLoGF
eLv5AGzd99gAu+pheZNgO3x0Ne5s0DJ5E+u8vXcQwFDLcd09D3Bo8UTBnO4xm25Q
73udEdCMuKJK9n/aYn08H/GalY1Z5s5Z2XR3jVYxwbvkf/yaXq10C3AxEj5aZpBh
NCXOQnKE1NxdB9sBtKoDtHNol6azEqLiMSBy1dZzhKgRoGn0J4nE3SKYjY2SheHW
4LxwXX9PLQe7DKW3oI1772DcgEWwxXt8O+WtMfYEbaVWeDbqBxRmJCz/qGthEaZr
XKN5zzOGJTK5yCKVelsR39ukqyhF89tZmA0F3Fx8Cw2WULuyqtKXlrs9aQvSG8s1
1etBtDdGybV/JBvtxSUTUu4bD7ODDFBYLExBmAJaJvoHfN+J3NE0hGMpI51vRjTG
2gkhcCXJQEm5ErBz4bbHxTlFpSccByyGC/gZh+Xp2SmeBDfC4+xf+RRLrNA7cDGK
19H8Qxh3UXOoONU5WcfIbt08dXfBwRLYk04HTQdrLvJqnnERzz/2NxKO3NOvCOxA
NRbgZ2ll3C6Q/xb6Dh+CJFwZxoV+g+DaQle2RF+So4hKHOeHD1NjEqsDMJbwB1v8
r42MQVO6KD12Pr/Lob/w2XjS6HGpIsZvW0s3fl/POhZ2GSGg6pB+LtrVldidhs9M
Uj/++kLIRvyTFY+gIh6drGnui7mn1o+boBSlz2GPJgnNlRns/tXb6LZ2bn2qDVCJ
9qp5H/Uv6zZAwf+5f+Vz5TgvU41LPc9vrPATGXhshbzjbzSSHDbvGeFxs8xlMS0E
iWTMVf1M0517T4T3R0PL6QMGagipJISZVMevp83lVzkVAqbs3zS28ONCGDs7gIif
isbiUAVN5gTdaOVzhdgiYmClhv4P0Hbk7ZYOi4kuaIAdaAhP/UV4lmzpjdhhEFbE
5NV8JPkvBpSZFbMc/aNhMyfPLwUsXBW9vM4JKDfVHYd958LJ4qk/gOVNyj997FnQ
JXHoKCwDt8k3XzKH8AakpkhktXaeRKwhIKHRJMFWeNWuUC2jyK2rDqYCR8nCp4pN
+vSPB5TsGgbAUdyDizF915WZqj10Fb6ppwBljRXwFu5woCFij34EtP6fggRTwK/H
fBAruKgdzfN3AYketys5VRQB5TP3Rkn+srHYFwRErMIbF5YeANSseIy5oJbs6RSi
0JHSf8AIFQ5EmuaGF5aAtXRl1h5mjnCXpEohZpEnOWCzQMTNanMnUollGLnpwKyp
8+i9osVGNiUvoWSXCpVEvI4A+eu/aiZB7oOmDdvQoq94Ag1AJMZYzWHMmHocS5Rh
fwbku3FRdI3QGwaTIh8HV4KKihaq7zsz+XR17hzAkCf/AYX/56grNCxDMh2nIB8m
8Ljjw5SGu6Il0L7hRSfykMKKlGrOZ7qBwVYSAvMBBq5IZeyya9CG8LtnNJ/W5ot3
M/XK+U8xZjHgyLU2qCHtWvVm012f2x+C1AtLZlpRDYorpYt9y/XcP9k3lS+jh7an
aO2NhUCb4Cknj6bnfKZECN/I/hBCdrsslqfqshSOPefKYZ2/bjbVn8ApP172STka
9DgwMVLU7MB/7THm6+qdm6NODZHbX0Ab0jJP0gs7tnQfqo4dES+5bXFDobT5W0ww
weKAuv8J0fn57Fy0M03xaWwYRhD4oRf/tnCmxk0Ev4Y9Y0fjkOTtIEVVLU/otNPN
OoZpsc7B3Qt+GzjaA7XZbMIDubWqlRsAqaUkcF+uS1Uhls/mhQ44LOfXv3iiT6Z3
ExG3jH3sgahYsAKJGrcNzlYFVn9XXV3zlHPZ31Ql0jnkUF8A/jclaaJLIVDxKiC0
w3eSxNF1nCPKYUKC7HQILr/5+bvWR41jnf6mA6mzSdKrYQeXzfGoRabY6DmQwxIk
NWl1IlwsSOBomAj0rlp08VxrQcwB57ehi1JPIWeH8ncpTTeyX0uhL1Yk9eJVf7lC
X3JdsNMDKWerAAqA3OzdTnTWbudhD0VL7JYLdEJKsKwTZRX5aWM26h1XJKvzg9hd
0LEr8iuodOhKvX01ERkKclZ+YlSJHg275MiVzGLmU5vAVuwSIaCxKlalW516oRwT
MDgMGHlDiPJ+1wpidRpeLK2xGmEoGVoLWz2vieC8BpCLqC0muKvCN6vxv+3HKjHC
yWvh1RdOHKrFc7YPEvYJXlB/UxBFMjiRT0p9gtDApZa8bnF8exmyXPYVk8xJLnlT
GnU8huparkjrQ0K4LoqP7KyP+nu1X36ym2eiJi5Ye2Rd4bHs0FI7ZlyLS/SfYGZ0
YsMece7wBXT79Ll36kodvs7bmrQ948GEqktI9+kDSxZR1mD8K+qb2Hq1lc030CW9
dDfXyq155XLJ6BLwFCMN5iUba0zRPSyDkLi/Aw87JmTG7AcXJQGEcJ+mcPk9k4y/
4+YQjoyHdRgDqVxcPLdCmK1TnEbkWUbHtNzLMRo06uinIWzfEH9zELAFCq9QLp3M
RXvEdJ4HckIm1AgUvSqAFs3O4muPhTBJrH9O9WTCcicoK8A8saLwIqJAMPkK6tVS
ITnjnw+VknIL1cYHskDsK79w7He47sWJZ4UdM2PRM6Uezm3X2OX2e0omOPe5BT7r
85Ryukj7eY4RFK8WpWvAeifUtg2JebYnkqBCYgMeARHJ6lXmKYvmH4omG1ab5O0U
7Q3OZVXthhWQFqaco3ag2zYWv2wVImAHEe+4HaKH8qfn1nQMri8Z9TM2Snnf3Ng7
U6VssQ7NJOGeYzEZYlwMYIFi1UwWvpEgr6MQouuuDLsGu1x/H138YM6LvubeX1hr
3w7PnOittXLKD+Jh2OnmnutpdF7jrUp8rMlKEm4K5CSofz8SycLXH/TeP2OAMGfE
tJOEXbwT30iWxVRDuFF/6weK+fEpZpacdo8F84eiC43flXq4lBxR0syO4oLVbn9U
sPPzSvwP4ed1RiPJe/anK6bkuH9Zzg10CA9FeNRW6A9LlOCVmRwPR/X1MOLsi5It
BCAqJVNunIVuLLF/BlGzbHlUPyxTlrbp0MxeB9q4pInn+6LyyZeZRppVJep7Rc6S
nAcNx8dAcN9L4NvU5Wii9Q6W7AKQnYLXFCdHg4Ay7ovyVaZxAbE89Pb22mhQvuhU
AW68cu0ICJQ7k8mGAWZ0XD3BKcmmSYnmftvxTEguf6N1c46+T0wzdMfAE3b8IbHQ
MXpXVjXM+cX6EB288HkFMxSOGrPAMqIYlnpzy+QXlZQgeKnWGzupiq/hhLOz+l0P
YIY4BXAkCkGz0QwxKW3NgxW6p9L1djgOtPAbBACRFyG2asHnACPBwIile2AVOYZ9
xaZkRMl+tlmG92bS8o3962o+yKuAIiQv5res/FLeiTKm/G1yESPlI2HA6BPO7VZJ
7Qm0jNYmRz/vIjp1U+A7Onm4pfdK8Y3SqfUW/6lAZ+cjSezKAhJweuPu168iVdei
D+KR326ijkeY4xuTnnTiLP6g1ScBlnVYEhgqiXVVd+LqWkRDCaT5EeVMxrupd9Nl
pm0IV05qHBeCpfl/zDKI9+dhtEuqy3zfz2arxI7tT0cgXBTcX+dYRLpOz3DyMTJt
ubvh0GKzdLqHchwvcNSs19LJzYXft3vFLgsFgVS9gBWzBtM0glEYSq/MmUE56xym
Xjo9z66byzS7V8SkynhC35DWhVxkV2JMpqXMpnZlXuoSdTHnCqU1b/qyO5r5CRkI
TghEEEQ3F61zhF1n1Iyhd3Lco2B5wkLzbK9cab8qZGLqimmD2x3FJbNlZpnSaqt+
rz1ZeKyTOCdcBk3F8rlYXRsFCzt796sDbzP8sLHeQifIvVcomEPgTA612QGNgztp
aLO3rJn3hVII90xNCBaV8UUQlXhLone56RsWxM5+F1lIjsGd4d9pCpQTKu4AgE0S
uGeThkJJ7lr2TvDWp79VbnhnHtPlrn8qZGEUhkYVGhkrzbjqwjYHMXS7G2nN6hJv
Frp6Ffocy8cuyJFZ/5Y9hPhBjbPfNOOekRHuIFu/hlO8j6pCNsTJpZTMizWsCdQb
tRzcCPn40cIYRRCtuiZjHA5QkK058Vt/ftYT6VzEkNXt4B0ehuWQCIg1gPT/zVK3
3D02Ws+Q97jd1ssVrLQHgOhjaXUT9C+bKxInCDUUaBZM+tYe7LLgDBUvLVUxF9ez
3cn0ImSIGnVc4QTeAN+rx8gkabu9MBt784GExL6gMk+W5NGWTSuh0b7oyb7DCM0u
ZbuumxDEo88NcuMfdutjpQ6QWaBio7kWtt3iK6gCmz4PpNGtNut9jVWFMmLtueva
+dKKkmEU2EiQcjshjDPitoq0qcg6IpkGTbHyTZFmlkaFlYmLBtWhi65kHqGXCECt
xAyQKATRiM3Y13rH+CYXWa5+CkWt6hibSQ2p2h4Hzx9aTLDGshmiJ2TxSbkLpjGT
QqqEgD56eWFj/ziPfkgvdl244RFEnepCvTG7FyfclxwPDr3BvryWRMjEu/vIKCjx
xJtNm7l+iiemmWE5w5PnKSijjPTWaa/0kDYgthYXK+S7E35BvJoCuoTUk68xhWMQ
14cH/OlLW+ALPl7QATcqH098PpkOdzz23HxZ7GjOWT5O6XSy1pIP3MBd8lX5ftm7
Nyr+n+VLAxeU36ERv5Lo7xx0sUydEQE16zxPJn32RWxAsvrt5y+WzOIISA6g/pzP
8dboMinJoXdpInR9NJ4AeZldHfygIcISUr9pArhGdPcTh0NVpbLU3fLaprWLeEdQ
n8hKcTZRdeGy1ggOQJJBw6xEyY/Z0c1Hf7KNKpWOVR+gYLkPrUTio6+NXkSN8sy8
NmkxVEgic//TA2Tj8Yqq17TnOzON6y0Bbz9O+1kMvgEkab+s0H5vlDUutUXGivvp
1tlUyiy99MWABaU/yJXLSDxUzmtHt/QZeGwDYQxruUNZoDMMaJKRbB3977iqoDDq
IcY79zgxscAVpfcqz7NAO/HNd7CyUT+moV5z3nr3mkXmVRd5hHnRVQcXhKHEsitK
CF3AyMwOXfBnqKeZNuA6WqPyqfzEktRX3ClclgoXGaYjLc1YADpNHBYGF5D5vOwt
fA6e7IHwTPCVkmvSXrVGJj8kQP155gg3KMKfUOJbmca8xTboAyil5nadRYw4iBtb
5fBnQS9ekxjootv0K+392q5DOL0rFGFXSza36UQx3KP7ciDyj4LhbgtzvHzr1/c0
/V+MXyIsL8zUGTdlDzWBeVHcf76CCmyK62oGlVrSKGPI7q+RPst05Taxx+x7lfuF
7b5Fr2AQ4Agxanf780RoEpZTKYI1aMqWKv5cc8L5xkj5ej/yjW+iO2nAEI+glbbn
Ok8MKytLcX4qEcvI0Fs4K0g04T80KxGjK0UcWQuXCQE2ox7T6aFZCb21VM74sZLI
sWdrjb0LHYZfO9lk24Ai0sAA5RDHgW8LBh3qQFU0XLyFYL90WMsG8k4KTGupjy50
046T5kkZqVLc209Ornsps3A7V2/OqMtCCA3/CtJw8le34mRfUIzbjiTEqiPMN73O
CJcKjXmmcEeRwpgIcDfiqa7PkulK8TmwG15faKkxyz+zLOeNvq7ACo8FsxyV1zoY
Vjh8NjJ8SD+14WYJiqudDNXaZ3sgP5nf1eP0a9XA+k+jWwKVWCfwaN9R72CEjfSX
5jeH5fTJgejR70ALkWmM2U9PQ8JagFgdPE3Ydy6z1OzgD3wDfw7UhoSov95oSNgk
+9Bm5MT48+n8cnGF5ZRm+p1era64VS0tdGg11fYqOiOZuhoCnGmBEYViicgTRP9/
jUhDvOK58kcKi1syTnK6FJpn3n/XniAUyaf+Ya7BUdNTfEzIr6JMYlEO971mtSoZ
ANnqFniy/Ql+h34oTOG2zPW1jQKBKKVHT+jtGrdjIAWHCqm5KAAA7g67/iaWdz0V
+PC2H3AliGTR7IU8Jcx+RB+6/xLOFxYjkXyLxjgQ03msvDyvB+Wblcmq7bDzKClD
93VMXiuw4ruhmTQrBZ0mqokusjBC2cztv3HrteO+Gz8FU8/RcB4URnKw5dH9AwUp
BB629ZG8OmbwFw4Lbp49BYhxd8UPthEAsWtEuP6S7njvTYn8StRnLgSxzl6BFB0r
+P+d2UTVbzDMtrQQ/UMTAF+4EfMAjd7ST6C3tTFucyroM10H4R8ZFNxrffVPaqLQ
KhPCvgXZfdJKI9gPWaan6an7rQF35AYropHWlrrfw6FRA1Rv19fnDdUFd893ZAS5
ieVyc9sLwoKPTTA46mt0oY49+JRXbdd0xuhCDR9tC29r95BSH1GjNp9YYQlc3Br4
4g4gfl8Li06LMCAfapdprLGwDFij3G+v8+/GpBSLiW2ZdVv0zx8ZlIR+Ay+9+Ycz
cc90SVnIKTb6u0vVcYTJz6z0ylGo10qN6en+kSWGv0FzhLAMaGCQyp0Jfk48y+Zm
8VMLHWf8Q+p4X3wQyRdgT6uzWCLqIoT/qxhhKlKBhQnLsa1sleIpH2L0MExbge3z
z9gjAr9V98gl7rxcZCacADPKZcNUj7S/8DsT6ZuaQhzlYikoiwxDFx7WzIvdA+Vp
kfiU+TvHaQ/O562POmRcDHxNMA/fVXucPmcdmBbsrjJ/qa9bt9NCN3kDZDBdpn8q
O5Uj1RZzGFwFDtvNdeuWQN7QiA3ydaZTJ9dmg7OIUFfBAkxlkxnZptELPlOJGdFb
BM+Slk+AruKCFzuEzXQiRjI+l24txDYOt4P5jNsBpcRGJWBkQ/Oo0gxvB5M4pwBT
nXiSTImt0d/NftmQv36fSdWxtXQhU+2NMq3xFe/F29cwruHb09YnI3u395mghFFo
+jSx30jlSuDr/U8vPef5ps6v4kgrcih0v9/oaeB/gAeEMix6Rgw6SKIBqkY4WJyI
DpX6EwXgLTBTSNjivNyC75oUJsAh0tBz6lFPmaM2IeE96f18IAVnARXm7/7ctyj1
cVDLqf3wwa1Dmymn/anFm+YmtphinZbvlYu5poFtJCoR6MlJLRdWlV0c4+vhXuOV
R2ScBInptxKtHk8z7rjQIjyE6mquBZH+2dagDaq8R2Gl5OWBmhPgkUObx/CzwzuF
RFgBLB1RBSvQxye5PltoEWaNyopWT9Bg0bOli0aZ8GYjFPsa4vSxsqBgul54uNGT
ZeEE4KhVSMJglU+h3UqX7O2osTckEX539KK1bCSU0Ck7BBh7RJKE+lxxGX+SjAE3
jrfOC68QKa89y/w75ODMBe9JeeN1t3BwIQHkQUMlqJHUj2XNpa5IDIn8S/bfu8KT
6vfzvKiV1RTD5mjE2672wY1cO3cNQFGeDnSLLpF5Iv37svL++a9P4bany9Gbh4v4
JYClk6upQSxbR6bcaMafphXgAnIfw5xbTbXotW68jqHbdU1TH1SdbuhkzLncvWY5
QYAIhHSqJ3FAgKrG0DNJmOLl2RUdL0oyoRvDWZmv2Ep5NiBffvBP2upqwhtENEfP
lt/Lg1B+IOGzNVKOtbabaRBGf0KZgMwGtJ7FqPmlhonC4UfEu3DZ4J5FRMnO7g2V
u5EaLedloovhIUB+JRckIH5i6s/T9kR/StLWHF/uV3gMeNo8yKJ7TXYVQkSZUqES
4eP0mbESwPSVbCQF4RiT4REkrZxMSQuOcYrzx0AwxmFY198t7s72WUbYxwd6rZO7
crbKf0EEOBonxKsJ/azPN6DeoSmMooLM6aYrIj8px00+7l5vzU/ye4roCEq3ZJcN
rKY4ZsmUCmSHjyF5qbJxzMXzckpf5dgv5O+oe2l8tp8ZlSwYKJsOmvuN4nCpLble
OmEMFK8r8Gr+Zdc5VL+4+KQz7q277nFHoEw2yIGJSNWFM+3MSf3iwSGlRgpGmBjf
dOD67Zpbr/cIxwuqhZhdwA2tbfls7gFmK31PLIk+9TcXkRPxhX3Ocn1O2RrvQlFa
qXFtqAcq+klR+MQBx5KSHEzJORXV0aZCFpTK9E6g+ddaa9d9WGcJmtIyMIX+fqjy
ebm0EZ5+tBm/CnRKldwusPEOyIuJB/sxP5/X7E9aQ29oGquL+nBP2i24bRwKF3yf
O+NHJFa0d5j7vU+6XptzyOtQPMXnUwfmetKJB5X6NoiJ/CjSpimcF2F4jz/iY33D
fLFuLXS59tead0j6sQ+3T/eAXabV4LYnKv74l7uMr/4bx+6vENebUdLJDnBT4yqo
y9yMw8tuFjp69p+vhZRvEvekTpZezlQWx8mqGZDl/hcm5LGlvCKwzP5qrtjj/MM0
n54T/04etobFbf/9qsIeD4I2qRXHghZ0srtss67peLSm8JvVnGNVPqZ1zTfk40nG
PSydvhn5bto27ntxgRManVUZmGi3H89XuJ1jZdop5sM8kCuN6aE1/sjn2V0RK0QM
blaG1WL/b+Q8pNTwNhWIHVjEbkdFm53UCkzFdzqigOV16dquq3zb6cgfpZnMq6Kf
JTJlSlsnRfmnTzevbbWSD+iHaSHgyfRstvo+5Vvc0K3HpzTHsHP575js2sD1wOX1
SFrSxpf7ZXgezOgbcQb+6NGSSdrK5E1yAfzwm47CMcVfQKdQBmZFUH/Dvz1MWyDL
AdAjtGLqQAVTcw7e5vJOzvXgxFYmQ33cR1UBCSDQX0zlz/tM5XAUADrb9qWVXeZX
gLzwDik0J3k/9yWrAnVqNB/gLDywsdjUCYnFeHB4Sk4e+/MEkEb+mJMdjVAZ+fHU
XnjU802vMjCOcaRdvMXGcJRUfzAoTz+qqa6nVKBmltK20n+tzpQ9vosqX5qDGZav
MEUQ77ILzvo5JfTXClMuQGA2DJ0seUl/NyGsbAmvzkF3/N8lz8iZ7Ea/BL5MK/DV
SMo/Uhpt4G9t0TNqGpU+lb7hdxHIwpHiS12jDg4nCQkA3068VxnqQOhth+H4YwL0
8TvfxABSt6tNd2KQR1LtodDqSqJtYDPYC4nX5BFQdaO9edror6IcjVWtdipn1G/P
qtXlLsTLRhWozqk53mODXgCFq316URwfS/sH0Dk1wmzzZDyiIRdsCElcXBN45YXx
e0zDcGCqNtYtxGCwbOvxrr42NF9U2i66R2Pdx+QZlWMq+YLBZ+mVbgmLeLXz8cu/
+5epKrmMDSIzW5OnEYXRhSMdzphyp6zRtoWmVWGzWyGjeZ3E/OcZ4u0wJP34+3P4
vxDE/joQ/R7W77a/PBR1olhTMLGbZwx6h6Yy2QNPed+okPfOvFZOXIEjeoGZ+fqh
+pYiOh9/eu6/P+dDZwKtN7Y9RrXjG0u12KxPJ3rDYgg3RvkE94UDpwCIJzfOuLsH
2EGnuBagAwGBYTvm5Jjkex3IZ8wvVGgjO9EojYTASooCfkwwy7r88IAfRwhf+kqY
9Kp+jzrFTmUFwqmRETw+juVr5KvrXaGEHsXuNkgyWiKC0GYDKdYgJSivA2EB04lK
aqbnhGKtimatvHVjZpW3tQkzzxWKly3b2BmlLUkaIPhsAUjkcyX9AEO2AbDKpC+E
h20Ug+PsanDre61y+a9BfLtITSSGjAJ2ofhHEmYeztoGFocVrUeDQwNUdgUd0sHb
wPxJhjstK1L1apNa8TWcblLfspOXoQf+Eb/U4omEI7T87qxg4goPB5SeFFkdxESv
lLEs4hF0ptWmReVe5d9fUmbrlGGr6pBYWThmGDZ+Tq6Qzz3tb/Swoh0gvveWH5uh
mLQHnf2fN1ZM/qDOnGXTCYO7kOhwQ7UKRfm/0UW1OLUx0OK65LHOA0QCUQuWGryu
DyRZhcKiaLCmRfbQYeC7Yt+eNdubLnxZanwuK6PnN/xy+XpFkjgCnd8PnorJ9vee
9Z5HgntK783AUj1AL0rp3fPwiKA/bc7Fne2u8zdanOZxXqDALtg8G57Lv5hdgLil
9DVr2GjFgVajVasPkSUDq4WrcbuV5PhKb3np59LJ7sXA4+LWZCSEO3pgme4D/Rvl
Vm+/YQEipqJT5PpthIW6nAkrDkzl9hsX+dw/d4aKg2mjLT/m1X7QAHkuwpPUPwuP
8aAZ0+KNhCPOQJ5BopBCYb1RTASuV3/qdBJrDOmDIZMrVoEJbfTtPbYEkzyKNt6a
fAZv5ztiY1wRAGWpGUaSb294Ml8O1CwQKArMKT/BFqznIWqYTvwZEW5oVoWpLfNw
dUUVTKSZDzh864XheuNjOTq4opmEESQHzIa0+TqrBHWzm/ISkSiGLcinZaCt58JH
8r+72eVSPNpU7flyIb6wQAyirCOc79InuYqOO4AZ4pbSWoWSpXbSvcDawCFl4F0j
vrD582zTx7cX/B2J9jSTUoS/OqfiuIw6gvzXi6mSyir0I4Zmb6Cy1SNG8M/OQQKO
1isJmIEm7a0aUq27AHBGXlKicLuN8GmoCweLbCLBdkJwfyXhhc9HEOI+o4KQqIe/
ko+RNWTyKEbt5sN96syJ7x37Dsu3VvFvRHpqMjLNhYSPYcgvr2J7nfq3IN3i5/gX
t+SlmepnOe7ihiq4jKgFQHO+7GwtFyzdZxzuEvmPfXqx2bsEePd9XLH3ERJjzWNN
tmRp3RtPtESdBf5tH60iV23zryUfPS1xWS68TJKhzPKWRXxNVa6ivFvhmV0ul/JK
ekCy/gpQ9Ah22wl90JFQbnAI9FgZS+68vMVFol6Hu390NNGz8JZ/WaBg4NSvE1Sk
LE+9KcJYKI5lig2cqvB9u2GCK+UW61qend6mFnTmglqhPVMOMw5cTGXWFBkaKjGM
sogqcG+L7CIFGDqUBQEX/aofgPPHPxl6pRxmjvYSfoFHHXnF3Ud0vF5P96b80GY9
6cfmOytimLyMfq3iFhzQRxY/VtljnRo5+tcvF4JejEx987hzs6bAzeMeLClOhaCJ
Vil7EK2ULb7IIscYP0fyCI0QZhQevldk5flnwaW11a5oVk9qf8AZ+DAj2bG0UF6b
RGUg/dhPVu7QAHKG42UO0aYr+79Nm1etYPonkTn3PxgY9ypA6zR8KV0ftwWgmDI7
huIRsx0UiYLC4VYHcWbEDVUhFytCdLJ81ZDVCt9vXNO7I7buVSetBfs5i0dg+O58
B/yIDMMQeCi1xE/2nmgTui6p8Lo+ggPoQ2URPZ6JeK+ha1seZWtLznMy2z/lP5gL
dN59zairPMHqbkiMCZFhYdoZP9n+kjpN+LN96OaVLJgcUU4Nowc/mRMjJgbWqVsu
eDAUeBcAryOgZ0BQ9Qpun2F8XdpDkrF27BsNen4RQsp//wR9ClBCZVNg2Z39euWF
8gbsW2sFejYQ9OLXfk9UCIZl/2pAxOH6bqEmj1Vemjgte5mOjntVzWP4Q6oEQx7X
fGDG86iIDXZ5SUA2YZNAJ+GpB2Ocfo1Pfa3xH/h7/+mUor7ZitLGIPwXkdfILDHe
7aVYpj6WfMH9BMXCyhV2UT+oadlfnTEH/QNvycBl7E0N7XtjP/ZZKZWI8W6RyJiT
Syc+qOlQPdLpqcSXlqdqQGMUfyrxtBA/82hT/Bj3/Es6Ju3zbGXX8ySO8XHj708C
UGC/UBFM2Q3Mgl4xVuJ17WttQOAjlUbxg2ZApAQknjnXnu8JnCUnPXR2xzV/bIL/
mA6J3SiUMKzmmWBwmJ1XLNhlcnZmINcLelfsPwsKSLkwoBNt/qurpwN1xADt+hY5
2xzrb4GLr4v1t5JBopcjx0GtDv09S43PYiVWzsZnqzzIo/frMN9c2wo6IbbATpp6
/a5pMinVJ5dKp3km1KuL8+cZY6cEiCvBU1wFTWp4E4MCQSAB28oFAdg4jKXhNnW9
ZcjIiMnQE2QFRyPpThsrk6AR2BcdwPDQLXuvkj/kwYI5ReLc6OAgvENR2EMzFA9s
kD/8xkrI3HhVcnNdpj6y2K756UhjtMP58XHGGpr3yZ48La5DzAknCj3h0KBd4mTJ
u0WLCUtAVlETlNF/OM1WaVRWuP+A2yGTLawyhLORCjre5pCnYK9DlSpkkXfAkm7A
KlRIrVGoGyCSjn9b0OuAS+yO+QnQ4H9IA/HaW3vfCbsMCIHo7O4hTusgdp/U6ByB
YARqy2c7n7OdCEMZw5dF1a5mnJqi/s+st5g9lmLHXQc84YUfrwLpMovqmqU6X2P/
d5NU6uVmiesZqrQst1NCRts8QpP+F7ld0p1vnpGhV7dCHwg5xDTRSRx14cB2HV1g
Geue8pp4DkwQ1zrRVKjz7Tfl79LJQE6+4ZCgOz2cZa/AG5g1aUjQbap1CEi6q169
gejBLGpNz+LvZP4qIvffNA7n+5qbxH0WK5VKct7/1mF+Vj1+gRgW5H8Tpq7VpVh5
Y2Bl/7/8snLYuFw33esaYE/1OTAhI4fxQQi7wEmDJGfDL1rMW8DnNXYHkqEZhLOg
9WENIe+4e7SRxJ2uz+woodI9ulnSmsRppVTjD3o9jYpX971v8SCHsYoY6LmxI/fe
9KbfA3ojT6vJ8eupUjyh4f+bMzrmEc/OX6gru58/dalUJ92Kh5VaQi6e8rtarecK
M52lX9b5mvQ+Gqxp5go46HmeVG8ZFqheCwdelY0PorbPvtfS6EnZPvdNhXMfkn5q
qNKM4fUWCFItzD1DvL2ruN5OkVrMACCqw4FiSi5oBGcChgXIHHDbP26aK+qqrZK/
aczu5cPh4efg5cX1kZO62ZQLx1ZCJxuDzwjOj8829AEYUKZkn+CxK5wZQlkG0zY8
t5lafcYOI4qo+ULF9GYGnDW04a/Y0d6ECprHrJzd1WZbQwV2WHVaKJc1pu/eVAei
0HwGz7/fxGM6qDvZSy6ovV+JC3KmJo5Qut2LyagiDKQJy/Zw4IPB/Chc+I3s8pHA
nsG9PkGIA8oRgH/tCaRXSNekjyUbj9gx7K43d7flvAd0oTKhLRJZ5goLOE/SUl9E
2ZO944H6uUof68yJv9VXnrWgXegjqCflDV59ybIHOLJWCj5pVKHsLV5QmVrEAFEu
+LMCBzD7r91aVBuBLaSoH8xsxjD+zmh/6hMckwqQAd3Wsv/SohcyM+p69348bVsP
Ixe4u+egX7fYIIsaKgJqUmU1/8uaRzLarGYwMXSEMHrGqJ99yLVhj2D4mBAL7OLb
+x4B5yMRzhpBQkz4A0NB7It1kvRyr2JaXoLsDYjYmBVsyTeCJpL6zJ44QHxbFxgs
K9Qf+uKFEAYRmeSmqOJMVyr3b87vCuA+96jSS1A8m570jRKdXg2evF6Y/OdT725u
yBaM5IkTIODrGcnPjZzzW7FUhymLBzVAcwcMt2dU3sP2DHhaFa3mtP5bDBdrzUY3
BpqfGX093qYuDYzWnbC44q0LXKnWNGdrQAPI+KAc8EFVUtrwooqeWUpom4SMewjp
v0koYp6dWDqdmHnjSxN+0/3zD5UjdFcNIDQ6QaT5sXE08cPMX5hMf3lDhAd4nTuw
HJSBNmUqDs1joXwu3nSfzhFJ2qyKDiDz6cEHTUF9wl3xT3KVGMNW5mVK3GE1Q1Oz
sGFYLwSDOts44nuhRg0Kt3pH1B0Fg2HOF1EEh95aNdCvVPMpyfFo8mI3mVD/4GjZ
7tBR1+9mBPslBrfyA5EBvPhhbDdv4q74ZMBb52sSr953MT+ljB+wKbDBE9USqIzH
xT2yC5xCsodioEpyrbvc+88xnPLsMlyY4Pjm69muOaslmntzWhHs/Owjz3CEYFQl
Kr5VSA4Vu/Hi6o0Uk3rl54+9iSxnmfZX6VUqpngvPfH9yLWATpVZpq67bsmUa910
kML+qDpb+lfQPjH8i0lyjG5xWOvAACrM2SfMtPMGTxWZliqqXTDtwWvxbbfz1bo4
j/ElWppnkRmQvXSEfbiHlQUhPIJ9i8ywRFy9WGZKXWim2zv1hpf/u4CnYhnfc0s/
iObihCBI+DlLmD+Y7lRgwTGLCSor5yAOKy19LYu12ApbX5GyF/Pm/e4NXzgQU4uh
MxENspj16eKl4USytvegKfowApHDE6sPohPLk3RHD4jXC/pGROgxV6sxY7mdgf/n
PFXeUcRfOAyMhxIZE2Hk4SuGR/T5jgCVTzVYYCHe4MA9QnF/g1Qc9ZwS/72SXXXv
3+95ZQR2XOgR9JW5NiXiYtjXbL3NJNdLjNbr7wGND62nKn35f5PMSehHcquiIBJw
tGd19Uio8yLK+ImteZp5PgWRgBMwEkU6QWyBz+9RtEOVEzcc0QiwDVFEm+fHRc2E
Yy/EEz9wj8RHHhuZ1b989nb4zl9bEWL6xfFzxUneEgjinbE4KMnbGHF0Dxq5xb34
k/5XHHgd88On9Ubeuoq/+g05C77nddxgnpY1Q7GPEpqws3yTwe06WlazXL/0Zkox
C2hQt/4TQ9LXrulMRinizrGumBJQTzQ8xw3zE62sBMGg/pUgOou5fdsqF+Amr3DG
qws5zCfwd1jcRPP/TP11lOy4HcYIBEyQKKxCFDydOAeQ8LKA8KAvi87AKD3LRw1h
EMhB7lX0tVXbFdP19KdeUVvjV+JO48GquixlI+diB1njvQtOn1euE/gb1h6/vOvI
o5dOtP548bMtdPwz2r3KBf7ceRoAGu6W1ktUdeBIDTebs3e70mw0nkkOVDMYbENA
y547v/Z9SZXn6BEceLNcrOO71uoc06HnshSW9MYKoPYxuAv6CVxD2twyYPusvZTM
pCKEo3rhBahiTZ6QD1mI+JMFT6OG7NNUHXq9P1yXBeoE3itSO46Rq7W+35iesR+h
eU8qfxwdNfCsuC2ur0WTQSN22VvpGJ3QDVDxNJ7jz+Q+BtpVwFViIDqeIKlLHX4e
8//gfE2M+1CnHNHCt32EvIEtwa4daDawKjBtV9Yezcugf4LFV87WHo6uTKXiWpWj
9NFWpHSztd4dMDMtZBPkjXpU4efauDHT3bsQTAMcl9wbIuyGG8/xMtoYexMWWXaI
xOmvS5/d/vIaL+MwYHmKSUSQvmTxZCfgtD28ibVIlQSD9EXSoIFy5AVWT32eES7n
dHciC7onSJpr/RgPA4e2lqzP6pVgWABrCilfFiT1i+CFAOO+dYvUfRHAl1s0rlgA
tW8b97ms8/9MBcQgFOze5lPGFlcXvQ+N9YZsRXFzhl5xwWlNmJyWFw/wnG4OPi4s
Wzf+k8UQL8Wm1qHU7kH7DVvId3DSddK4qIvjsPhjnGHw4KJQQOlwUsYRoXNTZl8b
K+Iv1fadNmOe729vRuG/kB+MefVtMuBK6YF+c5tHijJL/9dMd6bbjPCf3exHT+nI
KvqfSd/rB4rx+QZxU0sYXeM/SGYs6yDDMKaWxEAkzsPb9uNTS0cbpcryWYpHTrOq
JkG0dxYKCd1ATQV5QYO+jTeOqT9JPBw0Vdn+ivxGWBMy6WeVQ10ysDqOlwt0r4RP
GBZuFiMZstQVda6oC7bPh/ygMS49cgnsq9xSc6OndcGE7x66eTz2bYpsGIZIbwz/
W2IZmIuoiUdl0m74tk/wUqbfsCaAVfS7qtNgf1Uo17+Y7qwtGQ6YBa6CyPGw72KK
MubXrpzWiW1uYvvLjh0znrlIpJPs5Sk36unu9JJOcAyGT0c/q7zgUs207p5X36oX
fATtduMNH2WHKITnEYuf2YUxoAiR6OxPdyIyw6lcN0RoKmIhuG67dpRxZlbFxeO1
9+DmuDLPTQlLADqpazWl0a16PhKCUI9ZbiOHV2Av+IcH3raBQ4EQQQas6oQPKjDV
nkAMblY8d7waQOH+PW1QBF7tWIXAg0+rzEMKc2uYDdS+CUTs/+2A9zLCxnVaBlYm
2iMRSL3RDffA22dWNPcSuuVSFyfuqa8842FX3xEssb8cWHsd+bShD6Godi+ss18F
Pzf+ltNg92tAvFEewn5wB9pPPWIwwhJaPFFcalWvKv2YaxhBwxceqXOKbvhJEoIR
l07/ZtHXx/nnICPAHVjuE8eq4JiKsqLGlM4i8y8dodCyeRfZTar21HSqViJJ/X3X
8KooQEX1SFvYkxcUfNT24lb/XdgGR3cbXsyKgy5bAfXFPDb9rdV7EpkRYb19a7gw
gZ/2aMlq51GFKUqT/hjn3wE6EUcyr65q72VXeb5i5KILeW+9+6L3hS/4USRZbKL0
31UccMENdXldjYOgGYv7Kz3+Ep9bCZEd33dQR8K8XZ12S6ZpBERlqllVbZ7eyf2b
qM+ohA++5XyDNtyw38TCWWUNsL0YjfRGk+cLLKG/DUBEqclfHO+JeARbh4/FBr7V
PelgLKlug1PSlDnNrqkHAxY20Eyb/X2Oi1Yhh5Vb+GqhXnSf43nuTMDpq1duzWYn
qFWnjKiIVJ/8BD2HZfcle5oavJLThMYvPA321AGAqQOBKdm7fzHLeB5It14hTktw
Q2Z1r6j4VABWPk6X/PS7D1r9UFvmwoSNRgc8854pWe1RKUpmIwxcE+qGgEkGCHhA
1tJ1SW75ubSFScItlLhdihAdsZ8tHscNHIsIQNBixIxqqQAEaVZCJ3LpYxRKoHnq
p9/Ol5T+KX5X29rSLzXJmBG/hpj6cPtzOe8rwiCGEiZIIDjgzAFZaFWhkQC8ZzDM
NQX7PEjzMFF3Zj8X1+ucb8aCtBXvZNrIJ7a66YZLNXwfL3XLJ9wur084uOlgDvkf
kQ96sxJ+PFIj6dNzMjOgpsuQoYRS8DWrxzwOixkl+HFDihuL/wEaNHQ4bBvKQu/B
9qe9bDQUuMOsHIW0orkRYEEHX1swCKpHXKYIxDventoq/RHebJRF0+BK7EubzLjB
VXDLH4Ly3Skmz939hrxERP5jFviSm7epKxOTqMgVcdr86YUyFrMFSKYIrTqmD6IE
3jK/uazRF8dckNWcf1q+YAfpS6nUR8NQMBUuT35W5/ohpJ+pB7SL2oWmnTx7rhdM
7b7AoHlTeEEuRkUiCOiR53tZNL1/FAuTz5490mFGS+V3q6t0LOo6BvwySIrksAZc
IWfv9GRT6ddNEKdg/oV2JRqng/guDMpRxa4nNFya7kb1pBz0UxVn0wAS48SveMzc
9ro937In93SEozofGvpAAz0irgvSEGPAcQ1Q2M5ZBc08RFsuIFVTPJPRFa5VhZKa
2sjFrLAYLQDFE0WQbgbliPXIZmmcie8HlXcFgmGITss5/Ic8zTM0LY97iXpVmckv
IDpAh/fvX2pMRvQYZXKG2RF/10UZyCIlfzNDn8cp+l9T9SNnEx1SgQDMUV1/L94V
Sy1p0OKc9n0/WdNFm7iuyDwDe8AAkbF1p/tJQY832R7kmBG96K4oa4bk20BwDZQg
6iwaghTIMJPS562hEgYmhhY2qk1z6Imphqn+sNzc9MQ+IjE/0me2ZP9ZW90Mpc1L
fz4UcqDS5cr+d3reA0Cw9BNTJECQ7gPZn9dAYb70htZp0M1kaksU7YIWl+80nax5
Os0NosxIJz11o3GUknjoeotxJWG87KRu2c6MmnUt3mGn+KwqNbeSfoVY3/JDLMXM
vVvMJ17MAfSEm00gIJ85sDJ3m+13UR1vedTDvheDuGwqTQUgQxRGB7L8K4IPU4DH
8JK5f4K711ReN5FxHnTw6yz6lNkNJsmYRiYdp85yEaGIydMJGc390Kd7jT7vxotO
DGZHAK0ez0/TXWIFQSSbYcOJXBl1B8tDyuWB4OnpCu11eSXcg0mPOKmnGSR5E5O3
f6ouslOg2ZcCuSwCXMtLO3nQDb+2ZZ7XNGIjD5qT5UcR01D/15tPt2dF0OBHWAk0
oQt/M109ToPmd6dPYsXqGfPU2b26DvGZe8iBkSiFAKzDZyz1bTQuNT2AxYJ8MGJq
Bhf+dwtzEGgzsGNZR053tmJcii14MzhMNgzZGltPWbNNs0rmBSrE2QYnBl8L0jOm
my/N42Z1BE2Pjg+lW+N0BTvJaMG5lTmjYtNbTvtJ1eEgJIGUfabyIaFL7Pin1cac
aplRixCZB0ZCZNj0PKvIjYQPU7VY3AAfiAGox2ZEoRYH/a8kj2izS+YWT+NZPEDt
Fjk+jSjDpjRXtnZszqkQFiPEF1ZM72UoxS9wxFs1vAaPfKdRxrWICM2aLVMHZPdT
XgTt/btDu3nmMQReqm0epfggEHcDqGI2Ao+S+crjN8WWAWUdqxxZtiszI3le8tJw
etytHwak5Nvlig6qgdWXJ3kw/V6YGyA18iANtr3fbxNqjzaiUEhA5Ej7Dc8EaYFC
NqCstUDowKhBRBW4lo/lFTLJkkWiHfC6lkoNLlf3ntlv9XBDws4DPOLAu2W61b1K
r/01tLuEbxE81+VhJvHC37SiXrqYvlYQfd1bOrzjffI9PZcZ7p0Q6payngUacpx+
1kEhOzdWPCjWaPIW3ZtgoDKgRL9EUcSj53WXgMtIL8shtqEewM9zQsMxivu1iit8
FGBOqDUVYSHqXf75w8Hx7HH8KLtVGVD3wcEiJCGmA3ygxSp0MhQ7f8JolGu6l83x
xXN06Aq8nZpqWCA6jKwD1a92WZXf4Y8cxqCCEDKnbVETSuy44zMOhRsLzRSL8JjX
UsPJGvJcoLFmSsgyeKw4Zu3yKzHP5PrVK63Dx1OOVUd3GKhdf4YCvCrppP8nyGws
8jP3liafYNMYgLEDMqcHnK2vgAql9nfk5p4q3+rXZkAeMEyjRWI+B4Uegs+IeTdN
Q7I7JF3xVm4kNrDnsYepRpoc2PpGENN9b9Avq61PA8X2oNF1B1rrdkJQu/abWVBp
IBnkD/HnjzK7cvrF9oL8II89FR17LUC3lIEqlCsWKkowaKy+TCXAx2S7WskTyje6
bqmtk7KZh0hsqBBsYiJUNhJgYrgyy85scbCDIiKge0StGE18JXlTGXsXt1FvWK5W
VdDypqksYgARy2dcNcOyXVHDpVH/Ti080GwQp0i7UXZtS574YisFchF+ABh+9FOj
GBZn5ncR5Zgvh05e/RT0a62KpQD8Rw96OSizuR7s+b1/j056B2zgAYE+lt0MVQqv
utc2fjg0y3BMT9JnGgKhBnoY3XUct41kEKQb64GgM/ATwWFaDpOtr1fkuo0ZO4bH
yBRZc5kDE0xmf0zmG+BRNfSZCBBoqQklNPudsl6SO2vn+3E9/R+YbSTp9E0gZ9B0
x0ZpNlrF4+QzaMRCdowp1+Qwq6bnyxp3ZZnxCDaSVvblJSGihCbxQyWpjxIYDDcR
ldr1UipnHH8Loo7EMjxuk7Y5x6ET5RAF8ryvLzcZbTjx728Njvd5Ityd1v2fTdb7
lBt1jBya1j65KSSYCJDg85g/QNGfqYkZge/Td5z6svXWmoiH7AGESC8FX8+GM1a6
3kw5L1FxPVyFfQbzPtVGluDYFJzur4dU4dBzdP1FbdqEmQek0EPTpWMNKjNW41J3
cNWV32+OX/gQ43XOqH7vdO8rtirvDQcuaWIR9F4d9yKpuMXutaobQ1HsGxjPgMZZ
ezFHrJsRcEUmwdwIhZBUMylbnFWub0ay4TxCB+h5nAMWmqcijyTpaKKDh2PIMGRT
okvB8+oWPne8NOiYkRkep7qkMtXPf1m8vLfVXc9ZFAKwdbZMxTSv0keajgj5NaNu
8gdv5qUU4oX9LxCzL0UahkC1+o4/MLPQfeRoCi8PDa772wYUwh1/ldR1GZAg2s/V
eD7jGSdasz89/a7yumRhicdwoavV9PerCJE8wrM5liszOTH++EktPGBeFEVdL1Xz
CIXQVGFGQ8mF54jdRXmroZ1DnUYSqw6qulqScnJnDJOnvQiwyFs4bOt9lZu42lTe
4dCCH8iAFGWwOkqGoKGwr3KZRmR3kSer1cSinBi0RpTpFhxfj6FedqQjIH3q7KDe
JBYqlylGqzzc3Vcu4ca1ggsVqx4wvDYaPseQc/H7wRNk26LeRO5CUQC2qQXo7eXh
zvYU6HVrlW/H8KE82jEkoHsauFuyk+JasgD2IjyoUEHQD44D9jnD86JzwXmD8nn1
/X+cgvQIAs8qHF3FpznZp6PRhNmTWoqUA/TDnJebq+DvNN23ftbbXza57XRbQ05c
m4HW5qW6rcAulc3yBfx36T3UCKtvot43laC1UOauVtV8nr0gsTIA1J6K7aSAbwti
00nT2i0qCLbnCtLAKxXOcLoGTzxI0da9LKYVwXEtc6Bo+Mht18Qi9Xv50Iv1c/nU
pGKBCjoKlUl9PPtvBpEvNwU08cg/4j4m0FfBn2Zm+x4lgpg8kmNwaKOXu7OgawVw
CFDtHWK+eXa2T1/qpLjQN2RPdjM95JsWx/WFbNTaQeyYJn/AuuXtQdITiv5+Q6/f
mklOa5f1MuVG6VSwvbna6apdn9CsrvqHzjlOS6xge59zIEsS6Tj9I8d+VP6cClMt
MWbG5R6BaDMG7b+PabSVuZ651b5W6ATGA4f09oXE5ZHBu4IXaqDrlFwOO5sN49nW
3IL1U/FMXKRLCNyN8cw/Zed/5vBPANmOGgx26mFOCHNjtviA2iC9por/8AlO0Lla
dObuZ9JL71ghCGDlVPqWc26m4B5MjLO5bmx1GKSjZIEdaSn9/UWmc4QfehXA6ZWN
4r7lbaTHNaGN5bCpRpJ1g98BeI5fkAXz/ti0te+tixbJ6DEfsGLKet+wq4Ha13Et
kdE8w/PUpkBJPNRFYWc6y804Ck/2YgUMoaM2wxcmfVv94geOd9I3g5FpKbONB7DK
Nqe5HucKwR1Cb9EkP8ag3R5ZUsmcPYCVIRVjs1J+HnqWTohYguqX1nrRw9nnkMhR
pbkmNl8IpA316B4AyNematO3YcyPO1JJPLHDVSIOB0UobPaWlIp+BBoCCnnJeI00
2xRZaN6nlO/0/c6I6dzbdm1tpof+73nBRq+4GFeYzJT7i7KQKwZC9WDi6UqHGkq8
Qd4EXCZG+IbRijEaofZviZ+qZ8Tf2+wadMwQxl2m5yzVsANHrl8soC9tWxgoeuR+
EAdQwmobxXtt9yXh2fPztmSI2c84u4UFFONYc9CuhxgarFbR2oxDXL5CXQU4C4MZ
YlUliZ6QSNt7RPonjFmh5WZoIKpFcQq1TXPg3WJk3DmjSVdWj1bIEMFq/5zmeTNo
mMGQuyW8gL+eojRR00Q4BlblfGH75jdWev9/5qOrgvlnnnXh4Ia8uk/d8cRgUl2Q
Df3I7vXd2oewB0Q6lWrRG4llnRwMvqh8LPJUyd9CHur1FyJSoO0EMz2HrmBxbahn
Ss+m4DWCbnbsUqeI4luz0dEJU7/XUd/ulNS48tX+Qp8lP8vGjg0T81H8ofkf0vLK
IP0sz3T5thxx3qvFnwH4YOaTBJFDvO3qvDr3b61p/4ZfRAtBy4vGJ5QuPwKnOua5
Q+d6AirYIfsk6prMDLJmK1tAg8sEKEYC9xqOCTRTFYxfRS6qiZPqgfBZ/+r9AfJz
cmLWEWK1Xj0LNe5jx2V7bTAVorV+/SZf7UG0JjUaggCc5QnDbaO7IYYKoKDKPr1h
eD7spas6J+XX+ZAde40jCO/7Ho42rZIlDPJLDuAlL3SACwwikqxstSvMTedCOCfU
whgi1ghY95VipEFjqFcr57Xwnh0XFr2UU6Btz3KC37Zpkytoqi7+qWEElGcreVMD
9XctnfrVGZP68ARCrLSDAaDZmS37QQPFJw8BLWJA1gynTosoXaevBHjE0l3FG3fI
9RUz2UsBM8uywP7Oh66nirXjTtVuZLy6v0MhL04mWBDq93fWDpnfStKDq/6ymeqB
RLXQckHUaev+Lg76nvqPCd2ohBbSAhnhY5I6+fdRkvW/BoOrlHZft0hUgUVV/mGA
jAuWvLAcQu9Eqh0R/NXwyNesBqpoeegy5FahziAOvHuwVSio1HSfZu8YEMafqzWB
wJXDbr6zv5YE26O26BteTgFtjddI8Koi3TYNzxNWMsqxsRMKzurhpVhYFSoLPA/e
a3aFH+I6qwOPEvgPtRTrF5k8cwW674Ur+FTnuSDCPD00yzVNmDK4jgZpvmI2YEL/
paWI1HUyguTfyyuWzoA/ATWLnE9DR8rVxoERpf4nEGDrQDehMhP7Sxhy9Y6bQ2gd
eh24cw6eJhMT6+YLj6hFcU3Fyd6+Ff6i1fyc1vhBwlZfY0jVHDod4h50HbiLwJ5F
hEowYKyzFPGjqgNmNxhiQDkOCJg2235JdBRBjWUgCFm0bnARzFYCo3llHUO0y+jb
XY/Rjms9c7QKL1gobLTOUOiUeBb7xBsQ0gm99odssV6hnk6CPNzOxo/H6CjCQSUc
wfODWQhGGBAAJXpQbkO2iR3KP5BMt/cZB8YmNtKb5I5e2ihpr7QZrGMZ+bXARFvj
NvzGJ92ynhRBMYBsd/SQyXVg3iB/mXN+Ae8T/45D7wVUpC9Q0rCj9YAQGzcoy0W4
5Ua7Pn9Mep2maOvkimZPSdOTCtTasrCbUGlqdPDqs6LwXu0i5orZusQYeZDYbb2x
hddgEq1S0tII2tK6ojrixGBOZYA0JbJN9e+GU2NONkJ10R5B0i9egFdEBj9NHB0d
ih96NCGaZcgMkwVj5KWeH2ECoQPzvSIFXuM5JIk0ouqHByEsB+1/IOknRlXvgLsr
YDU2ljOwf14pFOpGsYG92SszhbCACCYuquM+QKQHmE8VzjhQXZoSNuL/v+sdKxPZ
OSVLqAlscN9Syn7M8hz1PI2RaDWC86DecA81Gp4zW3AIFnKyGd/mT+43jSTf0h/s
tkK+IAS9RgwQr0fm/QXZsCKzRIkuiRkz7Fqh2eU18//vy3kbI2CwTWsIR8shYlk+
1+n2OVBmfFXqAN287v8+zJarrJ/8WoQVqTlOdj7F2kwDfCPjgAd71MZlPt1/6Tqy
tF74OzBlyoJuD1JzbTpy2TbgO1erQZBFhXnsbYI9C3xXy3LPVAWCgFE9owlPhVKK
bcozrS9kAmL8YbCDwLtNV8G+Xg+MW801/GsC6HZGSy6ycVWZ207OUAv1U0UBq2Oo
4vOP5AQBuHMWxhryVv1J2Eyc8tG6otrWYX7CqR1amCOQInjT3dGgIZD65DYju+Ae
0jZ/t7YtIe1Wpwvc4hIEAo5PVDnebEpaiLPQkjrQ+tRFWnHiyWA81F+/5KwmiyYj
WUdR46hAtRkegSyp9cW0uq+8uzxim3TXMZb1U7T/tMZIKYqTwB61L8/U4QkNeFhb
s7QZDWwebRFYPRpkT/wf0A7j3xxpHPBS2Ygm7LWb5aH1+OIIxgEclVgIYuSrTf5X
bbmgPYmoml5YlT/kXRBHdN0cPLr9fzDpx34vuJdKSGfEzMxlFlmHAQt6SQScpqgh
j/THvDAkAZ/EktXcWnQ0ap2UQy/sjlHqbeVQkNKhauRENC9i+yfhNfp3TdNNuf/f
FQzLAuJWX+j+iYTFLtA/djvBxmyer7jOqpZnyK2OAAFgaehFO4I5/pexbv6SDfMb
2b0teU4s74opMgJIahY/Olnf7zZVBFSzM4zDwNkA7uXtWWDiX3iE0Vl2wkHY0CkG
gTBpHYwomwsoKbfT52aM+HhRnf7WL4akUClI9/n69/AT/i06ErDQ4kPk7Gq8HtHT
tiNUY0/OdP0tuC3SRr3x/yGlTL7B6EtWtkxTttGZweovvulCpDSNoEM4buvpSGOs
IH3T8QSOyyj+tA54T8any9ikrGWPefTIVtdkOAy8VckRrEOHiEHSN5ESwbYlibbd
DaaZHMZl9MxzhFXlrUEzmGl7pnJhtB9P7XtObgm2iBdlPFBO1fQvZf6LNx+Styca
85osVyblri5L7ls7Nn3bfuAOaqP+yLPMupNgHWNmgwbLULdJJbCgoGvhVb3iu6k7
UYWSdnduCIOPsZCykms5uqHOS3sWudVn/Z2npclLQ4MSDRHoXfeNKRVYGSNVkaTi
1yclR7PUt/qE8x2sTwvUKAzr72BR1oxTycssTs6ciib7Af8nLv6gnTiIU44PejsQ
U7hGjFD8UzofSKljVDKpQycjCm7P4ly1l26w5VjIvVetLsXVfLjbNgX8US3f7fhO
jbYHB9N+fjINT42PEMZw+sPFJwsBm7RnM+t46a32VrQK+vnkPJ1M4tOq8B7C+D1g
blbgdx4OwToOD7OIEBaXzV4Q6JXI3pzilmkPN2DTIYquW1FK//5Q3DHGERk05cXW
viQNlP2rWdAwfI3sIbvE0fvYnGerSLXi8PuedqxUahNYLGGuLDYF2C7rXdU53ZrS
LSxWg+hwrZegvj8YzVMeL4237rleN/zxBK7iSCkeV56OZEDT/MTyLbnwmwDzu9lB
4Yvf7AeVPp0RGeTMpY6TGLjg7tAgNje+JfNocVKXknWdh6UZF988nAb2oCEzII8q
50I5S2AochIAIx4mmGwoLQboyIoSldyklnyhalr0NsPF/1KNBMlQqDTvPYtVUopP
llNP1ENEQDAlUgQl08TxXwNbvyWQ18cRJmEy33nwy8iLyl2E/cpKHdmGOEoIZaPN
GGx5Y3nGomnO/ea1bQhEq7XqnOlV0H4A2OFmsvtTr4VNKUjAb0JxXkBnrQWQOQJu
gM+Rcq5Qr2r1+0OKgr1b0DeT9OTb/ZePS+THhzy+IToYSw6CPyC0sgjs+Z7PGYEg
NzzGsClgT4YPlEDfCpEgpWd4Cpquib45EHyZGGONMF5cbz593nOmWNQ3amrrVIYF
d2E42FJzxawkqSUJaIqkZ/nL0RyMOIPy5+uUi3JNgxsP+6GqA0QGf9A/yZoCLQ/P
XOzrpprB+KSb4JB4/sOCWLHr1TY9D9s2UYDdSYDf2RLbYSZ0UUFoa7du3jluCEnF
RSCkUIdHFI4xszNiXbjfB82g+bImcAqqLZp/KD6eY0QEB3jhEaZN1F49HH7m8ssN
MIGvwixucW3W6zgy6MNhQl7nUxpTx3WVWcbiuiXtECzwYDIV3cKa3fMglVCeHYFk
D2U4xPXpfKMyRp3dsn+aeTC3A/cVzWDLP1H6trarmhRA1CfMAVx7A0R9hseISkg6
EVsOFuPrRj4bNQYJ/nw4iniVmxvRDGxw28Mg8LW8+vf++2hVjixHuH4x8gyqRBBP
pO9gWGxkpCAs8NRvg009l85xC+TT2JK1MozgR3LRwopJbWTAbnAhXzoRdghIx5dU
+r3KEX+yDnOsQj/NA9iy+pD/iM35kbCgdKEJCARe494M4eQBuCBBjj2FwuRaxdUb
DeRd6LPzF5LL0eblF3iExDUii0c7ygE2bmxx2+VpLY/G9/RleMKRNloifRBHg66e
BEosfm/DblLUDGwwqLSeMUcdJoH9TupuChvkTCr1NoQQQ55jMLpAQhY5yUO3y8tH
MmKhF7SdFHcuySBvRgHFvAcrW+UVzkQyeYcBt+68bs/WXDzNNs+TX5H0toyokcmG
M94mnkJ2sStgo2+MzIi0UshAiDu3nMicP0LCRW3nOd/OkoOllYsnlceNAwfafZPi
2QFf/4eQxPEthuNVOe5jjDFUwwvxRLfpY0+IBIQfBseWDEGCCKsJKJDi7Gi71ORT
DD/hUs2prH6VJNo4Xeh8Bipi6Ra4llIdYS84vbuOW0MCK9h45jBA/CWgtuQDZpra
M9nqn1ldEVVB2QYYaCU6puYqW9Aq82BmIDNtBj9XGH7qqGzwHvaYMoV5cyELuoiW
rAx6eQ5gqPSrVyZocGOG41hB51CZNNPdD1HTsYqbawY/31pltouHM9G2I55/j9Uc
FlFKWEYWAP0hjYcd4msQnhDDaDQfFpf2TTUwpyM8i9l/lYsZIQXPj/Y+Zk+q+QP6
Pbeh8QMWZUChuhdC6tf1+OjaW3UEyR4W33QFCYIGj+KI1vy6iFIj/5yPLQ9gveFZ
r+NjKFplCFwGd1ZHHC8Os7d24E1lr2i7pd3++dSJaT2v4nE/Vep2qATswQS63OOt
JIlmSHrtliX3qFKOI7v+N2qnFUygbZ7VFRZZS7VmVvn/Mdjesv6o/1RBqCyczKSl
gdSZJy6/knMQ658Vh0p8PYzyVwhGsHREh1eRBMWaLx6B77GIzpSVHa0BIG9OphQF
wQ9Vh6ZdLRL4eXwreTP5kM+Ccgwh/1hWJQUV8B04A1PW17MfeGB5blchm80KDIlA
dOebaob54NLhnOTD11cuULTF9jMAl0pGYxDWpuIFFFIH+u6qwe+zqomlXiE+dnOe
qQB8SIqzJggmc6vq9Z5ZZ3FyFU9pdUqvlqCkCUTKNEOO6hT1QnoWhyde5zHyq6ZM
sRUSkeyIvPUNDZ+xbT/D51VVgrabFja1BU/5y5RTnYYfbZpwRUGnvIRfNFgS1Y/s
im1Gy60TYWEAKN/Lx0QYZOQRwuKlMF4C75U/UsrHNR9ETwLQWW+euZQOzY5gWzVe
ZE9y1kJyAstwMPUdOWkKqMjoPqwH+l6T7+V56n4id2yRI5V3dEZFKUVshEWz0/jD
8tP0o4RIeJnWm4NvwG5E+G0gycTHQEmaA9EwNtAbuc/EML3Um0v2rYysVI7k2ICs
naCeJ9/ruOLeg033IjecjuFiTbPeIJQL6BB1RS1zZpJt2YZhVOQ002yANF708tDY
twn2kA87DukrQ2UAsRURPFkvUyrzoj3ITcDSgHBlQOln9Y6zSDbyB0FZJr0Elm3O
FVOp8ZZsl6CNmTaqXyM5MHeqo1961dV8sz44v5Ojzm3BqxDSTSsCrDW4gp9ckrws
vnWcUQhXyeyMg5kT1DCgq51XMA9YEyFtG7vRLGV84smnBULTda7aQiO+D9IxdIWT
/RFOLu38mabagMWwBPheEr7Qf/gD4NTACco5X6M2PfVwSk5OEC7CVp1VUrGP68Ux
Slmg2DcTvob3E+4kaji5P+O02zusKEDXe3Q0ZNceY0x8VXg128JHlKGvyKPDvoD9
cssRq3bjbT37/WXgo4EmcCk8XAvYFVTmrf+ngD4a5UlvIJFx5J305vspjZcJ6zF6
UHexGSYuzKu+Yh6TA6tN4otYjZrfB7xMR+gidGfK6nXJ6eYEEx9DfuzjV7xlVqRt
04CjZjAczJWOlJm+sHYaYtdf7BJY/7qdRUhsrZamCxOgR81jlJjY7V7Ym54IA7Vc
ev8hcPyq0tFS1MKuHld0y4syrL4FLaaIcIeTwu2o62YCQvje9dUlegqi44EWCxRa
W1eeE6Dmlqk1IFSo/26ialDAJvWJok1rUwq/4GfX4mt93TAi5FmBqQv5zJqxIh23
2mPLUDW4oax0mphpRMdFUHPu7mbVz+CcIAEW8WS7LiA0urHkL+p4/7t8UflQxg+R
NmrXnKfUdG9i36Sq2z79BDumTbugLOT8q9sm2sagYUb/ZBcSK9p380Wj17MuVDxJ
quhHvcDEkWjJ2L7BK3xc33kmNqv6gRXVk4JaMGIxpBRMLifzpjAdPlXI0BAOcE3V
5G+rEmXIhOnPRjGCUC3DnMjdj/8MmbNMDT1lc3l0KtQBt72sDCKrYrietHAosqnp
3DvdGInVuK+v1ywXvHbylK+J7VN9Ws4ynRcQNmIn7J74DRDwr8Q+6uP57g5jK+Rn
tnyxfOyjQvo+iszrRaAOoD7LqVjuwA+ui6rsXd2dw97kdLWeYVeJG/ADpy3pwubT
TKrdyWOY3GOyvkJXFM3FTE9kTAjqK9fodOhk6KxWi0g9+OTvp3bsKifugsgSfZ25
MP28KnCYy32KSCsu5PDaZBtxw8Zd1fZmWQgpuZTH2JcxKpoecOw8ru6YErUHXTrG
kH3zzHHF10ucYiA9KrKG2Ej+pOBZREsHNM+LVDofXHZbVrMcc554/o67WsVmAM9j
BErzvWQnKtAvNax1q/fU4uHN7r8bb/oqLGIt55/NC2uweVMDMtvYkif3OooJOiF9
ZgSME2Oku/arEM77bRiz80fH6ZJkwcU7tADPbEFboBOYlAGtA1VUg/4NjempCMoJ
eXHOdrOWMFQYV3pEIIjxbgEu2dT7lOI9ZJNwPDnqBlmFOFBDKghPg/qx6KM5qzeS
ChLu1tGm2/ygI0hoykCFocQEMU0YQ9zmEmHgmhMH4FJhwyo9dfrYlV4Aw3fQ8gJ4
LaURSaKcAzTdJX/KpNY5YkvZ0uUfH2k8kTQoap1H013WY1BTstjQc8EAHP9M00Fq
svxUjLJvs33u4q1NtZOjIcK6+PMzH0rWNut4rxFYKTcs8E/BOHJJhuBN0QSBkwN9
iVpVMUZJkYg63Px3Ylz/ykfyW0yqVfe3xmrjcHmaPQBkBknDBca714d2HYmRA6PX
vro8dr2xflS6W9VnniE1Nq2GNY8P7+j+FoF0Qi4IKhPzg6hSbOGTmD+oTa1AS/Wq
xaltTCO+DwPWtwzyAevnOgmf8dFO3CeWEJqDA0yRy5O0nXPh3aLQKgRWIlpA3e/z
veQ0NHidFECECx9c2Y9ylBqWDnOdfoLgsQ77mlIZuBxlVhSeF13w218w3wVUIxUF
JLTWh1CFVfCc5Zr8mQrZ5pTtCbmsJDJI3d3IZGgmq74B0EK28ndRwEBBx3LqVdTw
EKYLWR0xIUtBspWtkfUKhEynuoai2VJ16AuuFVl5RzoAP0/jyb/gjwBxIo5Tnz/n
Mu8y2GT4H2AwR9txCjkjuGDk+ER8kYDeXXORniW8L2eK0sfIxucr9oqjDbrpB8BA
HUB9tJITITYn5QrIy0wrwsFXVxokGwAFGV6MSaeHenz4TOC88qVCOq8pVCcvb3K5
6USFlBR2M+n8cwn+h8lH00umfbI28eumlKQSr4fcNY/oOoVjaPwaRFmrW9xMmgzr
deuMjhJduWhk59/1I3dc7Eo1imB6GWxSRzMwAVyaw8EUoY5dZRVX+5B7CqV9yz5b
JVY6LBq/sYpGiN9wlgYMaYMYBcKU4IBoMh96C81hzDzK91pvD/2BtgzniFSnUEe1
hu2rJcgl0qoPoZb6tLrbkNN92WU8evQ04Il0ThKqg1fp969QlRDQeVBbUpoJnwS0
OWXaVvgPK/o4FTOuXop6AlgkxS2aPmoIhmCGt5vJ1sAOJfW6KmjM4nFulKKSCNfZ
B0yTBY//x1Oc4T1ZzGQBwBWAu9DT7WWCcXVxCLE+TT0hpkF4YvsrdUP0//p7M41o
og9/GaqQy5/qM8h7P1vS0yM2HQyJ7nJ4QYxId934gvsOoT2R9eCdcotuSuANlijL
R9lWybmjwWUsnRj9gvBepOFzPRXXSkf2knnQV62a5CF4W7wQRxbxZJUs3/8nUOsA
ez2rveA/gQl4Pi1GGK7AMibxTIARDRND0h8iM98rOySoXOu5czhcS0gy88je9YNM
cWp2/g8YFHxY+7F17e41fV4sSDGhZDd3NgcmaS2lLrSM0tkc664UelXAt81nUgiG
R6/FxymL0Ighf5gkM8pkN0FaYASRPxubgvEGQ7spiTDljkCTpVLNiEpKi7yTjjaC
tKw43BxI5SSs59mRdqhHcedE+03xXbLEvJhFXCw0WFvnlwJVO3Q4YnQ45USNrO5B
FCMy/pfwcpTZgT84S/ZNfgee+fuWSqcrZEijh+BliJXzR1cLfqAcVhaTPVBP8DTR
gYqtqM6eEi9l7K0pcco3M4TtoY+/c9mR+9bQ9KqH+/VZofdn98AU1Ba2xdZ+4ikd
LGH2/FG+7mc7am/TCJBvBPkloKp1y/VW0jlic7iFGu7o/x1EfnH7KILIl5TNXM8u
lfby0OjGO589fxlG4NC98p4Wt6P9ldML9mfT7WTiV0TBYtrRIc/Xp0YhCm7iGN4X
2g00d+Rl0dTJ7N1qeaUsDj2vl+0X3Z00rWVuTVGCjfEyIyPo23JY8SVwWj3o+xOo
xDFItofZ/NwiipqJy2xnodKQvCvq/kZjZycKCcBY/rlmrMv0ydnw8v1bDb5GIzKr
3bYPIwPBVdV2uA5soxyfUsLstaH/1rhtu7/piwqvdcXaC1kpIwVMLSgQRGlOK/v3
3chqJazf16taUpAlt+znkeqt0ptn5rA5chY8TYBoczLqGjUJvvPa17a40/hx+6/p
2l3bTLrgf3h6vrwqobxg0KivVSTmuL5+eFmnRNRdpFu4kJsU8496Hblj3zmXrYbd
/DnC7tLa6D/QzTbxXJe40hVAjGnJ1kQu1b6gIzUtTOzZ3RASrQGPFZXCEQf1AcXT
47KOzpA+9csnm3ULJhb3jRluzLDK9NPmiqfrSp0vS/LaM8isrMJh+W6Fr4RrYH4H
WyXWzGUxOSA/8cLRaejPbLDKKZjqMTiX4PjpRGUikKfDABBqW9cYL98k5qMCg8B6
E1Vmkm8pC1OioXQFmsndLv24WrkN+i/tO1ntBh1DnBs1u0RpwPxQuZf0lxOSQEnW
mf+4itXDauVO5KPPm3oqOiirWsdo2b9qng6sITl/9U2HEEMB3wYXspdqzr+2avsZ
zfN579meDCUSHx0vDgoY7cpvZjydS+JYuF4H1DyctIRB8P4lCJYUzIHcSHg9lVyv
l9EfGlAIebOSPA+ZBUWrl+TdkLV9zPJY4eet9s3p8i0ptYtYk8EeMGYpcBsVMOT9
JDGjUN/cbNrxl2SzhmIkUtrQo/LsAoRodNwfxXGsvXwKp1gk5zB95FC9XUMIe1Ue
OufMuZfbPQniQjo2AF/6MJFxlViQ6XM4fGm5DolSdhPsXJs0LsqLFR01BkepSl7x
CYDykbkperJekDne6ZDbpD+nvVhgZStBnefjjB+9JacVYrCltbhCjEXHjkGIPo9c
nahznq+ze2/pbDnPbhSLVCtWEW8lpXquKLjjqWa43w4Df3fbg7HZHGkk9AFkICGq
9yozO3ONOg08g4Jt8olmvDaPGwAVsk9ZhvFIBq5uRGGaCYSPUKWu/zgL02uMmiX3
y7y8DTqdNujndTOyzR6QuRXh4VMB4TXoX8hBXeNb3lujzh2jYsJhoTECGh3/+3io
J5x8fIlfjLjcByMlCqGjwDaekRKqqga7cno1odIEDXWK/my+Xd1IO7N7ljGiGZ+E
G/j5Rr5Yq12bc+QWYktLoabsW60u/uG+ZWSobEsdYssjZaiFD9CK1hlR+uVic57d
ECE2+YzxRwXTlpsPgt1STtB2uisCIow0MM/YUM3W4w/LOxr6NQlXL29ZQAZa8mRE
xnTM/MydFFXTV9PyKA0qOLoc3ds6IBe0DHaNmHq4+0I+g9k8puZl0T7GdLS4yenC
LpIPnll63GWDDpk1qyGurD5MF8AwPpnzc22Bxf36dT1gsVVzpCM58jzmWLfamAWg
wAXDvDLQKhy1NwXwg/FFN0iI6Yt5TBIYWsXs/AFGr1JlGeauCZrbRexXjLLorF2q
4HsshNmv+/ztEKs80FC4PNgW5v0wISvEkrW1bEZyKr8dSuGg0ADrzasHg6LFVMhN
Mms4TK7SOOaRAKuCRtYEMCyinJgZ1g5LD+bo+HDWABayWcK6wWpOtVwktxVFqNl9
57Ay4XWdaAKhzBRNEXByLaQm6O4v+aQiPOnXUcVBn9FVFXKGttj0Y2keO0IibCXy
XFlupLb1oVp6PpWAAKKkG68Wxw4DMvfflVV97UrizvALROn34Hr0lmrjDIz59TtP
yCHWbCminn4gYlPPpsfqAXPNlJmpO8ZoNMaotnI5OHKf5Kl9EYO0M9MJjhyxYRyo
9vztB6E8VaAt0Jihfa7EgbzFrCCzJaJDn0r7FCfXNKHdDFGsPEnCMZhOEPj9M1AZ
pM8AkQWn3sBlRv4UG1UXfigXWvD1IdIX+A3GiHlayuQQXQshiSvm3aqwC3Etsrbx
wJC2AW/juPS/85Po8rdZpqTLQbtB+Zld2SeoirUgPfF78esI7Txbtt7iPfLsX9yN
zCKHYaGQXAWeMeDvFPiflV0we8ug0ixUe4ZWKL6VrZSfYMs4vRvto3HCt2WNLQgv
+5rgAM0OcuFmS37X21B2r++euj8FNh79z/uGI+jRkhbacHztAf17/ltp/VXEYXjx
B0Z5/0up7twEfPltw3JWjhzex4TmXWbELmbyyiUqszlGuRazHR2BV9A1dkBsoI0Z
vN0prVQmR/+Q2uHMphKKE2ampWO0jIBKe5ZGzxQabKh+PWsQEGICKuGFOd8j28Li
z25GyhO8vtkgOM4AtpguEH2GElfM+KElgrVZnQ9O4MHVlTMi+DUCjhgq1vpmgWqi
+x3JAHRjPhPuzhhO9l8LLti4TZO7aSUJdA8lQLv6CGO+MLYN0iQqOeHmuw4eTBBv
iX9u3LcsfwDqhbwbTHFnuBmzN8MKidw6wucvcGk5j4S7lxw8BPE2WZl2rcWFY8vQ
r4SxepFqn0rsm+hzHGCAipHVV8TpjZKOaPmJUnvCa9uzjzH4Aw1Ld+FNr+44WV7C
YOCl0P0eob0DNk49q1y0gr0XAhNEfZSqJppBcFVILMBnA+5orGJmph5TVXA2BXAp
UojikyMnExHkubQJpjgNvoVvtUBEri3KRtUS0ifmbkhy3I4pPTABfttHOy9phpLd
vSDYkFTjthzvq+XC7r5q+2D0JrJpDqPk2M7/ZbpGDcaoZkhqn+T2uy3Fb74ICL4j
iTbklqELVIdNAJuN7twbA6xBAzBfhv6YEgangy3sqBnNg4N8nR2K+/wRTlkTm3Vo
fK9uIIYhXWdssCzjLkp2a0nIrQVVjG4SN0iuBX2fPkZLcV98T5fjGomE6ps271Oq
yT3X0j+ITvwMwITZ64b1WKIZQBGQY5El8axgjwUSvAmwwKqAM12FXsIKfyZv2Eu1
I+Jy3eJDxhVJb7ZGp6LTUFUwot6U2otPeZUEgosVm9ChwBDLqDV0YfxKv+CHzO0x
LahDZvNOjUn8kh/aDa0kVCOCc4BQ0XFATiCXIy/HHPmEF+xtRFxj0vU3mXYJ1vmK
K92bbf2e5ntMnxKJRmOi9sFC5B3wCZhpYxw2begzFVH1toJl7P4fq1jXaFGRPzjY
YJIOWKWbp3HUBIbelZO+9ixxBNWsQ8cZNTde0iOTXJZGvtOljIhD/1Ze4d4iMylM
qzFYoNNh+eMyiKp2qP+gvweCG1nIiI0+sk0FI2JCcaNddeLKn3At7cSk0rHWsUCn
gHezq8svL7ENtzCx1aNluc4/A4xn366tMg2p0/W88Wo307i1Yf3DHIo/qruvZ7xE
gJKNI2SgQQR/73BlAT7fmuClo4z32ajPhS5QhBtZ8psyU5WIY9VuCcYEqH5jivRz
oCsJPFat5YTeFlhArJ+MJfRKboyO6/nD6AvARlDVXBNAwRfWi5nvG9d9aybVNunh
ugGzkqCuHqH/0vPz40AP7Jf3tJ+3wV8fj9ko7eGFbNl73Fd29118h2hf65vu9Ugz
PMIRFzBIkM0xWqwUw4R1PjmZ1kwRVb3yemhUOtTOv7Fl/y5piNgVOi9PwJ0nwzc0
p/UVUK5L0nJcR/W57a+5ZyTKPZO3er/JbsifERmet8UcpZqICUGiEBUHBUAoFYGM
MZylC8bJNkMKXb+e9cP+InhO7NF5lG573u1rJVLhMp8rFP8AjIj0XEfQ3YdsWrK4
h5Keq0iggAnFRzQMhxMeZ/Jk8L6JUzWdrnch/zziU51pXttGKVicE2h3xGOTGElu
wgdq/Sg3axYFbuIaM2KW4Y94qRpByiSDQeVcBPWIr4E4ZG+SD/QJVTzL7CB3hRmg
36uxZaMdAy5DfmI3s7N+sSB+jErhSudCpZuMK94nlds1dGYl1DoWoJqERD19I6CN
Qs87Ec9l9z/aaj9Sfmegc7ed+Pg1OvqISMnUlksF4zbKVRrZroSvpkc/hHwWlU2b
p22lgBoy3sVgalfWhNhBMd4pUUmD2fu/Qff17RG2eQggSPyJZ27JTzNXWX4ysKat
KLELpd5zwGsbK2VsbhdvDgZmXJcXJGvTZ+bYi2zMffW3BIpFhcCqdeIxReU7MRxN
beg/M1+AyeskFPMwViMKopkZQPedZC+USrm49DdA/Ue4Ug9qdNiQctFbT5zohOvf
6SaKi6fUfwl9YHYzoDbOb5TSbt8Dfp2gtkWIm4LDfJ38dJSccA+TFPU9FLxu0cQD
dzZRjiXQfJy2SLIMtWfizywMRQ9mi4qyizT4tQCpAg108vmGKrj164/VivHxAyKd
Ko0TYbPOTPUpmlY5V5PAKBhUQkjLGJPTB8C9iy5LH9vshTaR8k2ftXJVnMyrUXYr
+MEkTbOk/Hm6HKtFGHb4AFa0qGOOMB9o9CCFbumxtvShUsLusrQzTWZpVJzO0eA4
p0lUrffuMTsw/yGQ6H0La4thlWXzojNLZb1zsgztdSltTidJYiNwRG+6tac4o+zK
jQG+698phR04pi/VC7InqxYz+cFnsBlIo+IYN924fWh8ro0m7VW27rvqdf8MfI5c
xToLFfZuEZGzMr2Sq8EiXJnJt5Zj80IHdr5cjgZSdC6fctnK7uvUR3JUA3nAAqx4
h09HRrCSggmN7sLBuWLdrJ2EWgd46QWs4mjrVPWPs79PLchcc6yx+/4PfAXoyWcx
G26MYNfKBeGeLFIiFBn6j9ehxjKXZ0zBIsRX7BQwmjJOMLbqP6TxZOK1Nse/EMrA
Hkfqv6uW42COIMuE5ZzlFvHUM/4L96/IlsAJf8ioZZC/lTXpPwuYDwCK2yyoXywi
L3KRID7EaRPuHnvXDabonOsK8RZ5dgeckqJ6a4S2xSlvf5VGAyzb6QClvr8ipkho
xebMFQ6WSN9Q4oSmgQ9r1+RTOwjQ0xVeF1RNSkKBmnOPPjlMUv0akA9a1unEf5E6
fDE4c0HjjnHA8Hgcduupz8LPEpbsEgFx/gKycJaBtAx+CHyHAMsFZj4+FlObIw32
tHMYwJett/MmPZCA445QPAfa965KPJM/0FLu2x5bsB6Evh269AmepI1JOoGSm1It
hfOJbq7i8lmFqEy4P9tWxGQ/pdt4jLiVhLq9qBRjUWuoTbP9jvK7CmpSM9KBAZag
DPXSJuThN0JGwTFIQ8rmZNEsG16AFwdfwNZZgtEB1v2yj9Xz5L5FJlfBYVpUef7n
B60uxGxs61QJwmBkiuwcIgsDu+juxeTh4xtgLT1mDxCC4BYutQC8ErtzWJWU3V/d
yJNDf94q6RlBiHvp19aX+HGkS8cPcNOUcJq3R7Ow8I0vPjezx9HenbR64WJHfaIh
ddtzSn2ntx67cM7NTeBeHHA+tyeQM8OMBHaOAl/xc6V2Sizzrq2Ye15s/W5o6Qxw
D8aKfrbSbiMtd9V4iONW2u82lPvBkOeuTMC2sKLTlpYJpdGqfuSbye/o7wv+JyVK
DedQIPSjo7zT228m4SkbY3LVaEJ2XbHTgF1OZFAPdc/YGbgHTaiC/ZNQDJ453yTr
eIfWs5xwzF34oyz4KkGB6dVJ82qk0zixA+k/sHaRh3t1Q/3UgQdEgmfpfi3ktKKs
+r8N7V1qI8ht5B1LfWXqW39cTOZSxIZ3VvVFRncRtctX4fWFil0LeJyDFfkmB+Kw
Jw4m3cEP6aLDwZCCdLGl4kWqo1pGDgNz3cAD4S8e9wt5KtXb5Z+69mUfAoInrGPp
/EzfdWkBQnO8YCE3haorlGqR8eld802BVvpNpJUWN/UvCEXb3a5ZHa1DHcKci+fQ
N2jXTiMugZ/8x97VXclbcQh9HuI/W5TW+ap2idQZOyVadHo0kC+dG1+JQdXLACxi
m0E1jGgTPUG2iBvicF0xAW9A++xHj3vp5sUMQ9J1hXMUvR6oWRM4dpBeySUSCw0/
Vx6DxbY6TFVSICEH4LaIZjqcCvejOQRKD2xuZQnn4dJGFOkkbwvOZbsm5MR/s4jm
KeJMf8uD3SUaaRry2Hpt2tjpBSdWwXISdiPubQG9ZWxINys69r8m0mrczDYkRTNu
t1ShiSc0JOyUKXLY4lAbWtsjEEME7Gz6dSzcVqPUI3IFWIVUQYK2Fu5M8EJYAHjt
hVtEII3+m9zm0BOioJq4BnPM9EBLe5EOC/moSvAmEhyUZAOmAM2ZK3LcePeIAIOJ
Oe2lqIawd6bcuGZNvS5v6HvbIBeKFm+bh/mBd8AlOkVw2m9A7leDxqSMqeycFJsf
IpqReJkQ6atIXb85bRG+KyfUbWugom+GORKT/B31Qz6BSsIUSEU8cUsDa8TUFpxP
74M40OJypURmPubnhacf1UiM2i06a5L1/+sz6mwxPTCzJb9DVsW4pXiybPYx57p9
Ug3KV0fyd07iqtj2J+bLiro5lZuFO9DYPmCUG8I4blmWODVjZqjUbmhEUMc1LyHa
//UH5wvUhB4WjRpbULjvXYFWaC5L19YsE7DipvdT+c4PSm3T30FMo3wPW5JgIj8S
NTsk5u8gy2PiKOdDlSZ2qIfGwbytqZ5YctbtozhdcCFOabian9UesmrmItnwuS8Z
u0EzbyWBbYs2xHUL5K3nuGFtSHbQ/a69zURDGyDbd0omZ6Bdm3GMEiy6YrXuf/gI
Pgo+VFR+t2xQfWdI3dUc9vvLjuM8Tax5deiJHhUbLctaXlCf7irZtVFH6sio3zeZ
6lV9Gur855CLVH1JsfWys2vtCrJK8D2nK/lqT4FV5Odc1FKP3MLPjYw63s9KrnFw
glJmovQc3xfhM/4dlKm1RkVi7MfBDZjFHFVvOqxyXzU5KL68EJCiXODuTWJx5rMX
u5221FD0vcXoHQJ86dAGZrciUcplyjVhUx7aT/QrIOFUEq2e4U4wVASStcegDnyg
ddBqxWr+L99Z8pmvLXTaFAepG9r0LuNpLIaF4s4kGbXdJh7/KdCDFmntZ9jWTqJ1
VD/mdaP1/oMMDnFynk5LdbarO15lGRIP1sx2unJQSZ516bQZxagcI7dogaH23T1a
6tZ0ivZgcmvddVDhW+Y2LB0qYHjEcEtigdxqkypSC12rhUp3H2Osho3UAF2UlJIq
2ZwMTj2QxXecE98VFI7WIswYMNhW0RTiIyCCjpw62Bt1fJqXGQAG9WT/TKq1v9Kj
+HZsjQwqmyYeGRnR6U/vnl3Ra4fvR/jM81rzOK/BhAUXGlEqFkhlsrEIOvqUdkiy
Frz1caQ9fM5xZuHWRu5VcPt5nGRyVVBCopV1KT1y2TH3ILht9pV/x9Ki//BM2Lpe
8pGRupTldetNNspdSYv4Kf4NOTYVECnF3UNvBXNA9p+Yc1akOp9fBwBGyjh5XAIq
R3OMc5tSdYVnXMPJ4w0LY9DqVwnvTjU0IzFTJ2vFw4GcKobrjhInMDxQccIor3UQ
YyYiBrnzz+DrV7R2ZQqkJBC1E6U+2DjcnpMdwbZJFFKJMePrMn3ynAqJrhbU7NYz
05IrMjc8sqgSQpx/d9Wc3wP7WaGnJRl0u17jLWKWKBIz1aLbG4p96YHhim5jr1m6
OmHQ8cg6mjHTtx3D/bMAbl927sP9YQPjLO8uO7/WOj9olcoUcbrbqnb15uEuTOe9
loeGh7T5QpBnno6NWqZIs64nCjFojSeFY81thQ/PxDb8qrsSo2dTbxvsOrQbXyqq
62fGHNqre5I2cxpTDMczAqro/4lD59r+CQLEpvi6u3tJhCdj1NXe0diNabmrlY6J
RIC85NCyeaKf4gqxVW01fiLCQCpY1C088zyMUAG3mqwjJgQ7F7dgAYDkvUBuLukq
pV6/TKbJ2toUzeHuFRRjUzGbCrBs1fH1YTLp9o6Sb2vHZzla7mj1rK0h5fhLZKym
x6PnCrqioj7awXyA5HAmsBj8MfS6/GG7uShG5wvxsLafDpve3HYloODdgD9AkaQ8
5TIQWgSkFen+8RreQ+F3yYMENJaDDiUWCxbsFS85f0SWjagjiZY9Sw88GYiyXrQG
GD/PzTS7xpFWrQhkkz5ZFekn8u5J04ZoI5ajJryWkHSYSEQisxOKjNApv1AUQmFO
q62AS9VfBBESzrXfWcCEIPH5s9rHiGRA/3PSDtBfxmi7LBWPMwnKDtc6TX1emhSP
59vXDQLSXEa890zqMHjAV3uKHYlT9wxsjIMwYYHLdIqs/qtWYNMFSvrasqYd/77A
G4mRlVc4nrX1Cwl/1U9JlcaBePqvaWRLZyrM6Bqr/ZpbvNSIAcZyaoPvo2tJFIc0
4GSEqrIFSu0qEh1tKDgdNJGRSNzigUXBCVMYfu0FWKFxIr2bmFXxmfEcP3wGDDpV
k//WhGXV1MXeY4j5lRNlaNpy/3YNnpj9ALyfeDsFdEPUFbJjjqQiEabDnZWi5sBC
9tjmAO723FRfHPkDFfHT3tdu95n3IZu9Iz3iH8f5OqG+q6bOp+/JmyZc5vtp0gL/
mEFLdJd1spux67b3ZOsrinLVnWfXf34Z8TeS/Yab2zYjaY4VIT1Wg/fMqTsmGdaX
zOZ/KdOTWXCIdO28hXeYV6PaqCErebb04oZVIusuH8wxEzc3QmO8bJHjulM4Ofq2
RaMfQ3MQYgWfIIfZE6rcUSbOCDnL/8RL0cYpBSsitHIHciyZZhOX2vXu4uf15OST
5VWhde1NRDjdxbpsR6gMbq71WIj47kIviMEQn2xMh56DW2j23ujCDa7tkkqkqNdX
YqXlahu4k3vJ7Dv/MjaEShu/zXQ/2fK+2J4pdNDxQpO5ZB9yilCrmUo7SpZyqGvn
1P02HXjBUy2gNc209BTqOJco0sr9mSi96WKb+SDAItSsIOqiKB0It/xb7oqA9CEF
ntFOLthsu6e2/8OyZWvYnbnPqKZz8DJyTlLtBGD7HNDGp+3SE3wmzKOwMAJQmrrF
xmI8tYmQKgXmlJaL1xZ6bMGFYMlftF84G8vKoIjuyEVzMjo3/1/e1M/4OVY9o63A
X66u81EjUNWuHjA82weRv97VRC3v2uot3YHq1Zm3xAkgUBp+P9LYm44e7lbM3dAs
CScbPUyJ3bMj2P9h0NBr/jkxKfO/4ViQF9RqWTx64MgjTLqLObrGq75ZV3vvceKx
o74S27oJcNqSgdghDlliEuZovpm/2SGRutCGVb20kW7siL4Jhv0HsRmcsGa/7QSw
WKIr1CA0BR1gxOr3KuDxZislLZdhw/JI1jNnj1H/wGtQkvTH6+lFqpjXkiBqqElB
ryzIC5bKwOvOeoLPON435dL3H/Z13kmNHKfgdaYqVRGocwrW/pIDv3IIP0/G2/Xg
lUcshwPHrwEgJIXOu+trDG2cEeTI3NR/yWQTtGkCBWSpIueUe6iTQ80FTHyP2zjz
wlc95mylO2es0EwhYZsP9quoigc/7uImn3s6poJQ+34yQJbZ0elLFFUYbYHkOVM2
BJ5R45cORiLY2oMPyP/W8vqP20fgjLiBuimQj6Kc5bKx+vY2y7H++qcYbYmFAxDN
vGkDRTESSkpOCXf3/C8UVyNN1AI6Ah1BffqyhOhMvwYeVj4y9rKn79FT/5HBtV6X
bsiYzBUOY6b/hg9ZHPoNuhcjY109bEmgHjMkdvXttyQTswzQ24a5jQCaZGIn+lOV
1nMvayvRMLuVAjDW4pb8cgwhz4pKCLnd56nreGXFtSJoMN6Eqtnq6tkUAjgRKpdv
+pnGW06pnC1VHhAOrPMyZn41JnenOZCTpCOFBMkUdnWmMKC0bXWbG50LWxyv9zl6
jWQ43sziRjpGdf36dao7BHn3uh7SaElZyApwOcsjXXtR5ZGTCFItHYBaF18BxGn7
tUqUwKXUOEU2SFlM7pK78DMVdWUdHv7TujbSxX3XepArbY9FX/HD1hqF5WcK88vH
QRPjkRYtxVKgnta+fr16q624pgXrWHL/5IfEAXHNXsXqGRwSHT/+l3esEpufzzCk
2NZDLUvN+jaOojr2iWmkNSCHTmh90anUYWffUyjjSTbwOKcFnNQCsSyjtskSGLLO
Zq5GVqtSMWuGxClm7gqd4RoO+MJEs4eKmV5Xfss6CV0DM59AYaI9ag5rq8rB2WFX
Vl7rYV9ghP1rqZfp+mftlr33VTw/88+RuEaFxVF9WjGBt99Ho8cbq9x9fAcxyo3M
cgXd+YjPa3LYRxncM8ELNu/qhLSPedxbyjslHWS7Kywpi/UEVJf/Sbyaqp9OuCXE
Ye/oFlKUxXzuzwctWtHtmMYpIHdgFuuJe9IBPI7xseyW/7K+UGV+iAW130OF/a/V
4NJUei+NI0Qr6yT2ynROjfl3/vLl+k2NFa6wJ0Ul8T8f6/q5zPps8uyrS2bk289v
nBAlJF6V1FK9kohTvmKy7tgJ/gze9I/JkkxQhDytYtcBVQyj7Q8qMIL4OaCmKWlb
1AsywC9kz+iUB9l1IWeyz7XTd9VoFrGcxN9nOeNxD0Zk+GSCp/RMWc3Sqw1ozIYN
TOZuomKVTkTmHvG3AAYm7/3iYuywowMvSxgamirb/I9ZXCHNV/uq2K+GbnPQ8PIb
9hVfEDWTpuydaxSwQDSAmiyxDZqb/oRuLRlhp2kXBDADZQs5D3ZNxSMBxQ7JI9kB
hH4XII3ABMsRByE+kWLjVKfxGdzpChHyGeLif4I3XQmJcwAvtWgRS5P3TkyZLNn+
PT0qRNeuyT1Nunzix7TBRLQTPbcV7m4moox+UobAOcgZqS8Biif+D/JsCtqtvZTE
qp80evKplOazLzYbcaU3F5x6vRk/1K2bL6uC3pUwWv+Xri0w+B+ebUU88hFjF+Ic
gx5FdhLhkaGuqdky6ItXiZ0aWBO+EhJib7T0vO++AXINdDe+VzJEStNA0UXyfn5a
2Be+F7yPGV4Ep/+aFsUmFSfwnHxqdZl+YvOUJNNwdQ0WSUa90nxSIxlGj7dKh8Js
qL4u4btl24iyCKXxnxHPbIxkDNRnFAcuY4FIQ/f0lmm29IJgKiJHsrX9Gd+9pJsV
+9w2CbMkaPgxmldw4pQ8RWogNPy69zzgy1AvnqqC7L17fYaeAlw8YPzTDQcgvilP
hy2+3sWNTRuPdephvD1Z85/uulpxEMhafgRHmMJoeU4YKxeJ3ZgsHZFqPOwwKfVF
HUEKmdJ6qQOQy4OK0eehY9EvGB/c6SFux/hOdfiyXHF2ZcTMzjwi9mCUUanhkJsx
KntBPhsHHUoQ6QElcIPp9LYUc7Kpm6lUeXt0kmWCXNyfGHYkIO+VVWy0GXlfEZVH
2j32lcuvtQfdgsrbI6MpsDQu2JPFMn3dEqJ/a1TlWgm25duzcBqKqu4Q8Sj9OVYj
PRf2hPYmrUUF7vQBxXrilPUf97Qy6c8VF7uwi4dqmLhbeKFe930LKRsnALpOK7Ig
FmrllO5m/1py097QS3qnkSRWOfHM7kb+VAwpiVYc6nzXNIxOt4iGphrFHnzTyrVc
Do/wqx4p9Oq2ynSgzcewkRK7zmE8Z9fmvJa1fQeBPGk/NodinNqf6qJZD8HtTEs6
YChMdp14VJLcZXViHLXS/Z8v4tu6hfSj15iPmBFDO3rNwAtkBIRaH3jB4kHEtKYZ
rUPFmVU6WVGTKe++KX9bCCIyeA/Lq+U94UAXJzG3BSr5ikHBF3WfnIIjYmjdzsDf
8DfPs9AcYmPQq2usavHPGFRig26W8mYqxHjIgnHv4PjB9gziIVuVsUjP1i81Zgs3
Ao2YEouOSlAGTeWDbr0e2uQdmy7VtyxLmue5eeww8BXxJLSNb0kF59gvpKkwppz+
U1+GufAx8TFab3Hdt3wsDSuk3gQmcgJinTLipjBRb9+loVJTXQjyXe1or8x4b+R0
NvEbq//TyNHHgUa8G4lX+yfkC9Huxl15Fx1drShT/KwW2FaD1LAoKCFGAZKl63t5
t2HMcdWYnqTlO2kigU+5khqgb0fw/1bm2J6KJ0Wby7mGkkLt0XvHymNqXYg286/J
DoDqqWxKPxqVC46bxhgCfhtcltP9jWaN2OvpDgcmY4LbYkvRRXT2W5RvTzJcfI0k
LoH0YgB/Eedt5zcmeocv60R+l+dfsUuEEEa/cFpUAhIO6UaxSlV0MoraDg8pnoop
mUn68fcPfEIIRpaChFn0m9eRnI6+2YF7m9VHcrhfvcnvY0z8tDK5VCe6AEHxZeu7
2DETpDqXP5tQRK/ZMNjCRlmmI7FYHBzhCOZFgs4SS7r62inVwD1K3Qsl3IrI2ZUG
0IxTWgJF8Qaj4PHYU8e9MnLMH2OrkvEa3kz4KSNqbuCRKXcuGcCmcvOKS4+y2UWZ
4JZchvUAvgNV7kzbi3QR0QBWYGo4gw8cbRfGnZDJ6H+3tPhRpfCRyt/bru0lucLE
T9mX4ydUUkRdU8f9b3caA3qK5mVKwFPdpq6y2BeAQnWZLILScyh9roR/O+/u382E
jXE7099CRgswpMQgJZUZxBQH6qRxm/XqpnioUZ/gxKBW62zOoQO9wyx3CTtf4baK
bvsTowsua2KZiVpXlFTpCKYWzASLJNeY68lkuUmTR4aU+BbWFm0NJ4OO+RHKlUQZ
PzDxjjcssVX2Edwpj6oXASqSnTInV9P+9b6fuUEyJ2xCmQDSU8b7OadOZ4e9dVws
wFCbAdSe2iCjKTWPpJquHrufzXcCWku54PFwG9L3XoaZb4uC+CyKZuH1n1b7tpI8
Ig0HfFVSG8UmfeGcYRTtbvVYj1Z4x1WHSPd48biKdy4THLQUVZcW1K1D5RaV2Czi
gkx/1RJj+k1qFu3dZ91WurjY3e+JnJgWcQrsxGtLaDwb7oN1LHj1OvKUwuHxBtlu
wu8vTW0GeeQkXzYpHmQ5YHD2ywgKDSuZHqYGX1jSEcdiV723GEVl5GjTQ5TVX4I4
qXyBPQBLHldc1qOHr4Hg9fDbCrCNe3pN8BQ1Tk6xgethv5DJFnkKs/Sat5vo/XOn
boHLLO8t38Mp+bvg2auy7uTXaobtUiaAnaQEoTmPZ2YztcajXv2/wZ2GCpEfYFwb
a83lk9nSSim+4xFxiHOTbdzfYrLEzFn0g+Qa5fiMMW47DOczNw5m4knnBSZ9RO/4
tuluscnii2Jtx/uhtYzxnNjpcCB8sR9f3GtfdnxlxIfX2IVkhDWDEv/sgvko+Gui
sbdYac9ZVnUgAt4dZMysUDjP1H/jQY2NVhRRSWkHkNpqQPSjT8KMvY9bZephJMtR
jW2QoWCQKS2pkAG7LBevOznZxZ9KbpmKtQ7BMlWnDjybXd7GyIZjhqPsWf2D7MIE
FtOWiyO8ben+np7R0GN456TqqUb/bOk7SpfnSarBnILciblSLkZVuuyUyVS3Zmp0
Jxoi+pEXDdnSDy1f/EH+u+EeXLbfrb0VCOOxjEnuf492pGVt9RN334sZfj3HSXVy
xmTi5gd00hdT2KALlqJHNjtCjZtg3501wWOVJRRbGPFQPcE+crPoBqOwHAgSfR21
bSinhbFEto9t7cNLJMJ5Ts8EcWDgyHk3HaZ4c4PvVOp9HayeoSxcAZIFsVcmrhn6
PuEvPNORJqZEHdKx39F3WdzmP5zhV4LXlS4xbDHIkXQGQ8WMeV2IIUOJQ4SGJ5uS
0897+Soz/5ZKZQhzMpCENwiUrgN0plYGzxDt+RwfiVtoGfQwd34kQTdQu3V1wrxB
7oo19VRwN4ByxWx1N8G4+oog3lLdv1IR3IUMUXv/Lery48SXh56dIpr2rWxofB4g
/+nmngqh63qcPz8n36YhgOZA5KCk+d6gBHh8FcmfTiO/AV1yXBiga4WnI1IUavhM
HPmh0dBISni50kB3h5x6moOsK1qIPkWKXzvNrtFwITk26/wRv6utw6XqKKHtELbp
pCoEahJMMZRPpZKg2Q3Pqr+Jd18XctSUvlHlkliNrZvj/sHB+3e5Ej98pYsblYaI
r/SOuXZhWgtU/G+EaDeavwJBmgvs/zkmq3fsOT2G8aTsDdpsXjLylgmUf+7zuWLG
6fm2162chYdoc+OmCsN21hhH9eou7PuL9rdCgp36ADYBLddYGLdT8vctP+J1cqWU
eDHhctAFbKbQCcaxSD8RwwrfaJEe9ieS/nyk8Mo3Zp16jccSn+vUKb/Dr3j/b3Ga
oD555qzNzDDiP7pJyseiS68kUD1jDQh2m2JQTSx8q/HfETaxXfBGaPTBFG3R/lSQ
WaioiF8pJ/biAnDmVANJVUBRHlHtUyyeZsdKlC8ohbTdcxwq9KBUdXprG8z5fR5k
m1Xr3PfrhQPsBB1Rdfk4Z+P90MsJWjFu4f0oJpIGZVaTdbuafutDPmuHyRiqhvKM
jnRetFNHK5l3ZHi3t0aR703inBzO8xRM0PLYDUu3CplWz0lFuuTz9Fa+c3rTIsyP
Vn4CM+Jw88lCShdrd0R122QCmQIgwOey8U9E5Yq59gLNRVuNgr033Rny6LlwxZIQ
yN4ebQKAFV09+PRgi+dkpEBW8g7mIEKBsEtPB2BsyAu5qkCN8vJczrggjNVuwbu2
KsRQPjD0S9yG7mCCZ4Ulghk9b/oNK8Gg+OpC+yrGXXobxWR1yHu1VBruDnkvmG5I
cgbPegSRR+HKMAENBXrlgA9tLOPSP0a+zw7NGd+yvPYowowpm8k3hrSbH8W8TAwp
h8i0nDS7KHeD5omvdKuj2rF7Iwfz/TkkNtxMtGYvrMn7Qs1GvpMVbTsOHfVO5qRK
yg6NWgDctKh4rq8117vdZfWp2tfdHXp55F/B6aHTzJdEnWNvRRwXQDc8XBuqdOFf
FqOedJBtDgXCa9/3K0HRjQbeawfdbeMbBTDXK8zKTGJmWuld1DSt8tOzyKJwbzdv
7V+5lLZNsiJz/xBJWmoFGn+3DJYaflmkvKf2BaHT9vJ2RVT3BWaM/lHmHxu9sZNs
MTlNo5DUdN+ZDx0FDP0teH6pp42CfI+jjTQNJXwHzdN3XAHeMtXTB8XPft3AUXH2
1Z5OjF/QHMbFmJSAvBpUzPLAVc29O4F42bBCTjhRsn0i2oXUV14SyI55LVfOCRAH
DIFV+9x9J4kdp3QfpJzioHImVIgeVyJMm3qKY63XqrKQzANn7rhZpHDON98X9P2m
/SZyM/G7h7Cqxcwbm3J6Xh8MJTBrpDJZK11XZGSq+nTrZ5qt6tVVeh64q6SZm/jF
ElagrMpeckQdPiWiUYT2KABuuhIHbMfLn1kT6gMFaOf3FVLYVPsC3xivRTgkgdyC
I4qPNCezX6pw2S0v+VqmHmjMMJMzwtoHN0he4GyCVtpBxi2llr6Sd1T3LQbTUpcD
zQrSyHKCWrihHAy5zNhKIIcCMqOOPU/ice2lTGKF9llgjZc3rtSykGJcp6sk53w3
NOsb2u+poH/1aAEyqzv8gF6zOKtZntsxpfdc/06GgruTO1A3QOmegnB4JCXR6Qlt
rGyO26AASx9BYgd74j8MdYKu0Jdd5kBnEGS/ifbTDJ8zkv68px7yVkfM+5w3COC0
lVSd2MncQRrDwTvyQdHBx9s8u/QkCllZn5Q4Cji+OpNCZfowAku7jNIq9ufPGDmO
L4bSWggalxRUoJnG9nCU12FMDHK8zpec8i7npZlt+D+brFEjDdP54Th6duQ529Gr
UoTl29O69NT6azO9jS+Ibdb8snZ2oIaeFtgYh0HSAvkwha87g+jzy+WshG6cW60e
EQVHi9gs+m+5s8+Xolrsv4fccgNCAO0tFbmswGrtbCk7nSRhUjAWe96vlXeXsDuZ
qX9RaVhfupW3tmqDw6t9ikYEaa/Gv1WED7fg1wEV+MZNBRScMO3LZAEYXSGF2uaP
shtKdnM4rkfTtTIyUqV6gPUry0FnoNyymfVPPDFRIDfde+lgmr4+WXbAWUV3k3/s
O4mIczO/aWR2kDvpghj7f8Fd8aJOmBP5VahhR32dhKvfOX5ehrCT0azBb3+B8Z+J
mxmKeWJD9fOj/amDmmLUj0yW0AGswmvgevX86mOVK3efsZGBFwTjF4s066KlJFVa
nZhGwW8Mq10g2Jsi37zlYmAphfDlAKd01kx6haR3E+nyMiJiXhKpRH8QlJuZ+TtD
L3t3sZU6sKKFTdyvmvwfyXCekllEhUqGlpdXAjKfjy9f7gh3xa8Hsv4r50LbK1GS
pXlBY417uAZ9vFnG1WGfYKYCopXhpIDUve5sHYPpjMmx6HnL9wBCObwLfXr5jT8f
VgEaAcQlqAixkfQY8mHRX0cDRbvWgalFxwjUCTyEr5/LJjmS49lv5c8JA/W92MB+
LRmZDaxrP4hZBJLt/UYLwcasf7p6CZ/kFaIAgyBUsYmxpgNqwVV8F+rwK4HCuPQ+
D4PuKZg7Jkyzuor0geuv9B7qsYuodFDYChqrEKp1F3vhhClQB6QWzZ/o01MPsVqE
mn1WM2J3WDTQx2WSCUmZae9PWnnnB2/lSMG7mkeFLdJ8K5crYNu40bj8U+krfCqR
9atSs0K9XaJogL8oFy/x7rMXutD1O2HYoFZ3lJ55MoqfOhHrLvgOA5BFkyCBf+FT
5UUTj+g2XjZi2HMCy3gIb+GvpVsmVjXap1l3Cz7EbZpv9GWyvZJ7FVlOiWaa+UrZ
M9wrMoO5eUBIHn+VW1JDmGlsd+sAD672+Y8FCtXdLV0VkiJb10s6SEIF7y3ILlLM
35S8n6fLrYVWmQ7I2Z1ptPFjOj0pNvK0t76PBmFlppHk0l9W9h6tZx0iUr0s8F1k
49IcE/P7itCC9nUSbF2Ynnbw+wRGi3b6SI7JXVHQE/e2NLfD8xH9fidhlwdQQsNn
1zUwUocVp5Pq5yGb5baLrzIn7IPEAl0+NbT2K/91wB22AHqcVmDF/EsE5oXQPOEC
aAM8ilRlSQYvglUw9P8zKv7mqMrDcIuylJrOc86Bx7GWFzWn7pLzROZg/JR+yPpJ
DvTuX7vHUFuMw8e47mSIHU+67jABxVwyffvxxboeCQXC+ubrMjwWQLeW6LxCgmDf
MhEU7kuc3W1hC2GUhsgrGl+WJ627Jl2xAZgQYYUJYCWlC25IJHb6cW2S+5Z6gdg9
aPdK+56/fMT0lVWzPC+wZYlRTAGWqfrOperrycMZRu/npHe5mvWRlagYJZWJi3oW
9hDfNTlkojX1oxtEZVWQ8QVnvCKIVXxvKJsbktzObfPdtNzH27QGlgy7j+b1u3Zl
CVAf+Gx4/bWuVLvipV8uDrYw3mZcewx+oWH6Q1JKJsDbVm+CPgvGST0vBkO9ZjML
Lxo0wHK2rUDHkT7tL7wqExwHVMmWVl9avgWuIdj/wXq6UBNyDAhLEqAi5V60xuJU
qNDBJZzD2DwbCcyshhuJAroH1KGmFQ52llxSQo2o+3qYx3ZBrSx8SECUh5bMus7M
/b7urNGEsh/dFka2BZprGqpwBa4V9fFHI51sxeV6dZ/GafYY2ouBV80JZ6I4AB20
+S2VmpqTKn8HZ8md8um2aSgmeqUji5+gd2XjJxmkhtM57gxMaYOXxiKF5yjUFcQ8
f5+8yYbFXSZcyZJBhkmMbymwpPisGdmUp+I5xX+NZcblgGE/y/ECUa3APb+fWWNu
oaOcXAMTe2MNRPa2/fkLO48BaaHv8sC87fwcNPceh0JvKlgyQ4CkZ2wzPic5UnxG
obJUgEcAfREOwH/6yH6u7b+y08mrSwx/UcnfrUfYNJ4nu6ZRfPMLwfPb5qkQ6WA4
d9ulzBVqjVURg+6H6FwDUQiMxNqTjt86pkvaxy0llQd3CcrqCSbaBlJj50+eqgHn
v3DPmqWjf8QzTj7XJrGFzdJNhB2sx4W++96fTOY5EXu/fPDW5v0ouyB8Ndbj6ezr
UWnNEJUNw4gc+/odAUWvfHV8kVn1vIvP5k/CmQOJIgyaW4XeOm6KrnOkN0JChNhk
q1K6ofSdfftWDobIaG9CgXv29wTVn9fJj+gXg/MRguijDIU4zpgUnbfSDInebOh1
GWMXE+7FNFB6uLNZVcQ4B2qkEZaLcI8RiMmfSKz3hCqv8qNkkHdOFguZ3ABHIahI
jdID205FEm3KSAlXBktQYRw3X7X2rWDrbR7ExrMkbF5V3HwwtcAfqtTh8mm7pZGc
v6P+2UKV+QJzOybvNcMWc6UiNnsFF7B6MvBgYaKClaktic6LkMumJdtFkapJ/LkX
NrntyElB5Bw22O+xauX/WDfvQFrrs9fjqEUL5URkPYpluRZUW/Zp5xtXWIGdHO/X
fZ0CW5H4vpzLqbIzQ0eZ+6cs39DWHINNygGjbN7hfc4oDLPckq6OLV/Aj3QdAFA+
D/G0+lv/mXBtwZ5wLL0yVaVC65byg/rH3tws8QfgRZ89zODaxpTMAdcrM7GB+fHW
irngHgMlzU4ap6RFI5j07stmAAtEgp5aVh8WmPuZ90SDnsPw7whKwDxpImK97hiI
VL5ER74B/vXLMTqxAA0AISDyvN7RKxNNP2rATI6smbI16iO6N4Kgu9z2yUjsDewY
GFy9rei/q7RpKA3a90d7ruxP1NMem1/cp1Oo13VydsBQRikGudQdboeVbWaUaOzZ
2HdT7Uv3wH9Qq0sdRHWFQBBoBxAIeOxA1pL/OzPPPLjX0GmpJVq3XEhf/Q0a6xWw
NvfNVlXo+ymaS+0JKp/Z5UtyWm8ne2cX0mToXUKLSVqpZA5h/a9UC7mOxL20N0ZC
pY55i3MnKMXxubOM+ZIGmBr8jwJPo1DbNAPyE+zRcb1JaphPG13VsIosJPR4p6J0
7dxuF3mxM8C4mqOj2BgpqBcGGhu7m+6jfSQFZU+NVIOMAkNG09c7VuuAnoRQjurs
xLoHIey1Eld7pgT5PfCjENeNhzngF6p6SjM/YklPt0gVrr23XzNUMaE0YeXxGuHg
8qvz+HQNYDYPbE5+IC4pt/FcZWxxOV4IpK/0Ul3lw8K+hiJ53RI2yJAI0bakxG+X
CcKeNnC3oqJYp4/kvzocBEut1HWfKA2Z9Idt8yQsLY2x8rPainogcw5L+fPk4NQu
bVJsG9TEmXpYauxVVaeaf49rpeOsvnC5K8tvArtTwvrWzRUu/lC2FxDIUwW+hBAz
eNgFc+tA8RY83ivE1JLEZENaz84ardjBomwGjyZ45RBQTBM8djWoI5XeIjP3dB8J
9Bhwtj0QtUdtsSV2ZeTm+VA+uJvhpJCDgCMIvYEPDfAvUB9vOngmy8kHekia6zyf
1aX9n9wAMEiP7cRT9sxUqyYENQJVFg+n1Y1T82SDuVaGUodJFS7zRZM+5T/JXRZJ
d3/DkkcOmO4YYPCC1dB816rPusfTJB7c2kcEhZUqZFc2LhXLhuHTwzWhblUNpdPk
5ALhfuEelTejAJJSsDk/y3ut+HVeS98dJM0Vtwno7taSbUkMtD5nZwNEg+eAwcsD
jAfMftratNszky09sU+MvhV8pLofIbfq66fVVwDZJXN7fBVihvlDAmx9RuJeZYnk
CCHC8X5zWWfiCMz4TYoEa3r/Z1i9gfnzD12Wosl41TFvM3I44W99+uOABNrkxek+
PHOojmMwIPucFDicgx6FitSyj7Qs1gyumqF6qHcpD4Ek62i0jNBxJKHwEru1T385
V0E+DbGB1K4v1Qjaf1JXP7izfhnRUXWJ3cnEiLJIrsh0Hip8vlhMvELLp8Ba/aD4
Yula4/XBivUHHhAc+kKX2B2lIOzlglCEcl0l5U7JwRJBvLWNMC+fWAbIK0JFgJC8
tVmAfR2yMywtllCgJDDuI1XQsdoiA4GHVdbNBpqqkhnqldU8CoB5IsE52qURAQb7
eaGM3ZV6JWtSuvdPPWTDh+iwyuuXb7CTq0FU58tuF3618j54xdj9vv+HMfcvcWvp
KZHutCHP+/nHut5JxnAWeYxO24aVRYeax9W2N0UCn8KGNHBUnDgCoLKeW3LvCSnM
hu7OV6Y6YuFGt4u6KN1Ag+Cdp1RSViJdzQO9V7rhp8LTJPmODzPnimjACe4H7NMa
kT9gT3+lZN5zS9ztk6GC4ja3i4f7XnyewxGDuopDZ3fSGdOq6N9b+MktMaRe9Elv
8U9jVLXakba+iFzq6m3u6WRpHo5WsvdLdVLKlGy6j3JnMfKYhaWkHN3xs+nVkSTU
i3jiXsXkTbVYRzYgYj1Uf/hB2Dianve3QcJ1KJEr4nWf6twX9dx7+RWk3l3nRRcI
VqzZUmqLmViSPjuCxci7eWdqWj/I98SRv0hunk3nc3xl1hr/6FL1FulXfoMftzNZ
0j1n9eI1VZWptuwXZgyPG14EGZOCzYbxvFe7kUM4NQxHgsM85+jFD4ddQJkKsb5d
YPzOz0QtS7D9AEYDLJqPivG53FWpovH/zaZK4DOsgfdtuDwpGpi0uUqf/fVZICTX
bHGFkMcz9S/tHFEiQWtywPcSYwntTjtfMM3ibF0UPlIl18T27PdcYvjtiNDG1Wuk
XXNIYRca8K+TtTrWRs+DzJ/oTGJf8Me2YFdawGVjacYbW0fzdiJs/bYNM0SsMYpA
bOR1d5/Sp4uxKobPsSwYBXCW6OFtieFZJfFbEb8t9dNYqTEI5To691NdfI2VwtAx
N3tgRDfFtVSaiK4cAAq/NmqMRZEdmZaxctCx+udVKXE2Pc7HYIGHVfquOnMhLk+J
nuoDhNFbis2C/yG/kqeqW1CypVbNjJGyOvSibj9xLs2zUxQENfDmPgAWnfTLCmuV
7S8MnTXF1R6IhE/Gfx7NLbpmb9oftlgGqMG+gtvw/Q1nEafrgmOZF7QLWYyigAo2
74m4rDxrRGCLKAHujMlM4BTKmR+MCmWxpb5r7cplrmxDSH++8B+4c/h/Q8jwW14H
Q5WjVx+ojPC7/9k5Znh68X0NCktQn89/+TA6cn1lSqjcIi2VxtzKCvFiuje8rN88
IqqlDzrRBRlkDA63/eqOaIRtua8+Xh7tGAOsl31xuYfgA0qn5KHrQx1lxE2K9kxB
v9BYf/SxhZOj5PrPpbzG5OBRzRRdzROIDV235yht+HEEDiQgL/24qtCNpNqRZ+Mc
iaMoTTUhGPMIYzo0HOOdaHLnN8B7QxC/ZWSx7ehn121hCSFCSM5ljnxY1h1rnRhY
8cINuAiCmpPdOgo/vK0Pn+XQuB3zKsKKS6xmgNOVxbOONdArErBS1ZyF3NOumXMK
5/GkkNQx0yzlq9polpl9NxY5N9CaJ0LdEJsy2ex4MYvJE8MdH0T1SlNMqPHAnAbk
UzxralHFfCyhiAPrmyW9JJoFwMyGJ/MjsqWj6AcOMecW7fNhkGlN9iOHtrmrjk0e
JgV/JaxiRU4O4In5h/ZsSwUfqdRIXbJyM96zFJCYN4NZgeI+Pu6h/pIhDrbgIysO
F+MIDuKJaNX8e/cyu8APNP6SasNLsSBMq70Ntfae/ebF++RC6Jqjj+kz1o6OgE5q
qwtW/oHv0LDfH1cH7SlafzP3o6ffaXtL83zaSZuX/XrwrS79bMWsY3u3n55bPQeW
QSVmOR/AeO0kuYitwp4csh4BTb5KOpZTDsba03yYdOsSI9u3X6ODZI5M46/CXX+V
Zt4OdEDbsWLgIRhC5KxILEGikqjQ46VGxI7el1ARObMtqVh14QO8ICjeDN/KMKzs
ecfSiYHEZdkJJHm3R+O3/UwJylTUvFwnhiOcYV7XGd4wT8q6wci/jXkmFs3GSfpN
lYSTM0QNaOPzhWQsZtjsAd/AF02lO16GbNezKVzE2xGiHxeMAZAKFoHK0/1ZYfoH
DDYQA6/BAgl31ONyp8aKP3lOCXYdTMU0brAxLqYriMRz8G4q7h0+HejBgukdeJvv
ovoSdtkjPu5+iBNMzbwagbvSIXglMt1tC4u9VOQ4cOpChCoaGsSH1xubyUCuOmJ0
UZTo+AaeYtBEb1S7JW5tpPOkweDjRvFE0O566atw4eq1GEyf5e3LRfgkbz3ThqWl
T9zUoO2+WBIch0JuNUp/A6c4CrMsgCXK/xTDF/P3UeyPxO58fOPeN8JEFIIzhNSR
TpmlNp3/YHWx3z/nb1VfcYsuxRC4iL05gBGK63DtbWS/GcaNpnnM44yvomWySnpU
ohMj3LSbNx3uT2ijmn3oRuxdmJ5FGhWJFHsL0wXM8Uc4HZ8jsJq0HX5u6U6wPruD
+J7GZwxfwHjt4eunpo+48zpoGBG+F8Np4yDLtKO/WrXBN+8pDKSL6cyO1h0wOkCU
kBz4nCRPJ+LY9qkV5/RHrow3r0A+71hJdjh7gWxXm/xCp5dbYTo2LJXWXYo6rfLD
dHOqTV6IVX0yGY4XDtxQPLytC07MQCQCl4trbZHZvSNnyaH3S9IviC/TLlcosgA5
2YwsWDxzeyXGdAelt2vnDO40/StvijHxaTUh19u6vMBNi2epeG5qyN31WVqlYwIn
JCKWYMNJWwR0pCepGSrXBudEdimjiJWW8RtGzJXk34599eawt7XprnZxfCh7RVN7
IToj15ro1YaAhGO0J0HuqX0CLeIb6BHw4Z24ybysuyvTfwS0epLCAlyMc44zotA5
m+32qJ84elcq/VWnwp+hm9H/h1EAuSa4wdXu6QTrt/1w4V4xPJ695rFLAhrxu3xB
ytyoflL4G3/lqnRZ+99xqIlPWLKfy8M4f2HpYVyyVpufiE7TKVUsIkfTi8nJTxUl
aymzZPBWHTFJpFb2TrHeGPqSTi1VvRzIIdIGMTG22TCXhCHjHAAUpdQPb8dtt3vQ
Iuqj00PGO484lNlMZbh09zrqRbbE8zmCIZhyeVkI5qJs1dxxkHLyFuVqeL+2/bAK
ZAeIFs06WeuRvmCPlise0/unGetM+VgdGgCY3nEaD5VZXbsVe1PvUvFE6XmusHyx
LkfFxoDKMFiwFQLkQIOkAFShq/San96s4gap99T2MbGrHNvoC2uflp0LK1UO+Qb5
goZ/IYvOTZ9dM7eklxmV/y94REUdFdUUNzDqKQefRdG58DpqcGiVAK5isLzCkb1d
kx6NQL0Ddttvzh7rjBROB1cmKKLwAPcbu4QvSWOqxDCym0SsW4/NxhkW0Y7J8Vzi
Fg6Kw8bX+X/azjEu+hxbn0Tjsg1o+7GhTw8ZsZgQJN1cfLVHXlHJHY0WDSVioPpf
CjmiPf3qJJsKOr8yiD6rk1+OpQxJbaMtr2GZq38te4bwf8QHaavZ+PfCsbOb+D4k
ktmCUPZz4NqYDTLW3fyT7Af4uop+vbN4IZrZSCgWSnCQ8OM+kOFB78KNVj0KhJBB
YehBB1GPqQ5cCt4b9DRrIWZI9HVq4TaiEg8ydCSM14WxuH9qk4q+v4G01lBenjTf
m/SEDbIEoR6qwrKximWnJZPDWrtCtE2B3ynYD5hef1lxvSoCf4CoVIN8V/WU6joY
gxFrtXRTzdoCStpNX/UlLj9686S7Ks9VzRpkroGa4s/nlrdI8JWni1dCkCLvjt9x
Lh2ySxLmBocJ1KdrPmF5am06suuBdmkhS/Q+yHf6/WwgGcVEQ5KS764JE4gKf/uZ
US4OyAHKufJf7oGSpKtV4gIyCnkSM2UdfWpfo4xsEsGxeXrLyL2/yOF6MEBtQSoc
Q1JZFSDTQDzB5hcbpCCM1QwgIvYp47D2bbwC63Tb9s7aLRcksXWiHbDQj5x55GPP
6KcrPqPDPgbCdQA9I3s4wx0QEZX1UDfld0Ic3i/B6jYBgWzHw9ZVkRnpJlx31ciw
n1LkdKO3mAVH3kbbGqphX01fMZe+JKqJhEPeQx8PrxzqHAMabOWyCusOgbgdrz7x
MmHC1B5cOBUIj4WI05LEty9qKCDz4Sgz2xqnjzLT7Pzqa8tLQj1YD53Zqg8RQaGH
KWdRbnXZhgc6t1Vwia3iuxpzQNL+3bsuoibvgIG0OZVU5Z61XEOFMdUeddTU2D7F
L+MvirZmT2hRU46fzdF5di1FwbZ6N0LSJ361KFGujUBz8mSJBxdFH8Ur5cMZG/BY
/mx012YFjd70esWcqQSwHboOAy5rAmeX8VMSt98CuPgt1Znw/BGfxdx9d8uIcmFx
OIwReX8WuZJ8xKdPmGuunm4YqKP12MEOLyMu3djkUILj1NsvPhI2oira+u9uKnJx
byS4098zGUNN36ZVUEVZ/ftqvF5AvRRUdgVPJzmOAtVsO7lmAYWtVrQDXOhrL+cv
UsAbeUwT81ke/kt5up2DefvOcj45DafNsCJ+0Vz1Bo8Bts5dcERD8GujleuVMg7P
6VLuONry+iKxDpCcR0noGeDTEhbsoN7t8iwkt8GuN6gVfFSAeMFRZ9++3tW6pr8M
W8Nv9ACsSw2dsm73QUcfH3/Y2hUrE237rTsWtldkQ0HeUgZwuq96blaxz3hEirQJ
VX/yHlirGgabnH1MQzbLmJJE++9JnEZ278tzW8RNGFKvk5VK5KxWyTxbEM22P5fa
xKlfnaC+z6pW3O+3wvlPDQSVZ5XJHrjpwfL5QHyX/JLyYpnZcXKOF88RmvwJ4que
NBLsMCilPdeQ0iUppmzlxJbVp0iuYlEKSsC+bF8XqoOIV1FK3N6RGD75/Wg1ymbW
+BT+iTr05x4H8XOKDxAM48idRoPsCzN+FqCxqa2xtTqAAlXsL1aG3DfdafwWrFkg
dmLGlb5Br5O565tT5yt5hzQqdxXCKOo3VpidBqKbGgTtlj/skXrCQ+IqP/dJWhje
O1iQMvvmS4VhhsJzsN4pkZsTs0RLTYPU3M7Xj1e+Cd5a444M5CjD5ko6KErL9113
pVEAcQVX7p6jXMq4P+gaTKklHvqW23FewfbnOPJYllbOzoAu4Ul0hTnXr6YSt0dN
5A7yTRQtoMd+Rtkm+OXYco3vEPJqNNpcOfDmwK8vELLrFrmBYrgyFt2OE8TypRK4
W0daZ0wU0FIMTFDTWL+FABieCbCURfk99wI5byhCZxTh93WAf7medsFdRGZE06Zg
7MaOX6UulNJ9wEm5Unp94mBxHgXgmt4LqjmKklm4TkQa1px3r6LBlfzpKOpSpLhi
kSsUE6DdIxOdHZ6pDgdG0lfQg/nVhtas524csazRLU++ce39HBhl9qIWSx2Fiplb
EPQ/NfO+OlMLe8P1bWA6gPOyh28fOhz3eNYO/awSGG3MEE2K8F0hIbWEyk3ff3LP
gcRZ25RjJ56+4F7H+NXc+R41npQ1w2RFWM9m8+F4OBwz8RFPVoAxLTa8qEakCxNS
ig+an9qkZH/qWHaWrTTTNKQfOXn/3+DcsJG+IkKeaG6/s8sgPrurbpnG0NwqENpd
6l6fr9K/BPN0SJGZbz1prqi9LnXgcI8W/iqhmgVi8bMrtGtjIHpcKImo1yZWj9DK
qo6ow2/RO3mcRvL7983vCdDbzbzzlj2MlASqe5+5BzUvwwptFCf2Tf5bu9HLFFV+
bqlCM5uBAlcPX7bAVKJkoX1CBv3MnC1pKSfqwTSkcObxTqFKTDUfDPwf2Hx2/j1Z
49U4SWny3oxWxCT9KaIvCwg5z2nbPV+3pVCYxDqDS+PetulyHAAamqm4R5n1HeZM
1C3xtrWgJ6YA1whkqCjw8/5na3P0sJ1nZ9CvvmUarBEHZdn21zJ1B4zEQXVcJkKK
NwETT10rZrjkhwMMV9rUdHaZluKFJLXnPMIgYnjmbl180CULvQVc43sZ3uQkEAhr
4oVL+AIP9p7LLk7soy1tdMDfK6RzrKEXsEH+eoLgurLFad2LfZWcP5/K4ANW2CPZ
tZZixR591u56ur4okjGq2m3LDB9TN6Go3BXul8eqRatX3D4meW6I5Aqoe5lyJ4NA
MqwQ9xhJHvzi/xcXjGTU14idk84ZsuUVuPuImYFQcR8EEMdM71x+ih/1JkrMGYi+
D7MFvuZm4P8KxzVuhdX/G3yrx+ogyXGxdX7TQe7ACVedKXCumZfRhOA6wFobXV3Q
rtBkQDMTQf3RKkzrHeEpFDZ7dsAvMyjxvVB694RBfuIGxAd4wCUHAV3qFv2Yaj5a
BfsrdL/rIO0g2DBo02sLCcn6IUWEpYb3PawA8huLwlN/giLkYf+7vsd2Skyfr/AG
ZQRBzPVMzZ1Z2YcQYvZagg8r5o60KIVcsXaBBd4DE6YjbvzpdRLWqhXIIFaI+e60
4cDBmmUqrev8Rdu6KpV0kXHio8ZfyhNIIqWNoSkBleXv8XANMPIAsLQXvwsGSqFI
Vgir+iZHfulxkWuhFxwGdBFCQwD6LaoUOObAMLTtXN6Y3TtTD5StPZSwTjMcTHB2
9nmLBHkZYNkbCqlsTMpu0UzoykBBPx8RVlCXJcVAhfAIlGJkm29Dcv9BcbmuKsea
mmJFCBMGIWJN0GWyAynRdHf3SH8Y24hQMC3qCaDB4JSVHeF7IS0XAp91BbAmI75S
F/DcBMRD8PH9GR1Gmo5ApggwBPwLLDvTg4NPL76hbgEefVq7Jj8Nm+3ShK432VTP
iErVGmT34XPXXJMGK3AxDMvSTZYNdOpWcJ5M2x4Mz3iBYdW64IyoBlDTT6VKMUIO
M30AnHgeWObBJLquRiMyUDfTL2r17wolezvTku5wGXA7xmOYUrufUIrCB5ZRRRf7
p16Bj4TDpQ2oJtdREhZY2CtlRyTJlOOwJ968Y6fRjZZTbvZOKH51SDxWtEHeb8kS
pYTSCvIYpH+9SD7RiOcaEw2MrHKXN4epnW7J/uOhd+cHeLR8z8OgdUk8ZFDW6LsY
sqZfJle6q3fZNFnRpTWyVJ4haYvSTZ6opR2PGRbG+daEYnSsMkpFe5I13vnEtURQ
cRqELy1oPgv6m32BExJ50PoVhtqV/YYn98I879QWazZ/yY6wBDkxfFa0sL7rvtFE
5JEhr3fTIIpAiO+OMMxg/hnrWKhnkaxDDHrHEOKJVaea8/qBsGhuaGuaX7OZ5C29
cmmfKhxNayFHSlkkUKaijZjpxGCuSdt4rgGzjEV4/L4Ws0Jp/XtwIgXmNfTzN8yH
/PeLNZLEca94mEKbjwrlyhGAXodBi9NHH4m3dJpo5dyXBm3mhLCPpaFD2gxwwbjN
YIIaVM5wNySlAcKcEaW6rdPpsy7VucCvFw73o2DPZR1TKZuXwvQwtP/uD3m3TVOn
5KMhIN7CEZFxzKQr7lkyVpPw7ZY8zf+3qw2Pl/EFHNL+6jnQGvLbTUtnanzW+DWa
f/cPJwhASdW01yPi8nlUnnXdE1PeKu+cH7+s03vmrUtzG141t80jLFRBaIuoKvdF
OmAanaZ//sSzUE/pyQ4ofuiZvdYqfVdCHHZbpS/ZPu5AtLHPUI0dLNiO/T00rbDD
rllxQcvhwS5HASEDHmqS7huwbRBMNPGpC09HTHj4LEl1QApZyItcRUNWjM0IuBfe
pmkYLEhJGJ+8NBUfVbObxci1fxmL9DwgFGe/1gYrZEbIHiJh8DYXIj+SU3/qRIsp
HOAH+cZQuUPO7nu361i9c/QH7Ny1cey9FXXdXUBNjQRuj1GCJ2xZCWt67zxESynG
J+sNhUm5toqSQonnoKQ8S6Ns5aRxoRwmUteE1gg/cNaCx3Jl2+Mgt1JCMbhH0LiO
Xu8IWCrFJhiBpOTmhLFSUyhZ7AJRS6Q6j/O+Lq4yxwHWTfRhIZds6i5y8UBc7msu
9WGBRSEqe/yxnz6ByZA5A79amfJHcxaf39Og3zMpvddOIKFJaubyHXP4mlIyz9Pu
dFD24EYmKl5ZpyVTym+d0l4m2cFAXhuJbZ+MhHlrK3PZ8oDGKuCdXnqe2nkcqyO7
IJDRMc61yXoyQty4Qj+lgwpnl9N4cm1/EzOuf+qTf0joh9rMZfIuYBGKGcEe6wZU
CEKBjPIEI0LdtSt+JrItLssZhzoumCy9CaeAP99Sn4hcIkmAw81F702sqvoinFIm
qeMUgTbCGdLtCFVYrtPq3rE61mKlPcG5pTlwLxVsWUf/rICzqTWTCJC25N0od6hc
uDfMOijyimv2b8APkIQ0qz9hY6xuMNgITqw2csEnBHtrHoi6qiOu3uCgJsJ3hkc6
zHqp5t6K0PifZKQWniQCANaYB5ky4+CBFxrBcyUJmeasTi2x0dtXwVFGvKeNT7vc
0SUtq9vA2n5kfDZpa9iKX3BRQHbyogI8P2X5UTkpS0g9+UjQm6hgwZLdAXWsV3yh
DOm8UX+S44l0vku0JWnk8Qrvs5fxmuLH+hrZ9K38sbskKivxKvStTLcfq+TiCufQ
5Ys7VFWQS16tInvy7Js5R34dV6thzRPC4UeitnF4ZQtSoZCYJSIsWe8eXMocD3Tb
RWnoYNGcbCturr5lTE8+HMHM/GwbwoqS+ElIX2WVrGg2+Cs7mO6JraHMvckqWNmz
iqTWNUe/KOWhfVgjnN9Ug5zPXyyOX+czP2IPWGJ4iEM+qXCZD5GD7CvJUBPwxJ6w
U2KxVDMDM9PvW6u6XFwPSmMHQ3s9ykiX6aw1HbWVo70eG1r/clPOOKzQH/9dpW1r
flFY72OlDtXZ6i5SGmeFwDz2D4yj2NhxKmWf5jEWmaAiQXPxFz5l/Y1bEIEpuERQ
PJcjgReklhXlNO1QfJhc5HJgQLjk9JsRdE46llt2Xj0SrOElxMnf7Lfw+Dw0Kh15
7bPdhE7mJigoIoSRE2FGs8aWjeWiKyoquSNb/hfBUzMmafUtygEpFDxdv0vFGhku
4gqbGwvb0MbuV9hDW/3H+WAZYnkki1Lt/9ZJOL8LpX1lO6y+eDDMxQu7XklJdMeg
mSF1pnefZgplHV1jj6lNFix3u4A7BlSUqo7PS3FH0fiYZNMtqsKxW8mp1T6BnwA4
vuezIcgfkGIWxA73caCYH8LV9JBBwA3Fj4nNc/d1M9pKvFL3CzvkE0KyGaCUbFxU
W04ELcMYc2PviK56VMAm7zf9C5f6c2kGOnxxPH6p4ro+7kH9AGIdQDaRhlXLTGfH
KupAtEOheMhNUYQ+J/nDqyeGUyKJ7GMTT6EmdH1CKB7MTXCrCiY/Kqb476HYa2dz
XWCEd0oQ1j6esju0lU0HbjmPtD+Im/jfFP5UJrUChr2vdev7sLGeotis1rxxkQMs
jNCkHLym5i3MZrtT5tqMY2i2rDgvxQxRaQy/ZlVXoiUzLt0AxXpYc/qERuerGvuP
5ea6Ow3wnW9ahd+feu0ALWK+qAA7F5WnbiMXni+2GIEFN+rRdf7QWhLf1zfmymgq
Io6aTzJ+3vNJXwcTDZ/510u/w4JTcaC6r11/Zbvtmw/WZqcRToa7QTTvjs1Bf4j2
i5A+YPnriinc2xn9VAjPtxix7PwvaSwEfrOreONUT+898qFfrtXk3HcHuIObv+Va
ouO8uzFh1kasxBfvSTkzbBf1hlQHAWUXSBxYhUoWqv8xNdliIvztdsc5QwSXeNGJ
ocKAUtWvLcOz8V5W+mewS9SW0ILQ/EEy5kSfTWLpZbavdrw3+2wloC8y9Z2+k/UO
RtBeLWq6vRwVG8/wMFR/79kQR3Ro+xJzD7lRpb3tHgYM4zVScIM4aSsxDipRJSSD
2Zl83qIC6R3km1Yauu/UwH/oX8buiBZaNWZJdVF+u1YHj1jHB0K19ghK9P2PR6aX
C5RRukac3TZe9V5UlEjeMgGD/bqZMjMEO5BEsyJ1tVBOn4FAqwXqliBD9bGNLNwP
ZndOy8q25UU476Z5cElFrNXB9oPdDpTXA79cOZcOotpgLiCQbfRRhrGc06relyd+
yW3bKampxe3ngi6WzeCk27R5g04bSUyGMNnioFXnhMGwWb6xBJPKlBl5IVYIrm6r
Ukputg/0B27H5yZ2KYoiaYLgk1XFVrhCRc9FJH3H3+EFn3VcL99oFiW7DJFXpOMK
a8o8q1Xi+0skvTQLOhRS98+qcbgdhMJ4oOoNahLqWeKdibM5Pr0Yd1kfQduFYjgE
EnwixE0B5MVxPkzP6r0Sc3ZIWA0P7ueLro/3fRXSNMdQD6u8b3cKCI2N2WVPcmmX
QIAyyGQIRvUpIH4qMNHQsNlMqCUBgbllVdcn3C7AvHo/0JuvsKzWRL1yhfkomAug
GtlnvcDfhjew27k0kQ6Jcq6k1OLYAsn3o+MYWE3uPcRh55Fu+02r3uAB1JimYZcI
BepKRaLCT/rPkviv5olzlHHD4C7cuG8kzXaBxgpQ5Vg/6ghsPlcBQhkbD4zoo31i
c9/1c0XLoQo8xDJOc4wTc8K68IKlez73YBZ1Tf8s6ImyZvHxRHmSJUJUPdYTQeu5
96roiwc5mAm+FywD5UNM9+sgj93CRaRqPxCwYWKDYrlZW0EhDFyZB6TxHLdK1JSn
jq1rvUcXZd9K3852HDcgIDgd7PWzgnQYbMgit5Yvno8WOTiHd79J0mHABqgy9Irh
EYefMZN6GXRZqDpctB82c9QCQxHMfnnS2d+BkUt4ZI7s+vBOFT7AtKkAUBFZbI6i
mrvx6YzNcxETyqu73YfIvj6sorSUc3ODRInjzP0NyBiS/KaAxhJ+wZ1xbQsWpf3l
zjrjcY0WGii1WoE6UOLsGHOKTax3dHZQUD0xPKK0Gso9WJAzlHiiKExS2PdJRXw/
8HQ4LUMaoWyrnX5MTY/F9yzpWh78yD4hGJn1z8mAdYfr7rK4j9SVlrncBPHIWqgg
6RgMMSe8SOEJDOxzHFmfcWTiQ3bYLd7ZHJjx+VbE2ziogihaBVuEljVaLwOdU5CC
ZK82wi6KLsS7e7Veg0jmRfu/OqEVHXT4ASEwfpWWvAYEzwfm49wYYRqdziQzpnmI
1JF24PIutlRjfh6rSloeV8waqkCOOo54qW6vbLubh3Lr82N+Rsyc8f2xGHt7olUg
vtnhDqU/Pd5HXOefB6DnNTJgosYeGkr+S+61u2IMEoJc5vrxZz39hMntT9wCDHjh
rgtAo1SXVw1e9gyQDo5htMKExEgRzyqaebZh0DiP6RDzOd0XBeWI3bRs0yAIsonV
Ie2kOY0Slij6vveT5EQh+4W5Kwci09wEfqkl6MdU/3SOC/I11F68QX1MJ9K3pFy+
qIU0ae6EOIbMTqCNWA/jREk4DumKfX6N9kpozdtP8ryuac8kMwp+LrjC6YrGRCwt
2BKqFTyD//gxhV+Yxgqrbc3hfWukQrDbmN+TNHVbcWV2urTeqc/VceS6kXvlsJMb
pJ+DAoIoNkm3B4tnCs2cpjRYD/VSK7cbfC1+KXN4U9dAwqO6MBkhvnCdPDwRT0wH
pRW3LkjXTIayCPsQCis3c1tj3b5CQykdEx9CdDlGSb2xqUm1Q/gDwY9abpN7GKx6
0mTyQP7M8jaXBc92nJJWDGA2jVCdp1+dekcPcQaLKolupZEGeG4oJYkcKDhp2B6t
IUe8lZiABVQMDjMrBqsKeFacQutI7b9Xsm2N7yOaY7/1MKwWxKXBRhpEcUjvTfvL
8BFizbbKaw3JTU5WOGczi/wX6fyxiJrOtoRgMEnN1hzDdw0AFwBLh4bouYFb/Tjj
sXLaqIY6GWN7ocIQpUrMy+zC30YsqCkeTgZs2eO6YVvpHJEtJMAmK4yVg3kX1lL2
OdVq6hu+O43rvD95WPJYdAhQ+aoObqqjejwqtjhGVuQnACTzlMxI6Jy97YwRUUDv
7vmVshttWRjs6H0lllWBu4a0kS1+ho6/BmIYlAaTftWTKSVQQe0Mz8O4wa47ViZQ
fFdaZ2dj3zBE8A9mmGXhSNXsVGjfMtVW6r8BgM89JJO3NkT8cQxUcFfci9aOsh6n
xlaHDZKoagO6boE7SaKb/IdVfIFOV5oWoX9zDDSFY0fuDtOmGHHsSeOe6RQrSBKp
QsrJ+iwNsLv58sIFgYWyV0zQWAblbONP9UX5YDDuIp8F5h47aHkEY2Gbn2N63Svz
6kBIxCgLPZ4n4avrIBNeFFlj+l7cN+t2bY47dQE+9xECVbUb69kJ/ZU3bUULLsIv
Ye2omB69RHwycBeaA5oFuheO8h1962GsKS3k0SBjFLW5axG6crm+EalC9pTb9VT/
LzngZTc2f+LTFSQW5hCetjjYy2vDgJ3fQzYpzdJVAHeUISro8u8vOgg5VyELZ5X3
o0W+yCROKNE0gLyLYBDThed38982PH2WDOpRjE+n6a1ukAmwuUez+vWBbsCFn4V1
jLxFlL+qpPfHCje6TP4cEF7x5+8CKvJycECxAdaORKKyuZYWbtMbamhFkXKmPD2X
cKDFYEwG4KHrwBWXdxjldladTqHC8JORsTPwFCH8fTE62n74kpf5UgU4za1tNgBB
PYZDAgYdOMiBpyLniS063husnUOKq/y2V0AsNxZAbYAQk34ZymiTerpSf9RZkc4q
qz4WckEXOoE9r8bJj8zyL9R0c1bpDru7I9mmsUBVE9A0p3ZtSbvIYvcEAHHH0mHg
fOW2Noolq9fNcTGM59RPH+WN67Id+JpTPkPfPFRFiLRqoSpCTeUmxu4Kx2zwAuQS
BHDBXFX+536EXXjvstDWHGho8DQNWcMSrsk354mkvx4BHu6ZsGtk5xRdtcGDmqGw
iLVKMmWpoL89XEBHgkuRrX7TtH2sF8sNWoSzUeRh/kaAniupvzoyMe3hgy7EWS/x
BFT3GkFF5HIq1bt5jQb6N6OJPpEqWtlIID7iIx5mPlH4TCXHi4+Zcs554cBRSLqu
ieCNL0FHHJA3AQEARhpJGDBzZ9/eP3Ne3bd4JBDinZyqOq/A6NnUbalYc2rvSwKt
cZOUrNriKMRoajUxgveL2oq9SyGVsr8+iccezhrNY2GzGczYFounQleFslrrRfd+
iqFbv1+umsmGs7v4zx2DqqTZXgbiRXS2JfAX9hYzehq/XhtKvKkvdPit7T/+FGSM
d3xQEEvZEBJwjSEfQk85sBQb09rKPNkA8u9duqzpHka1n7/wWdpbTs0f1wLUrFHI
JA54Sv+9zwtwC9Eypd5+fsbGbiE1Y8loFvh+jb3KfhrRV1bwYQbUa8ZJ4R5cQnnV
JYRpYSVPV6TXWQH98Qzr74Y/jejLKKA7UGwkON3MzOAEp5SXZCdQwNG8FkoiogAX
BfRYGzClkkk1FVzyMN1Va7lqbxdHJfy1J3pChq5EiWIuf3rOHGVzJlRpX/o0/UME
sP/7f67DEN24h2ir/byt7T9HFdGGeUM7ByMK/NFeWQcytOJkzEUit8HaenEZ2455
bCV18rfBHO8wm0uojavp9kTIsp9T921VuIHgRqMLfZvIxTYqvC9fU5SROzAcvwcO
Y1mIGRJ2Wd3jMBDsg5l3Y+Cg5kZenbXZvMJhaTxjOKGC8RjwLNJrfwnG4JACsUqb
BqChF2B/G81HZ4xRlygfkwXuxKdflnDksc6OVZucwZJSyL37D7k67dE7o9l+d97Z
fEqmjzbdZfz8Yfa0GmIWd4x957r7/38WYuPa7OqQlXMoUz3iE5ZxPoCOELe4hATe
FEqxnZXpuvkxY8UwiOmNkcfXUf9v3upN12BjVBBVcbv5XoEmRfB+NlRHDHqONfVB
d+0r4TbUGN0rYj98g7fMmcFv+heGgDuCV+Vl9IgTKoDYzs5kx5wld2CkGCBCb8ju
TiEbvYBGG+9maxkhqncybQBpLuBEfF197UDiMl8i1Yt3lzxFDhanfEKKQj2GDAqL
gK9S9dX7amULNL2pRxqzdt6HlIhP66u3E3nLUW/+aYm2GYS0slTQKaaFI3/ZG0cw
xLx4RyojvR9YysFEQc2d4XJekPVfLpZNt4Uzk3lOpZS/uYN0lT6pDJB69lI6xgOu
V7ORGM3jtsZbBOaG0/LejhRnS5at/3Mf8IF1jly0xLsE2MGsxS57KTPQssoHwp1x
DBlwpFPTQZ3DzfMQwTy/aJgooay4lYjaH6JHr8x3OTF24tGAopzo1TK8boT0C+qm
mstOCw6DHr6UZaMVihzlIFXw42CS/GrEp3XsewF63vfYAtgL6s3BUeQ3qA6kS/a9
a1D3SxITpigR8yUXm/PggYkeuFqJdmoh06PJESrY/07byXfP+Rl9qc9cHxmQPQeK
yJRpQE6nqKEkABOGd3fSSvWuz38iQUeQ5NvkIVek7WkIxj3UlibVODMTjh6/b4FV
QvlVPY2sMOg96Mb8IomrislpPzrYJX9XRc8+NUwKB33xuIVJ3AmCaK9DzPvt5AFz
CZay4YTOtmFJeCCKjs5NAe6pBupXCwUQ3UWP0Za5Zxn888CIxvqil2QEXXdeGlCz
Bg5fAV4wNC6B/rl9WN7JHriIVZ6xL+NxfphcLXQpOvtgpjzQ4GerkCZpOL31NV4C
6uS+eX+/TLCQ9tvBqNYJD7bnFficGyADrmWo51W83cIadQ3C1+j5BbR/5vKiErxy
nLGM6L/g3L5Sr57TStr2SLbo4GmnW1vel5ZVWTFch4gdVo07K0HESIS0O1pLmnDn
XEbZAzVdC3rhPr1IrqQkbtfzfBGhQTnTAlq4u5A8ZdSoxtVAXnJUnxD/ByZ7gUs+
BcuXS6oiqHeeiChBm4fXtyBEQr78lMxSkQ7e2ha4YDOsugjLd3kLt8eyN8szI283
hS58XyQbBZ0Buv3Pr0d7MAdrZaxGsST9w/fGG7m3tbmjgXNNeCQd6O+IyWQ/pl8F
MjvKwzP+SxgI6XXeugXuvay7JRsMYVzG1l1GkH/3li1LmSE67Sr8w8GJYkUe7vur
XTd1XTmd6qiAyQpApiwYhpA2ALk6Kv5nebu4IYZ/Ak+HAGyb6vcyIdPVg/V/sZMa
yd3gsDlkQ9lF6KppqbAO/DypD6JuMT3lhE9I5x6KAbx+kvWwAPjuwTPc2zYdP7RH
MxvZewIZztD8cVNCA+94YbnvI/Pt9ipMF+9A8hhGHcb0US0sV+P6sOaxBUarEJm5
r94GHbAzeaQQc2fXb4siFDLt5+rZubdNFSJ7240OBm/fVvfLbAWciG8t11pL89Jz
a6ip2ES3vysvRJDVh0BiC1mGMm8nNPNzxsnjPk/R+Jj2/jSmNiUbU19W51Y0OkzL
YHqaAmbJDVe+9FXRbAvj+JWEbRCPibj0cEzhN2KCWU/wFf6vNHhjXxzRqrw3c8cN
Hpkgj+WfMzzQx5fniTV499QJX/8WnJv9vQplO4DJsDFN6Uh1cPp1CVpp5q0tjDpg
+WhLK7HH8LzhNfyl64YrSFXhlCvkjEcTQJrOGSQlAh9xFmY8PswMiOeXequlrnoR
ULKknYHL4E4v8I3bxUK4eM/U/o9fvyrjEaz+k767KF61ue2B8/glY8ibC2bRt1YU
RB98huOpE47LfgUUFq3PIN9PIutn6X76ATjaZkMtJH90BEJDcOM+GgIZ+AXMqJ1g
ONlMre+ftYhjcfgRZsqzLW423nr06mRk83RqSFOdegyAgo//N2S9G34x2dKU93WH
4KZMQ3/8GK13cj1tRsL8Tw0FCjoaKLhqThuYzH4NXHhc+5t2zfEXybRPeDy+QpG8
S0NJKBtP3QtZqN++FlqyWOU+XCpKL4pr86o07vCD2PvfjzgKOyqVoUTwt4rc36cJ
1qL7a5/i4ls/G0B5QwkZ5bfNr8Y2viubTitf8Cg2H2gbBzNgDxtm3GEgHZg+5+il
2ZEzBBsrmLBVRhbbpS1Zg9sgro1jTDRwncfB3cJYBV+TaxL+Y4lqaNA68f5k+mow
ryvO5nlckh4yAdDab70Uk28IXTdZkZYs3PDtS7sYomCRLy2l+AGtVsxSbovjJh77
be+rpXu4QZoMhjyy5d/WBgXCgYLrS8FOtOzHI8oL77LkwytYtiVUchAKD14Az35x
NAQhK4/MxEnxle4Qx9sK9nyoSa5dp1UJz0VZsprGmdJK4JyEE7DMcDmLrd9MX4W+
IGT2YweD06T8sgvAFcXuvBILhGgLV6P0iaaoOTmD7y6wo+BRDVVslMC/o6CPVhpf
9sOCqDYzN3ACp9f+70Wxlq7vosPY7QtkTRLFUb3322+k3Fsv6Fzlvm94ytppWG2g
VuNPWvGj45vTNMZORqgCdRk272F+RdfwLpdpl+hlZf+6DG71u4uU3gR7D+GE5M7+
JfbcCUGwrczCjXod3sqO0o5H4IsH/cTKe0sj3DbkQu/q4nFzJEIq61Uh89IRuK+1
TuJxYgIo8JdrGPp3hTx+fEqUt1ds/U+PFCkyBSA1tMhxf0Ku/UKmB+dHU0ErV2gc
E5A8Z/N/4Y5Ijyql1baLWWPnP7gP+MpK1JSiT5nAa6gwu38Or2tJ8MwNTJOT1ly9
lBkXxTGycC4+PMvVimwvEDwybjfzbSuGc4+5FvuTmwPiT/vbLixIMXxBcYWg16zl
viHQnNshkSxRFwPBmprt4aCSr5OkpKuCljp2ZS3tzJY2Nxq+2XrfjZ1LSQif2Dgi
bX5+nxLGn224P305gyLTqRWBMWR7grbh8oCCUtNE6yvtsxF9XHnfjf0gwMxOa2xx
HAE5/ucoluzr3AnBPdZNH8YthSxiM/aMr6v6ghNONpHgLRmySr4WL6sANXoLdr/5
rcL5eg3APTdJD5uQyqx19iRzZlyNzxcfw8UmCG9ZyJhr32vSz+aL8zxRWJKvHUu8
i9mGFYp0rOCMCqq/9D0Gi0nBR/QsJzHIV3Wqk+gZRj46GrkgjiLwJLJBxFS9FG7O
k5x9u9gOLRKRfgBmBzu/qT8tN6dNW3sDCGXu3S2Ai9JbqkYoO7zjXqaHpsZW35mm
QVBJN+tPxgJD2J310kmtPntJx90RxRrYk95tbn4FJ1QJYdo6uQ1u71Lyqc6IpSLu
F0fSoQu6MK0B/KugS+xl5UAXBu7aIyM5mq8o0bgvSBiwvtLyY0gqCIjrg70/FW72
bjUTCRTMgMAE63P4lb2DFox7X9hu1hQGLrc8lrqs3Ih4T6fiCFbDYSdSiC32EXIm
VR1cwdG6Jo7X8WIrvwicpgcKxskwCrWW8cQ/iDz1+5RePJIeB3Q5ifb4yON/bsfQ
jEWfCey07PrwIaEVuwU69blyuORpPdajcWdBI2ExnDjY7cSEKX6BHVvny22fn/AB
k0fX781dpHfnK5HBeiYTb9qpWhQltEThs8WNSF3BxaZYkG/rqQQWt6Rj18HUDXTN
hUeq1+iWL5C/qHDfA3JDk+yr+HwhOJEmXtPYUB+2ezi0uIyJOBYqt+APnd+LwYku
OKWfkfyvWcGUkPzwa6qw1Mzg4KJ9+/XocZ1030NgwwivCOe4BC0DgOy+KaibBwPg
fixiYUbSqmOqje4ZafSCxUHCu2G5HY4KXmFDcMNauhoQkLwuzNuXKIbhfRQXMU6a
awvbuev6sCmAOw4GM4gSkylSIXWTptSAj3bHTScnoCxAb379EHIum3FkXZUUIvxG
n5qjlNGBp3jbDer8mKr67TRPWSz0tGCxnx95NBx9JzYNhQ46FOqUu8zZxEBf6uCl
i7KGXR0TWGpFnboXsHqbWmQc6vWgT+ijg/Oxz/bVxDeUy7bn0uBaVdbq93BqXB6E
U1IkFLaGoXchLHG494z7fZRMayzB8g7HH8p2Jniz1T9qyGwMZL4SdYHqgkscs5dC
Vi6M1q0SR+HkVAbBEIoqAsULCRronhxl9s9lBvnszwX/HKCrlWOtE5M8dPps/B8l
OTMJadadfLh1JyBAb46326alklhHXtdT1yFlQfYSRay66qG7gjmdLUhG3DvQRlV3
ouXOJgvQZllnBTNDjb38U7xluipqJz6FSXRYGgr18BPVsj/kNSas7oCGuYA0LKsf
92D9xh2IE5+aDW6fHeXQRxQFCrjCV8buCPxs+dFHL81D733FIYbkmhsjx5Q3yJLo
B3lrhei3+XN3CRbZDM+3lFsdMrDF0QuKRjmyLqvOHcFhdTpaceT3ZqqDLzk8uQVd
vCUeDjZ9oQqoGQf9GzUP3vbLJO10kY4/7yLQrbQb51wbuVONEiumOY78jC+HiWN4
5/7zgxvTceAfO6KS+2Q5PMYp3ZY1DZMLqh/sSQk/gCfxVJQBVZJV6iIp5u62py5u
oZ2psuG1SeEst+LXqqZm220QdB5LxyeSMH0A5BrCot2581jPrSJvWEntwR+daapO
HjAsBBLRFt2BcFO694lMDFrFDKJUV8mtdZQ3hrXZU1J4UxHr4Zcv+RJtUPC1S9Wj
VpG1tdoe5EDz66OV5dCwE7EOs9Uk/f1j78aFBGE2rhkrJuVFPtuU868hqn7Ov7U5
tjd/C8I7SMIzQpBQl8DJuf4PI24dYZHl3org7z/BZXf+UhkjYxFlGC2lLoayimIB
lpIN/lLM6dlSVDPNzTr93mj10v6wR+Ln2mi94fJs+E/WHRcXYb13M0KRJXz/Uu7l
bThnJAEEE0zV3U0J3GAdcCv007oJMOKPSD2i5YwIeACTIjpNNz1331rpG6rSUfjY
kV5SiG8WCW/TklJMofNhpVOVd7jOkoDeJEfyoZ5hiFX251ZVE08QgCi6F76ZpQzD
Wp4zZegs8M+oPMydvTbUTYBQNemLY1Q9gmVzRPAF4oEdBUOPbFEypddTCdKMhHaW
I5DgKzMlXvzFgMjXgDmQUankJkvamyHDHr9EmE1blsOoqwwxUpEnF2l91kE0+76X
zOjW6BNjDk2jb0jTdPpx41qTpED8nOipV1Fur4H6G5QtrFi3PL5/4E2r4y957oDZ
5G6epR/jImPy4oQZ4FkGqHJEr9Ph+HDGPp8xZkbj/2SHdPaGcZ/jFl77KYq81BSM
C5BmVHQA4uoprDQmXqPEUwjN3VBV0bshx+tp6dPK3VCbyDDBTyoZfcOdjuAGoDKa
iu7tGlqRs+QcswOwwxfYuYZT6lRqJEBXOs3B14EioECyghMz2jHqAFpGeXRtgHsL
1BCfY9VGZivdq4FRlsSTmLWyfoEs12tz/jLV6VYEHdYCsXQ/n9j9NFIkM8Fi3cI2
YRdVRwS2MMJlGWq5VGZnqaBbfEVmqBAojMzIUavNt2kuKegPgYuWwDNCSxIW+l11
b0K0/tPDehOxp3fYxhf/Sh/ZtyU6Bl8/aiBzJI2NB/8rIPCXDsOpnT89MV51slVB
HPQSYipp1xDienRM5XU5tpiU3Z/sNMq0axA2mLiKJgQxAhc+Tgfu/SeP+uC25C/C
5MBRAIDAG1OCqlrWQ+6J/+xvQ7NhccJUoOZb3ZSN8OUUnCu6agWzOHxzlSTyPo8/
5JUlpVV58hUgqGKvUOq9P4ukZL4AQxtF9TKGIUGNx9Ujru25P+USvXKjVvhVPQg7
mnlxB5jh5tkhU16jQg39vp0lpmMLFfegIKoD5D0kWiO0nU1vEW9pwsBAmtt09/XM
GOyaVKZ6KggTsbuUkBiiXTe3PUTex1xBWAVzW64RPD5f6EnMz4FaUyZAn19MHHzw
z/s5/7l3URMlNBwpJ6of9LR5YBUfGQLpxLAhXBD9JnDgIipJsFQPvo3mUrJ4qNoI
Hj920KJlSXb6/3rjeUjMEkpUOb/s/08AV0qP1vuJ4Bqs9kgVCPQ68/H6j/ag6XX0
p5ieicYH3r0TzXQQB42JXAzM5ECEN7pYoNsLIFNk18rrVPQvxE1Tmrx/YAMe8NnK
UeHBBrAOtvfdTtcObVz+9hS/hwHU8g8bNtrU5JgR/V9idicX1DTnRmNhpLv/MBIE
EEP/Yfkoj6515y1Pg2HSCDd7riwJMPZvGvt2+HO1iq0yIAD1NQENGRaH0hDyToVT
OggFXhC4ACLIS2q6UhJgyGJr4yVjdkuDpx+v1qjdyEjTCpd+ysDg9DOsvlT8CGtv
01l1YtxSKSYiadA/7rhGPCAN/ibbPBhDc5NT9ApOuATI64qGZKkbMoHo/At9EGsl
AJubCRgCC8cevBFq1eKvTtTHom58Zq6Q7uAfsynKuN80NkdsWpPn4roctIRJ8etH
WI0eCyFPMd9KAizJtlaffBMOEEEJUvvDSshUHsfgssh6V97pKFAvARF2sfYOMIRv
wpbmZ7CHIt3rCtXc/MPWTgaxhGRESrF8CRWjYSJlEAmOQnKgbLGil3Ru1ZQwRK1Q
GFaL5YSgBSNqcZRCAtTgDde6hI2p+j9vF0SIHJVNlJfyqEeqH393/l8KaRMLGKvC
6hwRRTxUHASGkyBRHUt9pzy0WCc1G+gH+suEDIR8ph2Hjec8KEdgVLhafW/dHbPe
dLNcyaf4XCdEg+Ys6Q0ipaUKjDrWYsJP0YC5VtzQVcTFckQXbbi7n+RIJjJMTV5X
WnuRr7HStv5jO4U8Syua/r1QxZUj2s6EYsavOyftM7iIcQM5KgRnARBMr2ANAtbh
KyfScoKlhmVLeGaiG+w9toPsrHJOe71qMXMua2WwvnE2keklGB4qT1zxa+A/RG33
sDV0Zers78RnussBi0g2JdWq3aRM/pEMY9eQapc7w5dFyG1CNmitmFp7Lkt1ChSi
Ljgttr2blfsZ0iXUgaxCMRfXVmliwlqKefAprCv5PEqhL8mPcPsedYUVo47zxCvY
SWeLeo0SdQFbHLEZbanCqIQgJrTeMJImAbCboNRCoMimwDUAU7txY4ZBh7a6VVEk
vF/ABsvwalavOObY83ucrhSvKcI29soLlrBPD0O/YKs1xFBW7lUzpksy7zhMi8Q1
ljF7/8oHIBDHFXc2cfm2ulIeDN8pBivcNsPkN/5uLOWUTH62NO4PYdVG8oHdZVUL
SIZcSY2rkehL3oWTAu0g4MPP0CztvXSXyIBx0LTbexgxVocVLmHMD2Ir4l2sAQiF
3ljZG7ghIzp0G1I73+O+9mySowO4NNAB50qP78ODjvVgwg4I/p0Q54cM6r2TmjI6
t0EgEsMRxC8kbGX8U883QmMeVG4ezyKvgHtMWwwbeGrJ1eiPs1mpjWTKH7+vlzG7
ATaa7vWUrHFtEtR9/IpB+r2f8Gishhp71S81Hg/iSV62zx+zucD5gi+jo2MP+tfy
X/7ybmZyEjjKOUmzQ1ikSNG+X7ieWpPA34NetoBXRghRFyWVjPSUXTzZ92AOi//X
WZchLhxEvMxRBz4JiVnNRNkfgE7yACGmi4Xlpa/yUnCwp0MhP1qTESjqc7mT4MNO
RkkiPWtx+dX9UtwL7+0Uw7HVWxdKQyyMJkMChr6a1frmphuRTIJBhr2yB7UrfGjD
0tXcenU7YyL1DCfzqA6m02omVOqXEvgyKNmsnOWSyiWDwWBHOZxry6B8vHavDDiY
cGWlzXbyWsdVwels7rNwcA1SJLVrF85FDfX4lNa3Wi9b+UJhn1L6fFHcfFdjRwZl
95JnhfOs6/u47CNfEhpxuyzWJAx/Y7Y91TD9EdJi+t7ylE6nPFQMVI/vP/vlXJLR
rMDk8Rrfn0pigFcRSfxNmACkcmIuHKAptDHLRDEIfvVyfJyoBp15P3gFojfUlZbI
9N8pFn2sorSz5OlKP4+zVpnYqKJpg0BUhI03LpKlJL4qMabfyhwgCYqa7IG0u05U
v9WUKutldUrZwvI35Q/ig7ZhF8iMo62AF+F9qPrjn5zP3YghpM8vw9xSCT27P4q+
FUn+B1pvXh+PEcJvi//kV+PliIwmjX+vuEmr+yp9+bYHFe0BW8nX+KkT9JVZbWmT
Qafa+T9UEYDRQ4eb0pyqBVf++wMwySBKcwlOsEy0FDk1YVVJYlhhh54qA5MDViBs
d8hCCB/aZtYcUa8RPAqh6ccDPShDNN86LkDTQefBn6wt1xd7csirWhurjhLGiRrB
rewasdPGfa576SuP49AmQ5O7Buun8lhFq54pFJM/6vVE/UFZtgk5udNZsL5gB86V
oF6BaTdmxLeHMbBOpKbB+haRqO7u6kjQzo9WBkOWtZdSQUBmuwAkyMHCRh3kD9iq
Y+4OY4gyIbq2Ad9aZgllwNDCPsq3jRuic1FmPguwv8RIOXGqG6HJ/opT3VJxyXKk
XNZY+ZpY307pmPH9cYc2ZNgQhAmL35AsZuFCSlnSd1i+qrWRmO1MxgXqTyeKQ/ha
WWfBPCDl1VOjZbeF78pHWNfhxDtqpihXW5KmMDC+/rnG0le8DXnPAUlEFVqSSC3d
xfzEPs2Kf8ge7/4nF2XfIHfgbBPAndaqXZTIusUuYhmq8S4jGYG1NZFn8FulO2dg
fpGDZlI1uXoJOrRhSu14XSDB85FGpQCHTtJ7JjJ95pIa2/c0AwgG/80pssEYypXo
1DWzzK1umRFbPSjN3AYtcz17fPvaB0pmQTrbnLx7VYc7WF2jt3LdlqGk7dJQRBse
fOp7JP8m1Aj3SMH3RplVX62hzdYKJ9QGoJHUovYZ6udkPaLu5h+3EeTGT3BnTDun
YITXsl+dqIPTlRGxzxPhb79lNDzDnFQZo8r7D6a3EycmfzeX0xyqcnwYHnlNQPvk
6lWHCa6XAfo7+IzGTa0qCMmmbtN5gBl/vWjrX1zwuAQ27ccnElHAi5/UDCOSNUnD
X/w0QsmPjPuMo2sOURxALb4g5D6gzwe+EYfkCsla/hVAhnYbB5tChLFq88UbEjbA
2HzwBmRkdtBxG0Y3qXsBQX1Duj+0wJproyw/SliuCMoHx/kER9EpzAytvoKS2sfN
oKfUSt7vrGuTjpyXYcDsViexTDhNFH7uxqmkepg0trGWXHG7XO+0Qwv6xrh/mTY+
ke1f3Hfj1JOjrA1vbqKYpZ2qO5Wut4qg5RehoBmJ/+IjE5bO5l4VjxTVjGwiYyho
oR+YwoEkaSt9MiUYmR8kFj0CRkTcNOPazmRn3Jnb74k1qSrRCwCTda8PnQyv6uJa
MuI532xNGEC0uQ1ilCBY8EZoCiBJcYFjUJIzHBU2tD+6UQBAKL1EsDBJ1+5uMoit
elc1cfLYpnQErR6WiJRKkDkOSJddzcJOUl9Yy8MpTK1rgoHy9Up3fHVJMzCWSuOO
b9QhLaWw4/6EW8Wb3AiEX99MMEnzzIVeL36Qhwilzg/L/wlvA39CREjW25x2vtSx
37rRyUs/Gldglh4XOo6thxHubidUC7xI3prbjQmbd30wtJLP4VVpMlonHo1NynXa
Sl2QSg6BmLecWrR/1vS/BNf4mYwCnvuidzyOwIJTyUIkj+Jcq10y4h9QghgztE1q
kRj7PpAY1uas7mUVF4bky9rAP5lqqsjnyBMwEXfpZgpptxYidhcWwpAWcb/7mrj3
ApQTAQ4o/2Xy1rNqBl1kAdhq9o08hIglPDJVvT+2f3d7CEk/mtqfEvnP4RHCqMh6
lHIkDBrAzwhO8FfxfDwQFkwW7gNbzuaztT2KJ8SXq4Ms012Z0oH8QR5QttMBxxJv
imP8/3qj+hMRbDgLK9jorugaMOU5pdNMqmtQU5XpYn/VIflechUEpOPoKELdRN/b
1u2SPIP70htx98LG9AcI+sW6Twq4HCXmFNPR6YXRXmFkId1Mk01zd1DZ/l8eXK4C
y5znIbKIO3RSaS/VjliPIx5lOUL7hDg4GJjsCM16ODkV3/9M+kymD9oN6JVw6oKv
I37R+WBFAVOPBqnGZ73Kkz87//0sozZDdp1iuwtYzlGkCquZb6F3hOYJDDuJQtYK
PhdkMxCamjwVKv3PSAYG5z/xkdadZhvVQnXcskK/SqY3yQ0eTRYUbjU/T1IqWryT
hx1kQJ4TIYnTvwQlFiAwcj35KpTOkMpl9WS+LZfKO1eVymK0eG1DduSMB37cJO/n
GQ61sRe/a/it11jhCQDpIaDn1C34e9XBZeAnRR1UmljMyBUv8jWCRr5Ttvc2Ltse
zIIaAodQcC2f+ccLloGymMGOcy4M9hC37bCOcbvz0f43miiQgPRWxOFzCHOzZxgh
/x16XLhYE32VpsO2h/bCmaej91VQWtNZE/6VjtHm64E7+cESSWVWmmNDSrk46/ls
AkenIn7GYzDCGmct4IuHcOCBmxP5K2As/x9OVXcAgtk7+04lPNf3x/bkUdDhAed/
BVxR5gzg3yaf0E/TgMhj1VnizUVoNa8tgINWkVl3Tb6lTIwQStzs46cfEeQpaKoH
m6xTKoRpqTynJIxOp9DB/aVYQ1nHRnA8cFlBc97D6K3mHhIoYCuzQtIdLNkEylVb
brgCmsL8RvN560Jfb4ni57AfFVbgkUNCK6QgpGmZHlUDQ80j0Gig7rpnVnlEA63E
A3LjVrpnWk2dHUI/MY0rjWjz1KFOA6oIESjlIPTLL5dP3+Mv3wWCyKvq7A978rQc
mz88C7wCygqu+hwDWlf2os7iJC3nDw1lB4lFjRaNTJmbBtEbc4S933/ku83hGaZ2
h3tDKOMfe7GpdG9NmBnOk84Ya7cWoSwS4giB2yKh1ImilYE1AR7CoqDHYugSFFXs
6iqdELKNIf7PWyclHpbZ0O12yQeHVbG7BzSWNB0G+9sjxjlMY9tnDYzIO5RwQKpa
6VZV2XsWMOonCGvvAyYywfyN5gCuahbTnEb00vp707+K+VaUxItMto3I/prKhdV5
aGAF1vnEwQstxRfJCGFW8jJrEjg48mmlv99U1fokUpJ9kSI94KXar1XVnmQvm1ET
HmQkPJ7LxTBTb2W347OP/O9SAiADdv025cGvGkV2RhbASzYRdxH6ibUDDse4HTNc
3TT/D5ubRIKuLoMLTtzLBypeRcj0jUWlbdGEiKDG4An46ZqCBhLh4FsXx2qLtv13
6bJe0r81n6HB3nyrkrz9lISQ9xDiL7wPkMql9CrPAeFMxPrttr8n387l9oXrMvto
n7ezj2RW8HxCLZY6txtKgNsgVbK5b6EEJBPSFzMoyziuRt/CuN6kSw5ED1Blxt1p
qWwth1Jhy1XvKq77AUkHLUMPreADvUSdrK1FjI6TuN7vuk+tnm4pWQi5H1xmT3uP
a4zYRPIZA4kK/5PQHTZaby5lOCpPmX+Q0fTOeiFEmpemEK8wI7mmcoeOldqktH8t
Ty70ATY9PHArU2509x9G9jBGXjk/tPZz/AZFeqWo0mfucT72Mh6WKfoAuqTEY3AX
SSv/8ezeffPNRicorc6iSf5TxYk8FZRi38HiYAK607qDQxCpiocMkRsnI/Pyv+wA
VtgdzxRNeqbM5rqFLfwigBwgW2aZh/3iA0oxK2tWAqtcfeXrkEwbGsVgCdvzFY5f
S5N/NSOCK4M64z4xXYPa6ACnuMCXZCMhGPtvM/EtnLjBRUOkikvVfSDjpTlcZEZT
SC5BV7zueKZ9bphw5DV+lx8B+owboUaE+tg21w5nsy8tOU3IhRxWW/vC7N/OQH8v
AmnLgrHY530UUAlexdA1ZniyVaGDF6TEUsMPQCP9nOchAivGPV+CGm3SSoHMEb2D
wgiFouzx1fvyDUE62iJhuJuBBh6T9YI74XEr8nJ957doiqgO3v5YdA3al6Cywr7P
TlNzMaSGX/rUC3ReJz5GM1n9cX84HNgjvgd+/eKW5WiObu+VtwU3hTgC+DOOBXY1
VfIq5KC5SdAsvsb4dgLcb07ZQH2oc0vK7sU8e/JlkdovyKWAB1Y43cH3kLcFMftN
CDl0EzDWDPwbnZGYv0zz1yOJLsXXMyTQ1KCOUt/RHnvvLOCFKMVxb101R3pokAQU
EliSPvxB8NJNQ6DE56EpsfACdqSdnt45xfiQh8cYuTvJtzqHON+LzVj1TSlvGANl
+f1h2jH1dQ+y6gINI1IrOuEnWLFrx1Iu9OABrRM3R/vou03wfA3b+wVT+lNyE3UE
nFteHXGlBAAsMT9kIZ2sI2u4JbV1DnBNjJcW8C8sBtmnLC2hlwQJJUxmUQBV3Twb
VWxfwtdrnblyKk+W1vSr5u+tcuoS9Xi3jfFUP7aigf9HggqF3aLljYyTNXt6FaWJ
mSJKexlPKrJDYDSnhv5289fvxwWYY9e+8I7dLpPMPCNEBh7jPRaQIBRJ6/JRuIF3
TMFhtlJSLDcVl2nwzmJFanFQj2RMYQFz4nLInXDmNRRclFNsMK8+fZAhAQEjZ52z
lACs4pS5g7TK24d1kCVovNt13N/g5/xirC+tOdrAllqhLTg8YvvkKTdPGcatRXsV
YlMtxX8Bi5mfOHnhSbRyWPdJs0k493XKWSFFrjHy3OWTfQ2J47sRXejUM2eD6+X0
a+A7Od3jmnn6P9zDSwAhA80LfvgWxgcb1kyi++thqZpNubvNXPiSvjcc/gROymsd
bWg63TH7J4Nf2BzFSEcoPquJxdvXeWiXpnkqdZ3WfdWs/KRkH5ZeOxUYrkFP0Az3
0IKLBNaAP1NdkPrlH6CH5PUJkXVYA17wz5c9/+keH8uxCnuW2np9p7YiKIIX243e
HHq79Pku5SnPeojGzQbpUxj4ZJ365Jyg1/jCHe1tC0C1rw+9WzcYS8pI2NQQ8r9z
XfOG9Re77wUMywsMIKFEvREY1rKhkdEl9xTqREXv8Fv4I0BxJ7kwJwcwcEREXcyg
V6JtuxwRrBBC8z+nhLSkde0He5+xxEf5HHCUcuPDAXhDoSxujb+qmpHcdw1fhZEP
vF3CioY3AQT/BOcl1uYi5YwXW/hJloTOWVILqndWX9Wpf6NrY6+xVAjemmvbbbsX
wcfeXpoku0x0Us0N7GdWJdwqy2Pqaq2iRnGLgbGap6FD+WN/oWbdhbRyZ9kRu8wl
Xd+o9ca1xBgLuWAuw2eUMwoRbUJWyJEsnVSNAviTcJ7weRs79EoB0b7qKcCCDyKf
4d0tkVpZXkgc6ReVCh9+cTGFj6Wttp7W4jbyR9A9pwTMLOPM81oM/APnkiC/J11S
ETZJs7fIliinedSf6e+8rtquiTq+ROm3SVHX6dFKkz5dmzZakzUSxbMs2xrNQqyL
TssyeAXfpU2IVOW/6LTFiIhkFNKMgr8lDUVzBa8eKC0iPpAgkGI5TzS7si3xprnw
fph+C6kxqK1D3tam09Ui7prn5sad32ZtvJ+/SX5mY0zVBbpt9G4TZs8JCYuMP56i
lcwTyXqe5IyOHgE2SZzUFuJ7g8atimj9SxWliecAfZGuK+8WP/CkzmKuH+ufr0se
3tW+ETNp4KE56JLIxBieu187KHbuYi2oGn9hpjBKC2qH9ykaJbDNugKoUwPP0cBG
tCXONrz3Bi+KRf9sXY2Kg4B7jGeJZD88sGVQ0ZnlABLd74zaE6WT3g3wWyyukJ/X
NShzeJnJQZinaUqt/PtWoshJbCU33EjBxJ/EmGDygU+9R9us303AgThDCD1aa4FR
bvtm7w4F/bw4M9O2Gv+Gt4QIhy1GT42tkFHWoKl5WBQYyYtm4+7XItgyfvZaD7wR
MdI9U5OfoUiHYxOy2F4kK1HrvDgodUB2AC8t45v/kfb+pbrU/+H96jc5/Y2lkgQ+
xL49SpuXGcu104MXUFJ4rt6DjOJnV7QrKzrXd7S5pSiDT6jKiJXuTc5eFeMZGoEe
WHakGb7Orlax0bf2Jx1+Ir9YLPLhEJ9zhOuiRTsYXOCAsLXAQOVCnpaKgkA7d7IV
UPpdZHOT1sn5gkyu8MMtCLPN5lsob0looq7ogxUIWdcPZZVeZRNDk7KbSA0q9cbd
ISZ7ZBcYonhywQfEw9nja1gzsvWaVnCFFVp0mqQl1DeixlD/dsfYLXdiqYZpeJ+Y
yx3RN3bqlqDSuzNipK7F7wFSCZfbHHf78NevTaZjtdxOhgMH7RCAcXcsHualKEmC
oREXt37KmDlLWYUcbdHexhdv5u69u+dxhdTnxWh0Go+IJsdSPj+fWkn9nGIkAzXH
Xbef3t0YHLSqIa3Jcxnj0mC7miNzAcsNQyuVXcNWIx4hSxkeCPhAQqDC9bEEcjLZ
ucqXBNdiSyF0tM2J4YfB4B7bbu+ThPcfVx619LPCNplhl6TbptdMU5jRzTHqY2Ph
vuUdoEZgScBUTYGCItVSV3DanPrVK5LG90Q345OLXNXLjwIKh7F6p53eWAiwWppb
U1UnOFwAmS9C1MwGVbWEtgnxDPthd/hfM28GZ9jS6jiPVR1CA+/YGODyBlZu9ex5
qWJ6rVnlV6qslz7p4/IklZq748PlkppitrcANMP+fx9Rnki68pZFuwkelVC6kYvj
wG5qQtkMlG7bpuVOh/pFzC6ptwSEvOJyfjqDhb86FnaVlei4bT07RFe0KncpXmuZ
zKjgkSp5rewAG7kDxkxFH9Huf2oP+95nnr7UMSTs1Fcqn3KbXAcNk866oc/TTvJf
5MarLsNmGzhucRbvGWVNnSmsjR+CVFmLaPmSuKbgJ3bDAbhlt6R6bAFoXinqGcJ0
BfBxQ8ymUZ8ivGfilJ0le78pOMaQgAdELInIEfCGuhqfbK27gu+xplK7PWqkO7MG
h69hELwdz5852aKyEk4DpRFthwo2hDVRTUoSH2VU1Ctu0J9II7jpOrPYsC3P4SH3
3aGZ20f5CC4MNVHF6V3rcfaMFJ4Kepr/YXPEzjX/D8avT2A/oL/VwiqWvv05ReaF
1ZKiRM+uGMDbChmClOrT/HVwzyFP+DaFAbpQXE5FI/v592i0dFqS9nxBiX4T0NiB
odDhTtTJmW/Eg60Fn+gQIjZRm8RDzRFHW3a8bvexPjCJOSsizINjRduEoufE58Kf
UjqF+O/q4MIK3px7A7NYYtA6T4DqmLW135Jty1rpXSVQtTiKl/YHktP1ql2mZw3A
C9rPU3FpSatCAeROifPOF31t4S08bZJ07x8Cp5VuBca2+9OyvOgb8aZg8kbhiDt3
KO7S3JJtJtmmLeRausVAz9iV5Vm8WNEwZ17Q1esLrutyUzr0j5h8E7C2mS/+nw3t
rkhLb9qdoLFejUD4Sjk+N3O9SV13DBGhnh1ed1Uxdp/SQpQ8wd0LBKS9twBUYIFC
81hL4em6C3Pw33n+O1nQ2gmsV2XN62Dnt8EghudwKnRBwOXLV7l19FR7IpflYDh4
DFF0AGdFPn8M7XGkxOSkUJFygL/N1qL9zvJ6kdCPefXcf8459bbiX/i+OnvJex0J
Ypssz9Y1m8Bmj262X0fNgIbIHhEYQ7ZOIFiiYpwGD0l5CpVIQ0mgAKm0XtzQaRn5
g8FR+CxBxIHlj4zPjELRaS/C8WfSviYWLS1UkUrjWGryqPhWesBCxleLNE3FhGDI
YSDE3UBPPsx0JGzOctwRYzMTL9prXUcIgQIAiy1XQZ9L1h5SrRxlF0ffdsEhihva
5XSjGlf3J0L15EdTmZ6zUmPA+tV/z7/0QhVFpkLJOTmm+GiSSYyPdKUaGNjCjgqe
Hoz1AI94wrijzRmHOva5NcrM9sIso2NrfexsEKDaVvLADsIEDqrCs95NIPhtpXQW
iz1yLg3ri4YdYmPoaGMlZywef/idDBB+W+mu1kR7uUWMkQQR0FdRcg8Wdi/Opp2G
M9PwbR8wk/eThNi+d+tCb79OI+Ib4oRGjML+OlZssqTIAc9ZSd4ITLbEixtL6mYB
KyBYr1H4iEkf4DnAQks213ZvVgzPTDDADavNrStVLHpLSvgljiV+iQFVolq0vHOg
pTqGm0/zrDulVRpU6T1JqHySfEKoLcF9j4zZSjyiydPshX2nZ5dqx1lL0IXrSlf8
AMDopjIq5WO2OMuxJB+k9DXxeLBCgjN9ZJ/pGWUZdZdtE9atS8vqiGlpepWFN48Q
/2/pMng1hPrSy4silo6Eq8XNzpMiPk65AMOF8tyRgDRNXv9Sk/qDW4Dl4CEIeiiU
cPbBhB1tHQDpawJYYHONWjWwfFKnfNTuSmUg8WrZ+Cs85VWjTPinaNhPe9KO2sPO
i/56RSQR9Mlw2qhOidEj0FWuAz3ZCtSCB9/btMG5Iq4b2kD+R3bOstehpTv/cL4r
AN1HRDmH2lXj+Pa1vhFTrlgizNEsmJN8SR+Cf5U/RnPm9KjlO6wV8oS2vbT7SF+A
wYnBTRMPVImPwnxlarUcwzM9iuYx2hz/FSrFvgpa1logYm3ygGfH884jvgKe2mkM
tLuGQC1JfP/8t6wocouXZg9qODpzdrnVd0fk1BL2GTyyyvwYpmScHCc+XyF/PJTP
UKKo9G/CCSwEk6Rkv+HSkG2BmMT9RtjMsYpXokGMz2luqexNTEi5BgKxqS9FHldY
sDdVd6oypdppKMNhgHdyCC/BISnDVoVxEy3KjFjB+anWDsp5aXN4DX93AtWJB0mJ
EFj6qZPQ5VpsJhFcHLK+mn1ROwnpSWeJ4fj8myjXJY26vjnOwR6devTDEmZWMzTV
4aV5XmAoytm5cbUYPtRVJ6rBLpQdqZ403LqQI2h6Cb8+jpgC09PLvu7MJD05hSp+
vuDwtkW5myYopGzkrM/MKk8n0komHcg/sglAiGDzbUUZ9B9yR0qLnpY1LQOCzzHD
Sj41iJ3iRuM7g6FzoHqQdmKU5mxy7dnpBJjSLvVXxlOUmAfENbpC1PLc6CPG3Mq3
yVah6r+SmoGqxTz/XpHpnVXAWhCjkK52uf29GK/vBJZ3vXvvwwIv5FveXVsAu58L
q/8F4EXO9dIIRz6t0xp6BKGXKWF1Q4jN9PBBZe1xdPBKu4ojvmw4s0rfwK+b3JM5
duTTXshyfLcG8kftWmvPuiBx+xgeMtrx/jUYW5B/jqN8vt0gLiegPMrfhwmw+bgl
9Hi4Vhlj/YmUEpOqIMLQhpDcTlXp0bqG+oPqPO9gRdwdb4L6tV5jSD0M/eCIWjqq
YXaVqnkzmK8A8XUvkTqi6tv6ZPxr9jSK3U5uowFQWPl4S0Q9YyOhFJ4hUDvV1f0b
yXIGDaKiR2CimwlfDA/10/T09E+Al4xee7F57sR462jNMLvLr5RwdYhuqwKrNzI4
KlpNMNqdYzsLH6j5ZhJVsLSm/kH+ZRqEit6ZkEJnT7zVF2SLwIvAKf5J3wrpd6EX
Fa8Kye9zknZwwgrpmqVhB7uEASh9/7gct2LuMyUQJXKXU+06btAsVoDUQjiSxPYo
pZr8puXxxH4KuP4o3qWlKMd5MbC3E9uPVcMWYWvVXYjOLjCYA53aR3OrmXY8Cslg
pkiCsmcvDc2x+hUQIx6WekLzLKjsXMaZJgLtIRMd5P1tL75rP7MbkmTFnJQSZn3k
9ay2YNpsgCnO5135P6tlXlfD+lojcUk10OMRrKceomOpwH2ib5QdnUtjrB69g8LF
kA0o94ALP+/tGCAF89eFTyqYoOwxrDPIXn/TtT+BVT+vn+Kvc9z6bXD9BAyn4LBk
N4WYnFkQzPHH0JUMZksUvI2659/ECVLR/PLRJU20LxlBYWODMubDgBe+4n9lPKqX
BAqsHSs7NlAQc6XCNAy/D5N14fwFmqR8J8zmvM0r95FnGMmqyYZXLXsE162TdEnR
7z/VrJaDpxdsRuslYSVNdOZN0U6op9TTcoXdCcUkWGzaL/l0Qq/TdVTWHyDTHBLB
Z5Md0wk7AEnT+U62IgnavajpCxet0JKFfHkIhWQE2wGUKBsOG+P6flO/NZkFTor/
mjIJtpvxc9Y3Ba0hMZWRnLM7p9Jl48m6xBLGk/GEUBA+ej44xVe2mMWYlbvUtDaU
Oe5kjbI5MtrWBT/SPHDCZ6gZk2hgdvPHMuIXwLSBmEv4gm7A/81cwuX2hvoQoTY0
r26n/wE6xp1+v/VF9UurqrDO1DxR2NraSUm0aV9yX/8gphjoxFiQ4U8FeaPwZs9P
NPWdNIveG6sLmLVfIfIBJ1Jf8PZK7zTOw0xsVj++CDyK3mpHwabC83+WJHHODzJU
qit5FVsY+4Cmcm539WcqJbiNRxHDnbK9U0fpinjycK4LaUk2IIgpi0LKueDvucIU
hDTtLUg4MVb8sCeHJYBMG3y5iwXruxO6UgkLfUVLvPy/B7iaYD6TkurnQDmoFwTe
gfucOk7P6O4MefiC+mIEkhUhjTeF05tjMuUumLHoGDp+jnO+HGJsZDaGzKje1L48
tzKpImzIcjB0pqP53XceClxcTSgkhqzESoOe43yu1Ll/UHC941E1LFwLLCXN68Q9
CAEJdsGztCW5YElTlOIlIRTtWlQlaaWMDShH5NwIDIjAsbVA6w2WhWFawdOs4CZc
+MuiS218TcnbZjIAG2Yxn6BYc5z83XbqKib9ah3r92TMsDN/UGE4ISfL6apRIpG5
bPWCpGDooprj4gjisqKavXx/o6mhXJQfproFBHksRB07RJQKhorU6jsWRFpoGTL1
PMxTJyfmW9p13uouOk7QVoyIWPwgllKRQ7be1K98NPor0KDW18OIld8vk7hnQgVP
7eowOZ4lVQhjogwPuimmLS6mVo0P7iIiA8DA4nX6Gz8JOn0MAPTDYEwN/nKOg3vn
3fXAd/8FzOC2+bGOBa0P2RrVhKXlllTN87JFiWJEnhoj1RU/ORu624kh2q/fCA+l
NFp7Dv2tBi1JHVdJggmwWIXJ+cOF/VGhN/YZ4mfZT3zsjCpLHNlLMkBlP6zsd+iJ
Pl1Cb/riCACymP1TuEmP6WhQ3UQ4fp1gZDWzQkUjIDRpRpIYT2EAU1Gknwr7GYt4
sT9x7tG+DVX8HMl7wmhd7FnCRPBgBMJDQapIKv0Ip7muwjIBVJoU/TKKdQpEwirb
L1MbQ2Y/k6Rct8sNewRKRb/WPsu8zp0rt5qX7vsLIRJkpn3YdTXS+RzBJunWZ0dF
iMZTlbhKwfeR2KNZQxWjLI+sKI3nyqsTgj8/8YE/d/fl6p2mvj0mi1IaalGU8UQy
ZIVPci5Tvcv9xSM0Fhfk4cuY/hbyMBHGKcb2AezPjlrzeoBUm/6P8S2vi9DsJ70R
NbeE7dClXSjpf9Is2SGm8S6VjAGwvj/G7tevbKi9e510Rmq+QcjcV6rfR0j7yD3r
iAy4S1NNjGCAyJuVubvWLv2LLqbv4+Vj4G+0ToFlB7/0YmtLKdqLvwQL2bPuH5Tt
jsYbhp4BXqis83LSy8i6Gwqsa/yfpyTL3O5Qk+QpWsv/nLjQwq8ntVN0DCn6Mv0v
UwhzZngAtP4JqzIev5YmIr4YdL+f6unYhIr6gbrqjCYu7rYH7CjpLPq7o7MRjF9n
qBbStqy+eYCtiVAqCe05ha1ad/MS7Pww3ZSsZL58tuLQxVIANO2QNtvmSmQna/VV
MUMETeD4DTHht9c/pJJ9/mSne2P768Fb5rnEzF791L0e5lDdulefaTlb/HDEcLa5
26p3kX/GUo7Jz1/LS3In5CyFwWXOUzbVwrznz6ItfxqICcysSWe5cRuBgNrOUfuQ
stf+GodQ6SLCeXvKMoUE8ekc2kjrL5Y3CLLTAoR0MuQxPX6G38tFHOn7XZYcvWi4
EBzV8CjOojf0uhp7kb3i1HwYcdrEvWGq/UY4O4/0yV6ZxpRphZ1VaUEd0xezuJae
f3UujhS9p7ptiQMBezzxkyhwCF82dPYauIgAMcYg826khVk2zmX2/Lr81Bbzvmn2
xl7fRXDbUquzFOVoqidZMA2N1WVTcO1KNmQyKX3fzInJYpjKslwbsViAiz5cs0jZ
0Cw7n1WRQW7Kk3JqmCZmiImqJH6CjRee641AzaSAnLROzT03zmZ9Bso1fNcL36sK
md5bGVyGYAId4kJRCFIGxbVLDZM2UpCVBaFo0NkIDH4XvMeV7dT7BRb1j+wEoeHu
Xs+GMYJpkk0MfaS7tW7RkAziV2kKagsfpgoK+Zp63lckLGmn8GrZVlKP/fmBr7Rs
JVafNfNiR6kJdfoD4abnJSjXwgGur9AOw6uK9MOxGvVAQEmlsxi52wSAphBhLDT1
HDtYnBu8XVZjeu7snns689wxJNShbQRUISEIqf7wrofYFDgqgjPXueFSSesP+8tA
2PcKx1lwpPhftMKA2le2ylapWlwPCOhKf6i+4MZiacyYLnY4JTVfKJ6k0nVUNNBi
5Us1w4gywOdgWG00ruoT4zKndLhHMToEz80aasFck5zZW9b9VaqZMgrr2X77ojHz
t8VCScFVnedbmTY6T5JrgHu8QZZk7orCn5mbpPAMFPITelCg+dY062riMuEZdi8E
tzZ1I/jEBkApRp1N6jcr+BOpJifG+Uf2/cgQQc4AxdgtpFumrm12Jt3FDXJGVD3l
+GzHldn6ZAb8YBiAL4ervBRgz0r1YWRplaaMNvP1H/b3TYC0DXUhtnNBEs4XRkdl
tA1ou/sbHOiAJdeqerSI8Vu1CfBUibdStO9yMy61yJnNz3fCtctmUupDcmXrcQQR
umxf33Jq3MXea6cqmmOTgG34gxCzkEp+Mug/x7WeffG2W3AuVRZCIYL/WYm148rZ
qQUNHMf3DHy9UvlC5Hwh2H37448fBca21CsrObmAoxwTOmEwXhuO9xdb+H98Niwe
DlKHIqTrNU0YIppMVl0TO5JMcqbDRyKzEW670tYVKWGkTL0rGbhpus9CvG7LLL+V
PJd6eI6BgOLObGbij3uXO7MysOdNhj+qfzllMyV1PwdlnY0/LWE/idOaasmmo1cH
KWeKsCDFjeF9jlflNNlb/ajG4oYF5LHaPN3RYDzv+h2S9WbM/iCSnfOEkgzUa4gs
gsmcB52CexAHsgbhRH2jHoW6jFdKkHwnW6Ce3b/nypYfWZcg4H2opjNaIr2BT2ZD
Ppyg0nEfcx8AbfvaTS98wUjsQAaRrjVjLWhh9MLMVXdHTSGUheV6AOAKB8Za+NCa
/y3AZLk9mkp297QxSZv6IpYfCBsUt6YpzLvtiVXJ2XWWPwZLmPY2xarVNFBjWnud
uLuirpd0fgL0//ivbCXWKWfBig2uc+1XS5V8YtEcMd4kzGOKFMfVQqK+hXQSOoIu
QXhNalQ8aIQWcc/1j1gRyp+GgS7uyf2tosIR9/kU8nfc2FYh5qA6ismFYwxaxhfQ
335Y/eGfX83CKSdXJUjOpKBaqQk1oPZmUdhYquVKa/NJN0HoBZXQh6Akq9nuNgrU
Z8xOLF+iF9GkQ5OmLEZ+pm9g9quuXV7J9OEsnK4xTz1mGtuAIRUUFvdOYM7zwVYX
x3mP3IY9Lk6oOSOC1fDEv+b4+DvcEzPqi5lAXBlxXQmDd4oBnuLe02MUQ3Ul0wip
vxj14PINE/s0kRsX8uljI/VOZrlO9rQxyJjLTXeUQeS6//eXhuQEMRVl4qNNOTn5
9Ki73NSCDdMq8GJCPolcEpQUNhdhkYsXpbDMI+2Sf+1cyfibKlPLsdJebXSEPICm
CyuzXkVHO3s2/oAsdqW9xTh3mWeJy5lknSw72+IOI8F7HiuLUb30q6DS3NMl9Mj8
h/QtyVZIhFbsQPk0xM+F71PzK6yRb4Rlg/YaDAvfoV2H2+vL65UPU8yeTre5jv/Y
mClNUTcqdHmFzCOrJ5PP8g+V4hMwst4WryDz9r4hwgh7czKHTiSF/VtrSZxP1lpE
1hYJtzKn+CQWeZ71tzow80fynaswHWejFUi1hqZcHz2YnzqGEq5NHlZDjhQFaykr
tGGZv59MFzQdc+zB14E8gB38NiZ/m9N7LH53+BuKJKm04zoynnBwhu4mvixizLOJ
wmByuTnID8HgoeG1ryqWOf496AhsNl5DRjG+yiZ6f5AAQgyuybcsJ5YXcJrVTFgM
hqCBMWEI7+/5YrQQZcu43PJskNF5x66YfDjY0vc8QTRkBcuNeG91rXallVffImnD
UPiVSF3ZuPhBEFnuUZFxCgJZg1sW6vzUXdXpF0/S/tjuwXohUUOnt+SWZr8GnJtr
Hz9u2UTSD0C5ZEUf/IxGsE1TA3czXJowOIbXQVqR2oy9VQCLKXtbF3A+va55q1p+
5NsXNF6L3Dz2KG53dqkAErUDfG/32SABZN7NdFEQ9Mp8ZijzPpZVu31q1XrEEPz+
s5cj1zG/WRe29YErz1ruoxRjZOM4z3A3Lsx0NAPp5bbOgUTqH0I9Qeb0ktUE0/SE
7uP+ci0k6hkjBts7Nj710rxNGmax3cgMqtTDtB+XCVCq+UYlhHRuvlYhUbn7/XU+
c4NsmDLmtXTLNBP/xLYVSg3bWL0/9EToipq9B1rg+/So2lzX0p5YXJEnHtjUEpUO
fOtp7q4gBYqJFthKJ2CTXpT6gyUZPm0rVsmSnaQJlEUCRBppFZdSL7BJIxtVRFnh
PIx2ERsn9TGTBLs3MVoNtCaMS/2ZWl/HuxEAC2m1NV9FSvgWtW7LtBeZN//EwIwE
hKcOykV6zKVFZWPi93cGgCr+bLzQiupokXUNK11hEGYAZ6vbFfrX5Cu6pgESXC4j
43EetwteWL22ovbbkStrekiJkXaf523CV2hkse/ppDDcOVlAhEmozgIENvCwouAE
HEuk+yoQ38JwE/9n7wSGE7hCU1xYaq18o48jicXhagY2dxy/C17K1qWUygkqHQaU
fGalbE8uM1pZo+IydaZIefVfzpaP8IYhKtxICcqMCl4uDuz6IkNz+Um6pXuA8lbj
P/eSuHNL6Fn/e3a4u1SweuIjnekYb+qJlAqAph0UVdWE74KhKjY5busLnkw3ZA4L
Ml9vMSOheMF04W9FMDIwA4wjqBsf/w6kAWPRRir38PFRkRpKB9aNiXkZg2bsZ3G1
S8psGZNpWdOH0HZyxLa/ndkc9obw8EhCjLtC3MXlr/zjPkGiQkjI0W4pxTAesilY
2cxmuXSBTsheNOiwYlHqFaeoGsLkzbVoQL7/CY4qe15z36qaUpsKT2p8drZxARP2
kqxnOiYydzzgjI3yFBdTtpVf/tXmvi9WLJWnKpbatmVOrsevxyYggKMG67b2F2Cy
Mq6+hxC1iexoDMIGMI8Hm/qEYKpB8UWkS1kcr1N3yvU1oGVM5soTwgteeQTEn0t/
bDI1ZF+EjOxHYmVy7LlRTBFEERd8FiSEHREMh8okPhzLilWHs/iZuGru6dE/AhG+
Sh9S7f4mvgP3RFWwPO4MWgwC1JdYUbaGdzXJl8jM4XcxT3YySvykk+8QWva4jJMD
dW7XM1oMQTOWSrYEnUOBrsWR09aexvDB8tR1pdvBzIDMJYThEysH2Lz5jNM+EOef
oYSDRuCmc2oVqCRGCciBRGoXMpOBOTC4WGZ0w8E/hH34DmRwgqvfcthE21F7OJua
Qrk9oGLDA8QAOMoH3HLeW9CPQTnAiKwpO88V3JfuHLGihxcwxlyY0MgfL1tFTdwx
1KS4BUUA+SIbcpnRmsaEngnIDiyPul3LannATuFvhnktj4tOgasYZt0+GoGcUSIs
DTX3LmZLRVAI2IT8M/l2pLKLLPLJww3x67QJaTuksChobZ5i70hchBXHrvnvJeQN
qE1Xt7UtNSgQ+Zaz54zyHjP0rpsPOUElDi3xFxze+H9rOsRuztoLTOmMuHU36gum
VcswcoMrdHv0cQXk+0KQTAB3u6IWr/L7rVKuIpUsmY/4RklvHSJ1NbyeuY5UF4l2
YJYR/9IPC4p5kifiF7607yTaE46EvHsJ6UCC66o1Bx8u8vfe6HfOcs9nASfDgLLr
YyL2fb/ZfGyDSiEesiQw6IwnEJUiWoEooFDXCwxh7Mf6PR2/U48XVQUNq7xav+OQ
8+IcfMMhL+a2oY41eNXVjqRGfexxnHDoR3mUlWtcn9bbVfEk5DsqGfri2k0U+B7A
AZN1P394+1nSelhgDo1hRqAfQSIbRbGZrkhUBbTPpUiqjjtOxYBlQAiH+2O1VkaZ
Dy+uz/Ai7VP7b6XElS1zA8F7cn/omi4F6fDbvdpgSqilufkCqRQvvSDnaXMRzJtz
ljXeAimQpwvwJjn+K8uzsMG69TRMqn97TfvWJs/6kxl1g2W1NoMdV3ZBb1tCIMJn
eI3nrKMA4MNVOVSieqYLLRoD78s4f+jwIYd4v9a31ZeVlIDOsxiNVUUmHAUPRVzP
PlouFJJ83cWJPRcph+1Qor/6fZdYrqpGh49Y8ToDGAZfgqgGsM2QYghPEk0WBG/7
VZSTlZPonJlqIp1tvI0PMqpVdUeEdqNNcftBrZtIt+axTWaiod8NFBGsiY8+P7CX
vn7zwGQgNQujKjUoNnYpp9nguBpe02qNBOJ2sXAPhnuAQtrXMBAPBjnKY6Bv+PAs
NYt8P0R+8iYEcidRJrnNekB5f51SrKWc5LNNFc6ta7fvYvCRYTmB4sZQJuEMwSdn
XN7f88C/Ia0cvl8pRa6Ub1dW1zwBYy2OIO3f/6ZqAUvbu/4bNzE5xWa4LsGp5C7a
xXPa8rsAmIARJ4lE8ct0pz2sZrqtWVnRBbV7zbXxdPdRGhqEZC5YgLi8c0l5XTap
0zBXDqtW+AxSjohG0rq8J5CiAODMfzKkBzM/dr26RImxOFdXfIS/5RLCrAwc2Kcj
acom6Jct72glqSwx+GFnZ4avRfjoN4y9v0ta13o/Th4Zjup2aqfcOV3irEBjoW9u
N9R72OPvZH87A8wjin9iENB1Y+7T+GkGNUkIBJlq3vh9mvo4d5HZX3sGw76RZUWF
TmKycdCaxsYHB+ZOj8cl4Df96pBo4vggrivcPew8HMaFJpv8EmSavH+n16V9FxeC
vEhiEub0NxHLfksCTjQDVNmPW44MHiaf2eixWAP7BgVXEZeIbYUXyuNWkbFzKeEI
F1mCmpL2pksUSPwWXsMFPJ2D2qjAxBalO9RmDMCJBLEOC6gVYK+ks1wuVIcAX4DW
oL4GIJvnN6+c+beqmjM7MRpp4RjKINZszggGZdXEjAt+xPa+SEfzRgx8bvq7r541
kTtcPNeWVT6So52JTCb18lNakog/5NPDe01bycyXejBifN+ZoQU2AU+aVnfaOvVY
BAVn9o5kNtIbt18FKXWNVCWbTLg2k1UX+xJDzpdIt9xsWD8bBgTYxODPLzLQMPqO
CRtAkQm8Vc2xWexY1DXLQveKUo+PDiubFEeJLtBqcQIeChnOzHCHnZZGuZUCm05l
1ExWp3RFd+u8zYPVlPcwq5sTvGro0OeCzG8Zq3bx6FLu+PbRrwgoKAfrzckD8oTT
uYAcwR9jGbBxPH9buPvX48icF20U4Jvk0jK+1klVtq8KCPt2RfiW8slP/lGPh8PN
PxhtZ2BDtn107kx7NqVdR70J+Gc9wWCz9olYtiUXGbPeIcxD8VoaYwtv1KZ64hxI
ETek8HxEeJRPqR+bXuX44XjRgbY5ih/Tey4vo6wgQag/DmM9ooVRgiJn3bWS9D5N
uJNuDYq2kbbt0uU6i0TjPzGsvYAP/VLVRJLoa4MUqYFKSpIDLMPuf6w+XCFqlmhy
KJ+DGZi1Ql/SGnrmeBQQgQZUBZModQviZhwQZw4Fq18UNfr4k7z/8wMAbBNUdjKH
Jr5cmwCiUNyWDzXwkePGIf3z5LcEFqkMBrngQlfTnkjkBKN1IHQPRTfeE8y0XH6G
gk3/XjXy/YE1H30atlqq5OG/ZrFmdSBMpSRUNRlFB/zlYQqMJ8fa1GHpG2wTuVEP
sxFh4RgUfDkWPWd9TOiUF55dCYABUeAziCyiJQXHBOs+afvGKJ22oz7VcTCF3nC5
DS0RXqyEWhFpNLO56htFtsplcCPocGFq15eawsDQipSuzAnpUp/FtX595yMXmjp8
vAIOcwElFYkKIZAfhdeWqd6LJh+U23k2ONnIQHSCnTI3TkKjha8yuI2Ih+0Lb4eg
BMv/3EwLb502ENCTREoG5D6u4yYKq3Q+p5wA4k0TVCU1Y7n42XJKKkjHmIehw4k0
rNgbWbaPiZ+JG853DAxq08uI8JO/Be+LSBuuxQi5YyvQfeAQA3RJE8L+5k9JIMix
1Pp0obK5/pVcooboIdnkRifW2V/yBONIchngPy6p+X00WBgGgn40dOu9UCGOOvbf
BjQCLLb68tXE32SvF/TkGrKHmYMJNzJKRAGgae7eynqjzyx4hSh+2hoLt/ahYxvA
AjKhxljmbNToMKAdN6V2/LhcRbg0vTXiqUpAnOHlQvE8k/FOAhyplzhVZngh6hxM
nm8AROFi96MqRNevR0OP8VGNS35hr3mjUMViYywG43PCvX7ODEj5dKrd5mivHk55
J1MblFZL22MTj2+HMmDGAkmtkL4K2T3CleEGXkAl0l/UK4G853U0MrhAbnvqaZmI
tipmagfMw+mzgwArlrXnHZRni38p7iYJQBjnGo5Kf0m8kWJX/4f4Ga08xwdoU9KZ
qBTpacNKd76B83J9jUB/ZWgc+I+Ua5Su0ILzYaVfXE66x7eDBgxZ9yhjIEKyWgNP
64pgv962oFMns3EYXmbkxQO9V3TTr+7Cx91g3MTgJGdgzcBJpHlw4bCAfklGcoCB
Ynj1wJjN8lJKo3Gsm8JlSC6w5xA+C8kEf+10zD2N+qxemaW43yAlrYvxRCsvAB+T
4B8hPbHdW6YI6ASeMolStFZQIAWigtoXq54laM1KS+PNB5eATkuaDtd10gxCcm68
8RrSoo50s7NqQDB5a6qOlc/NJ3veJNKXgcqKfNXStLE0Qhgeona7//OzAg2Tx1qx
jjeJUvcaPK4NwB7HYj/O60cpVE5c6Vhlwy2n46HcXEOJ1XFRjXg+r3A7sFDVoNfk
bIezExBCX/2QoxL3Mzghbv+dRgwZDhHuVi0rfE6u5V1bM0/Z8iDiLwl8KCJqq+iU
sRb7qJsBLDTEoyJ4/jBgxDW2UxxnNxGlJhX7HLoWvEFQAomLqVyCRyv9iobA4EfZ
GL7+P2FkN27tBBlP7iYu2DfZ+edzfvvdknVWB6ZKU9iphHg6NoHEe7LozmzBaGAV
F3+N6sbyahaGVo+c4UzStQH9KArNGG/dNch7AEVN4YkMXaY5j59fIdNTDNQ84TiP
HMxqXA2yDYEhPeaasIV1DkJCm3joQPgO356giJM3Hc8uZ7mcBAyRSNVrVcx/5SeB
aED9zvp0bfdD/axBciDRMfkV/PO1Wg6zwpOPxFDLhPBfEUm/7LLYABAQ3YnDdyE7
CivKzS03M54YzLvl8g81i64gA28c5h5n6gNbqvarrlRkpUoobVFIAE+a1g584mSB
+CBnqhgeWiJ60m5DN+48++ox3kRLD5T/u0kbdWU7pLyG4F+U9rkX00X2b+TKBuAK
F/LC6T7QgKezRr7Ycde+Y2rBkYHWaHyMSju8sL446fssD3Aoqu6pfPgDtURrwr+R
ggV9Z8MXyseHsR/2oJK+d5SfAdGV/ZAlhXksFK8rkbJjlcsCAEYGyyDwVpZRN1EF
KJiPru2m5gZQsfv95sj+gY5y84LjcPGVSV8rHnfwRxRa1sIKRXkMm/ivUhKnJQbx
sF7WmESMuSheh8pob3PUIV8xk1Ivsf8e8QA3rS5AeB4w5BDPeGD021lIlj5oLwck
LQK3M2L2NWfxt3A7jOkcHNwWrCYOkEV6KO0RKjmVlrmiYY7b77kjTi0WTFy983q3
uaNwFcopYXhxZOHslmvmxWniyza4gpn/prIH5vekdsWCqQEzpWR8d1JA6BJILOFP
0XegSBRF8Md7WmoGD43+PYyAjrxaHb6R2Z0PuQTV4Hx+EQ+QiK+N+S8FPC23vr8W
4avqlpFE4goQSNDOLjpdLUUi4jdZfZ1Waw4mpZKJ6/5+gSTHoEr5loanUx0mV4w9
jBPLjGwOEC1dnYaSrguC/jqR7XePTz5cLQzcGw8mJ0kxHxsZM9RDT/+QRZnO0UFO
A9LvIxfWakQ/Gzww2IvYGdPFQaCr5f01UZtYa1jeLltshtYqMIIx1CFl68MNIpwN
V62EQNGWPCF2CthUM89nL/pJrKSo677ll75vrC92UTQXxqjYNRGbbxW+qevpYUp6
0rKQRL5qznO8XOeJb2bJwAbNybtnysVK3uCk60n11rRSM9Vs8vDfgXis7XjNuAWX
tyo2IjNmjwTumNLr3mSdmFhEhCpz8FHzfNf4nfpW4dsSon5WuHjSgE4Vzh1pye4j
Px89qYNYP08ZEjErIh29HR3UJCBRyYPE6faFz60d0xv7ge4GIJE7/XxRO66exYM3
WwkaX+HYUSsYq/tPGLtBq1A/WHvTtLFRc7noAr/Cx5HxJjYm3TyrLE1mnhJw+T9W
S2zUoBoUy9V5NNGCWC1z2MrGlUIZse7UUo+0MWFMTh5wOCtwBOD72byxMU9IBkI/
p3JlfzI4p4NylB7HSy4c5rhxQImC/yDpqJRWq2GMR9cFIy0VjkS15t/1oKJuv+LU
8t5opFobw0qk2p7SX1C8Yy4Knd73ouwGL3DV+QH6A808wvmafGVg1hnSJMwkW/bJ
8X+vVDSkup3jDeVuLMkdGzQvFqZQWciAYlr7IoR2Di8qMG9TvrZriDypdA6YkAVa
cEn3W38TOLvl7hxrv3E3/Ugj3TNDekEy6iwwoBKWZKRErcbrZ57PSDgMe3glXtiG
Rnkj5M4xcOZrTiAoXtfNsvVvCWygHSW0SDNW+Od/m/MwY0qilzlYUUvogfvbFksy
Y9/JhnYjIa1SE1rQCa17OOcAnhFY8HmjCXEXoC2GPuwlVtrn57v0lyXnWl1DAZYX
dh05S5+rMeDajXboxQ0g0DC1Daj0G/RQnN5aBBuqZr0yXFjimK4qnps9yszQZ6hi
86PUDeHH4sgfbQruCvFEj+HDgWwtBelZBdL5/z1fR32TTUQ0JDngAPtqTtUfGAw5
oiHuCqOZS65jT+Q74jAT/nqerN1lVxqmvjM9D/fM7M9AcM9R4P/e1V54QXCWn/WE
d5bCJczgu0VkyzQja4nR3zKvtWGN2G/fTT3Mm9XsWYl9JL3RJZbL+BK3pZihbi38
uJ1EIdYSqMgHhYb2wAk0gc5BL2xVpubekLW2paCzZ/AiKxxla+Wb5UOPyYe5DVkP
udw4Bm1eJXAQyD4QHbYHDohzBzZ2wdcLZvQQXw27xjSsFNvGw/x50FVua7wTk6UC
tABgg583f4y8s1F/Inm5UE8dgPV1DtnguXQrhejphBiULWVlXq/HW4klNVmhaeTy
+tCNKAtS0p+6tbfsR+0zWm0rLLWstTQm1mLKk0so6c8h631MpZkWq/E1d8Io7Nm7
avED9/1XrDqEInS9al5jHTIIDmC9WZVo8Cg603r7jidnFle8H+Dibb+NlZfMEkLo
XqXy1IEtbwidFOL74jU3dayjmXqa1Q/MofpFh6NGBdAL8okfBQh6dOoeusCQRWKp
oTEVn46FDkpTGWJAk6J2RP7CZsiugZvIBLrq8TBoDlSkbUr7AYQhVAW+SAta+ty1
DHt9Opa/B3LL8jcJjB9O+3dBgfupmSesbIx/cL011vSgEZfLTVsG4arUGraZ4sIm
HUcUuDnoptiOU3b4MNoMAqrFaQDmCcbXFlja9qOqAe/uz2IPpPJFA4HOimjW4O7D
whedS9s8cg8ZJE1SbUunozH4H4f/1/web54bUv2OyWZOE2btSdB3ADfOvrEcNdOx
9KEt9MsZPOUVf4ED6PPOnrJkOsRVi20I5NAH+g85QIiWiS75Q2fCJ3j7E6v4Vlgs
AYCYCLRvv4yl8bWjiGEQ8kqsguynAavyax9O9iw3ovWP15qV4yk8AwdK4XomlCkW
2GLLKMAQ3uXsnp1xqLr2AOg5WBe0ooNCgpq/NcRSfGCJHULtMW9B8V5eG26F7hLs
krJ0O5Ws5sj6zvDvPhINy/DvBn9ms7IgxBJsuTRYoyyFemFUnXBeyGlN7wd/e+rw
0ixUhqzOzREyoMwOmTSmLyD7cjoD255dVMu+MIR2k3L/JXKRbkCc/RFQST3jZ+eP
16XzHyREkdPaSONYXCIZ44/xpbnNOYxwcVycs4Mt2Ay7TEa6HPowMJlUgL3iTtNU
PDJaWxIw9WY3Yq6yRJreW/5nKejW9JI/c/7ZBVzTNcwWyPtTdnc65H+JxCsjbk63
AsaTPMaBHpM7MTdPd8rCThr6iyWFJOzpbSHNoeFiqqmxLzL/1Ncc4KuTvI9AOHqq
p8LIjNs/YpTCQOYh+l8fa+7qeoKgYDQM4zYdjNi6BGA8xnppI3QltzVTIoU14+j0
iVgQaUm9NQIZFKpTjizCq5Wc6FWVrmlo6wOQRn0iDGmDov4qA0IOQ50W2TDwlfcP
04FEShxuwmglRwaPGvkXJ89dPUm7HCtoJ2gjoYgLG+sQL5kPccJ8POAJCzXuGoLe
vUt/Xi+Fh05aOwSBinIh3RopZt83HhnxGwEV2qEqWQrwbS3TLynI+yQ9TP8f98Ie
4/V/BG38jcoVCImZSTWC0nzGDbl599tuQqT9cy0cj8j9MjnwHkKJIoblgNG+QtMH
2kxsvepWpSuUXsP0SCBPtYA6n7mZ0+dFkAbkxlZvl6oEL923WuYF8a3BasiUOhPI
ilSv4wcvsJoClhxvp/vvCUTcTgn8TGXeuv3w03slTW5ejBKJDjG2jb8pAEhgftvw
/XYITRcfOmmXQpYJ8am+rcyP6j5+3AfeSh6i60/X7er/CfRs6mQKHHRMkaZRQqVF
9jLNQZQR9m4emziiCEUAUyMWzwM+mBsUSyq9SdZMRd8WHe0cc++lMdkzHJy7WAV5
xTfUpTZa0pJ8q/PmAmuvT+Hl+XoDoEcI4yNHYDOJOreIbCCgjkZT1f6Bex7uYcfM
a2lxHEpm6e3NffjekIdgdh389vifYIlNkVveZkx9QfaaLoZF/QhyIAVQItkFgexp
D4S/m4nwhcB2wNlo8iYp67tjr7m0p5WkELgZxzXAS34peqfkqEMGH/qpZL7YNHbp
p5OU8rX7dwUdcnrPBoE/4r+SZm0hTCViEcCQP5f/Xekne/mRtIiIi65wo6Xgh8N2
baW+KFQCFDtFz6NwqhUcuR065QmKiKfbqWUGVpWdcIUyIyBpbWVNgWnc2PpxBKV9
hg0b7ZLRkHbuAecAp6c932SzSwQfPjcMJGbhBvzKwVuv4Kipn8X4pq0vYrQntHXL
WkcwFrTGQBf5nv6PgH/hZiTfeem0km4pemEMMSCRdF8EyLFqj/2waWCniVNlsIdw
1X+Hf3xZEguzbIsHHO6DUqc+tNAtmMYkmnMXME+KIvz943n2i9DO0EhzOj3RDoI0
UKS7WvBMVYmGuNkb+X/rsoaGwQ/ER+658nbWlCQ7839iYC1/eoVxX4wYLmG74nla
zVAEIaX7F+hGZRKdAQ+mbdLOAcXV1+slZmXqNhuv9u8Gtkwv2Z7mBl7jyn5Y7/JT
8exm1L5yuDQ+TkHp9MX3O8CwaejlFvKmCxw4l4Cfw4zszbf1KLXooYZIqJlaNcXh
4/4d7gZk62+hsyfP9LRMVp0WtoNMOll7s3WxYgKXCBjXZJKsx5pVeCDeA/WyOams
m4XBGzLasHPXjvyhCdpkTkM2W/AfoBnkTzaGHzEPnGWokoN4UWzZIfVIHc/wZsAQ
AuoVotcWnmvA8+O7XmdmxEKQ7dNVwYf3WOr7BXlvKNb8NXZYQzRsFRhz3AdCdenG
8S0D+h+CjfMoizvT+Xt9U8uYVkL4wJVy4vk0iwA7IEfibY/NK8gT2DvgdBtm4t6R
fx4GrpJ6e50iuNCQOy4wREgNT8Et4a8Oze2xkmfUVMrwLb8h1Dy4ILJNQ+58esqS
9IxnbhWBZU4vJWemGpw8l6mo39ShXGZRp/Pnb0jkT3+r3Tx2aqvPwDW9N3xxOauq
bbt72NeGX8ldLdY8+l/rktZin2wiI56fuVSr6yah8KO8P6RJt9oTU61EsG58Yvvm
9TVfLQtok4g39Sxbo3A/WFVCEJP2fH5eHZXtcllLijPaxhNpKjtArlb06nytyK9q
gTKVuJIHsptCWn5Rms/ffMl8gLi86LQfDtSivlYNnVoCW3ji/7YYxjrbDBxBLmto
MCfsnpyrO/FxRXQtsylKD/5UyKNR3A2Up84pI2P82ao8MLVgnYqW3DM84nAl2r3o
Hv0DeoAFAOBmdg02rW3tawFHx7XKAbUd7cpPEDOdB6aIFUmeDKCiBcNdLRy7EtZ8
o9jXgqkDjMbbOv9D7eTlupDukZxvuVADM+1jgQYtN9j9J9anjLPlBYCTZtEVuLVp
uBLCgOCRpezkevN8HXadNV4l8/ss6vDKtgpaI3dQlUUMguTAEOrdSzUqZklGzrQ3
sVh9ng2nLEWkALuhGg5HPt51Z/H1w+3qlybeCfvIxl1FcI001/9Qu/V8Ms4F5K0a
PZK8VPMvBVb3n1xB2nYmymZqBkp7N1bXgkdY8c2z2N855xEI+DBpqIMJnIAelzqy
1L1Nw1bMVSBv9jE94UiuTvCWwE7yn7WB4oVKsuEC/DkST0nbwan5hZVjdj5P+NJZ
7wqlz3gD/6wZ/W+oNLIpczX0pmrV+pcjFY2Dh+9p9b5Rf4XdAte+x13tTUlyq66C
pPSBlEL32icBwiYsOg5ZSF/h1kvzBpRgpugE7bkbL87Ulvx7Enzm6r2eQBnYHb8G
RjY6vsC/KwZ+jrG/Py7ayMc/KloktLiHg9uTJGLILMJjPAONjhS6L2U2tE9aooz/
EqN6CWB1JoaxywqScPdNDcl81qlzxnwFYpgcvmN4fHUzl6GIYzYmixPYQbfYftCx
fgUi85auXEquUJOatijyQX0d0di/B4ClmhWZViMzy26wgGzLuq16Kuagc3Ej+cV5
exiJh2DbK1b3baAyDODRxdVhzglEwbhjggK8V4n40aNwQ8L09S52UjstpU9uA5rL
It8lls5e2hwaPnTjPxDxq8emVLsR3/g62aKaiulpSlGItBlxB9TKDWw3lPoS6oyX
vWbqt9HBLWhPeUSoQiTcthQaitpeuSS7s3CvxlbvMz1n1AUv3zO7CFHzvsxyOd0T
lzod2bpZ6foNPA1qkYP4c4FgHXZTgSQ4AQfzXfOfdLAzMusR4BJ263hJie4dTqhR
OWDo34sau1y1n6AWzCNSBygXQkMmCR8jdpGv5uArdT4bf4jYKotXPim879Yp7+KZ
UcITpD+f0x5SDN8J/KyYyuJv7NPupWKhWuvW8FN1psMzjinJoMqZ6joM6fhCbgVM
RD3xCZBNCHobJrcBlIgwo9Iw8LdkwKuymnyJC8NclxNM4JP19igUKvci/kqftIFp
FuktWewU/qzeLNmWk+mZ6f55flL3/sJWES0YaQAeKTA9dmF6ak3LbnsTDgc7eR/i
dhk9L4BNfGM8WcFS9aAm99keYb+aogv+wpzh+zwEF3uM0zDiiL8M3kBC/a6fXp6i
8/WU/jp7ADsYflggig+urfAHWD463fSZp0UIxHUFsGz0xkpBw/t98IRktXtBX5fQ
vNkljBw6xvcfjEYOy+WZ3JLmWV0GhkncXAmnWiXzm9oYqJQRNngyI2Yw1X4m1rqw
g9EQaCNKjJjFEuSJ/vtF50vVN3xNk0OEOomj55dNjpvOwm04Meokm57c1wGVLXVF
5g1qr3pDzJxaM5Knu3pPH5RZf7fNRpyhHejUlzb0TmBtNZTT4zNWQFzqhTGxM044
eS98c5laZ+zWXV6ZF2WW3ejOb2EmLiOg43LeYpXvnPMvAF+qVFgkyTv6ZYpAkhJg
0N/m3XN7fHGjJIqahu1dqxSP+nZJAcsfIRPWCO1nRhv9J5bHmLpckJOTKWq7QFwk
kLib3ZBS55yhWEPK9c2uLH6OjCdLnCE9r8XT5rjGnxUS+B9zImuLC/CRuRoFCzyV
f7G/eoYUDq7jUcsKFfq65A5WzjI6WTHh7LweMUln32wK+E/WnaoQiOfELGCcl84q
oeBWcvwS9wd0VzBgz9eDL1MF6kX3heDC6kyweT9FkB5vK1EM2EDl30VFC4wQff3j
CSVAnJCuuuacZfh3CLTrQl3/6KtwD6HGzeR9UgV43tY9mjJOO1gh9IWiTapYzgCz
rm6A7hVtqcwPDsTY8VYJBcXeaXhY/tDweycL2DeHnqa2BQFz2t/Ee/SJcgzAbCz8
fIHnGHDvre+l5hyrnZ4PKXfXy2ohjHMILefOfdOspdea8ui6pZYQkwskflCr5w9R
rjKJV/5nXXWWXI63TvwAhZlVsYzMfLPL0a6XwO4j1VGjnwmUdZ2LHyaFvE4aeZNX
fM3ZATdLbHJDcimF6sVWyPgHHWdraLVPKsoLelaYsmiKLyhWUSZ2Lo0mHxUrIJSM
0UcOhpPaXQF0gwAaT0/nOCUYuAwHSQ+WHsvrcX056B0SBbYGo3oC9B/SNZ2VIwNS
wI1vuQ3ZbjZWNL0jCU3b+95FfS32aV6Guka9sbXXnU+phDh797S9t980GEDNVKQQ
ER1vpRVjcmeVuNULi2QA5XJbEuKxzlyRmhdPQW82I6XgS/tx7OdyHspdxy/MpxlW
wHztw0GJ1gfTVsmlnkqO6m+oOvjtPVf8+SV9tzo+ynSYIkuyinUA8W2FauGnmZnf
1M/Qw7hUfX3jakuNL1uhq9W/z1EKWotHPpixZ16K0C/+HjNkkLxtIPE7y4MwFpdD
bj72d7y7KFX7eMamrjDH8g2L2zgVD5n+Q27V6k7VvkyE8o+PP+FWSJOrbRyNcTJ5
A9lC1ZOM5ozByggDh1zjPnpBweaJXieCs3EacG3WqGmtpHikVbDIkeqMQkqAa8wk
0iEC7klNPktfk/vKUBACeqebJKm5ym59nWNgM00XmW8mFN5OeR96OAqCjwIsp2Zu
ypQax7rH6S+17v4q7fDpAFDho/dxdaPNrFw55UbehhdCEBeNGnB8SMXBZL24bC+A
L7IF8lejgev00sCaxqLUZYdCgz/6lyJHNXmlpqs6uT13cByykKXaguhWRG8sA7Lq
PBXDcCIfugG8pAN6dbTQ+jFyPq8l2ZUqXb2VI5Qk4vYceF56yFoq050PAqQSq0Lf
f9+mk50VenPTB29nOCJnyk6pU033YVZsGfdmsIu41nCJ1wrqHvF9d6H6NJ74LFKP
UrPZQ6WIqIwwtkYaFqoWXFKP2VfBHUYUMdLXcJvtBCqROwn74t9hOpMk5yHxA6HE
+clLqQMnLqyYdMU6gal7kiXrxCGFld0SLA8t+83iDA+czNzBIeBfiPQl7TnRg4ro
NSMQfM7fy1XkbXN+hxwOwCzaufJ3oCADWG6nkMP5M6Vy8rzMmdn5pmUj+EMhGUt3
T9qDOeFKTp8AKOKHN7TpaORE7rZRDfXGq8kl/fCL9mZCAXt8fYeWZeHNu75IvOQS
u4/8snLvmQxS615+Cm42LlkYCHVHyk8mwOQe6UQuS3nAUKQFclLV4eWTkQhR3mtW
xY6xTFudoxNb58zLYHRSyqtmkAnPszQ+STQjFoc3dx3mbaKXIpMrl0OkwERtFsF7
Mw78zsZi+7Lta9U7i2lv0/1jdy6HeuvYZis/2dbuS8FkWaQzG1lWKqZaZZlBeBu2
OZWny7yFuRwaxYyqzML5KrVlVW3Fxjgjo0f+5otmTePfLb4txPg9cOOObm5HBVZZ
eNSigz6k//3nrOckTCDu1CcNopWDtN6QIFdyfgnCbC+onF9mKXF/ZP4OGchtH168
i5ZcjGbbPfOfiLLUt9klIRQsHlVMaTdEFSK4zaeI3R4wKcDt7MWRJHxQc/VyT7xu
vuYtO50RzQqk501tOJDYsbiAwdfKNC+pHQh9GmpoWnis0BhZywReerNhGVoWupl9
Mm6MBRCGZqlVI3BElnkf1OfxCPio/yudh97pz9S9nlUTiQEuvWrp6Jbt5gNK62w/
3BAtg1liudaaK+ha4W6jmrxoodt0NiWGWWOGLgI6P9OGc4gCNdD662hv/ItbN8H8
XAXjcMN6LC3YIQfifJQ11jjRVeFXbseOo5nUUTzXqacTKsitdrKBm/kZ7AxFng9e
nbf+Lloc+Ncr0HrSc8tQr8swxTf32nV929baY84svxjvLeymViKoVCVBXuSsk8PR
AfP1sVTI6hv+eck5ulC4UDN8nSLR6O09KoW+Hlwhh7uwf+pox/YPojswWz6NjTqN
R4RpUJdiOYOP+7uKKWoMUYjLW7vc8UL/QaDCGMlyGmH/H+Z/C+uJubeNuQW1W149
7ZZkzYWLX6lwRSz6jhZv5/hjwj8x7rcsEDvW58Tp1jMvutruC7G5v6j86kCJJ/GP
2uz/wAp4HsP5c4bk/q3J7+SdcmkqCdX6ikM4JX77BroI/yJ6v6ci+5nIwYYGWNPn
196BsPEPArFiaWwPYbi/poPar+cDX4gucCeZyZRu7R2E/24AHLnlsLGfOz7Qrtuw
wm+QkzSu+ujBw6FFBtPlsjdn0hY4h0IMmeu1c4Xr9A7RpxIMyElIOBAdAPYSjcxP
GcR5PaxfQ2t4Hv93xGmBF2TdTcZVdOb4HTAdaToyKCly8mf/qO4MvLYfUJImNzqB
kVJq3Q92Ad75pxT3jterdUZFtgk4EPF8Pg2jiZ1d8L4dK0aPv5VEBkut0ATyMfeH
SCZpFHkrCvI2TiwObUMlwNNq+5LAhj7a0focxng6+p/0AM+2CUPzUeJTmiI1QHNE
RhK+3TEPvMJlL/ctPErJpDN40UJywyjvCx/Am94tkB7GXduh0nInpm11NS+ubdL5
EAGC293UMHZf4eNmB54bFNjv0I8ujF6bFxwi9mOnO8KHCGJOjUSsX9e36E2mdWa7
eY5pL8epgcHTKJ0LYZE90FR/cuF/WLF+EVyMrldSETyawLuGetqD7NSoxn0+2dVm
yLcSCgjSsSB8kkf3SuI8eTblqw1IiNSoBx9cQTXKeE9QPaiWc1I1fppe3nvEIjEC
jO/k3V4mf54sCQvYX09MWQyr6DFx7Xc4ItMK2pQiFDJ9EM5f+TklotZ/mspUlxZ6
OuZsoIuwxu9HUtP+lznVgKRhsYfDmcmj+LTPmch8RsbpPAFPlr7mT71tRpfEDigp
QxBfeeURcPuZt4waemnNn0vEqwCBoBFoQ1tP8WWXnb3BnCKu20lpjv3Dvj7b8/Zt
rkU6rNOeiaotkbqf+CWQrpqFt3wEif5YBo8joeEHozCDq4l0vEOE/WqyQg4in41S
SSLkc0BGBw4LA706FZ/zVddy/uYx8+pzKhoWY8pmp06g5GaG1ISHAhatRjKrkLd6
hgvJooIv53q7UVDrcA0rslBljoliubJzx8WCXmTIKwmVju73WWWSTXrKTX0MM1LA
IaB+JUjuRWFsy6dVPi3jAL+bp1o898V1m7HBpndRoNtThwFKvix2FM7QLyA2jll/
m2WbQmFHWvNr+j/sbZILhig2q5wgkBLxicVvMNNwupVJyOBeHjYaERVjHma3AGF4
hT6DrUkzrcs3bpPioDIR5/qIPb/KBG8gHRUK+gXhuwG9WT9jAjCVe6WxDwJ1St5v
RG4whCOSjPKgQt5i6jkdQ2HdoF+smbnCJtWPKtvz42ZuhKdpnJJtiyUyzq7zG11B
QBTMYJGrD1k3v6hsMia3PPICxkFnOnm/2yTcDAeh1A3rPXWRJVCypcv0haqroLrN
rlWSJi1I4i1kTgJiv0QQbi74DOVvSLnQnl1eQL0ncARMSjNBJbgB1t908YC0Jwvy
yCGBDflFZER4YaBakobn6v/HX6ZrymlnfNjuKVBNb6842rqBH2czoOHPWezqyDzo
yNWnz6XagOBGvnNmZe5P3o71M9MCqR2fOrWkBAucj990TkE3gwkABRvQ/D/Q83Oi
kPfhOiK6LpCD/J9j/y4OchHhGRXZDXiPUNWx7rLTZLChcefJL4E1f8o0LoNY4YT5
tsqQcU09ESHoCAmAGa696UmYBo5sbi6e2BdRDXGx6tSTPDx/TULyQkOeq9zfA3JA
uMgykhqlZ1SzJdg4IRUXe/KQsm1aslHdMDWbdswSt0zQFUyRX/EQhQljhuLQnKk7
AnpH+Y6sFi0kO0687Tp7i5uEr2pkWhHWJDKX3XnOxk007COfI62GGqdINRr8wvI9
tWoHp0K+nWqWtWrN23dNlMoa0/9tk6JoPLjcvELw4SkIR7iiYH9DaDoIMX8zJSdl
XG/q1qpuvbRfM73hetS6mVw8b1IDwpB2fUlIDD7IhPm8yG9YcrLqXLOrg4gq+kA/
5DYXQ/5CPHi/DL8kOXp1U3uQvg1vYF5vK3OnGacA6aohAzCfbZzapM5YQz+9R1wQ
FhQ1OcJfwt8UYqxBpJkeQfAeeq62n8soVB8dE4PcOOWXu7Rbx8tnZV904wBrOIXj
TVHkrEDTejlwVi3zBurae9Xby+Sb/YR9evNu08XJCTVqHjpHbcu3IFc2eIXoVhCc
0UHf2hDQMdRwJKYH4wcJoin0VmG5mXUfNHuVoPsVtkf6Tg1T9jbHOOlos3E/QTKF
riyV7Fm7OJMwM16CLqpc3+QW69dhkVeI3D2quElGDggAJKQK8Le/5B3TZYkbfQX3
xYfvJACu1MfS4hp6yLlkCarZ3ges8y3kvD+Mlr+d6lH5JSv3c1qptNIiUXvMp0GY
+OKMYxkG/trkTfyvzSauBet+5Ww9y9GhyM7p1k7Z6AApvGg/BkE93/wwJisUPPRl
oal2/Jcjd+8AmBU4eXNtLD1x7FhFC/GaWFqJ2BBv3MrOehNentR1c/i0Y3FJbKyO
Icvuiyxr88jWiufA7FWrUkkQKq1GbnFBZhMf6G4U43HbZKV+KxwOi+RSVJoBry0l
UeJWFZ1HYDn2nL2pF1amYX4PKT27phiV1Bgv25eAeJmE5VmPZterad8H9O+pKgUM
YfYqJB2HRp35eZc9XxjbCNWVPfL+6ADxS33cmZba7N5uDqEXiUx8DhVPVG/d2qeE
SRZkwgA4CrgEAPIpvC9bQz1uplYUYZdHr0q9yxruVoaFs3BTcbyvJkAOk0hVzUaf
S3NtnobA+F3taY0SfF+/YAj1X5lo5cgdOW5p67TkCHmsuyxlDyz5KQDMMH4Qk/T6
Hf9fq7tMhHPrcMuiKSQqBdvi0QLdNaEtVTtiidstRQcss6j4Wna4hvWgI9UIgxAt
M6mBzq9frdrrKBSdw8rUPYc3kZxKbELC1YjpgooeiF8r9Iue59Eh2Alypg0ktTxe
Stsg0jDMUzHnNNlOHv5iKm+1FRSR8pmKprpCc3s3zQvMa/HUidZj5RhSSmNkFAUh
G6wQsGVS/fT39B5HHxiumFs/GiS8Hw6xOZFx7ecT645MoMUD8H7DzBHTN6h53cNb
Jq2szXNae7JB23z4mb8ODD/5YJrGjNXdMw0dFn2mzijwryFbYoyY5tf1a6cCp1ey
En7OkC9JGFkP9krEru7aYvf92/f6VQGb+Al86L39DyjqwP8NVkUDoxc3xERfOFhh
V3lNzXHPP40WN2mPpPpCGBCzCKbwnjBCIYihtnkJ4okmCpu/3BAB4SwwfvfIN/Rm
l/eRYrU8Gt9M+rc+RFkjEgdGzZxP8cxJfiPeLl5gTTOtWuTNN/9b3Se2K25KcnBu
qflXudn33fJhCy+zjjO/f5zAGx+zuSVCSPhXgF5S505gtxQeZT1Yy8Gyg33uufKL
JJaCb3vxG834yDm9PiGne3MJZqd2PwdzO0HpCBr4xTTh3qNKHCfO5vvZRZ5r4+gu
gwtqQ9TZHRYq72Iz5BFymDkr1IZ7HNMKAgJ+X0GiVU9m5+BNiBp7G0UtfLb1Biv+
EcWu8S570SEbn+c5GJ7QwJyNoSElfMlX0/6OvBopS41sJ/84V2CD9GFWxxuIsPXF
3sbawlGOm3mK18Utb6grUm6JvpFR4E0CktmZyuiOJ6Rb8Z68vo6+MoC58iO5TSLi
lwYQ47cZgAMx3RHax6AjCyS+UU40DcPAGUeeRQPjbacz38mtxvjE7DMn9Mjwxr11
4NATbBmzXU3/k6SNaCG5fQcz4DyLygzIlwaQHO/0v8ZMQp8yu+sIvXo2o2jMkeDD
L4KOZYeSdpDmO5JWXRfE67eUVvIE6oYn0kWPrPrZbIB0X/NWM0PyWfnnbBuomqYn
FjE80AGnChp7HgQ+1JJmS5fLxeIqWNmuN6U4+Ulf2ClmJFKX8vEUkWba3sfTqpi2
EhTCnFuft0jeUnpq3Xj8xCnpNvWJMpGRIehFkKTtUau2NS/nlG0L66pOrc8AjSTe
UojbAuNzSt5NZ7SxOShl4m4HCZ23kOIg2ZjGH9TmPUn6sSp9lMC+KzKNaSzumwYz
HCgqhL5joJpvwiZjKm6tEfEwqrM56xINn3dt6j6K+L8/IacZCLIzY/ZJWqp+YEOK
Fp9rio0zID+QJ5WmutUtywfb2UG1IfciVD7b0vLEmPAtQk+j+b/1hBlPymn5ew08
pDj5WgytzqN9I6l8NforrdCeNgsQyrumVi/Iauo1FMSPh3PxzbEkDyc1nQfZZGvA
393/3ob1MRdm6Zwqq2EALYqYTMas6f2b8I1tIs/WCmAhzJB6yfa97N8lwh9LiutX
9c0xSgIUgywG+MqLVJvAPGUuOusuzHdVCVTgwvha4kzOg9OrNMJO8ika+E1uKQWA
AaP3w+RP9SpwBm5tF+snQHI8+VbW3eFxcbzJqD1fLnMn/jcC1LRjYfOHZlfWjD8c
AdkjaNp+kuxM8UeXBNE5Im0pm+3bgcsANNH2tS+igQIy/LpyuWj3zs/XCnUypdIz
yQzfXwc8HX1DmQnke4tO+Zanjegkvk656k7hg2Ti7U+HBH0Haq2Gx+L8AX2pNber
xI4DD8Avq3U3xD9yLNh5O+Sqmlt1jR8zQmVzZSj5LCFoDrwWmPaI22gpN734WxjV
vZWNw8AB4NMsy7PBPgbZcXZ9msbfY7+0DrcSDjkzpcpdRauFpzecLer2jFl5AeTL
/4IawtGX23Vl2AO8hhHDxUUnPTSKjTDTL4mM2ux4A6gHGUNgqC9NNC51Jxz7qL3P
dUlneYyX60jeoxl1MH9HRa65Z2YY5kKy22fT4uWEF04jU13fUJEn17q6ZJEnP76b
AnwZzUaLjQ8rb1IHiii405tt4fo5uy2KS0ux7w5mOy5tkF8mlikr4nqDi2W/h9+k
9itg5q8u5TXBHHR14cwcgq9KUIT9YQt7NdhlmoUSSNGninJamon7ERRHYqkxrs/S
743W8X2UxGvxz2XjwkNKVku15GCPnzeoiLKZ3XwBnGEI7uLiARm5aLiKBZJ+rkpQ
NCstWBJm4CMzaoQgJCAHY6QOqjRbfqvaaPsn84leP9fLDo0bnyJD2kbTJyEdbF+N
SnMgDYO9y/l/kL+7EclL0grE9kQbIpIUfDCvtNrru6P8lVZGmq49TBBbBkad60rF
xvnIvQAJFab6FMri46yWhw34KtoY/tSrcbLFvHsz/m41pRadx7WCY/Wz8AyMPDXM
LkPsmiPhrmPPonZbT9a0/zlFpZctEgqv17t87kI/vYG0PS1pboPO2lwJrhLQ5H/7
gpITr54eyvomAVNH2REEdtg5edQGOfnizVE/PSszpcZZbux9uGswwuHqMl7HlW9H
oXA803aemfmnD2o4fit77Y+Hpuz5ayXYTEFEiILnjXBnlczCG8mm3mR+znf0YZWZ
ZVDMXUYuHAYWYKGFUptMuvUTRUBeClepvBaKofgydlwS1+7pJEHlvM7GZ/lIGBvX
qCwjzV7PXXGbgM62gHyhmW8Mqe6PBEBKj0G3Oc2HaEwfct/cCzDQkqI3eY4iqqAF
DRxTlCBw7WU7AtHmieaOM9W4qfP1IbhVEtmVpZtgHwgSxG9Vjvqtqq/VgWqT8n+A
sVMO/t40lrfKj8oKCjp0YU0WwJbAXgVPMkB5mgiCZu61XSO96QSr06kui5ImsJTd
MNXvzNv86NYZhlDvvVcwgRhvwcFTdRyTGwV2zXxn1OZ+jAGGtYdybn/6HoAZLoao
YgERhlUYFo4LbdZIYx7X06KxblwN6J9nrIK8QcJqrf0uIR7IVmIww38cuzmXmS3M
jrcONBVJ8lkbqYEnqRPW5gjYAzMtCDIWax7b6E1AbffGGJRqI1k7pW3X9Fs7KULr
mLAnPA0aaJq/s519eYQtQoUYcqh+A+LAcXbvnDahQWvKfewYIGsxbnZ+gPoiDOkR
LKD1pY47+V/W9rqPcwva2K2LR3b5EKycVM+AdNrHUwrW2zRE4p9k7VOl2M54t+tn
vk7KvWAo3+nyn70NhZdSbkoDUOy7oNBIs2hhb/8JVhTcaIwSz3UZfhkK+nISZjbm
LVfs3CqQvjy0WvAt2bo2H1/sqww87mFmLCTW425UIHRlRt3+I0d+Hz73TwfeClz3
E0JEB+8Tue9huuRg68LhgajCErQxpDrU5EUSRju1nUhpgqlDplhBSVsmWXTkzO7V
bg1rY5QWVnPixiLbAR0NuWpvAwPdOo2MMYHWZ1PLu0J4OoEM3q+8MmujG8If3fpD
PPMQkKPGGwrYOU5plEU/VyKtpmFuyJape3AO5+jCL0OIFngUF5PlKx2xXubYEknO
du10GVip1Qa1BuVc362qjxTGc1Ux4+Gq/tLd8/t0AW38H4Cpk6/Xy7m9ZOWcOnJt
NuoIxmK46EDeYNlPSMyueCM3alhyxBNClROsh/QGGtfk9LgBACn44qwKaXIrY+Aa
9nxVnxHawUqPZGGz3MYpoJxi8m/z1JCsU/gW3s2QpwGL7FdzkIKv3Li0okzrzJiJ
JOUcY4N06ieFhun1WbPCbeQcLwI080SSBmMUJSHlrs9EKwW0G2oxL8wGqxpnzT/H
eTpccbbs5VXXAGPYcOaInYqTMbfjhyquh540KReUep3NJ/TYgQ5euVfKuz2BzUXE
4c9RQe0WF2x18LD+i7FqYv3FrlcmmBGopPtr136xKgO0kjgiaOgoefHEdSqzKpBC
CCd6fMwVJKhv94Aq8U8ytjtUeIhIpLysEhS6gUgDRHceeGgsIKbbK/XdMYoV/VCA
szeCvlSlf90SBqBGwMVNAHdf4NGK88PW2X1fYVK/b1X2H87dI3G1SVvIHtL5kWof
q+OmNLf+7NNjE+CJEHjpRHXHUuDoZzj1Tqx20vBCrC9nNjOOa39/6ZUn85W1YTSd
LRxigzR/P3x6kfgVRZhpYgbxNvzmp5yIlu4ZjvUtcFWn/IXyoQLcqL5QlkA3UkeT
iO1XBOVsvEouBDhgOoD0aVC7snekyK8akOtZ+5ZwFdzFMb/eWkPiJGre2lBzK/kb
fu0e97F+rXaS+lHg0QECJQ75k4agKDB7l2upnoFfTrRb6+gKrTI8Em784g/qg7aa
y7m4cG1M0XCNjmuo1wYndqGMz0I1zIPPT5W4J8nU058m7z3iOvifM/MLQz2BFMmH
/J00gJNpYUYZLUB0t86FKz+t384o2nZ9aK0CE22snEXoey3/FCKoUJsPLI/TEFk8
oLjHRPv/xZrOiam6BpUHiZ1R71Q6FbHP42BusC/xJrw8C/j6bCKZnIqKhYfbaC1w
vWsWyaPiOvs2jvoSf7uqAY2lpvX2DojDLb1Gxwe+FNYj6+to7n0J1HRy4UPNWUfj
cVJeSnXSd6Wb37oLHpfAU+K7GdIg8NA6U0KYUFarMOw0fa4gJlZzVnRixaVUlrnz
5ai8ZL5TZPNyR3Hx87eNdR8h3kr5cy+za9cNBXeBkaiFfmLcg+UlruVOrgzxRPwP
3vkA6uVsDVRI6qnJcj/GyeYloB9HAkajFhF2Q21KbOBOTT2n+B1avAkfqNZwCCe5
23qVSm2iVKP6gQ1V4E/apiK1NuoCA/yBsZnTJcOxw5KtToewpt4WnjkTuHKF3a7A
hOMdZ2Mwf3Ppf7QpdUQmD8ffqJEym1yGBopbjw3VCPVniLGvhOmH/W5LtZ4j/0a2
pZwntYWtFHZp9YdslsnqyxpjCf9phzkU5GfHympE0XfFZr288brOQ05hrnvaYBj9
1QlXLOXn9it720pKUmWoWpnpxpKJFPNE1boYTM7eoF+oQolvsmzaKIr8T7TSa+uf
4vKnz9G80odLJrErbJbNculd1GVVx8eqwWSD5jRi2yHCvuruFSrjJkDKULCTLMss
APY0hHPTwvbu9HYZghq9F8vlJyCSl5sxkXh4WTc0fki77qPnpxAUcu6goe2RbjUj
EvA6H6I6G3NaRnKSRHUbriIrJy2RBOrfzIJOCgmcBmlOTTV/BlSz+zzRW+t7JoRF
RyZlUuI16fjJlxowZaRjeWiCoygoIZAeJ0LbDHQ7X8miwmFhiVNtowY0uBXvyqbM
aLdhq9oVuUjcLqhYQ0x1lGjN3opwZloGmPGBS7fvOmzMHP8G0zDPCeUKhLexgeas
hU/fb5Teg5hGEW622EADbuSMdMtiFikO85rPDjy3VVT4364ueC6HhqAUtaV0wyLE
ABUXUFjeoo09tqBW6N2b061uTUyw6jiC53XKctS2/DQe0U2LfJbDmiEb6vgo1Rko
0o/i2RL/peKI3TphvcMDpNeR2AhgXA8FEoANMOKcZgGiCzPRIvzEde6i4giYMLc7
VSypTRtGg+ByVJ7qeJUE/bb4yTRA3YqLxLssLz98IA7Hq/GqJg5tincmZ0IDhdL2
lmJYO0fvXyKnlFr14UOQrm3ZJUaVjJPS9z/ElzalSZV3hdUmmyj1fFRcww5I65qp
V4xPteIWu0uaNovJF5Cst0kUEpPFibzSbAUvWUzwN/7aE1AaR6i0NZGoy9Xko68U
w/tg6ozZbOQG8vOTJW6U2Lla26HQtnfwYnKi7LbJjYkUjAtzUJqXsG0Ft1Sqr1Za
WKEfekBIeBceKRnF33qP+Sl4eFjAMMvN03FYqaacatqmkWdkQ9xActdhb9cGN4U1
+HvHSIoVHdeuOui20oCXTDGJe1nOwQCuxSkZXoJnUuLNz+MNurCoWhLrEizMTMMv
22qQDxi3+6KWEj+kFjtoug4OTd+3Vh2TuXcUqyg0KMByvKaU6ZOyirqBcNMdO20P
C0xNRPpIN9JMxwug/MmPToXiHpUDxpL7dnigHK8mhwyMxGezM8NI1YeSmmzyoV1Q
eKjdr9cX2t9HWmNqKTZBGTkjQZpdCnM/kFEhvie9f3kE5p58zBbRDI1MChBCSQb9
4ETbJNEDmCFwoFs46Vq4JoS+BwEHLCGHZxL5Y5GnnO7UexNDlxrwzzzmflh4i250
xadTQNuTbi8cKu73z3mlZLe8mRn/1kxGj9FOIDFEb2vrwkq13pLL7eKs74jHb7DV
ka4C+k/gT2GN8V/P6/RkpkBvp+ORULaYJ7Kq+0DW5IpdsJgbqG/OEj0Ed9JP6xxZ
UkUaE/rWZ2GTYFIZzvEQwxeU5Nmp4e/z1sL704dw/1gbSP5zFZQGYND//Ykddcur
1P8hE0r8efsUV63+s4FGV65V1P8WKYWnjznTR9s0hFu0C+8xTpGT+ZBxHzkzuLjt
Na2yAZQqbWTvLA7Pd33DCsbvHd9YpAImG2LytR8bgXjBgF+I8DtIC993w4Cp3HBw
0Wz+JS5bTYR69MMgemlaeyhnKlHfUfJbEWdRKPfolXaGaK2Ns73inpeQWVjjrG+G
w8zy9ez7OINE2kec4FCxkvaA00uEM+X0fKG06SmmiTpXn215kUIROgYkeucir5KB
w1JrMXdWVwyx75E5MWedkm8IR+pryRFcxo/GgRBQoz18Fl+vzjqZGsm8SRpqY7p2
01DGOALy7bs0vYp4x6EWOpH1zPFfpJ3EynLIGAeITA5jakiLV+08Fm7CQ3Bgevdq
yLoawgPRlOVmIpLP84ccNnO9bByYF3UAunzonkJ1uq225sgV5Ty0OP4euRut2tbG
WJ4H0cEqU/8lfvShrgfIfEWsm9mOkU5wpTTZC/vs9CfffVAsjMB9ZqySv/l8Mo1U
p/EDX5mOTVtF5XdsT0LLJm4RzqIrdFuB0gDoYvvHQshQNtu2USA+1gCPbpv7LMRv
Q3hi9QDU2xYwAaD70+Fl+hVKVQc5v91Dg4Y5UmcZDJbFSTQqV92gjfLNI/NXVmoE
bXUiw+bPj5OKUevc2CZ108G/lkp8kPN2CqmjTF1k3j4p/fL0uega/jQ5+rrNSsx/
8Ao8mGPokL3QYLVmJv19b6NHuidorZ02qjXaK3TFGxA4qlSEG1fb/FBW1bhspeGL
S3gMtKAt7YR96O9r8qPqwcZ+jU6dYdf5trPvt8RQTcgtquGUrROhc5f6nrqQNmNI
8WP2wTToB1yl1iIL65Wz9oSHAk9Ke2MYCQdKTrURC+WPmtGTc1oSr9CqZCrHQM5s
gbNeKC7ypzQQAohyU0i7++mnhjyd7MaBSI769iTcd98M2vVWlCx4Vu8l+V+EZ/c8
vjtqLTLi71gXNk2sCGDXAEPWzh4T9ZxuzLltZyFua0b4JAUtsRWSHlpNY+0/ZD+u
hYLlE6YP11SLAmjhQknMuQGc9DEI6ZVSGaHCIqCnYlcSuplGhTZZudDBKMmD89gX
vr2B9DJLmadE72CI7gLIFbXGnPSLAzT8YxdsmupfURPGHE8xI1H8UnTuaiBgpMhf
w1wdL0qpTOaqMFW+rZX8UL33lYqdAH1k7OMAmr76P8u3NWXJjArAGPtL40I7Q5Gb
4qbs8PhLzqfTjchMlwGTGx5tC2OvBNAk+wEAlY0pjnKOMYLBFjP0HNzuGLmawQzo
RyWY5nCuzwPOs6Pxo6Gb8LrPKjMuq6MYL61DlJApHL/UeqlOFywAz73F6AxAxVHN
eBe6lyZJk++d37/07mZWt+Z3zKBvTW00DGtH1N1NmJFBK5g1arGDJYL+C7I0mXBm
I0cwwKApMmHH2UJbGQec6spQRmGp0LDRhltHEpdUy8sUjhJiWeeWBUTz6ofO7d9+
DK6kEL8EgeMizgI7wxRgFzrKsSf3fs/aRceYNcPl5ykXrhWuncz6REtRKlc8BGCa
RiNEV8IfxohlT6gwov9inTPRhVUmo7aSJZDMkLTufwk3gOA2KZNrFPhnFYGrLzkB
fIgPhRxGpIDdvnAqubeaV7jQVmf6266xkI6gMGZ0MIomnK/lHAEqpepeQ2hzdNyh
Jib86LOvncJS/fqaSHOhLVsP4oMWnQO1OboGXH7+3I+/xyDalZ1J45XTDwAmPlwu
dMdtTnVXRBV835rwP1/DnFOGwA/Mg+qQ49f/f0epgeakVpg8tfH1s2tl51WLAinZ
3shrQszVhvn/NjfrGNg0EvXR/tRMYfCIJfsCPrhWOnTuhFpPxtZM4omy5UYnl8zJ
C19MvWaVwKcO+S9ddjji5Vczu4w3MJskMiUn8xz95a3C4r76Qa0uRIxGON61a8lF
mcNg5YFRoFgWokZbF0uVtwGJlEirf1LS8bDCsk72xlXMxv7drUXVrjtdAKWe0LHX
0y0MWxr99W44iZxMo0GJKB8pwX7Y9aaO+aHzKa9JT1nnj1PpMuRxMMG2gZ9MIqx3
A4g2O/ejEtkt8003ACsiwxJNu5E5f+7EIjSEs/oagbIaKED994+U+ZwWiBaX2liP
drUuqgWEji4TS+b3XkON4DOgFo+tdn5t4XEbvciCjZ55b4SMKzmMp//3rhgh+fDn
8RW/nzFzjDNiqOW5Xiu9Ku7UdmF8Te5Ej44YmtxsYs0dCSAQOjmjOgeVVaCg5/VY
E7EuYd7jEvg3atZpk6u1wcFpz90NndPMr2uHVY3aNXGdh5+Y6KY+jfcm9DREWypW
OMS1rVM9SbayWYa3a6Cie5Cnjx2h9ftb+7yovoC0qCI/6eNZ3uj26UEnhbmz/IXX
lVmpboChR0yYskkjgJ2lI0ah3rzcRKf4y5bzgUXRxfbX0iHl5Fbq+V3MwGgD8G39
XEKttLgg8FHu39XyovOv9KeY/ecQ7O1W+puU9uA1cFnBNEmTibUhm5UmxUA3PTpz
NN/8Z4lkj+aXpsBygDQVZNXtcLc7zbAgp4eq2iWeiiQxNnyAcNdWJsoGB0GLWe13
TIseHTUGUcnBfwRlBG5p7hgzyasn7ueb5fxHjXuRjNjbfmAa2ZAyvias8xirCHTV
za/zRjRc4hp4WkKvJrteMfQ3PpDdPMg7WJTAUWplXoq9NrE2w0fiV77BhtN/KIZG
lCMAR1wCPfICpeVaW2puXmVEcRX++YUbShScWK9cnxOg4C0yI3cDBujXcg5G9QVJ
Oc7JiJsvcQTVVinoYpQkyTfzhMz0R2qPI4w6xBZ3pi8NTjhRwA5PM++1svEbHQW5
mGN244ARQUuOS+UJwGkO33nAQuGbhRukw7aCJrsPWx2bYyBY29s9nQsE5yQeGLTT
zDmW53XkJ+SSRLR/OYWzvpetUh+qRiOLoVBncMbyPd8sTp8qUtFT8QZhP1VE94lL
iPZTZz/5ULuALvGvGMzSI2jyRvjkC/Ntmdgp2O0WansPbGZsRV8YqA7JPfv8Z9Da
/2YGGtGLkDCy5EUmKWuS761fMYkCZfu1XMPdp8jjziD2dsFD2528bBU129A4ho7S
1DBbMTvV397R93W5xJbIeJsDRCnnBlMFAWkhurBEMIQB2/Jpv2kb2a/oRaCq6CYT
z2yHUBMbdsNM1CaDs32JrJxLR5iq0BCMw3sdiKoqGotzEVPeVPEJ1ULp37VJeUF8
u+YKKSSz8XAmeJa8BKYc9PXD+LekTja7I6TyQrAvwdepbPGic1h2vAb91MR1+Dfg
gv/55+5AyoyT16AGFxRSGHVZ+IF6Xfbk9LCuwLGSHMsMSSszS97lhFSsPZZzvDLu
KecyqyuzZGofN6/M+x4HMczYH5xcp20JoBhwoY0SvG3QDC4uy/A0LCyUgPgjo41R
JR8t4Si1bZSIyZB4IweV68iSjIyAzwoqd7F6JmHzT/iVs0bOF9tbHFX3rF750nlM
PkNS8HZzMOMFeBQFmQpm25ei4ik5H56mazVB6va53P+MIpBhDQfBi5lL2hlSqzqE
95QtBv+Sqh7AcfQU5pitwAFSAS73o+sb+bsiIDv7+mWRaHu6bCl+zmPDvn2cgS2M
V214oAXUmtWGQ5Q8yu7OWtUki3w7sUyobArLW3gH4pvFnkokSdU6LdIZFsu41ebf
i6Ih4BDKjuOu0q9RcDQlHlb4U6zDp1dSFBp0ibqv6YWd3r5Wj/7wmiJhfGxS5Bk+
rNLC4PXl/dZ6pteQOjtqi0p5dinsyW9VVL8fsccGflr/7jAw+MBwQKORAv5WB+uG
j8E6RANUkkQIsZRcCQy53ECk0pWmmhG3SWE+awTuzzIw4pqaK8l7ELjtawrElu6B
JYSnzyq8HsjwRYqjJPOx3SDiAI5GDZ9bPdMfIl4OOEN0+cevDNvcIo1F0qspyoVr
O4L+8tM3LHpHwwMJr7FGg5tIhVRpUgWYDRL8cCYoZ8wUnV7fULa6gOWpFtD8DfJo
rrq4tBm4Ndphtri+EL1bVOm36YNb9P5L3H3ZnLheJi77tnRWPULxP9zXgTTVdj7G
bnpQXp8RX+uBo7XvIkgupilmuw86b+aK9Hx4oz+Ft0M+kBP6eNzpnFDjr6I/y8Jh
WQe0ug+Q1954J7lpDkcaK80U4ZAs7IVgwwxhC2sDqHnv0sOQfyk5QAG+808xJUji
/uyNW5z48sG25K3arBZE8rrV7hlSF5x4tNihTJzLoWDJPPpDGAzUyHQ9oZIDqibD
RsNMUoOnZL0uCbUc5TJafsHO/F3w6YRQ2M/6/NIqki6JiVJdhYAjzBOm6RYjISOI
cKrqi5hfHXdD5CXfE6YzvTZBZsWAXU5+KESiv8hz/FJvnkf/ArJGMSDWIF5jylZY
HJCMCUNbiEcH9mYh2b1n4XYvOavxT+JjszEyRsOh2lTNpsu6ZApXlou4UNGxPeJN
cluZ8xq08b7IUJrPAheneyEG0KLrogdEFqB5xRiDKZfwUK2RgCfyNNQL3sNg89Hf
DKS3o+9KdTI/1sTwkVBYLYlBL2paTwP635pdFls1ZEcNw++ibY1347ZK4tlkJBQX
F9pZLWBze4QgyhAG5gaqLru0hx0m2Dp85UOZb6E4jM/ytmB7shyotmQ3Srq0oZxG
sexxmHmnzYouMBzp1R0KYq48/nhBYt0dPGlklDEif/DFaLi5iuMEuUrz+rHMBuvH
rBnSMWfx+nwoxSOIIJ+MuQhMZCOYBpb4oSRCGdV3JAcQcIEqOvIQ0/CyZHgyZ62e
r6/hNsBHYTs2gLeL8nD/8odfV3yb7ouUmAUAfoZvyKqRwErFWGk7eKmihbII8JYx
CBd1/sITzMpCwCughG2eZNrau6Wv42IQh3u7oeS5UZJE66HvQzb52a9jmbJ51Tht
w6VdcL1enuhD7ROysXKMNKeZuhHBkZrBToKcfryeDv9mvDMCTeHCGzUqxNITDTan
J5zYeD4nCK/J3l6eJiroSl1nv3pE6WU0tY2DXg2e6a24e9PijHNxwESetui0+kj0
4I83afAkknN0jdfn+Q8y7xJKDTha0nx6GuppS4CfkF7jxbElKHLMu4lOtzVeTi9f
KaldfDVstPmqbrbWeyJi8n7TzlFcrF3h+hgllTF3Q6vk3ojyuhgB0sdr3xlIQ9I4
A2ElHUaAL/MLlvdQHJwwn/NzWTHdmIW4TWjTG6Xb9qJGGvqdsA7UdcOKLKH7kQ4c
57tAHM3/Hd/fgCVFLlONoO/wTcWRrDLrv2qw4RpyEdXRW6mPbJzbqHmGPGRxcHQj
wEgQA+mTvOovGt1pDm2kX/TIy/ChFi8QSZh+M5XTFjl8s9MLG+yeIXr69GjBDJ8p
tH0O4zk+uYWO62vFTDBCweKrpq7KaV6ZsNBOqAIBkR11BZg3nCSrxpMbJcWetS7v
e/5a1VbDyiwt0Djg1kXkuI4sez8xi1KBe2gl4dvH6Zj9yl3qjYdb5zuN1luxnbhc
VTaUbVAMgLUiYY3N+/7wTqT/FHw5KiF18B4HPcqGHEEIL2fA0G1Kn9vlhuLtED3J
4Iw5eGXj9EpXM/nWdrx8i4GO/Abco6dhfTq69XAbOEcSJsBHCzsJo9NeuPoBS7dE
WfYd01xF3ylU8kZGPvVnjc+3XgP/rWaeMowNEhBVNG08yP8OWJO0H0rTKS8fL9Ki
A+NoZkKO+u2bzWcpPkl9rfox8srtjHUEP3L2uDaCrs4gWoDpVfDPE39dyHdkaYiP
NChL+L3/lmYVmbLv+D+At/DbW7m/27aVaNRUGHEUhLoQ0BY2KbXopWUxLOj5Az8y
9ndUfbvAl5Tp2f3whJ9sgFveS/ygvfHrhQHyjQbT5i55CpXvu5AscQFes3E5p/eg
+ISWAI/r+LezmTl39WiK/KA5H0Vz+mkHiOm8IaIqycEf8AITmP/sSIW9nKArv54M
0yYoKFoSA82REXhjBMgJe7H50iJvFzE5c+xG2xo+jjdi8ONIpqUUyu0E9K3K6hJo
9XgAEYsIFIkY/eURUrsl9Iy4TAh5ln6z38BleiT5/Z4WTbAUnxmaHNNv2IkQAvbk
O3nUxoa2k3bKxZ71NxOVEzRNwZ8HqMuhngAc1Pr2ztp4iKPxEUTejXnhnVkx4kOk
hxKomVhDl/frfJqKcyltrb8LZVGPwD68t5UOaxHU74F4eVG7qA6klnM77HD4lFRK
ECUebtQIWna63UEgDIGssDOCUBCGa7lkZTs21uHm19YYjYUERHFcaTZJ5Bc2H6dv
G0s0BMgvBFqXKtZToccb89zoFctOQVOSzEPKGs2ZmPt0kzR+4Dlb+lha0y0XJmZ1
j0/CgBKRl4dO7InGJX7ADXhhFOzbKGoEPfIpK1+Fc+dadIfTwAv13XdUimZdaBKH
bIwwHzACpOye2lQdeYxEFTKnX0ib+xMGX5/tT8H+DpEuFoftWweAys/wXAL1RKwS
QPb/YQFoXLKVI5ZoLdbhVSq/vIyEXfelZb/sJSdcz+sKHDOHpRNtqQ6kwZyhcrov
ev8KPpYHOB9SEb+Lfd5Ld07RVcawQ05hY28J7RQgnNERq/vtbSfs8rqZiGm2653F
CgCM0saN5ehDoKYqHajk32wTqvuAJyCxn+8Gmxy3qk/zH4+HQA1nq5oWHbunlu2d
MIi3z8zXSTLOr/SAJaWSjI4ygns7ch29FTxGdSxNJhT6ybmme0bne1SdBw7ztQVi
q5x+ZntuAK3n8V5CY63hpqkEVxZ0AwSZ/ZrWHcNXuptY2+XcZtHcbcDJuIA2Riu7
97CbMeOHUSuUCyXL8IEA1uElQTH7jmTLt5K92Ck3sXYgea4DRnSKkV4TmOV/F2U6
FdKjfQfhYFNIdGmfve3wRnQ+PLAdtB2W/lWjhmG60p/NB15b/KtD69BYGv4Mpfky
+4LlZg5D+vM9nnTe1rxyhboWTPaPbEoeKQVqB2yoOxLqJuX8wYTd7XGViznvS2tf
MxDiUanjVJlYuhvg/nyFduuPHf9dbpCkZUPBccmWPAD+Q7s2rCiPZEk7QYbwuhDH
ZDmVh7hxf0oi64UorEfOC+3WWkOr1U6tfWmNJkPTdYX0mXUQqqJvNfmV2k5Ng8h/
tps8Br9TWGnvw4BK/+5OozRaDLg7iBhVWefocgPZ2UAWxGldBUuycEW3U8DMNuPU
Xg/KNQAHCrEeeV9aE9zH1+bX46rLE49tLbgiecZfQ+RNCy+l/N9U7gwjBdgBWgnV
KaGv3x5aKSOEQbqVu4rEIjRcWkFEPQtXccjLHLu+n3JIVPkrLfSKdbVkh4EnR/sG
+UGAObT+tNsc7JphsCEmAkkIihFw5TqTDxSCqXAr8kwxeX29Es0l/7qg1fhSi+F0
yt53D/sSG7DpQsCoRLNRPbWTJni1ZVlMwWeG7CB9zmY4FVIdSa3iuNalpx45pnO5
Sw/GxoT8AEs9kKeuYsgzzG0eBZqWaC/q7Jwwjeom5yjtGzDEynEAuxBm/ef0rynx
fVHg9rABMmydhIbqDiEiEc4XddWb8KxZRL04L0CUQC4TY6nTId7NlkQFXgAYodJ/
lOsYHq62nL/2b2fQ93hlN2vI95t/t+aVgwQf0MsIKP27lHH8ETHmJHdC6mqAu11Q
Iw5SS4z1sT/xSncLgnyqwKbfG3d2a8bxAJ5AU6MxsUU9JWhLzkdrZv6z6HgdMbE4
Na+xLk30hA/XARpuohS2JS/nZXfEVJyhMZXPfL4i1ub8fVyWXL5IEWXpGXEmNk6F
UTBd/wjWyJHa1SeFrjMgEr4Kw1ZOuLjqfClkL0gcpz0egkwrEI4d8ilYeVIy4xdu
po8IwBSgwtXf5QuZwIVxF6SwB2HwQzsfcw/wxNvNwV2X/bKJ6pmJlmcJ/5sP0gDz
BZAKYSboplUR+Hbv7C9d249wBYk9rqwDjNecuNlu4taWTYcCmvsBUdmhZW5QROgj
TMYsKKANoNshs7bfyivYza+1TbnozULV+3yZbLoTY47fTN2iC7iOUPocwr0zycBO
20fVzYWLn6aFzpOttOcY9vI2a+DySqsqwHA6iI+bNc6MKDvr7oFx23zx5FoX9Ciw
Gl+wN/bKsnucHiDaWlUpSFttv9HP6AXHa55S9fhrrMlYid4qpA2h8pbwlq0pcaI/
btNpWryuPCUr1q8h7Aeoy4auJkeqxxwHBQJmiSzPcwlyAey/puQEfzsqNe6WrNos
1b/wDOO9pr9QN4xMB1hqhXre1ukh3w9ymdXE+06fKDly9g/SazeM6ct98s3Idh4o
/rC9aRHlVPaiX9RVqQm7GXnWUZE0GyaATgz6BVtWko+uGJ7z4IGpqClEAUlPYYmv
1StHFUPnnM64AIZAneJasP+Njrj667zu2YmwaMj4GkZ5q0WCv3/JMcj4TLhr2PLR
SVj+jsnJzB8hiL0bvajVzc41c1NiylXhc153qdwK2Bs781oeh3xR+QLgG6HoqHgq
Z7yujdFrqPaO6XDp4L+HxQYVw7YMD8u5hk5XSq/JQxkUiD9PXTZYz1Y0LphDv02C
IeRIWUEXW7k+ku/iWJY13/1MJKG4Qa8E/hXg+Xf2aT4+DDOb9PcnRKFMsyveb46A
+HmaZIGxEcannxdfGP2ik3Y5Wpsy4NcZMQuS9celRdZNE49G8Qi5/AnmsZgZcmw+
wMIUYZtXodKZr+lhyaz6x7UmczTViCX2XWm2KQGhq39ely6PNq2+aghQE2dk3FzO
l845q+AHazp/rGYg+XHN84ebXb9WPQuSjze7N4pNGc2dnQMtqZcf0NzxCv57Fwt5
tZgCHN5kQK6r+lf882lgynKal41AeVovqEOB5scS7VVNBIfTfhvmlwW87hW70uLI
4J0xGEgpDtgkLwXFj3CAL8Zo4oKasXq8I2iJrwNVlgiJBIprS+WBRp3FLaO9aIOJ
sKvBjCo9mqaemqTryE7WBTmCkA0DyKqWvUpsagqTlVSIsj8icxEmWexaOV0t5gCw
myt6YvmyubQ5vy1w1z+uA+fH9zQ7Lnp56+SgQn5HfJe9tXg+M4uihWYgTj1VpBIW
oaPpcvovsZJNE+9+B6g9l/Gz8e/PDfszRsOhT/ysFTiC9fEywclpQ34BhgVtLaGR
JvSGCFQ9NXawyIHdPKfZ8E5VeflUDhI0sUKR512g9p8FN97fj7yZTzrJJcXsZhVr
Pab/DM3LMcF3/eoAuNmkA5k0dqY1PhsYYdfsWMzMT6YtzR8PsRk+vPcZpJzoqsES
3+afHCqqM+wPu61JbR2iUS4p73IR/akxZF0zQHfGboB4ovDCu3XVwp+u2DmMUN4J
qBWvIz4hmlnlo033wU5g0IZJ72UvNaD5F2D3hMrnqBgvJvtLpOplo63WRceUxpqO
XtZGTHhbbtOG8YNNu/kW4OZVV/iVyRo0UmnHYO7MH9UoYp/zuyMgZM1LVEU+ZSZo
NH7kyVQ32RJgxM7caP/A/a3/HnoeSLaIQwYsS2fInai42dMy9AMfBfXzTeO/QLYw
bUFjSavB83/wpdjVZBmPIW0emg8Rj8CZVqPVevAV0p2nrTUziNSar2Lw54XfYH4+
Xg1OAfD5owmNyI9R1lL1lBJVYCNMrsmHKOyjn1EQeVqgX1vpDnzn0yjdxsklFgy7
NWI4l3LIUQ86HDkUt3BmsbIDQReb0zrUOudtvQhw0+GlSyRRGiJiFdTWO1xwu39L
xozu4yGinoi5UtLWtfhdPdkhW9cZSn2GHICj+KSASNZq4L+5qhv4TNW2CeevLmrJ
Ahn9hhCVkVzUsHSuX7VHzbeYoeU9xK7r89rm3GmTjE2r6eYgQ+8O5sg6nfRP++ka
TJuLmFecLboN8DAeceAKzbB0jlQHrDE9NvnHDHcGDCXEiquG6zKPmzXz29j7ZHQY
KFlsoHnpSBKguWb6l3DcQx98Y9JtGP7mdW7Rm0DxFIGEZnDvdVjn5juosJlhkQMh
HuzmApIlTMfVID7HYXhyefNSkvWIQjH/mYCiNr2kRoyoo43Njnl0GdnJSEUQBTro
NE/OOByA2C6eymix8+JRxkPdD7O8lLg3Fv+Ed7c1fatINktdnTmhNQg1h+ZRZ/bp
LrJKvnvV6lxiCUNmyNQKHosBp/81kzaJ1fDIXyWq8VpT8tr3pY9sb1ljpZJw5UzM
uhdHypFozn5eQRl5ERly49qQ8pvovkqV7v8p+3D/vazwOJ3hOp0GRPw2FEGUG2HS
pQhZVGWKWTRuEUQuJENr/Wh1anm0e9kGSZX1/N1ukEWoDo8lGAKcxOMNP3u4hCto
coDtB13AO32f8jTs/tOmYAFJjSA048DZm1hD5lUwyWWWsQ1SNpEKoPY4vQUtU79n
qn9+IpR+dwPpRtwhueVJUCD/uhZZAH6gv64To4O3402uC685o4sabtZrTd8NY8Y0
pBI/Ze9n8w25uvOhtUXZJ0ZqjqCXbLUwpFHekftvBaIEUIdwuSa/deWyvkbC/HVL
ud4o3EWZgnYm/+Kd9fZ3GCRnYLCBjTN9/iHvnWTndIgTGYMpZeO0t25YJNv/OZOn
leMTlG/JpkgqzWLgKMuGrN1M87yWKtmQlNqcdzVW5qqBbV44xRX67K9seNVLhXEE
xAcKO/S5qZQWC2mGJ1FQ95ujA8VcyCqaweEiPcqUjngknpda/9F7uOGc0qzwZHUc
MLAnApwoRMsEcwt40aMT8pLRPA+SJa47Fzgic6ltaxFUvFWbgGz17/QuJehFbam3
FdBiG97jybtqVf+kEV2A81iRyGcJSVh7dZ8o3DEZtIhVq3V6aFXwaA/8afqxWnN8
Dx290RfKpp4xEC58Z/O6MzFF7HdVlA4Z7cAEQme++fMsF8y2ZA8cxQrVeSsktLJN
jvDYadoKZ2dhTzywj4pBtU2SENM36t39wZ9fFbcmpcvJ7SXIItYMzjxIns1nthx9
AkBwHH58bXMCCAxxkfUnXmobWR9EaRwKKDEVhJbbOhdwoDTpDQMpnxmb3wd/EgQ6
m6egGSPTqYEJeLvlEPTtwSnlJ1oGznqngFlZv5nSC9kAkzybAsxVcMgmX2+5MxAr
LoWh+gbCkUuJwKWBnWXf+EWsdRgU2wCZFdFFkD6HVlHhQE3YQw+rv4rbvYq1Jzax
RcwMVk6IvRVH4oB95mPZgHlse59IrYUYQRwUhgw1NHQ/XNKzE8KysGjvaX55D9Bg
m55eJcGJUXQ23YyWafYJtWISgLCFhMz9JeDTj/pIrn/y/YClevvzWgevkskHOYQa
mvrcuErdC49iVe7xcx3ZvKLc2mCBgV53BPNRWd4MB8+/cxrZ4Pw3ifqm5inq75Rl
IlzL72i8RrqCjfUXiTadFXYHTslNjb8UbuJC1+4yU1iLsGW4R24b9xil3lmrUDN9
g5s3OrJdaZcmLwyZ1dTcNOZu497neNR6+os71Zyo3BoEr3hLtaeYqoh97tlz1H+I
AtNgfX1uHNbIEduN1Ku7J663zDfdU+8yZTn0UI3BLIyLHwNa5quj9kSoCce6cPMt
UWks8rxIY5ykSAGkSpp77HNbo1HJeDdw9pOsQY4UMX4DBDqERy9bkegL8e26pfII
3fR0FT6crfIE/6ooOLYvGc1KBkULYHKKcCUcJXSpjdXEo3QCy1SD9iX+ojPQNLZm
A1yXFcS5GNERzmdUaG03R5F9EEMUOjMiUOmhnfTjl49TX61BJHrjSOfVCKqH6W/h
EFoZHlACGvLwXv8XoF7BSdKFbqDrkMIj5OZmbcwlKQ9gCqAa7TxbSH8/KTBA+m1B
BdBxkTGkp02KNZr01KIEqazGgFFD8xdII+ay2QN3ivTE8nOkU92Y/rpchWHyIUjA
Ch9wQzWquNDLZgU/FlJvXhP3pQho1MkyD6ft7/cDrIKEVItQgZRkgvAaoTyJ6njZ
ZG0otNvYpFErGRVbauMrmxm8/doT3cQkDK0irlu9VP3cL1+pjtL/EV7FQFE+VuKN
C2i9E9yuzPOX/RINQD8vXpZ/thMPyPzoaB/aakpwmWG2b/EtONyeJMUNAiDB0mbj
r3IOnn/INtABCy0An2iD0Q7DaNaX8MkQIEfvohfPvJ7jm/sxEmlacLP6uVOBdup7
bXIVa3l3NICRK592UaG4O1q/HB2NO7vz3X0lezv4o2wzkQvkh59jc/SPt/6mFHa0
vNnG5XA/8QTVIBCL04J7ATXP3ucy75ltp0HbZz4NSVOlo4QTiBSnEj/NOcgzhSHv
4ghceIxjTOuSTQ26MCgVC3D6fFd4IqkdNmE7Glsb1UaB5xJvOpFEecdn8SG18iE7
At4Ewr8C8IDeDe/wZhMRHx/UMwIZY+X5Tpm5vUfFiY4jVCCucqFQCKWoTjdFTHZx
tqzC23XRhKqEJo1b2P4gHOSEWRNhDrXbzs8eVgeUZagECo80VgYRCe21jXnie+hn
/BxjecCjNXCfUq/iTW1h7pPqjsjhR9K6f63U1kuCDZ4GS/fJuqUpgvmd+3Plv4ey
5XHfh6iwTc6XbxCd5RDOOzvdvFBIFTuLNtA59U9fsP+7y4bHy7Y3thby/GmwhgJa
aVLLrYZliGU0c1KwLtUtLlk3XS4nrmtjDlkhbyU5QM267ft6k9X+3cKrWTdtBdTD
fYhq/buGlmjQcdGeWSZNANK6KgVTxe7BpOY+F68E88YO5GLvqUdZBPtj+dM0OTBd
S4/vFz1pCxtOsenJu4D+vwRl8k0G5fIR+11ZWn+q+pbz7GI8x99Ppyw5pigJZNJj
zrRVZ+FIYI5Exa6c1+wrh0jcpjOdrXPZ4Ah6kZdVxVe0mAA6dJ0XNGQ6xVvbthd6
wD9vN2zr3j44v4weqWsUbzuf1gs/JcYyDNdkREzY411MMEZqJnqC9naOHU/kHZQk
+k8g6I/Sdekvkc4nHTQ4TKBjaK0KTUY08M8//Su0VO2og2qwrVHdgSXoC1+gFYuP
16mtoJeVsok1NCGTRYj0jmMMgyFJGOL9z8HUa6ZNxEOBkiSNGAqm/ndoLEbDJMZ6
ZHoRJJASSk045fseTXEEddI61U8MQfaaSp47WCnBlki5CGoBbPThneNyw57hqHZV
YyaawC65ydHsOn/em1vnuQn1IyPZVqUmFz76/M+kRNmZbz/QOXUteC/Mtrn5xzFb
CkrHXaZygC2Afj2HZ61yuT53JrXO8P0ZFqYa4J2DUUaqdeWUBPdZpLlupWF444S9
GP9OnrhdagTwOwRQut01YffrY9u+ooxEV9LAodkLxuC9vBoviVcfUWJHywnRs0hH
OSKSUg7D04qzwkO7LN+AqyxNFiV16v1D8vowbP1T5SixeJ85SOkv6UhDKmkc0ak8
pvGdc0c/zciYvucCX1+AxiHse/DNqaOzRtsTwVKGCq8Zs+BdD33xjwlCvnhtVOLP
ydKGRvIDeCzfqTrRwfy4uHuwLmqjrIWO5o/Nuj3iRUSh+oulIBML+nAaeBNr2ltE
j3HvserPiSxZsul54CcXfum1GS8ibH/HcXjjZ3vebTwmatgOYY4QynWck4cZ5FPI
+ZRa/+nohPo0ZtvqP84zLU4FmJyFOTQK99giMHu1jhqBkFPpTzBE5pnOdvtRHejq
USprEUwoeGz5RSCRv9H6Oqf4RMrPAPraEyVP/F3Gk01X0Ccc5BQpu75KgPWOmnM2
jGiz86if0p5omxtnKRP1tIrSiN6McVBoE5vmQyXJY8WJfHpICrE376Tdw/4Fp4MG
tuCDXqX0fMuPgs1J17D4VdaxPxbidzuadtjvR+qoGh619W1c9UdQWjUMh52PlxsC
LiEr7/B2kx/LCi4vmOu+sK3wP3sjzzkJyHbs7N66wjz4iNhvLeZjRhOcvvlpL4kj
Z25VnRn/smshQnZ62Mag4rU/6rcGW/gO0PKZAF2aNA6azJMxoY9bj5TSaC8/xBHO
YjCiEMixkewz7H36So/sveCqfsUZqVNbVQXM7D0cbD/KxgFH+HV5bCfs/AF5E8HH
hVlF49hY4vnWCRFM3uVGp72rQwUfQRMFXX1e6OgURk1WT2dxGTtu48HTUpopDLCy
A+GGzI4iafP3HvmIXMTFRKKEM0/xenNJl6B5eZ1XrYTuKN5iBmw36zXkpQKyfS3R
egaWqMrMioY/bUw5xqsB1qrKibE+HNmTShxNbGLf+XfbVbxZfEJF9yKhi+ecOWXh
mwO4IVFcTPPOmDBvifMqsjRNLoTYVShHfzIDICs3nvjC7M2gf3OVzlZPXbY5RrH9
N1ygv9myeBAQ/2FSwnFc6hsW+0Q7GkNlLN3uiQKuOOVLkt3tH5zN1kMehaJ514nV
3op2//WVW62nGaAWK4XM63ZO+RuJvTJbssC2bUrV8FPO0Avd19RAPdKyB7/TUjTC
PEGbU/DPHUQf7qm/gMa2Q5zrKpQqHttx27+clU0/hjOayUrbC8gFocF7cMwfE2Ti
fLnnkcZRb/mhAy2MhGInscOWTDBMT4oyGcz8WHS4GX56Jf5vypV8NpkjcEaXV3ND
JyZvlNvtZ5WCT7rCG7GA8bIH1vTGQjpbTvXgdPD0TmudT11NpXBBNxo2o61Isq4P
Lw9ZGsUIWfaZqAwLj/UuUQSocFZ7jMwfzwisAq0yVThfnOKuJuXECV+RwmI2rDXa
FZMO8qIN1ar+N7adt2YHPzEHw3+NsFPdYh9zUdNJDxLkGH4bNg6a3AwLvkJ91GFH
RH+nkluX2CsiIo5eF4TBpB0Vr23DkIULKd7WjH82veNTd5plj3GWoJAccig+I8B6
7fGhYtnp5zdQb5/Ze1bm9sHvCmwdYuDOvsFPGHUIT8OT1EtkM1htp0Hi2DMpLO21
PfPDaiw+XZ4YL8EnZcxqWKO5AALyOz8scsSUiy3Q3zXEfAgqOSJFwUY1kPYeVleQ
vznqCEr+p9kAFq4SbbC0zC2cdS09rIbQ2fONlB18Tm2LS9KPUPYmc7A9BIegDHKb
TTG2YDGAKK+BCkI5qduybvYYZA08ECB4YIXWy6IahvjdO2sFurq6tqmDetDBFD2X
5pe6Ovfeeu5WfUf6es0eUmxufceMjVxCd7eWC4MTR7XsE3CexZ/OhwVEOtnb0yUX
oUdS+8G+JE07zITSMypAS7xbSoeoCNow9uXupSLz8aqsWJrqp/mZLXrLe2Gn6iDn
0+t7GkAykh9czHcunWgaWA1lTxkFsSSp+81P/UpnQ/6CeOBp/53PU3iYh8VYVgpO
1AeVvVAS/WLiaW5431pWit+CT8ZQD7txm3qs0S1+aKPBSSi+PSJND4A18WbtPZrw
ykxsM7AUBc+rVurAB2/seYbVMxSsDK/WhqrBv47WW/qRWEnlz/3UPfZwEDGyD00w
TF9llG56TpH5o63z94MaQLEfFNh4MUdhbaaQJZtWP5VGYBhH+gDdtSbCtLolKAa2
BQ0vDacRvanOsKgFIP+a6N51GlHtrcCTk32MumFH+p57/yy2raCITbwmBPx/AqfA
ZUK1fcc/GNNie/CSOtikV7uSiKxLe4EQ/R0tZQ7h3Nccc0Pbqp8+N/wrc6CXNH2A
f9zXrsVbHShihy6vZOd+FPF2f0wLaHuraVnuDf/znpwOSXfFmLRSmoqdkILK2a8g
pIKKhgm8bpbL3FfGdp5DL1fWD9z3y5+2GL0Fl1BEbt4IZHolL6f6D87nKBxR8IG4
gLSOVkXBS25tVys9VtMenb7wHg8fBIhvfKMQ9iuD4U4h7Q/mvZG5CPvagBP5eYAz
ZaZWPRf85JfBkTus45Iv0aqbr7YjuvGe0jfYoBLyubl7dhGvuIZL+JWUcxtWLodN
bIFWEU0p09wxoV/Sczxfalh/jKrOsR8EcEoyir1wGfnQtYLjXb8XQ1wAN8sX0bb7
SBRyia/rPQU751kN1k6i0rHh4PT0BMeRuCIb0WQ85+MgFgHRGRuTh3UYtF+wWp62
/G461ZJYW2aWWIUXvGNWcYz3D+prGsTlxnQjvJOwTTxDAousyDnkOdLBzhRtgpTA
1diHKdWcbb86OSQc2Q71stoEywG4ZFsr2zcFTMqqFhP5qFCr0d5HNZ4bhHOjfBAO
ScInWN4WIaS0bmMLj88SvrusvTA09bnc/QmCffCeCBc9+vr+teExiNwZPU/E2/Q5
3uiHaPswFmYmzHeyWUke0TulgsRpi8KIuS06sMhkk2EkcR4Sv8eQVAiyZ9lPMadf
aKbB8iX+T0+F6PV2NOVT/EnUCOC4/Yni5H/162uGsqWEnsgyxajo7IjZxBuCM3Q8
wSbcOsDlZmemfN14frOHxcBMu7EItut4pUR3Vb+cBxkQmIiITJtLLRU9zHmD5LWj
vKVea/QY8ozfzhnwumo5jv7TTMsdW3xdym9ocnFDj2y3quuys+oBxyJ+/SwWHVFt
h7CwP5fqMRpdufNWQoXuGEC529nwbdi40M03tZ3KrFW8Dx+uviLhgsUUw9qwZ1oE
xuWJ7a/YhBcGCnEa3ewT1D00l5/Q/O9uxfm7wVv4prK99rZP8clkK40c73qb/71Q
J0rhxaDhJxPqa/HgQoswag0n7qQfMYIJbDWqheVPQCBeXpoL4Ung+6x3Wwe95usa
JYu6/CbuWkoRkCGP/SORtY0LdUN8gj+qbnsdimpF6w1ltzszhm0aW8f15x4Jm9sk
9H4zNDFcShLtA6t+gjoQWF0DNQtwdoxaVV3n/0KBFLg3//lDYsYFNmF4/oxeP8Z4
x3Oc8f6wY6GdciUW6ALlYJczIiRuleO6viveUo171uF2uNRGnFXXjDpdvfHkEUpG
urkTvI02+SxJ74B1K1IbZRUAoNQ14T2DghjlAC/ltTN5RlxOdq43brmGPe4P0fQC
IFR4NUrr+ib8fAVp8TsO9EPhg+6hwu80e06cwD+qdq9FAgd27NeR36eyQNxxbW4i
5Y7BaAXQVDlq3Maj8nqsBWhdCjXBxc5xeRh8kr7xveeN/k5uTlx9adppdaZ97UWy
z23qzsKN3jVw1J5akr/U/P1G4HOCAPu6Q3gTObXFkwURmcKwTlgWHlLtApGrln7a
1RrvpT6+ylUCwdLyzMqS3ufI4efY3QHpYF5EN7yKDRN3hqtEQ5efLsSuNNkPe1jb
sL7wHAUz9vkR/modGU/AbNjXGDqzxSjNHSWDZFqKHTujsXDPlM5dsNFrNCeJuqd+
1dKOlAl1f5fhKp0Pywup4kKKgyoYA2Od5WCaZWC8rTW74kzOSBiL2ZmE8tsIh1i3
ZdwTQirCj2dJlocuu5SA4a1HovG7u09sMIgBSccvBGfoWic06cviivQmh1taG1mH
SETRkXqxZA4q2p8uekryZ07ZDLIOmWrfu183/SXCa8UQviSrpk2eYTT4WyrB+1p2
PtftwP0QR2CAGggfU3LQYGpJ4/BZ85PvYXntrKN9g2/uSzb/WztRRpBEwSep2ii+
QMCmch8SmKLdBbaINJ1SZShg5ugT3RvoCBV0sELKRQnjQ1EFLweTFxkM3N3/FSrN
5p3Gzue66LHY74Gu12ereDrqPrO+VeB/XH9cfUI1G2eJluRCC7kktMhthZ7BpQ8W
SHBwyaN9d/MH3z+QuPuMlxO/lQnjgk+eabQiLrvJFMJi6xqZB2kwunmfCYLfqjL7
CnzE/Pn4I9x6wdM707xXh3Pa+x1ZbTNjor3jKs72tQSu/d4qcipXBQcSCRXafBVe
SkM5Qsr+wQSIyNHWxM+ZswnFtFZLTUksKnTKhSmnLrLP2weSwXXUYiy+bSuqQ3XZ
rIvMwilPZzM9eBn9CBQGWhO2tShZYAdI5eAfOW21xi2OsAdze0femZ/T4ruE+BUJ
vlUpnbZo1UNXblriuKlIU+y6JBUMB7vcDTfkFxD147jGqmoaI2T4cEnF5AVm2jjH
f7rFCjX0NAdo8JmWEkylv4haHIXqO7YH41TvYWwz1dot6VDzgCzsCTakHqm9LS3x
snXerCIjQ03lWbHIcYCTgTnIXCAQkIEzUU28VDdQHNC56JGemwdIUa3RhprgB/iv
oEHT3Fl9yMSJvD2FthurYanUCiIXFniWLmnPU0bd8BXwKKGHTmV/IYcng832kV8B
JbShLzsrsDMoRYLGMBL2WKZjamIdlgjXOABup2TWX6wtswYzyGvgdWTxYi0BQCf7
R+M8ulNvn8up7WZExqHnZELk/9aPYW4/MyAH6yLOTA1Jbv8hbEFbsfS4llWYgdEL
N/+RQcMItCkHddoMgSK3ujz0eC+vFzNLr+a5t/mi7qqQtL+jHTwATwv+zylzY6S3
6QZ4aPKc38/YHEp7PRDnOZX8x58SfhsrAFx6Bq5R6sTHlHXwT/zRdpx9PW/wm/ID
3h653L9RI5/wOkfxhdhRCQ/AJYgbkZ4fBebmAn+ZOas1w4M4KVsrb/kbdLWYWxDC
2/k3wd2td/CETIYEn5OX7RixoOlhc9vWqON+3JiR7DP+yONm39DVDgVNgbk+cf/M
C7h/XAkjl0+hD0dEMTG1Y9CMZO0sbbFaYSmemVIf4opqd+lcNLoYtIKKvy4Ah3Vv
w7Z5nst7bISpZyTZdtGKmOMAe2A1+Vs6FtCEA4X/3RV5JBJ+xSA7cLkjuRbc2XVR
gI/f+VyQTBGugpHOh7ygjARnywWnynC0q0D6SP9YW5lKM7AcKfu7E98RL999XKth
ksyDuWT3TMqaa9mbyTmabAjd/05+yhlBQQlPxmrzG5wDWGUGGnswJ2rTo7R7EP4w
NfO/liVpYWYsae19yiMhS8qvBBGBM8PtRSHsCT1JClJ2uMr0jkuafLceV1m8ct62
WkOythw23i0YxZboZKkRhKQNxAmcRsOOdCuF0KAuiHPtH2rHeIPserxwb59xPIt1
NuvtW+lQChdrVOjjvNziBdFGfFNYGxuJwnvC412G6L9fUqqo4oyupHR60ck1hcn6
ImE371EM/cAeFqiVNL0ip1yd+EHEMdsFPitKSvnCC89QEwOe+GW7PhxFBoi0zqHt
VYB7MjmDOspwsao7MNrfD0aAvmdwzNeYf7e7Z4+OLAv6KL31ujoX/Z6YwZITOyZI
V/TLqwDnn/kvop23a0aG2WfM2PIekIz+UmO62HctACU7/lWgzbMECYTb8XtV1L3M
f8SpSnkjPfwDGUZ7GW3PEjRhdlW5vRfN4y3z/a8oVpjBzy98D89dPCNUjhTVf3Z9
qS9UXBzDk/K7xvALVD00J2sdyEwpOy8zFacC1jPn3b1r9G5IoT8Gq01Dv2fZCHDY
9N82+8dX6rDbzel62wBrNdQPo2brDPTMmcHKy6qTxiMwmOLN9FQuE/x2rr31Eo9d
iGZRW8UZ9glaX76if6lDgPv3Fpru/G9niUXzoDnxCvZ4PUFFur+ZDnZF+q1TmzMs
LBhVnMlQ7c09ZD5QvjhQv3P4oHcR49IEonNhllfDrykIYxhYPgiXs7S0aqyTRnUD
WtCQBkT8zrFjEBPLPUqTEOzU+x7GoHnHsBJMVU2rleqluYCpsoNor7oqBlKVr++r
YCIk9yDZwxkZzYVAxQb126bs7J7jKkNGOjJdByg/vsW7mp6nnuV/Zx5aOL9D9ndp
Gy5GsJygSSShZzvpY7LKfdLZzLnRfonFJC3zquE9RxpOem1nZ8vd8evve67X61Ry
oo+H3/k/k/42Omj65Toh+Wr4FigQWnSKnlvtKLLhEfUfWaBxMqjApp5jnei8r5HA
w3xkRFNENuu7pecds9ucLSdFp/AOV+WrDYk8slkjVIFJKJ+1zmotnXaUHU7mtDJ/
Cl8oRz/3GT7qGNAUZxJ3biuv/3EkC39t7hXfpJGeEW39otwWoJiyKR3+uGXEsWLe
mJMooCWbqIbOd7Oju7UdYMMI6E/T9EJNQBU725LLztXhHKOpBqx1/WAwsHi0Ye4n
k+t3lwuCgMCAOfESS0ihud75e1eb5E8ER2RnykIqRq6Qc8K8+kq4oUcG9PgEk+6E
JDJOVlB6r0LoZq6xzVFCPaUvjfmTsPZHG4FeZfRyzfHGwzkZqFGP90/basmCWM+x
xlbi7P/wxmdy2lB1hTOuWoC4dA3w81MLTDcEUQXtAK+/jbO163cGHhUBZUZbbNGt
S4cGIaYh4VCepX8+MoyPeHuSXfhf6oFcQZ579VwsQ0HXBKD0oTjPeN2WDjfxZwZX
4B6deUD1RbAwnvfQV+3M6aM5LTVTiHhHUNpzeG7qfy4eQ5goabMVl3HCmAbNfCPG
p6Adt6JN6n26kvpcVMuIE2gq/CP5sXB5XfbNCtfO7m92lDHheO0JpI2xtdOp6V2/
mVbUs57q0Fkzte9NtsOiQfqMCEznxICVeoeUEpw6cBJwihz3IN5NzBCWiK24WwTB
8iHAmNEOSqLZxN4rTOV/kS6mo6Dpc4BjAu74wqibaRiFdW/GpR+LpJy7x2BgyVm9
vX60/3OcpWwHUbKJKSnkhfJG+1/Oacu5q5TffmTmvZDRekXm1iP/89fs4Pr8UuS9
5McPOGJaKWr274Q4BTQ4daAgtrIpN6YOT7q7MtvG6oOUWm73a9CQxe9XoDBDlwpY
chGDhTvKtw2FPXXQWSJrJd77rcIdtZexXTiVlvkUecGYjE6c8bH6pQeOmXeQrpsu
Xs7aOs0ic7kJPx4sLIDH7gFq1P+SExc1ObE/0qm4Oix9ZaVDI2AtMp50eBB0iTEs
uBudIUfSkeIZMToP1JAXDzwOUkB7+V6ELAvgjru9TNUyp/7hVwwub7OEPtKeFrCI
mMi8oLxGfqbuD7//6Y+jl9nGt51A/9ZpO08Te8quk4MBOWk4pcIi7qFb5CEtx6B6
wyHcM7LAlEyfSPj4ECf0IuvKBWNcjhLcMtblxHiHPmp+oKwhYFFHih41dtiPn0Xd
2vuragqW/kyKq4Ykr4O7WiAzF+83ILqzD/w5O0J6Xf0IXuOnIiDOTFIwZj0HPV2e
nvAWdr17h6S3cCpY6q7CtvJ0+XVulTpPstIPvsg9OeCvMGTw7/Qtubw8HVd1nrKc
MWaSPp8wK6qmF0VljQyGBOk5DrC3AS1vygylPYPcvZ0wrmSoeCzsEg1CmXIqzBvJ
UhVlOb6Nmw+77iyMXQ8qmCvT4E9hUIJelziAtLo4OCFA8aS8yomRzlgH0rqy0Hk9
9soamHn+8u+zzYeswf7TC78R+3wCTm37CZWaXP0dz48tPcPMhyZRot+AcgFCHUDx
r76MMdQlNkhrgAsnRwEiaFvxKEhz96WUYaIzwWZyxkU28gbTwv/TIYTYhW4r7V41
aCTlojeX7KNKCN+CscPPZOw/uW98sXSXw2dBJL+N0q5i0W7sGkDn9hAmWSQhH3qn
Vxns8myYzfIflp48mqF09owl2lNo4zKwKawfyZ9YLp8/UtoUe+ewvNyCZ3pa/O5U
S3kYpqmOLpWYRC6o2iAtB8GjKSHsAfcdocSfVWffFbSXZuzOXQnE674uqn5CAueh
KzP0reXpkwoIxgrgqcXifmyZem3o4aSxg5N4aj8NcAWEKWnOP46RkmbqPaEMcJnb
yomt3AkAn+4cBHLvAePfm16Az0CZzUTDzVxZW9S5L5PUeRU9kGVM9YAQO5hw7bNA
KpQqDygBxEoOs4v/Jlo3H6YAyGTWrarKe70PCa8orF4ef2kFTA9z+5aeqv7gqfc5
Aek4UjK8mCtRDxW6hx+RryiBxOlmxderR9pybDvCmMC0P/Bl5Wb2cL98Ceq659ur
Zgzx9AhS5r9AfYUECzyEGNeIbSXFQCL4upo1qTreiN7jABE6uHL65NENWaEUI0qP
/K08S59x3UWthngFxOiM9AapNxwVp/IxoRQwWO/UWRU5P49OlnAd/O0shxkFs+ix
fr6j8Ox0zwcbUofow4iUTiDO+bk6OH71WEYZlIwMsuugiSd+OMohlFs3hSBtfVTk
QDNLFeTUb9o+cKkEC41rX4KvsPDwDElClG00Js6KLTSR1F25D3J/lFJduTuk2ZNy
yXvF5x6M3FnaUfvuPDB8h+vH0nZSC8d2pC5PXy+ZqZUZH9BMBRFYxk2HmGgvTUcl
+MA6ZifbvBRv/KJLiQ3z+RZA4fcNHSbC4FEvk1Cp6M6TdUv7TzbSwjqpmuA9Kfch
zJY5P8VHRT8f+hK07pWmxJFGHtTHKnfP0GH71pbuVDoV7L6NfiGFFyostb6hFVA2
9jUHMwfn3Pj66WOAWnvzY/K1YFGkU6dmCjWHyAdotlZIqtY6jkpuTmYFWKW/hYT3
p8At5LRJbgNGst0FEpGk+2msuoHnKiBY2yQUOz8ybMAVTM4wAxrEzA4Y/wgTs7VM
ogCo0nVMBjFrtW4pAuaIRtHv9MxSPo2XrlVRf4gtdVZ0Z9KX319ep8GwxVdAKPM4
CKNRjxiDVXT3EEqvC6u45NAAm3kLR7qTmqnM7lxCxaP9JwPjADX2YB3nAHQBDVgZ
/uWjtL83uYhcn/LdLMy1g+u3r58gV5GK6CJgpyAYd7YO028+iYRAlKeehuyDsQK3
5HgrtJimgzkvXZ1wajISt4zSUR7GqoBfy3EeioatcSVva7d8cDeuWhp37qzeEsxu
BwlR7zy3ofaESkuvJcYSE9tbF+RV4Szrw3WvxTLCUH1IuhDMkUq7TjVBMcr1/fyf
Oa8ap2uJrUentqlceZ7eOJv9mD5sSdxiC2QxoSi8W/R4Gx2xA7cFZGgYZrmleovD
1R7QD3TO8eC9hcCTZ3OuGTmrRMSTsLPjpbCT26RydpYDCAxW8H/H82T3TOSpQ2vy
3YrCX5Zxck6qnGOcspiKnRV4LrqbmDXEy4j6A5QNpNnIwj2J0KfncF4+hWcy1vZv
M+UXJkuiUvrfgZVim2oy62O5+55PYth9eWSlRYXowY4m5a1iYWmWeLFQF+M/3QOC
W+HwY6MzZerddxAmeS/qyZHWkbsoVfUVsX94P9L9umaXuFB6YECNHhXaBXc4Jz6M
r9kSQ9F2Hz3MFct5oe7rDReYes0XoNKJ/K4rHevOcaSqZQPd7XlXOQa1CBrkLFTc
pcvw6zoG8bdtPDHsRAnRSW6glJPQbkXyBtzxnQ7hSZWcz+r4BRKNCTAvR9Fu4iq0
M/sVXfHS2UC0OtCa1pk7ADYl6kDtLOC+QtNdiROGnKQpjFmKQ4NQ4uRRJcFTg02x
Ri1C+5iWypAPbFTOJQsTsj1MgeRBQAh0SkgDj3OHJxnmb5Tzf/hOYwdHNO04Dunw
F4sV8uSk2mGtNon5G0fZ+Et6YlE2hOitPptv6d0T9B3t8QLoMWCvI9FpFUkwloHC
Sr7NOmcjLaQcYF8jLSNU1oRD+l0nvVWVOcqvp8NFzadhBXWAmTp5dGZUKpW/0H6L
45/1FWdQiXqZd1G2tVotMvaiM3PfY+C/Eprikql3o849mHvVTV55XVH9qAOEzI1z
BP6gDD1ICsIRP/9rVzlERHExx3lCX5JM0eCX9GHiASKZs8Y85ap+eAVbU1EBoj8R
Ia9ICgg9fB4YpERu6RpST8cXo0W3+7xuuLySrSewjov69FKsmgcNttolr0bgb1ao
OJf1hD/DtWttJosEEcD0yV549tmGBetQMj1tVqvyhO7G6+Cl+TtQlbc3LHAbusu2
G9nxEGjrPQo7Dx1qQULkME65Dd2Sjz8kGqj6f/x19ujmPD2BnfI7lZNxqL/puZE7
ix8ZbNfsuW2iulzf69T3Vt40dpL3bzGFrFwhzFHU7A12WpENBKDD1Qo6pspH7ZA1
6m3dtOWA5gKMPCC5zh059A7/gZjVBe/mfuSxgeqvkn/KJyh5uHICStFrn98Ocxim
qa3JnJRF0yATfhpxAxMdBvUH259SogobUz+qYV6ApALw9Q9UnBg4S9TS+2S9n3H0
qFFEKHDZItTBaWGHhR9uLbtXHcOoVoS2xP3YAyAW07x87iWingkLWOCT1zc4oxpg
83Lgmx7/eN7jM6X3C8g6VLM32ttT9a0oC9s+6pAEmPXYJMw/00VsL7TWwhtc6wQR
una3JSCNbteWGzp4YTK7AeeuT/2HFyNlcB54hOiAns07Z86jy4I/VEZbHfX/iL6a
rlxVDwMU+545WeFpEYugqEvan6t3Dw+eaOikEACgDeq+H44sAycb5/RDjh9qwIt9
QAElm/QQ3ZQFg9W1oZ8t1RmJ2kIu8+vbCKkY5JcXPX8eQE1IwFipl6GF6osGetLE
ea7mg/6VoIbD0bbvUna6RYhH/oJYwY2rVgVPPGMwJsAOQ1XA3Dn0VM3+NGKDpm8P
8j0Ny/mOCC5sdONHi06XdYVDjjQPegCNLEgTuvIzwdM6yTwF/7m3flwQRovJdqHL
Bx/kh1XU7Rf/mTGHxV8S7OsgDP3d9G1Y5PMP1tibxanA3nV1FhLwo6vkDITnjDF0
k7IQArB0baOJu+1svvCqCr3Oz7YincoQoEpY7laaTdLzl4GcqpylZmOackB5zJLM
Sn96do5roHclhEXRW8ktBWiBmILlifcQypjC+Pms1bpE+nrvWUErmj8huvfPhyh0
AUI1X8mlnHJNzLOQZ643cjCkTQTku+3Riz3CClAqfpxXISoZ41itqb+L264XS5/H
5XRPOIOF8KwfMtCSdqLCA8eyLtsrYgiS6UjR2ivqB9ApwrT90YuLpz8+H2yWiGB0
SlQDtig6hF94CEZqDCH2lf9WSKe/qn97irmkZapzCTUwhFDVGgIcRCo66q8Id18t
n1S7TWZvjX6tCdib7IXAwuZWB6vHjM6bP/vBU0ZOH063X4OO+H7TkCYIo8oMT6Hh
kIhRCKxf5RMGSS4Ce8J7Y+kP/nWk13ks+idra0laiu3f3f1UZzGGC4XIYDRY6uYU
yvSdfO3Pfgp4WBF8gXa5OWx5fTMUWFlRPBufkR36zeYt2DlgsLrTrQxG3eBW9oOO
qQfxLD5jdZi2cqXJDAPazKT3oLKUO+DXh38gGVeqZBeuJdApuylsjxwG+sG+5wN1
C1/i4qwT4Y+4OXmJhQg7QdtKf2feQk7zAqLAOWq8wimHrjWsf/mc4barlitBNkjF
hxKF6S+A6kvo2cO4zUEMowEFx4NBE7gqa9/fDy9f1EMelX3X/k+2/dtzksB0DbXr
+BGOXaIzqdfmwSWq39AXLs1zlAwKV+k9N976+niHHixDK0waC/3FdLFwgUumDxL6
2Rwmh08UcmqPH6V4q3GxEYyoUub4cgM5ZwUFVsJTSEX3yw2cwl1ZFznTpRPYybvV
Bcm/iJTyjLMX6cf+b1vhQsAjhDddbH938mclUyzP7d9O8i8jxj46PBBZa+D2xDUL
Sx5SCRjonWsqHfdPApk3w2Wo7u75l4SN2cZHLiK3OfU+QQFxwLkjLi4dH8/cRlEp
jnbpxPkpFETrzHrQSal+p5MwHo88QloNItRaLsv3wniW4ZON08ZYNrenRoz9f5Eq
xcCkv2t79dB1fiDVmYr3ILMeF5/FEajFIlNCWbz9ejreHRJilf8/a/kp2L9YdBlU
aoVpyJYQe8iY7Qo+xlHO5vjMF+YeAhUqaTtWbGwEDjQNejaIuPu/2VPQEFxtxXip
2tG15r5E8cYAk3u7MhkcYHlFfufjFHkQETX/Kr4nUNe2GUYQBYLbf8M5IwDlwIoV
w0K2L8BWaLYfvSgEbA0+lq1LP+bpb/achmEzj+koChYADctFmBLR3qLYPjgRO9wZ
l/gbRKRAkmOFIjqoXJsm+AXsh/sPIe4/1cLX3DX2qaNsRUSQTyB5OlUXllzyTb6H
H9cSeNe+TR3+nJ31ydh+7P4gtMOMbJNljHQTDFTa2XD1e0pyJ7INMTdM6eg/HKPA
0hHQOhHP0rjIuwhbexz2FISbpMO0S+Xl1Qd2YrOw/I8veVUU2/nOr5RRkiXX+/G4
/xbcLx95lcpPt/wpvXzSBhKXqSMrDL1lBl7tG4Zzk+NmLHEnYQbb0vD2RRyYQXCo
WueqcaN2pzIwU9LbvVyVKqEm4+ZWkbGR43agVwvHmedLgaj3niEIdjlKG5Fxii1N
9iMe7odePlQvmK+hMxYrhKJul9K+SrcLALUFlImuTyzDnfXKiyD5FGUHEIUP0uwO
TlquBVbN4sUw9OBKlwn1Kf4rawpQOwM2KUbLJnvSh5hjY1tdylC5cNTsqH6+wotn
tkOa0m3gGJbqphDInLqKVgNalpVNnb+8IYolPWxaKdGOjOH8pdRMD/WIoqPD7xQi
wkkYoVhHyb7i/cIGm7J5/Mtv8zr1XSxczHHUp6J26PIBxS3xFy7PgSuAvM+1/VhR
5NpS+BX7Xu0oP+RSLRGbuoUbM2ZhjMoAXhwiAVHA8euK626WYBJZVBOmCfCfL+my
IPa3Ir6YPO2+SxmpjHsXTRE3EhArs2uXxrzV+FQstFNFwPibYatxfI73G2Rv0vYO
P5X6GdLmRk1fHrlklX0MWWvfg97tLHtubQYi1pg5fEq9iAqoDpTMELGqpobmCJUF
oQZR7Fbl7Nm4yQnbPUTCzlXge2cgbsr0E1xdHFtKk16cTDz5yVsDneMLnziQWiE5
zJWs1lRxt9e1iJWMfoweWq87xDmUStClZmACy1hfE9jckbV7Zo0FdABn6OC56zxr
++5DZI6wp4Yzsuqa6rQuLSOoXYNNSSoh3jJBDOl55l7jc1ZAzLkaNRXEOvzKIVA6
fI1f9KKdA9u/wiBQZl+N1kzzKNndr6IkoXPxgtUmzpQsWcITzWLr1DTbe0kXzo5H
S2WRfSppNCfqtCNIYe+8YupGsFxeIGplwgoS/WtQ00P4UT5S6fOgqqCaU8wTHd8E
t7aSI07Xn9LVmgd1CXm4FHz6424T7JNUEFE/zbV5mt0vLEJhWsy+CkcObVLxSzJV
4G0amHdHislqmhb/Nu/9ULronF+tReprHOU1+kkpsgiTr0625SDAz9XjcVkbKEjw
7igFNvpkcrdWQBBn9jk7w6XUY5ChjywlrrTSdi4dJu6YibUzyu7YAo+b20qvWUzw
wJdC9saMWc0PR9f7/nVXeIDvCDI4K02yL3TG0LgA0yn/Mt96dBd83tbyl14OgVUv
Y5XTHymfvRaGelQMIf4uG//W/fb4+uhRgReI9rWN5PqRbLFp/MtlCAQNFBgv/TQ7
+YbJS9SreXX09aYkLZmBnC1Bu+JoRbu8QvyKEF+vCjXKToXsLeGPHyjI3vTnCj4X
efgRsjvQewOb5REzADTi28LHX7tVmFeNJANdxK/y5L5qYl5X6XZ7mgTU0iKamJUC
dPtpQ7P5GrMSoPuq+LgmKW+DOI/u+KtGpgn2p4q4oBNh1tk+QFncM6u+FFNbC9um
PaPBXQI2B7uXTjdIW1nzOLOG8lkhOb5/hNDjVCYBNEY6w1unTm0ySMVZclEGjvWb
s0PZh91ytl3wGAlEqzoBGyPoHqw4ScVFf1yPlaLeD7CzwEqeD8xKpm7jUTUhw7Q/
z8LQBB7eDvJ96KqJlwgkCdmui5sob5ph7lD/5jRIRm/YOCyrKFbLh++gnV7NOuWI
NfGTMpvmHZfIUGxHwA85eQ1MrAz2n4b+7OWYYOvWyflVgIpHwLflpNwl99e+X9Oq
LWS6qLI89F+An3rvZNbNZhv4mSvtZWlV3bOtKnPmGZh6TKq4Z8WXS4qWQfHoAP9j
kfJSeY0anLgry2bYJ5sNt7NQ8uq+siVSleJkUkBCCMMok/WzbGnG8bszHmPogWDI
GCJY4WGbHGPb4HA+EBXXwh8McPixSfLoc+ZdldO18yVDyoa/yvQHfZiFc9vXYhCV
xix6Q7C9Ww7y4pTbDclC3aOtJ5QvqYsWPrcIpkvQWT9vEgbfx3b1xGTSDXgQwF9L
qLmeE9mTPnsIRu13Wbur2CuR7i1hdNrdBaK5zwwQnIXYwliUnM1wCgHnwNUTstaM
9YS4uejo4QeJpYwTuTQNodvmfFB3kfJ1WbvVHANRB+9PW0+JDzkYHbzGpxCaKT5W
gI5KJVz2j1rpkwO2s84yirhTUT63EM7K8bpFDeocrVVmctDa/WDhqB6lOdPikQuJ
z9LDQbSTNmGlZlYitmI8DNtUA0+27oxPG0Jv78d7ahpVy3XXjhIWol3pMqwdBVP3
E6T8jw5KSdLfTcOk/ow/NpQ64rHz/I+4p5WcgRgGMG58Emln2wuWT3HIOIj/0mYR
5VHqr4GLBzuVC4e1RMrqO5/pG1cguPszDaL8wB3OV0pbBnQxX8mu5xi2e/f/M2VE
kRodtfjhimefx8o3EUZjnUpLUefcWwjg4oyYZhndBpUrLAZUmHLXuCFPGyurnss8
tHqmRBB2kGedId2eTNCSaIUisjouhUIyPtgVjCjrkZyU9p4lOjwB+7PiNyN3g1Rj
A/TtkKdUS8ai6f0E2Zeo4d8CM1iBZPidFWIHQoQZaisDJmn/Yrxbw55otzKV2OdD
D0FfauGlzzFhSCF0KmKIViUOcwCZLKnrQ/xZXUPwi7HS71p5jfpt9Q9UfGfGJxjp
yC9e3bgl3/1jhvJSmRavF+yAhlzDo1nIVoOhfqkTVH2FYMiMrYUuUeQzWenHfl1C
bzRSE0PrDQDMJuI8e3WMuyZVpD3ylNk/0vuB7wlsjQZWS9rsRZFc/aAwNjmVQrfT
Xy6KZsJTsWkDUQ780084YuACTlVu7wmDz+5e5hAzPlpAASgLqPpxKalsp1unm8ba
KIO3IvcTRe50gXQ+2dlQixEuNac5uNxtRunH8KexKTAYAhIhIoNUq0ItGAzEj4aN
nsXcAdOh5POz0DSFMz9WErQoVwzbdCma5Vm/xE5rTiMpo4Lo82LjyKJdqTDKVuOk
vYHlUJgwlXUG08E0jDXZMiJI2/a9Hjv4sElSLPHdjrBiAg4NnBZCG1ZKwQzqp+OJ
JiRs9KVSBiZ5BHnqJ5LgSv81ENxemXVOMhuLbp8g2jjO1M6StA3/+fjp0lLxNFue
g8/fpZgmcVqyvjmQj01DxF4CPchJx1aipooaBIDnMKYs8mWL0gMc0khCNwRfmGAn
AhOFz8BbDUtu6PTJEG4f9NduNLn6qWQayxELjPvPmgjJZ8BlYs6+5xZILKU6slZN
KOd98rBxaJIB31r/6QdZg6mG4N+mszw1yIUcf1iqC2gFniCZay/UxrQ8ZqVKroKo
RNUX5kzzXiWuzq7PzYUws/pZSe8HUaAMynVdW50TuYxYDGLOvxNm8oxqcYZPNJiE
GD2YimLR9tVhaIdHmf0ptW4smYBwwbMFqiB+QrD+H5xGQSV7BbqvKTHF3ZSdfgjA
9do1NxwRYa1lndLRNpPH7tN2xVNeWqEXcm81Zuvn50KnO+UEcwLqfqeINyxJUh/9
yTPIQVxCtikRnGi0IbYHKBon9yyXsEhWLFYmiwyqP8yo1hpXFz9QduLprS58iOkX
zd5fmkqUYXj9aTou/p+s+iyMjGfEbNhqjeXCcWgBXu9j41+MbCXT4hD2aMZsNzaT
+5R7leRvytKz2aVSItQRMteF+AJrceOhtr4KWjNoNTMRFPk/9xDKy7kVVvlDx9JO
2tvOk7lQjxxudcifMj30YIHMie8ef3TuCEsF98LtfClIkKDILr6WIZIHNZIzYQmg
kxtr+brkkOui/SubBmXzS/qDdD0eoZhuUrYcsoZl5c0CFGZ8grzPdCnKeFgv7d7s
QdbCLownTabpz/x5xqSnoI6PP9ZeJHNywJaoqxXrzLfifSH7u2sDeCNsD4Q0qWjJ
tQlBFiZXeh4yd+Afs2EEJ2hUgwrl4rYXhNlTL2VME+oGik+JyXS2Z/yx4EaBCcal
aVT3J5nnA6ffKbuaZBguaimeGh16WUEf5/rTvqgbpSmf2aoaUZlEpEuUKtob8FqD
OIbQA3vX6Rp0PP5uxXupUCUCMSQno948McwLkOt06lZqrbkij1RWwpgmKE0+HN6s
/lIffsULOjXttu1xeEWaEP2Whu9cMKd4nXWeexNVlgc89HnreHlT+wPEsXZQbndG
rBV6eE9oT0s/i/hO7H1GSFzPbq9Dxt/4HbJZB+owb9lhQ4KIFD4mjtMjkhXLu3CO
Z5UB5v/wV/wzl+2RDK7on4Jndgwupad0pYRG4nMl54cpZhGm+i6V1DuwInS+XIo9
HokF8PRb9KW+TaWF813acvM7w7mIQ3Wd3l2Zxx1qCGmRNvUR/307LUG6HGWwoekq
cUwUMKxEQ+IfCc9tS1V98RVjURiEMUqlcb7PV6vhKEsArDK1wA1IsPNN/20+UxX3
739vJjScTLakWUdcTXTAW59316DV/BcQ+CItt3eYNjH8c1LesB/66qZuLHoV9KzS
VPvQWFhaguaQo5h7iidFjvAV9JsBFYItEKFs3pDegcR8v29KumDMDpWTkHjOPx7B
wNb3i58zDXg71sedSSfzPFAqJgLNfbedm22g/r3NkQYV6h12NMoRjWGQkO8X4BaB
uKxeF/SScqGRPD9Gml9NKmMvBkMY8EEZAoMFbXUamF11ECQ0RyVe2+aXJYIj28Ei
HLbNFuvRXALc8opFruB1BCGFyfgmQVtW0oGZUKZpZ0WAEYD0VEpZstaM23BjJSmp
exQw2K7k6CYY8IktUU2dALHIi7exYLI+xTJEvvJpTziMXZmGgGuCBI8FtzLMMoqA
BNEbPDsemgIhk4vI1k5VQDSdlicnR9zOwCgQ8bs1FvRtLy/pGnXEM2l2ElcErVeJ
c84MMyX5jt09n1m3BlGsHWKgC9jfk7adp+crBW5IwpZEhGX/FOhQLrXmyg4Lg24n
L0+XWtMjCWM21/KOb8NseX59wSnuuntYJ0u0iS3FJybhDomgXm/+kC/VViDgdNuR
U6D7cx1ItTGGpbi0X+eS+Wx64YCx0TP+gIrAgk4/+fWF3vg9kn8l6rmp9t1w0gal
1/wbo8KTL24Q20miQqlR3N0N86KOeAi8/3z/SfWgoZ7VpCfDP0r22OQ18qU0pQ5c
lrwvzi/PZyY2CR28t6v2bD1Ww3/pYRGB+tirhbFOCOxM3LwgXp5zvbeDZ8M+l5Rs
GhVjn9GAt3GEZ+sYYmCDxZVbmvbN0LGyxZ1up8tvAz6wa1fCtksJAjMpOk8dXcsK
GA23n5K8bk8iVlfAFkVjhAHeomhvTNAbQj+3DIU2xSvZ5l16zU8pJNwm8x23a9Ut
EUr2dEXclsiibXfkobcHSnS+UIbSKkfDOXF79GNm+LIWH8Yd93/kXCqlcDwnjJao
9RAg2iESwWYBpO36Sf75/Ru7pyg3kYnERdjlKSm2NmUv34NXo1gMQpWBJbTSJatz
Npq4l0+BWNzZIzAG1pybvpPglyuX6fDN9wE32O2vLh9ldD58RSXK3wkQ1ZkmvDVR
sHgZ19I7rW+jJqN1H5841io4uNaC5+7iJ4Clw14sdf5nrFMknJ7IO7x6FtreHkwn
v5bbInaNBXTQ668rTHbxrNAh96Ht8pXQHX2gcjGxcIcSrDTt+FLWFB/BVmPPdtM8
Gf+YgcBbFFG+hOEtoTZfKWnUXsgxp7fQAf9E1JH7H6J9txxHHLkj0QTQIRYFztUv
Fl2zno0Y8qCEVPAGlV1SCVULvlzyOfjbIYlOeOSIPw6G+dj4R8bJbHMUBEit7iZk
lpk1eHXdygoZmqea1LSysvLaHK+SmKHzY1Vhx4GW7nG9hevwnPqKhOsrYegFdF1/
1lqlro6umZMlqddaJ+8jWaZ/ZbYXYjeLLLe0pGR0pkXC7Za5XQLagguS+RQDAL27
nLo/08qe+yeO7dOelthWOsvJ8vShwSfM9ZeUo3k4lXEcesu+GIfxxmE0F739Gojl
3H952GvOEE6N5nUrZMSBPjDbclb0QkP5hMHjWSFcvcpC+Kl9+rpudDkMLjcSiXC0
cPo+UG72FAAqHSWw9syFVXC6rUWZYMWvBvJ3Z0POtAJEAy+HvWmZoSDHBt2DKIQc
EH8Lb99b6z1hkbP83Lh0B3UNuxvG2vThblBt2zscLvtNVAwh2fUUl8JqOCfQDzcv
U/OyHObhh1fC37m6AdLlVxiYUh2MPG6QNIy2HwIQHMqtdURG4LnqKF0Xab1roSCj
uvQWU6OYuTuhIUo/p0qg/i1vOjYwKKKCVxc9+idbXCtjoUf2G0b4Ivi3QCRbaCh8
qUlknshVjuTWLmgmaqDmj3TL+tNabx9AAIjF+LRWCWJU3t3P6ehs3VK6YRTSBZ/w
Up9mONU6rFVYUoxsHRHIYhjGSypjZ02HVoZdJlo8kxxYP901dJWGHXvXqKiDCAUk
o8nkaXwHKD3EXEJKqza+Jh3NIbdsdoae2D2QKGVQFPj6ZM6598euGHbwxeu3e6Jp
M81I7S+Za/poywN9bN6N7kwFF59c8aYp5KeRrWr8uo9M7VwizPID28UsNVNkYXVe
slLQEDo0jrawAVrOLVRh1x5K5WFqnUs/MUGrm+hpilO3GWRkacAlkgFacqQrI4li
x0fUVMa0tfd3bzoNxbIHpxcHocLIrkb/ST2xaKdVt33J1d1dhc3qtdxCYmHf/bYG
8ywsBsdcxpzZ92N8O7ZQIWUZhVpXGBnVRwAaSEWYvfb52e76SAqFFvd+CTKrvTqD
WOgykhnOHYxULyWQPRE+jSOSQh9Pja7PZPW8JRvgNkodNgIMv8Nu1DxeN57gzzAx
S2L/FXh73Zklc2x4Dhyc3DuKhhAjCl7FkCfcNn3gasPvRDO0YE8zF18PZ5wy0xaT
c6pUIQJTXT8z9d94PPbC5GGNvH1TOaGR1SaunvDPrKdUnDgBxG0m1tobsfQmjI+r
zuR7hmGZVaSe91TyDDcTgFaniiLhxuDUcQ7poti04ExgSRGY2K7Kkhsea1HHFvfZ
TGSRzQSgwOyR/1cgeCt4zT/mjc7TApAet0KIss8gyTR/s80JUIiD9rTUvRxSw4g3
a1bSZbVdtWBgad/To29R8QP5VzPFypRfElgchv7wrRWn4Mhz36vCMh7GI/3NrgDw
4KTtK2yXOuWriaHlvEkDEG43Ri9r9EU6dfgMAV9vDONZN5lgGQMuoWF5264j61lK
VJqYa3hne+fb+tjVG0aM6ldCfq48p9RuLIoU6jc2Lny8HQtKH4KtJ2h1eEeU0TMI
KhHnW4CQeU9iQSIjY0CZGqUt0u39B/J84MjsPndKkauZ/jTA0gukdGVdjFt4QBgj
+f6v7zuJLnTKTGeM6d9vEPhXVl9tWV9/QULb7lsJXVTA/XsyqtUaHSDjlRMKnPr8
YtcUvtOnmzvsqlkm655oOjyrxU8Jw/n7LdkbUazpi5aOkNF2ygYIw22qxq+kPQsT
44ABvmPv1C2qWEsCc+lA+QMxR/I5/VuCgalVx/YO5SajNxy7Y6yOZs9L7HyZw6tN
dlzwfr9atL86cAE7+ThpXnHaswl7LsEUseyYL3NiPXSvtrnOlZSFDPbAR5XtRZFD
H+L6I4HZxWDGREPS/MbV3u27sxpjIC1MW/EyGuwvuygb2lsbmzjPJgIbPmxRlqW4
wtnuYVFp5bZWGvC9dG6c+Rk8+hxVjoZk9HO7cnhdO11Q8X7++H+/eP/KPGW2p0mC
ev4CVZleMoOkDtq0Pq5EGp9k/7KWgeA44+xWM3LrT1/cBOehc00/kgWj+2B0lHAq
YtiA+jo7BveLthFMVgHGbFfqcvfIoE42459HkY95pvbmcUzStDtcS06PKuFraUZ5
kWG477CZt+d6IvOVWEwwFAXfKsRk4HfGBgQB7fpEkxpqPIDa0lVfT6jRNybc8XqB
ei3Busmk1eQj9FpCABpc1clBeXBaCuxuKSLPHEZNmDvxnpaOhv+u3DF2AQLxwP7x
8Ko+KQBb/FqDMBikf2U2iB/w07aY6kyZ7KdGGZqeUm4Tb4NcEWwEhoFGKbIvgoNj
fXpo/AuJXmquyKnC6B6SsV2mcNPlf7gLZj2Aytpyy6vm7zVirPa4e+nEO4xOtSX8
PqXj5cGFAiVKRhjIdoD2ZoR9yVe8opjqZYnynSjmyA50sbehL4uSqOIkkbzk4xfh
KOWctisLmOPwudQt+Fq7N7OBqREuVhBq6KrWH3hpckHHFzAtmsM0B7I/RJ3jO/ms
BbsF5PAbF8E2xa6EXp0KikW83fJdifbc7iTzWky/nZW1svwnZJY8vyYCjERZQn0i
RxOaYSkcyrjKhYRlpc59F35re04FLX/0+t7+O1u5D7cmKtHa9ioEveH9e0Xqjwrs
Cm1E34QvrtPG+NmKvvprGrbEEOdCHOGHJX8m+6ULIrEnHR4TA4w5+gpRJr7lUh3D
ds9HBo7gRby3GOKySeNcdg51KGEMRQG+MFQLkWwYA+vS9NIgjJ8nEYdA01x6LNh1
yoJzl5iTIRKjxsLY/iq3J093oV4rszWbMsI6QCS1EEPYnHE13wthW+3vg01W2BFF
pSFCTSSKPgG41r/HRvDfYnXdSN8PqpTGjvuK8pSc8V/7XV3WFok7Qf5SjiVtMTfd
LoT2WxBZNLBdMXGR34Dw9CaeTx5E105cUTKzDWOa3MgSJMalhwhJak/efLQ5o8Cz
usHrZI5hVuHSX+tlicvbrPjukW9MkioJmekRD3stbRoGm6A8Iwas8k0edjwDn1y9
FQHMpB3GHBP8heiJHYTGaHFvT/+O/Hx4C9swtt0yVBeh9BAbdmvhJMeKEhnQr6Uf
cAeGL8MCrZpimXaMWQq94BgjAXtl+Xkegl+yMVmAM2zhNEd8QcQ7kTgKd37OB2L8
p3FMd9cyB8PJ54A0VnVSiZFuru7VhBlfyUUZEjytB9Naj3MhpoGZ5BR6lUdMFVgA
lYE8yqBvW5UMS3CE9Wo1cWphojSwu+CKfMVuNelgdy3TcWjglWL/5oxklhHKfXXm
kozozl20ZbBEwU5SLc0uPNgcDzX71QxIIsh5klg9796vcCd3Gq27OUahYkEfy4k+
yv1b4JB4QT4+hXGiDCGwXv0rAblvF5V8dbQnzmkw31fSuWPu2qdPsrm6iXME3PXS
hesCqk5tnqBFK/h3tPQLd5/LT0J1nYtqXrGG1yJd5/SBJJKlvdqwRykHxKRNRSSQ
R+ATNFkcSN2hAcVjCP6ughQu1nTMheC+LH5rv3vK3O0r2D9/GMRjUoMC5MxZO8Ur
ynl4lWWm6dnm39h0T1JemwlhYT+4Rm9yM+plUFMcW5pglAMQO6ebzOsfISZcsQjB
w+17uQpE++yemffSB+zQ6/DEAYzLZs+TzJTA2dtmMNahSLMxZOptsJoas24+/RjZ
J56mgO46rHT8c0pqtRpCVD2zojJkzBkQPgb9lQ1CmAuaUV2sKM2Ta7ZgXxh37F9f
Bo5gUGZymxV5BRTTL65cAiD/aTxDRwZaQrqEVX3+NBZOB4uVU3SumLdIWxsi/Ny1
BHWPKqV897KlpjJvYaX5gxHZomvLgT0tgzWdggvGkTpw8Nmp7O9KGPO8jNMvIkXC
uLY2EkFaZDg84l8hw8jKbVzopUR8vFD5iY91jE1Nb/pFXvV7pdwEi6XapPYXCZH7
6l6RUiwwwzVi80E0Pc4D140TPRenYkAzbuMpMzqn15LrS48dRESHv0qv5p9A9A/b
OwaNL0Y+JssVIfJNq2t/ej9x0Bl45e6tenGYzDwt9LE+sMdf2nCMQHeQMv+vdmv9
dLZ4kCpEaNzauaRgnPJ4sJAjHhRFDUUYsZJ/HAoTmNONmYtCT3BqjpFPWwNEaTsb
vB6ib1TW52eJgXtQHST6BUVVDAbTdrfp+ed59reaJHMNLXd3hbcpd/B28LnvMLfB
7kh63SUdDEGvdX6MCM1EqHIWsttgCwBoy0hDZZ2PL6gTR0haFXXpdpLNItcYGUFD
BKaOFemPPeHmoaBYd7PoGqS3QuKJqvKgz3P73nIAmcE6XO5qcvLYneyqgwCqK7vh
y8jgC5AloUeQzB1soyAQ/+uz9hTQqhKXkKbMaTEak49nJUpvpAM5OWoRJG7j+eWu
a0UlD++FmrUz4OxAPQsbj11CFLTRNKzqXNixg/pGiwJKwA3NOG7AnR5Q+CAcrtwz
KYvyy2O//eyspT2JmZ8o5dIzYcfGcpGG9Gnfiw4N+88eIdn4KUohO4dQ65wjz0OM
CyOnCmn4okVqwEMRdmp1NDll9OrYNd8oIQSAxtAH6LIFv9MAAHT6bGcpMg4w7zGv
9Y3j1MC+NkZcMkzeWNuWj7wvQPIBrOw7TDyKivp1kPWfdo/fVqozzDBbw4stY1gY
zsLG+wUBdCAJwzXmr1tF8Ry0SBdOBsq60IsoJR83WnyMnYZ28uBL6Iw5GoDl8OtG
Uz01vyalA01yNfJPul6cgQgYBmWsKZyKf2w+zgq/4BqCSYKn3juzXNZso/iyRE11
qik5rFCcUEig6VAxt8NF+GPG90ALbS4/T6CcSYaVPZpyFqIXvkaHUDjafY8gqSRe
9AD1pfaDE6WMgBHgqn5Tke45N7a2+7XOVv367hlrl2zgt+V7Bg6OtARqrT7Gv9c0
Xk/mR6nBPV7M43fpKs1CCYnO4wkofhv1x+4p6ompnX8JjjKxSH4F7+mIE84IpCQs
jXp9Ri3gnUyLyNq4o++OfnLvIWKaqDURkMD++Jh162AlR1a3dVQbZaxUAx+0w5M2
sN4lk03/kS2fbmZ5s2Q/F8QmRapFJTqZ4O/cYqvpZ+b9AG9tWu485CHtXQ45ITbs
Fvct7phfG4zZxh/GGi7no7F+8cCrTVRDv+9YiajB7ISMiKJSwZlhs5Bb+3Wnttup
fPBBtuI3R7ySTM5nqDy4umZ3GQy66fG/pprJQUD8b2Xj03gUTn1IXVCROp6/Hf1q
9xDM3q+/p/ai86EGJ+jhq0+j6Dvi5VZqay9EE09uduwEC4oTyocJAbSFy5narEiU
Du5onxykpL4s0Y63JRmM+XzNTwzO7DSolOrFVnAczTXF6Xxxdt01/ObgSUmenjhg
jcDCO+D3Yx7WXSQ105TpxhRLaM2M3xlB8HeX8YzFkH65Lq4ErXEdA3G4fOxHzWkf
4lCwVcdG3PSmPTcuo3dTnlBPjRuDRAOBN7maswhKCRyyYgGzffHcfRh4cn+2qovc
RPJKhZPJhmEKCT8/6x5WbVLLkyCrAC0jmH82Cqe3dZZp9pnSphacyJqqoitwywYc
IxG76CY2ymsfxqe3PY0Z4mZa/k/xl3DL5kR0jv7VTzbMLfxmBrdYo0kWd2fzwsmT
0kSMYPTevJAsHgqhI7Pjv9S5dNufa47zX3Uc66sFjDs4QY0A/0MDuj+srYRI/U57
zjUkLRoj4Q4tJL3LdSyMtLjr5MEXjcns04SLBrAiM5MuyO7wdj7eb6nPAGfOQbWU
7STYZdXx7PYftbBK1bC7hn5zJyrSoTXDI4g6fHJnZPQZbE98o4XvpTvI+Vk1JO1t
YcywWdsf3GycqYVE41zU4jCaB/w83KHG8b13tYOPMjd949kfcQtUv0nqiR5HmLvs
Ar+U5I55LjCTuznDOHeD7bygqliJhruldgZbGwBdRl8DVNcvxAsraM+AlsEjL1ys
saGXmriVdSKBAUOsopIkYFmQ3I7doJcwSFCfHd6zQYn44ub0iyJ+ZcJ2VW6M+o7G
yZI/3fhuVFRUG/8Cz2rz1W2JTb81nscZcSa/0S1Xv9f0CuQr8BjFcubJYgoNkKKk
/ZrsL+BcvGH5Pw1miHnHgy6Qo2s5/jevGYu9b0GU+PZygYWp6N6CMXp1EemcB8Bl
0C/cIFXBsmMNRYhCdWqke5rZgMIWMDoFWSyJ/fVRp5p56S43wF2Vsa4LKj8SL+pc
gjkH0QrTuucsxoR3ZpypEq6cbQtdMifgWwokgZLjWXYdB9MfnDKIqFMk2WxDZSUG
tQ6Q/2nGYa0RXcOqTyWidIVW2gjXuZ5l7bD5lqmpVCgi5En3kaE1GxOXvLm3DD5t
ckxCW1pyJZhueZkKLIT47Iwd4IVywuI5/5G3ema6+7Q5mxsHaQ42HQciMThUlCVZ
UIvjSHXP2pgzyLAktI3cYW+d3Jdcqc7PiUIwnsfRmqFjQdoW1gdREarlcgZbl6OG
iB8e9Xqe/HLu092RazUMVhMbbstqhZKmH0d70ke9J6vZj+pvtuvWmFCMOqyyUBny
QHMEyH8zIE9mPO7z9XnCWVj008DDTk/eojGKg4ovbwODk7mAARo9zNjQLz0Af2nl
4z4H5U1/+3RWm8gzZ409yJeL97BpSlnqqQxdf1hhA6ma7mgMdTF6caXN2km12tHA
R65NIQgEE7RPQym/U+quqNud/OsV0LWfpEg1Eq9wLEF/cGKd1rMmeby+ndnlkIiT
8sj+9Xder0077oLLIOb6goDkY7oy6D9yj+3KE7unjgoC9vO3U4cQgnunJ2MQdT6w
qO7D9OWFmWHYv/sq/fEYumOAEsUptfWbrC4nMiXRJykM+XGoP5c46ra7quTjr2ns
gdvzNp4M6gouksWtVjY0AZmJoxe370Zl69nr5KT73Fe9e1klvsAGhbCSNVbRauAr
eXy4eIena7ks+zW3GZFZhSt9qMraSMDQ6HdphTPPPIMXML+ZA+h4CdZ5TKkgEp82
XZYg3JBrmbdnlAtQCNR3OIEuOUipvYE4u5cj5id7bmGuluii6b8dJqq1qgN9pYXR
oAfPMM62lLc+03ZFAp4NYVkLLbmYOKK8iovgNudJWPYZj0eHwZgSgMCdVHcTwiji
kZeAsHz5aeRfXOZwFjyIhLjcoSS97YLoc6zTwRuboUWo7knPaKOd+h6YxTW9gDMy
S4enQqF8PkvBoo0W49wxk4IssjcIuY2A+yLD4ApbRg11PwBvcPvglGsYj9m0dEtM
LEtl4pPlUy0q8OCMkz8tuda6MbeZrTKbucCCAERG12voprrAVkibn+ovMXCTTfHw
G/BSOm8VHjHpCOI2iRibPItVo43et6ZclbSPPKKpgXJNLfXe+z0tG819x5l+xyna
u3WPq44PeTUpF9D8bsiN9X/FrP2GMJ9IPLDCMOi714446KUszxVl0Di+x0N92cD8
aWGO88VJPxQL6r3Dm/zpW5NkwK1EXTD3xMQBZoA5XQo32uJ1JiCoXksPHtdEXOxl
qF7W/GM8qfql3Q0+5C08D/QE0O917djyZd3ID+S7/Q5SfWomAvNvehs92wX++pZa
oNrsTNm8anzCR3jRjf4ibPPtYtS2uc/OQAqXggmoPMZWXjOOgYHp5E8X0QBcSK3A
nHrOxoHAfUOppX+JGUK+bmjZldkOoupwP1uYVRbuyN7K5+Lf9BFAUiNczoTxh/p4
scw7eF2iuxsd5TORceFDXbBpFR1dEEs9nNCfHR53PGqR8Mq2IXCcmcgo5K/ljOan
6cYxMYvq5BOsBoWu9XoppWQONDwgB73tDrB9TCd/qP6sAhuV9CufmArDaSyfwkSi
jmwdV7WHEhxwjB28wcZi6NVlD+1vNCj+wg10q9sn1YvlhV7uirJgD8AM6mE+1Ray
hvi8CtHpmxHdKPFuDCemgm3Mri7YR/YLTK15uM9YjmfGiN0Qki4Vtaf/ucotmpsX
Cc/9j/Fns8WifGWlupysuBx+tA55KlDQyH9VbqEcT8BqPVDY/DcGQQbsLsO6fuop
eWKc2+fqR+OAo7PMf0u/WVebSernCbH2+M5bS3qczij22VD1j03Xn6ZLifZ6oiNA
KOwJNwO1ou4dXx6SyqiPiHcanrVn1/u93Zk0KPFco8NZwkpjkKQstqac78y/5MZO
5zcXDnUSW44gUztiLOPZpLozL0/qyoKEYsMv/KMu0/57eA5bUYrN/I6sB6t7XvKS
CbuoJGC09lzPmtzJnKJw+TPEd2fl1FApB5k/rHPJ+QB/1fR+g1JE0MVbw1nIlxXn
8n/cMl2gc3g0es9jOKGDERxWbZ2jsx14ntrXkd5ZYYap1qgIoxchRigA7WrfNQlx
h06Ea8XDDf22+Maf8bLo7XD8aAt1B5F1WYpAbgwuNcIbDE3nkCg3qIPv7/Z6QTo9
yJzu6UCIXDw+Zd/eLGQOTf+f2s3qsntGrFOzAIDa/KILSFK716fdYeOyiSPhTC/k
TUWkTbH8pW8FIsDHSYlF83A/OSs62z1ge9FlHyXhWO55M6xu3BTWTlXnIx1Lp/Xm
7i0FX0VdYKGktbpBw9CKssJUR8v64HKh+blnFdIVpcVgIlp5hdnI5fvTvgyTnqEM
75Aaaze8uL7280ENJ0Lsn+hAdn6LKHoCcyQUIe7SilX/mMwj0rsBZSulYAs08PYg
KD93wtpg1r5VQt/cIFjTGW1SDd1S4DPxNBEtcVlwxKhDwtkGKe85WEd6ux1SmNUb
eUPf3qqldNBTmPmc4Ff1wR3cs8soCjPV2H39+Q4WpHAdoDXK0XgnFH2O6RFh73hc
DPWNB5tvk1xqT6gvxKaYUAIwqldnKOSMJwtN39Eskaqd7O2SJsp24HW9CXhqY/Cn
c3/uykN+x/8hCkHcQwm/mGzUXcQDbbSPwUzi0BSo9ok1+gVppyKouTRzCg5/grea
+89fsOBZPsmoTARcUZ/uEWsIxBVz3H2jWQaDBA5awf2QxxydGvG09nQSlLhk8iup
GFMAgikv+nmmbeBabfx6iqqcJaWB5aBEPz6LlUhPVPjSE+Vt0HTe4MUWDxU3JBrj
3BlyDnX+1SxfxZBA2HHLKFaoOIZTq6Ws8VLzTxq9zacP9Xl0slnxAJG7agniRAMB
cdHOok2K1028LesFmzNuONXbsTVLQH3zSYvfoagLN4tGFSPOkrj13gqpAMfpNzM7
G02eVy/fcwApRMzSMMCNZ4bOxWzfCarP9NKaosH9M/nQg2vBGH8qT6sqH4KufWmj
AP3pfnnXC54ic8tet2r4Ydm9tzIBAFkFTkCIo+ymI2yhul3UZgX9ua8ujm3PQRrp
oIEoo3fuNAiR1O/mTum4nsqOH+oAvdeMdLwyl2C7N9dIKq9jDchBaJ9Le1HEM5Pc
5caKdgF5R4RpSViz5wQ8WfFxZC7nQQilPmzooYYGpugcds+V4ptsNX8EtUNLqdqi
wXoQCFz907QktQGpb8hvyWTCbcsas06FsYOX6vB7NC3spkIRKm9v7N3VCrMFiMLX
Wpa3lRG7QpKw5yQevdFdcDTjqZGVVBDTtuUr63mpRGzsZAGbtOc3PjkCxVxlbwCH
nRaaHtG0pB/Kknmz3VpGRYEJNks7pIgub9DSnfZW3KGXc1ki8LOa5N6tS44ScxO3
UL1icgxVwIZvTipgAxg+u5tsrNYpoYOp9aQNBW1rIIpbUdj4Sz1H3qN889C9JXa9
L/uw2/PDiwbfezk7i3AnlaSLr+M3S7Qv+x59YQHrH3iFlm9eIzxm6H4OpgOWR4Kg
w0I6dsQq3emfwGymn68jsd5nhDMYdKn9HJhLA53oybG2nG5gHTZMGAnwzDVlIOri
LXMrWuMZ4zdmBz9Zc6Ed9glDpKJZ+N94n0a3f4XcJ3OQwnqqupCM9Syb5Q0yrKMC
HysFlNPw71zzlaW9QfnD70DUQBlVOrUQH/E/9NGwfHnfZHMWZjtEwfcEyqEqhUxA
4F7etldcnWmsvJ1K8eN4zBW6UHxivDB3tLJJVeTIL0EbU8QZFqIoTfa5HVhZC3RT
RZcRdnZyBQLaFKO1p7IW3aYnWDn/TvYN6GgEqJvhBS3JROafy6GqqIzC62fvEnha
jgYTvMO2B763nAtC/M6xGgAZ0rfiiVRUB8thL5pXxH/tvE6CLHMzcjxSJkjMgIR2
LkEHiiIQ7ouWef84etS8QGP1wZC3rRGHMmH1VktkwkoVMsGzypOA0DwUNzF4at0o
JZEeQSeDZCOg4sWC0zw823OH4Zj5OtyHVUP55dBHqzR0zKFh0B1IOYm/2BA+3iqY
cdwd27jjK73iJP2t0hVlxwYOV+SswdYGaKn9WfYuGCodpsAFJRKjzpwNBd7O9GdE
TxSnmOLQMZyIw/QpB4/fu7FRT2JhqiHDPm1+u1E3J926l+A8oD+WpI3x0hwZs6rB
zF7VrORlAxOPLGt7ttbImDbY+PIuHBACPbvRvhlLIyAl9Q3dtfTs9FFvdkU710rb
ZYKIxs3DzrbHzeI4g9GZ6CsGf+7hfA50jE2cCzDaVdvy9sPm5+mL8GnGG9Y5wqUj
P/NcCrjduWuabw8y/W2CWLgQYCsYdewy78eaa76qIMWpS97EsTjD6CkmyVuF2WNO
hZqpLCDbaIl9P4thQoi3ZcKzO6c9SRWqSQoMoRMV0MntxP+wWvk7+glrfHNBCbP9
B6n0Pp2kCQGaN2DY2ZW9EeN1m01zxpdwSyCg1F3gelSpnOLdtYveHEfEsFqhiHdd
KC0ilW98ThyT4a7zN2ussPXWB0U1t6isQbUIPzzlxMAVzRlBCvR0KvC+Y5Cxi0mm
lEbPnNJ7tHpvPmyzB5P13Ex7W8B05+ENEs9EEPdXOh/LmeWDsSq9a0GrlSVK4xlt
1pt7sOS8flPyn9sNMcRkww6l5CLrs/oRq8QhYCMNMecLVTy1u/jeVhzN6VLr0Vnw
LUSHz4YwKPq4U8CMsrstUpmmYkTz24gYXFCI8XmFOS7/p9ZVZK45W80wzXOHfY7T
7nYSrOMzWkGx3QWcKrnyDpCdlK0BnqF2cHV9DWMqcPLQ+axRp5n2PlGE8Zl8u6qT
fYLki/9v/u1VcgehIE5evKlqE6flWXdNQ/+M1/Lljyj2vPVZcazm0jHbAp7MSlWP
HEhc/R170C4U5mYIU8hKSxXj6k+eINrjBvtsrguaY0QMMWVa1geZcR9V8w6k5ApN
FTcdNaW3YJ8RNab8fePyJv7xd7AN7csX9+1zItp9rj9NAl8KiyHTGixELul5ie/M
pJaC6tX2+JhrrQQYASp3WgJaBZ8xmSja93s6o9NwHclx0DNAgFM9O8b72XjXaJEy
z4wLl7kDQGjiWf0PTyNwBZQ77xLFYNcI+aa907rWDHWiba0Ybnt3FCznUM5W5Sw5
JagnBHv689wPL7WFEnnuxEfaYty+13+WtiFPZsZfJiqDPvKxOlArM2AYqPPeVuOH
FUbCFenpFkdh+7JQcbQYB0Ejxc9MhyolDbKX0Y2ipEjf4PLCY60jWCgL0icCMkXj
Cmh5/fWihr64jA9XAlpffJeO+9cjD3DudU4jP91RwvEb98wsq/NKQ7lOSpuyuase
J3Z9khmarByYvg0KbxG7oc6Q8QX7ZVnWsPShFa8jVJ69dZUg3Fhshjqp86B+WiX7
DiifAquNq3nCdjAJnJBldoYoEfztn3fbFNUEuR6LlH7zRg9NIQzNAk532WK/pQ8k
6EhQJoLsqyzkfXG4t1NEj5YY3qJ0lka2xZxf2iWvpfWCGENegqNymIiVG3Pv3NEq
0L2YVVWmax75AUagy/4qUZk0AW2RE3C5Hs32CkZEz+itYbKBW079eRlRMEaSox4O
vyF37EgU7lLvTHuBT0wVPLwBbIUDedYz59W6gMZwAvMtf5MwHIPHuCxTHz1FwDPb
xnT1PwTp4YKpi00lkvrnlgZ+h0C35QP5ylIgaDaBBq9kiZ/fFV1f2LCrZrcWPr/a
NXkzpV3sTu6uBwd529odoy9CE8ZHqLgZ0sGq2nMs1xBDpWB2Qk1ylZboE/oyCNH3
SNXv3EUZpOX5onanNgeTa84e/0ma/NA2hTkwnbhV2Usmp7lOONW8FItud1XrfLEV
EBFWtUbaMTk6uXycIVqcgEZcqQ7d7HxzRQswTSOy33oYS5qBiohRYcj4JYcJIxL7
Ei/qUWTiWkrB/hHNn8QY0tcxXTk7Q+qEQ8ke5TXPJkQSxMiLWwAKRP28GRJbRWLm
prWIMLv4oeL4+vI7+ua7TnJANrELZNLnHSCpAeIMc2C9D2a+mz9i/0ygF8O+9m1z
yXapwEajRfoINXEL9qrnSTIDHribUUKmJGDMQAGABdoqi7UOplGHACXt4eJEXuCk
zhD3mMHJMq6JthLJ96RUsjQFbWZRTxPXNUKYlXBAAO2AgURbbnz9Bfom5h6fx1jO
Dz9rJLpGSpvEAEWf82cRmiy18qyqVMhgI3w19tVoIaAvkkTJekIIpYjZoIlRlO2s
NG9zPMUsKq0Nfogh7ucvAy6vDXWFOLg5g1h6/cRckBWnOxlU1bUi76ubMX/rmemz
S6C+fbbjKWyT98kV6lP3z6k/21ypDtrP6UyRMCRidIAa6E9W/6V+ZkngMG418sTZ
bDDJZL0mAal0afBKwLM64C3VNRmJnTSl56NNiD6MoE8Qif3epN1wei7JfWV22atO
iAEtTO85Jh2l9VVJ1Hr0M38RcPZiJ/dA/6vM3M/LSuoRVe5iSe53xYuJSsTm2Gta
r9BdYbtK5mxwu4qpcf0kplB5gGIPGVjPyAmpWBFKbFqkxmBaOVmA3w2UPj/yg4ov
v8oNgT9kLup0TMBN2uAT8nfofQtRhyB8+8sA5RpryGAGve1pXH1YHVFY6O2yCrlF
0+lQac5MfU3Fd6AK3/BxmO2XMhpLtm71ojvJ+UZzrKWGwWxt9SqIim8w4peejIYB
n3NUkRu2xYpn0ytfjNxfP9htcASERDx8Ja7vjpbpW8LWVfVFdKu+i2haJD8yVQM0
AATzZnPYJVZFd4TLCowcrPtFv2e7RhGMB6r6iUoFVloQkv3kYZKdvCAXyRpjloMX
m/6UFngQWCsvphA8PyUCQEi5bSF96kmOL/Oy49RrQ/5jHqEmS20W1uv9oQrmcGoX
r7viL2al7myUHGAI5C4Duzf5uuSsiDMo6sYgDgIZyqSYL6R5qUL7NVzzqhC+mv9h
AadQZSi/NcVDResq3bdIPxJ4GWh1/8TyLkqSptq0J8dy//AgtVJR8Kxvi0UAHue9
SC1xASvu7U1TlzR0H14K8Ml3KjGVnHUmXW35IP5pRtbmu8i0J8Nk56Y+UUiPBrpr
VtY67gYUtWTCjZ6JJM1udgxJI/hPoPGB4WMPN9daqKuKr8y5ZE9s+zAqX1forgP3
9o7QjxZoLzNJmb+nNb09Hi+4mBfb/4Vp8rZxtV8z9ZZs+CYyXV+4m1nlEh7sixT3
mfsdGOtR/Eci2qHIXPUVkHOUpmofAscyVWAPIvkbCDMxf8brN+Aey44e+x9sf8VS
8qppRNlJn6gI0woXbZi36FdNN70eesYzSfc+X3c5GT8u2fSd0dt9apwXEVoWZ7gO
MPkvPsioACTdY6REI42je+z2Ny7qVRYrbDZBsTTf+Gp8kNgNZ1UwJpHlWJj/Q/Go
lJxnrgKt4KqVua7DFmugOEIWymFVUN1fc/wgNV07z2FMJ1JEKYBfI48NrqugPAJt
++SzigbWBAGyv0Hx8Meg+KV2ISpBhiHnBJ0kZbMAJ3EC0aegQPs532fvcQpd7kTq
z76P8v5xZp0P6eU61TWD2webLgX+4MatUaZnPdKiwW6cN5w65fymK475M44v9lew
ZJtK6BQiJinMnUePMVgaBFiIBNngUgDFzg60tPA2LDOp8O3GCxF3ySyTGLoiHETk
KYtvd7lv3RGc8IuEJGanJVT0sBDoVdv3LvG41mwqNQb4CEvUZ8T9NjDm9V+/J8Zc
kGWaRt75LDC+tUE/9qTn0JBC7VYe/5IBCsT3wsIAKwE+AtNNb4T5mdBHeN7Ph0IM
irUjTtDLXQGB8yQkmTKbkxW7t9OW0wR6KLlRBIh1v9PRbIv13XGqKJwL37Cuyvmq
FkJwlZya/nvVyqUaeCGldqZOHSigfXtydrxB1LI7XnuCSs6d+l0hGYeoXSZiyoCr
xGzvfN59pbNME/j/dq93+zMDeNYX1fuRPKfObWjHfXYKgJl+A8h/8fjVSOzxxSMO
emmmwobjch3KOegreXxT8zhCiwvJg/LzA+4fcBA/0CKt2QvEq6uzwtzROTLx1/E6
KkksSEhYitqohrlD2RPmS2eYg1yTnXxrG27viQHTOMcF9znv9EOMNjNTOHI4MOlW
4WASuS/8FXVDsWHvk8JBJuXW52467v0mFu3XgMl/hSa8X8rrcHQg4Etey2uR0jwx
RPUCddf35f15xNTELRlhoRcsYuUkkcBVINzCbrlR2JrtlXAY3G30xICSnjOkaNwT
WqtKkL622mfatZTZzkAOfHc2fsA7cjXM6M7tgL00iRfnb3x+I1wCAHZWgvqKH+Bo
1Omq3g0WT1J0TxpLYsVxyIQsCXO0w18ssONqpaiLe5rx1ILlg8SIQK2PG/9O3nd7
kubhf5kVMQgP82RPSqWG61wNzg/ZsrwUsFDlfaQEYCTq26jmuHwff+oS7vSj40OI
U9dxk+s0zJxge5UIA/abICBgEBj6IKGF45pweymNmPcLQCUkBHRTJ5FyrNg+2QMs
2ohCofS7A6lC5UqolMl39p9yO02U/Bl6sEcK4iLFL+cF4nyaMZHNs9q2b4Guli4c
5v1ppMcVjtr62xu5eypUZf/0xyxeXhd0xPDfwwuPT9EA0ETZHQMpr17THZgHd9Jc
uwOWfNl6ATKT8h8uDl6GgLdXcNuHyrVbYcjzbAduREf1sgjfO7xDsoX33Lucr3SP
2VrnELaMJAloGmZbTab/Zuxz49pN+wBbNZYeOG+H1amtDr6pRDDTNRj52x7crCqM
i54zx58RtsF3rWotnm5lpYZGDHXS/TjaJDZ4qQM2nhIC9Gn2XrPORgvD6ww5AVyi
VSApKtWY8RUBrlQ+UM5SSU6p4GI88wjjI4mZ26qcMhRRuZLwKhbRyUfxt+9uYCjL
+9EI/KXtLZo3h1eSAzEtVyHidgfzGAe/YF9jYjFJ8FENdV7AqsoJC9nTZdT2k5T6
3hzfZ5192DVecT/im/xReoDlAhHCiHNlJm1DXY9HNJjup9a7PoYvNKLI62LAI41s
cIgzzr2AH/a4t9kwmDZQJeVy7Ee3IYdiDZM75gQ4OdDUt1GKvKnpJUFGNRXYKdMD
46FURdgNDTrw3JSBCRRA+19/Cg75uFviyJbgc5+XtOOkmK1Hw5kUVlo6m6bLUBa/
CQGLfXGp0fJtM8PauX7G+cBxWYwNR/6oGevyF4j7SATXatT/rC72Iuht/ALFSLTB
dg/L4b3dgl0+aOvhgMOQB56oTozq0oY1FBY9cqJkd/RV9v5/3CY+4ZnP7pctINXy
mVmw01yRw6CrNQWwB8meoN7t/Yj7c2pu/n+5Ihhc26TEXuEvE9sRAlI9iCYg5nAr
+0SOVlNJ4bU0conYyBQTuRAPWBSiLiT4oTAvWAtAko3ib5vFgt5AmuFf5PGpDY9n
KAvowkOdpkCbrvNdY435FJ+P4b52Kl+XqGXIqB/B9Cjr6vyxl1QX/J0zDp8iXio4
B8N+MN2LujbMXX4spDmotqD4fA0ihS6VYPWsS82ChiBccyJSQ4495Uehu1y7ENZN
GbUG/I3+yHU56z3BP1PkQvXeS9fksZccoPclrPz0ZWdlerH1jJa8tvIhnLIl3U9C
50V7nwcWnJe3DZOTGKo32ctbdAH88Ir1T5VQmyeuR25TxFIs++QNSulrzWbccNAa
uq/deh7eCVurLdtdshSWBBB7iPUmVK2PtoBcQ6WR1R6hrXQc1cb/drS+jUL+tWbE
e+n995OQ36WGp6HWsrSw2QywxBSMhSr8xHsZaU6Z4idXvEinElm4m8h643iHA1Kq
nZigzLgUE+6OIQkkSrpy/wLZaWTnZz08ScikJ5Okim0J6hDIxUqPlWQTpfCFH71n
t3MUlkj1zXtiCTsgXbJXMkDHPiDHGt3A96xcYH662tnFQjK7viBno/lbChNDGPIr
xHa+QFzxfKKZKtXkPXi2NrQ6fZWrtUXqdB1q3lQHmPKwJb9sVXoPXa5LG5i5RIgi
Qa5ieKrvlXeS37MF1jV2XStogOicwxAhepmU7YgACPjSI/UhLqqsE0Qs/fUNN7uF
l7b+jJcikjYnWRP8GQcTtIe6afdLAYLaLpZ5jfK+Va191nrKS2sk0DDL6cw1IAyf
X9iMl7BE7xk8p85O3duRWfcpuzH4rxQKqSEr4xcl1GUQWd6LzGNXnlfjfDsRCdzV
CJaFUXP0m2MJC1QXB/wCFNkZvg4wyATwyJUlAa+Okoa9VspRGg23Pu3M2uGawHNv
Z4pHwDSDFLZYl3FOA/WbX5f9mFvRzEhEA2ojhdJQvupwH5w/zc0sPuHDt+T3aqK2
Xl8zZGImHwROIZj+EREJt+lvcnoWU2ZuwB9P01w7DFKr8Uc8hqegwl6p08EmNHCX
ZwkxSBiCkqmGJaCaJiQja8o4FjZOjpGEG+vOMR0q+UFOPZ9EVqpg4bGZWj+tNrGP
3wgHlUVjhy2Yo09DEydtU1TCFdIP8Il/LsBhxrX0BucWsFnc1sr0Y3XEvtX35Gpx
ovdfWl7K/39jmZX2METaWJzvvhlamBRUplj2OE7OsCdxU2RlsKUTAAht947m6gdU
pk8YFqjzPexXhPmFWNvTsIIP/ymAD6oCPeuKY2/e374hbfrWe/XQ5oVkNjHOW5H/
ed6RPMy7OgZbxXa/LVzXzdwGm3HlwqyroRwmBIag+F0tvLNzq/DOnD0WMx7UAK2y
qTyTnfFvlcbSaCO9LxQkscX3zeplSoSHzsIEjOxqOwB3Gknakmmf7HBv1SK3Jkot
Fis6vrCAiHFf/KX998nKN6PbDJEFuMUGkUqqVS79+X1RcVow2qM/BCS9pxwL/8Lh
FjgcPFFEyQ3RoHDmn5oo0eA5JzlOd2+iz3AdfQvir4u04J8+NixsIZNTMYDCrbLe
IuWMHc5psSs8uVzopX7+3lHOGA+8XGwThKaG8t27UGzYKXkP7vHqtlj3IfGO0pLF
3P1zeo2xJuesDFAoMXwNb/ZRZ0VGuy/DkwDJFyA0WDUiPSPnmX4uDLZjqPyOypc9
sQ5XugH98NtfScEscCheQIzKTFjDUpPZivBb6npy8o0JV0tn58pks/Lk4s/9a9W1
4mBH5jaJ+thH9yuUwsv/NYkdXIOeP+RzuOVFT99/3oUvIYfqIAvXS3rGpIdek2+6
8hpWexDY3nkSMMBejsIbGQuaOTlS+Pv/jPG2flUz+z7/Z3x4hC0+yFR6IYt19D8M
/gSL/RK4pHeH/neUGA8bPPD6LeZ4zNsAc+5m+B286UR+HSVX2lgXhQq4kW9sv5VR
pcoGXKMAakjsoZhnecZ50G33USItp3b8U/FNY0iNoyTxJitd7rcXKimQM6lSAyGW
7Z93Agn5OXuIOrF0hb0jlcG55sRTUDlf+aeTLtQmVq/kfRXuwZhgf9DQk/sadQzt
XNyO+03aU5vEGtBCiP8kROUTLlm8oF7pOlj/7Lf2yJGxqEeuBLyUSp6dVc6E+fR2
BS7IHl0NaJJBDit3HCYx3+IkqK4p7yrd0Z0A7NImvtQjC21ocaSb8V+S0/YmKrPr
YIi5stLVl8bOwaJ/eihHgl7oY1Tt223wri9PlkSZp1nw7EkOGlwzJrx/cd1kMqKM
B5X0E86z4Pei0RXbXmLy//CrWetAj5fqvF+LDdw36x0jn7DVojgSSf075JSjg9ck
jm7WjReqPCIKzrh8S61PHrp7tqdIs/K8g0d3adMu3CrOeBJZ/rR5cyZRFI6I+e8D
/3PDaRBFL1Pd0copaoKjgOPC0u1Axo+eMMMyPAinixbZ/0W7Vqqmr5XWFFAjoY7T
XTVuirgh4eXoqo+DjWEsh/M4UxBIwo/0UjO7g2UYlGaj6EhP0aRFYXgSfe0uJ+nE
XyNmLd+4IAhLGp7A1/69Syffvn0lhwI/sKtyw/wQarFLBiw8Of1RKmJfpgxgRr9c
vgsEfWKqvGpu+W5RkHnjugCVgFbhfsd40lWSk/nfUetQWbrxFZJAnmH03ah7sG2R
Ooqupx7mgRhp5ofvBGTx9LaAlRVVLGzzZoyp8J+ZJVSrf0FYRb3bmZrshzm5HOGy
jEFGWCYbr/24PW1c3N3jhH6bG6zGwpUgg+KdgcZ5t+20H34O47o5qivGiGo6gv+X
p6mq9UF83trO/hpgpc75ADMhLipE+pfR417/Q/BXZFl6/fqMY8dQr95uvZ8Q7K5E
4CBr3oROm+Y0k5kCxmmf4lBFslwTLVypKvSn6l2USmItxrDOc14ZRj3kYE2oX/Y9
ZKb9MOBeR1CSbrXiIdyhNVBMzsUpWIpPV/wUi+lo0yIZuVUnZCY/2xE7gennNSQj
L6PDbsb+yfKG/Dl1zkckZ4/nXdrsBukalM0Zhfjop1l/WWhzidxetRqW34K2vlrD
emHDzVtUMnRreXCSWW633CXGighPTG48UvElqnPIDmysIwhEhRurLURXV3wKD2ES
EPrTBuT63Y9zxGMlJY4dB6F5ReYW4VFtYYyaYBb4qzucmAGR+LQ4SkMu7V2xoUDR
JVx+rQwAx1iCQcsDmvDhBb+wz297xcvMJGE79b8XzlCXIyQJkFM/hCihcfIlcHqB
JCmjS756VQyxMELOTu+dqa6ndlTJOKXibehRrNP/7zRC9u2XCjVU2fvFDtMC/waC
TBgVX76VYE2majQP9l1E4wHfT4szzFef/T6XmA/e8FwT7gpuWaGkhg7FmrYRKrOY
jsHn0HzLSIdZrNa5q9aq0jDlVzAz409zFhYfedMr57KN426rxHghwQot72/t43n5
9dYvgboKKoLif0AX/IsQd3uvpOlyT2RHFfoY0ibWtPlocuuT4VEKC8HVsSRt6NnJ
SlfgrSRLkp45dRVJjnHCTvPVkhW5xS+USvBgQ8NsVTnMhaqX66IDEdiZyULQ8D9o
xie9V/Vp06MSESWkQ4tZFB6O49qSj1XxIHGkvkD+Ab8356wSf74oZBmzDMDWnGeh
6HYQilAYI3zFrGIb+OSxDnWrUJ/Bhq2vCb27u8HUULzJF3G4zoUSaxxHnF9zLLYp
Rxv2RaalB4IiGHrNlDhBfW7VgCC3bVm/qVVS2tsIKtp2W0Uk5+AXao7xzcrb5XEW
kynIwVKyg5mnHV7D0yhC25dvd9AqgthF8b52h08NzWQC+Vp8SeKt9txPA+MDNJfi
YRlYNXhH8FIHtm0F1NcdQtxOYG75PptM8iw6ifKEnhJY4qs7UAtSkbCxVL+Q/E+R
2EU9AIjQZRY+Aqfv69CsiGohYEss15qDqXbUEAPE6RrmwQzHp+9c314Rbcpwlt/S
LclaFCnuWNvjyjxkXqZ4f/KgOEq7xDieC9KgknqsWn2/0scjBF0i2pCIMEfR8wbS
X2Fw8091Xz4ODdzuQWEMFNrAqTG6PET3iJAy2XQtuuf5nDh835dSY6rOj8EhSsTU
ktI67asKDp9STPjMQgWszVPYHZzg69sA4PJPVhDjRw+FcrUob0+5ZFIDiII7bR+x
FWkQDwW/XWGIGSEEqnmeGTk4e2aqYQyFHTLoiaMWSvAnqcM4iupMwGejQTQMnD1/
fd8KNnk0wMeRQotzgutAOrcV8/v9zpDfc05NHGF1syI3DJevN3zWAvXbC3ZIpMYt
aAdm7udZKkZlzw8xf2JcWcAUubfWK0DfBLTG5RNMtBbCljzYDbGuxxZfqqMZHWAi
YwfY2E9ulH5+NlF6w/kxzoBxk3BRzogGq+T1+xk5JPdAZjZf/iFgAI8DNIzVvVcl
CI5UD+Dcnq22YfgBt/Ve82yEE8uZ+BtwBt0NU3AnUeLXx2zKA06+ACQUVe8+huh5
2Kzb/8bHfHT3nBr9frCZFW/Eu9BRvWmIftP/sNLJzR8CGQEJlVMVaFnw1Okc1I7k
HYvQPtYPq0L9uQadAhks8AbaKDVoPmrs4jkSHCr1YJuiNBBUyNTEL3njDScguUTv
BWnOYs1Rd77lN/dprmBQJrCnj9FBZjMY6DqzFO4+3T5j9XRWCgAWStP7+SgzaXrB
ycQSUlFrCpqLRS3l7Qnnv6JbFKtXF4MV6duKXWDQ68YhHslOLmZFbTmQw/MyAZsc
q3NtJdXq4okqZ2a9ASyWE5YZIIgq01gJcjIJ0NfVdEtS0MKMr2nuUZFm2LEdk7px
DzaA5fdrgw87u1VbQsRS649iPGIWxn8xdvAS9gtpydqgXzCwthJ7malUPIBXGVzz
jEBcyTKbuDYXxiWrjVVa3CRhoI63uazrgzw8pYLfIAjGMDNtK1zRtfsiQRt0oaA0
zg+WCxuaBQ8OrqPg/yfJV1aPVzz1sr1fp8+eD0w5FwljM48MftszqhhHLqF6isuT
t5qoLp9NpFJ58BIvvomDHBpYwB7nU8j3ML6tNFC5YP0UI54RHu4VoWV6oJFbMUvD
oy611Jq23HZE8HxeeNxtB4QuB/6OacAG7v2x+6EVUwqoUm1F6xXRWKcXmfaLqnDm
b9FjBOs2Vy0Tm8brg5tFURsvl+mKbvWmWvWglPK2tZ/lQrngUW3AAKOKcG3X6PyA
HMtwlzu3WY/mHfWlj0phWn3wjcmghftribS2d1NhkBzm5Fs/UY2KJ13wppctQx8/
fk8HrqRfeCkWbFIrwmcSIUHdYobkqLx1Lc0ROAckxXlk8ylmVjioe//R+eUklnW4
gEa/7+Uc35T93jiR2miWJk4nC33dogHXnzP2P3ugyu6Ym7cTqSjsHzBoapwYVc0S
ml+KwPwHTGaoqf+5iLJBaIpfixlRPtxQh3T/rfYyT2uHDwaaAWiwsKwPb+lYdkiB
ibChZRm0V+QEhIH2dqnANqAKs/mbnnpEzgpLhACyG0o3ImouzLvJJt74wc+J/CT3
f2rBIlcQTfnY2oc8+/gMz2uXprgguL4AZKbkrfPK0lSc6dg0NaSSPla2uBEFGPZ2
aWEJlSrMpY12jci4XwbNFYm9d8AFZOtlcqAmEkrV2L7eGxofUq87tS0rPKXs6mAz
aPLIc+j3HRIcZ7jEGTVaXkQUnKEhuL9LgU1+6FzVsFLYhJz3d89ez4IPlcR0Jkv1
j99ZvpPRvz9L248pK2Gt97O2HuzNQI1yTq+dR6M3ahh6BfOcM8A0TnCs8ZEk3hIt
oFg1Lbheqa8pN08AykVKhwU7/o/IRWLeyZDDDgok+QPPbfjNM9CDV3KgSYsa3CzB
f9MpFPxRhGlad3siSk7CQCazJJTCu7SPIgY+ejxACGMF1dvMhOX5tf6+WAQqtI9Q
es5d6lPHd3CkRYPy7DRyQaLM3UwsbewtXsbCWiW2nuXOWQT4QEoqW7JBElklqqMX
mLZ4utazhCMLsZ/u2qC12/7QjJN5Yu0ilG3Rm0hV9PTHlFOjcIpvId5rlFPuk5FL
jlJCigNmXnye9VAy/UCWVtyxFFxEUOL5HiyZ5EuKNo3Z5oWDrZsfr6JtwOBJNBh9
iyvOffdoWtr5L5EloWqm9nknJMbqpNgvNaIPl/JC+irqHN1SgLE3jtjDV9DM28aK
4ANotsBvNAMH88N8x7vtJLrFI8yH22sNHrr8axEakAJm2VFhDlcYH9cD9ig0SC42
bOsJkoMqZqaWhFJ/2k/bBQ7asegud2SJs58xP1ZhfAyYgOBIZCly8c70qEMmDPrQ
XWFWHhh9x1/LYirIUSLpJmmFcTYq4fnmQirP3/r2M24+bZR+Cs7nXGKBOFqLP3ka
m0Jo5lpianMZocdZOIMMdITkEBquVaXfhey3PlaWlNCCM4/PtLCZMYBLLqNljhTl
5Ommi6+DZ6r2hiz7SlNCpiEbRzlOS5VM3i0CQbJI5mmmWN0nV24AfpXAu9zdDuLu
j7QyuEcJZI1Hu0nMENgj1M08PI+laiwxPCnVPJGemocdB/Ao/9AlpNDm6ARdNj19
NIlEXGK8JtROcvyjvYpwZXJBRxwUn8oafzgw0ShCbGkBDlajpfhcsziFLgYBXdsD
Y36/G6Iut4RZLxSE3GbtVJFGERhbbpSgnt3HlXJ/+gg8U1IkOqjxH07Y0h0A7not
G7pHwl5CWpb7uG1qs3TzuuS+hOlv6JeWy91ugWPwdYmdr7qBQknDJxqFRhLZqAdA
LhzKLDnkfkdV8MGioKL3rqiWSNKMkN6XoHL5ZpKDw0rRfSBwAmUbMPRCQi76HH8z
myprEdiFCGRqLI3Cv5AZr9iAnZuG1kfEQzk729uvSBgYtvRSs7iIqY2DgBwLq8UT
5Sjy9XzLXhx0mpMa07E9EvRk5Uc7/lLE6Z0csoH88i33bYfQGtcbe0AnuF8ddfZP
2lt3sReUM8ew4PB+j/00SZ1o+rE+yWBpU4ipMJbYS0bpQn5Tr0191SK14HQdvnpk
+h8UMCn5xmRMLJBK1lNy6/EYuid0J75Db6o180hFpGQofNpkR4EEoNXHMW2J63hf
N96kunDnACMwSUMYI9sR9n5Deyv132c9S1GJ4h75xBwKbMN4lOl13piwobgkGM5g
FjeEeyeyzVAeWMpEMlcXzfqiXKSnNrnAn7NdR28jQVUTWFbyvrIaGMIgZKIiOZGQ
xA2sl9p8ORFKfMU3nsmhvckV8bnNvofgBAY4Vcjp5QF+SwRVVtkXWXUBOqgyiOgw
1Kh3P0mIDE0z8iN+UN9qfCMbBm1lhmQ3rPCnYgpy2Hk7sVuucBEnugtT/BFk9Rr3
PNnKpNr7vF8dzOOlwtHmCavPYv+j4xRL9oHmvM4TVoNxXKUOj6P03/Iiksf6SYte
8ki6HdT99mcKel8lLKbKxQsiN0esPkGZ9EAK/9wQipWAgEoyehDereRXtisGIl6p
gQnysJRZwQDRxvJuaqlHhKqomoOkJVgjwupH95uvvq+qG0r8TeOsMEJVZQO08xAb
a6nhWygsbdTfw4Hlf/IeRFIJxSU2XBQvs5uk87tbicOZOAYM3EjX/SXb+qBroVLz
k3pWVPkHPGnaSVltrVxrNF21MzFRpD95wamC58JDf4evt1Hk2kIpZra1aYhK9Qal
E7tH3PxoDfGxTeaWEdTSkRp3nTPNVYEff9bmFGxeuvXThC2uJiHWzzptczRaVKMd
xi3GmxL7lmpg5epWEUh/Huw4uDWO1FihWEjOW+SuGrYvxQi2dHHQQ7vk7EJ/tnPh
m5WOf7JOxv8L6/NaKhUTqOygxQ1IUNixK6Ok3eXtrWP9yrF5K+yvsGhBGdfoB1P5
JbXEEu62JhnQwgDrJ7eaaggfLgWtSP59jL0VjhjZnh6v2nq+SNrnMx4K64PTQNl9
//XmQ6DnRyLt88HD1dVkjg5YtQWknjJdH0WXr9z6Hs7TJ9FAWQoasZJtMfo/IqgV
slwtR+e/t1LNxryWol8xOYHpwi5thldrQyTEWCEpDANzSV45KUmMzvQyoQawxQev
kqPaoL/x+MlXAEz1MLR3pbE+YqHnaG0FLBT8XLAcuXIyXtZ99AkNdCOtpsAD2w5n
+PFmAYLYtf6/bTrFOEYkqcvFxYmsw0gRgER/RshRgoWX5gHJ5ZbyTaoTlRfUl7vK
4GYcJCbRsKukVk/En/Qq8ITsOQpIB0bg4qEDGuLVno1i4HkY0pN3SppjezfmWCNF
SJarUAbgb+HrScGgGRvpCvOi3Xz0CkCEYCRI6HsXwRCJxWCIv1LVeLDOvugii1Bi
rVEjzxnajbUVIvzc094LjizAoBKFMzyc9CZRPSsCVKh4W3PwHpB4jq8tQwzBRV2Q
qBMDFM+A6c0jB3+KKLhGtdWzMpOXUrzWh0tdH5+deSq2BTO/fPuL8888OuOBRs/u
15ph0wXor6riyITF4/5KGeeRqTCb08f8WPj8FaegjFil/TsVXytNtVGJS1KZROex
DGvD0DZ1Egvoge3K1E2N3JVzsgrjbQuiu1GP2VZJRgf/CV5BfHhVg2twuOOsIE/Q
y8gXTQJKoU00eGYiqhYlfkg45jxbYZpR8Hp4bim2sZF9afAKZHEI+pMSgPm8EokU
Q6RCQjA9ldDYnzi3qlHWtCLPc3NVH+DTYShu+HwrWlvAISZCEp46+0jQkAqIjfhk
0scuapne1tpbAiVEKl6zh4SJKy0cZM+FoArrxjPxMzQUeGRu25J9EsycR2pkhO4t
TzC06ZB40TCsTXZhWDGL5xNE7hU76AcM4II2V3IPYyfOkhuxcN7hyI+baLeFaRC2
BALrH6Wch0n20rrS620XkIgbfFLLU9ItWHCj8kLw5ZbeuyXmjGZUeAtRoCQ1Fb4J
jQd+uv/H5PZFgQNAl4CSrh8ByRVAeDFMbVkdtc0YJBZNeuGrq6tNNgzGUqTDlZp0
eHSixxyn4zkESwoWw3RNqs2U97OTTL9EDcLpD5Jquuhaw+w6d0hccr+5G6KYB3IS
xW5D/rvEMxBEZGMKCSEKHlXAuQiwGZxIzzLpUV2O5EhDDAOyjp3EBAtJELS7jd/1
K1gUhIJHUZqy/EN+/+w0byflFkkvaks0P+hx7MLcNzNGq1SIDuGKAoW/VhoknrXQ
HvXJEXYbsAcpxzvROGtf2F+GsNk+N7U25i7VjsJJMr0f0NSuvDjl/9yrsn5M0Hmj
M2MHshPorR0l16s8RXC+W/bDSnBgj5tw0WESIfHWqwFZIkojq0ma7nC1llXQMAcd
YEbbZneIUkNcmDzLb/2LhDmhFLIu6Xrd6+D5IpccMC0WFWgxWw69kPIpKhjWnhBq
v3UYUOdw8RCPlG+jOreLJ+mCwrAO6KPja8moD67IKN8DAUl9OsD73c7ozxWIzKvt
4AF+x72Nj7fQrfkqBvg+nXQImZQGNG71ueahGiNwbumYvha7Z4OHXRVcI3MbVZoP
KliPwMH0OH3rSBrwICdKPLMYWc18O5Qa0InbC6IGJ2171tfzuh8ZwZzaHBEp+saM
CbEqkDsyCcSOm33egPjsostlkKLRuGGPuo4hURoLIGedd1kwqweE1CaqvrLB8Mc8
xx43yq1GFfmRwll5LOnTTNMs3hE8o9rDPkoV/OM+2+8Nwu6ITt6hzkl0E0KikAA2
QtC2QDEEGEvMatoAB06jn5xo1kuxaGp+IlmJxVvYLf1HkdS/3EAuALC71M3ik6wO
jSVtlWpRHK/WIZdUnY7FzYFX5QczN9rnwGzmrIwPUtYoskBGZECXqt9srLwDM27+
Ju9v5W0Z1iIKrqGLkEqfaBbiWiQuicKv5Q/TFcygui8Lc5Qmlh8I/DNOICMbblvL
v2DDLLof3CBDBt7M5Na03SmQOH8tLtZUwvZ0CFAJ5lsXyFNxk9StUrd7mv+pGBBt
gNf2BmpY6VE5dylz1skzxS6GsdlS6VTev+6ALm4fy6FzGCMxmQDwUxS4xl/YHVFw
6qG28W+7AsARG7+92SvBk11bpAKRcwjKLQLs8o4lOFEOBZvl0b9Qupm2e7fqAyy/
XPyd2RzfyNqlyHV0mBGudGjCVZ1e5L89GCK2NPHKJIHVdpXhd70e4xOp3ISZhBgN
4tBoL9RvNwBgotaULVUY+G8VTg6riW93ZUNpXBQ1izIAb3HBgQy8TLQnc1H+2CcE
xdjtmG7h6mAAeRJRV5CC8STXJ83i6Cu7nfxm4bOq847kTDkByt0F2Fb2V2610t6v
pa3CD0Yc2wuPD9kTBbUlYbfLxjB0VNtRbXLyX5LBLd05BEoCGzhs4IhMYOVV22oH
nWSRGhz2GsmDCAcFNp+I3O+h/YxWd7fXxXPx/9fwI1d8PX9a0ZmG99LhfLQo3D0k
Lv3vauqi51rE/l5eHxpISTBx9mX7OsKaz1fO2VgWTNLA3r9//8/y9hON3NYiUxrd
w4qwbQZ3dv3YqOvqz169GIYo5gjxy1WBgiiuMTGjQqbiltF9Q0WQztoNr86045bR
IzhZeAv/+f+mKmfgRJHQQk9k8MG/SKuVrgoYCnxvLvWKhH2IeM341aZepGLNZd2/
xDPZ5umaI5HCklJH5BDVFx+P0yYgypqV0RmwnM4GohhiG7eU0K1snCmTi5V9ajsR
B+Q2XBOMdcw+wwZLhw3z3vUVrg4mjl9ZcbohgVMwnnSSagTgp0xFDP/M5tDNxPXo
aTgbP6N8vzSCtCkk6l8E2Sm+jbOVn1fZRSfJvpVuqFdhJl2OHoSwf3X9/MdNi6gM
9DEK/icfKlHwx9loeiQXZWf6AViCdm/SQcS/ctDkhliBy3vlRT+a8r78LtQbfZwd
EtROwkaCoO18MR9Q/osiTgPWlFOsWXR8pEeUBlzKijATVEwxV1/F1lSq/LLtMGfX
kftGn3VJQ2LJNKP8JsxcUgzJkjUELvxxpp8mfbEM/YCqy2Jqv7MGwO61VTqD9Y9C
tDJp727Xq59FtDbk3JVYFTtiyvLEdhAHZ3saVAmrXz3B8OfQH39HJPcF0b+MqUmg
J0AW+SCOQcJ7X/9zX12CqJJCLhwL4hloslWak2NlrcaDH+g+k0OtpGof9yWt5riM
TdJ3l3jJ9nzzpIp395kH7YkNBMGFG+76brRVVlvTb2j0CJVrqx5BHZT7t5iQS0Pc
wkM8WRDTk3R4HP8+k0FTlei9Vd8NcdoTicXgP02tak0zCdQcg3/HniCExB063whT
bNNqKlSkAZgfno8ouYgjp1iD8lq3zxUVFLUoZHGSikpJbmiEgyu/8PJ1J3DUbWpK
vVBJzfiw/wG83970M/jTPs1NUzp781AMOT9fq/4anPhMYmfIZY9gKw0Kxuj1uQSu
mYKwOP1ETy1B7PmlqB36m/rpiPBa7FB02WRHgd3KkzvxXnzODa2dZlPhm5he4hZR
PwmD7T1dXZ+6gtNuk3y6zoItyZTq47nglb05GVzOzQtcoFu5hZNQ27KG0Ha1XER7
ti4huix/CJIySu1GruBQGkbeRt/zAOnPKb658u2GIRK4+5uQAAficx2eQ5iACpx0
A5/LbcwkpbwhuH+C0HyXn9C7aO1GeBfkRAIiu44mQzfiuypwtFx3mlHiso4PPJTJ
vUym1LdSKNeQ2T1h6xjwRGyTHjy4JO4age+Oj5L5pzjXiCfDIwkgcrOeDe58xwKI
/m5rxvFM8EW6UoU577eASABSzz3auDNp7m0NUFAgb/mdrGfNNRse8ucjXCwcBe7f
4j2ULnDc5WBiZRIffV8pCr1yXy+vNp05mh6ZNvopIu22tRuUcywrVcKnux7WtoMV
pWIKKdzyvD1yZfmgwpsMdr/1OXkRo5OakgOgbLmm6FCS77M8PdPDSKjfNSnAKj41
JDktr4zJU5LX210Zkviz3AqfAOjCGkSI8AQfHtUBPkBHnNv4CR3pFmzOQzwjB9vj
UzxzOkHTV4U28YRrCQMyjUm+xeDNypMgpHrMdsTUCdUEPy9aa/7jzsL5DLGxtrVT
nCnXhTYT+aGiIAx6zAPQUC/FEhxdzanMPsWYUdQwHj0lQmhz4X+Sv7mf3c6anhCb
BCTRVIUrIW04V1tqHJNmKASvWgFx46V3AjTaVNe4zOATOgjxGq61x9RgHG5Wqni/
Z6qumPNW1qSnhRyj/TXg1eveYJVzCH2fSQW7OAfc9xnNMkGhQCZcjReVG4zffy8R
1fZyJkfvBNYQou/upsW6mRXmewEuoVWsjJhQK1zzhjXOX3J/F07zixGONKTddrTP
xLqqTGl9QwZrRxsjlJQDd9pZO8U/lksgfrdCdCUlQZpTflwoIQPQSX62xMRi6dgy
pguhvnzT8BGb5a4svIr4gjeHnV09KwlmKRtNMFZwXTSHFsE3RIrh477DjYKp9rk9
pFM014RDJoqOwvYkRZ1hWW9IA7KsWp7wSRi9pVWavSHrqbF5c98v5vmheMDylawN
L31AZNPqAjM9ecSMINyzVSY/Blo42VS1tP8K/WxLXTfTSA+CyTt7U/yZNCAt9BKH
6W6RExNymkohmZzjKxTPP8du/+BCMQsilP3Rp6dk5o09HwwgWIH/WA7a2PPMWaoy
/yCbhuapfaGo0chuYGvGSBLzT6V9TIgYcWsPOc3qXiN8IvGV672c6FAd8gsFfxqb
A1qqtRkdp0wY0J9Hh2gI0csP6VOkoxJepufaqiG/vktVBBhtNOPFjDV/OLFJE+BD
8DA1E4z0dyPdVxFfDm7+iCHpa0Icp2gq9Bbfm5gN/e7Abqmzy2Ld+SoaezWu/Fvw
596fiIhqN8QCytJlWqjQ6M9Mxx6Er43RtJUOLv6/zwmP55q4fktvnmeMblUwPeki
LE/68sX5PXb8fhBmi2bM190ADAjccIecRPSWw+WcahWBk2EmXV+ZK6S3bDHVwJkc
ufvAWxYbykiEJwKJZGPiVM0sQcUjARsq5EnsOpY8m/Ab4l6YsS+xu07mU0hE1toU
9YvH7GY4Im70+7NhbkmB5ZcqbKIfftDEUguGitsH6XoP/iVHXwK3yHRm7zW8gSUI
A42nA9WVjH49UH7+ACDN7C2e30zmXzdzxJBrwwoZglFx/jYhlPkXMOXANeZhNDiB
pqVMmXBfwKNbbX240bLoJm+fE+QCNe1gDlX2GaqR5f1flUopNYmKfFbmGblM2Dt6
WhpCPUplUg3eFvIgY1uU3VSX/r5c5TC87rIVxXiiKcgLyeKnfXonZHEH/cGPIMll
V512a3/ld06EHIh0OAjv88kl209s5Msq1JtXnSLYlty50qR0wRAkr6kr4cq4Kjq7
Z32Y65NQOo8HP9fXQo42JDjOCARl7eu8dhykBTL8GGF1T68gobubRcxPEj2NZWmV
vwlIeLT40MEA4g2/fCo6gNimq/SwjDKa4mC22ig+8BPml37awnWYqFzIAy3Qk+Cr
s1VVn55GaIK2Si5mrMD6lrlFsE2qnyspmg28CVP8wVZnaW1kvXOlhbtQzQjXR0BS
KrYMEHe9x0/2GEE57phMAEEkRQWVXllH+Ud4F2stIk0zc6fAkla0ZN6UWWWmAKZL
mrtJZIYKzFimavPUd//Lv3c9I+/aYADswUSOmzqz12xzzGT+1GnhUyM3IlUZsm79
wPsetUp7PZA3tplwCMAhYm8A1qLFWX/eXfxokZ4M43aLWuS5HbDvk8UI37uC4XtG
2jP5HRoNrR9rcT8bJZnH9HitO+IDDbYcDE0n33E0qCQ5RgHsh+FOV+d1OHjHtRMK
scpng88Uv9xbThC058H0OTxym9dA9QocIgA30WIFWrYAMvLcZ6ETn1jv9uLu15W9
k8L5oxVetlRlZn9tb0VYt+4vTJO+pYSGtg2OYjO4RtWmyx7jFalgT9utiUQlJKrM
uStzmftWeTJtYQB32gb/DIynq5JFSZTPBaLbEujFJ5uMd09oV7XWenbev2JzITU/
Xt54RzH4dKI8JLgS5Lc+FQJGbLa1iMR2ykexTMXQKQxqAsH7ZdPrp8376X8OmqoB
XifL8f6NtODw52xAHODXPCccaVH71gQIsHRQidInMtUM4JhR3TK0iMohn+AJHPJ2
3yK0YmvtWpZG/W8Lv1EBUzZnERQERD9eicg6gO6Z2cZCfzJ9Je67bcynTOQr3mT6
GXAw8Pp3F6w0YdA/3Fubb3Gr8lVvn309LxhD+Y21VbWRJm7RF38MF+efNID9huIt
7xVBNwkA5rpmS6keDcL4g/UoPbXSFRwEAWeEhC/xaL5CS7PTkj3YGRZXf6RWl6R1
jqSM0n/VAl2mBV/niEqQixdluhv5cp/BcLvvGBT3KfIEF3ZecqDMQBLOiWstlFxq
nM5DbuWFYGANZd5R1PkfMuemS6QRwUK5kwSu1FdgbFvjJkoFpYkXNYVaPgLqUcVo
CtSvdz8Y+Bl6ud+ChWjyNsYGPuPqzpuRfkVr/ktAT3TJpXY+jRIeMHgl+XpcSrKo
CN9mR7oVIoufrGpbBCgoqFOx0OmHywKa9PmdHjan81phKL8ZSsydirtj5jgqYGwv
vIBJhqZv2/mlGDEYwuUpi2micXKtUug7zhUGtOwKlDEZFiLXCM7130UPqMT9d9dk
FJKRDljjQAV+rXviH2VE3yQguRe6Qu5LMJI0IY92UNvX3zJe/UUuP+pcU+DlcWyG
HNj0VabuNX0gVrFDW1MEqPJ9Ux0rPbj6gj7ev/Cp/9RBre3B1LOLVpDUbsK1SHUU
4+BiEscpQbcYsq29N849Gs/cgcOGHe+JKbIgspkjefg7Tv3EZEzQ20dOj2lU6GlU
bp/qbUMqJDo8nHb6ydNXkitBM/yneUdjH2OFCdWYZM9OvIZEfHwdBUuaiPC+Rupe
uUXFURDfNlpDMht6bP6AIy9+s+vZgqDWfZARbPSsx+RxRhKSJ9NJoyozMUZKJ/fe
ddTuFU0YKaowhtZl0It1SMvpCYFbefslM065/HDDJYTlg3PXhGZoVveSVEN9tpI/
cqvjxkuNwALmeXB9fwbHgJa+t7ekGGHru6fUipf/AU8MjRjIygpR+omauSAWGKVt
waqDwnbB6ngvt3b+b140IPJppQNMzHUzlnhBFUK8YX+e4p8r6ctD6QNfOowbQ/Eq
ks9cauOUBfsx9YF5/cOZHGOcH3uVTp8OtYf1fl2IKsOr4b83jM+bulk6gTpaJYvL
WeQQXWsI4Q5trq5zG4BdFYdC+q/ulE6jqRFj4ph5ajATUKphBaIhZbAdDBQexE7F
i3JX6moxEmDWjZoF9/G6qoFp6PWBeGERfBq72n9NsMI4MzW5KrmUCVTKiixLFX79
fOnXkueNM5xtzVxRm4j0aptEsCInBPFFHPUPlRS0vOyIbvO/4Rnsxfh9Y0Gwbrxv
2TzxFE4FagAGSgmaXWKK/GAOWUJL5o0RHbqBJbAtHTrcfEnbXcjvPSYo0g8OVfdq
8QBA8QcAu4Ig5+5/OfcCNxnztl9zPa5rDZE0o7NiBAAmc4kGRPQr0MEXjQvFRHgN
XnVOxBfRRTcJBJi7uxjni74nadQI47Bzv7W4kIznxyzjDNZ+6nurYmblldaW3Cqs
GM3+5tQBNHb9F2tT2WI6KTLHdjUP5W0RTU4gR9ffYvA0uezS1T7oNRwLEbiJ8SD3
0BUc4+thar8XcEBl/ruw/npNmJEuKbJpBOPFCEKO9eDLgdd3A3Yx6E8rgEbjLm8O
tOSwtnDzs4W5UQn/VZo3SaRiYt+rC9mW032rRhI7w3Ws7XOfnC/RPe5lb0U1W27E
5CzF0S/PxAPDQtwqIBXFImUx53APc/p6gFKzYSChNUbAgxH4HMoxNK/EFgGQYmBz
kgPrYHaLQlKvpjngVrfde9TYTdeuM8rkd/HOYluWNMl87t4mDnVD13rGajiFj+2R
+Pk008JiMT5A/tQQiTTmWyT0OjWoAx/HDgavHoxMVte9nSeOQfhtCIIXoYQKYN41
NETn9qlPWdj1EU6zsHufvlTJsbViSoDs+785tQ749O++PfzNNIWxrQPagS0hkh1E
b6zeCUj3WdSU0X0E03MeDU+W+eqS7JnpqTYr58/Kuu11gbMSpTy2L6MO8yEkuMyc
FZtQfwGuEGmLZhhhUv/DiPVuQlPiOPgIhs+hgiosIZF2NWpO41zXP0NOByHkoaom
/ZaFpF2LmAhr3G5qJkeTUn2SNuo98ZlBfFvdMCdw9s/3s/FvL4HTg/1V0P91qsvx
KczAtwwIdblYJG3HFijxkZVRIpl5TcbY4aIv7EpirQESkZZEbFfK6zyN7p/SufK4
hsXSUnjYAq5vbQ80qq1EkUV5dY8wxVnVraIBdEB++GKEjW063pQOIxoMpDqNeHWE
+p8DtXz5eqLu/9wUZOUFG2neiff5KT8wnKiiGT7ks8hlPze8wtOmDj7SSMchsrYo
QEcH72j3ZQCXRVVkFpa8VAXMPTgZG4muS3HV9Pwp5vLzh59KJOqKct8y/k4lMu+3
YHPF7owaTV4/ePfffAdHuz+s+P46SVJ44F/5Bg/M8GXMbRYd/87wl2GTr37qT5WQ
QP5NGgxeAlKrSdLNEI/XSydKPFW0r8KmJCxzrP1oFUGygU3qqraBCzvBWhlJ8Dl/
UrttHj42SaK+2Fm+QGheWFUvDbT8dvr/COSS5OEoJTNIXOzp+k+MtuBETFfqmj45
sUyOgudwbjsVwKqGv57l433hVHmp3Ui3wNEHQOU0uWr9kO3tuv6UH9aRg6VEu4lJ
oK+kYXUPFTXvvhOYusIwYIRQkxwluaWWEoc2r4ImMnHSN0ndz7p+9gAs10uMk3Di
Nd9KO8wqnPWie8NWBFWlUtHV325MitjwR0hLdLc7GvR9XnCzFCN+i9iBSq1Yy2WX
vBvut/3DU+xnd8GLPq1qAsY+jXINuuKKUoA24MY55laBw3nG7qhhvTqM90nOzY18
urEff5HfJpmoJFe4qmX3DWoZ+C5zOMGMX8nqDtWzcb57kmUSHbDooKc4hHgAPcKt
KQv74j76PDCkSTW1RP9l2/FWeR2SI59otQ1YKT7mH6YRASv+DChRHNY7hO2Jz4Ks
Bp1Y3MsNwEJ7ajVdrT5Wk77o3f+i6lcGVPy+j8zZSTLDp3p+7E8Qr+EZPOGlvqi/
SGlgW8FC+EQlJUjjCWhoel7nODXXVjlxPVbrGjmmUbCHqUANBGHcQImd9ZqB1yDo
Pseaqr2jswwoPIcwsjTCIZirdVKeLPS8Uf0+59B7AYJgU7CX5vgK/7lHvyTmuXrV
uenNtz+Qqpv1Zdln1ggrOVdtG66HshH0Iffp2NJ6iz4XvtFnYtZaG5wcc5o2ZWrV
xV3mUoSe7b1Y7q0whMoCYYHs78nAMO7l70G7+Wjh5IEUHjvWntthRz4HisdjPq2g
wmKBY78GS96tOnsA/DAgUMjQd//b0S/nBtlSV1j1Kbwp1X07+wNLSB7xTzC9Xw0s
lkL8LS2XU6j24KJfrmKpcRjd62Qr3sLZHbgImUZSzE8ZRcb2UjvxODHi/AJvursz
I/cSoK6NYhPFcoEY6+b49tt6Xq4Lqs1N0oMGDeb1+FUVSkOOnaQGJlCo76E7BdS9
pDdePjiXCzQa5hzIeAAJNh+qSft2Pa7ISdCmd0J/pzLa9BVGZZZwXKt9UXVdl4Vv
44M1MozOzwjT1XZo4e/ZHE+ynbL2tQjW9BZ/lihSV7/GatMZQfOn1txDRzvmt+j9
o5/OeeARzYRsIhHnUtIDp4ck9H/CVCmxpVKx1cfqSTeZ4qc32oNu9q3gM0+I8Duj
Myyjr43nCsBNObieA4UAoYdnaQKdhAVL+qV0zmx9/gZAiQ6TxZ77ZHBrOLEb8Fvs
UPYY3ZqPZnnApCUfuK/QMZTj5Z/YPGOJohh7P49cIhNAxtH9oSlcLJ0mJ2Yh+KJU
bwjLHPAFxV6NUpZ+LWlTpHRQtFs+d2RH+w6G9pEtaLCCn2yH9iplSQrl8JCNWocO
XnG42NJKmwZU5RDLJJ3QzDolzERIPBxBTKe2Gq6eXAwg6a/tCdiXX261c2v+9aTq
HwRKIDAAlWBkr02HrbUoanCpKp+EI+eeAmW6kmTkR1ZAbj3GlV8xsyS58aRR3Q24
akhBpeENVq4014JZgQR4X2OOyhB3yXvpEmhy3lALXHU66NZaqPxNPCFr8R5uaCV8
sKSNBxTF6yN7dDb8GelwsQV61wHGSRiyfArz1wgifh6vKec8tykeWQyMNkMnQaKI
gm5mPXpaIWZHhid4HQifxqFi+JTie7wNjNj6c9Vh8ZNaE4LPztZFwCNB3nBBdwP5
txSm2ETYObxwdnTxlX8awpbdkpbXy1Nn3sdwwiblibflLDnrRUZK4r6MYcIOJzd6
V51HWli0Qj8UC4lQOEeZWioWIAXmMbaDNGXNRyNYduYnrXVNe01gcEsEArVdv2Qg
msl+s0FrgatwmL+grSL8SU4MSb8lIBiTUgLeHKP78+n6Lw4XxhfdURL9jynXPjxU
VnaJB1tKuDK49Crvhthh73oAWxk3KkPuiwtCRQCi6DLc+UWoVUjSCTsgUU88O8Xp
Q1iujcAcOAG/NKi0ASuIgXDRaKKbTrs2U/FXSgKv+ERwFNF0okUQRVbqhRPrxZGM
YhNJD9frOzQZxmxGG3iFgvrCJPtaUdPDdmke3Lm1gxAxQ0nCn9xoOUwnBiqJ/cP4
8Lp/WqJLQLbtb4dsaoJNGInS1jcVrsFRRjRxoDoLNtfC/+20AS+7FEgmIVND5KTM
mHV6oAMnshwjgDKaCJ+9HCWTFpNdxMcvByrO+Mj/YlpzPXypC9iUo6MG+v+0aynY
dn0ITRU9VQux551KYnoo6fYpho28wkA/rXuXaT8clYqD5eQlg+g0uLMiCuoLNrmt
q3munZVjzYPbYwQPMtGpVpKUafq3mAMDgdTaZ6OXuyVE89ZhXfOrk9ZsZ7TlLw+x
GLlsp7lS7LeN+ZZJYhfD8cZiGDpL8u0m6yAMxOnWCFAkBVyn507hlDLbIHgZhri3
EdBZn8lR+d2wJIDiAkxv/MHKrb+ahUKbF5lllQ0mUyYlUIUq5IzEsmSVuzanksLJ
PuvjmptTwxTeGRWF9X7Ct0rqms2uMMmra34X6LcFv6q/Encdcjtphqo+uCjmuO3L
0qKK/NHT6mHMFgMSnbGCieoM+C+jr6qaXE0mTsTvQ9/u3X/ZJxlyMe1ATD+DmNfR
t71O9tBsRBOzObY1x7y2kKGkv6HFeiHL79lvDUgqKeyUkuex+1jmvx8dynU09FQz
4rgxBiT+hRywIHW05Lq04GscX07D4oQ7YnaYJB5a6No8IWoulXTzRnxSzoT767EO
nvR1TALPbUuyr8kmY4zm8vEShFg4P1ZDseEkPfUFlJIvwxO2OSQMA/z3atTzEHwE
qeIxax0sUJlRrVN30G4p8Q/EaEtfFvJzwffvvv0LP+qR29qJD65BTUb14VDD8jLn
+jTALlqEdWnCAuGc1i8W4HN/qoz0kF4F+MTqO/6bAif8v4SSAajGgQQgV0yGSYxQ
7+aaU5f4EwpV10uyIntqLjH2MFveJAN/bdrKKJB4qMvpBlw1LgeO5SGsBXI9p9ri
yjjOBLeiRV9Dz4PCFZevazZaEhj0jDDWfwQjECKK2qNOxur3sMbGk4woZloS0Rwa
fzR+TiIuoTsDM/HOjE4jS9hrrbbhEw8ruTH/re5RgrMK6bSIN/0yfTL780mxp82c
KUC7DiVbnys7VcWWbp8bdow5Z1ScMA4fbJSawPAR2QjZ4KQWLWSPeBDNoWivxmyx
F4xYSH/leqAdtsr/hB7odFq8X/3MfDMI1tnPAfHisbsXEaHSoib9kPKYhHt9tMQT
kBgNnMn5HBfR2o/z13PjOq7Y3IgNuQymMjLlUKWIxLFLLCdOnVjxrKcQwdNrXhze
kfA9pEFuDzCHZ2Kcy6/RTFORLFYzJ6dnq0F/uqVBk7T6EjS8ciylw8VGJinMs/O7
w/Xodwv8V3a4aN3L3YtGydOVfIgK0E6W5fNBp+jeVGRGoLiBzbzYisntPP6GfQ8L
0o44sRdBPQM7WkEKT1flyzjMXO7zX+gKaFLwrlbpHf+Nvpqb8NJTmf2cv9+HnFN1
avWLNAVKhQ095TN9u6P3oN0XUhcRFf2esOEuDxnkk2uF4gddKIOSQZeN5cPVrcLj
CNaGVcXRXfDeCpuIqaWyLSEnH8tGAQnyAP5xIX3Mij0inVAcAyGInrbc3kJwcV/a
WKAQeu/JUcXD0Y0LPAlPEO1xeCM8ooAsBGhfLgRCniy2g//t1eQ4ucfewpZ/EYKB
7JnO8my5Sufsc86X4vJr/HyK96O4ld4Opv5+v1wWGLsq4jRIJr6RM6359EHsiDFx
AhU3+qBQbCEwLbKVrcwKUP6R5eeX0JJaZFKCz87jgGzy56v/mgE4reeF55bsq2+l
m0VNigxYJWxCx0uCJ7YUXfeZqtCdxQodCR61fL6zju4f3IoGB9osCJQsvbQes0ci
g1ugb2vPLLlODq++ny7DRt1hG/S4pLDoGyxYie3rZJBxr8JGnYeA4k8ECPGg7xQQ
n186EOFwJ3wykJsYxuR1ahFiGc0TwNgZRgo1J5qRxi7X1RraebDO9mQgDUySEYWI
nsUezQ8IkkKYkw1TQGIcNqY+aA+sdIwmjgfv5oFB29QwDBc6NGO5ECjRkmHXlI1b
1dUauHOR+95fpufWyPy/8xHEy4BN/1gdGf/PQ28+OcJ/G7E9IR2p/0qufV5yGvB1
CWRiaFEDqsKO2cbC6lo/UWD1rEVjQXOdUtPrdV15RDdC986dPGZPTYVyF0hbtGf1
aEDXd6Xkuv6ylvSoSCIjUQPNltMQjj4wHU88LdSYljy3QwpVkeyX6UEs5F45QQbA
50rbx9Jj42RhfR9UViL26Vfv/vsZBFAyNZBJaYzDac/VKsB6ocKZ/2xSUeMEt/p/
MeTqjtIP9aTOS12UhttpFJ+j8t8yrse9XLhrTdIlJcFi2F1fGUaEgFKs7P58HZBK
x0SMGNF/VHcV+80LM+TWcJOsb0PvBNoK/hurbPmJbTqscj0laxXCMo9+c3+Z5Ty4
bwhvQufD2XCaXkGwJ1+u8Qr7WRz3NsU6EEXx8Njr6pgI0wmnDtPvrJAnBG3w7kjt
87tBloKaBLYA7zWuq+/DuGyppwBJ3423oBk38Ooflv4atsMk66YDRfudctk6fyxV
PQN/hKcuDZxRd2yW4eWpxxAjvY5Ylq/rlPJXLt8FS/0TwsVPhRfBo/NdF36kTw+l
vuHVSOrjp1XaYa8d8StzdTKEkNAB1pIQoLj90S2LAc7bLcEoAgY9/xzqfbznPJZX
uPs9HEoK6418J9eXGeEZM7Z51e2wAB9Y8lHvhoCoHS15ePzn6flhxPTEMJ0ttiOH
z7NvYsdXBchr8F/MZzFqyuJQuPEx80Slidpc6ww3cM2wYvY/nhiLXkoK4EF05TMy
pUXSwNlBWzJP4AhzYY68mLWIcaMgOaPEt21WzxveAvLX9z8vo30qshfTm9mlSdh2
tStmJmz8GlUSLTwJjR68fYnYLsKuFKbhDli5xFAuBGwOtk9PhwyXktssWQGzq+bM
agR2rcNJtVsarBQEW3cye7FDWDvfGJEhfgaezbg5DiUP2F2xgYb3lFZeJdrmvkWS
EjkKQW4hTSAQXMsIR66UgpBt+y/I1E0fdzyyN3BghDMY2/V7NAxfGqffW+4DHjGK
JD67Jc5zFicM5o1vTRenhVMwYpEbretDUnpiUbLY+ZzY6eo145zpypECXV0kspB3
vfGkkrR+E6MFwihcSsubjxmkz1ss0Xhy+TSAKA472i+FQumn5lgNrKxCsqfQet+W
iy4s05QCd1EsQRY8YzKe4vOf95FCaw3pW/SnOXV+tz7Zw/TMCDiztTJE8Byh0gyT
cqbNAGl5oN/1e356FR6WjqYEBMWWfvSC23QirJuY6xEhz3jFREsS6UtGHCnKjmQi
szTxScCnnWWTzK8lTyQZsc/N5F78GVyC8lTzcxqxu9yU/o3lhErsilsmrq1rEmrk
F7yQYYlCfbM1brIDvlt6q0zs9tQ8tpkiFNUSkotbSdp5mSTToPFPGYd7Ll4/RjWN
C+slVv/NgBh4XKc0ijYk8fhkV4SEFG6k85slF7HXamZ4t7NKJZcM1coQ9XE7KXN6
Y0GMJVd+PZnhBSQm2ZioHHr0TEd9Jf7yrdmVL2Kek1k1XoeHoRLN9Q9+AzJtbklc
OvKDq+FDmWShu6iQWXOCXXyMYkgwnzfnL+qXs+K54IS6lrLqJyZfufnfeYE4/vaJ
4VNSwOsDybQe9yud/xVlUKjawmQlCzJ/CI+I9/MCqoQzVz5zEd70E3ztWTGhbH3U
HssK6Ht4h5gd+n9Nq6XHXTvaFLujRvxf1mjAE99B/V4p2pTzuhv4n2fRKyj/U2uO
+DWcx4/PCtyaXri72PCMefX5v//4IVkCijcq6tivoMXaQz1LAAZu+yrELPAbq2EW
rjRg63H2SFXphw1fgP6AOa2MhKcWch2N1cKgoU9XNuMmNljRbAkBnzzhq0ph4Ib8
ix1cbzaK0ZNQ0DlilgPZXyBsx09PMQqJBxgaweHYyFh38Muz8ejO9zrfMZBZZ5KZ
GNuI9w2yDnGcGP6Q5luyyvQRGVn1yqYL8KJUvKtcC/0ixA4mJQjOgX/jrxAykaCL
kYCVU16Vu4vKR2rAJOMv9E+xx7dYeKizfTBW+dxEz+OyW4WmiZHi//ePLid4EkWH
uWIyQM9vEFr5FAUjryp8UG5dHp0s+cLXX8DRtBhxmuRaDuw6gjkEhm9J35kPkA3j
BFWwvGVDE+TU3yj6h+z3AlXfNDjjBm2acVETking179h7sTLA2penUbL50e+JosM
plwaYQPMPb6oLL1FuTOw5D5/JRH+CneBgLnalX/rWm+22WmrWJzVXcKCDcBXtu8M
AKSbw5SOD15mOVahBtJNj3r7mHNjbYJEQ57tCwhYrMazWmV3F4qkb1SP/dNtClQy
PhT22mzYwbmWXa/dteVo+/Xz9VeXdWl4adpU0RjDj1bANtITNFWcY3U4jZEh/R9M
V6b535g/KbSCHUisr0Pc23cQoQ5DBdRKwsi4+zaTbGN1Nn0wCQXU2/RYUFV3NKBF
bV/y1eRMQpACJjDMuwD5tGayLwTk/fozjETdM3R14Nsf7U8rFccr35zIHl7jmtra
INun5yG8KBmCr1JNSx4+Pwk0lI/2W1sQub5VRqIxc6CTQeDZP2zJo0OWS26cIq8u
HoSLTX+MZiK4ZPJKWp/IifZ5gv36GoRLjC4aPsFXGl9qezhw0XVdGydHiO3NC0G1
ln+HS32rtsomAA4pus2zausprjKclYhzIQjG7yjrlscYYaeiP5mph1Q+qdgo7l6V
qFN7J93mJP7/uXyKtcXS+kmQKCQYNbyAZ3kQIwEu8cMrD2CTX24mONYeATvdMpIa
XA87p9C44zK934Kly8o5aP8ojAwqUV+NAMhMECmU0Bt2hkDy2IwU7QYlH9BikQB0
PwFvDOGIUC38OYvKZk4QShGQsMiqNvPehX5scwR3+mxAc6Bd0ialLJF8z8eefTZ/
cpzCuYtaWlQ3z4p4jktrxAtg/wpaLagYEBu2DfBHNNmK92TdVSxy4QJt0dsJRRUS
noyNqZw+WRrVPrXZrUaNKyLGk1cl65egqNOKXgvE1uKwMl+WygXvVffoDQ0xXurW
XdspGx/vrjaFoPFZ4ER8mn5SkVNP+zOzGQr8LjRkP/nsJpJxIDQ8OctwULOn/mit
i13tYUsxL2jtYegIqWL6GLuPgkSTLIXovUfc9QVoUZPLq1zoOpSYqfTAcb34fW/o
kNsLxYbq1ByHF0K/pv0afCceZFi3gA1LgLz+WLhlwH/+TaXH2q0aAjwaPtJGU51+
RMpUha8iRNvY2LB2W88KufNp36D6T7rS//uxzPdQMC9dIP4LPjiw1lVWxh9l/OBv
tHbJgV0MK9jXQqQsXDqcSiilpQRM8c6KFOyJC1tT9feNGqtRq2cISMjP4raenOub
Vh7mkv+KM4AdgmtWFUI9pITp20XB18p98e53xxlcRjT2uvWpvOjXSvnLutRZSHk9
1/OjfySkBWGpE470Lo+XjStIM1Eydxa622A4XNmccfxBitfAGJHdwnT3aCbui1x6
zri2CAenFDlll3snGt+bxbWKEkw2WX3XVh4hEWm+60s/6R9wLgYEt0vOEhmTlYpr
1kxRoxdI3rs/fm1dLn/BS8pkImeZA4gwH78qEjfA/Px1sBLX39qOhe3u+8Sa7kQx
YwKaQV9IDmhO2K0MOW0XLlJ198pefzy7HQZ7Ck02hmN/FkRnAcEXuKC+bVpelh/P
ZPAasTY6ojXiFGxp18sbIoWK6tqgTYPlivrhUtUmIdrALT0IW3WkTdryAIrvqQnD
lSBCcZ6S4enjB1+TOk138wPZrx6xQa99bOWNyU6vb0ZrRLUSmjyasE31123QeHF3
y1dsEulUZeFyPr5W1xkrFQWX0Ii0Cqj1QOyOx7xZG8xrG4ID0aTuyOXxkuj61OCL
IGqP1tycdvJ0YvGoX/3ps+Q9PHO/lvMtGZC9XIFwh/tjCuNzdcMqU7Jp19lwfrVD
HwfzEtdFk8FfY2zF5AhRsz9vRoNTM5ENlsx9gaVnvwwxiglhjMeoog7EyZg6+7MP
XC4R27HkOHqCbFvDzNysrEERp+4xnr8t1AkETNgcxfo7yR/vd2uJ/efLM8rIry5N
mxpcFnwMHKPLGaJsAIXJJuIV+TD6Y5A9NkKk+ORy0dCIQp7IQ4vxdmfn8DtN34oS
JPNikZUuClXa9oI8EH5B4AX9lH/IoyLAKrmqWqkYUUlO/S9h3aPL1DGkRpbFPOCT
mWBK0fqS9CoSSi2iIYUsZ8BxZ343UQIUXf0kJJafUHUnzXFcuc7C5MTP0CxDZwBB
/kw/2rioRD95Dkc2ThXVtXRorPw2d4Ncn7M0e5790iW9m5aEk2P0SVtSZJpwimz+
eIGEycz9Zd5pqtRivOpEXgl+eLNJqy/hgJ6MbW8NPkNxNLBxN3XKQiuZNfUD94RZ
Qei77pADNUsDV9ntzuUl3FBtrDJVsFqrCrWeQzGDstBWUWtKOC+V5sIjzDMaSy1g
FvquUAlYqVzSCOeZU72811RmLVfumuRrPDFlmcYdCZOtpqraGTQ2JLv/7jfIJu+E
cJnkcCofyq1j1iiVwLZ+nBL+8/P7nKvw0kg+iS1PMZHSLnknoq9H5GdKEKE5GEBu
zqERzivr1L/1JiwTDmFWNZVg2V4rqkbK8FMV57O81wsV2d0hZKfzn1KvvhquwgWm
C4oyoGccRJchxMxAHjHzZzMP5QbIYAq964KyU24yw8hHlVx3RSjZy3YMKiSH2Ewr
UHiEIhEQTQFgDwXsWY+n87uwepAK7/vLGC4/TxPtJ0WAF4LBTjF13eXsT2XH1phM
z6QHx2ASxJSJCmRSJRt5EifOiD/ag0+G/GhMnXriYPTQHW4jz51h5+HsGbA1tqjY
TJTgMLK8soQut4WDULbLMUI2+9Kw6R4OOOBCIWh5iDzxgMwyp3k0A1gMbbC5Oz3p
Y6JfbDjimT3D23oJjKszlmsY4RMgXpBn9e+FDYtdhP1VzJhkXegra5UX7RV1hZbL
/TCKzfayaZzj0JLFkd8mWF+CPS7DMcwkv7R2GoPqT/zT6mdzNoIxAj1TbarfkzOD
PiIHAVo0EMcGfzoZgTNS9mJ0h287YZnzosUFxzz4tOxmeOavE6EssGq6Stp/hRlv
DFDCBba11laq+q54WpOl0JSB68Bovd1j/0zDZO9ecNWglVB2sPN71IqtQ27Aa2iy
pM5UamKaUzZraSRsb5spuvAEhuw+D6nmKwigDrOFiHGPVAn3XC7zjaohA0FYT5z3
SC6JkIO55cejsit+VZHNY9b5xHdj8TIHnWImndm5qNsVelNUyLf4DzDeMh0xz3dp
Hhm8NwtpwCmBTl9Yf0i+TBmprCiB2Qr7rehVZPq4Zhcsu2RDIUhgKaXzEdeaiohF
wiZrjqP1xgGmodqf4VfyeU5vni11Hr35Dtsd6kT+8yBMvg7Ed0ElrLmxcBRmmnqs
eYSkvNUA8SQpyfS+ghJsartmvCu6a9rrwqM7hKjGvzhFlBorCKpTcAO13w/7FZVL
7z2R2/ZTofyU1qls7b/ghZmQ5dyE4eNVXPoADFuw2mGRGOiQAtPDt/OMiPS5/xWE
L4EbE++ADK7pV1nfgxsApi19LSazIgh5URBGnU3ESTh/U7HzKAcIjgg6rfQMbFxg
hnh0pNQmuUtn6dfpv6Ovm0Xjn0Xoq4wgd3uSG9zIe9hPRTpp0j0J9DZcjWdGgPCe
eUcrjY9NA8ZBPo39OJ+j7KWtdQBvHvow+7tLsmnGPew/WZmIM/MqcmSx4+hJKaMe
uQ0hQL9c+Z+nLqLYNLV5QEFNhzjl9HSCV0sjDxWdBddRo30ewltLv6IyP4GefD0J
uRM574FSFVaTZGlpiMYhcU4YVJHYKokUHX/YXzszP7CvUTXrlMq7sOEzgEc8u5ZR
uS66PsGNGskJGw8PGPje0EHUUROg2uFkaF5v1uX2NsRIrMGaSbFt/rPuUm1XNX00
VM1bnmEhW/HCeUmGmOtKBpJuXZvIvXuHoO9a6YtFM0/948H3Y3ZXqe1zCYiDTVJZ
aSM7g/Na/Hkl1tDxcSy9q306q0qpVt3ndjEKcIoZOERjtGbUV+YDWLu3M/sj+S6V
ui8vBdsuUxzCiob6l2ojUZK/kcHczv3e4N6q3tHa9on8zrVUHdePDt7R0jD0qla3
pOEP0hZ5cYCYQdNDxlO4X9VTjGRDJpaJVGJPEPFyr4UypD7W+MOBUrdfl7FDU+8B
WW01Q17NUprkL7l/t57rr9vS7+FIeSfmRjxmH972CLKmuWqtaqe7F6XSLToXQJbq
rtGynAPrmDsqqDwToHrkyF8aOoIojPi9lsBtpIv4sA9ry6MZQaG7PpkTM6xvq48X
5DIKfFT1LETbckyyUgEmofYQWNP6zwcHarsRyq857Iq40kUQQoSOAbvUmpK6Z8s8
O8V4yZ2Yjex9Iu1nf8Ns1Ya/gNIBVmVJ39OBE/yca+DKu8W+ovnaDBTkqJijg6zs
nxviMEQyrWHAOxhtPqWTMlXfD4/QPVQdTvCX0T7d1BbYGR4yctK99rVs/qL3szIh
LV+eqH1ooaxDyMXGZQ/lkykJTi7r2IsAeh+EjRJDaAkQ6L+v8S7uAPBg8ySvKSZr
M91vqtx99JgbSRSd0uGLqXIRDfvcwIw7hBxeicBhDjl28BT8Qt9yWrGdJQGpyIOF
gV6DhrJMVTBmPDuNwTv4RMSHRyE5xC0dGkdHb5gMpg/jxFReCf58BQTj90lDsiUJ
Obw1SsLpnHbKYRRjd7KUCW+2oZydqqiMrpUGJqGzZvJjpnEjgFJTRy1dV1wl+lxm
Vx77jtHZ9llLby8qe/lCizlP7IcJOOCVYkShnOF7ksrSSe230leYq8NB4FF7aVDX
jaZcm5Nf82ognjGIL+kAMnr2tKe5wXTUYfJfhF+E0ZztF0iWmn7xZ+l9dk6BSaEa
PtupUHopNoNHkJBJqZ1nax6Qh+qXasLK08LzgKwpXD1/UyfhrsN2OEeUmDVb/AYm
hyRfIz6B5X5XubHdX9CO4wdnMAPwRJ3+6bxPz5Mb1tv9GNpA+eY5hIfTYR+VTFLP
AnNV8Uetn+v4S6iH1IociMxKFK4nb1eITvE1YjpUrooXXKirruYR4v5C7eqViugy
LCoufnpXDWVGIhYwS/vv+7UBwsxbogDc9BXAVxzIRxXA4iLRq6hZVhUf03eADJHU
0mMFaKZEkEeo4Ym6p9TCFUffJocmJGkuoUIp1D7oN/2SlHI9Z4uS5pNNnBcQFrLa
qql6wL4D2EyfQlVPdVC/qC1JYn0xASmNqxGXSAVtFpJUcLXwVNqXqqnWZUNWqVXz
Xz9UU9+xdWx7utNqEPK0gx37lDscS+jxmbhSJgWNDYyHZT3JDUTzBQYa6p22DwzQ
32AuOvmxhy66sT9c2vC8+9iZB5dY8cu/yjfwkZzzbfythD8FjLa3YE/utKSjcmpw
wpxgov7PbXggJ+oinrBRPCTwUI4WW6p3cg4Ry7JzSySUxbUIPNjYq3eZLKPNzKPi
eyZRqnz+oC+cf7Ml7ftmPaZAdWT6/u0PMGSpzf/BvHgvXcY5wXiXBrxLglK7KOTQ
xx5kYo7+P6J1MQK0iyCttsNRLHaaBWpPQRBMm+LB2hLlEf4k2sk6LrRH6Ux8/zA9
PscfZvvBEmoSOF417FwkM6N+IIIUBUp9j4pLs+Uhi/pcoRBZAv8j6JOxds+XmVIK
enqQ+ZPe3/cTs3T81DsM4K9yMDtR0ZYKTt2pRMSQDiETfsFJO6zb6TNySLojMD2n
hvPRvP54eIgR7qquTQaqY61y+SxvqSbjNZ3ps5NKmn+6h5rR/O7QIVDzg/y1bUXV
OIjClt9yvLR6ojZkWZQM60SPNJppvPDSCLdKIcss5RpBaxciVxLd8WnyL49471lM
Ju1qPCRrLQSZzMeHVKJbUpGfyUSmSt5W7ZYKh1YZQz8M9RDQZPsd89MQPUYzLlVI
qtXRb9T4CUxhHa6F30WGW6weGq6vkR0ptMzjjp3AqVDOyFOlDUrVmrdsKUKqdTg2
7iZoKhM98WprI3XaISQtLDbbCCZN85/dhLW7I22FZ2zCu4dJfmOh1NlgqID7bN1d
TT8r7jMOOMQnIYnA32+tiMnAbUNuM4/e4kgHFbIl1oVAsv5fh58HP99lsZhDeySj
xM7q718nvWKN+rjI3ewt13AlOsUUfVqzTK+bdWg/xTjtthkyMfhDoIdosZRBYnxy
t76hFR7LTC5PPJjiT9KdAvbPp4L33NGzvXlsi3kTz34kbEeBJPsWlFqgwQlUKeUL
pFqrgIOFxNqgxfKze29/VFyJSuicuo66/Lq+VTpbL2hvQ4np9D+Y2dVLq1Jc6V3O
xIPtVY8d8DFGpvgTtFVr99yAmblJFAXkjleHY0PhNdm3ZubYMhfFtWaA6Zme4Qjs
TadVb5Vwv4e/gEydkjKGh6ciEHb7Hlc23bHKM6QUQaTJnkj+avoftTn1UXh3mFsv
yFCmE3eft7XNFouwmiB+D03VZrdLnPdft0W9YkpZXJ9ZOWQS59XruHh1ijXcV4NP
Z91RQjLtCkY9JyoXJVAJqcquuv5PenrJquRxNPeYzGXNK9N5FmdlqlqVm5bAQGFS
Zpg41b2nzDfiE1F256mABLIxOY+VSfXxXHAzdZXoO0ylsC4WjY36vVzKG3lVOxnQ
MXf7epa+6Qc8EKcI2FBjjH6GQUfWMGeLl5YHc6TDfElC4ZjBguBgH6qMIvx6nySF
z4Pp009GN3TMw/jwnY0dUs9oEQrfCiFkxux8FVWhJDd2eG5awHQGrdMGrc4JuiNE
MZ3PEdHlCbwoo03nraW+q25B9qV+6aQttmfxncVsr7GinfRcLKbZQ3aKFx4PW9IC
NCAe9r5SzbEUy5192wwnxnZXkRg1PUpRX+Lx0Rtg2i5CqqfK574vZFKBRhzDtkX/
daKdsfNEjNssbEAa7VF8hWPKUt/nOmN0wRAFmG21sClsMwXtGWNPTcRwec4KGz76
BsWv52A9Bpi0rCkpzqfRjc2QRSRYzdhKwR8W9sg9Osxvipmn5YPnL4uG8ClO1P5W
IQErpUpEaBCQ8NkUPgDCLQSZ5sB2rfvPCREPToCfsZZheCdVp0EgvKpXgXCN6LI5
CoglrsThGmXW4pLDeqV6i8WdyxG2zW2wNN/EDVsWh80qLXS3Qmt6Vj4PDmdRqejc
Mt1F6fVoFR/hIvCVZehmfID5lryuSLUVJfOJavUJ24WSyUQoa4jjpg2nPaMtW1vi
fAgZKnvcxuN9VMgAQw9NDjlF5F/2rm8Mn8dzo7XqT0+3AChhub0nekvn6nVEb+oh
gS6XzPK/Rv5iTPnhtneRfU/kNaOBTXrWvG8XGBFj3bpnW5SAW4uP2MFljUza1ol7
p8ZvKv1151IogNUY7YaMu1+Vj2i51tzoVjDBT4Rdm3r97J5mYjjc62xcJRSQuNPx
y+CngBMxwxnt+k1JOGoUBVd8sqKU5jqXkb4ft+q1T2aYaNzvxZPlbpnZHdWngdQ/
cuK2V+ov6dNIeo4DGm/1vLNVto7JcE4MdfhuxdoeTYfGACsLSExrnfsX1TMQOGJt
M9HB4vgrlSF5tRQbo6taHdVbeg1WiC+KhHfNygRtU5gIbPvMadCFlcySawkRXVOc
mp4im3BaJXL+lqc6s1ilwScET2WimHJ8c7Pu9/wDWEVY+qeaLI2u+RTQrTaezwnG
rXwpaqIAMbYRAR2LBz7Kq30r+ahXlcbl3qvTZqJklFrQ1ajvcRz5ww8KeamJnKAg
iz1/lO7bi4FdVNfB1Y+Y8bVY8zhRDw+d3jGBv4F65Sk1FzrYtHVHDMCjN1iU5v/9
GyO19gyeWuRcBI84EWEtGJFXL8JTkavOg7pD8q7q0eu4wmL7KmMwKbXdtFBXmebC
dLDuOmaPNeFizKlwMhwPULZoifyCIQIgm/UKMbxCBfm3HaWQXkI8XpMrDhBTcL8Z
8eLJt9YyZQbMA0sFzb+p+dj36n0KY5TlOk4tEOwIBLRk89ApCKrYOSAzbjiLEr+z
5EsJ6jd/qGLHjD8UTd3LlphTVS6S9nM31jQ6QcgDa8nd7yD7JTUahN2p+E6c3Q8H
t7St0SfdpMRA6Pn7CnzBPCu52/xFHFznHv1uEykNPp5MCiEtVE2DqpVLvwKe8fhe
g/lokwg/klsdD8qY3mjFO2dvHDeur0QVoGbomL4bBTkS715wyhnDqjKb74YJLZyx
nXHCF6isvAD28RNYXW7zKTby+ClUA5glas9de2VZBi019nsZk9VfntzBtCWg0cPd
H10UhUe5Cmm6ycVkMSRdbzXQ6W0EE9fovG76rsNLoq6J5lH7WGksMIDeg4htM3P5
R7WNZPmjSUZdApt14gr+zj8SslXajYb7AM3sjmXXptY06NBbxWxhPYFLhR+kmsPf
a+ZMf4+nLZmxItuIzQkLC3YFRtYoN9ZioDVWodbStQlx2D+vcuZgKbJ8G5FAsaL2
N0ktQdtzibKEjJ8RJxxAPQAXk+z9g6YqUxTCE5zDEoGz1FOkGsFOeqeGahLE1xL9
PG+jr3f+GVMaFWS1geR5OVn1WOdPLN4w8hl4F7EBWc7DFqXojEd1WDyQg/eMQHw1
1KfTRWZEvz1rsrbaHO2+52I3D6mkrWCgsNgkTkY+RdC3K0fAsQkcSsG/N5zjw1Vk
XK+jMEyE1+1kqQv200HCYhRiOEs61bMrwc27YT9NwcCJ1AxE5eXLerG6t/S0R+94
nHlu5BzDCkWGpmISJz8jrun6pEqdYEDlkHK8UPnTpFWdAsYpoARxR9lx6Q5lLQLa
8ZjlqhuEEZg3JlwSYejWPZhORC3OBvJnIe7uV0x0a915g0o7p15jQvc9uUTAVpz/
XH6CwNRLYiUzzo1i8ye533tcvY4saqYzWyyo0Aejmt17wgtyQPDrrCmsFIO+wYvX
9tcOc6KQRN7Qm8YLl1gCqLzvpAK5z9BMg3u7eB8MdVzECcBR0YiYLy6eKrgXelBf
ipZ3gBd7q2rMXa3PNSojreJJhtPMijhNEshXdbnaAmimsK741sEwFRl4kcn7fzbu
ZDsxFItv8RK63LTiI8MFXBVF7vkHIQWqrOu/kVggu1HOxFOrEMtMwSx6z2eblb4T
BKXngzQoqjkY0vfyDmmBQHzLuUcoAthWPFXZxBvGADy7VVnyJ2W/b8a9iETkcIBg
O/udSVsgcphbvzjV6IyffKPEibHqhqp4kyH+L04kBTNvhmZqvj4modJCi6vxO1dx
ASjg3YNtmQ2TAzH3Z/fuCS1ztC24iC26BSAHrvl5umZO1+AAEkLogEd2d3j6RNSq
xnXRaSjAWgqqVEWVMIHNwvOtJGt+32gXc9phc/o3Ea+pxoki530JzCo5my6sPPjs
NPnEOk6CX4890LaGbYZNkACZZ/vqodRLyGQI3Z12IULi+JNm6dC4Jy+2qxqqHJr/
VJRj8DyzgwuBqqcHr+X8Ga6xD/nSlH61qrjPf2U5iUqIRgcQIcnIpytIGjuf48Yd
6QpamnsQmkR2vrZYUk+G7K+M+fMnh2a2Y5gQqyVzd7dh8fXuqR/F+23F87DdeAZ2
aQe49wDco8Kaz4dc3mCre3hHYzc3YjtvqhIF+N7EHfTcCGcdNqPL4fK+SDafZi8m
CNoJLLo7xyxy4Z4+n30glwS/Y3ftW55OvypNG8juWC0HmzWd69mTY+GncOik1hza
WyfMvsC16EGnTlhVaaTNmTYikEwRdTajIE51OrPwRd8htzg7hROHUjXBRJSX3HT8
w1gETN43kYUBKCYo5ox7UYOQ6DGYwK4IhqEKQnvn5KgK7yWHCZYhRORh4lJ75fmG
zwm5RqWk1zG+s0It8jNa0PD0oYkTPONDU5oAVNnS/8fykl4K4dbeBh4Hk0cmdegk
HdrCZB9ayGFD7VFsV+6IBwHIf/k2xgTJPcLPB5GHPJ3S0NYlYSpsQMrs3vggCnbJ
AkpHzX243mcV3J76N9JSkG3imVA3ECFXTKXa/obY6lgjRz1Sb6ZY0+yeCsTsUBJB
HcGfqXY4bZ5NOCRyK9JUOFYUdKTiIq+yaGhezGiKmMPz+Hj7wNGj+xJYR27gwQEx
hANlecZcTES1PtF9Pe1EeFx0EPpMnGlHsdMhmuFBantMgz19KLUCU8H3EDDvJdc9
DMr35R0jl2r/70xKZbKF/0f8+81fAk5UYWdd1kcILohNXc6lTAlW0qYt66AxYxQz
hVJDzYXPE7HhgwRGOu9dUQeliSwI7/XP40Ale4h8ZFyVeV1lzjPL3m3ki7Ykufev
vlVJuE5tQZuAjHnUlSh/pJ+YZi+FPEyPUgOr0dlSvK7C65yOg1ibNjyYvpL5cK6B
WDcPqAk7yiayQuSGDPsVnV+W2K0fRY2PDRnssqgxHsY/BwP5xseZCyxaqq+lsXXW
QqlxltaVFPjpjVip0vDNES95qN80q3lBspSIoJwUojB8GjLuLfLOMcdiJsF04JVh
pAOLrCatjWp/bJP21YeJ25+14KBvHvYQJIVIMJh6rEn//wOeOREeK2XZjTCgAHXP
h19jWeHgULaSUjGeA+Rp6J+4+1XYqFvC+54CB1KQVewBKnECfb/6ipStFaPTpwAm
cf9IDascGP2goz3kfFGQ/wHO6iGMB7BLdIJYrnQK42j0CgINQWFDje69zaHfqylh
ySmNgQgNRXCBr3JK64RLnCQDCPyteXLkEXGbJK5KRJ/yif0z0XeIvygITSD89mup
xPOPI1NKxfaTd0T220exogRzjbwOBVmcWziDrjLWjONQH+kJjv1JjgHwjG4E+aeY
FDnd47HC1W+XjbFNMTeRDzqSg6repruRznIJCoMximqCbRv0qojqhJLnSIJqzcSr
iidYg/xvCNc8rLBv0+8PQl/NWZB9p1KzWYG6xtHRndKnGI48GYVrDtNV9ln1bXh1
pK/yVoaqHrOfYo7XINeArzJLw2Hzn0UWHbSfsBaw1DEW8NT66bbi+PsX1P3QxuT9
RJsz0RbUKsu8rdSqu24/UMi/0pbQMQr9EkCrRwN6Nc0fzzEaKL/y/GQkKBPyywSe
D6q74c0RYibpLM1CBYdx/ej1snVZqTcblha9TPfvfO1FpDMBV2b7l4x3XMYIi+JR
O+0aq6Y9wwrSpQ91o0N7imNN06WrB9Po4FzzQStKfnqeYYkgztD9ugDB89Xcaffp
St/DGStQUpL2ZrV78bnPDB8pc9QpuZHQ4+EhGA6UA/VHEaUkzEfgPy5I9xoEPD/y
k6udEhed2NUAyUovl8qJ/B9SCXiy9n4JF+WnH5cuvTv6wKTflst3YASr86qqffxz
Z7+xuG3w+JWUwcl5iRlD0i/fHJQ2yC0n+1erJJX/mbbwKXSg8QMBOYiLr2zAs+rz
JTCW9ktEvMZLQh3d+La2HZ3m0qwJMGYoT5EfZsiKT5ZVHClXVWYu3vRm9WoFaQjN
JgZnnFngqPD3hEXlRjdBFZV8/RZb2rru5VcBC8E//5CTC81teaChEQRR3qeZNTgW
VTRNW+6aG2o4xEYxNJD5rzLB6OCnUN5mLu54H/ZzhKV4hUXCI9MVSM2x9uAVfWYv
dnGpXMEzck395EPC+ULB2ao1SVBmUtw5PwI0vdJK/J+ryCYUpz405/ZMpX0VBuNs
0HU6wAchtZ/bM5XifQ+rhNzrmpBl2knz+Uep4syR84rdrUqGjLh2N7GrBw+Upobk
zJXLrUJDJPNLPrKgOsqwJP6GaZNoOW5vQvKAJtfdL++8i29WznZPHuZXt2rbeVog
FFtZ+eOFBuLBM1m0mNJf0vuaRvSt/nTg1aZitSnB9XJxPQVBrP0d+Rkwz+SXcF+k
4XK93qj+zJYZko06LOp2v7Z/vTuQQkZvV/DQcHl+YToz01PpedwjjmypZILUmENI
m8LhusJ0rlhmfaA3xaQMgPMGIuOuAddXhx+waVMZkDsVdsDr0r6RQTBw5FytUPBM
1WLZbRsdG8E91vnED+jp+jCRjp93XP3FdINYue/2UsvUgvgMhQWGnFnFXxL2ZQoK
l2ibdVxiv7rPUlrs4sQgKBY9f+/cIZ7JdNywjzcdUttCq8Teh2Ryk3XfTe+brqSs
jPec1yvqozVGqeSuUarLmzuKf76yjBzl55xejHDaXNu15tNtXVsfIkQ4fsRoLFm7
Go2JemwlSChNu5a8Ia0T6bUFJIPtDDHeWB8lLJmWS57Vi+p8MP7yLvwmpb4sr2Ku
8rmM4Jlk4zmBtGrlEx6nhIfaPg7O2VGT7QCf8ohux+N3hVVZA+rsUr3EMvPODzL1
QQIvomddgCeQxfQpnfLhDvw41eIOKm7QDK67ImfUdFl7rC2c5IPIJQvgkHU6Cc/8
Onn8ftwoUB1SzglmrFXn7Qogm7UyWu2zWB4J0zU8P/IxwD//4oL02suIrclPaULZ
XO+AHEcVqvEZDMFmPSmeXT5x1PfmoNruO/kCvvmsn8bIHvj0/DbwruryUbQY/ttK
SnnfxOc/QzwP0pfFhr2tU2Du2bbDlDbSmx9pneR7QEAISrAF+Np6idLeAyd1zuOw
a26felOnMUPg+F59gYclaQGa2/5ta2BuJ2AGOukFoXLAb/MZKWsGFeS630SwthNk
avSWyH62ltBFvWVVuHG/H8wJ8w2/oOTCIXnm45QGBJu7dAXqKTyoqMLObZosiZvN
3+fe64zEmchxDzGg/IVMWi4pApb1T/hgDzMSL1ZlJRow7HWvBgGcmSKwpqKmOTej
Fp9BYn23GlGUhH/gqcD+PfBVa2a5N3MOxzjlaeuu3kNi0x1NWDhz5AYiGdIY2OJu
/3PGAkF9b1LBR567owkbWk0jvnJva0UrnmTmcSDZ/O39UGz+RyCphQsVrqoMy0a0
awowzLTY54NKB4/gEZDQ6wF3kuV9BHmcKZ+TIDRas0d7/cIRBQJ6IEj/38P8noYk
Jh195u1xaZRCj9J8PEaRuLA+PbWtlefCJQ6skDsbrLIvg0DsefGcVrWesqLpAJHC
ud2Y8Mld3/H335c5K3gcbTrdoX8QGj+2XKVpB31qygEhJemmvm4xINtUafcz5dWo
CMJfM2KgJCC4rONRUAKKHZcKEtb/Zc0VwkGigHzw3fG7iWgAK3SFVQeqSba/WXuv
m2LyZr0qU8mYxqz+uIN6qRclqnr9Jd4bi5Xryd1JmYvDnRgKO6AUaRGxE3F4hhUq
KyVAj+AbUYONYRTWPF3FyzyNPgsnOtbf+7zbJodeWMpZQQGfMIAAFiolHFEsIq1P
/bdJJXdEZgW9eu0csC+krHhTKSBCITBBvNEdjYwuwK/ng3eDGY3O52EIlqcKwmNT
mZ+7boREqcb57hOoH/F/Gy4dSgROB3QgFS8JYRNs9FYZlxP27pULe5YoydYq7cat
2YwZGF95gXYtvv883ngFh89XGrNzbnFrw8dSmNy6bkrl73svF8fcWF89jcXWMFlL
+ToSOKxn9srZ0GgZvlASrymHtAsgESOR//m7xI8bK+gamb665b6QESJ//Sow4vW7
YoOdihdtM52Q8FX4A2KjHOmXRezt2x1LayCZ29NP+n696uf34Hz2kNR69fudnWTi
ekyYJtvwEsFsy4Jn+J9OEfPccaued0QJuGO63P2AVogBbKoj28MWXQrV6YgkPwHx
dFU8ZOyjkS50ktJB81sNgycMwO5apWsXkS1mRy7E7ngL2NPulA+U9Qrakg1w1SNb
eHMDoj+wpmUXlQHzxEFBVnGd+gPa2fx2SUYA20YcyqNOiweFuASnV2HFIrwHnjRY
xseSfHB+v1zlwdGK4INOjfB99cjfjDSackXRTMwGzxsly3RvR/MoZ3Ob/jUo6mmH
fBRxsRzGlIAiHMjIPwS9YyNAykSq3bp5ctvuMflLZeymj5BnFrg+irYnLP4iTe9g
D6wYzH52fdEIVbeg/3JFCFG9tkiImTOarfZDZhChKYk1d1Sn8IcV6ZgX42r8RlOq
Qw0TVbSBcsTkVnQtmx7CO07QvBLXYHDQLbKY06lXkOrIDHDefHejjQu1jjmzvcVM
DiMKDLFZGPOu4wYmuNGy1xXCsJmS7goKrWC7qf/Hz66zcXTpszwrtUzy/8MHKINa
YFtZ3d8Zth6gXVXsXRVotHifaAXBf19V2Cbmqm+d8RgMUewm/k74Mc/3KffhTrBj
2Tl6dlXqYbcgToc0lSvdfOnYyrbnCiv04lADvGbvBR1WU21yf3lcEtN0kl0vSExA
HmXVmTkQ4v5U4fn6QGCdrm/5ELndcWtHed6/kWJ0PyBFDDlaJwoTC531Fxf2SyJh
tcDalV8a1pmxEmAnD1sZXrzCe9kEHBn250heGylcQ2kYMTDSmemF7R4w3Jtyf565
MsS+SZtJ+KiVEKqbuM0PUxzatdI36dq72vM0NMmz+IpK9+hursuIeu83i6aMtnrR
ljPVZpTMqAPCeTDv+F8yeS7B03AVv4aBUoCeaQVEiSHWdoApkNhdkDDV77uDgXiQ
g8vqbOu6u2xHlEP/lFnVcLaBDIqKNIus076AAuXWIpj7VlgZpgqrTa1aLHHsmCqY
PbY8LPfzSJYw7uBWdLtQtI9u1+JssQ51N6OqCy6IizU+pnI0Pg9wQvicYTvK6lEy
IXoiOZLoPdGTTUfthiyj2jRR4CioHHeOCOuBgHepucaIiwI3Lx73LeIkyDx2DOZ9
nBKCmUgsZRESievUhdlmfvOV7/If0zqBjMs0T7YUx+5ANNwL8MoaIuPdQZZK+s3b
iDw5L3Qr1aPynh+XBlcYnUS5C2fRsv6TXFqWVRRy+APVNiRBF1DA7WsMOcNaArNl
1j/jA7D6wJlDrvDJahHXRPKBXWN/vUIwLqyrKT27ds6GnQu8cVxKGgLZ97H5Ooh6
fQNXKOhUoggv93TvIRrjfbOCbuwpW/1T85Ej4ukWlP9Iy+MnXNSRQpei9u+9JJve
7oOjYuj9mcjw+qrDEUgUdHadL3cdue4Wkm/UzbQC8LPgppbqulXBhXiNplQHO8GV
nadZAiQ8svex4O4NlF3610pC1xgU5Pr8tzr/FvOuVbCmD6+uc60UPzD+IyjskKj+
8ldGITshiYiK/VaPko2YqVlblOZvzJwQTPRHgK6WxX/l2tZbwHnJKnTvTXwwmhP3
TZf0gyF3+RdIyV9PvA6xqM+woIm4VjHQnU1TKcWfAkSlqC+aQHcjQ9BgGf4YD/YC
ltf80bxgZMfgsCWCOZeBv1BRUVuOb9qV+Gpudda5nmlwIOZ1T0VvXerjU+NLaHl8
+RPJmVIDePyddVB0AoGKHRh1XBIo4wb6bMZ/RpQ3zBEMyx0SQKs1oaJi2J90d7XA
3TIDFcBjzeojNba5QGVHLfkDTnEO+/ck/4yhO7hynp5aF3LYMFjmzkNT+rg6NjJd
JfYdbzilaREtPLIlzs4oeKFrtd8dxTqJNJkSWhCZkbJ8TT2qoBYHK0Fm3jneik1W
1QsJ2ahHPbP03Aq9z5rOAwoHvAg9Ge3dOnkonTClG69boqzWJgWTW0/IIpQTLPA1
ywG/puLa0OXjNAhUGtzT/ptp35gUIDwEFgwXHWcscoiINX4UO9xu10Y17Dv0n8cC
xq06W96MyEB/GoPBS8yqW6cSL/KISClHZr5KrGCSWVIj8u/7Aup4t6TAfJBKXRL+
CYx7m1Ct4DKgxIx1HLOFVKa3rYF3N/xEdvyIVN+ydSEVKzkfM28feurvg1K5XmF/
Ql6k8pcUGCMPv/uwbuhYNGKg14bxIaWDtzc87/pvYlnNNNctnFi/O/RXkfS3AUl3
T2ASGrs0FfNoUni3Gm6May99N7OaKk07laNZozCI4KH+gfopP/RbOkMoTpszzFVc
twcDTT43hLTtz0krPl/HTQd7hfidg336J/m6+rs/OYX2oXLjxDubMJJroIKlC2w8
6uvvCHI/EhxHfA4cHHTF9PC3t/UrjXqbCrK2CjVRiOzjQGAzreijKd4/j+wVuGp8
uSgNp4sC1R7dIqg1Zth5A6tzf0G1ALjfGjGVotg4Jrh1C+/zVyYL5WeBkFA7NRL7
JXIgGmxUxDouRQ7vhOFUAitrAEq7OR1xUY6rUqhgosR/pWDMMiBqJ/vW2IfNN7BG
Bs+pg0F02RwkYlpybA/uJ8XLp/rjsdrAbB+Fr8Ks5nYvV+Y4wlZx9uqzXB+btISo
gGaytju5m3P3hHHd3XB1KGsV8lyAtm6BhQbiKR3hRTK5Mfv6VPxs2EjDO0d05y10
B4hvY/gMmxuY/9uxQgKAWtHJd92Xw5ayLnyREsB2qtcoqQ1XxkzwUkHaqt1XA2fx
TyoISpHEDVkEyFa1EPd+fKWpHweG0ov+znTiedy372zUciV2x52z8bn+b9VuKHNa
V7x/JhN1bRfjZd12kMz9xWJD3Vk+uD9kS3rP9LAnlON2aVHU4FAWKnEHx6ISja3P
mTVwOzWGKf5VWy2Js6Aa7SUijAUQ8/xGlpgx/7UzzH0yE5PjNRs47AkQgz/pEa6Z
YDI8Z7Nxsos91OgRU1NgRdNicyMY9BzbvLgbm6a4SIa8ZhEhFxir6QLUTEqzGuOV
smmAHBR+BN27sdIE19+ze3/VBr4wy9FDCYcolc97FCbIO0IIjU7a9mH6sGMJ8kqK
I+9bDWeg5Xn2qPYGZnbT7pYahKi2M/LImmWfzpKo0QKcXxh3bXzS8sygFtUXY/WR
nVFhg2XXxPAtzwasdL4ycBsIkjcnZBWdQQsWirUUmn85zGWgd4y1H+yCF7/yWRIT
+ZoazXTMhbrmlPFkWjurhfDAkOTzYcGypIXiaN2Lz6eVaATp+EHw9e5bKcfA3eY5
qaoOr2oTJ8Rt/XSg+dCG75T3odDh7tU7Lgu+/BK5J1w72odusMEs6McrszqnBPiB
hVk6qiN0Qaz2KRPQ4CtnfDbqY4qp223EsaPH6MckfWoJtagO2y5yAtxCC6E6omUI
j5QfaqsOKTbeSGbLnFsz2tnujEiLdprtH4PBizrOGQbeD3eJp9lxetpzTLQHvM2I
lXMPZIod1OHbsukd+d9S0sAaGUEtsqsLoVS7kHTLE2787XFzDLkANsRKyAsa8Qc5
oDO5e3ZkxqDnyGiRVBS0u78zm+AAj1581GGhU9x8t1lmpfIBIGTkzPLc33OLvPk7
Y1jdHsD9mgCSAvbSoNov2WuwmllFVBjDdbcIab5zhGU6+awD0/sN1dVwcX647mV3
MdDAZT5zqporoKWLOvXBmPjPv7t5kV98w+K86QypkQc80wHQtJjRxbDJL6fV3Cgy
BBkeaXDkamOIS2IqXnGiiWzM1jgOa726hzjRV95IVnoPh9kWRvJG7v3FeugRU436
phrxq6J0W66oVfjJmhid0RO2tSEA7sk7+yqbryBieq03bUlRVnZYp4cEmQY/sR7p
KY/i7BGGGGWzCTeiMQgp4CYOeXbjwQVGYZ9sxKgeEX0qQ8sePz2v7j4mEAgYVh/E
DTvXpDtfv1zNWNvc+cItsbtFeQV5owTwdKC92a4ky8emLM5QlgRW3KPdt6qNDXiC
vRMw+ZkdDfp4wz/J9APstdsBMRDRld+5rDlO5h5E5PhePeTT1zXd+sZkZxyA3szd
BtPhqZloqqjMXtX8f1Yq4MYBDRlJBgX4vP51i7QaNysBYktB3xTab7Caou/yJ0/S
RUQCv/jwP/9JYSXX9voMOHWDBi7jEbPdsrVn+yMaN2PQBw0lsbrfyhQJicC7HaEz
8qtxAf9WQ74qJ2BRt0EPtsb4V+sm0C97QQM9ePqSp3lYAwEXwneIbGZ20+z5kKeA
I1huL+GWoX5GmO2UdWwft3Qifan+CdWDBomA9cqZaZQnQPw3U81437s68Vh7caJz
zZbL4NHH9763ySI1QgHtDzzAvIYJpcyia5ydTmFT9eUBwQft4XHwwDopyHJhLSju
hMXD/x7fUBV8+SpWyD1hp0XtZ1gphwU2i6AG/2sAwBvwGoNEVC1BKT6hmwKPCDEy
xhq2ol+flBbryogTtheTjrsyv+nPXoCEEAYZlfcIe0aS0a6p5QH2crGVJjJR6mZb
l3GNR/2g9b7uBZyaamwiRgGCFpUTjwCLUNftOG6p0tJBymBNHzmNVPFfGbcMSxtz
sn6cud3KB6EaTRPi6c+iiUcenGib+DUBq3vQlHLmDWAepXE6frmcjvo4tyqrpLKC
tJDqAN9DYT7ORmdl99BG+X8swDZrQLxo6mohYXi67lOnM0Ee+XtEnyNAxGzuR7Jt
dWLb1wwL429RWFtJDuxUlASSvTR6cseXNCUNyGutUQE8k3COo3XjbS8OPlZU1BHT
np000SvbKycP4kY/awuFbbKTf0jHQ19bgBp394NJ/WLTYJ+hcpDr5mRWgd4U2mjE
JqZ903/JaSJIx4L52LMbplbnKfK75WOghFUTUaJWXc7NcIYHu6MldJR9mbX5fRdh
bUffYwviQ+vPWOGS4uaMMbi/ucsbQvhUcO9E4lYIRJYyjRCl87ahU1cb3vPmbuga
kUI27a6dEYH2xlkPly6BRReAByplcbo58Bju0NRq4YyOGfxSqa0/GQ5g/pJM0TY3
ZaRjtiFJDxoW4G/zXrPykua2P5R0sJdnNT4zOKh2sXo1txQ8YpNnmWoZfAyeiT1r
WfEjx02ckEoSViWiwVLpJm4T4Gxor+o4NKR1kA2YFsioYgUFUCwzQOk6QIAOsSll
THOf0Y09FVeqHXG/yHqNdTSIlz30Q69P0fECIne7JIQAW0jMYV5bK0IIBvoe+wYT
5IiIVmFAW6f2mF7v7KXthCIQWky99PAlqWt8hf70JSUpTf0tDQx5ZmRmVSzsxCci
51ws2bChEu6jDuoedJaXOA4ogc1UrdYDshAH4Zb8HmYTCUVXoDa2GvF5PWDAncZa
qEzQ67fyQAP83B3+PTUpISKXqmQ3HDGAAhExsMimiINS6AChd/9LFBvXUm41x57S
VbYNhgc7+MXanAA2RuYCbmkUl3VW4wxxTiIUZHKDb+x/+yjk/DX5qUxi2ox32lpx
lvIDrmPALPBAm7MLwCMu7Y3c1e3bK4P1Okm0dHedxgH9tbf/hRXVuSUdgoIuwWfK
pel0Q6HPH0aRstcAiEfCNxM6DSKVubiJ7t3xsqhM4pme7crvChtz6hLIRj1hmsyQ
UcteyQwA1NlI69fKPmwHfjEdKY8NuvydlMaH5q/1khe32A1+rg5sgeS1cKzqsxSE
1JFZATBUmzxnZnixG4XLtToTirDtUL9eyM7HcMP+JuNP0S1GOpScXyXPgmXtrGQJ
+TuQWhW1aHKAnQHc6g9jq4GVFLofe7bs0Syo4tsTwXhW41wdHLrgfmLgAlQ91cdp
CKb3pogDjuQK2Y9AMQW1objL2ZfKPULJXk/TQXbq/uSNkE5CM3dwZg5YwogGFNCb
qSvblwgsgGyKec1NNHDcFoM1Kbe0SUWgqhdhAWCUM9Y5oC3vS9UbsWuo9Dtp3Nsi
fxljLx1nzBWnVdvj1Lnrqmr3cebnm13vPgqmTXr2qoveCRQL0dhtMiP2EEZ/S9St
suOjs+1d0TzyeYLUsr3TK9i3D00lf4eZ1pTqVpFEItgRKCWKBZF1oS9Za2gQILil
AZCxIr13x8l8kF3j0CU78KHJOll8EP9gAB4j5EMGGJhhxxzkKAvk5lBlYLTFO3hx
aTyct8MYlTrW/0sExRT7EBVlXbyVCgDYifIU7ftX2rpUatBkgluaR2BzWnC/41qc
cmz8hjzASsga/G0WFaVApYhd18yFSREwS8BErYOBTNQu7bQejNt/KaenrN8vVURL
dTvb8I+86CR8MBeASNwtzxcd75plgTlzK6P6i8El6HXDNTgtHiDEJYkg5uAnxNoZ
r/ZIeFceAfyE2FwP3fN0TYEC8S7l452Jq3UwGPbDNZFsqWbAWHa8ZN8+mtCoQ1hK
w6YxMsGUhOtExIuTuPoPkz5vXCn1bcXnv2nnH5wKO1z6Z6JXitXvV9re8EzJVwUG
y8V5jThYri12qkBKc2Q6zIfVg2qLg2UJNGQHULltG3CFdSQNvpiEMZfQhXFLceQA
giGrqElBpA65/4oMwcX0iOxpt8yEkRTTNKm5MuKMs+Xhm+G9dWKeW/QigAJcNvva
9qm3wku8CBTG5Joovq6iIGV7O4UWYvHEeNsaZ836+IUTlh3UlPHNma7L3YDCohAD
+HCBEyMkVUbLDZcix7RCT9CWoTFmCEOLRxufsBcF45G/jcNB3VOBFUsxV0GIOMpr
XzqahtWrv38+V67ThuUTuNMjJjVAwZPAIaVXm1Y48SRirJv+AxAWjVo4QKUB3zFK
/ltBYxepOCVwN1l26o/pyBibYL/IXkoEjfU0N8E8OzqnA5ITS/Vx1qq/BvKr3UGS
PYDeAmvzVjoyQzGY+SIiggoGLKZSfiR975+0obmBZxTYhj82JRPjcm1Rqlnlafry
ebqnMzavOW9hU6M8Sg2AVAEVaX0JR0DrUE77wHHE1u+PmA4Xdoyr0UEnPXfvL67o
/MZBnQUn+y6ePU3e2u5aUIxJRbHIK88ywElij31aXkjvWcwZKcvRRlZA2/E3M+LM
vhxHPQdCiitRliWayhEQSukB9a1kFsX/ozSL25lG861oC+aOKmG961lyaFoAWrXU
DdkHTMEtnIBy2xUVFAVNKtYgjnhjQCqzvyXaDXjnsmPmZZt8rc80RKBJeifQA941
nxQG74Fn4XiE9gAiNP8oYSuTma81lITV4HAbyrKseYYauQp+nPYVfLshmp5y5bxk
FcApBtFKG+tQfpD2Ezeur/4S0laXqEFIckeKwoIHFj7ajAyzzh00jT3dapjxQFNZ
T7TEDeiBIZMxDye4cdreftjLqS/bA1hX0hMz7F6AOKJUXSDCllBJFgP1I/bO2igS
Yzm09T+huWLQzf+k3klFOVHruN8lfV1vaQIh6Iq/UPu/158K8c4kohaWooE3oE/c
3e006Fyp/IDEE/hh5lYoAPnETLjss0SZqTioJ8TMtEt2VctLwp13d72TwCOB1nBG
MzLgMR9vfAXs/pBI5aL6RghFQ/FJba+Vy1//InhWVm8z+IgOCssScLaTBg2Mz0OD
ik9vfk79n2Bd0Mgy68bDTjK2RJiRWnwJypmv9+aDDl0IBg8tXM0BrHrEWuU8LL+f
7QGvjusOKeXX59dkL+GAaV0WB4QBuuylJijBnAikDoEXPg8Q8pdVQuZT47W2ltZc
RVGyJZVGj+JlrxA+hDpwItgrWGKSDoxKaCXEuZFUQiVJa5uc1j84KvXiBOtYiEUC
uz9vwyZaSaGL3a5ywCuUgi4+OXTRKtz1EVdZFYCwQ6cg7DRANYMPPNXrhMdjCJhE
BH5oqtQ+aLbW6E/Xn0pe74XnJmtBOl5VamaxC0yxJdEnGA9U6iNPPo4G/0enE9X3
Dak0US12hTpSHEmiL4btLCUcH/gNd5jQQ3QJ24AaZJ5Flb6d3aR9ROh/cjVTOj0Q
fi88qQfgxT8dD7lRkNaW243N061nC3U5nej8WlIB7qEQh3XXgXATr5FlXhJMdqCw
ijWra+Vw0pXxE7PATJGxEuT7/QiNIZbhfUzNuTEYKoyJ+hIgCjJS9fgqxhl+ZKtM
mtVLBZdlRtDfptYxKA1lAIhKkrZWd9DWO77Jmpt8tV8i8zg3jVDaK89yojn/CVaj
8Ks3NkFrDNSUpW503bx5BNti1MUijTISHVaREJ0vFWR20w7GG9b528a9GYZPbxz4
I2qplLMO0gjfEOWwDDMjT5tVwneKrJxqOV450GkVwscO9iybZ676iat9jYZ7dgUL
JXzUbJ68ALY4aW4UMSVAJnugbW92HcU1AO/B7RCjgNvmUUc/75EkTnV/pXnByOBR
B2JXB7tVTlkTgLp0TIo9H9bxyNiNF2KFEo+ZZtNsIqYUQb8HUspKNKHAZJda85lh
/6ZrGI+18GEWSxi99Ju9NTZ50knpz9AYnedDz/1g5Y3SO1vjbcVho8sITXBjQ9xc
8DTRSGLqj+MhX3WXRLu8bxNKsKQFiIPoxKzFUkJBlSaioBgTUlKEjnJUaEk8vTc4
C0oVgkOHiEAA5eVrOHM5rbpbp1KUMCNF1h9ajIOP61qjJ7ljf9VmJqRGpWeYu8x1
x7DwDNludI6iv2Ej+sa/K0/8Amuy2OXRZf82kBsl/Iwx2q5dspbijBv6zR1nwapf
WcH5jG6hmg4yhJWi3W9oBzyns0t2MO7y2hnmMzfiJGGKBkqPQaHzo4MwLnNlLv2d
N80GUlF8YWbBbiLbRfFXLHfmhk5Qxmj+Tz+8ACRAij7datsXGK/i3slDTcUdqwTP
ee8DyZ7P7tIIMVIJWrdQBgWkVBw8rDdZ3kV0pf6gUpgNf/2REcJklb/P49433NGQ
B8RE3k0G6tO+iaIsPP5mNoYVYu5YEPCpBiyOJ3g1N7KeWnJwBr2gdIWwqUixpBUe
5f2w9gmg5dGJVP05bhi0/uOb03ibURrziSV2lwWBrEYtTbGKCzopIWMOrmM1htX3
/1VkH3LIoA9xw6bJcUCGyb9TT4A31JxyNLo+ljRJU6xCpM1EjkD7erbQuqSBZmvn
t71hS6Td6kfjlYOamPTzz+Ajv/lmWqZCN+mJlobSvkmcusvb42r1/xZL09Cwx4oH
8sDU+X2a9HOUdOQr2bv9KpfElcT1TL638gv76LpJqPq4fqQLML4QhnsbWVL9Qf7g
msKij+5+9+o2nArhSxUfbO+SOUaA1AWmRq7h+UKuywyFbhljv7jSBXJ9MoI7fnyF
syySe5HXdCrL7Vt73hTJ/KTGKHSTKkynQ/MUhVIUfcKe/mCUzU4JVOcLzo3NYKO/
ArsU7FhSSXOElyNEMUPQSyKCTamI472SRkEkBgSoyE16Rtu9zre7Ht64X49CSJHb
xgTKcVxW4XOR15b0PNYVSZF68NTrkLPWpJJas/j4tMqRsfgfW3IeS1/wcqGcaDDV
DLU2n+bDyAwgkZmwGjiZSiOfDjSwBzHHEbunkw/HKnpEX9ZXx4nudtKb7aWLXnWk
4+fNkXVxe12+CoIVjkdrl2YqJEg8bPCPSCXkNav1B8Xzn1y8TOGK/jm/dpxUjzVH
0h+SIVSQWCZ3nzfBcI0Eg+Sw6PA3+bQdpT48I66KgqbDDgAWk11FO/JRfx4+d2pq
T6wmnnFcFRYvJFg+JePHee9Ot16BZx2gVRqhKeFKhzMEjgyMO5u2QmJPZCYvsIo6
17uQZS+uRY32ktnZYJ4q+3cisNQap8jz3bTBd1y/qI2EOTHK6b5bgC+Y/aRE7rZG
3ufSGmcm08feb1rdEfztiNAe7svD7u3P7ABMjvw2rObYdsoBbz53Xp+1LBnYNFXx
iiAQsepuzAFB6EbCragAtzm9j2PFr1c/DdQvnRu9x0ekr0Z5Og7OCpIu7aCrlMLS
RO+UKlzE8wJqeVSWeBXB1YQ3vqWniPjC1r+Qm1TabgUBj6ODQ6LuVGnHgafH2XTJ
w4OCghjJnQFdBdizqq0hN53pM+/GC/HjV6CZS7Y8xvfSRgH5uIKSH4pdy0QxKZ51
1oNptyex0P2FyquRfHQ3aenwcVTgtriwsajn28rUJSmJST1kIfZ3qTymq/QjBog7
Nrce6o6otjJPfeSgV4IebS87rblu/GzoOprQv1Z1t2qmJLqrktfRmKgyCfAOPJ8U
r1y8Vs2ySqZ7gj52Z3OvUysIz6H5QQlKEI1KFJlXUmVXMUsn6ydDGVeqvnxS44fA
iW09m1yfqloPzXEZ2qqEKVKiNNG3tfJ1as/FdTdHGlkPb6FPkEH2AjA6nctejpAm
wEluUdLt4yXeTO815cAqYUvBqPfJuIkRCo3DvUfb08XXHQEJ9QeO3HJk4KxaROM+
I6yzNkquzUy7/b4I7Rue5U6sGLi/Buvqn2F/0SH0IARdWhmAIP2QstwfEZkOVsZK
nrxIVzA4FrKbXlyfkV/pzzkorQ1XyD8kBOPynZbo9WTIG4VRVXnEffqYF9zD8D6O
/YWvptrAJ3M1IlPyk8zJ39YZzIv9LOHzEqm0mY/YGIcddKsHb/5PgR0yksKUbBnw
51nXPFRIrQyrrCau9EtCffAEd9tNrb2O6v2agpr9UbVNPNY5negU4N/4KR0sosJn
fEpAYzJBwn5JOqRcnpYLiBI4iaGhA1e/j4F6G5VAPDOQFh3tWJ+iQR+8o9/sIDgT
zpdauuy3mAJyCxlXQUUbSJdw9kDR5KwOe98o94HNQL75QOHbOJVRawyRTAPbg5hL
iRlzpNxTL5iQ92kk3RyP0uu5PAWxGQaFZ3rsgS9rzu0wwgZPPmi3FJHJaeD62U4/
aQwk8HPGDL7zb9T6bN7N5s3KJwklCrcv0zZguU+Nj2doU2FHOGKi9Z8PhwvkMS1f
/rQ34lOI68uRW+GjuXrfhfLtzTaAd0v3aks4VT0lX5f0kkWOhK7MQ2XDshiu0Wo0
/jx/fFHtBsCzaSd0/L1ywJ0eLvnEkfvWJT2KRUdnpGeeQSp3KRcyNSM4+3tqrtQZ
1Q+xeXGkgq9PcCzUU1RfcXUx7mDimQSA0aPcC7nQwOstuMBBMhUVUzZ0I5Fg2Byp
PQHyDkABG0FUCPZB4NT7/HvUJ45uTUs/k1gadNt6wxmXp+Y7ukLc5VDMzpmvxZi9
b2LDcrFdI9gncH+jFDq9053S/11BTWff3aaxJJCD+6ZGplNXil3WvgB00ynwrsbw
Trh4UC85CHcsycTsIvBTNS/pQHqDLH98OfxThAcPwnZeIhcbv6Ri0u5Ch9AQ65Gc
MhKofskRoTQm138bKzWbbsI7Fad84OTKtgoY+cNZ/vcYxSQqftIiW5qkjD/HWT5x
pKWqQg5EkXChjBzAgdNOZF81GOZeIUJCVqEOM2uIE6qYcIQtsZ4LufWV00k3gDWn
VWaetar4kGXDSQX7sxMnntuXj5BxEJ1SmoM5PwATWHWcrZAXvuXEYulfyyfp9m/F
Ufk5R57ym2S6/lDJIp+4cWCVOOUqoUmlzgwmQ/FoBxIP1j7KYtsvCQRuqHybyJ4e
B9N5GC0FY8o2vn1RF6wmPaLTxBW+gpc8FuKCK+QwFgwInAEv6Wj2FxJwHOKiv+Li
smqu4uwuAxdpAXqV7TtrUco7hbDUlhBv2SVXsnPljBdMzBVnbwzTJ69cySyj2BNE
h8kzFfCKb5OIjN3MuPgSj/iWLP6bATyNbENbzwCEkhpDHj0Btcp+kFpvUaGoD+yj
Z3g8Lk3qfRjPCKZdI3cDhw2PrFzS7Q4kccycnCAV0Uz2NS3GhdB1DIE15B9aL0dd
0VzCv5ej07/mo7x9gg0FMpg7xJ/Z8VOw/8cXxfDM4Ri/uOHsLXSlX7pfoB/DTnIV
0uvu2BKTDI4f1EBdpmb+dO8lvfbrc0226hUVtpgQ6A1mN/Iycn+BP4Hr3GLkZdrt
UOHCopqp4RYVv7ViSU0Kqn2OaIxvobnyBYy6Qb/5JHSTI0DP1FoyUIJS7nOfnMAZ
ynvyIukyY1UGCpnp38WKuXLGoysqDOCVgdbOS/bX4f7OTgUJNRRhvKsqMPXS2Kgg
77t8XRKPJ6Op3kQtdAWCfT+kyrlQuFGZ5XhqFPQGJxB2Zz9yWuLIMo50O2yuU/bx
u9+qr0e49zjzVe1EsTKGcDqHmJE2QxSsU71RHneJtEV43V1Ry9c4SPbca8hcbaPX
UO4jLR0MBHC4UBp+ifOG3i3ZxHxHyP/kaYNyTlXKzFhzvnGCrqEaQC7H/SF5vm4l
ko0dFEJlcqn4ZL6YTY1kvRxUqMail88iWmbr1AOjYPMWTIXJLRu4QVaFXJoHpSJA
JJfxzI+HNaDzuwlcZUk0iCFlOnRjuEJwr8ioOrx6NAcNAXBZBsZVLunpcYtuG0CL
64STU3SP3Ajsib8A89IxYnJB5hKExs/i5ySkMhnV8y99OMRUzbhT1rwHGPnHymFu
MtMFn0Cmpvxl7X2sBGEmNP2uJqKWMZM2dMm1cuMAUqxVdEdP1UTB9yAJzNzVPos8
QtND0YFjizcOotoqX2FxiJf+er4qOAVJrmlIJnY3wmsnurskDmgAfE29NH1smObQ
0h5W9k7cXSAGh/g3G/XubxhuYmYvZMy0H5xwnX9T18ZYoEWVBGp5zJKJAJ8BB/x0
2GBOiQKESK/MV6znR+rJHR4wKHcEaZZ3d2rmnuTO4mPj+8TCefAji6ozIFYhEB42
Z0XIj85aBbj/2O3CBTa8YS3TeN0TIDiuzJ3FNdI8HaCm9+ie633fDdlqPJjSUeR2
e3wdUVk6muiwUrd0QxSKtHW0FV4XNAjA6WjuAeddjW8/iAaZhsZC9Nz4Az+CjXPp
I+ogNLzD5UcmSsUFh8ESw4Bk0Bsjh5Dsd1EyQCO9VRvQbL/tHfaZbeMxI2B7ymMA
H5nc/6425clFCJQ8wQAjeqQ/DXrbewaunKOYa5CLvTQkyQ4XdMY/WgfG+s6CYMfT
D080eEX+zpIRJdHRNvdDG85Gllf77iiD0J+he/LVf6wuI0rsd0GGOgEcoA48i6Ey
GUzPOhd8SaID6dny/GpJl+eWJT5J9pU4UTbIn7SRlLQsPWJGysETPwbYzsI8RvE6
MFZd2+Y9me7j9SiHF9VpnqyiUtQc5G2BWnMcQoAFN1Rb7WmCxzcYDV7C5jGb6h8Z
Z0BQxftr1QiBWeSWbSqNeFFpNtJvr+ihnbD5ce/7coJzqqjdQ5NNzDusjDNODEIx
96Om/imJUbrBA7J6t+Hr2E1ohhbRhcJy42qqG7lz1Uo7wsrD14uu6yRUO/scuKLL
ckREQTlAz2mP5hJRPiSj1yrKjT4YmYiR7WQOQ40pNca8wol+W5jQB3IHt+qsqP4W
AlU4Zi5YqBEp3X3QbVI7h5vmruTdJUTAAZsz6mwAkex2D7xWkVxvQj+TAAJBa4hE
AsxK9mnFt6v0T7ebYtt8YUQXqOo/iHyMVyjHZc7Xr0E997xB5dhUux2xQUAagXaL
kpn+aqyKMRrq4TNvxJRl/qHyqvFsd5jJAJSEjZR2ch62HJxlz33MeorAEgPIQ7dr
Gg8eA3QhUkcjipH+M90g8ELWjCPQu8N6U4B++aLVy7VT4CIfBdGQd9uSuMEivF+e
SW8SE+p/nXpNjzr3euKD2cLiGawM3C+so3qgNkMX5xbc5Ngy7Zcovu8jxAdzKvev
YTn7w7pyWQjVnbqv+QrJZCEKUH0NwLFFVLIr8vR8aaguGJ5UXNb3hxhTZzKQ5CoN
FwSOSPmJnJWNh+A5OB/TnjxSjQTFsfcrb5wwrdHGbp7+fAojCsM9TGTLpEFFSC6W
Z3ETjr8PLP6Ur8D2FLjegxPu/zpQ5H33g2Q6LPWmsbud0xVDFCAe8C4uNcDoRzg4
lHDE1lQKWEzpI1qdTEHnMCiMBtE0Km9TjhZQc4mwOBjyUKlRUSAaLQmUanbrsqYw
CGTfBXpzETK6zAKpgZkrfB41fq0nxwSSU76ArBGmcHt9E4yFb4Vv2kw2nlSLDrob
PB82EgSis9rRYDaGLN8lZrhmtjaDCsylnCsnetfCRfWXPHvsmsZr+LsQX8ew7dsX
q8/fdYkEkiTNhJyFT2QvOJl8dyY4L0Z0gJw3SgaTzmeSt8vz4LPL1cYEb+XQWvVb
inODWfyygFif2t4AxazvPYV4qIC2/gzhNKmt1tQfcmBiVMDfTucSUmSZmczjdrHx
Xj32U3XXwnnHcj016SPvLK6kHoPhw0EfM7hxuN/I3hf28LxSAIUeEF5YAR1WR3z7
YiUnONRTCJDCYreKoWne5bQKJbTKurL249kFvbY3yU+1hiz2gjgo9FXus1yKaxVQ
kscu8SdNw8cQUKJlmIvvneDrqhPAqMBhup8v9WIn+SjhYKdbI8tvJ0GhwUCuXNXs
FRiF0Ti6gUybpJeDJc1KNnu3R05r28gXmSgN/0tkkf2WjNTFUfEdoV2CxnAOCnq8
XMJ/0bhY8ofHsX/rk+e25g6LmLL4e3yF+KzDrR1h5jT+JZBUHaDKSjlxiYjWIaTD
L5slZA2WtPp4AxN0bxkDQSm5xlSCTL8Ai0no5NRf86ak8mgkcfjQlZLDWtGkNpCD
sVe/+YWZSPor7iQp3Whsar9yL/RbM9wotza9y4F2vj+83fVTBtUb1WVYNSzecHp8
Nj/fBMvKknS1Nadh29JuYoLcA7e1gSfq75mHmr9TAEDxehSj8rP3tPDmgrmg1+mr
D7LZ/P05U8qpEfXZl8nQ2njsGzIz1aj3BHRAdJUFneH5CvRVo3fvlvL/osTw7hsj
cXS0s08SOGc0dCy7fZs5VtPATdhlxIT6NCTHkVsAobH2snAPUecVTSEUAfDNEDuZ
44NeLa2gAWcYkrvxyP9qGRhxMJ3gPEBDMSoLEEqOOPqnJBcz5EedfQ6Go2lQksZA
fIHJxGQagHrHYbNLY4BPLLHcLETl/1wMe67OpAVCPAkssXlMsLVsBqZX7DW4Bd2w
WZ7qCrmPcJkEERfjrK1I0+tg3pZ1cCzaK3/rES6+1lSL3EhXQGJ7VNaYmQWlDQTw
E+UM/Ze3HMdU+kOqPMxIK/3qN9D64SuXJ3CCRBeej1E7j2+/io1F3hc0/IO80lCg
RXmwC7qUrmacS4D3iBTXzC+EzD56Wa3l4+bZrK2Bi5fs9AclnSN9VSUqmuADmGA8
vkEN7V4PKrs+iGWiSS0PycG+6Yg+cEmIq9sQ3oqihuSluqRXK1gKO5cntPyZ2gtr
NiKhR+OfUQ+Npyjq7kbh5rR+uLnM+8aiCg4+m1X3NKiqyDkQaa7JZrRGfK2/Rni+
YGYbS2q1OhiPOb20NNBtEGLg85BUAuxb/ZGWWMenkdRgT5stum9hGS5AslwST+Tb
xrcAEatv67PfJzCWjyGuXIps2ed0wleUrn2u6sO6fnGiOge3bWG3zZ89iC69MUEs
A4MGS+67odFYig8urNV+iUIQt2xK1cvfbdvJIKpPwe5/YlUC28TCxjVrlaslxAtT
v5TLUfZqyV5/8Jr0UxUL+0KF/TiLrGNcVaCHahDAocu/G5YG2xqC8M/WDdx+dR5N
l9XsWJdC3jrkVIxugzb/hJmaAdas42njq9pBmOM3csZz4oi7PxNU0FxbFQaZ1kLF
BhUydZ6edBNspnncQRu0gSCnJWnXso1wF/phWddXDt/APOpfGuZOx+FsdEhlb+fV
VufeZrFWE2oH55rE2bBxt2aiNVywYfsidES9hLHtObx7ltOJu0uAUv8POT+ihK9x
x6eDWdnzcIXQOYMUR+M2siAE7rYUprLKD6atyP9+G6YaFQRuVcojik7hkV5aJc8w
JAD1EHKV8RV5H9ki1nxaDRJ2BJeNxf4Yr08iwMZSOcgwi33GuIxZsmkiJAwM7x3D
kqHKT9f04+JCNn4psV18XqLBH4UHIOQJQocim6lm9Etvtg/PjesF7d7JOyJktgrQ
3n2gqRm/RJlPM0IU8S9IRTEgrim9+n/ysC2ljJgjWrjRZ/EikdSNZ0ZPIeZcRtSX
j2ekZmOQ4qKZMfcLt499y6i0F5tjDMVHMjmv1ZVzNx5r9iI54Pxte5iIfaYmLILD
v3datuhdGL2Lb25JJ7fdAG9hHGIXuDw1ZUwQniz4HlZl/Bxa6OUFbHJLyMTbgvkQ
zkiJlAjIqeRiEvBOHhgJZ0wAWKNuCzpPHdY2f47y5lAGFTQUnQAw309aWqYFrDAR
Kd7qpfABzsxkk9YTVIUGpjGRrzBjZnDVQ9/T4Xluyo8YMrP4ZVYKDBvcTMqdIvIL
XLUuQtyTD0HaTr9PUqwVgSTqktCFEmHbJ7+4oUGDJGJaSdp3PIzoKKhJIu10Z7He
W9UqM8pKj31Venr3XrRM+I0r/Ir05B3aTg0ZCzTa0mZmsUyawfsEhMPYorqyqb4r
W1A+oA2cy39PxVLYCMAqxqarWFpjSXwpKRuK05AGnTnW3XOp41f+jK+6ZsPBK14q
DwYJn1kFodsUJLcKmzI0CNRPUVCvjHDmiUcYVsP2HNcHYJlF9cIRy6J/RwhCqLPX
wMmbsocReuSS6vV8ZvTW0L6p8ikDAsDh9f5j1lMUrji2v90LeGeqqMmu09ed4Z9l
ZEKOiN/5tw8IDHamvyZgP/xyJXiUc0ozZwB4Fw42xhiRG1QtutaP9aTpIzpaNb30
U/w0NkNDu9NS4C/9/cbllmFRXj6gdTAi9QGJ9OjzYm7/tTsDB7sFuxa+YPoeZYO5
PxP4jE1eVjNDP8DN569R2TVg5ymoSQ0PqLh/Sv9Fno9QivMEfNS2w1h4rpXIlYRu
yMxKnDzPKQT+Ht3UZQQqbhttuA/i/+y1AMtpwl/5JWAgz/UvDXqUhqm43OUARTwl
IMA25TWtGDQV956u3Bui/+RYi0yxVIwJEep6o+B/KCP0AESkAhkGnuqyu0ENWKYQ
W1lAb7UFbiBoaVlv7+UUqaTI6i5DmXMhQnOiKHDG8ORGyDqDfWHsU42Y99dj+0lO
Y/70NXYyIuThmiVUPcS99ZfWznwk1WDkGvmhfF1tNH+q+4Esw1k7BpSyFAea6O6S
tWwMZ0jWwIYrowo/gYNDm32L+IeOrVGJu6fAFpPcRUshzImKgYr73g5xRpZD4NTg
LyNgvvG3yrhU5xbUth7pnd4cHfO/k7Nm6i7VMJCGZrq9CObws0xXwrlDggIIB4ei
nUIX/CMb8fR4b0BqtKgI0magsh9iXi1ECSR2oUx5B7LWNHzgoLXzI9JW6jSxpz7J
2hy/kaetBbKibZnPTfUc74/JDjSL6DLhQMzDWaIK3RmEdyxCd8fwUgH+VuHjz/MI
lYvyihcJTKm+jOhM8pFsgXaZhWoIcd+IzgdAPcwN93ysDoXqHLx0dkvdCvHKLbqj
zLWLX9+U0CrDPtWdoJgKJ0bDkoZDwKnHlQR8XLB9/GirGP+ydrLD3kz7xvvcYPAC
x85vwU34lyQsBHcITr47OTANsHcguY/xYnlGUC5eQ95SUx/ogAgI7Gg2Z/XCN3mz
VMN4KhK64SamjQcdi846tKKBhMsG1v3zuON1E4D6dIqfs1f9DCfDQg41kqScamic
wZYnLxwhYavcxbCIUofvc8BdXmEm1DpBo08swkNr+B/mgWtwXmgFaS0jC1rbbWPc
LXslL2YkB1jEIE/Ao3n8g4eupYTaDkQoAg00xZGMWUGsSQQ3TGBEBYZdiWDVu2QP
0f5/luX8wuTRxuvpcXgzZVbnD9RESVuuhNqoQN0HM28Lc+ZZ5fWTuJL8q7pPbKn2
pETTWObMchphdqaa0dTCtPBVFz/NysGEWiiHBzh2HN0EhOg4qzacuongiH5Wl5SI
AEpwcJffQkPTEc2IkdDaKDYAOD+DUGwUGrWUfUVULm+48ywBAh/LmmCl0U5L2kHE
ZoUMuU03rqvgT7UoRaeJLLx+Mh3tao5OyUQZeKhJSBuh6ndkXjY1CZbuM7LZV+DE
C6ZVM9rToF0A8CYDCTRlALiDYpcwedNhQYepO2xgTHe9fEbWdKK6AeLlH55QRldo
GTvqAI2dJwK3fCphxGvNtIC78DrsnCnyJjiLqujK3C8Oe3ye0wpMYSPciyGdzNVX
AIUXbEYoFzUKNtit5oiL5H1xLjc0+98QUJKcatLefAfHTNJokjSMsWkGk56jpK9V
VBIc/oGnMqYyq7U77n3Q8jmgqENTplD4qRxAAPVJbT7XN8Pj+z28BDNLYar00i8v
Zir0P7u5ooAI4mkzRao9qLoTbC2WXqrEI2yBGQfyLQXzOw7v/Yu+WjI8sLUWbVc+
I0f/40BFagLKjg8DA/pxtMY/y/8TAMOqUoaZsmsziAEOHYA7cHoLKMeRBC0F8k/I
LszIG+ALjS8Xv3GBsqJ4vJxDjYT5lk/hg0G21Y8JW2hPS0S5Sm4FHDgRweXmvWj8
ln5Kvv9kgxb8uHz+cH0J2nzgrQA9GuzJ/afQKEazZ3VB3TpijhuqidAgqz6ltabz
Rr7is3Jzhca+fgAfpMfOFaxwNI/5LErJHa7OJs4m0QHyYV0jL6cDrfbXPa868J3E
YoyLrO9v/T22X0MGLkAjluzEScefJbV/u6NuV7VHHQsYvUFD8X7Eo9GDcRcwyYNy
Jkav20MUqC8R+CDl6FXir5zbeWHG7FTJ9MnI8hdpMY36GeoIDBzmeXB5MIkRg0V6
LPk0wPhiXpGlrk54G0HW67zQLNd8rMQZ5ddoKvqd59B6VoBDjdD/TQ9Ishf7RTui
npvLBnUICVmnz8T5Fd59XvMGvqzjJFiLY7EBjQnHP0ipv10AT7ytpon59vu0tpac
loQj6edIw3faU1lVNjOEx20zFTCvQrBdMRd1NTSCXKopKiUDMHyz0Lbxbso4A/z3
Vc+pguTBWqbBAXE+JJtcSrCpbIrc2UQwoOGaM+3ZZiYO/LhcHYlT7L2FrY1Dt4aU
f/pt4QdcM4jhbhq9rm9vbGtlLWIw6tIz8y62pVF6zBOj2Z0gbjkNqDSsDU8hbDGI
4o8H7zGCU2p22AB2d9+RViZjqft88nF/0JmJCMyHe9wrEizpGXcaVWUJpuja1g5t
Are8b0zG5kE6D38lBB8nJaNur8xYuNyh3BBhNnq/86eBm9BkQPZvx63+KPJLB3O7
4wuXgs8UCLv7avEx3IKR7B1KG2Z9nxtOtMTWgwznBy7QcywAenCATGWAib6Vicy8
pjjnErIumLvxE/MZzY6dj1YZ6EOMJcnrAn0CGkP1/lHt6luWEDMvkqZqQ4g7KkBq
APbiSu0hhB1O6z1S4vqlQY7Ehgp+Y6gaDkzFdzEU5sBxq+aGD9gD9uj9AcvyC2gH
hCKftUNn40pLWgFpkJxN5H5qTzE2sPNWQQpY/l+Qvh1+AU4V/dpnqXY7xOBRgM9E
ejUtIAELmfwBwyq9fhp2wcQP9cJ4VYTVrdxEENkL222yt42qDwr4uKu3qsrsQWWn
0zYBj8xtlzCGYZ1XqaadhPnaCvGOxNtePvZzt6HH+N52QsgO0LRaaubWMTg3Rwx3
yobA5cZl30+lEoEyTaw0XAbpAwnX7L0V4UtPpX4BiYENOv8BV1iLqJ0ynCxDiDR/
ZsnQzJiJ/1y73bmIkOyIwk2Kx74YgmQS9QMu8tyUnRYaZ12XVWlpPRzvEQpuWGEo
zjNr4kHLqhIf0ChfwB31g1yASalD3D8RmMCBO3QVFAFe2SBpXyUKen74rgu92i5v
DJ/rp1WUETRD0sJjKG+57gNQQriOqEpe3aj7FfaleH/PYXI0B1vTB9ps+guqBLXf
4kFIYniWeMdOksmItw/Saxi1uvzRceISyOuaUOJigztqjnWQG29jXpAjvRS5A071
n4De0AVVwNUW7f5yjxYdPIIuujbiwocYmpei+vgUZ757+0LvCuXz/KPJX8tGb2Ul
ZSHaimhAECtvALwPLSb+m4DKQmTE3BQPj1geYgzvFyBIEX+oy3CqjTeDhCx+gnK/
H+uKtLqSUSrBTaHZ5yjpyLe+JZTZx8zXI0gU2IzTpsehgdxeSWa8BTY97aNXrUye
5Boe92AYHRSxvU3i2mbAUuX2JFlCxq9g7FyaMk/Xs+nI3V7tgxw42UWvzc326JzV
xz07ANQC10yYvpZUOzLegj6vZzHSonUAaAw9Nr8PGtt72vSa2MWN4z0aoIC6T63f
gGTgqZA0crag30tm7JAqaAK9pOelyjKyiGLroUMxmzAu80+cX9dwXRtBOJRGgyI8
1enBxZvp4oKptxoVhCaiMeo2H7IcnZ7XMQFH9JDAEqa4fZexmJKnyGds82zXDFMi
RkhCLw+II8ME/1nVCmk+xX7lMIBg4uhfPSDMhKxMMds2PpXoTpEBT0eazwr+iSse
hl8JkE5ardEhIQcv2/5w6nhqpVoOEXp4t67ivcnqVPsnR7ZgBw5553E0At5eLTkZ
6S8tksqo3VUPm3dXWeE7El30VkxZcZfA4qi4ld6WG2GP+XuYvanKLoxvrfG7Ctm1
KQya3py9ZgcB7baT5AGga5flUublw0131ECgkH8QaFuDtN7O/lU2lIB319nQaGZx
+M2n62WpwLtM9SPOp+vRFbc7hnU1Akvsw661nvjYJBVq1QNtlLj4Gwub/fiEBFWX
/97hWlJYGrhiCIM2gUrjyisV0dTRIsfHGm7+Xb60APZR2oIBgeDzBEc06jLzMatc
Ly4FOuvi5jtxlzAzdb/W83PdD/Bt9qTS52GfRxF/Q0bqBlEy/zJLzFQAx2v32GCZ
eoXPyJPz6T9BwpW6s1XF2oWcujeqL8LvIQd0VEwvXzJNp5B/iB3V+zn8f8FLUvwB
hnnQw+Og7lrxbKdH1Qr4JzGRjNI1A2uODWOIkBXu1KGVbyr/vn05nSkWn/sf9uIO
lKfJURWt12bpI/ZCXILXzv1MuxqGdFU8Z9+17uBBxbqktNVY1Fr0M/WfKRf9wTyw
UtGdU+DrujMAIb/GTacynx04Uboan/QbBCxB0S63biNWGJBN2GRcrem3ZjIijz58
6RfbuousGkgVZTLTvycEBeYJJMme8VPp7Xp4nPAkGgMOlhF7obJuMNnwE0QBiZWI
ZJf2Hgf6fLDKntQWz2EZfCNdQEhWpZL5lhxNrj8A0ZBfl0vUYrGj1s3lGxW2tph3
I+VpN9QhLIuQ925YI5/TvcMPN5AMUEFXpR/MbtFZJnKtIaZFJs9pHw5o5atsTqIK
a5k4dHqMcbeNg7g9Qne3Q/8Fj7gl7CPnJjyRtUgnejPuaK+lo8r1YkKdVty8gesw
KGQgn/9m/6gj5AcIu0VqpUWTh4iHyJ0jYk0uErjvK1nnEEpe9gA8dd9uKB2RcXLQ
8nBRTicp7h8Mtyb+5y/+5de1iMSOSxLDkmhMiBwP4zdSi//PoUtKnhFC5SRM+kp2
7yCf69buWbX+cLt//hOaE3PC33MXMjOSBGqUwovwnmZQm26mRgHOhqLGoMVB682C
7ORSX7QtZ/+yMOjjABMKdO5F5+D6Moofc5czOmYP8qaFebmvKjTRl2LuK87PflYZ
lzGdyOr31HcgHDT+ohCMRTO8bIpoZbSMrhXR9WucYg2tfSi7KNSW+JlqQRvz43Q0
NeYNV75Fv9MP1O/oNAls3+8NBB2aorIb6wiqIhEe8LxZxTQIBBbvjUaZvHGOsshi
sbp3Yv/cdumRxx4Xoe005ArJifeFgIBhwbQVqmFmXPKPIKxMcamW7NpZi+fXeiFI
r0JqiZBXncHgcsylJqk75jAgXZE7Jj7/tiNCB4+SUK0nEYW+HOs/yB0cJXIGIiaj
wY6jLzKEBHtte2I7FEsEZbYWYOolBL6IEh32mGxBZKJzjaElXclFZKJiiYIktsAm
2aT5RS570U4hPvA6nBCLQRA9utzIZYrptZu/LzzZx9wtQPYQHJAL0fv9f2bxK60e
yTVM48JCGawbzW9kiRWxReGCqyr0Hwr6pof+EnGyozGtv6XWsrFfSqyluYVMbBG8
AgnkQUJsKRd5EJhn5g9CCeURTA+w8Bjp26juMbkdY1O3zf2vEqVKUWnYUE9yKXa0
NTvyxbnEeTxlCB89mj66BEVAJwmeRQhnptCpUSv86pgvJIpNpsvaStMPEysgENBZ
kiqS/3XiPXNN13ulw9s2kpskvgSLMnfrhTkcW7I1qtUTHwli4SLTBTMn/13Fx8lP
EmUxihisxv+fqlJYO5yCmfLkeKLkyu8/3SL5NbJEv8geKnSvjMn7kPYC4ooofSIV
h2jQC7S9ALV9+KhoPRQtZDja8l4d5EyfvFwoAW6PBr1DSE8Jy9RpLpjkQLqbuJkm
/4tJLkD70bIjn7csTozXN1EPENWkXsr/lwMBb+WfR3bVKe4p92IojKTRlc0cepIf
c3OAIBci/J/BEfIbzdbzKsTO+Ia2b1liQ/1Y3s29ABsGHezujSFky5nMLRMBY2QY
tMoWwcVythOjDzCSPRRR9LIezIH7npsLIdeilDUvEq1HTrndOn6rveo9MZCnXBre
dx/C/hXbie1sTEj9M9h2OKy4cYwasTY62EUwzNjtNYuGTJJIP5aU4oMpHIFsVSzD
Gfs7E+w5jCeruJ8Dc4Ns/ECWbHqNZOlgc3LzUbpOwywHm0MMiA1CoLauLQX/pvm6
x0LdJa9Wih3CUkbLKUtC1NWbEPPai4tYkH2Ht3C+Id8ZS5mo/soZ9Bvl/wB+IVRC
2zNpCkrUDgo4qbDY3K/xIds/IlL0qGrYheOh1JZwRCrbGeSJmt2EBmd2+OrEWo2W
+4t/Ild6QI4l7+h8rtXP5+9db9wj6nzUCy1OQFr9yDBgGprJXjMTyP8nXMBqNT68
4vUk2dQv/1B0poUM/Jx9ed2WaGO7mMwb7yBNHE6tJ1+R4IMXyLqiOcKHc7FLm688
z0obeFI2jYdqmWbyB6YmeEDr6y030zVmI3Ig15VEVgsd7UXd5q86CXGaq+gAz+tn
OJZg3Hs/lkHRB0UqjFT9+Y9AUFusn+EWbePWaDlcVSrxvDvZ/Qmf4tRTJu/+shda
TdfiCLO5VTFyAYBmPScHgf83U4j9gHEnr0l4vVq9xyqf8zqkxNKxs8zdFZXIipo2
0i0o5AgYo28GhnRt3ZdSSW8WUMqJcgAT0qjyjdcPawe8LyG4daALTMI0Cjc5qSZN
9ooIbKEIdOtG+8jhpPEMq92Ujhc6cddJlJUfPf5agWBDitUwXoZOqXKQcy9Y+1DT
9E1ps7lfVoNeq+A6cioqyoFHxplBBiGYjZnxG+paaAKr5J1q7gmbSvJdtDfOgDhr
c4AZuFfmcoNz/hpn5Ha4EzcxNKfOtjt9kwsTp23s8BeDjl0ghv3iJ5Lhv3v1CNA0
psPsFDt0YMrC8tfYXel0tY5ND7IjXq+c0L/23MkiDiU6tAkugKQXDBS0wQurt8KH
2/wXt5WUeOMQDdrLNz1LRF3zPxNHhP6/0hm4ArM/XibnyJRiZNYQ731IVTpFALSq
txTkyx3ZRegn03Wkl4ZKNnKLIUFyMuQL2fCs2Es8YdC8w9S/eeCGl06Wp+PJyyQo
AKXPF64LRsXWgIKQMlzCUl5alNaw06tFNoWbyoC6RsvJjibzf0u0u4iB2VZp2SOy
qZMX8c0Z5fosxKvWxCD/Y3WrnKiJ1or4/e9eogCsAo8cBjX4KAfSbBInHw8a0Fx4
f8Wq1EiDSRVlgJKhdl5A6Gm0V6l9D/yaqo44/ek2Epkwf8n+Zut0iwrH9swnnuiB
KRXOXucpIgbQ6M3QCa2KzgO9h2RA+Wv5rz9tumhNl9xHhRxYbQfNZKAQYW0BLTgY
0AdLjcYZoJIZRRMsbwGjGm4eEPXSA9cUZ4S+HZJlZn0u2/csGQ23JD/n54sh15IC
4hTnG+OBa/Ekvay3MHUppAp+K5Xw+hz4OvD/mvCt5pPBv6xogNNMeVLQRwzkAwEF
mHf6Bv+QjKCaqtf4lha3jlOkTSQFPZS/deZ32sTDDQUIZCPeWSZFuBAN8s3w+7JT
I51MEMNlkVp3yHFcLvV7m/rr5D7mna86jZ1KZbcsuB4iMTuRiRSl8zSHhBiqWwOJ
OSdamYUEVO7mxQdYqSsfOS++yK//Ey+r30/0YLzt0pF2+tjj3bAuP1g9fpdPyAe9
+qamarkJgyhpJKMcSfQlRQh4tt4vqnl38SjclkR11elLQxn10F6r2C1M2A2ishf7
VvCM4d0Cdtcr4S/EUo4+Svajb10JpUJN8udU327frL6kCiDSUfWr1S+2i43AZUlT
Qam8iGpb8BAH+tYbpv84nkzR97f+WO1VB9hWHamwDvgAb7odJ7d4OSijIbFzeZD3
LBlR5v+zNblEutahBWTC8dwpM09TcgASmHAQN9C1t2b3r4iO0jmboBe5LwKGta08
p5+UC0y/NawtZP+OwqE8kYAnmYCOGrVMh0xujH+jO5EDXAxUGvpBRjAuAByNczAM
y9nnVT2YoRPsVfBOgWGFpD+Tg6kM6OSE6NNkSf73eqm/qcolTUPSmtfvT2GZkrLt
1kQ8w4PJ/siJk1+GlCV3CVfS9SkKrHQpcqeNCArhEF0R6MklxOSwcy1rni4/NcoK
kWCOF2N45kVPKfvsKRpU2lo3uZWravnCpWZ+1pUlQjtJMMsT8mz9Gmji1uMuzgqZ
QVeG1/4dLZumNjbiMHXDauzPZFQ2J4VQMhKiCPgoVUNUK/bBJA8E9Hnm0aY4J8a5
ycytq6ExJgR80zABihr3wIBVfe3gY5sbnK3M5sw4jQGxv2AZ+Qb2MAAcsLYQU5CZ
nKnMkI/omOK1EgdeqCTE1NE85C11Tdd6biCfKZH/ZslJ0/o9MywrLLf1aXKGllFZ
6fa+3O0bgiS7WhibZXz7Qdtb/PgMDRoTTDBHLBqAk8WNRj6NPtkrtAEM1bnL5l/k
3gqC7umNuOQaX+zDT2DE2OnaYKgwcgNCW1BZ4lCaQHKBhUjuVNW5WdVB77SxdP25
qL0gkkXK9MCDaFBujVBJO+Yk/I2OW9LlFD/RZ32/KJjB7ioJiNAfwJYDYCL1tAJS
HnV8GVPcUnyXAiu6Zr23gEdJlFPG0t5oZVYwo+4Q9DJiShtSX20M94iu5c/KnT5L
jH1ILmee+iKdWGeezA/2ObwCFy5V7YicIcfPlMTbFhpFP2ThSlAURh10Vryv0H7w
pU0ZQDDsCrdAtKTLTNwtJRNz3ZPPXao80LikhcZDvDJzgFNfsI7qY5BDurrB2qnq
DRgNtVSGjURKOXHvjka8AeI10YIL7g9BT+bfCmCtsBszNuXkckE+28tsgyhwwknL
HF+e1/1qihLNHqcpcNXJUJ5ueQkdMFPhdq/c/zJyFYyShSFI1+fr+99CehctT/kU
HSgID8d+YuD5i4VQVjgeqQ4oujeWp4kYA0NU2dqxJJSZejxwU2oQtrWEXiIS4Iua
FJi9sXKbbuUJ1oCCmaIWHiFWFBjdaOjLUEBfuTbz1ZR148j80C7zC1es5cC40vor
YLm7f2FbocidKDbrZtLmuQmPgzbZAvhVjagmR/d7dRk1eaWR3BweujmwX56hSaj3
kuLuvnv2jTekGih6tio4BYWfWHEpJl+FehvEVJOLErPrdeMrBXlBavl49HoccmTI
ZkSwzJ9+0BAZFKjBxyNyk6dY1oaE7s/QUc4iM6HcFTwNBtRML/Gplkls/EmKX908
eUUvNPx7dpA4N5CqyLA+IdcOWGnGyLSs3KAuO9VXbeRBgUjwETHdDJotTfyGS/Ff
6ozwrruQjV6mivYrYIe1y4XRn2nM2LOPjZIQSYanUtraDovUVMRsazWcMsWf8y8V
zgQRR0X8MdVFKFpBRRQeB8j9COa1qJajQp+brLoRrhZkBOVs7Na5snu4gKuv1vs2
1q+e4qemBTceV4ipPVCeeCNy2PwRvzdNASdaUo9z2ArexfkO3HYCMfdVL4dYKZr6
KQOEyEkgDZZI4etb04tkA6p3v91EV7kexwMG75d0VAKnmjbu+bWWENFGpdapFaN0
Z+awnMP2k0X2d5hJ+d9lTBohNhwfQ043Rpxh2x6Q7stVnnnywuDO/NuI+Lxzot2z
XWzJQbqMiQcrly4qvhWVN+Yq4zyq+26Z2jGSbWVTkLXRhIt65YkeeTHIY/qhPnYG
+5+RsFGt1qqOYjs4NdNzZnb6pfjGDXnQ3fKdY//xAckWIUWZeGtJeKJQGuuX8mZQ
sCppbcVOq+ntRME+g6gBt9L+HBHErQiqMcz6zIgOiCO49UPJ2dCcz50uV1VXByJe
hOHcVil7AUuvkAdsgA9/M1Fyt1WGn2HcyExGKlgN/czMrjyfbGPARTwepDkuxrp1
mJlaJZo3stLZPoT4pkxDUkSzV9PxSQXwnN3Awxzde2uCfIY2FXprEYteBVryrT4/
1OwCbYLLNSVXrDkAhc3zY79Duhh5SX/sHhD5E8PrkeXRrlQLWMJeo+2ILw2+cO35
5HVA4ZHQswaKEgf/AklDEmvxYne5qKk9PIOtdBSFbB7G3/L/YgtlL22qVC8UC0Yw
1drOENXQQjWGLbMfiQeu2MZw33hecsgAfEJ4/HcWuYj0FHHvMx3qr23Z6RGmcKsN
wB7JduM1oso6aDm0rVd1Mk2KcP53GvY5l7Vwvi8jofZqXbxIqMOLGx9Nv9XjEfTN
+nQFbJeveiKU3l49oi2RMnfIWw7kOKj6VcZsjCWl9gSMO207uH2cfad4ut2k2a0J
RaMc5njUAatgZPxk23q9UquxhyZr97nqHlndcJCp18blTK8Lr60/0EnylflvCUdD
Jiq+rAd8q0i7yIyadRQ6UotrMsNkOb+37WI9H1VZgSyz1xjVx1vX9a/QmAw0OVmW
dfu8diVePz5RZPJw1UONBHxAcOqFEjAhp/kl3ObswASSNEOwnsaynnDdzfXE374S
l50iDZdihBJpz9kXvP4wwo7GaL7kZ771RAV39WZWHtPowTEgZq2pAlVqrS+b3+ek
NxVC0nZoRNf4wyikD/3XH5E7Jt84/fMFLk1ThOOeBU6NDARwnRxBvYDsKaQVG8yi
zmXShFF7o52tQ83rKbq/Kjyx5/d6T7iIuzwHSoutdGhpz4mv+Uvuv391nJjedGKD
PIEriEOqIjVdmrmIXOZiwIhTA9feZg8Dn17rC/DSiw1BL4epRGWmIXGKfsQZ41bY
t0Hdbr/R9Rh4bJ0q6t1INXqq/FAi3+qXM3O5kT3bFCzlTYAwBHeUsqYexDCe8X/2
dI7I0u7n56Xtt2uGW9X1KUb0BUsmYb9Cvasj2ROl09GYpzemSoNACEEAdDqObD5+
2hIDeKL4c0Ihe8M8fs4G/JPgJQT4Fd2jOkwctowA01JcalaDIrov2WvksIIMaf7I
DAz0l2eu2FE9JMfXa55VYPov9jWTK8lHb3hopjj+HhMSWJpPfw8Cq1oBAYrMxzCo
3pG8DZTO5YCvGuZws0yIIG7HqlvS+wxu3a/aoSP1mMdiCvmmZxm5U49vNoVb6NHk
0DUs7JRK/UVfKI5SwLPiPLkYyJS1M36jTF+MBgH9xMlPBnxgya79JreD2Lj/2jqr
MmXf9ohjFP0AjtBEc/5Xfwhn1EvUo+LKHGTXrRgy0v5fIZ0W+Ldj6SC/vVnIC/oV
OLfv4ADspqGrdRBYk+fJPFO4GdF6DNBd4DRwIAcyOAYWNG6wWVg7OoK6xxXssumL
E/scAjVjBWLbGh+xpI0bg8Ij2S3KVkpF8FjAzpVzKd7XM4ng81swdIRK4fcaRucj
M5jFxshN1W9PVOycBrKEL9w3shhJUWyNVN9L1x+gRyBNopwtL7jsIlYWaUknscJo
nmYl9amTH+nErMwrheKLS7m4cfAOxIanmxDv3poduJWahnXoKZT39t5GRWcKOdTs
nkfDJP5jwfzbJrHj4YOAhAIS+DJ3U0AzbYklWZjszZeL053zhNsciY18B7hOdHWo
E/oh+/nkUTC/LI9qYpAXZnU0k+MvH8oVy0LjS2Ir5m9XcIiTQfKX+EsKYquCQTnS
xtYjmXv6N+67t38Hw2qYqLuPQY6ZEfe/JMkcX4tTQfqnYgSVzh8ONhX6YsOVKkIV
LntxJK1TJBElQco2uYDdsuACGCIBeisg7v2BAf49nrtEEHqbM9ExrsIXkboIlNWC
2QEIhZFsT+dLn1u0x1ILzZShtJBg7hZWRsY3OMvubFpWadR/9fvUhBiPD6gmfyNI
X94VsSkGWGgoTJZ8yqBHHUZ8DSXpDjKX0uryo6spQ3gXlDjDFPRgIKD9mdy850VU
akE2VvFr7SGPz0SkIJZgJROxMlje7Yv+N3/Mg8n9SpXdM3VFkDfFg1VcYKnwLgVl
6v2/ZVIKtGobYc7kNKlRaBaaGSIx/KXDQmuy02R3hdAfoOkEOIH9SDyXrR951l0W
36/4w3APZPTycvKGSZ7snWJvs5P6Bw3rAZNAKLLybDS/ZyE5byYYfJF1H6eZgFXf
Q1pw6D+iNVjJCGP2ze/3QVbvLcp7b9E5dLBBS2HuSTw0bGSG4hbRuMv21NuRJuyL
g1Szfob5J7shRtlffqFvKTQVa+Rb6KzCV/SUBvYM8/6jY3l9r4lO3ZmHOb3quA2P
W2FrPUbMKiD0Zq/apy43lNI+BpfLFylaX8TnIYL3YByaueqwRKWKggpX+atZ8yy3
X9tZRIM6QIDetU46NalAVACbOawpUZB8+MKAQDaG+qJKFgadjoH7N9LZG2KAmoFb
w+XMH53ZHQjTBpvIEU7QdGrodqklNlNNiYLSdlFPQzQ4vhxdgZJ5Z61+Us5seKrL
g24KfgNZ3KyYXfPKIyrM77ziRQe7AhSf+La9I75iE5eCG4ZNzg9RR81XtAGF4YwH
N5YK8IE9nrg4KlHXK+y9yQf0zDm8axMMqhxi1dWXChgEyi5vE1YMcxiwHBtS4chT
fJodg0HTxaZEqfqNQIvLf/M3RXhbjp8r2YUudROtaByrIe2aiLj7ksBMFssVCjqT
L5Yv2EMZfif4zm9YibfhLWd0V5MO74RjG3YZKzN5FydzTRG33KzWx4HXL5b0ZM7t
g1m99JRNsqdtLUNh50tnJhYe9P2nAZ82y7tWcGfD5ZNb2rAa0WHRwujCAg5ChFSi
1MPRlF9RGKEDZjAZrjbFrKmpwbZOjrwX7ZSEb+HQw8GRXH2h24qCdVzot8vWP1vH
pbdDxsSUus7A/TMmrgFTWppytC6CutTvluV2Xsj/PwI5RSp5eB/KEJ9DUriWITny
hhKP1yhO+pY188AcZODM2m8KCY0adW2oRdGXCpnntho4UTwoSsrIt6TNYJPfYbEy
3ortbH2f8cN88N516VMoLlCCQLThCp1TFpD4Qmr9F9RopcXoyPuoI+SqaOMaKzMH
NxMwmCC9GcYf2FHT+ThT6msVzTeWX7fQ0KxJD+tRriTW9AUNqqSUQZzRltnXlw6t
YDxJZFDGVbZFAKb9Kys/xwOVqF/AXUcu4Ng4i3Vd4uDCfMlx+Om6AYhVxlh1f+TE
6ha2JpJWsz9QM8MqZa8KNxC6JSMDciVASrkJtzamVYtjW06cPQFVgLvtj268D0pG
SMifvm8aHg/RF1ejoeVwoIeW4adwfSxDOkvIOry4W1EdvYNF/ZJv/9JfHNdBp8un
FCEVsbfR+AX4ZrZo/1oTk6sL1X0VYlybEdSaCRJxBCQy+0dpvfNJD6oB3SWKo0/i
/t+cVnn1QHp9cFWRnuJyqbhjrZaG1MatoiKm8vpqceb/pbq3VKpK7Yp+BKI2rDS0
FLUcobQV8amA8Eo4bhEd9h/TCysyB20PJs8TkSWJ8cBqD/28PQ4WM3EI6SHYW5O7
zobTB5AFHUedi3WCg5S5uovl3CubJJl2f0BWONKlXhwmjVF0YVuGovzgpOvnRC5t
Me0kiAKgjqtgsrlvtwL8c1l4Y/yQMIeRUZXSltDW5A05NZ0HPvcZ0tq+oznYlcfj
sUVOufcOCCRPLH+x+ap7g4SlCzRJVvd0V91NXR6W+dWz1itz+ebhzmzes+00qc/6
AFCMfAf+/W9h/fTa7mbzJfSYwooy1Mtt/z4+FScplO0bHqtiXi+0pPTSbvb4qDe4
a9F4GZs73QJ66PlR4UJNYS18rhcLhmJX18jjp9grjzj1DOhUXHxGaSyZXc6yGLVA
e34zC0N/UCp9hIFE3xFm16NBlm4QZslUdFPPcHPT7AyBYuMhik/0oeLUIkwBLbwM
qIgHnGVELxy83YNCOPXyYkR9MVyRe8m4tz/HBWGQETEVEWfD+89ooSraryoDaWb9
u/T1LFLZ86jvu30ivWh5GfRYh2u9kSQVUvNuOkxSE3EEuoKLsxWU9iJG0GvXOy35
rOerzwaRPqzRm5QliXVNvo5Z6hiujogCwJPjoU/thuT/L41p8qRHOYBderjyandQ
f3DhKLpVH8aKarQwHgs1xmJJFgFoW/vnW/cc4L9qAZSsAWoWNsRcD56S3YTY8XMe
pyGMqwpDwOqLuHGpEy24iojVq5lcAdhH5Ab9MCjpFBl/TRtELuakpPeC7+K3Jzj4
o3jM7ZKbJ1ujpm2W99sMaXYBK34WnLBorl4JAE8+3UrKjWTiPKpLgZhOO2jcOPlz
TpOiMklFYB+PTRi2dBaZUJFpYFgxPUv0SdPtjLgMLOhYuJ8CxM905H0nBz8imtah
d6xymfJ1znFWFLlWzUPk8l1oUzT2FgLKpeyyzCBudu8ka2P1hDJLw3VnpQvg4WWI
KPE2k2HTh80I2WVp62OUZcD+/v9ghuaVWqFTfeHIbhXwAporgJ68FQgnYsytNyjf
FrXSLy/rTzv8JSKKpImCrRl9Flv0fXedZReL1LEW5r8SdNsWJu2CIT/aOpJvwmFJ
x19qMlPTNCRUDoPQoBo36LrYYS1iQEtyeuTaK7FHEapXRBW1fOPYr0cTVexLP5du
xSJ0MqyG+/Sk6MDcprSNVeMuqFTT00UTMv/hAZ3+RYswb/myIr0ycqA1Vdzb3PQF
69EO1AsGIg724nIBHniEZdL+BJ7G1kakSMDn709Pz8/pe1fpMpa9QcLaDW5UIUp7
w1ZJyNBK7rHyK0bNCzkQorHNqE2Qvg/weKPOFP1wy6j6oYUUktUNbcnVaatDrYbt
po08O0aY3vJFy3aNGVr3xjbs1LPkQ6AnvHMLWKoIznwMpaKxjdtbmZTaVRAQ5vxZ
2dYl7YUlAjUjCUuU+amxHaxlQdAuSR4HFjCqZOZZUN0NpQQpxy85jBXfsxIe11S7
WZ0OGd+YrXFGAAsmnNJWHsTCFCiBOdXi947cEFuzWm2rAlwesc5lgd9ikUku6lu/
3QuxAZcCLVA3Q1vp53Xr7+L4nqHiK20BmVyIbCP4qJbb93qLHUyN6fLkcafEq6Yl
7JI91iIcNOuFlWADa2J1gwnOfWfN4gzvUt4RuJkxzWMzWkm6x8B8ewo5uIFXQofw
6Ex1ROcdsxTONIGJh4GK2aYumDxj9JT1HVW32aPOPQkDsJ0lv9wGWxgotqoWOBmh
foY3zE5tOnysAHHFeGG15HUrAuZXyPKz2f1Xft1rA7YAvBJiqot59XVN/mBhKXqi
qihNxbwIFMpcksqtyCxmxg59QAE/wLyqDQ19qkcPAdN9MqTuPY/XQ5zT4jd2YIc4
U5uYxjILGiEJbsrmosWRQmbsnYlSrtSA+3971n2F98ro4Z4mIx9/OSwcQ8v+HC/T
5X2SwFAQmHI3EnDjQ6dlorXJou5R3Tp8f6Osd8fngYCqQEGHZoM6bXpbgv/ql8yk
5iZ3tDbc1/k2aZBucm9JDEQbok4h3ioCExnOf+QYa4tpn/Qh7cpfX31UYwbzV2el
0s/0Uu9D4oquFGDomnEzoxvjMMf+MdKFwaa4xvu3bB3/dP/Qw8f2YxzzqdewmRzd
qC40YZXeSS7t3LkaimRrM0XcKvFG3NKiDAEiX6XJcO7Ui1PCAjREmOBdPEFoqgZA
PVCP1ngaFXs7BRmbAZHtQ/5odWtalsWAHgoS5pQnG8jljLq4/1UP8hKXKy9LnNtt
lMnaG4c26G+V2EOl1kKvaSmm4CsxBPDbjwiNLPfJhkTGoHoDMDCd+6Plz056ZePQ
VQTPGlRTFBz6gBbGZfpRnypesNBATLhkbfiB43M5WapNeMLiLYR9wP4mdLqKLTGJ
4BDYSBgASUgOcJVWQQAaY7xzby3Xx6YkZrDJnx7RhQzPaX449WKVgvn2sUd0wnFR
FIUnbrlgC3ABrgf7bx7kEyAo5R0xrVdbaqFoNhNS2Ij7k7fJzZkuBn8rQmuy4F3J
utiRs5+H4Q0bgzaOBUl0IQFd6Zl68zmQFGBzKJW9HDo/6lKjlAhTzmPnZz1YSD3e
9jrK5pIGZVC9LL5dVc8h+nvH/cYcMi1AePZ4Xx45Vlh8CDC3+zeskSdSc6Ft4smS
q4RBMUBsKGYk4fvIwIAwc/gsgHW7xLset5z7fUR6OCzO61h7Hkt2DMuM9VDg+JHi
1OuXAaHnxNGRdmpchVk8B9lSTZdNAXkKO4dmVDJa/s8tKmHznaMORsPsRKVp9OBg
Hziv3gBbnvndvPTlduWQ6opmaNLRk/287Q9Vrkxv1yRgOlUyyZARl4zkqpBBo7jF
t4qCLGIINagDA3kHlbvyICK1FWYSWdIKVTIOBqzrjMbW6MBGHJ+saM3CwmC8/DxF
DGZPZuc6AfwkPW3EcUdW46YtfRvABZ3ETcxVSO6EevqriGdj60mc+gsUvqcrwa8O
j52vqTZD2UeNG1hV2gGOjFzZcRB4ZXTwxZ52kTcU7JX13jfgYuwYjEeiLCCoyBZU
I2XcRjL0us0lUBkl9bD4VxgU53dMNnVsbpv4riOlEqL5cG1iDo/UPUZBP/YZ4l7x
GTow82fmegXaHCK82FCyvxiicRxPOPScqv/fxOZaDrSOZKhF9HzYoR+tPzfTged4
NOVUe5BPSbfqfmkexJRnWBCSB9Zc4ub0vOFfosi25RwYHcEO64f0nW5vFf34UG09
4aGHcFquKzgXUVJaszhKN7r2DitjIlUPhFNI4zAALgs/1xCvH4RHI4u+RB5/epHI
iohRQAE9HVFY5SI0Z0mYJNHMAplHgrGNdg+HYd3/yC8SLa8S0v02rRWF3fB1LrGH
HH3gDkt8xTzjS7MRs6b01KZF66Ei/UhlmUdGqnK/sa/rDRULGRhMgbLZbWvheXjK
LsxrQ+rcLLcDavQ6AX6PXYaynMPeYLZVQ/WUB0Uz1dG8pVO0I/H40QEUka9gDImK
F24pD63w7qB2DUnQ09Pty0bnWE4lr9s+UbcbONScIQjSXuBGhjK/IkqaAoT1bQIT
p/tMmErthvAYRIzIlv4+PRM5xSwcEUrEOV0X78JI1y3iCDhctkWR5Yjb68b3UbSp
NKzqWSTnX+EzBVaS1sHnbpngiWJ0VOx0YXP91D5Oxb2UXFxT85y/IcYdVoPn+IyI
+VjBKuY8A1bUzBhXHxeg4AMO/4OMuWJgRngDNLSm4ekQs2tbTN7dIp78t+JKCAov
5IWdV9YCW4LKRU/6WpE+lvtiI9JIy5vVgQCzv0BJd5RO3o672YW4Qydp3jsIuXFd
Uzf2JHVUgbNf1a4nVZwh0MopdAKey7MfUbU/Rt4teTywsXKY/Jai66QaFDyT3XI6
1asaF66ynNK8L3gUw+apti1utGJ0gBnlHrv2amg5sSAGzDu7TlE07x5Scu9nbGOO
2koZsASmOlciE/f5JcX9ZJcYYHM45viSeWHPqXAPq8Ax3P0xh7w8/k+8Lg35eXkJ
9sX6Z6EgMo0Ch8p4z/vXX833HhysIpoCyGbeP48CafibXuSJeyquqraaqMT8qbAO
Py+iFgQFJZOTocUqqgThf43u8E4UxXBJICNUP1CKfNeC/BvKmqjlAE+odLkmKNuP
hSKLimLSheNkFj6fIsfl78QSuktt8HQ5+kkotzgiHlD5aLkOOGGnsSMH8L9KpD9J
DGzSPlWa+4AZy2e6Tv3euATEQlt2vvqeTimL6hb2EpzguRPLV7t1CZd6hl6AuRlh
4f/9KhzrThqVN/uqsmRai3YGxpvYuJjC0DzsHmsHHLUpkJAk+W22X8gypli8LC/Y
nJExrHz+Uui8rlrJ7mIUQgC8QsRMqPO+wDu8cjzY2NYP384xxIjiJWxEt0kyG9r6
Ad5LrwUuthrF96h4tsLxh4ksJKvFFgFxBlo5Bvlzu00guM5p6e41bi3ZYBDbqPrP
7HWpsORxBp6kFtbRDGVaNhFff+Qlw8cNCh9BmX2mQ7WibB6KePsbFxsn5Qr+wdKj
pXEtPFBqw8mKnWpwaBXQZhixAH66FtoOS9E1nduyfFsGKSrJGk3Rvy2cQX7VS1uv
jenxq7UdMMA8z6TLktDK7+eigY86zBykGWsAFjZuY7RsEckruVSDGsYqoyt61f/k
Ckko0II0P3ZOwxqZX6st1AprXL+nVh5hggDuz8YDSnkYRbhvI++twmUDtcsF6tyW
KIfJhUBc9FcGrLkLvThQu4ZTRYn0rCMJOYlvXzdhj8snOwCKxtkBg85BTcjps5Cn
r7JVAiNU9428pMYHnUlf0By9QC3JD9AIkqhycke/OAVqMN/n/FqalQJaC5WbIE26
FkJKsoxzh6AW28We8VLMI+wm8cqwUcMn985Y//R4x/JexosQdgI2Rznc+x5xtrEG
c8iNy2mFcR790G7xYXXZbBUfY/UAUCeactWNVOmBAXcXh46ZmqIsUiBgSgsiB93D
L87GBUh60b+x4f02IC073QeaCRJ2+kWWwoNwtd9DRy0IPECmmu561HXPJaEGQ6zP
ioteIz920FoZLIio7jKHmJhjwHRNq+PUniR6GbmdG08Bpi75yPTDLMbo6S40W13H
tuP6F83jsijUdXmfOfuDyhtBXfkZOG0Z7AWIeL/BuA8sSbw0DLyMWutUyGjp+Nce
ZHQn2SM+DQ8Mc4EWmouuLni0QGzBAa1rBhecY2RD8I9O3s8S0+LOpPqg9A568mWe
I87SOplRrbVIpDNsIxTxtjvTP/wt4HI2uWlQs296pTXlgbAIgIsuNq+zu6xAVlVi
hmwpalGx646g2QwSUsfVlTM/u9ChVUep7AUm1DbnFKuRGlAlHJqQjXz54CRmFQ4X
Em5fM0FaBzH04KjhsiOtmSw3xhmTEqrQD5QvlYm1YYtzsVbt0yavz/yCXKzaW3Bm
6W1BpKKdRxWsCfSNuywgbzpyQyZZKRx+WUGhvlTwXscUA9fy3aItKBpEPN1Do8Xc
SCyIv1w+izJJR6nU9xXQc0nRkYrSk6yC0XAoF7RlxsRtGmAhKHb3Sb+PtppULebH
TrjAWqirrGN4k0YwcfqaeqrJEmTxi6uJ4wsqGaomG2JRi8/NdnW6JJekjX02W5x+
wA/lJAV0s4j/339GNOIfZQ5h1wZsJ4YfgAi3OUfOqu96LkeVIN+x/NrQeIHLW/tp
1kqv7LR+/6+1y0coWMYV4RGd7bz9YeZjr5g77vbitq5o1uXIq+3fsHVLqSuvstS6
z5nwv35T3E/VeGVudeZPb7kt9pqcSSwp3dpx9GaqaXaXH354LM3dGX2EmiHXpm0u
txxdPSLFepgpq+jbUdWQTtwvRLpqaUwpp71hGJ7pqiPXsQGL5fCBZifrbYp+LB59
XuiqdkkHTXB9nd6kAXANlwU9+UsjOMS4b6nAxKolvq/tBHQJR/XZHYskpKYjumwe
2UVdmlX/xyMrXuhxwBVmDjKVR0K8eqz81ekpitBQHoApIAtywyrPR9ExsxDd2ifs
/HtAPXdIgZB5lgoq54zsCX2fuSxvp4Uiey8zC7hb1d4+jtDpUJaoMR5ZoSOnsHoM
tWUMViZ6eosLWVfu5DGltIrH6Y9FTYtc2ocnVp2uz7saoxnzkeu0mM7PoZRci3KD
hwHQf3n+O6qiWk39CemCGM9XXhHZw3ZhD79zweLbC48j9ivhkGVfycBGiVorE1wu
Dt5bKDvlE9NkaXSvJiYEUqNjFyFe7NkNJiFoTjaVF2/OyWNThdKMj867sKbtW77S
CEjcFf9RZCdthcdOHwHgTcEWW5z1uXorOl6p9LT/LeloDFUwXsLg0cWoY+BUY1z1
jlDLw+pZuY2gD9MJADDorAImMx1ZXFxNwx6mpGwQayt5jXtVa84VDxdOAm72Dnyr
xGnxktlhxj30ztk5WXgArWrLfKvyGrlsIyjWd1whV9mrjAvn7RBcsVvCVhrohEuC
SiTKs80mJL2VdNdVLa+hEoeHNUn4dC68DZmnokyoDW00VjeYdzQM/Jg40jHI1WBm
5pXAl6ORvMa8HQ1hRR6rZg87AsD0R8BP/PY0UdgfNBEu2/gLMjVDPXxyxZADpBez
BvJjHz80Qqcrv6swqZLL8q//zrNqch+io3XFO+dKqiHD5XV5TE0AFfCbNgLxzeM9
T+I2Tn69kYk4ZGeCO+9T/78BXwJauaxGVTrkR3Q0scKZXc357wGt5ryHuOlzlZHh
l3VNuwqd4rVi2NwQdy6RkzbSL0nQLTr1F73PfkeptqQNAQhJIgBx1Oj6dy84/f0F
9ummnRPjzvL0cBPwsR50uglcLuO/Hp+i7dzNieWqPGF0vuf/CXRWhtPXdR9A6rWE
eGEgX3NyTFojnT7FUwHBqfvNedKefWEcHk42Zea2hBdASxlSJWbywVVJkjre9mwE
WThKBR2UITxh89nTCHJ9yGhl3UxpOc26+fv7xQ/RMNizCQlOTQSn6wEd0VIwpeDz
lWQXVdNl5N99lJ0l+iS1yZX5wjrIX6rmkDxxAnJMfc+5pEFgQu04HTQtbZOnPQvh
gaoz/nzjW20O+4Cetru9FFlgenS5FRe3DHyeQzk/mH39nT2bewiFOQmcYPEx94lg
B5kMhnYd8nSvgCzksU9Jwj0vPABC4k4ZEbF+nMTyuKdBbpJAKJt+5VJFg0wyLu5Q
on0MQPp7pItiueJDffBELa+u3x8vAVpMRNhkU/pAOe3hP6DS2/hoqgL611QMHolY
iSCHoEgZtlf8zH0+ogGOxV7WmuC84c7GTuvCQpQ+OtaZFHV11OHkHkq0IYDsDU2K
l+3ZQkDtX++4EvgpQpWDWKjo4uxuFpdCvN28rTt7QA1ESqF8gSIIeYm/j8OaPIrC
Se7XcKxf5PugBaXbgBFLOfNBHSSftPSUxveschbWcqhL755ihl0bihJIKSJs0Md+
UzzoYbEi/yO0mCfRjgj7z8rDAaZhhY32lHtKSYDIUYMhOi4K/+ZLj2uzdBzR40rf
0HDirWAGNghR85FsDifHG4vkjFc6CduQyXjV8mu3G4hLLWPgF8kCasmUsSb1PRj6
TnuBI5PkKR9ZHDXxdKaoGbnUplk08wEVvGKrVzkWr9rriicks+kd7cb3wD1STpOF
9ITFI8R09XZaZxv3wi9xQcNfiufU0jnkXHHudpVm9XKu5botnqCChgD9hhYCadWy
K3IT2epBFYx7ehxazy+xZwarNTWU2Z28bS6TdxnYFMzddbUYCRGcdrTCZ8Gqznaq
fpDkXaBLTaCDNx3OHVEerCzbftWQOlR99fCgauDzcf5kSLOzHIDhXXLabFGhknXq
7FAG21/gQNIi1PayfSjbnq+H6WzMDz5c5g0AJAN4YQWrKcKESxrhVsIuUsnpAxna
tbHotZTVQGZ5YQLpz2wVTWDkeMTZdpAwMjQ2RPRB1Tf+u9OcqM081jxWICs/QnQ2
0u0hKw/GNnSSytgUuR//E42N1CmiBVV8z5h6PLD4NM/0UWRKQRB8IqlUJci3z7RE
w7FZnKb3T99tFxqIECIlyz4gmDAZ3kJb0U6OZUwKuiI8ifkgNkE+cIRZ+qKBKaKy
Z6oXi44eEcrp7+gn+ybYUyNfuEEBqgkq569NWYSWqgGzw3HC7joPeAfRWsZKs2sD
FxgCaTLld5BbZPTI4JnwYpsPMoc2zf8DjtePglkvfWxBJBRwXiRKJJZQ+dhtEt2N
4Wwq5Frhp41vtgsA/g9KcO9aTCsrSKS33Hy4yK9Wiy/UbEGFTy3bDy0yqllUQwn5
mr7XstVr6oq4e+T+zliDNYRLD1ve4RwNdVAs6v11K215+MSqdzsev2BuYGCxi+ct
BusERrrvgh5VAV7p5BAcbLOGV41R/M8BRrr6T2lro42dbXCIdhDD4qdO9WLwyOJK
34vcpg7xlbgbVr+a+Wgdxif+02nbHem+lxlywi2bphFQDwI6dYrwNaRbfU8yvzbu
r53KJNRq9S9aF1FL6oQhcgApCi4PLBMLlE253hYIqx6uZNniz6ig00g1qiGLSTMS
tn/5W9yUaO+pGvCA+Um0Z0NEDfLASSAGPr/Nx18K1cSXbRKYaiBExXBYX5ixY71z
KRYRrW9tDuWavi7btiAbV1vaFJs/Ub0wYlskXCPIG+8E/ZO+BjxDzuHUTEUalMpn
KkUrliRYc4U3KYHHserDIZdZ8nuIDCT5YJXO4/lWBJmELnQTlfonkP5L8ilnQB5C
n364A8Hasm3sh5rVN8xj3eO4V6c/OAs2Nkva+9YZtFeLUrQ0XUhOfNjCY0Yx5ow3
UHrVGL53MlYzZjCtDbnzdweDfAZJhau9NLtfdRutdxbc0O6X+Oot1J7cAK1IxRN7
KPAQhcLc8ygEjphvBFOdL5A4f8rMCkYzjBgNiTvndko5TV+rAyoQzKYZbgR4q8QA
W3d0J+JKfAsCAOhJHN0OULpBKILhFsgb/H8NlRKSpxYZd6YEzVFFiENcogqyFr1I
UqZ0ZszICtcRzqGfYodkT54MqQu2nYl1a6D27MUduLWemd7bz0S/uYnyo+kRAvBi
bOqF7DiiSXPQywd4Z9vn4JbKJ7MXGjTUv/6oQY9HkPjlMLSA/yjKM3rWa7M6+GCu
uoaNKWzrp5ldpufZr0wSTqVXF5bKvezYmu8XKwog9e8o9zSBPb1MhyhN6FG/MOYA
GWyCd4HmIBdHTjF3jI6LSHurJw2tpwcMnlOrXlA85CFSkaDkDj/tY5KtizmhXfma
16LBs0TEmUAe2Q5nkRICpwEtb+qQKdOzYxleuExHyVSxPqmTJ/2rZqtu+buc29kg
OcCobFDtp3D/W1L5DJ6pcgriDYoLN0+OuXzDy79BW2dSSi3AQs4MqAj/VzdkkRKe
mFAmv5R9XnoAfLZj6YKuo8jWCHfXgqo9isjhdZvO5ajKRLaGN0kqbsZDm3srAMAB
Xuf+gge+KqjLr7pBCu0zt+uTWSF83TtaHyc3CjTBBG4Yi/bslhZB4QbXnSjYdn7R
r6FVe9y6vhVfnfvibURnmxynPSCey6cnsP7ie3ttU1XyJtn2hQPY90/XEqZpHXkj
YDp/k3UbWMWToKVbeQQjvUZFvy8kc1DFaKW6UzRcaTOjBKroeIVyYyu2gTaS6ajB
7SnqzERum2keoLYssmkNI4Ky7lA/S5Bsnaz26f2kKLOt9B0trZtD2oRXiv5Ma0UD
R/gX4IsRzHWT6JtedmB3TsFYO82X0AZ6eeAiEWZ1SZKDy6k++Yv5zL5fLYSyEeAK
tX71eeg6gPEJqYxDjmjqZzWz3/ThaeEwXfnBKeqvN2ptLVi3CuInl9EnQehSAcTt
OK/exTT9wnn0aPb0WXcGsltJpc1D8OC+kSp1mOEk3lQW0YjWe1y9W3/R3AxyrE0W
B7zD2ZxqICUBTK4y/GntvnUZAQt19hOeecJ9YD5WkdAUt5VwjcWDSqHwFz0Gf/oo
fVLKsVsMzCssCYSiXQkn8WrCe3hTqwDc++CS8oU+By1ggcV6a8r05bz3nRe0V45M
Sbir2rMbC5hJq4/OsWvMXSXUwUzZSOx71R0ACDf5Xq5eelqsgb2dWpyhuOSOqB8Z
r8PQdmf37mH/kILf44mqIAI8xyETGXF36SqLRckgTs72X3pEDpvOxspxut6gt8qF
0NfDgcRPQPS6RvwIXm6LgSqYex1Js0XMjBW8o4EfDz4btSccMH9rtQXDMvHBLJnS
yQt4FQDoq8u5maPJ6tAP0TheyOcV3LWLHnaarosIFVOQ0ft6NBbAbwLC+8/n8YYa
uiSduvZN//IvIGTBNSVpDIZKWfvAMF5ZfUzSHIDKxQ1nbAtEMqbgGSeJ8sBCM0eu
imk9FK69ECYUnADuNzsW6h2vqCf63t1jj1+Jw1ZaPqIWxjO0VyOAjQ91BJgR0LFL
BZhzBRRMhkT9T0241BeW085+USvGzJfbQTKrPPIcLn4VNA3EYll5B29HTZQTMaZs
QyP5mkNRIXiqsatFohuC1NpO5YC2m4i/axlT16mbP/DIDWznADN5HDt4XUDHv/8j
dNeYE/52s6GkawWR/Z8iZU+d0IOXb+i5kH0D4+V75dKQw8RgG85Clz5GGL9burz2
4ccq9tqt00QhUa+AyTLJ+81gd41/IkxxNJtN/yS4zwgmFzpZBYCfX1SRZAaw8fYu
q8C/KhKspD9Qy1f1Odv9p1wN3+bh9UKJ8L6HFDhW19aU0TsVR0FsIoL8AXSLPPLx
Tv5WCIOgGao1nd/2qtsh2V/EMzuDdm9+uBRkVuI+JoAZRI8lGEygidK9pXIf4hix
d9tNdVTLmRebnRamxZtIE0KxQ6VQAJcZ7J2WWBPqtjVgW6/ZHTa7CS69COR0YKUy
a5XcjjbNd3OSh8LIpWMe5AmqGPkCsQE1lshVvD+LFdr7WzIX9l36Rz45nhbHA4Af
w5fojD+AFjfrCF+nFFzq+x6Pp/zKjlf7i1LEG/tNV3O//VNSWGe+MnEKb7l38UAY
PxSvOJ8L2YdRWN1Bm75DIQyKjk7fwkTYMYK6VZwTSU8QOtvCYOfwu8RL1GylPeOg
ji5whslpztCjfX9FlBKuBU1O9VVgBgZQFre5n8wHGWhugJTCRDlDrqEd9czXxPBn
4FiNzWWvzME+qCSm4/4Im+YXQKObUo4/UQwoF5oIFPbQh6FawCPaGR544Q7cX2q1
jy0tiCjZEdf3IGzcqGRLWsC17TqcxaHBn5aAJCLs4ijFpoKZadI42tcGC8z6l672
rNuq0dQUdxHJSBAMw6lWONwGSUekG6FuRLMoEI1iFI1xweOdZAJ/Vk2ND+SZg/cJ
mYsamr9iGMhNlxx30bn891EQCvlo7wJ7Vc0YZ8XnDDjUMMIRslfrXkHL0NwhmW2r
u8OlBc278rcF7Qk1kg6fdab4CaoNj52K46AmAMyjetVn6Iv+j0QxJT5tXV2CBrpi
URAhPwp2gTWHZrokKw621TWO/ReZwl8JMxRJjn4ACgXOScIxfPllyc2Ab0/4Nnl2
Hiy7mXQkQ2SLEi83CdeY908fOHixOaHr3WTNrT8XwzIZCfCGKC6r0hj+dgWc6TMW
I5rwWX0wSGoSxZT7e+QGJRM5MJa1KM7v1jeflJtQi3AUnifFWCQ8ZPMnAJznkS4U
j92OZYA1Sg6TqBr8lM76SWH3pqnjVkc/fV9ys4eqZNjrAcuOtW5Vigp4w+lha1J5
LNk9fL4iZ0f1jHsbhE90MKLdGBbCGOWytaBgKs8q+iOVKfm/Ybr/XtowyRzx24bQ
SoQigTs1JTAMARC4LV2djvqBwU/dbw3GaMHF1OUWjCMC3CysGmVcyVZuHBs9bUaI
0wrKyC9a7MUsZcjsY5nk7YPBVxmR+mIKrOSsziaUOwxYNv+ALNmFdKGPPyfNq+cR
ZkF4P5lJoWsflTkAOyH+xRU+4AST2hp2JRqYpfrJUvM/T2bjQVq4HMokHrDOlEMk
je44xArDsbByzHEIhxFplgZZkoChC1TE5virGsxfpj0yvI9+3HD/HM5ozGeZPscE
a59oUjsvIWUpbieWCWVyPlSrnnrBTw48c5+FEHResRwlb9XDv8PmrScFMS2Up6YV
7OR7H9rUyhziWTbxm+s1EwvY3A9jc9kKcSLYEY+WYIS4duHNJ1N+5nyhPrVCaxnQ
rP1Nvf6y8kE54Oube5jE5VBaMsPLDfC6Z7Mwoov16udmDON8BiIGHix7uQNj4/Ll
3bOOYL/otQ1OijwZs2yUe05M45jXRE8jIr3f7CYL0DX+LU2iqmY3/cU5/o5uZKi4
p75WIfUL/5FGJ9yF3yWV/sFP0l7spZAE86Xb4vOFfu4MrgRuB/evmaz4KRKuXob4
giRDuAyxDCKRiIl1ZdN8LcckC+LDuBzNUpF8Xmf/5TTAtDuwxOCpFEPJ/dcPcA/R
TQMJN7C2IhjyAnh4QjSxttTAYVmFfcfP+dJPmQo03eyWkonyIL1Qq2YHhtY4tQZc
LiuINa/U+PYudYcUCGgQ+OAXG/ABcOUSfq0HGg7SItQOWnkXPMfJva261rUmbz5P
PhSOncuJAzNp15seFNw0Sj+hWl63uVwWONMqSSEl4qWcZTll2lsxow15LopFr3tO
N1yTDWITa1cSAydoGi2BpL63ME/w8dJsa8iKN9BaebxdhoRT6UdomlNuShOWJgzC
gU3/Sxzh+oupgb407vwEW5g1i6wlpM2qdQbw1v/Xc9SS+iikEwRKKu+z1f97ytWO
edMJ4swZFlX5x5WIDtQdbFRQBD5o8/VPhfQQYwhe4lbw84aqzkKvP9w2R5l5d0AF
5zenkWZtF3DDmhmyIBXoqE4toUyGiCQClkO4oZT2j0lYm03wCQK1VQIWkwGf9/Co
2HZaoDZZqowLwq9SmQHkQ73WFNrJbomFObzG7T67eeQf/4E/kang8/Pu4//xIwY0
Xsj04gzCu6oOdBC+2MHudbUrU92f+14ez+Nt55jon40aHcjzC7hkt+1Q4RKH/Y3+
dGqIyp3x6KhZuvezdRCEl/iyZNloxCROzc9jzYQj/1mJDlzNERqlUxFYciFID0Gd
hkxEO2kNetzR99zqRAbI6YmwuQszYyAZpp4m9++8l+ZlU11wAUwiih/3S9kSElIt
q3MCfUEl+xuZlyy60K6spviTPKbMD8T9DEHP2J2pu6wIFMcUIEEnvPC9IbD9iv6X
e6xApz1vJkRzeBILqrwF23qvuFyLN5tOesg8dtlwX1/oH7vRdZpy7k4Sj47xy5TO
nS1WN6BGXFnqm2xsbXbaVTD0x3Fuy+dsNcuWgHVeX5vTsDjdu4Sy6Y/QKqQSWFa6
e7SPD30VfUYR/Ji+sUrtYwwEGYMDA0CDIG8+/PEKaCcfnnsqnDXySUZTPVu3tCPP
XKWy39+4Jh5caMAxRHeq4iO17aq37SowMXl+jObM/9LxnfqI+WxZytsuTkg+3A+c
E3pdd2TkmK0VVdCY8s3nlf+iPLUZZTsoI8aEY6bwrFmzcnc5/U5vZDVB98a0cP/T
e1wJ66h89P2rTi8AZrYiHGCbtpQwrbBGhJgjHfjEnH0zqmpfgh9fkGm3D4Dw9w5H
QaiDL0on3tPU4uH7rC7iO2s2a1/ujqvfxQB8NHhxh+jMyIc1N1CI1GE/RyAFDrNA
5qxJpDhXKCSX51byvwf8Oh6JFsCS6fP3kP7h69wuEvQ0CsfQkK6cLAI/7nYX1m+9
CLPaDsZaLeGGkPNo/JnwDQYzZ05DnPHk7yAB2YkDlWhC7P43UiH/zDL8oFfWVUP3
vYta1SJvm8dBoFQqTFpvzB3IobLRn1ws0dXK6f44jtv16Of0cHwzDtlBjsBP//pO
FKEoYbWwB0X8DX2EuWJlbiIXuBSwc6Qf0fGGL6LnJreAN9bPc2dH8zqUJe5/IGaT
fi9t24kueS+fiwXxLnXcEhI3pVfyMWzYdtOOiMHgViilJGKraSNu5j6QoXoTKCpw
aMbvmtFZkWcz8348HQ7LHqCZl7ur0j0Ihbbmu57s5KDAZ9DiydRdGfL4SJOQ3dpI
RR1WDXCW//LXvWN7ykhuG/4Bk4Kd791qpMZ9lWkplp9akfZb1oykt2EqWLDm45HA
UWuf+8KaQ2HwliGY1j4TtSy3gGnyIOqgnfSzmqxNi+LR08A3F/y0kXc73pGdd5Rb
BZ9yQ3xGmkH8B9qDDYBKbVdRqR1u+zSyGjXpubebMh4GPsN7ni2wPzQlYUIkoAIx
H8Gvhv9UImgeYVapO05/ZhtjoAu2yIFfPoaXIluc+Z0OdxEAck8nogvMrBIeAnnn
dfTP2TS1A5rn3jGZigfaMcRvNGHpOjDstCSsd3qHRaiSdH9YGQxpfsL8CSa1nmT7
VjSRoog/nGw+Y9OZU/I2Kw49IPsvSI91VSE2SINK9spWfAkBFL4vK7u1CeKdb2Dj
8rtKZERvifxOGdLyW8wbR5+1RIBV3udusj1RwsKruWXGZ5EmPPCNu2Rn5C8AJJR9
6DWeQDch9hPHPwp6SG3c+Rx91gHWA8/QRvf8xHfY2ow9CY8MpFbT4JghpqILAUgs
hI3ZF+E2N7eRlzIOJvxOBnqiq2oFnRPH303jnZ2u714S4uvA1NX9EyH89dueUvBZ
SrIehd1f1F0lwTCYzLtktfBpUdw89DUeCg4UHgxhvRlQhiX/XYVOqMz+gbPHheIZ
aNK/c3ncyiVJMtd7Wpwk+dioJbtE5s7nQWQnUOZEeOXjkDf24ieVd1UA/GLzl/3u
yXUS3LwN7uZuZMouM3QtOxoxGTwKLcA4xWAowoEe1ejYv68HoPsbYXOp87EzmHwi
ggXNgv41s/ZJApu+bq4A85VlxUpuPCrJXwUZY+/2ibMDUIpu3iMXpA5kb+bB0YDp
HAYbBppvJkDQ4ExuZJMK6JCvmykgOxf5nWEEDLe/N3D31DxG3vkwsK5YtQ4wZJkk
ho8H3ygwkcu+koSenMSrxrhsLIbexAdLaQZDP9ZEf4jtLp2DSCeJ49BMHnZYpI0J
tmzliB0mM1oddRpNrdS9srXGLlV40g7+vFizvJJa6j9ITNgLqCt9KdQctX8LNPz/
AizPSBN7/nUL9zrCiFvjxjbkXuT/f55ZSvFjFU7T79lVpTWe3slR0Tt6DGoynDHS
uRozS83hUgmgKDoD1ALM5lZn3wF1zmsv1hrz+hr5KEe0D884en7R8OucYr78OF6c
xWv8w69C/zLnu2KG9txc7fEuvtTMYqnQ+62v/99dcPQAhiQNGO+adkAJPiOekdPC
QzSUsEJF+e0yhAo9HZkmbv8bCca+Rctquq4ojoL6h16znXIvVSuMqqMH8CyZscb5
bjXdgc+fFU4BQt8pE/ls7eh3D46/1qeSRjfScwtR8076zhzwY3d/Qmkhuwc7Rl1s
K6hg2IYh/ImrwcCtYPtFJItp2M7/yxWbgyBydzwtIdRSRvZSLXuR974+VJ0StjRM
qyyNABqJt9fw+O5hnKS3pczlScAh7BvB+h54xoCk+eM8BOKzrzkB7qp/VmcuC/iS
b5uOpRyUgSQwwVn/NOuIqZx8k1LqHzlgPhz5Ix6LJ2VCot2hpgK1o/F8vqfhtjN1
5xaZmsXvQr0PuCRH32KqfY46VSZA7SSwPYfBzNdqOHebXH0BLjwGo7n3wujRds/c
RkDsIilNQz5i8bI5Bk/jfW1qIhooZ83sOBH2fG8EvVOBKc9yxOXv/5e9j1JSJjmd
+SyGLovjTZqHF5zZ/QiysHWDI0QxFVaN9TLxjdpgA5zchrweIwHp41ZJZD+0Ec6R
gBUcgktAgPhPDkA0r3LNEs0I3MrtyPWnvoUJp/+ou5fEX1VGR/t5o8UmQH7xk7hm
EHjndo9mkYqm+ZvTHuG9nIZb4ZxUUdCSVsC/wZOMy7MTga+mZPQWvthzG5S148rB
lz9QCXOXOwYdh0Ls0AwqNzuortJPJatUI5X+RzPQAXc5+nKr18J1zhQGB5I0wCbR
9PlcqouEbUjjaCQLxKm4nQpntu4WqSzZ1XrIjGUZVwoJm54+46+RunYCUqJG3zpq
Tpg3r60UFG4xSJhZvqZpzux7ceAso2UGwsZDLlY72HcPClxgCC7omz5yjsU9rlPI
xRk539LBOKVi2haDp5YNyLoUgiWDHvhq267l0zxoRBlQuZsRFa/YIaMkX/ne4tag
2GM11LjBU23cDnzplr6VO0KUrdN53u5cfeDcaUGZ0Z1ApjDNKhEw55rdtxH+rWMx
2vLpXouLF+wOFWlNsWzQY2ey/mF4CmDV8NjOs8pqZD1MfBYA0/C8VxHYOVNOYYpT
UeYmJcgN324koAUK2Qnz63+IgH8znHiGhbI3RdWjt9v7+6XAxrzLkBKyyx33Vjl0
CBDrVfNexvlQ0/gIcKn5yCflKdCb73m9fKD0md62escgmkeLpOV1bJBPbqFnlL/T
/Q+amxM7/Ewca4CHvwGmG7m70ExdCpYpfThpkeDoOZKlrXP+Vb/IX1q5EuXE70qW
ghjy0exMEnDqoKoTX4Q5u6MWolkg3FsRWyv3ILNpgrWR0wWrV0jtq7k76jzjnlzA
iJiRxmAop/eRn8lhqYOj1tSBGjAIevluP0iASt+lWPIy3C20kt4nPgnLzhBt1Kj3
v5KHhiAVbadI2PUNltPAAxjkVak+TvBdTThZ5/opWMi2bXwaQvWDHyRifBduaozW
b2ujr2nAirV6NSxc1cwe9KY9YVlgJo/Twm7R88Ym+D57BlxuU8MmtVtmq/tUwNtQ
E2wK8dnO+6j5+8CNlvwffkmnVLIdIuPsIKQxweugwWjAkHeSmCOt2ao0mxFTRWyX
u9WIS/PiGAWv7nS74LZtk3PoEzSruifTHo8EUbyhuRPD6nos4BpMGfcTHHQtNev6
BDRZJErm7zxtKSVF2Gu3zpuAHjxP+MDz8BLP+BIM+ZQ9oJ9aVIakon92/5Ttm87a
mCGnt7bG4fCXTg+gVHzZjZVqn0WjaYriOllIr1NuAquuhZie3J8VPn0GNIKnIS0h
w3qLGZ+prEn3yHktEZXf1L8b9379feaWZPgIx/W+PbOdX1soxZbIw+Gs3OFJ/Bus
TD5D604Vclx3ovg8eEU7sZ8uj+q464bHqSX8YV8J/MRhS2korRPlV38/AXkYdpZ7
LAJVrzYVbvN5ZnDM0bAwuEwbsNxW4tDoPwhGqtc7y2jsfjAYantMRcD/A/2jMQJt
8VxuZJgP6WEjZh4colSPVQ+ueFXHnyQhMvlF0u10mjrzJ8Kh3IYvEgMMKf1uBePR
EozpOuCNEXGQXAfOMt5+qgRZ3x72fCekBBeq2K2p9n908HKwy4Qg417quLb6OBXa
wkwX9qumia6nFXV3rIPS7ASSbu+HBuKecTfu4cjoWgfg+7DamJrf7r622G8zZ0NZ
DE8oGK3JVp4LhAhBl6RYFrXAaeb2Qb4dEA6wJPuPV0dhpi4somaV7cBY+ug9UKbQ
MeF7fcQKjmrHBhQnNKgRTt2/7YoF0k/idLYPOAcCGMCneLJKxelFz3SXTotC1Jjt
m1ZbAeadAtn57MmV0l00hvCYhiuDvfUvoZ6LNyEAKxAi+whb2rkE6Dgqm04EAfWT
ori4kcqYdzCD3d8eZjXbx578ZcKJxIbjnSZ7XKO9oId6xrnUJ8Rcn2jSd41F9HOW
Ov1sP4LR3Nqz0vVUYh/rloJOA8HxQnJI0+vV9vh2jlYOFjXBEg+emNXENKWX8l0p
ud3xuK1kw8XuYkPePe0SgtGKkt4IIkArWNiVpiIp6RuRCLI0hA8nlKjsmcF1z3Fb
9OH9F7hH4bamJmEaJlQFkjalH3miqjtElSzOGiIuJdv12LTTSK3O8XK8/+bCzt0g
PR2isBacerW29yxfbPif1wD1wJA3s7MP+ZdhKJUGtatwuXlbZix3de6pOJhWENJJ
fjDG80+l9hc5+NWsNPFgLGatVdJh3jJFcAsYEPuN8g0fY6cxwlud4JF8QW6ELluU
1vh1iYSXAH8LjmrXyG3pBRD3A9Q/mcpONU8jo3Wiy84IeCoEV++ZmljIEwEaDqMc
CCu9REEXDRxSBGCeLfE6AkYzk1kdiQXAFhtDe9+f2UciOqjdVCvaiPcbZlwsVyRU
/M2dKuJtc+fDRirbbw7qqMsZUFN1PzgjtHHpDR5h+YXMKmhEe8izCJMaHV4Yw/2w
5GuPeA8LTiQKOfRU0ALd3RtYUTOH0GA8BHVfzfnLSnqFgjexbYrbTynTwBRUeRhe
gobDo1OBQv7zSl2NCbgAraYtStuOQShj7T4gKejmZO+tPSCG1miY+ocAQmb1WJ3y
Aj/mnaC90olwb1ndRD9oNCKOpX5FlrmbWJ9F9PpZ4A4m0ypRzyDdRK8tixN5n7gn
C8MVBuxXbYHvgBQxOaYZrRMHmTgnKKgMF+GviPYoSZ18lR2nu6AWpM9gLKBkIAP3
PerATBWXrQrrD03qsurFwWtPHLm0Eg84DSXWrofiuQkefBiTEppKockNP493J6ZX
QLW4/B4OofCrofFQdgnh1PHNLGBM5ZjTSFZewOSPT+vR4zz3vWagvusac05YJfAH
Yb/dTz1s0jZn9UKIcPr1uO9iOsF4AEJNE7mO+mehkNo1bRfIG3pLXPvv+u7io8cd
vuaU9ce+ERUnEbY8UNDvB2MBMept++STD92W6CgLdzxXdYZuPB35JvPruDdm7cAv
a34nsDFn0SExTXkd4FjsOLOD6TnbjE5oi9WVpNyLri5fYmUta4E80MXGjdaaAdfm
27uMfV3GCT6b0qyfEw/DuTbr21G8KqHT5lJnoQtHA/fKKC33zcTVWuPXsUlNf9Sr
dYjhs9VUVljyq97MltmJVLRgm5zp/U8W3I/+foxQjXa1I1MZZ8tccjFHbaC+AYHH
trLpWwuMeN1q9n2tH0PhtuJ5KTxyNYByNLfhqhdD2sI3CsGKSbNS+ifjCzktzqic
EgRlGbccZ8O0CY2UgQuJknGpKYgwKipfIECYIqWonRJS0Ajz6ruT5ooQQbHptMl4
HtHaEbHLC7pX4iaekjdcPu1qWQ2uOSeO4sqnBRsQV/LELlEWDGAB/sJDawhKXNJy
sMpRWPjo9I+cDbZIpjZQR3TrxyFl0oXb8GJQKVaDQaIqBUA0dXOCGWQsJZ6RwAtH
GcqAsnGJiFeIshLJEE77pnxTuO+au1JjT8XoJbebp4UvQXlUKMG4vgN6ryYLUYcx
OXwhvsHenzk4A/c1I6EpuqqNgqgZamvRp7mf+M9vUNZbOvoEeZekW2RNJtBuGynp
l/JPy3Sos0O2qeWVHxKH++3A0S8lGCukFe0OFA5/SPMCr5PmxFfGXmbBclg3hEQ9
kpQfF0rJFmSTdlZUaauIA5L3jY/euzPUIge1zrLTjlIdvWMdf67VAfE0nhUi0g/F
NYhY7+E+FgGOxtL0VqvEhc1C3V8iqm3ZviqD4foyiicRrSuinMMQeQU5eBqBBm1l
gB8HNjLHUWk7hZ0CjLcamAs7EwUgSukicxKaU4IWZDmFkfY9u0ih531FuHDXsZOh
Fmd57pulZBDGc8vErJ/niQTpE/+y6IfMFiezL/5QcZJskiMu+oJD4Kc6JUYyMveP
i6C/2MILGto8pgUiNUHmBYwWTjtATq0slQ0fi+5hgbVHo20BITUDTeoWwU88eRkC
LdkRBBu2ElTmSFW9ulIFa8uBC2HfEpx7T4t3OPEb+yFGVN0Ar1vECyCPFvEhmiLG
hncRCJ0jSnF11f0gHG3WqREK3746sd+SdcXea/8IKhsT3w2X/ZCrL0ddQTtBH1Cf
iJswaKSVA3td2iAAMXdqzrk9K6iXURA/pcvqA7SLmQq6w9tH81p7LTyp4hTQRS7Q
dgxBtyja9V1G2adfvhgOJZrj+MGUHTjM0i5Y9GMoaQhqvNvqCYHd9e3QTgthvKVw
87zYY3z/8aKm2r6jXrpIfRJf+JIpCUEK6PwsK6roPZKERqFrfZs1TstF+XouEma4
OTxGRcC/4p7tWfNqh7mLG5SAVN0nW7fTohn8gm1H/ON4gc835g2qOUMvC4CT7AY9
NE6TMlQXlebi/5yi6mfkzKE2fKi7TuLyqB6HS4h0QZboUMo1kuK9wlU84+6cFNLT
ir3mSmrVDhksLtjYx+hwM/2SK9+2hhCmsI0F9/q47vj/W8Ls2es09kJuVu2B8VWB
+VvnLsWl4xFZ0AO1yfjr+qf3yEcHc9P1ohoflXqPD21ZcnQFzDevDVZ7ZvOD/m5x
Bd8SZA/Kp2a2iuXB0DRwwYYiYZeri3zTprvIbr3qK+fvTCK87WQVZ7NMh+UvH80z
kNzMo9eWHkJ9HWruh8vfOhfK/eL48CdWaHCasFdUdgke6EGXZiuuzeWq6fT8oLx4
uBKxpxOx72MIIWuC+hvLXy1U4gQlYaKVHLAT7MbvSEiyOOWrxxFdSrk1u0neJ4mW
Q4jV9e6ROeDseaNdPqFTm8nT/6itSKom3CC4VJ6ASEUui/PXVx7ErHlAhtfa1Kgo
CNRhTjvwmAjZp9AeI2XYSeJv+kqgLx0jG2QYFDHw8++cj8LWLUjJpszvJ4gxq+Vu
trWbrmiyNOOEsrtZLWfJggooEKTG6Ng7+uCZkIJPmPrpal8UoDE2eiaDM2WMBrn4
5S5wF8S0pKsGi3HQABK+KhtTvEDi2sAlrGg/FCn6TRZ4jYKkjdypWHRd8QTSp1iz
k/TIfEH7ge5HaaaLQAOlXKI25SwoyqFLX7MyoSqQ8wSgBAas/JfpU6fbadSOYwfe
gPN9XXTr5nMwuDKrsfj/e9BZqSAp7JmoVJ8IxArqG0ohZTv9WN/5Oayw/o8JdlNm
mMOoNr1+nRed12pjQHk3Xemj3gNfCrxiVx0Yv5j1YuRMM1FE8cih41ip/os6sLAS
BWvppOmN3vnsgbWcqq+9TVDnsIGSnxuobWbYK9rXDXwYNjnXyTkIbfPwzbzQcAxv
Sg7CXUqOqNP57y2iG8HFDz6nh9tKM+lnkobkyqtvBHBA2JPfwp8dD4PRN6Un5DMm
7x2/d6gqy1XutpGrBfWT1fC8cqwUC0E3M3ZdmSJv0nyU1MvXUQ8FpbusvljtaBkh
AQo0+tGAHHT+4lJspcfVL2nPwQZafaYFm6PiEH8NonbnyieA9gRDwGAIwoBStB3b
wn3v/6oVtC7Z+2nRz2Qg6M7YOiKb32h1hnGZBG/OYsfqO4DlIJv1fPAfjOFGqx3h
GBWFp49OVfeZt+bosDNpRFRSysugUdZWArv5Xsoaj5POlrSR5alYMmEFelvI2I+p
q/ChiViaFQDl+jtkExgKykFvJBXyIbVs9HVc7qeKDSEAs2MLvFhJP6RwexBeMEMz
RWvXQw1smUAQkYn23660YR3q7pSZRZPtnznJE/DNBSQcU0Gyq0KFnb3UZHQp0O75
hHUK4QmfQ6WNcCYhRxtcExBK3D8cB+izkNGKcm41VOvzxEdkUXHf2u6qJt9glrcc
wPDdXE1hyR6CFqQsGirbdaZTgTvBZ+cH4TUuRI1AbHB0GZrDS8WNJ6ygZ4mFm5/a
shXp/yyt19uj2M6EisGplG6BvoH4qgOupPZd02COurJCo4sQ38mv4yD10RBacI19
3cNUvF+DycVKSKL70uCdsmBBeLvsIsMH7nNWihLtI2eBf+UirImfdy+CWGHIRfy3
w4gHflz0jvcTAlZfj8soCYOEK9ESx9XaB8uN00QgZ03roWWo2hTKDMJusSMzPVcX
L47dpA30JP9ww/MkbofFjqcFrec1u0oaeIyx9IUsAcn1TlOEwMANZeRLXZZL8V1n
TJkyfIkG2jYO/IGTW60pWcP3wo+KJn+MnrWYSbohH4KT3O9S10rs0xdIvh1ZbqjN
hBTaDHTie6VoPJLK4tdcfESlr4V7924bNwfZOP5PAaD5yN7QPGN347025UXLxfcf
vvztzAsp9hCX5vzv7VkuQZrVDpRQ1Q5QgGD976//vOPpY8+ubXA03VWG6tM1wFFa
fXgqEjOy9g9UG1qcjrA3AXVeZTCBso/mCsAeWMzHgFn2yhI74VdR+4Lz8S8qQwUj
TJcJBUEyBiaAac/aGHrFKqmVt6frapWArzvA2RGu2sh4QTWRu/oGeSM6GLYGQWvk
37relCH7WjjTcb3qsP0JhSY3qs2j4zfR3SzezAhVHxS3XV1hsURgNiXp300yFcl/
NIzRLHre2///ofPGwIneFLOyMlVoBexY3OffcOFUTvRh8pBxOrimenUYRQvSpZqO
XgrdcFMzLZ2toXUlSj9pmZhrqq+EeBg+Gf8Cj9Blde0CaoqtSeBs7cKBMxJ1C13r
ozfHKKZ8YcEcUA1qP10cNR8kK22fhNRmwAaOGSzZuYvcvqC2rrEFNn7iBGFTdQj5
1zu9xQ37jlRF2eiDJ9OPg1V286BfDkBFPDB1SSxKAEdT6SxcdlRKyqv+9UU5DjH3
O3yppfOPplrarbogoAcPXXd7IP2jyk++OE0X0enxDJ5Js+Ovoa+Flus8TaD5TIgG
Hrzag8f4qM4KYqGQDafdjiyKZKpgshzNtM5Hk1OQ3Ljo2I7WedXfh9qPioLethc6
lY0B7vP3GbJijB/08yB/b58ddotZ+XL0DyINOUeZ6OunE934kwOvoyIychUmfROA
3ZkfSPFZhCeJJBLjJ5WyhDl5no08IokZdB4IFX1Io6z4FjADBz+IWjVZIwSZTj+5
VCJmXJMWIPpDQLw69BlyNN47GMQA/+3cY4Qzebha4kFjR1kWY4sPvqCE4QAM16pB
4aUAEOMfwtv/JK+b1WAyEDj2iaVMENdl9UEpFMXX0Y8eK8GuuIBSnsINY9uTqx5N
aQJuzhcE8FrdpCjh/4rcAIIGmNAizlQwrntIzO7Lz0hAfGmDdlX6CBW6eNWeGrHp
r8svyAP3DlsMhB3D6BKQ7lEqLsQ+inNC87cXoCXg+aRK/H1spCXc7jNcMfgNo8JQ
Mk2gvends3w7H8RpCdpIOg8hjYRZ+LYg0a0lvnBr3WtPasacxiMuXVTqyMt9j2So
M71eRK9sX0uMMV8wTxY0z4yYQiPXh847QZAR7FUatsKhcMD2ZiNkk2zYgAexWeFx
JNQwzEbSpWuNCnQOyY1m4YRU4OOLGYpF/Sz90ah0HoJQ9a73QbzKrP8Lo40CKbfY
6D4L3SkbmdPvJIk4AVF8mTmKHAW56gv3dNnX/CR8shZnoMKJZ3hwKvy4MppdWM3O
Cd2to5iM+7xDVw4u+YAax81lyu68tKbKem+TkOuoau/NChyaXc9fCywIFM25HaBa
eeVtAkKtOv8wBFz6tGpz5j5HuD4pOHi9cA7tM/5J/SUral9I7k1EtU3cbQmFFyKl
qKXDIdm26bXBV2NAnNiTVQuXB5oZ1px8iBo5y64CtgAD6+JA6ozyABHEKGRj+eVZ
EMNreSuMlIwQmb9Bpr1dqn+y9Ffs0pWROWPlgb4R4WVdm3h6w6Lgy2cgR4tM67hb
aeAliC2wpJi1m8Ry6NfYcDUOmCx/lS9c/0znVAXYYnlidC2hXt04cdY86/hhWAex
/G40q6euaa2NxWxHDZwd3FP3y/muJADe3/+Ix3UdkSBgi3DAVLEYj4q/0likrTdz
RcHsMKSka6DVsGuyX1EDixYBxe2LlQWlB4gUzXOd+Ocwmqsrf/Zf5v1Y683QAfVM
5FK8k4wxoNQUahJGkIz/0/VtnwfAIYSS3tpGyUJLkdTVc5QP8CdSbaoWECK1q+X7
mGogyq8jp7AmKpbkHmmN++Gmh4N2iDotCYiKG9f7OxiMrCg2ooYkYDV0jBKESS2x
TDMnKa3kMw02ryD91pPUjlyoOoZuE7SArlW8PwOuJrIoQnW+i+9TwqLl5XiwstZK
2FqEjhMw/kv/AOYWwvSHwaoeywvbQDaIRrHiAzp1WN/bXV17Gvw/mnqkGck5Xo06
IbO8FlILaV+7nonf7c3ekt3ITXu8LvDtQQi9sBw6mIUdS9A0ppcWIxvAOndcmwmf
xKB6ZOthZlFB6U97QOVVOOR1LrxyRIh9GlmWeFNNMKHS/FuQhI9fkKKsTPKUEgCa
kk0mK/fuNWPVXdOg/yR7/R/YLIdrbIikfVswN/PbTMcGgczdKdAKP8rx5Tn03uSd
h0fvySQC/3FQlkI4LY0KmAKWSxIZQuS35TS/WxkbpOYA80OhD/EIqa67paaFCE3F
q9FT0fpTsCFtiU76h/bB5a7h0ZQy8AUvmhQNtYRz0cB2FRi1C4h3a/MmFYvbhoI6
vIXjBGz6nUHTRIxUdMRiPkyY3PLjNsq8Zwq68sm7GuinVGrdKtaMyuR/HoVwxmG4
GgYuy4JR59iJNM7VOc7VeXDJKwut8k9ebZMsz7D4VmkH9w1Yx1E/Fatg2Yrcti7H
j1sQdeLlqK1b/yQ6KWjahhw9dseuN9LERC1Nf7kN1LD+YO2d1OQCSl2kTrxz4W2c
FkTLNNwAWZxWRZ/VSTbIxtgoq8O9z/4frlGc72gLgRjjD03dScvsMLKOndqSRD8k
JdpBScPJNOCwJGK0CTuQdkopP4Ww0G0y+1OvVw5r9cJVdyLsTj+JuI+RqT09SNQX
N4TDj/HYO22/38HtImhcSoHD3yg/84lXpC+kj8fJEnD9SkpgWPBTrWuJgS4HySoz
Pl05pKaydDq2kxfNU2h1v2v+BW4/S0eSN3DG3qGy1e7Byg7kezCdZfEkfP9Wo5Fx
PDF1QRIJukGDzJygcW2QMdNpqniuuDEVMKxu8hhZjVwaNydmH7tgm8YPC8KD3IC/
kL4bWd54G8jQjhJHZOkIuBW6hGyS0mHrjC8InzBb5TYZukj6KoV1bcrgneE+lXfI
6afNX5o6ges/YpDhXelns5Nt/aBcyPB94kzpv2KKmL7FzECtcx9SnzveuDFiyIn8
YSpjgK/5oiUbvoKJCb1XB0B+CgNJMaIAEw5QVgv6vKp7YMTAPt6xRgIppNNS6sRi
og+RShk91gwovLa3kOPMyZPPK7UJSD7N5tjx4+wiLvAiNoNElvw/3VFQ8TAHkjEr
eoyyr/kzih3ODI4kx0tLhIV2KoMRPJX1Yf1/WbKSq9CPtfa7yzALZNpgQcwCuf79
138mzzfpM3EAJPN08gFbplozyRmwBIxziVF39S8alR9fhLJjU8fOFRg9L3VQVmaP
EXLlAzicEfYy6ZBYZvTM1Y2sBI928Z+xT2xoiKTHKtP+j24dRTKXjzEns/BQUaNF
4aPHFLht5oeo5A0+EzMJbDxsdikC3Uw8dUSaEVHgq9MvRycLD427xVunNQu6tFcI
SJ27woFfvU8VYS7Y1yfjgCtU20lzy4+i7765Pk5vvywrlmv5flIJPrTmTskyCQ7p
hBKsl3JXxdXP4MGoGK5UimuUDXSG/JbNJ0nhSzm4Har8A49ZIRmnsuAQVMyhdlOg
8ZMENJVxPjBvJrSflPamrKLMm47Xw2COHP4TUMgeVfnSXsQub0Qo0/UuuMybUFPH
b84MTEL1oMbTmKQvtBHeSAaE7hE0KBPkhlmMhMBIquGoKHnsF44NaPGZL9xGmmYP
BjNV54ti6+XdPngM0kQawLex57no8YPT2emGkHx72G+3LY7kncMpiQJgiJfBZyZR
0dSR3P/Xh/GB7IHaQWSAdWGW6yhG6teBCfb8oF6w2O/wuzwql/PY6S9xLo3G8Gu6
3mm0r0rALTfvSA3+qN+SRqgCGQtrlnqFcG6H7JVqe+q9wjhod4PhHNVXkqsLoDYq
ZPSy062gt2PGCh8CQjj7IisrOXQ7trzyYnJrC3BfVurG1JZMz4BU/OcDhfdKZwIB
dhvEHb0xkl5WV0olFk3swzhBj0B4my2jjMRA63DiY2Tq33/p2udbMGiW/W3CWQFZ
EZMeN+6CICa+6jcjLARuMo5z3Hx/c5NHUQP/zbVQ8Nx41WHo5TqnM7JGoyJj0axu
RH080SgQGDWOoyaEGpOqGiqmjmno7tvM9H3xh0UJFV9MnwSAAEkaP8MVc6B+366j
PZVeR4aPYYFlkXCY3T0yK8hO4uvD15Sw7TnPm37IBwA5Jy8BGxJ7+xCrsiSYOe16
WmCxhZoKdCwelBwK2qD85u6/24F9pqeArQPxswQhvZu3owFCwsSeyrQumUYxbvO0
XgQY52QODAg30OVdXQoWKBauTI7S3JNkPuSKCw+/X8AE9Pnycqdl5rrFywpoffYn
RyKlA8FOTeabSaeqLbP8/AeYEDCKBSI3apcuSAN8QCgpZXlwQkHVX/RbeWlyvpJ0
EF77IAwrGLxdEcf8lxV3yAIkHIOTEL73K1mzwaCtlajSk2WnXliVf62nwbMp9AKT
cwpzrlo6fAqeVnbQU9Eb/+RKolwe76bTMPn+7aBtFHMmkvjQkQHpiHtp52DeIrPq
HulM+hYpph5KU2WyS799OBJet3C4wGF/D3F19JtleKBUsn2fPLOComUsBuVDnc4A
NoJZv97GXMBn7QAEoV05VaGly4+7XvIUNlNP2KTnqu3tHa/NcYmfKi5qV4Ls3M0/
IGIahsI9yAUg5zT1QLdZD2l0hULWJ4pWfAVckmFnvpNKX+Cm5qcbZwTRoCyupeA3
fR169jKP9xLN/FTwfMC7C134JxTGCpqDa6MQ2WjZ2r8PQRFo1HTIf0MU7z/jl6qC
M9U+wR4lFfX/P6V1H2F4k7gxONWuTTzNwPYgFiJ8VPGe6Kn3R4lVd0JRD8U0cphq
m1Cz28yJDOZkj+Lobk9rworTGCTqbyKxFHUHBTKJxlK9vBCVD7UXm/qDONDNzqv7
MNlOlv9DItyMA8wrkAWYx45KeIvNEJqtOF737vd0AiOSNdJoRPEpl055O6ZZ+gfB
fvNbZ9t8j8ZVTWWkxqYuMaH4nhRnCrZm1wnOxx1z7L9AwV3sxToirK8z10KVRLCC
4jtxZslNxs1iDl2iptsXglOVGFcHTJH3HHD6A6eSY/uIUoc/i5EYX9cdxY92V3eY
PqWP7yuIpx6kHZjxZD7k4y1AKREQmFhQOJqYLlAi0RCz82Dm+g/M7micWxcggnhv
TruU4CSgNPTqfqmmICIXmtADTtbDxknqFqGkKoTpK5C31VwGPR7jQvwSa9VmNbNl
7rEgjMFC+zR2Tfwqjaydva7uEHC1I2py8V7uqtTJc1jpUD5Mn1yASrTzGzlMuKrG
yPWSWL6jRumPOOkc4aMUSFocSTFOCskiD9exeLlLuueY5lDe95jfaBOV88tHHDxw
f4elKdKQBxPgYXFkSdfBvhrt4ZfulkoeVn8GEE/BswkPsK+onUizpw6GBc3zJaYm
a9oOS9f2JLsH/c0+92BTfeBCMVfaWnHBz4CKpljdnpliDKl8vIy9I1CmIZF0hGJ0
1+Y2f8eJ//9uVuiniaEDqne2zbxPBfOGsS4IfjPIjV6rueGe5zYuUYAWJiPQmTUm
7d3vnELEY17JVp3tGBpRaEOtMTlnFW8Zu9Z/WhD9/YYHywhHioPSPyt6WTfHraeg
KavXY3oMXpoyz6IxUYiIyxH87eXj6hB0shnTzefBF1TJnxGmibR8JGgukT4goQJP
094LOZokeC5yy1Kyp0Vw3CFFxO/d/pYazdZXYnpU83AD8HHuxAq403RFv04QC6aC
KX8YsvWA5pmtrQZ8nw2vvW85QwnRHwE8Nrka3EGcQWwUrlxNlWujomEI+pH++Rcn
eYror4OArNOl5chdYS9gj7mYcfdZqYaEHspLc+k2gY2cv/kxKdGwG1Ld1YgYNTsz
Kr8Jwmn70L27D0m0VyuNGFk48ILsbeJS6o1DySlr6Kl5PadqOtECPYApU4uDktMY
+qwzxpxzxxOlkkb0vkHWJlz4A1wzamM6HdHeKxvhwxbfWsfL/AqaQwkUfidzs7eJ
h9P7hTw3JSfsh1ruU/1jEAvP7QGZjs69TAImU4qJu9wuntBtNZcnneKutxV5XZ9Z
LR9tfQNs4F+sx1RcFJftvTj8lDZbCA27qjdZr94VSYQ6TjqvCXKW9qsWealLZLXs
QMdG/BoXRhWBj8xOr3TMyc5GeT25jP75A17LjAujUr3BjOO+kRDoekbAndtWnn6O
PQXvYT6wtb4pzPx+u4Nuof3funNv/ITxCkyKMQFphMPUrITn50Lai3oifYOwRLvG
ovkpWMRgwNMdA794SflagRcL3+MbEKlD6e8+duCuqT8oNwEFi2XcXCaVYqBqPlpD
LjHeDR0NyEyGGGCUmam3PwLyj0W+CIp+/rk4qpCS7wAKjLfbTU13TFnWrCJJ7Vj9
F0BvwTQ3Se+XZRb0k7aQIojCr1VLoNIXqzR7GUYleYuEbXs606gOSyfZconiVGu1
dquOxZ0HcA/i5aFnqNUO+PQNPee5oriAF/laAGE+u8N4YpYThWGITHF+4Lb0O1BL
G32vrkzPQGxiV90bq128zD3PbpmSGIsHvQpNa32RpZKeFkVU0VD5fNtlasqWp3Go
5bhXoc/N4YqmLUrR17Az0WAc4ufAPl0khq+GrQojTdXW3xiYEot12aZA+kutwshd
dYFq3+C1WwAoKjM3BgJX8/Na+CeqVvSZyEnxVYQXdvhP+D7z4J5Pad/XsHCZ/Jns
l02sgyDyO4E75SjHCIDBUDRks8ktTmNXpkAnXKiyRCBELNtkQP31l9Prza/Z+v3T
W2NrjNtGLNJr5WyIgZUUk4V/8ZkmlkiJo4EfKRVQxbOm7iAu+WX287EGcee6bNiC
xpx4qM7buduu6oa7T+JKwRz8NJbg5hWpwEOo0Nfg0IHycWtFL4+jgS4U98d7I9Qi
Q69NehJDzzTH4CbiH0QhXzMCPCnjaoKOJ4aRuh0A87suKdL57Ur51AAeEvKltIil
VkH539Cm61deYHBQb2sNvd9ahM2SuXkfxb+vk08k9hcSX4cqRk+2CBEL+h8fgp3o
Q3MjP7sAkji5A8L4aFi+M68oWJQ4mlJ1Squ2H5CmgXeAiQJopQf26hLa2C18XBzU
OJIBj8xTg4FSHh/mKxirqIIKUWnAiXfI8F/2vDbxv6TgfNupCBgPTvTd/pHauD5j
1HAZ6C4AvgfWitY3B/P87W/IpeQI6Rs0kpf102OWry3vgjuQIpSjQ3dcgRF8B+XF
YXK6U7+Ysm5PuuP8YEtCR94GzUi1aGcFPqVIi6WCrsWaf9Omcql1iL1N3HCcwvvD
kH1q7w1qFzONeerY4s96p/DPKp7CL0IVZNoDrY/qCHTM8B8j87qMJgf/bVZJtei8
j5+AUMyAi+3/JOU2NdlbLAd2YwMrZVNFJcabG1fQ5i4RjwRikzmEqg8k1qlI3+qo
ne+TIX+CxRzV5LJLMw5FfrPghj2B6iVuB4hiHOlLwyY6cGvZMoHtxzMFvlRGiKpZ
WNRH8FebiMov/kLK1vtK9gn1j8nuJIaIuLNzeKBTYzhTogVafRxaQRrnogz8tbcj
rLpePJDq7tMgCeuYiQZ1DPUnB89S/Rlq4I6rSWuLPhUvDSieqxXrSfq8rwGiLXqv
GcoqcsvtK+qZI59psW69rhki+kyRk/xA7xAI/Yj0RVjCrQkHqnNHuD06jBb8Xnak
5rVQaycAz/n0li/JEo7yMhJsGVsSEwmv+gDB8cqpCYBhB37jWjulzrb8EVYwWlOQ
uH8FDXQYMIsMc3SJDmECR0HgR2lD863G7z4g7HJ9WdgGdX3k55wSyBZ0PWEZxSAx
IiE+c/KjvjUcyQxws7nN0QllmOYyMsDs9PgnKOofBl+1YllN3jq8B0Fu5VSfel/X
AINs20FUgdz0sC21UEZdOlKXIeOj89coRv/TPpOcld4cheI63hsDz7XsqedTcLkg
sHkkKb40UkbouwU+cB+MfXKGP+JwlRpab7uQhSrM2FYjrI0HvsYEdsSSDlNx+Klx
Wra/cl6jU+uQ7J1A5DlvyKZe0JzvR01aUvti9PGMhcreY4wWBLTC2tDAffe35sZ2
KsogbzUXO0u75HwYJ5XXdtzMgDg8rsv2lVAa/IpwQmNlugKjy6usHuRmbFuNN/e1
uWUrd6hc7BaXR28Jhi+GrX18pakUiPK7jKWqsIBfPzDzlJHjDKjUn43mqmGs+4x2
TOzNmWFNz7v9HbfLUD6SmMCXlgBHw5U9GSp+njE9CbNv8tviy7TlXXvoZkvgO4ug
9mOJVmymGHzyIm3kLb54ac3bnPF8MxVxYhLN3+mokezsG5VQ/uMdL7iHA/Mqo5lj
LUe5QZdDLyK0r7LdWawzJp+zrWZ+xHqNBjhyVUpPmNBcIT2j3FA34h/8mrq8RLzO
lXMxdowijaws2G8Du4C/y2ORveXoZyvPpZy3KUNeu/BfT71OfRKYVGW0/Dmf6bH1
UhmyHSOSs4Q+8SwPMDL9MBF5GRdaqfvqlmVPdiux6KlRE7X5AiR2LoUx1S/jv/vI
u5G8C23jxEDzMFkrI0iZTbOkyLQKdA7iZUq1R0M/TjqG9Mn44IF7N/S7ou/+nbmI
JwjcFjgNURVGilJBQueTqTv4K2xHLkaX27G6ybX13HWFNnbKvo3OZh6K3FIzK5uD
cghoEDpZZOGY4JN5ySTHU1P4IoxZy2LXnHHjQLBQ6cANnRV9dXuhUV5bD3Fm6Z2i
7eLXl3negWVaNveLcG/yY4MNXDhhy6ED/ScifjV9uHOeDkOE9mwWnhW9vsdGjdeT
RVTHY3ef/ET5AZmfHfaVoPu0wbPWtWHMyD+H3SebvIn2E1I6CD5/EhNUR9Qkk540
1Mj+TAL8etf40pW1cJDI99hnNZcaMM3XErDgUi3BgWZkycim5qGjLWLS1+Fdb6v4
5BLcm3mEJwRQGwMxzE+ntd0ubyKKnl55v0YKQ5ZbBpdF8J532wUKI5KKEKyIbqbi
9R45iEsIh8BsdteFW7J8KAR/grWQnlPIvURgpkUE88tC7Mr6XKwrUJ6w7SSk5YQa
wDmhkNTCyMRrEbE2QssdmH3esq7sH4G8blWe+HIifdPepVblL09llB3pQkA+WUDf
6pu7nbnM8l36yWmH5P4Ay+hqmOhPUAtoM6GijtbU6om2Yw1HJSFrPUsvzkhH2VQi
OkAmatLjJLf9W443BtksNnMk3iUkrwBJPjcHFsObndcxzVGCa2tZkAN6t3lerVOA
mEpmrkEhSeXSB65BgB6vifPHbENHoOmMiVnIiFZG7XYVeOkk1tM3QNVH2XXKQAEz
W787f+cLsjECGfWyxoe0V+sQR9a3tLryJZI2ZG+pvwSMkhi0tB/5Oz7y/CoGWzr1
mvashpVO19sKkN9ncyeXeI0OS1CHTBZn0LAG0QSeEI0yr68p2QQfmhljvY+X5xsd
HBqPwSBJg7C9vaTrhmsP0vjdbltq3DV4HaS5+JrKcO43Jv7k0KGTRwoNZPZmJchq
pUN7MBUz3A533t4W250HpUig3dre2T28PLwyGIH7hdQEsfFrBWboXCsHQj8rOmqq
LgPGhAxk4zTsV/PT+0ggDo7jale7Gv2jTPd5++kfnOTkAlUB41qK6EHiNCbLtZ2R
n7mk5auRi6c1LGCVJwttwbwaOBBskax4wYPFrBOv8Wz0/EjZQziArlQ8kMWBOAyp
AcYHiwmfC9CUleL1iIuUXqYiZ0Ul/Lt9KXOabkDc7JB+R8mgPoqDbnK0kyalGZff
gvef04NXYptu9HT2oQiqW42Du+cmShf7fZxjiIaMYUP1GsV28qOAmjK3U/ejX74O
pfkVz+uKDH90VOCtQsJjHg8Qopf19PzlkK8IRZfwRgAI7tamuvQasHfy/1KPOS2d
GIVwACR8Y88Z/EGNUUqa5zlU2ls6BgwQZ9wc8omQaqUYkaXQp7UP2z+s74Eg5Mwb
U6CG9jBQ+BY62SxNe7sSAqGOievA3kEUCVQSUeT8KxMVxKSCQlpkEFOHhy2j1o9s
Ch47HlCVH7yeywxtylaxrYWVtplnesxQvUz8Qhww1Gt0MDYoeU1NBctx9ssTxGK+
2yeOAdSWS7yMGdZdjWbfzNG4ZT/ZtvZY0puDWp3+IUV3QyeyUoPGBr9Ui/xHuRKB
7zAB5OURctijTp3C0msFGKIF4LLqi5eYQ4m25A0bVyNwq+y1h3fzX7cxjkTCdDJj
M6hu0v1MiZFrPHy4SEq7T9fSFY2f83t4UzAbz6assPwuaTkra6MHQ+aBsaD565+x
Fh9iANUvl1BBN7O3yf7OO3nW0Yv9/G20J9LPTDUsk2VRXPyR383s/R4pgVOQa9Aj
IIW3L0MBdtBnTmE5ujIr13r2Z63S9PPfaDfLP/ZC/DzF1vuUgWB+HGxGFRF9EPi4
cqba3JnVWl8eqnyPKgM20lK+ZSVCbJpR18VPemFVpFH/b3LW1vGJvCnpP5wb13Ue
t8Gz63kV13f9uySohB1CQmspbEBP52mbC5Ql+QlW2n7FJOZGlJc6lBdL/4n1wc/V
7YL5iXFgVrQto+dhu55Z0CpeNkpiEBsfiUl5TzB4Qxuw5PevWG9BHOcPQ4ZA9mRh
mpnA4uXcemYsOQX+NvpO40TbfXCzG0j/ytKISZxhOni7+amuhMZRWo5WqSo6+cHX
rmLMm+xMvRZG1tFdadzAhsiQ6oauBUN/ePexG83xVVrO8m4CnfCbNIQXCNFBSAzK
lKc/NM1JnQCxX62MwMVFAfi0sRuqgx8RRMrvEGZ3hSnNl7rM+vo2xwvUcX6nsA/T
9pwRBv44r7QHYlEggvkf6BVxK/KfWkaWgRsDyZfznMu3lBsCMAXP1OAPxoaKD0OH
oKCQkPJhMdcdgNSW3TsjlauijnJB5kShMI7x5uygegs6ADvFVl+gDOaEp2Qihn4S
jgNtHk3BnKRraQ8+6AlwWPFLVLhPf3WhylQaDg1iFSB4V0jZxRPv9jytqFDifppq
e1uXEx0WeskhlXwmNQSyiQbt299hV/0iN/KGvYrmeF324he8AlghUY3gxwDwcIiU
LZjXlSoTuo1qfw/ZwQw+5Mx20GFGX2rWrk55OF2B7tV2IDoxZrPzrclrrznDMEQM
IMQAbW6Hks3ZAopd7iz0xCi48qZM8R2zD/lzaycSQmR2W5B/188QlQQ2aiLoAc2H
jLWHkZ6jXRYQa52DiL/4g6JaO0OA4ajC4ImCpT37plmUC+8fMLi3xuTpTIVfHpnL
vow1bcfEhtMS3BO2BC0nzybQbB5tdlFv5eiLF5MBg7yrjrtulU2iDentf+qesJaO
+qsIoV2twF5XDNeVRmENB4lLBkNb63qz2hIVbge1OObADIGZkkCyKh4h77ld1rZa
OPpWy8fKuT0XeFrYjGXH7VBJCRRROQd2kz0GSRnh4hVYiFWLBlQRbrMvuH99yDKf
At/ftlpcPN+zjgOvNumUNUWcKvWyK03NkmAoBu2zq5GvVjygDRWXC9p6xtBM8QGd
SDfi2D0Mza2xk8toX0F+8OBSR7osXrV+D7P/Q4icEMyK9uhf/oll4k8h9O7tEfLe
22ikvdxAzdeE7NvpJy8INMrFOQVL3gnDkXSLTnI1oMEXRqyLTH3XLL7IkMTn5Lee
K7AFBsVkNF5llo/9of31tecnBJiyJAAYdhBJPzludxuMvgmiJoquLQzHEm4ZAWnS
BI4zGORXXmp8PFXoy6o3sKbShC+9hB/QjgoDlkYakrGAmG6dCzls7wZLAArEKCCm
QG7YphWAEINPA2OvUlxrmczvaTgcOC32LOVHJnVeZL/ZxVxWUEWeLbcwxqJFKaxM
4ShwKWHVImLcsjF7XNiB8TosnI79i5govEekXwzc3ue9aRgkf/N1taLQZc4S5d3/
ye9ALQWyWp+s+r7xAUbu0pkHVuJAMz9DqqrrVWbwV9tnjqhZrJ/I3l+3f4wCDRJC
ltDNKjC2+ytZHAxgvwCdibZ1jsADW7tgIR61Yvr5FaC539aFYN6/5oWhSZrjO5Gk
5xRk3eVRYkhQ7aQ6Ze+H2eKXWhkC4vkRyQ1Yyj6eqWX11Pj0LflZBzPUEJUWmepB
EBAZ/03q8mBVy/nx3e1D5EvDXjQlVP+iYyn+zSi8lAjaGnIn8ZaKL6R3u/qKhFxh
cMVeMMfgnH7oFTxGmTC+Bx2Uzbav+3ksgCENfROl1TS6C4QE0/mmvLr6IKiYeeNX
+VsG6/qHgtEYgVAcfhbvGQYAAJ3cwvbRsUAlnW3xWbiIPGxszWOTpQfGspgeP3Va
xMIIHVsPHIsW+RsORVvJrm3iZkq4t3H9j0SGTZhdFXz2SnuDMqviOg86Z0yLOt/n
b1s9xLbJddKPMnPHt3ep7OqYI+baJ4Bvk+PzrBDc7thYO4xqKXuqpaPIrQpt1cuX
cEzwfemFqxtqgPNqLicn0RVYPprGrO2lw9EImE6ovjWEWTeZe9iULyTYzZ4Vy1FZ
Z9zdFW4pO14K6coyWRWOD73PwrF+clJCfM4CLvUXvCcQjaKnyR7sUF27am8RLj5Q
fw7PW60DHxI/rjfSESexUhxwbSc4hAHVBZq0wo806V5O0zetly71X5NFFHPnDEz+
gfc6jdzwQOcGpgkRJDgwsW2gqREFdKHk1pPOmQSzizvusrorjC4bf8CjJff7EvzH
Ispyszqt5Xn0k3oIklI1kdTN0/LpvY2lzVYr4EEcvMdGi07ws7y7cvQfUnuEGJdn
3XhcrdvL3lwjN+NGZ184gYQdOtUMFa0kKypKYyrd12J60KrZsWe27alHG20Kw/m8
ciWPmy2rxeoE9TfkwVL9YuuqJh/+J7AgfCG7F5BIFCv+xR9r/ncv+on9hw/GHk+E
ETqo581R+cQ2z/C6XiVm1CpLGrga6ET3Kkl0BhZ0OQyFGlJLQPMGVqYlVt0BS774
+cNaLSF6TziL576ogleeruzx23+46Vc3ajlBjMzOwHBG65eJQOiM5/w5kE7ydV1V
kw032/fKCe0OFpAsh0bnGVRKipVcR3NYOYt0y9kUkowBpdgdEtgZQZhyfTjo7owA
ICV2jSFCZdvkdxVqkSQzdLOZOjA09Kmf3PgO2om8+lTENVcC3KmjthovyDIBv7me
oJ+H+nMNc7HVzsbAy9Ngpyy41rxdTPNcWuCdndrlmtpQEVLqr+P9jIHrPCfckCi0
1pTKu2jacHh9xKJndEzWlNa8kvW4VCMDF7G/hG9tMtD3hDs/EWr6wh0wr/Kjg05H
6fNx7+jqFuaM5mlMaS23o2D5v+8BSZP8a/VuibBrdu7mQj8YOUOqpC7/OHvDMb83
B2p3Ty2SoXD7IPhZ3yIT/GdSWRdwAz3byY0t+LW3acv7Oz6QoxyiHJEW9Q/YqBZI
LlLLEBup5L+3lolfMo4h1b5pqNhbavw7WzBo1jy7kzOUE9qfN1hbu7gV9fqxDJuC
aYjrfbR7ggCPHPpKri5hGIEosS7O6GUxyOCzMA1DfSv2NavgbEgpWbGpmJ1SAvUc
KPZGVmbb1VnV3Z0qLUy0sLW0rjGCIoEU0IddrpF/KOXwv2AwgEaU/Z8MBOf5q5Jw
YPf2msf01yG+stp3aGk0DUNr4vIpYxrMC7tNbQFgmHf5E+5DYVwyB1gFKmfsrefA
pjkhZ+QRuurkHYS/XUIap6GbjHsxcQjBvGccHh3hB5ddt746inLeAi6tjyo3MF2h
bthOSB2U5rYNI+oPcMCK8sBdW5RO8E6GZrXKu9GmOefrEJmiFTkMHxwpt9UWOj5q
ziKxGzISwLqMfZK7smqq6zhzHKJuLKl50Q+1Jd4ewfA+f8W7TaoJDOvZKQBA3Kvy
YerIIUj5624xK7KRaJvjP/qTKiBU6QV4qDLggd+R+A4K5n3UzRq8XV/mXKpfknMv
L7KIgUm2tG2CvcHxwLX2kZpOZLcyvg+ZLbYHvGpM90j1Ir42wrEumPEMGLGu8s6M
hWGj0AiElr3VBQgjx1wTlIuZh8UIF7aHV6TbTBxSRgehFunmdXO59+AYaDLPYNvW
fdEL3xYjzti3XzuzFVrdjJkkiZ3SZhHt6LPKiYfFII3s/5wXENUTa1htrF6meQpz
bYADx+MdNjKUPuJ1EmMgTgK5SdESXBduPIg6h8Vz7CmgtEQKVtfLOSNJQ4L5fCwX
RRnR3FgIV6L+WqUkrXlR8PuiSGUjpbXtcDvRPq9MPpoYbLw+lRR321e7Zk1DfEN8
5SGgqu6qAtJmUFOfsLx/dcNSyZe2n03IlNg5XAryM4J7/103REM/4c4SYEzBB0mO
6V7eXH1ZXxPYZUYXlLxJu8LQX2kEHWD6smqLBisOvOLXwJYXFAmqYPzWqegj/2B8
WN6pwqC4gHv/Lc9kiw9+o8eFR/FDcmty7V4SDf7Acj1XOMeD+20TOAcAlYlT//SH
E58lIZ2B0VVtIs9QPpegNZftjUnFFFwUo+Ob+Qd4MS4U+neywM6n28DGa06VFf/d
ndutJatQ6fcRy3XZT+GjBzc5I1N6e2xUOJi7HTTyncgiO1WqgYem2Z6906cLVhPU
5WFeI4HcfNweydy2hn1keKJPjESBvEn15xfizASbhtfCMTcOKnf9FtAiej8EuRSy
zIPyNELNx5S/PXs0ClOn3LMjNFIwH76QNXgr1VvKua3Nz1C88VzVFxYggdIMLAiD
GI+VHR580XdDpjHjVMDLMe6HOBSVqOOVIOi5TWxStwZZLwA8cb3W59+I9s9eWHit
XlKai5KQ+aqmNWNlWu6T3FBdT1YoYk2hteZrCVCqfV0RYRGez2kAQgZ0qCqWBU/m
RE1WrxKznEvugrJ7c31AUMZiNZQN7+OT1ZbO0UMlvIOhLktXcnRxhUyzbVG0YxFJ
xpbU22e6Z4lhpEeXaRiX88JQfWerAqP1wfJwMFR7QPGbIXmWVX2sK2JNggFntF2s
oCTM3ttAHL/BXphPYXInNlqqsfalzlffLXUjX5ZljX28ql/TZUxkl5eBQ1TTqzcz
84nXHOyXJoTxbCd/bibnkYvhcheh50B0/yADLxasxcxlYPi36owu+HW6ALBN4wqX
xkN7gjZpfU0YKNLWR3ipFhSDWjAyp5sooYeIGATmCdKtZ0A9TW8wm/wcolo9ekR6
rTL25dx00mxa61JcDdlJw511BabfQhf0SEIS44qT2wzJ6Ae1xRauWu1inZnTlfTu
F7LJ7SUQjBagdn80Yy3gUThHrnhBJrT4d261X+ewrTwOfpgGv7BFWqba6pSVlYrd
DMFxNPyxVPdjAPtUJQ4lzjAVmsx1EELCb06Z5pmkOYQLpijt4/nDIQoddSqPn/ar
3niT4X0Y89M/7YvIlyKVxAkkx3aCBvRW8znbr5JU6xG0qmZp/66S7SCg3DczpXgJ
TTcvpMFYXn/Sz+L+hGHVakQT6y/r0ZdcpUpKsObXSI/AzE9qeGxa/wNQUNpOeHSz
PXyQSeZdAf8IYTmRKDNTUKoRaG3G3uUTX+Dn2tfPPVHXzTiFfRQ5kMOnMgPD4QE9
1iigaKgLY3GeFQBGTazo1WuYWvT97/Oo0ulsIjyiwFOkyqKlBT6OCZmosIUhi8Op
KVAyW1Om+t1HSa3OqJUK9oTxPoZ1xH0mS/1olMdaaqqrmoPD2Is4qsTCpXg12Uml
AdZ0q7isi7DcJsBevREmF8N6IuXxXkxoBLNdhVF7UMtOqCHKYi0YyiogfwrEdebn
n1zvYFZ9kwDcqVvMBGRSfkxY98YOnjV4UiP/g+CXopOVWXNdhaGEe/uOCENmgPk1
MjFZogFSW6Xl+yTh3wqWURheTvinnSDBz6+kENfd8D3ONuUg74GrvdHLeuCeTpNR
GJ4q0UnCuF/Hgs0B7f4Igt211px85gAwjULX2ZyeVUx2iEN/ub5/t1zqc8fpUnkY
uSjUw443Dqx7eETIsdaSQTWiQA1VtDrThsrPE0sjDlzpaEzypOeSJmxFqicO3MOI
WtBojuYBlXyQA5oWEVbbo88i4Ig1NXP6929LcmA0LvsO4UBs02RxOxDhoYMKa0de
HA1UrCbVU+agCX1ygIt7oJrgaGY1itqW0fPQzy2DHh3UY+LROnJswizOiqoEJYbK
u7GuVWKY1bjldx6VUVAEzKOSAJl0Z5Bztu9PWu9ptDLASfzqm4uuhljwgzt07vbR
DEMAQxSZlzb80zmfGkwMkoHhax/Ggwrhkd9EWDzDfIC2TTAdz0T+5wVI5EmPNSue
mcCf2ZJcmrlw2u31BzEAYFrCnCHL7cd6l1aS+5l0hSu40eKIxmAU5jZncp/lH6k+
c/oDhzqN/zD3o9Al4Qd62fsKvQYFt6u76mmcl5b6sk3RnHo4DR7dL6jQh1J3YpCb
vRQwyXcRqnU09xZ6rjMl9l3Qrf35V4vZs3x3VW7g9xqQwO7ObI4FPDkqDEy1vxul
7x8jyFxbzIrkIxKZqq5bud2iyJC1zUAByadLl1Q2RHyVX2mqmftfQUY8I4rruWcs
+f4lzbB/ni3O0PTlOmN6Fs11kjhvHInQFnF1fajAaG3bRx4zh8l+xAoHWdAtCWBW
HJ/jPVYIzIAk76PpFO4n1lgnv2mcZGvYDk2XLivSU6kvt31oXj2HkpGMI8qduLGU
1rVS98qLA1ALPA2c61wcDF1X7ESt9TfZmwuEMsyRjiiclbCQdYAbj1iobg3y1wHg
1KSMR8o4IK5Hsl8LsQJTt8+9WulFLUqtW5m1qkM+kJdVtS7w3DhIXbWhnmUMKrCc
8aLEsZWYHW2MEFgteUlg1vjNKu7jzLa1bR3cGFSiBHwR3VFC8XFgMPKuRBBlRMGO
nFtAwcpb8dSaZE6hCsUradDS++OylEmgPiBHPD8vx3XdIAsttts+ikIBrEO7ym/B
BdZVuIxWmioMVrhahJtMM8A29I+tvgjv3dHQEG8Bj95DphVEURdrggv9ILTlYVhr
CxIilsL+iBEv/TVmtUlMEf3aGq10XAHv64DV1Vvmva3qqzyMlO67f1kwWTqasM0Y
Agb3UYyaAxz98Nih1B+5gK2f/gX1J8FXoHkqLtjuPNqMZaop2XO9Y8fun85bouzh
bDLSt8AJFAZga/PV8D0hVBkYsmYhBhQsma7OitLRUlPsr1lnjLpiITcmST/QKtWY
kMXDBXueAtIUmtdzQQ7tkbqx0gBmP+bSZ+iRIfX7Ur9Ao8kQD0t6c8UzLMUhDTV9
B8ixctxZxU2GUpR03/lYR1ui/kgRA+koDhskwMRRCL7Flw85nIPsfv6+HmO5aA4d
jhw7GfAaKTld3EocuHzBwF6/vCupZfrl6lVPKusF9lq5cljVGh4iR2znINzn69Rv
gwRKfPFLkEMy/p3kiuGX8vLje0BxRF45EpygOlmAWGnL3kNLeVwBi/m1f4TnZpMb
0gRKD2wRJ/HcWjKL8414WNy9Fi2osaydmvB0G0oVrsWhCBB8VoOrRxYhTJHx6v1f
BvauSbgbBVvrCezaGBMqtzXCXY9iuBFRZVq/RAccEsLeYiAHrLsTNQmAWjS4/MG+
LXpc4izTkgMOK7O4Zfnwgf5NEuXJBCEUcTMHaPnEYonzRCvM65glAdPgEQQsGNN6
4Z2uICyh/mkgcPgGn+ZPETK/A00MXxtvC8X7kUyyYABI/vE7omm1s6l4qLHIHjLB
fzYVqg5VDJx6NIGeBTWDSkFIgT1quRH9Jc1ZSYKYRxqozAPhUHU9pMLG81eXX7bV
fVY7T9NpSo0pw2mvgIqKSJVYRw51nfKq82hakDA6Oa7SWNiLY/nDfMqa6y5z8PeW
TUoxT7IM8Hg/fV/2ZNy8R9JMrZo0XvvG+RFAT+zYEIeEOCcZFxmUjRvsZeTMdDfO
4B6ULG6R0UtcZ+YQzI1JIk8mh/RMx6YukQaabOYmzTNh2thAgCVjCr2EtdJEIzST
u0fNpIF8wFj91ztNraghsg5zn9VLep5YcjPi7awNtoBvYyocFqLZm5BDhAxOYTZ4
iPout6nE/8ZQA1r+t9f2YpsHRXB2tt79fakQuwVb46wtmPP3WtbXKhCu8fKMbOsk
gXpfxD+aZyB5Pg3DtsXkkDUb9O0xTWXAHWJgAy7TkyASUfkl78IHhdwVt6006jur
CFUp6d7Qw9kklZ5hEQSk6SJEa2ynCd5ssRUMnvQjxys0SU5MFMF97vSKXuRnL0kj
hpgVVeWDXLWfq/L6S9u4iXT743EBVq2gHRVW/EgM9QuuoaneAdc1tlIiCBOtVD+F
sqgTWmAT6V7008rjTsLVUVLsDaOrxJpj3ymmLFyWKxt8KKIA7rs/R3SiRyVJIi1e
ushp6gM01PlctCkwWZWQPVeqZm6jYwJXjnV43UFPxs4McqR7hyrCumpGtzlNXyzE
kwa6pAHKY5lRApKp/hkt72kdSk6CIq479R7iVYWZKMa13BhzEwn9Kg6ckxhlzguA
tyDO9eXpa14p4Kp7q6/NtpIhCLbie3ikaKb6mrV7fpfyz33DPjc8k1mnV4nZA22E
CEBlvaHUrpqfuY+0ICYqp76ftYB9M79F9eZU5LDXNTr+88wWa0hfb4ojVp766IdK
l5Gp4kA8NuuyySHSLruCRWrnAypJLs2Nrym4nYSDXj5nKiOu3LlJlcnbTGGohISS
iAd80kl03rftSgreq0MSe0Zyc4KO2vTq4gZYbS3jHjYvE5ErrqdMVhYFj5TBxHgU
p0u+HFDD/HA66iy+m5O0S71EGB+7e5pvXOc0Gk4gZd0416bsr1c1jTLerZ7qN3qZ
vnVsEryyGBNxuBZaaxjMgCVjJ6DmMfXjv/5LgOCFgrG9ipr1pGI/qF0lR0gZWClM
gguUSbFF6hPW9am5Io78aNgBQXszmv7vSD3csHbYNNa/vezIIhD0hsBe7h1VcRfE
aUvewHzbMluDIelIo66VVngkELhp1yIyej62h8JrhMDh498eRFQXSi5k+gK5WcLm
qGtEAnDRWsRXp0PMHYSdEdS1HiqhiUbqkCeSPtP05ORikIvOC0Z67VXJ8Z2S9pGu
n0XrarKSMrNZnMkrLgHHJ5RzhdzGKFHzht/+hY2+92aU63RINQqBJK6PsILUnbsP
NwR87rlbyo60+Wkug9dfDzW+rovYvzxfDhhS+rYb+2H7QYPMEDfnnwhhJRBTmdgo
6JwzVyPzRbGFihV+ViUufLk2kW1SUodPPi3/E9zJcF0/jiGb8JojSSYIFINL0L21
fT3dLBkrzeGrYhFc0SHRWBJfyERq4mWXaTbOPMV5LFUBco2RkmziZgFrBRp/f0Mj
BJqfxvDPI7nq3IARWPtrLdh8JZtHAiqA8Lgk9u+q3QdldHME6LkzUCn7QuMm+lEn
MMBp/g66ZC62U+HMoS4w4b2/4LLQBQ1dYrtFXuOoGlmcSXuphesH+1xETIo3BD6q
AYNIFZkO0nk74A6QYKIaZqhL9ecVkeMFC6zLAiUvMGVUrcsd1EyQ13hzzOy+WlcE
7uv17wn0F0E1bcrgzMhNhErXuQkhcyCqiLUSYz4KYHoaNTszRi4LONzoTzNiM4Dd
zNT3qb2of+UR1iRARbQHpsZweewL/93ur6f/d1TL6UiHoXFuP6LaPXsTRcp8AaTQ
eIJQvW5/vMKZ7/orDkTj+yHODxV+dln78M8e1nsSnzatOsowyWtBCdx2XZd4C2hi
6qCdBL99S9OynB8bhxD9mit1KWn0zLZmKWzOjclgWWXI0hfMCFj/0LlOxK5gh1wa
HTDOzET5PxGrll9dUkGxX3VaeEt5cYGSY3/evv0sNuWaAJyPNW8Z0HYyMOhdGIgc
N9Sm9Vw5gTIW1yJjQxp+ai1ziGpKmCEhqV1fydcAjUGqLK+ueD/kNJPedXw23dye
fmHhofzgb1vV5q5w7m0dAqTjhi+D5AMqjk35rttIWIOPIZ5fsBH6rb5XwdAGjJrW
NvuZ9vRBTv1i++wabALHEztJtOak9DZ5thD+AEtbLaF2e3lXdZBZ+Bekv/07j/Ks
LVJM8C7oNMhofDwYeDy8BkgD56gB0rD4K2kcht9ULUD65J5uQT5nMG/u56e4Qq2s
sWxCP4ayrEPy+YJg1b+DM3p5v7ktx2YNX2NZ7M4KvpjrWve5D2mj8V4oqSHqjIcL
0JNnLZZ84qKM5PFk5Zb8u2BcyAJKKWkPubaijxowKbfMFGOnxTrO6wMazJe8osNX
A+6fzLxYoVv8nvT4S8sYwyd8+cCuakS5vahFGflVL0pa+K9BF/xYUpBwd0gQXO+x
CMPqN+pKAtqeD+tE5NRjmomAAEdp99UpPMOVm6QqUmvJPDbZLcbCCJO9dMdUYIAr
oAzHUDspLyYqXYo0F/O8+heqgn6P5oudgWP1FgzGX14swNgVCpLPM87l/RMNb3Ae
rrHCSKQcHeOqX4ytPhwoNUoYqVAuQqtPr1pRKI7EuV6wqnW41+bYFHva5LCIOEsF
CzmVFqK9A1qU7GbqWmVL1vsegHOyYDttiKF52YQWWc4fz7MfFQlbxM1Su+fLpf6w
H05U/KlMSbZIDrnqukSCl0Uq1b6/guz/dlzM26rEFgn7GdFUwIC+wmsCry52ftcF
bz98OL2Tz/VK/F3OiFOh3cpyPKFmAE00q6JmhCO4g+aq6lw45Tdi/YI0bfGd8Bo+
61Y83ibEuVta4na15Xd5nFwauTdSew2EX7Gmi9NjMCaCugvrf4bEYWPxg6ObqLRd
gHrwuI6zwiSOBQPQ1RzclRu+rqQF2DYyEr3TlABkPJWK+zVscgNfhaqgBORS/5FC
/7QM8XQ98fx9FzZfEmeOUCwjD8+0HUmFuk/wXB/bt08n5KNGA8gSs4bB0dJZrMAW
PjoNUtxbQ+jyvU7MFyhzTuB6pgmd9XLfGzdZjikDuGOuWsfdnQxSJziSeqBybRxX
FvJwJDVL4FRLudDkQ1YrmTp5U/LB1ki9V5VzWrdhufXfdQ9hO1aIuYhHl/rIrDWT
QKqHCIXeFZOYMYvWCJwZ2D2GOuFwOfzCR+DaYFMwlzUDrtV4rINKyQUSUml+jZux
YLqXtUCz5VqFlg65j3a9pueQNTJpYUB9BaHiIecAbCuDGcS3/3Ug8ysraFkLdWh7
QMboxiSdtmFsZy01mp+j95CzFjxAaLsh086H2T7iXH5LWnkhZVPmefvWyn1ckCGE
vsGb72ziNCyeJ+2Zny4du84FR6TTyhXrdS/Cy310tlq4nPvEYYjUKmfNl27z3jKn
64UmoUAsWKigHviebnAKE7SqZyG8D9qHA2XNG3HB4ldNqomqOqKvKeUWaR7AxiY4
PiSlI05T+X1S/WOsZSwznWXjp6El3h7i9cxyQVjeEBnTF2F9wzAopW4vhYQlxIMw
f236Fd2D1QAJCL2BWhFu7W+QrPK1vZXMjHMTDRiXOpwutXUsvBhQI6IJqARxdCUJ
LXMDDD4YJjZhSjwAUwUhpS9iQRWgKOGUZ/Z6tEqrLw++RdZZrFzGMTXe0fU8LoC4
e32BVgYSs1uImliQdXJXyZ1L92YgwraFvAwsS+zqfBjw96znvEzgSTh5LcGdLoOB
rXGWeGWdb+H41CAJmpMRMeYYL5mEnoxSLyUxHOlYfqmoJCrxbpcmkNV/INuTwcHt
MqTivgtlCz1IrmPztaw6t+e8f+krf2i7BREGgplL/zh825VV93X4HaSoelVmgn5e
kLn8DSOFzqwaXh0H8wt7jfc2B9HvftoB/YEU5a7Ba1LZIg83zFqIYI7/0eWxW1O9
UyCElj5Se+ZjB/PEyBXdgMHvivmzPTRCdNy+ag9KXp11A2M9lPJY3qjKTG2ajpyL
NU6dgto3DnaFrQBegz7E5/cfz1cGQOOiVw1r0/eu+adY8gXZHxctE+D9onj27DAJ
rcZpx0wAnMHpJnJcxIOQYegDroNNV+gKLvJVq+bh7gJ/hEiTRWS1ATqGVDF3zv6+
2NZg1MbQgecReYO10IrjA7uZedBYoYhtwoIHOoLS8B2BYpcBC4Hg8Oqv4HaGND3j
sKCkO7sY4bRT8Upb9lBi+9xIb860Nb5eCJgjWjhfCjmBAwUQ7QpXlGF7M5bkpXX0
KuHdKziG5RKlCc1bhmtuB6sK8GEs4NQTGVoeLnC4F3mSxzh/B8cjLUeJRyUCQQl/
Igo5V0583R8LvCr9LmadIVdFPZZf5T1HeuzI7k14CmVmbtE4c+RvBFE2tyzvxXlJ
B1hhk9dg2tjtaZ+BTytfzp2rPwPatJVvSivuG3inkrC1mKQacnfvwEH1hNrnFBQu
qnJQMKJGnuCa9N2x5/fbNgzb/SgJgz/LRZSq9M/rqq319vvNxvoxa+PwicCXHYi7
vZ978ZiSlhGqB0fQY6H6gNf8WbvXDv0SvC5qYlKX9jt53pxtMjS3oBo54v77Dj14
DtNzHKjP86lkYT61U5Wurwj9VGCNle6QZbW2709SlDBdSA3gNWnCiF9cFkn9obHf
fbMwTOhwR+5sTpwLh9mdznRbRJ0j/Nb1zNFfwpBqvjG/Nh3uZhlmtVoI7yT2fV09
iVF9EdUGTdlumdrOptXUltt7pGqYHcASi+s8dWelmM9zTmtrkexy4YP1rwdF9QB5
T2To6/ONzrwmnJRKyOn9+qqckvL2gd/+itRTLaWiDY/Ox0W2WzsmyExe+Lebh4N4
LjMjJDREzoHPFnlazjbYaXwL5NaRvA/iB40hOOSXX2x2A2yLtT9FNXMKDKXB9sVQ
KsPAaemNMoS+5/hRg+EwFXSXheibWfUNyo0Sns0ikvv9PDkb1VypuOsNVPy/sPC6
Nn8n+DG+HU8VYnby7zJevWK32p9c758Zscv49/p5e9ZQLr8AruLK6+NpHEL6Cirj
jR2TfO6CB6l6+IUTEGur45F8BjWzX6MlqoQj8XrieVfu5GnoWonv80dMUqjOpkW6
nwwZK4AHCx4cxqHVdy/jhdjlzwROXaIi7t8iiyWyVZcOcWeBtLWP8balA55C69Fi
giR9ClZw1mSMjNkq0cFPSp4YUMW4FYX+QIMnv+icOEY1o9QVlpjRS9JOpSOjfg+s
eP64Pu2THkKibzQ6JAyy7pZ0yJgbPvlM5ljzxkaflqbWf2L357cp6ihnm0ZVpidm
ASwpugKHQ5eRzhq4u9z2uxyPpLn+cUfHOsTtr3MLP0g17h4p9ONipUU8e+Umt79B
9y1JDV4fFDiGu9/i1HaB8CAlBxm5lSM0dK7XE8hsRSwBshJN6906c1RM/JE4nFYe
AP3Xnh8jwv4rMl5KWRwmu3VzVsqqgRiNi6QZZje4jHajGeu20sNUoLvNrJWzaYAD
Fz1pojIkVsH2Lurt1JdUrlxc5JwjNj/Ci/mUbrMt8AkkTKJZ6EusIx+05ES4jUNK
L4Z029su/KQPPZ++w7VHX3Kogjn7fLh6xCPgMk9NtqqUx2ANOHBt+K0pqOGY34Ia
B7YX7Orj+tiBmdROk4Vi2E1a4snKppE7CW8LleAdQR1a5IbKEwe/N0ownJJ2aKqX
2GZDhdHpcxoMhkZHZamYNiiz2TdTZhFGMruNBkZFLoqQdsLp2fLYevnGabjuYFKw
aA/jKF7eQmgkB6O/OTYESZXpxB/RAKealiQA9HQvD+qw8UaFUHgG49nja75rpCdw
W0RZCSCVs1sRbpO41vpk4yqbP6PGfT5QdrIgic3cnerXwiY3YupRdpQq1VDUoqat
WGx0c4cB0TDddAkElh0QcgJICF+zrBav4zNwKbix/1+6zw8E9mofgn2YBe0Qyo9+
DfJbiaA1H1Y9BA4IHCQXoc23kjn4qwpNDT809x3Vwn+RFYHdLX6EBnQaEwooNkMl
jQ71nd35zRp7eYUUlRn3hcXLbGp9Nl5nddGdIoS8CgCcshdXHlqmhpM4DaqEkOvH
yXnoF4avtiNChumsIpSxPWVv8D+NMu43D2ubjcXG1XGGBOOmReWRo43xsKq2zR7d
FUSVh6Y+W8DxVx87gjyPt3DIuH04yjlwFSE5dYuhwyAyhCmAQIr05p8eaz9qoBLX
uNYKeShP9VHc39AxPt16oAG7nU7NzRZz7MXNJLIwKk5uphO5E+HUBoItMiTt5Kws
5U4ecHuDWTTfgjP9OdEedTjBg/vwYulfSeAXtxJy2+vVzv0rHeOfZYPgoMjgdazu
L3twugdmeowAZWSFkqklLeOZTPpId4KCM7jxB19g3pi8MQznu0/gqPCMxy7VaE+X
Wh/5iQjVIwV2Gx3qZu+IDh5Yx8azoXZdWYqN1FHbccvWoIN5CBKDzOjxtSH8EIXY
jt8gQ2QC4gd+m1/g42ax0j8AiJQLCH6DuRutwM8mhSrzHWLHH7OcQinfyawQT5gv
Hadzg+Cli434Gao8+0mg6z62s9gHL/5LgCLigBiAAwD4w2dnoKNpAita+u0oXoH6
tsuXOe0oyS9hPAKC9qluR5hZJBpLI3XPsXpBKOiG/bO9JRLYROWZ1tUXYWNQNhpZ
H9Tb5nW9jjNKOpA24SZAbwOA6ErcS9pJAmok3QIzInT/ymYb6pgmlkUl3xjDWPk8
R1AIMvlfnOsCNc50HfR+rP6E8zG2Hwi+aDzG8SqK9s50InIO7h29/Zvc+gN+OYDu
ZgdU3LS2LHi/PXNpzaQ/e4fiOVGXEgeWT6pYca7wS+pl5fL3dtMopN4Gqqu8SMaV
dwPHgCiAzVV3IOBZRU1EJ3rwPDO4bJQbSPrQ0JSTw3Ad/cDaXGwfVRkOqX54pvYf
tAzNnBEu4ZplI50T25fOvDELkoIC0W0Fuo5o2jnrsUVfuEUfxLiR3ZLryoMIqojz
GasKV3byd79JfcOY2c3RnupG47e2g2tGkib3zDtc5m/292eqx/qtntwGrc8MxTa9
39/qd/zwD4ggyNy4ehycwyCtEdRoLWVxTvCvzYw6GNzDoT/b7e5C0arE8m+3K1Ri
iDmCjJWexYiSVQxn2O9TDej1uBKU4EesJAbCDJL3ifA0xoDul8BcynW41goP2XDe
dAmspBBd6YZ5CehzvEvCg6fmdTJa9UmWgVS+XIA9n5StnIpiWGvkNnbj9qnNcld6
XQr0reHrhUqHBdFuBi5ga0aC7aMa63N3/rRB78KuZVBii7dH0B+2JpUxy/VbAVf0
VMNfR7Evz7R4zLKBOl7wAabHuYf3gtu4AuQmxClZUnk3QDtDFc2ooPnUYroTTBNg
W02KQ9qkC86L5I9GXcMZkAIPTG33YGOMQQ0bDjn0dlBNy/OIas9HJOiYnMyVtKil
DGs+ZzM/WLfzc5UdZRBOHWFjdkQ3fxrkH1JvIycWA0wkdPL8ICBNQeWZUPr3yHXB
YwmLvw3VZVInnmgC9LPXeJX195Rmv2+Ly9M6FrmX0XZ3rOo75I4Mg/0a6Bd6yGPu
mOZieq3ZhdPea9e1HXbmPptKEXi9+V8AySJjrBBF+DxSnEXuUv7VMP7pl47SUhMk
DWppe8QT3+N7DdWw2gv800APZjeizYTta3DH/f3tDVW1jheMAjwbrz9XOY/1LUs0
5Pb9Bm5F+DQ2WcD6ito9K9d07L8cJ3wYlCwHE3QipHV6Ve23p6Ormxk4YxfFCF9w
xyVfkE7JLY0Xp5/UbLbUcZxbNb71LAXIDu78SwwjjBZISB2uIafxEqA3AsMY27qr
bKGOLCwFrcl6Ooqy2xzjwNp8JDPm4mM6cb4JFkVw8eGJomNSIWwdB2DvoKzHcAcV
HGS5msFrpm3xL1FWeYKmtUEPDm2KnpcwGTwZAkO3LqkXk8dIAkWXspY82fyKjkLv
zvBM4ws+jFMY5hcuHD0HlnDmg57C8ZLeSTEQZytIiMTCGo+CNLyBkb4nlSMO0Kh8
FssxM2FiibEArI2dPWv/EC65spsE1OVVUs3q0vUHE2m86xFwI6p0otOyEk+2PFhY
COpMo0WqoCNE2k6vXq6t4BGxh8FI9pka4qXEzXo3C+0VnVyiR4YK1ID2bCHV3cWw
p3h7aHUEzQ4203vkCKzzxDreGVv71TOj0oZNOvQmOXZGCFhdertTZc7EoMD/418p
4i8uRCA+pWmaYzX+tEnMREm1qJiEnVtWca11dL9jf+yWip5m4z9T1PZlShKnHmGi
/U/QsRKA6FZon7w5tvnpMLbEOMxkVsxmbXvx3yuuMaSBJa0B+Rt8/UX4Njxjik3S
rv4Cw8GlYepbMkBc0D1vs+31uJjjx85CeX2UBNVTg4nvcYtFyVUWxQ9Ze9ViTZXy
JDJkt9H0zCz6Kzrn2QYcWecRuypwd+UUHeqfM624g3Qk/yPoGueB3KK7rCESPIyu
9TEJ2t+nplJ/g46SnvWR5DeihmLXDy2/TAK173Eq0lA8lnvTZM3NUqSIWsrl/CSc
tkq4Vp5dzkdbZA6rrQ0ykHKizRxcdX66EZtm4mS/9BJi/QpweeGXLd16/uamtvaQ
XGgXsEoIEZ0IUvLecrg7jxmA3qhzrM0vm57QecAR6uYyd8rOGGubvJGUAc7KT1td
spudG0Itx4tCJ2zOYlXGH0mVQIBaSTtEYnBolhbwxdKSF716U+ZoH8NYfjrKq7hR
TjJZQdP8Qb2cdUF55FvzPJQWdZu84/v9MGRBMQzQuSRk2Y3j7G6dPVRITQ+HXkPO
K9iKpjfRszX6m25II8G4ni4XYEomhpoeCWX7rnhpwKavaeSzQSXHzojhqYwBYnJd
94O45my45MZEKvwrdmg1tdMOrzn7GTUm0H5o8729GjJbUlUph1cxKpXNSkoYBgUD
6vlaFTv6n/ms9+MJ8u5lSdXxycCywyXG2Bk3fWvDHzuXF3vKryIkat/IWCh2xv5l
TRJWN5LH4RFFATs8CKZ2G89JsTKxQaaFHYGLut++ite/DT1zcmTAe2OK2JgYIfNk
44jbLvSXcFO+2VAu9JpFMESiy+8JrIfVe7NlUB1vsdjczwxWBoDk9cqlTNUl6OtJ
cZ4Xn7QkbJjQdxNwKV8zCikIRJnan+tFa0NnQ4DSa/IK62DTMwA5kJ93A4MJGGAe
lQcc7o9PP//52eO0rUPpgsJZoXu3Nh9ZBCvmKvnDl0B2Wq+eLfHcZhjJoKIztFSw
oHoIxl4u7rTPSKgs/v0bDbV1S+E+gSps/tpy8HS1YBHOyNut8dwN28w1WlCUVNuR
ekiQDnABWzA8xQj2VGDdgKcoxZuTK/8/n3U9mXgfIhAfpAjTK88mQN4hdAsSRXk4
jNQDWHaUDmWqNjYH93WzbV6pkle6sX8QjQLmD9rabVUP+zEUsIzCkuoxLXjaXpvm
pspSbomgEoF3Iun02HuOOQC7cXoHHjGMkAbPrPXDXOv2iwdVGJqwVS5sFpGeICxp
jR3zZ9bN++fLHlIzpSBVb8fleHdjyVn1dMnR1bs3FIYSCPsRj+863hLZjPRSRRet
gVWvmpQnyrTYWljY9+FukiG1y6SJ0vR8OOdKivgjuem+TLXreSCx80vPsUI/WNja
XS6wrj94sz/xvBBUojijCD28rFekpn0kclWoPHJlzQs/memCI9XAUUXIP+7eltcv
BaY+f7QyDJagxnyvq2XZ/4FXkojxnPnjV4kVSdbmNxN4+z6Zk5IsAUbeCOp41Qlg
CPKpUWEjHM3YsauciABQ/Zjr6SFwWFpUNJ5pYkpj8bAfkcCnMwwfyGZfn4X7/CD1
GD1aI/PXXTtZPcaJVKpRxazGkEaLJwNQlN3PtRABpQe9lwtqL2Pxn3ryOF8Og3t6
73e7fQ6wFVVQxRFAvbMx+wIz0N7GUVBhaL3JOuJL9362ZXVzf1Kn1zuojGnJR8CI
w7mUJbjOLzYwjLTOXuhioOoCN8ksFTmh4TzEUesKAfBve2hm46z3FQIbEG4xx7dn
f3Hz/QbQqNlplmjsAvELujCnxXLISG32ZFkrA8wNfEiVg5RszhGmY4Xjbp4vjUEK
MRr5XCAUaQHp37jQ3bEJTvbwokGx7gqaxPshRQo4RGPJMW/zZnPEApmt/HCrhXvq
+WB99ghMZBvvphKAR4OpzOOPjLw8qYdilQ1UqMxXiFnwPcaUW7R5ZOxAsWfxv+CP
paQKFiflj21WSrFHq/ibMW3gpddjyXWaPuUcF2ev8Szu9+B94bEMI8utnUFrfljC
Vc26reAjVnDlgfsv7i7gdaxjhJV9OERAwzq6oMTh5QClJvkABKCHeI28yNWjSbJj
ZbhmzfbPyCQ2gRiHD58ON4Ubt65mobspjOr4XwSHYqcC14qZE1VuIYzIGrwJEEwc
QtakzyMUrT+lPfuW2WnPCQst6kg9nAxWwjA6Z7fof+JMJxn+SxbzlPHrxfl2MSp3
QzK4JLktuAAk6Edze2SwQxlilZV4g4CbWdso/fRYl/bQA7SmX2sM0aYdrl/aOJUK
SbZ5A/pM0nqOmi4p2G8FiejfOYufHUFZhTQYEax8FjPq5IHvv2tNmUqH4vQnovYZ
AW4aoNBkXMPfxankuno5gqewfsFCfsw0HgmEawnvk6q3uD9MjccsVtEfsm1rj2gs
4w697uSFC0kPxhQM1xKW/t/zIdSmLzsaSYzR8BodZEG0m2wZv9w49NhGBisfuU+j
rR8Te0Myot65Yi5E7HnG7JlT64uGuHiPGCytyM1g2yb6/pYgUUw8fJZ5FTGyE5/P
zdz2JUz6zpA7MWerSAMF2IpCgITb0p0pmsdcVkpEXTZ806M+GVgC/XNvVOOp8JkO
oZlBkRy0nrOvwIPXNEAWicyN6QX/AtWro4T5uVxWJpJ6Ks/PRnRou8Ra6GL1Phj7
7RrNWR8j2HvibWBRhRKzgkLGNoQb1iwQAhP1hubZ+HsrxBOiAL8ZsFSNUgEOxoLj
ZGo7zVZym5BSe+25UDACgF5J8H50v5CsxuIWdwAav+oFxVtQwXWZaSgmYBL/8RF9
AHH938+IxFIaHJq2HiBKj2vHG592ZMmjp4BJkd/0oLIn+SISlh3qHwgXdyx8b0E4
bM44Pt3Cx7SLqnrfeCvWBmT9wcH1bMLB55OSxUu4flqBXQNBc/jKX4AJseCjMNvc
9LKSGforWC+z7yEurr+7jSgzCrF/+XJnr5g4ixrbpOjSNBrCqg0qh59DY028EBfl
onjNZdowMhpQvIKTBRdYvw/Pph4eKljyFXZv55wLFeLAa0U3yiEJkBmJlvqhEZqE
EJFeryOn/H6UJn5O+ehOidd2bRRpBuHHapmkOvoQmtEzap03+FUxo1HwKRqWGX+X
9Xtswo2jPcXCSzUdlE9ciIlhI0gPKLNNktl+GvWFdhlRisysw5orkphhCUwRn/rB
f1rM95LiJ83JoJJPDeejVEdfndAZTUw4QAgFjV0rIMFT6IPPuiZ18p9o10IlxGBK
2/xgFESjdTK0gihhZYc3SNWDEsooyu4/HhiRARDLitfeGcrJTZl5aIoaIFKXzd3+
z98Q9Y76Q+tcMbbHgYtXHOLf2+ler0aTP/2OdnUz5xnldyXDXFYrHyorjezclk6o
Jf9KvykpZyLtNCjWiCNmyhw+rxLTEMiHVLyWHBSRyzWD1qqP6H5TfnaxcNCnhy0h
qZ8Y+MGo0mtUIM0ztbeo+zc+KxWAwFxhqchFSryUcFmk7pRjQlxhm88oIgo+IW+B
nCmgT5XpPu79vcmMV3gyogYqwH2pHroQTSmDpOJ4RXH6NuGKHSGnPvIqBaLTkBr3
mIY1tLgceNKFnAH3XTkLhM93GgZNf/CR47L04RSdg0MRLidM3LnNDXYu3J2WhixC
YRkVF4IlMWUR0uqSCzWo4xWZNOC7T/P8BbSWk653FoWOOtSeekTDMcrMGqF1Xx0o
2k8DisUHqXqA0ljQ82Htq3ChOT/tCCDf8Vc9zTqIzAvJtnewKqxceEvINkcvarPR
3dTIpqrxSwj/pqXDv1sLI8h+FASFaGRFdtpoEm0hV+Ig4RMJugXWjyCCOw/OAIFH
iKq55+7P5IQKb4ktn03GdB77De/YyaGSlEfeYA/8t4hFiAqGpaOY3TlxLG/FU1gu
U+SHmPJdfhfq8PSAZMu9kDD3FHwrjW2p3+N9xRaOH+wswqBJtX44w8d1wKyHkUim
1PZGWg7zfnLi/Ar8fqzvVzddo6+1YLfRLpc2btJ6gYRI+3rwy79IqOpIfsyjNkWE
wXgVzt5NdgDVULUGFn6B4Px0oFC7FllswxKmKXjjFaGEKFaqY+1/SnqaJc7mOVwT
ETYpAK/2uMWHr1GOTUbuUdbSE3tTi2ykh1hhl2dYESbEtUn3oSprr7VrAA7pONsq
wgV5V3B/Il0PCaKoZL17rjwYZjKLVMC2ReDd5SNgcuA1WYaZvVLpdFYUXLYnwqIC
a4PsztJCLvS3dBmNVDJ2qYQkkIpjcDuRTAzN7sEChdPvZONotDrxjQcU3/JxGo36
/1Wo0OS6VxLR6CKZdnTEL5KJNbn1jUG49wDux6n195hW2Desl85VDgwVPQbhcEXd
k2bckvCJUQxadfXrNOyyaU1+Su45reGtG/SNT2IKm/KSU+odHhniqVurlMlI0sSM
pY99M47wkXigs9K3WxxYf3BOXSB1MY0cQ1/0sVcKwNe9NXT/L195Tb0uMqe1XQgS
TIvKNbjmDCDos0nJrRMGObR5Z0t1y6h7O/kffWao1logKTACozZvdIHWJ4W3y/P9
C5LNB/uNL22Ocnme2GHj3TlQsd7KTviOYO5uiOdTRvKVIJ5CAxrtdOk92h1soDaZ
I+iqq5xekmXYniC8yvcpmti1IQFEBCxjuDkoMv3kmW/ekcCJ7N8la3WaQsKPpjU9
wFXFQvhxLavcaZgda7tqXDCaecQXKqiXiTiArDT0wHUZpgD0JPJqntyzVkP6P608
F4xHCHSpW4rUnL91K2o9IOm2S3zW8e32ViuCA/BTrQLFqizQD/mBpVT25oCuXLcr
OOldylG8Jo35O+PgJkLwZYfqLj2VYJJcqrdRyhJUfe+MxsPPdFJLMdugL0kLI84e
cs8EGAJ97int+aSaa72JcxoUFaMHimFz50Hq7egIl7WoPChgLQxtR9f4mz0xo6wI
o2Hy7hirEURTEXrZazfLF4VPVcBVLK0Aop8/rT+960CnIS2ORVrwlqviaGO4H5rS
p7JSrnAUcLv12CF0llXGeAVeFdtzRBS2wf/G71Pe5XJUYA5pGv94j+GAOmT4Jxoa
r9KZgs3bV7JQMjBcY6k5zctD0W//VihqcYI+F4f+DL/U3YTGLFEW8NDtFBpXBt9B
H7ThpYKASOxuvOi17H5Mp7itzlfMlH8z/YJbNL57m/6f/Y8w9srsj/7wKLPCgPHi
X+DxlvN7OCE6DM5V8iKsQGsW3TCDaSRwQZ7kzjzQl3dgwsekPzrur148cGTcvbz3
SKvcoT933U/QGEt4pXssYz1Y99vqpCNpD6pCRYuzSFBzFL7poQtPLHq6uhtS/Nke
OCpWgHI+EYK6zSjYyH6pOPo7ruw36GJv6RrILXuvyav3JNmVPtgt5z57AnTXmErJ
v1dCMOCqfhKD1dEH45RBaIf3TuMrfhx+kD6tZuwziW/XssI55HOzO6HNrydWMnSv
W2ns+fhHL+0fGlSnPe1zq7h/US364cufsoWFLSrF4EJK5TgihdyQmtJ7DWPSZSK0
pyym9YuOhDzFGLsgWjs5BER42z8/tq72b5QD7PUu32BmNF0bE61zhaJixkSR19V3
VA0EaxmGSZDbeufyuCn7hGR966c8C239gVuN+a10eyVtKIP5JjlREq1tvXJ85wzB
3pthb83OCJ/JDahtGXwCnhhBXtbLUzW/6tonTWSIjD2DmmLbI4+k5rDI/iSBBX7d
x94eNz9lErDW8m9vZoVI7MYo2UzaHCLYVCiAgybhDwmpPGyOXNhPyXveFST4ieI5
WNLuE2QfoPml9bXdfXYHt64+2l9u0gd4HL2SJMrwz/fm8sUQbIwIVHbfnPCpiljk
IR9p7GNRoR+zH+YQp0hZoZSPuIcoHqZxHM9rLxNsV4zkgyGSCs1fQyleWjx5CUNc
Nx7TCJz4EOjMCjtYIQUtKoztOlgUu5wgzFJpMVzl1aiNpBTKAntu07Lus+7q1mRv
noVqXRdhqmhm9zxYwbQIsrJICDZxC2wQsimjWmlf8yZngw0FQVUSFgNUWqM8RdGt
7AeSmCoW5NreS5eBkVUovzAdMcILghhHAH8fC5bYEXPi2vb/ReaDxPhFbTVlNsAX
cpP4MFU8swxiRylQQ9wZONBYOomRImyDLfVLt9K1BAlkWBGLmJbcKT2/2zqfhURb
ADDLUDcxqZPhddGEf+RdJgR+EUTtZaP2gpW9IpEQA59WX+s+b4xMwqVcMCx1BQV2
mTMUnOHt3zmPfM2Um4DU/8bv53T2a2b+ITUSFkwNC6l/PVQM4ZUZJHEBT5nQHTbU
Cny2kdzMquDIyrksYjhvCAaxzSo2cSa2QbkA2A5NDpScVcPl+XabvBZAcnDmk+pe
CoTqPvdBfCKxjL+EiWVcUsIN13KuWj07hUX3xbj+fSPr6P+ckJ7mfjGtV67jsC6D
CsWfdEcKdHJD1xp05aEcgYx7MMGScgGDLWwFK3D2Z7QSJZb6EmX9LgMDTjgK0kXw
5DsnuyD6d9uUthCluyRovRj+tzF1m/Am20u10DPfPju9K6Btz/Rf0wK6eApSN6iW
2n1MUplqwowoTx4RCHTwAZ5+wH840g8ttyIE7Am4CoXq0zXXdyreG3oECiMc2XrE
Kolj9icErStQeHF1JkH2O1YLQwVc8/DXBupSYBSxYHroU1KJaET32YuvnFshbPGR
vN2KkKXZo4jXnDe5L8qBMikjDddKW6TE0vn6XykakigljDjwARJGTfBreL2r4fBH
APQb7rO2eXq73hKeUwtZfewaroi1zg2mMY98H2ly7FtsZrs0h86HVuDie9v6GBWU
pAayP0QYwqn1bf3KLKm8tDD7MJaZQj8DUDypjlkaBe9OAQk6FuSWN1MAjdSoNeUL
uzZ7aiM15VUe/cFL3Oy/PnQsHoJDPBOxmv5m2ZtraWMKVdd5BnSDWVNczVyJO29+
DqTrMFPxq6Jkiga/sMINAJYS80vz+A3xwiIncsEZunYIRnkc3S0UCcW1ld32UNDa
GroqaSAbzhGpPun56LjF7nbdPXPJwVgNFKRcTdWspS5VUE5uZAEgWKWvB0BCIEZU
2yeIiubFJk/eFVVBIce7XBNZBHp1cuHC/xUw0Wb1j8zD0DlKYQSDltoSvvYQREDr
75wU80YOgo8W465imkiPKgKDI9hGHeCQGPlXNqO9YjrlJtGIlTv8dOfFKQjR4Ubk
uc8LVBdvJ/JWzGFgZgQgrMVLbJRjwLTLv5ZR2SkppT2JifRgNiJD76QWXgs/yVWa
Ex8AeVEi33gU4YQ7nzoWVpLEaAg1/ugsedmfvNLbUF1moga5MoCIdeiMXsaeddBs
jq+/jWctC4EzaAp7f8t72M3H3QVtOEX1vcSsLgPXCibiW4cplz5so9l2Sb0xVB1L
YjTWuReFMVwSE9i4BBAO58DbFLh10E9h00X/A5K5XynFij2bQ/L/2ILvybka9HEQ
MIIavvNaEEwZ2kciyFb5TLh+HqK+L1UC4zdFt4nzLyFBSMycd9+BnJpP1v8FgXwo
uB4KZR2p+T9csb7zEF6iQHwPXt/FTgc+6iBb87aJBV0p2tgcjVNO0YMbtuo1WMWL
EpohXcOitj8Tpq0c/UOyZyYZnwO5ybLUOp+twUM6WAC6S2jbya982cSbFewVzbcE
rg9XUyeQ2J+1RQEhVBuT+btQqZvJPw38JgbO3mTzFIom9vjQ5sdG8d1599JaMPOv
1yW/a2qbGIQUEHuIHNhPseAU7DkSLx5Qo0jk+3ZRaJJtf2sfpP97Fkz+NSc7uqA2
STv438OREoGOGjuZpU76TYaFUoRLu777eiwa4JZV6bH4n17Ya6M6GDM/1enpxNXP
KdM8iinB/VTdtCElhN94cILTkbg1fCaRgcvBCYNxKaA1juz3CYRsTcI4cs/Lz3hs
51kwwVnRh7/HxIswF32lkenD6e6jEp3dO5t++LWkkctpv9p1dsBprGwnEUa3Vidj
Cu4OLpvhCdq/7kHcByaifL+8amxrQJv1NAQHhco4+iSBjBJX3fUy18iOX4VtW1XM
RcuW3AgqWbLy4jc+y7QCTWUZZRzH0y6H5HtpqYU60NCUEGhjB8Ba872sxjJkdBJg
CPBtbOxpPmOBtfW8VxENpOCrx6bTDyuC3xDDrPJHvj+vwSZknfdWBkmGfqLtl1gv
CUlpQP2iamO969Ki42SVdmxjhzulxnnoFIpqleh1tNmUiAPjUrNbN7VWq5C97EMB
wA66aLwo9Wy/RhPwmdwndlXksjyXgwGsKy0sIyquUnfDCTE0Z5ICJSGpaPOZLQsf
0ACqJwieRnwyNmuyvJPQtHk+e+WNQdZ9I6YJoECG6TJc1ZZCRE/oM+swTZZ+cI1d
DZYRLJWTHKw9PAnS+tvk3wVhXD6Bp2uDu6/0cO1UVkhMCwrktmB7iFno2l/1s9Ps
euqxR0Hrl00jEdmla/CJ45zAIvC0o+jx6Z6pG8cJejk8UKcLKumkL44Xwc96DVvG
qMEhENkdwMdFnq9CE7CNo1+ssGSsmfKqVTOWsXkKAiVCTcKdVrVoNYRMotL+wFTD
PL9fTwG3FoIfF9071zj/89S7mgUPmvPzCi5Vafd/6IDUGOnUVHmkrzwAJbBhtYFk
K0dFTY/vuNhDlPFDjibvwaT8KTNSqgqWKVEN9EQmHDDDAOJZ5Yhir5tZXjU4mY8+
aItCpIatVfGChyHd8Wo98Tye6UFWsfVGRUXZ6zraWKSmlu9le69/gOH6XeKrytYG
pnPucqsHmRQ4SpSq4nhSr+6doRt2udq41bGZmMxADSzYY+A+GulZ9ylkUA51q+Ep
h8pJgYCUcgLn6pY2kW3LQf0D8VxrivDcpyanT6CJe+Xobix1M0C/I1NtBOU11JHv
1Npxn4T8rYE3e7gojilZrL7KYph69jvGFHG7j811zgTuKQwCVTmmXU0BHdmEBQpn
GpUjW/MQNT07bCCwdERZRCCzAC9ZfelecR+hxGkzTeWftxyMhJEqcxAFWrsIuwCU
YZiKzn7OAzs0VeIW4iyyVChBm8I8sWTHF82C7w83ngX6K7SL69H4ysJ4ygg4PXNj
jn7beYziBx0ZivS3Xa4pBOuzSC49SRS3CwyFR+yMn/4EhXsl6EGhZDPRIrYk15ma
BWvHePG/1Uz1aE0l8rG6tSVa47lTHgFNsQpeLA1GbJxKeBcX+R+rwWMklgaJJ7pf
Xt9tLe8m2f1zXxwGzlG/N7oEHtPyTMRoWTXztDFKFFSIEyUVU9tpnrPpKzKOka05
Y/JEP8MNgveMc7t+acCqkw18O1HPqncNgaIDbo2shOQMdArk4S+xJXGy546991Dy
sHVlXg4fO2SD9tkrI+FUmVBeaEC2bZcq4St9UCvYVJoUYje7/lv7LTxqsIAVKq85
lqr13A7ac5lSf4WgJZg6yDdPc39yoZGLlMktX2nHXZx20axcxeRIMB21nUucxlBM
STXZIf0WUiuYU7HSoa2pXiAeIKgqmT5fFQOBxsq4i3XyoIQvBlwGYucRkJ8YKrTs
LGg11gAKdWo81DK+LA5TyxgWWNHVVmzXfBtMf6XM5WXUzzK2yWtQVt5eq1RL0xbB
l+8NWANnlhNooY8rXh58Yt7RsbRM8WhsybkwTKAUXKJgkVEJq1hXDAi4sohuP6hY
4CxOn9VRzTn3JsHIswoRgIeKDYd/8PJnZk4Q5V9pTq82zuP3F0o9VK6Wgq95SCC9
i1ijlaIRpIEc8FVS/1eVRYx+hqI5Zm8o2giXD5bvOE2wyNCbCTmwpp0hWGjbLy0a
99ANqDNV90L1JSA0QPe2TJtUKxh7BTa9yhrUbGES3dBlS+FPiEAbZftvF4MsvkSJ
PpG2A4is+oPQsYT/yPKdaltEbJ/lZ9CzvZQf5ZIIaPwAkzkcmy4jBukkaYZoMZby
Z4euDVRbHospP4vP8/pVqj+OgtcEHAeEJAKo+r1i0nc0KZgJbQgiCqsYtoj1OO5d
hgh0V3iOnvpFmWiJISADjeb2kksOob/QtKE8QT3fkBFmAYKdfLTVcaqn+VIWxcpu
g+KHM2xgWobgReifiSABKeQHKDaaLby9Ic/my/otlu2J1S7GgPBoj2uIt+gVLQrC
b/DdcqrwBmOkpS/Mdjfyr1eKuYptH84+U7r7Ba7ZQvB0x+8v+zscYbF+IvmU70tA
4/mVjWRGSy61zEqmTAXvMZ3Iwp1ZJMUZvwDWLt9dk9ljI8x7xjBybdMpUREiB4sc
HF+8R716rlSueGVb+IM9SoUPqNGuVTqk+aDmddmgEKZp4EqiHiB8RchwKSFqqauY
Zm8qguWuxTU0hso8HrWAcGCYW+oSYL2Mq1m3A9nIClUrqks4bjusCZwEnPijFrvu
b7Yi4pOz29c5WWLmW5O6W/7ahw02iNEjDtP76pF/yTmnpqTwjW+hi1fqz0zybHFl
5cs2n4w4CTk/5YEepecYen7MRu1yquzAN5silwOwwfY9JG60h+vj93kH+rshvDEB
PDxcLc/xZaV3P+PymRrJnWT2zV9ll76ryw0ZONE41UR74iUhsjPZuTspL+VlfMr5
BTs+WhFdKMbV74fQEpMvYd7R120QzQbZvkn8pw1QXJzZlwechGruXLYfv26ifyx4
N7m64uQpJMrwcPBFSbIOm/8m8fDUGQc+Mfm1YqHUmi1YPeVNrVZCbH1HZYZFlriX
rIcOy4gZhN/dVlaid9vHcupMlOtiQMNfzl5XChk9mEkKNBnKVy80W/wV7TIM6Br/
ssVBrIx/m3jEpRKvtqlhrUBaawzFL7nMxlUsqb+WJvALv0xq2BmYXgQwYy8VLprM
ex7mqaV0jpRDlXRCpWtUoZF6Z6Mo0urWColhMlg49WDEoEJedis9YAylcQPFEEVp
z4j4OE2DYQuskldyFsTXNuMDQmteheyOdb7MMFU9qq2CPgjAA2qF4DZOOOE+fwN2
FiZaPaZv1nZA8p3qadr5YVDX+J6dfSxKtW3qKpBrsNiAW8OSmOmPtCBx9JBN80FG
8fQ0LEEgIa22kotMsKGtfP3eyGpTxWU4tiViYDM4E7jwPXFtdqhLaYYWShJ2F9Xt
ROP0iBpMyHgKgo26tRkLd4hu2YVXIp6fhfMDRLj7QbTmuL4bu/VGdzxgjbF/r5o2
AdacVXsN11InP1u0+Q5+nL3ErsrE7RdYJ6GbPZVDk1ekKnS+A5AliDS9PIxA0Ci5
5EyA5hXuFKh85GyijB3eZivX4IVgcGct0pHbZYbPqvgm25xhvD0EQbQQR/pQe5sR
GFUtgDorJeT52QnwGpBfBubxiAIJWKaVh8t++2a9oPngEr7n2BrNyha0iu3csK16
1tq5SiWf4hdJKmDv1aCXkRNXhxnqf4LWNs6a3YPlUKEXGPKoz1MiEXfUPjER3nu7
Pq9ubAAAYtCLnjldt7yej1MCC5n2TshOItfEezVh5OxArgK8JL2JvpUe1SGXKRaR
3djQ1tr8K1Hl0Q0EFFFzjXUQDOfZI+PDGg5bgHOxi8RaeFyH0ueNiZhSYsZ+0eqk
TyRc9M1CjdZqNqgiwZyGh9cK2H/v86IehwX83msyNAkRmZ7uCXsl1vOOPF2At56H
MhsiwyiaaPnWN5ESuZtzfHhjOEYvYWOxUhPXDgVFlJiMRf/DcgeXFIe9DeAKFnD6
n0mllwFwcHxTHyYEx6vlbennBHncZD5gKcXfL+eG36MuRBzF1Ctfnxc80ABzLVqu
mGtu9ybe8YnU3aMMdYEfpifxayY5WnzS7SGXZq9jLNYct3k+poitHxOzq42FB1Uy
Af0eBdB6q6jLKgOFH9zgW1og2Jx6z7/irD+dckXAVucHy8H2z7h+fHp9QP6+3DDu
ab/Y7N7KYe2zp1oWfmy1uOwOrFv9FC+xebMMcgPBhk2N1IRIJCaER95Na5D9vewF
4QmdXUtm7Z7xdom0QEkvQ8cStakjX+ikCwdx+aX9E+KMaMjagrqw3WVKH62feExY
IZRqlNvZ8tlTeDNEd6FYoINO1qfOejc0Is9wm5v8mF1TUDBXW2k22eX/09UPsd/z
pq4QdeppmePejwkuxF53uMT1ySc6wBt1qD5GWuNx0FYqOwiMvrz/p+S2hS2gQGNG
LIrJtwpr2i1S3M3kfudM1zSlI6ZrSWL3FQ4AAxf6H3RADaq9WZ7nAoEo58VohUn6
/xoZB5BUaiYz8miS+KgmHGz0YS/YhFXdbqQE8TJEkXbjgf5cgVRjS4vC/geHFoEw
I2MjVm9wfMjyCyu3RFeVtIcfzAuXfEdSoQjMqx1JmFUUsZ4NFQawAqitu4KS7WtE
ESTTp9uwbak0pJqehjRnC6IWOmnQTZJmkgcbmxJHf4/Y3eIy86lmM3OH806dvhSk
DM6Wd0CqVFySfNEtOGkmmKadT5mYH6LM/ZIyxb+9o+lsL0iWfToBaDxyzuZf/Uro
5iHijtimqP9jmDQfViqOpggLozSqG+fJo3HYg/SML1ZgZkM4q+jhQm7I5FuXMj3s
YW3lJS35Iv9KW2QHlvII88KjhmQsXAtYxqLEBAqIzWDW2+L4Zqlihg8mFg7fEWJE
2UNZekO5fK/TvO6qPv/DDp40Q765snpfveAGXt9FlUCkx4XYFYbA1LHe4dGBP9g6
fa9v/LRx+M6WbHrRzuq8tedOPJ+egcbL4FlHDoHeCWbXzMrpdNuXWHEuN+TQ2sLl
OOQUDPZbf7w0OjEjpyQGwu5NfHvXKquuAgnMwxs7aQJg0TqTypZNUevv///zqi3T
XcQYNE0i2HIE6xyKGCyUfDjtPwaOAiWhy3rd39VSv4v1Rwb41+pwqXw2OsPLmf9k
pNan5+ujY7S7QNiv/wf5IpEhv8/2MgS9GQs252r4PBS3D0DOJsiN8k7UyR3rkHfx
+5Y3NxeoRdMP8jFs/OhT+jormJUKLVVMWGr6PO8qnqb+6ITVYwp4vOEodswuKAN3
HWdXMCxtk6wdEPxxjh1H49mn8kpjF/kEITMT3+/O+H+j8xVf9Zxs0FRbCUVnI3jx
oCeR3eztrqyUxrOfX5V9RrQ5qkRRhBzPzPOU/K9Kj3Cu9CiCqHm7LU9JOiu9tFzT
U2DdD/JpS7xxbkaHwN742DIt51RHKCgO9bJIeXt5bMAB7y0ZGozDkQYO4P84erj3
zuBC3Ur6s4aVSqQzx0UjVJ5NpePYyGY9onAhOSHDhyDaYoGj327OExCpSPqhAuGH
GIwkc6lrC/PVp61jL8gNXK4CWGNeMg2jJXKFg4jVN+uBGXLq/gkHKFxnpN6WA+Fo
uMseLtfKKtDKJmtsOIC8SRHp9igt8MjPGrguAC02dGbJ2K9bwzF7CyfnTFdlGHXi
AJjh2sKnajHx/V0+6YKHwuKzFTsUt7KMPAiNhPWABYjD5Jyv0fpbEbB6BuUJZO44
QpO+UZcpzIiVCP6LdcfYLrXq57yYhGAawfQTWo6istTdX3c0Y0oD1p7bHwAT4FZa
AdJpAZipWFCibg0WTHHyc3LZsK4qbVKxbGaWyOFNZ3PHFIU6nD2Z0kXXReMmImua
AK9sVUyz6+LYq/XgAQAkckoN9COhQf7AWYnlXRPL3h4bpeLboqJHrjbuJASl9+tl
w/gEeaHIsBxuy8ME3STEyBdOE/SUgjOsp/5Q7KVml4gsBPDPg6r3XJ039IYJW8Wf
BX+zDfZiy6YYq43AevRXcVmJ2IVZDG4LCQI3wCtQqpKuxGi9Hz6atYDhfA6rp8rN
W4q2+/Gz3FgB6bMFp9llYcCmfBoEHPZ5mSwugKyTNBJzz8RC3ciTt+ltYdEeqXjI
i8jlBGDn218DwNp8CPMogBMchPw0P6vJ16rEqI7GKyjLPBxo3wnVnXvSujb5IOpl
xA+CTdGPhWFQ0RynTyWNxFw1hPOjuTjcsFkgiH2DAaRTHlNE/I+wt8Pmo8BwkG4d
g/SuEdcQYiJ15zIge7F+cHh/AZ/rbRBNRa1qQAIadnXkp4z/lOtjpkhRTomc1gd1
CoeqEoL8QzUBV0svyFWweUvWV6LuiOgtR2150R2skunNJmKy7aSOMWmf8FBNZip4
zqgwiA/DLg4MDDpfAaFBPdZZSoG8IQebb7TgwQtD5njTcPZCaZ+VDcxfZr+qoSK7
6JsGqdFCTrsrQWh1NlAEm4PvJOT28ccpqfMf7g+52SgU8aAHIY58vYf2xibicQhK
9LRt4OCqydLiMk30wOQbqQ3UUek2fQMz0bI1qug7OhbBSrwxd7kLNeJGLVtq3dP0
JRtC0w8k/dow+cJYzKao+YUz//XFvrROqJdkQwfqTZi1oaKW6z5m2suEJz0Ipiiw
vWy6/j7QH/pxpPPK79vk4uC+0CjvjADWFzBXg24+auFcd6eMb6YyvlhbTAmiH7gd
cXeJoY0ZLKU0A/6XUQVt+VamifrUyID+Gn8pnVf5Yy6h1wlmlHJxPaKHhgN+JCWG
WJk/yJ/D8Plqn62m6WjuCI1Ysn1HR+KInuag/bwwA4eKw3IjdCPxPQR1L9iVvVa6
piVKE+3RmmeU3PpKEJ5VrZuM39qRY5fBJekZ/Y8vu8TYdTDlioF10WycpHBehaJl
wUrtuEU1G3UU2pSCvkdiXevq1Eeswes1CBNAGv19xJAXgsnhaSZmdBvWqn5aGs7W
Dcuo9mK54kffnW8IuSD3/UT3XHCJMeqLkaVGIfw0a30ympLoLifA169qYeqg9I5q
QvZ58UTQKv4Lzl83Ygv2KdQxsELSLKW6WELSf/fh7kpFw8qP+2RdQzJgzkcElpuw
NOmkU7cfczOHoABlq+MxizVANNQ5RLSSg2AkGrN9H8wVBlr1sg4YzlYTXsuMDUmy
CgK2ZgRN1KwHfSryYlW6ELJVCe16YA9w7Hr/DDrb95335eDSbgqE/WQ+OV+5TC/w
sDKMeC/opujtAxp1q8L3baM5pGmRzhul/3w4aoNsUDUJUMJXgdTy+XMQSVN0dzFS
bvFPJOwKfRNYvHZVbqVxj0rTwSVD/7ekiMBTHGknvQ7IBsOYXSM5WAQISH0TCFjP
lt0erEIEUJ56c7jzB30rDzy0euIOmtIEJFC4p6e8n+3F9AbXVtSBGSKY3cbku4+y
P3KhowPdmUa4KUQMO5weWqbH1IT+/JVL0tsGNOJXjKyn5OKa7Ht3LSUsmPgdFhV4
OPAatpdUg2bvD5P+1sQHZYo7IYU1utJgoYyx6E4kjCc8RKejCIOD5U0IwQUhlywT
kupwkIojCW0T6Pf2ykR2k7dRp+eh2DXIkSQJVj3fu5t0VC14dM6P96Sku0zQ9ZQy
W7ZG5tc0vuhaRy7N/Gxe64nBOa7bu12q8xL8U4htWlU2Ushz9VC7uYqhkYzXeFDk
3e+/BgkVCZ2w4AAYPegWimbQMPJw+jV3Nscsq1zwORBP8ADh6G4I+jwnZdEUR84W
l1ARszhVyRX8Fax1KnHkC/MH8CxBc7tWMRnta59xnBkI04U4g3kZQ4c0W7l+tgzf
Tf661VpsMxcsVTmXhajHtIXhp7P1xOH+u/pYzUt/fCkLFLLpSAX6om8DSlEGMjXk
4Lkzha/xAsArrXSwkvxxTQYTQwAnCmN8zOp/w2YLbJICqAZvJROXxO5JFnpkOrRo
LvX749y9FT5rYIT0yCOaqYB2OzuooDB/mTkH7IIu6/YMh05Z3/nykdrSbqfVceK7
IMvrUevE5tHFV+zxluaHgflZ/jKj5CWeaMkQ+bh+bEGUcCyEWt/0epNLpmV5zAGF
rK1m1XQYcn9kVvpnyx5e0c+EcWHVbl2QxCr+wlXz/UaF6u2L8bBDIC6wH4p8acMQ
VTpZ4RIdYvU7FIG9/Ob4v31mAVH104OLq70ZGneD1gfaPRxx2eDrd/X13QbngcpW
kykvdA1YGZeC9s1J+g5vlpnvppiPVLbSqIv468T4pI8FYuzAhfqZg0U7R508i+wz
rzmgOVFqeW3MoOdwAPA2TAJxO6VIi1CVSqhxlM2FoDmzE3gozM96L16DnI5LDgh/
Hu3D3uYEejMT7fu+8B2ZWNsmsv4r1jwNL99Zyqt2H/0aYO60YmVP7DyjdPTcXWDl
TB1E5UexcPfi3CUF39G88C8zJuhwcz8YIcGbch9ZW7TcNQxlW9i3Dep7Kptnm2ua
0fCnuLGMQUl46+QdZyh80s1UZAHbmCY6I7zYgpL3b+UreOXtHX+G52/CRlcocdPn
W1Yqt3vZJ3RwWBXoaYri7d+KFhBstpO/m9dqePgp0tS51JunvkHAG7ZO9sIYR1L2
88CUlTdTswlOXzXAed4blzI7gmw2ubJa1T6fnDnnn7h64k6QvT2SOjVfZD/LQW5Y
qv/IHZW3jva1NX3uaUTfJGXSSyNKkXOlpjNwkz60TOX/xQ6O7Xgdgyw2OBUnXUR1
BZ7Qz8hnMbEeAjUldKvd1rs5BMUbfFAqwNOaShzYtNS5xcRytsZaQeY+0IHi6Kgq
LZm3Pz3wogwlmQ9is0punyDYiXyYlXZ3Ex8qowP/QyKPJyS25TWZ2Ib/pYpmXABh
MaYbT0A10HXqyA69GH7NPve8S1s2vusVc5MLVcUmCU6/zz/qK0e8koGUIGmJpT5M
MWMR74LG29dOm4WWaooGK5jC72d//7vlsxv7l4oFFtIU72AtngZpv831dwN3TFeL
C9pFubVpoZYQCk70IfRCHs8UHX+RC0i6sJazsqSjI3ycvYMzyF6jl5pgZrYsvpWw
8e7+h3bPj7RpesMR+m5XivI+D7+F/D98kp4+ravq5Ctaix0XLwIu0d9VmD2co2a1
FSyPiXGEpfY0xQetZtvzruCSxMCRhMhWjcExdgMZY8tlcDC89qfMPwVbKReXyQyT
4Tj1zPbhIMzHuYIe31Y1yoQK8/NH6IeKo/ydefd+LjpqpOkZMw+Fjlu9U3D0PhOp
vlOJaNIAmGQxlIE/JAvjzWzAvSM6SaWGF5GEZMx4jP7LanePzGOocm0HPCFrhWn1
tjKFgnmMBckgICqTgsiow4dh4DmZjUuDw+Db72wQMCpH5Ry67uaVfM4N3MaA6m57
UvSAILUYR57HvumtbggNJHe1t5JZr38WLMeCJtcP4hGSdAuXn0+IKMFyWkyZmXRL
eVwxV54p8Zicq6uk0y7sAg9oN3gDYQZ0FJacIw4n1x8/yws2CQBDOnPZn/YKseAD
dZmrN1VpzRzoK/vHT1ki7U0z4kSREBPJ/XDv3qouFWVRPZ/HDFQnWzMVLazPulVU
fvERo6jbCpigbopWkcP53s7z9vuLxCWUWrlSjv6InoE9Pmu9S4+HokQ0zB+4XoP7
7IZPHeshIUnqVrX+ksfiLToOAvDCY1jXdmiTkXWbkqb1RH6CLU+2LxUNswdrSkhN
k51saamhII1L6yf01ygUfXSCRhXSNNCPKigpSLtIV6d6jfa8S8EQ5dKwR0UM8Atn
tR/p+uu3MFqlJaedapQYOYZ7VClf2+4WuAvX8y9+ji3ORmIzExPtIiWi231RzEor
KBEjWGQMvIQCKuj3kd/tJEnipuKxCxtpwsXSbSRevGTIjUQrIZqOLxd0C5VeXUin
qLuevxlVH6rhh6SWllCJQ1Zo+6e1Md1ZU0GEusrlsF0XOeH7cpRFjY7LgeOR6Ofz
6UhbhRtB9KrYqdS/UkTeeQm6XH9ytZVI1OQCHv7uvqmMyEQS/3360USvrq58i2Xc
CuY5Nv2X+cmwB3nEZq8gjzLw3K0dkgu/iL+QdEb2Z3RLjikMDBgWnh6rTgOrgF1m
cV28GPF3fZlVCOnYIOa3JWoLYmTGFmXbqLUNCxTrh3x1uW1xDB4ygFcUjoC6tRAf
1UZ6ZA7chCu8phQBB7RfQDYcdl4jCIxkmlHKmYVCdH3ApH+aIpTyvIsjRLii1Y67
JCl1x8QVxuw4vs+6dND1FuhIajMNIA6hN3ubvlhtXOCC55sp1pV7I8PyUqz3gNac
otsnn21iow6+/nMOj3UHRUlJ8DNAfQNRBhJn22KAsPATzQStWVULLvJaSWRROPIk
2haapWAOj2u42upLmqPSOLgfkobchN4szlYepgWUEVF60tcrmblHwEWdN2uZG7UX
wBDy4P93kM3iPo4cBksBb+SCLyrHFxBQgRe9OudfxyGfbWOFkW5irSFu5+ubFP2p
gHda5Z2AAvTQUwF/OhooFJcvaYtSgSZ58u8JzuPH0M5L+wCwgMYDXlD75iM/T+1N
gsIa35XFqvT3+G6E2tK0RcMMSOHqSWAc5OPlgvPdfEhPZ7+9JAYFqHzdqXLBsoLT
eKlVCzco9PrCm5E+vCEIDk816Wvxn91w9jfT34JgUE+9C6XmxJ2plp94dl7Ha9TD
wSrJsPdGfE+ovBA8TmXz0j/8pPpOs1Dc2d8aoj+LyPHvj29c9dJjPZG065iULdkA
7nP/PpcMo+QT3X0pjRKUKIxii1rM+l6x7POfLrYtbMD0W7CAznrUXhwlcGdHalOR
1yUmW51123xggoVt3Sonvzt6uC60dzxpNWnYJIp5ElGj4VghqUV8uIN7BFz8lJLg
XwltDGo2CRs1g6G5PjmMcs/QqhnNpNt11lnBPei3w5fSd5N32++00S9uZSjX6rdc
XeR8So9XmasSFaeFZtDegfPu6/p8fIQpmUASxt3oiDCVb8/TM4AZaHWhhG0MuvV7
mMaZrwOf1QjxaL2ObLqWMcxQUVK35APaUGv+tZV7iLKfXdeC4O1hdOChepGx/qGG
hUgWaU9xHwEUqwOlWRpsfs5iw+5MostvDy4l+iIgX5AoJGUjF4E629lpgLLzhTXF
aVRFcFLDemLN9Xg0iHT3udQEJy8wntbFkw9UIalEO73enOH4qqXxBDwgJ9+WQDS0
QMZCU6KRzikp8bZyo5/yQxDHqQ6nDRtcyMpNmmMnWRC2H/uiR3ls6ZwHJCJpA4W1
5Ovt26MQqx3S3l6MCpsjikAi7Cl8yw0x17kgZvQeXZjguGucKl/TRXlFo/wxpYj7
NUXuNZcJ8VrMvNbQH6cMzIPKjFCyuv6AwA5BI730HFbELEZi1x3cfKajM/m6jd1W
iU98HvQs/5qXH02PHMKztHqYX7eftiln5bmu1j+0No/U2YejJgQ74tcfh90Pj33q
Pfl+sR2kfxuNPlBu2Gq64LRui9IWDTGY408zyFybGqfCaF0Gj6krBBcioWfu8cD/
BtC2GT0o3SwoWJ/JHDI2/kT+bDHJZbpdnzgixRuaTzVdwLjWgzXdbXwBdSN9DMxs
IVYO4mxOuZoGvOdJKPyOP3tGwk7kpUE9W7Ra5eOz7oFYGSHKxmOquvQAYgCq8vSM
3VE/HvEMdkiZGSmbAYyd4Oeh7uI6jTbBl/yFJcMdtw9hFabUdEZSTmEtLpn2o4Tj
nurkjLm8VqSPWGjUSs2R5z2aFPUb58RR+ZZ/uuTx6mJcRVAfuEq7H+sxyt2KSAyH
zbVQwLRiq7J0mL+lRh1zdmMnSBTA64N2hIR9JxfSfH9W0p7lLjDUdUF+2J3ZTGMV
EkbGoG4VQQv8SLo9WAy3FeeRYeRcrcfeLR/1mF7XnMGzKDQI2gbi3JuMvjxxgNg4
LksC+j716jKWoy6BXGTt2iw29GS9lxeeq+XHCoIlU/sR1ghJFlP05g2YASKea808
gCKxQ6UDh3Um0O79Fcxp+MLjd4tIerGXc9/2z2w1OmRfRzqFunwllNp20IX3Inia
TjuRQZMmScxrNPzxKcAmmsVqAMofhGw+m3746HRfMvlLQXbZekUj5d53zq1grfmZ
mQxjNvc4KvuzdRfeFlZubzs0cRO8NAQeQbKBc9yIVPdJFoF53SZ9aJAgRhMnz0yD
br3459AxbM18qqPlyWO5Vtdivh6QEzLuMwoI1BiogHqs1W7QQ7blw9UI8Crd2/q2
M/Gy6Uv7ASpXrgQuAnfCN2BFpERAP03FetE5maoGocSUHivIfiK9w+koDa0xi2Sx
27dgC+MvZXN1VwXI3X5K43Xbwkkk3AF3hJb7tsnZMvPef6y1UZ7Z14yPvCZGKo9S
o9bP7HbS5mH+U66AtLQG+8asMmMOUX3GeVulLZK9G78tivcSBFns7EJu3f0xqjdk
Ti5iUhdpzfndnA0Toz3lu/WyGw/qziEJMt7NGaz5ZpGQLmbtVJe7By/xJNsbZCha
YsvtPdplxIE5robaSHcDpfvdRNfAcORiwlqkj4MiUwyaPuKVZw9I/ZRCwq/CkTKw
pIOg1UF7HdjrHV/Qli+l245L0tYqZg2z+ppSpTlJjIh8VxFSCdMyk9X/RJMDiWcP
L2Be4RgxXuVv1oHqhq7YsTMD4FzC1AXGVBo9R1zi3ZG5VO+M1/krRdk8tvpFdDU+
sa9d0jntPlKdDZYEoiNUVXRicE2BdbrH0F0fTgpkBwnIJ6fNg51NL/Dppfca4gsb
/1rZed0r0tfPj6Pk2Ic40qMU3VHY3z2MLR9zJb/kS0uAlAtEiq6zFfWU4qDM5wjS
+PDwqbpM2CDI7Sxus5INnNtbyU3XH6yUqWe1YS2HHHgtqmhmmeO9cYZH2ECP6O7h
p+yBwpQWK5P229/7JBxPuIjy4DmTtgDK7BVrNbvtpDXb5fUUYxY74+XSjO5uuAaF
BmxqaekB/pYUYQneoPNYkeV9t0Q6xf/wkHwBrh3rrWY0YhAF4o9zLW9SBDq6JV6O
oAoQDuJW4TBQkqKIjHyMZ2ahoe4e1wkoFqjlvK6zscyoGc9NdQVAvGElyBsO8lNp
Fz84WbFYRrcU3nOBKfA2dH0NpcBEt58HXZzrYYeeN3nRz3J+6K3S3wBNKZuJBDPd
+fxuCbCOax1Vq7k+dgFI+3nSPXfNABP2LwLIi1PvHynS/Q6YuB5OZqroG/EEw2PV
wMobWBzAh4bhoqSh+hMQI9WGI5C3DZvvDkpqf4qlt4xhexuSVKNE6dHNmit6GNTZ
NnpSzNrTjThBRip6gP80WvNLCZoMfzEDL78DENaSHyGL+LBhwbfJ/UAVMLCiG0uY
5hdQpgRs+jfgORynVJGhZsKGSnDg1fhZMsTZGfwptoeDB2AeEy0BCvqr+Pztgz6R
ITHQJL9Vas9G79EO0DCdJ9Ef3ULexsLjxPfmzqbkAFiSAQd+V74F/liWz8k/4ied
/NcP6e1DhVLvfElp4Sm6L4sTlf2wiVOLCjQP8hxEJ4r5lPdy8gxRijOieJfOG9P4
Slgp/HU5Vp4+a36JLRDjUwbwmNQb99iok4Q2U+msi414j8ihd8u2X6iUIcyhcenq
68+WMraBBZsZllryNzR5bVgk8/9R4P6mPbUr7j0OcmdvuWCq5ncABTwtV8FIMTF2
Di6XXrttDwTE9B4fqQrJqHRgTSP26gLXbxo9CTyDMZk40ODmO2cFzzv4+WAaAz2y
cyLadXFkMhV79dxYgPfxKmMyIsDW1Fd7R7gR4J43IxDLzbeBOPQPVOc4gZqb64t2
aL+7LpSCNoQ8e5FNpobsyTO0EdmAjMAzRuXORWSrdMRzdmPPIPTaeCRFqmbMmyy7
5JeWeBgydx1m2TotmizHGuxNcx1tcSROm/5i7Iicmtm6FnFGtDp3GVMz+K+1Goiz
1Dq9D/iWpRRwJcYG0JW7+U94zBPaZXjuJI709cEal1XqYCTa79hdZViw/ZSlX0aj
vmOMt86mtsnlW+Mx64U//sK0PtkVJylX5Ie5+UyM6D8tHzRTc1Q/b582b0Z4lSs5
OTaCl25cDD3y3+Eaf1+Sjv00GVT3V4d6F5VpLvJMDIEwBgUYqLCNad+ph1GS3MXk
utoGsekqja/Bkbfv9WS7uLHLA+ri1Ma8kWuH9KfgIH2pEKlqJra2ONgQxrngPT4U
4I+VrdsJORWa8kLWU7FkY/7CO2VH4XwCG0xTmSVvJf7Nubk9mpOgLMEqvN+zeAds
n7sAqX4rTqOD/MUWkIWS4wbom4TJFiKByWD9569u+rUwiQMGCZm6RhP+jPA11UfI
JILGmWuGEeaQZ1GqZbePckrkXxLWIz+wZQ3zCqheSaa38m1vjmBnmIz0XOcVTe0S
VmVEarsD1BzxIBxi+v3w+tOFF5adoBh/bQ0R2pYk7ce+HJM1cBU6pPW0pORsnPw5
hAJhltTW9YN5Sk1rJFTlV3lHIwNDv8bKlrZR3W/FBxus67f9QvebC5+ybT60cZiw
Xpss3a7IdZ5hcB5uw0mlJI0UJfTx+bfQOp5liLSWktefI3fO59VRyEfx1XHiucZ6
57a+nLQnpGa0QPGks1a8MHeibq4PNE01ZU+Auzo0pZRgKsI0eaAAyJPsp2R2kOi9
xg61BiuFMcCmhFxehflHQYm1LM9fDjbY70aiCmP1Hh5E6Qi9/KK5iFMbWWr/qG1Z
6CtNwr1NiBOePISxRg5resoZA5TetLAbYKLFB1U5urwizhCcWFGR0FTOjCyEFU/h
lS8/sUNqZeKrA7usq2rWR0JSMw/amVLsgJ6NyWL3dgi20voD0yi8a3rWg4ivX6Bw
OfQQb7ifFXYMZvd4UkThuWd7zT5j71KzmxqRZDvBdXhTThTDCgNjTzvWXjdlk0yW
dX3SgUKf0l+aeO9LPfCYw2+h1KU/JT95H6krASomdr1crXVmMZV4iO3VGnwBFA/Q
9VqkZrO/1cAJ1bIqJR2umyiQz4rALQgNkfU7cwzgzZCqUAE6DBZXdm07xzgTsd4t
iOSFTb3FT4rKfR2AbuNLflClOWBSvoNFUwNTdt9XXJz0goMesJ2FTg52x5pC4hD5
vkntyUDlnMHtw27UBh+tWWxvR86iQPUpxGHIaHW8AHoFX6SyZadpW0Jj02CmDGFC
KwQRZxpIJqDRlWP07+AKG0AMce2+nVi0OGeSwSZjLZDbLwf8kSD1ygVUo6mCfmXG
Xki+PVrSEoENYYXtqfzIR8JbKjqBOgTvlh+D33yqX/+gt65VUbWloNwITVOwDC+u
0rmrQMa5fuHD5Mqf7vDZmhrh9xPxkfu3LWPQghZ5ek6BgIJ/h8tgV0hd+F2oe6jk
1TcOm8vF7JkZqjdDBpG1V1T7/qKhAP97GKLgSn3bEj8tg32hiIYDNronMuflB72N
VXJpEFPgdbwuRnSk0/ZDlPwaI50jQGEv3XelTJTopmmWGLS2OqeKyG5b0NnFtHEL
Gg2oujIbgMEc6f+fQ2ymD4+KG6UrvaloN3hUIw8ApBOfsHyuMYu+j2DcHYGgfNiQ
TxXXqUpDRI77tPo2TV0TRi2avDOwo4B5UxTL7o97/E/DhzpgwPJ63Oju1kRorpn+
uPjByKAo08CRkWRD83BFQtXDEQWUKbR1yl0n0SLOHDtKUyp7WIZrvCodIO0L1Jid
7pxLSv0P7He0b1UhO5WY3R5sVxifdCb5AvAHVFV1hJticj9TFZDMxIHQEMryqDY5
099Z7inMt4KCR3QouYBmbSTxIze0iV1ipXvlDELE62gwktiWDYf6eX4Nnd3u7Q2S
XO5p7rvk4+GHbKjNFW0utU4sL3nSCNgbLu+B00umWDWLHw7gg78Kjzm/oT+LciSF
Dn6Jf+5Vo5ayH3Pya53Q+FpK8NSc1yFu1k+KbX3lIzbu/tNQ4lwRP/F9QIty3ltw
uonsbf4H7/ip5/Pe8CMaAjE1RT3LmI4h7RhElGOhrClqB6EX8V5f81uogXO/bfR0
ZW0B6qFYksH+hPfs98B2EeTxQUPGB/FKaYBNDHNOZ51EDjAgs7Tvw/1DuSmx0/Fj
SSa1Jqji/LFkChz7j54mZCaUEfJW/i8TCvKgKzkKeiC7hDTHwHWwo1u0uDtfRkoV
svGHNCwtmXDM+yu2me2hpNqMkmQhLOrCfmsaSu5BJlYVO/UqqwGymTFKgAfpX/IR
ERL7jpTed69obacF9HPdEEO4aD/rJ9Oi5PL55WWBfcBQt4vGkBgMnf8B8roGob6o
eO4XGSf46TcpGsryrd/B3qew6OifqshondnpNnoI+rCFyd3dQXdq3mmXSxiLyEZ3
acnwnsbjRKMuFEpE+NRAIUFI59swOZaA/7EHcpCz87wuFCysh0y68MZamoyzGBzG
DcpPXFHPzqO+2gcmYtBzRegXo36sxYI80TrnxfsAjjACGpOGZk8TZ7CF7bH51I2W
+yiQEjO6vfcIpc8jvSnumD3R/RHqpL2bDPZnKG+pfYj97y1IwdUuWTvtx2SBFVUI
zd76ube+qTdGSFrxRMOZix5FHr6N+xEiatuWggOuCpTBUrt3SVp87RLIVY5wU3Ty
vV21uvIyoH6ETf/AlC1LymOH1WYQPhwku7RHfnjAFm0XtUr42X41eEPJdNKbkFxh
NrXc/g3D0OkL1Dxpi/eBNTJBfsm+3Uya3dQGukziyN/EVuxDpQ0LStQwrvwGgIno
+BnpD/UBJyVh0686SOFyKT74dBal8smWXxEEtXKReG3Tqg7khkXzy+FD9Zm/O8n/
snHXZ9iPoR/s+DfUpsbMXhSmHxaKLIC5ZlbMp6cSi9DugZvUGgCE4ZWKCmXxhajG
X2/RFn3V6cEG5rewy0tikTuOpEpRj9zgkejeNQGIbZRhnlcHzTbfGwimduNgjjgX
p8gMJ27wcCABaXpERGler0j8H02MP9vpE61B9FEdd8kJUfhpDZ5uxHgBBRI0aeg7
ggeVuPDRSp2JyY0DLMyj5Uj6BwPr4/42pN+LjLV6QPfTBcKr8E4p7eEWFWBhYq1O
EgzleuSpTljFEDsv6JzOx/9LaPx5nXR/Spkril3l36yuf9f+NYqC0tFLs/dWzSkf
Ole9yQ58/l5AKUZGvo9IJGPTVojFf7ZmQzpyrCnHuKdQP4S+M6dkqZmARfIRIGvc
rzhlQv9oRKQO5iVUPZRsqoJaThwO7kv5Ccc/cg9CNvdZ7yNryWGNPvm6AiRacyr8
scPsTbjL940aHETK5p+E83IdeaxIvmtWWb7OzRAdYZBoXEMqFjEqxEsTUtLKPxuw
rpmXsNBOeo/+dn3EajIas6MazFiHQgpCDp93rJfVaqjpzRtkH7LR+uyuBA4Ro/Fm
vitoHTM4Qe/Ra8TEcFXFBCnW6F7JULwCAuL911A63CCDk7De6xq4II5AcVwxHhd2
l3KWQ3fW9wQZGrP798IT3ioDqDCbS0dtBeIEDpNikb2ugtN8/JKxJmI1GOJoeKsu
Dkuf9k7bVmXrzUPnWQDq5kJbb9/5lc0WvianrZQfCHZQYQYOIGKAKG781yhx74st
JrwauhcVp3EhBSAZZ08KfmSpnUttI4Z5fflqerzv6Vq9JBdKq6bicDkJ9R00m+Y4
jW6IQKcHOlMM8/BHeXj570Cu3mgH6kyObhm43YRB74PK+YVgsuiX9Emp0U7MoB0B
oevGDwUL3u+ajF3Qa3WTyuJqeiLotXOhHCWYo5H4GywOqK3HbWechH8qhYckGUw6
8IgRk676Aw6g9oWuDHxaG5Rlsv+Ml0q3WUtIquj2f9xMNcydond3+YhCva9DI8pA
uHI0HsqoWT2Ni1yh0zP8D8d1UcbitJoQ1J2NeuCs/5RbEiCTMy9y3VEu9PVStJeS
BTIC/tWCvqAtHHUR9fSS5ISsSQ13txhE07UKbdwwsi6mCMKnGw9hHzg/aXvTJxrt
wp9JaQecxHMKGzF16B5iEjq6l7A0na/l7TLLccBEzEs3vkM5t9imALTB07DiykOt
t+E4c3L/2zoriMfN+3xmQiEzDrXzBWnXQRxiRgurj26ZZMkscZ6WBON4EHQlH2si
lTdRDj2IJNhhb4J7KY1kIpKhWwkj0sKom4uH35Q2hO+hHAcUseb7plGGZngMjFSS
3+Q3Y4w5aBJdkAN+YQLgsucWJPC+J7sJFstBx8SdR1leyy491o4lMSxieMy6r1JX
7oxBqHq09ZTWZinqor/FWvFBYxFjKaGYNtPyB+7oV1SOjS/6ruTIdV2oWKwNRUZd
X8CvhMTuBE8Ru2yPNfCvJcbzxRw4Zp6M6Z79i9yvpoT6va5OQ1mAyRTU65iHmEVr
/7dmlTCLCITckhk+wFaflB8SKkd3ov4rwdMhkKF1kFB4D+m2EUVlzLIagAtZcI57
BskyptDjyJ6Lp1cxfOwCwSpY5mD+Ldkd7/dessKjKDBetMMizJ8HLUBTeuzyq87N
t/K3KzBdmEk7jZUghyIO9Cui38cYm43LOVlOMuWVxfVwOkTyxHRavUT7Mlj4Vtzc
IH0KKXHJu4gJ4TEL/6JlD1VlXbCgRgn3C094wOrg2t5rxADTfetDHmScxjdTlbPi
CUu4vuSkrYaLpMoBw3yWjhFsoBTtrpUj8mgt3r1K/LKfDHvcyqL7znZ9NS49B6iy
47qqg490ARu0j7Z56KIdiH4qEhV7DVvJsBBaKOascVKQ7AD1Vtnh0+iLBB5aRYa0
ZB14X7sNMOq/S6xbUuTHjqP6Ua+QQrVoJBXYsGYVZEv6mq0TebIaOsZVhICBCiaH
vnV6qx26eOo3JXUnIvvT0l2xBfFO/yLJEhkRapT5Oh3CjO6xVV6Gz3ihtruRZB3Z
+8+gLcY5cWXoTgJLp88C9ogec6cInEtLHAte4l1UIGauY4p4nHN2I738z3IyQnS7
C2Ng/HPAjB5CVfpUW0/sh9VVzC1FMhi0UUwlZUOfBMNecJJbz68JemB4jxzgTqyJ
NLP0LswnTU5Ic371I/2tDLX4e+9/YMTAFQpT+L0jjOjT0gCSzMf0KMQPMtug1LhG
s23hU9t9NBdjjOX826O/cJQlOwt4AOLTAbmz+KzKCn9zjc7+iOE7LNzy6pkkwzx0
xiIal+ZkOxKd0pTiQCYoEghflmsv6Q18v22OdlOTTYcH/TDf8Edc1UBPoE/s+eTg
4ENE6V79cFiAArg71RR9enfa1pR6HfhrF1NukgR8diEeLXdJOjcV9WsVJFmR1XQI
oqMhRtyE3E0/BbvjjyROTixvvBYd065T/6ulgdPgaX7V0DdfpDeywIdz/ciGvtCv
EcW2beqGAKTaubgaf4T8jGvGNM/rqrdc4XO3x5Ihyol6KFU5uHFlgUenGohLwGJm
tPdWPn1hKoTyiJjNwPjOMD8tVxD0qtlmgP5oFQKvAFO1yVcODoRudpymDA1dq3G+
bH8up/3F+XW9lcTI4zG+rMOWocnrF3GMi8wepx8xtWhOTsQQ7n6IK+PZT2Z489Ae
KChH+1IkvAbBNSoN1a133pwMHzoHcoySKKmORUXEQkgZ+VgcqYOrd7pW3Tu0Nd4f
VKQSlUOpHcQYRkU/2llbL13Gpj11o5R59rDIDVDtQSAG3w/IRdA9bNLKIkGZtgcd
9OMe1LJy6CjRU3xHb0Kkt3r2uf1kElzeXwOcpKvbRCaGZsUQA6L1a9QBkGzhuTG+
fLa+nlJj6G1wG5gxacX93Cb4ZD2R15+i6qHZR/7SNQhvreV+D78/4raoVz0eIIas
isRRasfH8G4CpC3V9y+Mf607n6Vjl8yRNtH4TNADb8ZalzVpg9LkW+AgwXrLoB3d
4dEJyT2PyYLHNvLzKqISh7mmuZ4YiAJzweIDPml0u8tw7XSCuG0v0rGTe9UWWewG
doxt4we3e3GKzakxKShI06cwMA/C7rU++q+ik7aST8KOnuiShwlsrdoy7bZrx2eK
5R5QdGmT4OG7k7gbJk9GCVRy2WZ7QOIQjkIYTg9Pg4CwA4sRACZqoPJ+YDKDWwEZ
YSGCiwUTz6bi+BSDC45Olgv0Efs6oQYdirVxC8QBQvxrT47QD553FwoU3uVU7zFU
kbrk8AOboEmkDm43xR4ZB8HofjgDHzwrkbmN9hEWRlbOxzEBFaa3ICFVsN9JQL8A
IwosXkX4DJIdxuxtk1YvjB3/L0az40Oy58EkvLZOaStxlj5FFQJWyviTiOE4ttWv
jDeEI/Kj/iTISp+Gq16qxYXCjEXrQMd1XwvR0V9urWpE/Iui1M337ijb+a9cxseR
4spa9cfu9ApW98B7McwlrIMlJuSGAplIg2BBd4A1UyJKnL1plIJtTVV0qVWx02xu
RjHyVQGyispPvyAIVJ2Kumx5rfqX68+TE59V4w1IBCR5HZsacaFVzGTTFoNE/X53
ETVg/jOkRBtyNhUedoXQmj5LtALxn2/FYQMwAokbMEg4mQ9oOd31kJgf8NVah160
0+UhHK4KusMoTVsbR5Oxk4VsrJuFXTb6VHA0/gDGKgCkPeK7agf0tgOlUBstX6Xa
UDRZW9zRj/J/ajwd62/NxAxvJ88W9r8LscxgvEb7YCcZAdTL+DuAwKa7c/LWVqFk
vgjHJD8yRRYeK2PnCY3mXvhqd/SjnUp8Se4T25gReYpBdo+kAxPkvr+XIIHyGS5V
guBDJ0M0Bz7KP+NX35gXFWmA+RDkB3v3xwyAwD7lzC80fIrL4rluy3WqruiFFt7d
5RKgi9zw9876DXfCwP2TPj+7NODo0+ZVr+wt2NwSNUteuk2Ojb+8Gqyl0Njm3BuK
/gWfjAQFtiUrpYvdEY6wU7X3Z1tJ38BM0uKZsD07QCbdOBJ5weDlv4Zrx5UltF+S
gdhvN679QFktTWCy1sjSl5VbBpK9BNtOEnw85wAyRr71Nzx92AyJ5wXiPvYXKYYm
b4ra+TxN+UnaUnBIfWlepbGHGwKUd8JFliWXE7bw53cTvzaYHP4l4aHWd60924is
QXR8ujx5Pjpt+EAleRY5k5FOPZByJhwaU2tHxNXJta27NJX89utU1HoVwztzoIU2
IeCnMtdmGN+Nd/mF5RLZVKT/tnByZ8Ou8oYZ65dYL9luTy44FvpbfgYop/x0JK5R
Z4D1PiRaZ40XpA6GvqrMkax0t8MyLRS7zGgO6+qFlkCSjJfoD9wsZFhzX4+ii6g4
zl1ScJTtoP6kJ64zADqujW/J45wDhmG9lHcL/3X+4USB/4KmFEAd0lsXpB3SK81e
zEeJ9dgjcdMOJ9Q91quVGCHj50UQO6C3HVnDl3cf2Rp3EJ8OUsB4Rtly6StX9eg0
GoKYn1lzNmgbN5hE3QehWlqFGRHz9+RdNQ/EUXB4AefjNgZ4NcG+BeeJhY9ATvJn
+YpQEsZ7WmZjZNjKp5rziIjM4BqZ+b/LrTWU+CtXdnIzd6s2+yaceWIPZCwtup5L
T+vM3DeBIkS91LFgWPepyTIFXZUkvnDF6fcEBqJoiGmDcqn5euGOgdpQttWa26Ld
bBnWbJU3FBf9s+C4I4lQITqe49jiIZr31obl4ENeM4mPwgCIDWZL3XOxt2ZwTLl3
kJCLuv7NKOzTc1NdwIvOQxW+PTK5HT7yJ2OYkNsgjylO1NU7YcYp9dbt++IrAoKR
Kt2d0rDOF1bFBUTQmTLcnHBaoFrciJeb/SDuai/n0SvFkBirKfmiWHbH9HxFFqXH
TUl7AZda4ddicqfkt2/JhXvdw7a6lYz15p0bqzDD/oseD092pR3qNNaqm/4MTkl/
NAFD2DJbx6dXOhnQwr5XdJRdgXQQCcTV5STqUxy2yH/DF52nJEMqhdWqlrI9tBg7
wb0RJ9kR/9LOJG9LQ0/GJK3Vt9HoKKBqGhYwD/C/5vqe+h4oDo08JYKrFBfdNbeL
pqo7Grg0GT2ZANIpfdwcs9ZSEu4jAjypPdCEUS8fNOyXr9cNpaK7FG69vx/nyuvy
EZtwL0n6TJ2SGqvUC/X082AqCZv0Ry5M/HO3W453gu6aAiAZD1a13HIBAA8K1Ekk
cJbZEj3oCEya9AxSkTTwaBf3laxvyqvEsj+UVk96XBPzc8PaFTWbacNm8ceA2iLb
NRe9pPANJ2z3JOzYvkEEj8Iiqfg6KB0cuqkAl5nnHj4GzgOJSDRalu/qyJTJCtny
ltqhumssCTXxJJwiHYytHrm3VaxAYv8WabXVbCSeTZQ25yoqGsDG8QO39K66oilF
BG0a7NomaUk0ZWlrEf5NF1H4ee4tz2o88vA0qyxZvt9+xPg/YTA/DjtC+JN/9msN
VK97sm+bZyHxXHBCgSmgQ9UEORyt2jq+MRRggwdbQ12b4e7iGxBfgTnFgDk2OCCA
4Dl39aPubjDuWkjVtwtH7dT8bTkanL8ruftgp7VWd+FrskZOvuQOvGhqiNXohoT1
09RDWFmSyt5ThnOPHyj/WWGdnqSFMQaRDRMtaXnfV/0C7sbdU3auvbUFkmet06Nz
X5CtoOU+N7CKN1pEAaJPlT2YA4BC04J1AiIgvkYvmYkohOcDjgGqXq0nfH8xBOOp
IkBT42PR1ReJNMGqcWhS6II4RxTuQ0dhJQ0v0CijCpW7xYG72Or4RBSmHfSLIJ8O
WX3M+4KTBwOO0qczvBPQ648zvaAJNpANuI1E//qd8cXa5w97SO07jUAeyIXiot1d
H+LU3scAjwKf0pdLIssu2lN1Wn9gdkQVlBJPJhTfxnQ8Bb5EoGYoOmUBY7umgqyz
zGedp/1enjwxT4YwuPsSTWjB4V3WiRMDexRXFafRna7RLurw7P5t0Yz2uErbLsFm
8aCHRb3/Gddgv32dil8/TCmajKuvyO3yS+LlOyefQsffUpNNVl805kGywBjUlsYL
Wwd5HvDHKqUeV3fgYSKOMYRcofU+g04Gu/o879hMNXdmd7KHnNq46WsTJpmjFBVR
7sPXsHclwf7GnAZc4+VQygvCeXuNo/5XsubXudkaG8G0pTgOg0Cek+Bxb5zFEBmD
+OkBKTGGx4u422tFD7H2syupMW/9Jim4XcdLMWyrmGhBjyAOAmKf0fDdq2Q/oA6X
yNYmKh55JOLTyh6lJWgnpxpU4XCP0HlR48CbitEwzsIuM4NGOGRs5de8F5I6X0Mm
Lb2SHXj6ItCGMkl450Zvy14eGPNDugiA9P2XAs+dJP5XxNFBSy0fqIh/VWi/1636
qclSVDjx7sDufwfEmOC7gK5crgp2Otu2psleVkLyyVaXDCChkJFeXzfavVsijAuo
Zc6QNHFGp+5IFJya2gZ7/6jaYqMdITqUvUgD37YULkvOPfDJnq6s2pkuRvdW3sCc
0Jha2zKYL3MPnf+VFZeOTqOBQuD4EHjdu4sQ4Gdsko2IIodP7BEm9T7IV8PKtMdV
4Qo2L4qFTR7F8NT0AqE+Q/wrnPrwylf06XC13XH2z8ku2IvdoBm36eW8jxGBdE9W
cutpDsHDBbMnSt+n2mqYMaaFD6JZ/h4HOO87By01geVEETCmd/AJFIMaynAMfpKd
3dAC5nSJdgzx2+kqVMpeehDNsZmKb7SbABWnNnv7w36oB+AScJB88byhDkwwut/+
giRYtrI9OMmWHSAaAiuKwkLLVfcAijm4AGMLDyssryeYEN4nrmfCrfjDjSUc/UZP
B27h0iElIqDffL/9eaUYY0Sej+XTc1FsuvekigFqujjrx6C34VLkk7ci88mzKoJJ
ofqJgTMRXBx+Nso4ZCK6MZR5tf3aeogcttz/wYmkKSNXgWfcFAtJFOmPeceN9gs0
/HzDKJ70snCMdZ3Gwnbt8SLpzB+gnQ5TRYqDsbk9v408ivw/DtfztNgw4O45G7ym
nE27LMhVSl2x8gcVGzUC2JhSaVxE6YUaCfWUZ8j+c6Hbo0+ZZ3LysqRcx3rAYj5Q
dlk658Ciu9GhBIVbbIHORKlz2CKbszoh/hqBsswisaB66NKiMfM5UVdXNbnIiy5/
8qHGhDJvfSgBAn8ruwUWy8uApD19Knd+tO2zBiMLCpjTvgUd8AAeFtf0Wwoyiipr
3e0Une/EmQp3wRFnFVnBH8gzLw4CD3eMgDbsBxcvurWiuItfGJ1mtEW1dhjcTqHo
k1EZZNXFD82N4ggyZCR5gO2zE1GksESTI44jJOsr2rVAZkNZp0V0WNazEzV9dgjc
9Ro5K535kiceKcbCtlTgU+Dt0Vkbeo69oTpacVCIfIojP0F04uiPlpKfm04orqVY
dDhy8DeWrfWnbAVLa2/7/Hlx99S+NMJG6FEh9Smugw7l2fzU8RrbnDmAghBqANVJ
4S8Wt7CiUvYg0PV7jEEXof8nQxpdv2LwzUEuXK5vHwC8x4YcIDvtAdYqZjQLuirl
bTezreM5DBDv1k8TJ0AU2TDAZkKhvY1s4FubWkAQL8t00FVw56l6OGL6Gn+IoKC7
XL+LpR4I8wCgSYwBWr2AkeJ8QXfxHY1YqUv10VGEK5wTVNQt9T5Hp7tYa6OZNrk4
/L8AaHASRwmex/Yr45jYoqQ1UPDYt1smxMvOSGOpRXsd4aqcGbXfb25ObBhpjCy1
FhUdMhYEQXYHSA0wxojUrhNRvd56QeUzTTQDTF8JNoCqLzXLMBNjxWBxc/d+/yNB
1AclF4X4qc73laADwdtVUCSRD2Q8m36tzAmERpsp0Hx8lTb3+Dur69vld+EDeSDc
IeyLnxJHtsu40H+oaoU7q5ZdjFS0oxTzw/YhlsJHiBMGnzipvvj5cMTgt0Qnqn7b
YM8wghY/owwR64c/cdKgb+H8lvLEHVlmyW6omnpGmbj2X9unAvJPX1jXWk5rMILp
zfMTm5ayf30y05ZMqcNOe3AtUDgnncW9pL/Go9Mmcf6zKpXjZjCFg/zrARVXlyl2
PLTaMjTboZ/UDeX9NlQJo8od24lyAHaSXAN4oPftytU9sSlKayVodvB5H83b0+p7
NIJfi8UsJHodr35AOPcAhCJjHh+QqIO8pmQ/ycLgq7qm9lQ52VfHTldfC2WbgkLB
1sZMKZQ5PI6J4NKjyACgnEZEchUJ7lySMYefjjXfF3WFI4gYdmh55ZYU6M90exDs
q3O4ddam/5YmLuu3BBFN2vH4oHRcV1yEJae8UBe7UMsQw59ia7pL9nzrCODegNkj
LYc0f7ib64T8evudkujEvYUZT0sXfHTpY50iOK0yhVX0xd4BSWqPIkCK7fqrOQ2U
Q8i5+Zx6a7U+2ydQX3B7Nr01w3NF6knNiHAGl5QYxRpOoCDcR+rq/ZPLO664cCtZ
NilprwHqw+1PoTbKkoh89Bl5Y44G4EO5bl4tYtX5Kix7L+Jn6WfSG9Fuqasz6pbl
k2AVQDiUzrND/+aDykaJKhYFulusKikdma24bv7ZmJj5Gmf6hYsoHseYpdPLkXNu
k0iwxsAsyje41a/IHDf13Su0278HtsMWdRkWT3W/6XaJMRPEEZf+9JxURqkFCI+R
wsmIq7GuCWYBQsQcQkG7r3ZVpdYgjMnUS8TIvNaSdDQKijWqkJg2ealvMRVwIWZS
MFHs8pA2oyrHtCbPfxO0fNAVcyrkYlNb5LvvtIBg7qo064IvKV6rzltX+QMuISrT
5hl8r625ZoahawRGlfHa9NdPzjQuEWsylzABnLJp3JSrc8al3AqdkQIvfISqZeQN
3rFQ7ary34AcrJ6f3i/mLs627AkiJfOs1X4IF9O0EDVVpj4+4zVJW9FUFNXdyPyy
zDHW15xr9B4JfHojKNiGFQiK3SDNSQDEeZvadk7FZCVpAd3S6W1/MbrVK201DJLM
zHJA7df3V17nIbHgDALtrEQpXxkY1TWkcPxWJqqv9b9ZhEDL6kSmJW6TxNHw4/+G
iHQoLBW2stqgG7Jk1udkXl/yJW2K59AXxw7kGwoPKA/5MAyvN9HZvq+xbcSmpxj5
Ky50e+rnWTjkKKnzlm87UsLqNKD8Ehdt4CpcmFENb3YH80ryn5Y2wa1sLE0fyLoz
g7Dz9EYuuLRwu0kD1LzxXfz0R5j6Xkr9sPLEube4CTl2Dl3685zv3ghJCEMNzFPQ
gwYLFPo3JNSgbaoDw5/Nrf2gCcYupBVDMORzit9j9iG9alHTMY2ZXDvI3+ZCPzo0
aMq3GrNUiIqq3YEkQ4HpHhuTKcVlb0Y8UykORPfv2E8xBh1CKR84quSyskTa7XgP
Li14iR60VYtT/XQSs01IjEEvZr2jdMpCbnWgUP7UN1E4iOEqIFzSSI4mQxwsj546
MSEeZsQmRuMnGCFLEVAtuNQqCsSyuwZXz1ekAtUiJXp1kY1LrrY4g1uvziX9HAEu
KuUF4Es/TQCBIdIxSvBB/pHUp2/SpRpupvwimcWFe5AS6xg/FKhfenLEoTULKbcr
4/1arxGEe+GWL6HPQYVSSVHuEq1oQvKC9BxNBkFBXDHEC8rKn1pe2yIrl4DxIkMZ
48AtD7e3kAD61Jn9jEqssO3dhVFZNQpsfISteLG7nj0p1ebeBXD01z7n+KW8oxl0
d7zzRGqJdypASfqrJ46GMskEGvXTxzl6+DEZtWsUbZSHplqZD6+ucznOxcLjshaa
jH1pVYFm7bs/BK6VRKWoVTkyO1fUZmqQq2K2KtAc4yVjqKca8AA4Gx+LrqxyOdLw
0nT6d+v0L8VZU0BvxmN370uMZZGzmSgsDhQ3X6KsEgDYarYxxJH43k1N9pG8acxX
rgXe3U6gq82ndDkNgXpSm0kTLa6b9cWe8jKsfEmR4ZwW4rkDloTjdljoID2rBY1C
o5qkdoXuueep2wDqalCEJ/yaHjNZ5mvRlWXGPlheyNwM8M0bmbhF2aKDc9c5leKC
CF8Ckr11rm99Rz5MEIJOzDY3tQj9Ht7IUmjlO//03jFQUAduvSaSjOBhWEv8t5Ld
pW6OgErUN2LUKBwCmJqjf5TgzJW7l9nca3gT+jAlVKI8D9WCJ4OIXacqR/F0FOEz
N75genuPbHrQ4uGF3zE3bAHh4xhH6pF/qUYpVWESJg6lv/n2qfEqL/LPeHnPuX25
8qNaOJimlaTV0rdhvQ0N3tz5FjjuzCzQsmRdRzNC7W9bSGmraM2XMu9Fd6wwjJbQ
sj+ah3vO4kbo/zBOUBrVG2OkW4IqxesGjYUDlOdiKV46SGe7vSWQgEmesjH/pmnJ
gYScEqZ5quWiPRpGqr8F7s539mIN+GuDmoTqi6snnqq4Lm/V/VbnfF/m7XmN7Ror
n8NkQuySR+hgHAuu+9oY/t3l3C99kTuM+Jb4GVa7xq1jYzWRtTpyrficU02r0OLL
4RTBggQKLV8DmdrFaYYeZDuxe005KWzCPwSwVmsQzAgoHKAfCxByEvEqYzkevii1
BG27uyVJXLJdY8QwVFwxPfb03R5GfV9LMxDcPlYWS/vywyJAmD38eQ8UKDa9fJEp
2JTf6CIo3r/7bwx0lC8wh2VnJeVXDxz02gV6hFiC/ydY+rJ42Jl2m5oGjon5Cr4h
SM6Uo+5ua/iZWVVoNf+A2nArKwXMh9ptC30hziJ6iD+tpg63436gN7m+VainVxBz
2vSa8jjUCr0hqBP95XyY+1P3tgdRWBIjWo1G83ZTJiNjwrjlxfRpjG6sJqg6OI9n
vRtZwmJwzl526wKcHcAbJCznVsGj2bFEEPpPt1mMFD59CFDfwZTNUdcYOARC4oTE
/Ugzw4Dq4oAyacbykMcPyP+bM3BN/4JTeyYvGnVYlFv7FjIBMAQPPS2wt/n6IcVn
XpwW0WgqE2indsoNolOZjmrqjyECLEJnpCV4ELsNOovaA8frpow+4fAYHyklCMv+
F83jK5NFQrRihAUccBKaASwAIO9UOuwO878gPBRCadh7RohEHsdbb35vTAOEnBF1
2AFntYYvnuxxFMdmnI3n3WK8O5wcAX+OI4s1PNJprVgVImds1At5rQxsjyvcvcg6
FAhCdigkHnVsvm3x7k5UNl76SxzheuPp97tFRAx/vTAKTfjjX3Q53KsucoZ+jZYI
bYFxzugYFaAyhlpkjCGzAXI7hyv25CMhWX//l8BbKx9hqjNZ93MsUmiPohNqa0Gm
w5kv28XO1CKlCjOXcAAg7hyOGwz8jP+uEyeSa5cShe/L/rpsip+mH/7lkOQWt+4U
xcPLIY40QAQnkpLgVceqiTUZFFV/g9Jxk67AVeG6t+o4s3kH+mgm86XikeQGMqol
U1rHXNOVO4BHx4vqG9o9BwcIkj1QcHxWiriOAMvCuuwcZHgxFkb92bfwpWv2xfFE
ibMydcGEfLL9weenIJESxaNbvCRE0KS1OjgN6ppQCfnrHsqle/urcdNRt9F3HHHb
6lhutb9UJL9OOneZ/Ww6L6KkUzUmdIbSdPG6TMItqrPg+iM0uiMVcZIFoEBeiGk6
XBrHBSNU1QfOzezXkIt5Pr5hQOMpZQhelcigqa+b2CsEqwUCQtfhD9xxyaFRMCYP
WhEaOa06ZGyV1yjCD4Qy9LpmIwOyT0j91PgTbWr2NI9VrSkxpNPd1myGx6NE92Gs
MHK8k9m4jDKGcW/0TGO9cRkLeYWHDs64qKYfd/rkt50lGjJw/DflIVU1OKBcx93L
AuGRv9EF7wUnZf8P72axQ5CNlpznz/NcLuyHTEA1Gi45fmH511aAUejwv/FSLiuC
WImNkBWhDZl2lJOH2zEVK9YBfwT0Z4zcUyMaKybjAoFh5iNYM62LNwxMyLFPb7oD
xb4HkfMUrumMT4gTj6E0d6L9ofzHBgHbxv4Nkb6u4ATKcLS1jZjYiDwTxtmyDWlG
TT8/DzG8XCRW67emhGxnHB/Ij02Wam3AgKNfbbAnl5AsF07siCFdZzHWcwb3Dwen
yNRSqbcRZEuQqOblrB19JRrh31lj4Azp55nDyBc7mpAV2GTl8DYNXQdKGVBuLc0A
uUYIlsuZl/Bk6ZTxAWw7d6hQcPYLD0cbQEg5xvTEN2ZDIjOpginU771B068PMMpu
3kGY4nKv3oZ58qW68+9ayQLdKAWtYQPbnvQw0RBRmHatzdU+O+TdrE1t4tSQn6bA
Ck7b5yV0YKSW2fdgmQexR01F4jGvebQF+mMYFjlm9PoN6cveBLhsJAt8qfjy0yS3
TGepSu3N3XfQVSHoaEhtzPzUGAjnNVj2eDAUqh8nasK1NmzCu7ozjbmW2mRTNuqR
1Qq4JVAlw2vDVnead+rQEcJxH1w5euGdSZlyfyl0GtfAIx0zXII/56GvJplzLfNP
MQAmKWXJxFOOLiUYcJ0LxLny2hYg77c8rzuyd2cM93d1r96gUDjUnezY74EZWA0X
yYwaFcxJ5g4JvTb3W6LPO71GHWKfULuxwdPT0/JCKT8OE75sVCl4MCKYAc3nA8S1
47zJcJ6HoOp4B+owXOT6u7ZZWrfLythgF0nVXSdIDm/VDU+DijVemFcClQsO7fRE
jyPWRcEJbhrh3WX6KsslMv0wljx4In39rZArfg7Jxe1HFBVyxRbnq3LmgyrhuzEb
cEjpu8seJAk+t29lege3agOBsnrTS8lvJCI/tul6BC9cQhiQAY6oq0F0RhEPog9n
NGvPezkrTIRierhZ7yl7vqq5jNU+1edcpl1Cp9eQPfn3iDxpA/E0MjJQBndx1sZt
LcumUgXByXbamk/AzHnso9Dgv5sUJl0jYrrPenZhnJgKvrGOf9gTgqXrEEEWPFmQ
SmYQrnt6pFWxLI38cmRgK1to/TUh4dH1Z722zHgI4qPlIcB/Og/vqkoQ8War8zO8
j2v3qoQdqa4IrSN+GxTUUWS5/Fg9FRH2tOBCMZUqAvL4W7R/LIjxMsxybqGRA+Q/
1ZenR4FWP7M6Z/OpEAIylQZZIpevJEWnPZMJ3TpFL/b1QxDKx+2lrdZq/gxxfaIr
tB7UfyYOK6vDT2WvrjCfdKNgWUXN1IWoz2aW+wzoepLUn6GAr6KuzAcPxdKsW61c
XsfyjlVg+AstvXH8ggFW5RwOIf1qbWgYCakykNX4bmQf4aFC3u1P10ShsRW++PY/
QNtpJwOSr9Gml4TH6TPobJQpzHpNqZUiV/E0L133UbQ/m72M7TFzA+GEWS8hsxNI
883Y53/squzfbc+qfzi1fPDPAMGx0YVDn5KDI/MBhiPuhxNuqHC8ZbUL1YYyHMDS
ObNsXmP8PFuG3nepA8bAOeOgcelJlUMQSwc+SN6FbMGWawzOUsXDud/w0OE1MKJI
eRIRWUisUEfSuYyEyTCPwjynpMGIceS4Nk2NEdDXrEqXfdG3qut3ohCwFD3tT45G
dD+aWRNQ8/w3jRR2OtdRPS1GNkHQ1z8NCk/LOhYlMYwdUEp7EpzjOIZQq5Pv2PQR
fXWMxXzxWpnMFIUc94Nlabpp7D3nCZHeAFVklNAa5kE+xx+PiRXB89d9MpJLzO12
U/EoWduTMHJPHgMQxG7iTFqcFtYy/CCNXR3b8k83xtb48KH5+17u5wjZlaj21xup
/l7tJEqCaHOeBaHmD9PBJc50C/M+lpexpudB4kFO1FqjdY8ZQ8hNat7c2mKbPrkY
Lv9qthPI62Krqj2hOgcPCIaCs0GMeD764C/CFsGf/qR1x9y5T0PrmbjllfphltIP
JtCuKxSN5Hjx04Zw0WanKk/9r93+K9A63tx58s0NQjoJUl9/VmTwhTHYP89RRJYO
qLDX8Jvbdne9N7KikFQ6QNExa9NhTvQBRcVItxzwSOu7YUa6kPrtJGdg7Llh9jJg
4pxzKfiN0kDVCGWkvjwo6EZ37p6o+xynOp2kyfNELb0sgFPsWJbuiSLWEU8+QKxC
mcSOGfGiQn07+l8eSUbS1LTkM0YhVyaa+I2gaAmNKSbbVPKiA8NoXVluRkD8FBr6
5mBat0quAcXC0UOKDQLG6nbWZbq5oWcNPWxSpiaQrqYw5DJqVsflNqSqrcg1Xq5I
1+bhm+X3L2c/NRiTPUNNxA1auwqnAl3MYv/igPMvMEBbmJxZOUIdW0qDtpG/acxQ
zUJjm0+Xi+zv9QBdTOxT7KFV7Wu0XxEI1RJNRmP3/8TOWM5ODkfBKMspcKhU182p
cAXFCGmqxQ+JcW2B6IYdnipCIqNL/510RcRUzp1wrcz8DQO1SPmm+Lpio+8ee6ug
lilRQ10Zr7GF9dZ/tSMKxVdtmFYUrZuGHjgYHGx4mB1OQTUHj0s883sIRuwdtEVe
NNhJkKKfbuZdkeDSeuNHsITslnrQFSONnbwgDXid5t/hUodZyhIk1vH9HEEGcr6a
lWgRvvkOOuxz2a8hT59nXGsvXCL+rEbwApUGLV0qSkSYtHZwMtx5raIAKKSagKZb
OPteeXJMDz42D/XPY2wlMdILRj7Bt3TLZEYBE2DxpnNhm/DrNk4B5YXqwn0kWLQ4
2g15QDbDziYZ8QSmzPA4KF5UZhlCMSNdfLk/qBN9Tzi6veLJzjMi931XWm01P3te
HNF+OAxk/ZmjhLWNAGmwRe8UoqabtmyT7q67p883Owm7x+382/D+vErJjV1YIHxV
6H9T/FyRbREAj3wXFz3qK4mlsICRgDjFKVioLWkc+PM8JI6ZaL6O7jowNbJshmTW
DQaOJDFsvd9nZZjRBFVJ/NEfkYq+r6JvJfXHQEVnomzK33nFezySZR/CjXY2neoB
fAxvt0ceZyXkDHJTiMsYzhjfHSv5xWPd/vmkk8RCCa1gJoAUpVL8OpS13icqZsjc
/9qtP6SPGedOgRKRbJU/hehSU1S98PJnXT6cQWJgJGcYCCGULxQA8LYBM7gaomCg
ett4uizv8ZdmJ2QYUe9MGGRkEppvAHWCugE9hZgSBQ95oU+sXXn9N8blNMqs3rH2
A3DOryvzfX6Kvsc7pOTFD79yKFJxbs6Mt2xF6iRFDlj1hAxqTnfxrsVyb9DOy3Sj
x8iQ4IuQrlapVIK1UoEBEyXOKX5wDEMewh3Mv5CFdbcsCr56Z4p2XnMoiqv9rAa3
0Cy7FwI2SVV3rYsf0knnPh/L6t3t9tW1g5zQh1HdxbzJUezS/cuL5RYd6grWND8c
secTsxnAcuJ/FvioDF0dRAwXlvfHHOtZA+nWJ/7X1myPfm65P/Q6zcOUahL8Dw4Q
ak3uXQQJxkzLAAxuLL2JSWi8GDCO9Lp+Kch/wOrG3d7j658fM2lTy8Bbwv5p4h2i
WRDwks3LROS9zynk9dAmlrKKD6wsnVGzdjzTIvsC1l+v8TkHP0XibbmCqzB1s9l6
UIzTVepJU2ifKIT1A7m/O1M/6TPlW3u/kEN1NXHoOtutANS+yODC7MwSsVqkD59J
9oJ9TCVOtm4/QdTi/WnP7nW/1xi7VroNLgE6YdkrRANxHJLEr4eqThFkC1ND5QyE
Jxao8wzUpROHsPB8gQG6ilY3oU3KShBdt/KF7XnG4NlH8yIhlIMxOTu/gFcNwClG
AsOKC4N5yuvZGFNnsjlRpyyhaXVAZHYhyiJKRWDTSGR3Eht87olDh49AyRPJY5EU
RjlqWYB8DM8A9oVrtznTzD1R8O6W/D7zm4rAfTgXStpIz2Gz1emnHIpTrbGaeefT
zEVGAC9dDFKln1xtkynq+45KrdUI5JXK2M+z0uyTxgSKkUenhS9v+L56iH0Ffxdo
wBLJ0gnMjlTpw7k0T93xffe6dUWyoFG6k+7YUmdCL48cFumcSeJLAf8Ds2rBRRu4
A5Cp0aM4QeoXytXnoMnyGVSvVqSZ8vxBSysyCYoZcU+pxHU6thiifElisJ3F+vOE
zNx+63YzWkWeFvyiRNemLM371jrLvGzurrtEGvqkMvlun/ZC135imefljIAJyO6c
wET3P+ny3dT4oT7f+i4YGY/ismwgCGX8CDemTZ4O1Zmg+VmHDM3v+7/k/MVyucFS
9U5qH9GdfmKCx98KBHUQcNO9m+5rf7mcM0GtXegVNGZ8tWI0e2eZSiFqINUe8ivr
5sJFaNVbCLMIMfUZgYQAiSwnU/4Ha50xO0Sar3B06twrNYlsbRE5t+m9bHkfbQtt
i0ZdJLoAsb+cgGgS/0FirYqbwa2FdfK9vOvv3U++i0fU4SNhTfvIjzKHoJQRWsMw
uHNIAf48bfHTBp38jZJeQXX2440zjGIeSwNx+Hj9lZs6yxXsJWLXpjtxCHBUZztQ
zOqohBiVZzztWBLKoArfXuxZGJHK3jEqQUfYog2gzLXtD81MJN5tLUi9+t/Na/eU
rpD+fFYI13LGcJ2QBitQ3VV+IUdOgRJasJ2zAmbL58Z0izncBpecwWNoNuJsnNj1
Fn+fWPS3DUQlBnOmiMmz+kI3vnXO6VFc224YHBA2Sm3IrPoDzsc4AaJrUyQRvdtR
AtHQj22V9DptxC+xb91Xni4UpJXKTKhSFvbM507lQl4IvS9jGdFiggqITB/YSyNJ
gdgMQgC5/TX1NJngMBH0pUdXCzmEW/Stk1qM8S8HKMNUHjCPLrcHoIJ1Tsb/hMV+
jDFx/DqJmqqrLJTTzyKuO9qzjsrTz394UzPwWIwbsWdzQWVmB6NKq15vDLSpxue5
zifB+DRYLbkP38d8QIHkAS/TKjiUL35W+Bw8qLJjsAbM/CreVqf20nefhws7rgTS
CF1TqkzNfGkWG7I3891lPN6Byltk3cV1YX2soCxc/p4US1MHODZlI75Vwsd1CJPT
BZOvmQ+9pK5kwKxKrXH/qx+T7I/Hrp3B7R+NoSneew73SfLN61wAslCKgZoPAVWm
2B7W41dXWMC3ywarpbcUyTRZdcrbrGiz7aYwQGLDB5rY/TywopQdJtDg+B8g4tj+
FvGUy/dG5GH2wwm7oNz4iY1FDDXDXublydP5Rs/fpRJ+3eide6FsFnopJa2rWfT5
zGudFurCC/tkSe1B3JZYcnnjPaRo+erRThZ3DVR71jWzpa2vS5RyMkPmH9urD+mk
WA9bI1U8Kp/NSiPmGhRe8/fcn6wyQWCIvw44LpuKMKG0yazid1U2SMCxzAdvh7Ns
lIbf30NYLNS2uYvy/B0Uq8GDx74ptO7IleWunrA9OsD5Rxfqbr47On6iXh2pwGgu
MT12SdYE90Nvw8VRzz7NwHpdVIZvjsbBnCj9KpIFDJQcpwVK501ybIKkrJxmd/Ic
19ox4BQdkTqUJc5FxF1vWloYgCY+3e73e2CNI07Ksd1xFm0++mPFkUx527jwF2XH
jpzo/fxCaFuJwmEUra0N+z2UXk4OCH8wUVJJHj1Yw7qWYOt5QZsvlzlDiBowMJX/
Zw77/cBS1hO8FQDBNvHxZqk2+kuiMjT1KLSxXcbdjvSdhM+27vD7peWqMnnTjHYl
BSmAE+lAVSwB7Fh0Xrfoz48hnHoP9T1rZKZX3s2hcu84eP0cFWPxDYQpWjE0ES6H
MnGPIJ7kHLSHYuUunZYsSJDaeV3ZHZBmfNEx96YC+QoMTlXvfbTGx0leoXeoHMKy
GF++pb/t5AF50I20D4Cqg+wVIL/hvmuE7IogVEuA4IsdnW2FGPUH6OKFKwhLaHTQ
7PALWtk5fgogg0Yb0LnY4gi/3EsIFK1rn6U4JXwsnhjV21cx3pb/5//PFlyuOAd9
ICSThdLzCQ0TuWxg/7yjFPXxUQ98X0zUTEga+yAPzICDynGozqFYj+s2+HQyaxu1
yAmt+ZM7zjc+lEjNQ6uSPIXz/qaChOrCwhAQKtpb2D/ETzMQN1OsTmK2crntF9D+
pymqsI6vdgf/kWKbHKccPegKSa93anr/SUnrAnawe3WpySZRACgi4hxqeM8Gz5Pb
9kNfANi+cdNSOmY1WXNjrT0ljG0YcwXO+KRZ+D/O1pSrTY2vga4yiG0FUtAF49HG
1uFMZFbq3D24lh1hoQhmpmkzp2S7T6JuHqT7kyxvgSemxtn/H1wqEN9303ZoB4oi
CC6dUZ7l7kAtnNEz7MNnnz2z1f5F9HIMvlaWVJS2XIPXV2VUGvX1LejH3m1OREAj
bRwk2SeUhDQLi6+FNzGahmT4QfPLPwzzeUmwzlmc/rCArh1fgTw6uITPlEQO8MuL
H3RUOm7Oeo4bg4mOUDOYkel8Hx08AR2/VLs+2Rine9yStvmLYDWWU2LlOEBHIRW5
WsHl6XrP+lloy4oRjhdSIs/i2Wn+KecEo/Ovy9+NTUzs6IarvkgV6XRRFIXsJmtU
Se17i1Wb3oc4h0JAe5vn9DGJxp7kN6zj08QBdUwFc0dnOzlvDb0QV9zvi1/R1kNT
7yMJs/CZVtVQARM2+/Mz8piWkYIOxNsNi0Ccw0x/FRBxM5JWBKo6OM9IDoy+z2y/
3B/qiPySQVzKneq5QIDHlAVSdp25X0noJzApaSKRGy8b4g8bmsUlFJ6dlrIaj2Dz
U18/pbUYxY4SueptUi+Jh2e6DXzwF2UukrwwgySYxFJVqrISX7E8SBx1xJTJJyB7
WV3t+SpqbKka4vK1usXmGtOJi+5eI4olirQkgq9jc+i7u84JtB9U3Pt2Ah8tsFBZ
KhQVLSi7gytGrhpniUe4D5leF4x4cpsuhz48L5qMaGenERYiKiF7Xuk8mnHVUpjh
Zb9Wo5gaUOVL9RaKsEc1tMpsJ2TOgX/CtcBhjseQRLZnBkOiCH+YoI/xY2uBYO+A
JcpP/73eTePmK9BZgcnA+5TC+kaJToXSMHIufIigaKUt9rBZMIsYf7oWdntpBaJO
qcqmxHRLTVdZKwMz2OnRlQquFreR/5LB3KhU+6eZzH6tf8s1hg1EDSzohI2haHLj
1HBKIef2PVATiH9H2nWS0Ho9kKuECSpsEY1Jv1RsCBaFrPWZ9P9u/ExjigtBfXXr
GHYHYGWpqsMR7z1zyuhN9vCk2q0Cu00yxk4C/OPo81yF5SPGP9rUcozlhKGLJ6lv
NgJCEbCaZlf9A0bZ4hpiU/QiraZo8PZBeYYo+Kk/lce8BtHRNMkC1IH7R9KOBFpR
hiwFlVo2eCHEqmZNWsa07/qjkfEDBo9gTPHtgp9VCqn47eity5lqL2dOCvw8LUWZ
32RzFIQ0h7wC/k+/iAcgO4dNhaoh9MzryBYLb2R6AHKDdvpCZ+fQkKDqPN3L+U1b
VjR4hmrkHoMwmcYtrgDF+FiqeZAril0iKJ2DdkUtuWDQg0BlU8wAbT4yUICmSKi+
/jhBQzsc5MIpvOPq16Ifmn/4TySVinlDnBcCI0Ng8tp7D+wrwg69rEvr1GbiA6ML
rwlaMRAVC3Eesyrmq6KJPxmRmKGbrUM4GgKQIZxfRh0xPbQH2I8r8ZOOCSKj+GYY
vk0ml0W31t0hECBSmfqPFktoDzLkfULfKpCCaZXissG6Wja1h8k1EnCVI7YVc0w/
PQ1peUrVeHNs6kCOqHVyYhaYvNXJtwFsABZ+sobitHwT7U9voK1qgTL9PmXo+Hsl
MAcxtvkUvu7UrsreCNTPBWd2zkzt3aY+blQeBjNVXUDzxxpZG+vs3T81713fs1eW
HLrmNPfvlNaFRSxj990QfpbE2JXFlskovtoPFwcnfbuBKZ897pJUU1dOAcE3UbCC
lGHV10JVoCm+2xFToA9sC8nfma2x5uGIsg22ezMDS57bP+TaEEtXW/lczx0cYd75
Pr39z/4kyYdjNoAw/IgX4XoRnChcTcMf9EP4fWcUBTP0TGh8sMDQM9fA4PRCFH1E
KBNLJcLvZPo+WMzF+8HWMIKpM+G9e+ArriBH9dgu/uBEiWS2vyprPzIX2niqiLTl
+EacCiGaIovmjR+US8g7X9K4Xtky2cKwPe4FHZpjeDH38tcG9aaYcSKg7JWHlyZg
RNQZWgYc05c9OyYaje2a3YhWtrMtLsDMUQu/spT15mZgu/arxsK2BeVvII8LbsYt
xT6iR9gKPZPxcZ6My5YOOvEjxIjIidqwG2LsDu5EdH+nUWrUK7t50m+vFxktEO1Y
0yAlKviFoeKTH4oxPKOMKZlLrVL9TTtPok4RJwM2au6gKPX4PKpxfkltBXo5w6td
A54NLDzHu6IJAV2oLbs+3Egl7KIchilrup/tIjbMAAADLLTbpTfa/Zmt6gPCz0ML
ruJCe3JnNfIEPw0a8rd/1NHdfN6AHenIqYYXa2olnbTMOQyX6vwS3CSfkfx4MT7T
6AYXCTNPSsmDes2yw2UL72lZuXPDaIRlDQ/34BES4VmD2FHokGlpR9ZSX1BW93Lp
uTU2bWMmp2lichXgCWOZiCqrgcKkPHGCIEmRW6v7JoS0v2jP7hvhZ7O14kiFIjBf
gm3MygxuVVaIroNlTqPCDHtXV6XXEGfSyckhzQznzCUDqdYvKdzjTK8ahSOUp1sw
X463kDykIytHi5oaLXZvBoda8W5Ajagc3JXbHgUwBCbv9K8jRT4OPYX98V+ydwAY
9m6Sws5yhhnE/CUaU3ti9/tOGgfabFiu/geBSp1SscQlIFq19UgMqbbBKmyWWJpB
N6obSOaEatGO77HSpCSa8NZi9Mp9z2uoKyLZMf9pSeKgIBC5PGpB5KMHENuoP6Ny
+nwc09g5FK5Q72iSlPN6tKmqy/vaFb+vlO6xjk7r/8LNMNwRLCnx/8tSkjNxn2rr
I0Z6+jI5rtARcVyKpnsdg/oAmIK3D3g2FVt+/4UOuR5jzc1J4JfymP7A2g7gruQT
7PNjYOA2/r9dBq/RzmgO2R8bmQfzAliwhFABeTa92dh8gpjIfcBn9hLvzVOEXoFC
9a9ZlgxN+5e/2+Kd9Ir0EqcM5tpT3GM+H5Ele7SSNPDuwG/K554WrHqF3cITWqeL
lMLQhRwhPxaIzZsXAhXIC5cyHDUq3IknCb4Cowt/CL8KUyK5jF9pqjbEGivNRxaj
9PmrZFjMZugBGZlLZPRiu0Quoo1MRQJwpKmQMb6T2H+zJuV1MEnc3IY/7N0nCZNJ
8s+pE6c/N1V4XD32DuMcSM/i8vfotPHcNSuTH1o1VuNQfvvaCN+t6j0geOw9gXYJ
Z80ICfwNSG2mlBXBIr96HWboqwnmszlT8dnhNH4fnP53W0HVoPlA0Nu6d8EMjm+d
uSylovU5AsmkQCNaNsWQIAwpuG5HBmJx8BgEiHOJ3q8I81LlQB/a/Y1G9Fyc9mtv
YVGeKgwSlq/eP6++4pNpwT/EnPWj5EGeCaXmND7G34bgdRPgcsoxL2SpIhe+yqtZ
CW7nuU+1YBTTxoS9KkAbLi3XOFizay0SxHKMGMoRu+A8YsCMadk9dh4LWN/PSRkr
la+PUUGbvPaKrSJ8s/CVqEUw6LSfVV0TbPITtKzuv4Ji7XaqfuYFoAWbPjA9rrLj
4zLukgafcO4K0NTsADzDIty4dK3e06UCqT/dpmd+yZDdCS8a4NFzljaWHt0uLDJ9
1iU/uuyL7P7WawuIKcpw6inrETGwoT6trE3HW8UaXV+u1L9OWe0R7ZTxi6q2ZT01
aSFN8Cx03L4w8jooyDdQbwBb8A81huWEuI35rujKLnLElgMZjpVm015opDQEKGVQ
c4iMbW9BDDy4DvNdmWI4TM1jeXF42N1aI0JToFBkhgtI2WXfqexl8IdGZeqmwSp+
eigVb3ggWvIIi+8memPCULW+PHfxxirb4pd8it/4NRwVRyNf7UANuaghVQOOWH2H
kms/4DysQm5usNB/F+wK63jmKwtjYJ2lwHOlmgh02JIIOUKBM2QttjoEDUBl/WP6
VG7yXQwwbu7pSEJwH6cD14U1cJaXcXITFIdER9BUJ4RQD+slqiBRgVC5lN12VRBW
ijf74RIWhr7o5CwkbrNoOGBSbq9s+yraGXwzSr79njTehb/ayR4pJYvkI4p3rDWJ
3uyDWYLrN1DvD4/atVMW3kF22dlLgBbp58ykFM6+FyrJnFyIq8fwOhms4qDzFDFC
3a/PLw/FFyygtTZliWtPkIsnxOaa3y4JCmgtvPtw2a/YzQ1vTF687h3QCFyGXphd
GNneLXtul3DlSi2rZs7niSbRc1J58ztpwEjN2tNohPYPxpSsoudijKPLwR+2Nuk8
n3HeWndj1i/dsCGcfIacql3OZGxXNfUtjF7wdxpYg9kplCowUoJmS6vIzbX5616v
xilxPqcGLyBFIVm2TC+rtHwFP9reCCLobWCoPD3SczPJM9DNzaCDT9lS5MrhpieS
XfHzHAggOYo3r0ofAzMsrAbMYcB4ECBQDiad3c9V5dzciU+TLCvi8bVvNOsg+rOc
7DwzhDaAdkne/KOqV5miQpJkx09WDatfAPRg9Rr7zp98c8oW1t37XJ1DWE0Tmmoz
h0kS+50lbgPBLUOfSLnIEVus4mfl82GLRyu3wDu5Vo3naG68+L0ilE3Tbw9SriYY
NFQpLqAyXrqmfSeSkJMiuc9L2/y93Fwbgk4K2l2E6W+WKh0tUnZ9CBPmj0lbeMhU
10peW9LoccBqGbMDOE1UN2i/LGXuwZECTIN7FzVQ0wFPc7Bz569BWEa0e7FTAfQC
Zwpa8tCUhNedvZze7p8AA3acGMY87SZbdTMwrSnZXLmHVBNQc6NGN8JJm3jKZC5n
kQ3UaHXVh2bcmfV95SSxd3v417JNCi8EFGwPO+PcpLEXGSdrVRng9CX2x2Yrz0Vz
4z5HNDOjFJ3du4SCHm20dc9HBI6MAkbBgfHw0fuMXfDsbzmMD8ldmXfoUpM8BmDe
RzVQ09H8vLYRBEIX6IJZLk6NFY36R6vL33ZNL4TOATE2mXFfDDZr+XsoxT8FdooK
byTphW8Z7jmXH400ZWs/FYPhPT1MS6cbYGTTX6fN4b4781qtkKCOlKrnK7kAtk0b
b4e6OK/KjgL3q/AkdixRiM/XBLKggCm2qAzTM/PwI43tiZ8ll5szgoDoeSPf4xGk
DrTsLJ2yAQyxqX70dcIVba9GMo53aHPdBipiE3hSfBF1nsDHLgRUpMebn6pZ0Mc/
TCMBsYnSw/3eQTkoOV1WzW1hwpGWFmWsnpQSzD+PSTgFF+BFXmrKbay88yM7TAzk
Rym2QPM6uB5k6bpeg00Qx78XyrTQVzF7GW/y6j+jTNPCkyDripG0kiNgWlP4IePu
kR6qfPhYzAE3MJSfR7aL+EU0y91VklNjdvScRsEcSatbKwBZ0IASHqF/mXaULanR
w7CK7++Q0yykQ5H0JWL7jOJGeDqE4GjdQOkTl73aWPM0UH6vWvzd7YCCQP0aIqI2
CUD4EUulqFLSxCzqDokRcQ4y4tF2VFPYkCmPZf8c7jVDLXR5l8t/5FKifH/Q2g6U
7Zt1zmGkp301Pv/gdmQw6+hp6/Pe74NBqxHHVjCNXwH84PsNZuJAPycx6mBknNKx
FWMZwTBDJWZpzCh2JPGgvT/onQt7FE4c6UqG1Zz5c0/V9IXd7MsaAOjdkrpmAw1m
n2mSlmi+8gzY5UAzReilUnZbcGR7UZTfskDdeZjAoE7OiruKIBYVDWRu/HKsq1vI
US1ihZgZ3vEGON6/xL81YxTyE8RdUPWpUoYHdW4I4OnkXVcSWOair+Ntr3UXSn7U
kciCYPa6QFjPuSs0ANJQOJelXT2U3tbZJH38+qyioMqgyK9RnGJlh+iKPzHpVmH+
+Mo3k2HRmFvkRjRY2SkXoEIBImYBlW92xEMWOn57f5AaastEkgzZ5W9RSG6lRp8y
KH5RKFudLg0/l1HyhxAcGEntkkSIT9Zp89R3Mw2bSDwXaON+fgNnt0WB1njMtjeC
4JSjUqyrr6Wf4e4Jsq2yyRusQk5t/fzE5Hj7VI3ITmWSynbt3B7K6BaDcrYfN9WF
u8/VqPehYSDpCn2aYyeVVWgOmN/8zMmffVPzOPm41JWhzdRIupy5AS+CQYBwFU+e
1NghwhyQO/WigejmjbgtOeb08GO0Ypx+pywHtwpzEDApHqdg9chvz0046yeQdj6j
OSB+BWx26wRHutzGWPb+tCFntonphpWlHk/1lXqsUYA+lAVmxgLs6aBHtiyyWq17
k9P44NIEQkJTdwyEiJy/OUhOGMilndakuGNA8zMmhYFAUd2pkr07zeMcDoq2A6zZ
/JqKK/+URlsIn1Fe9cdxThlDLWq46IzVEnDBYKzkypRl1dd07BS5OhtBi9Wu0d6T
cagucuBspTEA+cEEq3fxmn0vlfXiCpE9QBUq978IPfui3z/IAZwMsuJTA4Om3FPD
NczWwYW6oWapEoDcaU491bQiwtRdQrDJjqIHJH8SqtS/p3SOBVrMzwllyvN99aKU
5XtXk+pGYmr8QiaWMmn10h8pe37EZgoJcpa9UemzeQXomP1CvfuhCHSSHt0h5IjT
dTAh0C09gboNEtS75hIFaCiqDLaKWKSZ9MHUMaLOPSDsJ0sjjljXuGyl7snqwQG9
xtyC55fvKu/ow1wZ5+q9Chv63CNLIMWRjktVC1DjvgZN0PdZg0eO3uw04MPN7+gK
ePydtoxVSHQbX/6SKOS8a0oEvDfOv/knnyIY65nCMSE8k1mXAZb/v4S/LZ+LqVUf
jK8/xpC+L6/ApTVn6QjIO2pgqYcMgHi71jNdUrUk47uoGTC6rHIqbfOvbQ/8AePU
cfP9N9YZsLwu9agGuZtXhCdPXBl78Ea0L/xDQRZHtJs6bHTnoZK/+PzkouvIgqLY
4WucJYRhs9eo4ytjX1HaHU52Fiiy3gpED4C76IxcbWA3qbqySwyYDGOr9DzK2YV8
kKFELZ78mpD0L6E9cYPepDhgasonKWPejg8RqKGQrOE0DOdhO0Q2nJbDI/ogSVyq
xTLmU8/xghB+vguPg3L+zTXUN5pqPixP4fhwzVfPE1GvwMqKmgmtC18DWYmashcL
8rNa9GZ/F6lh9d4xBSidG25BNtmLH83l72jj5Uommvg3r5d66Z1mcekHsxa4U2mh
6s4lylU48Cic11LK6+8mwqFoiLvTmsSxNquRdLnT/wY9v3TYZcQ2PuCOA9bRQBAn
GJzJLPtCDp1xPaSEogNQBibXyLB/iJaQ1EM0lyJZ8p+lMNLDBPk4lCNJsGnltllr
NRZ98ZolncgQhg0h8yxpNhKO1yPoljcWYmpJ4c41phTFH1jHqFi2F2lzPoTtOcit
LxFC+uxr6978YX43sTb6WHpECtIe57BVKcd/WBMHE8Psy8uOPYoowNFVzeed+bxT
fUDHwGefz7ARieoOM5TM4JLvFF7E7wPxdCRpFDm6EzQ9BMTiXZz9+9EgkO/XJQ9a
FKQfWcepYN5oP+QR3MmkWittBeGQn031hw1TLqPVdzSGjXZ63MqrZfVWNx7h+dSE
KpxWAcb4NsfdoIuHCB9VFG6WzIP9yh9YtbhTDgOwIouX7bAjaB9VRCw9Rbzpr5Za
tE0aIdqPnkW8qVrhAjz4DcKtCdemnGpBh4nPjzoA+RfApPMWEaZSXNM/Dvr8nqkL
+SLJawwxhBrSKeZXRm4/KsmmXB0zUOXtJDQRf9wr1p18SmyDEIwQSzeKB52BcxGs
2vuyZTW+dzIwlYjuOi74HvSMwsarGArKkvwdFGS84wYuf/MVVHg1NRnSAIPX7UI+
iaAusk1/1x4C04IyRVy/ofd91Y2p8nYcbHjlcDMXPiBVBH9tBpRCjewvshWMkzTR
Q8yxOmA8CxrOlqOunCWJM6SaiqZbrLt/5vrJPtlM1/mCyFrqBWvTQ3f7STsrTGZz
tfWBHRHvLWIEbcfq2wOGP0Kpz5O9kHHAujoTW6krr+FQjwNUT/vQ9qi/jk+wUOWQ
2r3zH3KRtyhdkTCQ5/CvnD3c67eHSOhG4JnGbPA/PUC5AF4rcjJv/WVifoqSVBXz
/uYOaulgR0II1y79bYx1sdcR3awDXYbdrV19dKjTL7n/mvtyOePtTaTZUtDcSQdj
O5Yzm6EUMGxvgrDjrDCHX+mTJhDLpy0KjB9Plrwi5Tx5UA3OP9EjCvchzrR+apDC
WvPSi4rqmdLJ5u5+c6a/HE4jnZZVTu+7jHrat/44f4hB49+7qiU/xmmYnGCzd8j/
pXdVVthN6I60dUwa0IX7Rv8uc0K0l2pxtie/WkwvzOMkE5UDEkBfccobfiATIEoq
eLdcLcVKmeHsqEuaZ1rib0rg9PoYT/xnfewmsuZw/p06dyHA2H3kvvIjphzQ7DfW
JInJw8FLu6+XRGH6KYzK3xqAp1Xq0ySXOwV0B8KGGG0I+exUZuIuSknysSU9rtYH
YLfI7nm2wa/Jn7KwLzQpQpnQ/DNKwL+L/GZLVeWJ7F5q6TCesD2eYeeqIiU7yytx
718GH7R6O60yikxsqeqm2NwYSiHNKF+T3zsskwRdyGyxemufBDKQZFgX5OVWh/bm
wlcoOJJAcReTHm/tvwGZKw5zT3iYPKfRxlL4quq6QG+0khFWyF/6p+IEp/u4zxLi
NwTsIJWkFmk6m8mVppLpzV6Gm+Rg+Ws6ybksYV/PfJab00P1nJPwSQEdbKY+31rm
V7pW17EwM1Foc2QVNKqmQa3TB17aNIYJZjIwQ5mubI8LyY3lnpr5Zz7CKWsSoN4j
0TcBZI0ij+hOBFMDDE2/B7PkAhcZhxHw3O/107NfcDyt8m51/ggrlUXVSmFi2kMG
WcHfJOruuNsLV7VaBa5GE1rleKMCAmMG3p/yUI+GhbizkS83IekjGpQfjDx5zMG+
hPhZzF7Cn1cHuxEVmzy6NvvUO9YJg5lISPzdLivNRcDzl6YBvRa2NKf77/KHvwq3
RXttPPBzIed7dfE+FUjmMezqJ7ge6cMB1EC8FFvJNiUxcwNcaNad4HP4Ks3xaRuO
lmyKlhJLJt46JSz/q4RKwBJeiUKqVB8yaJk9MDLcqFGDUpmUThPpO1RZxKuQRtnY
PQS09RMZKKEHkMPjza5Ojyg+RO6tndaqaAixdbKI4NbzdGUDRJyWxeRVkU/b4nuk
g/7rbezOMpnYazKXt0Yk2b+ICX1nlQvBPjWNrtGew65RqXRHwCPl3TeyUyUtG7oW
uinEh4bDIgFN+PhkA+5z04aRqgnOSWCVgw3eBX6RZZx/KQzygDhSUVjNgCBoKQCN
weX6uCbMXSWb+qSO5aOBJwjN82ux1DeTZWZVK1DnKRsVBXg5KP1KbEex6uG63RiG
0rZ1fHLvXmxhuebL3SgW8H+inLKOeFmxlwLjp3TlhEbWlBdIUf13R8VXBjpV2vl/
TGMylYCSfyh4RKQbEa2QVgE86svEwfi2o4LHAXdt4kogiX3QJVs4ya7qjkVFDabf
l+i6CJU+Y8sYUIeMNOLcjfMBTYacsd4L0wqN5BMFOPxdpue9THpjI9Xar21ffktY
20KFB7BB33TkudfMMF+Hfur4H+WKUuOY0lqYdYNGY9R8I9IzvDfSwJrte1K3SII5
VPnKhPoEjb+QXedk04KJ7Qyio/afOZUa4cAIlCPPTUAX5AynKJ85DJLaemRFc8ZC
saAO8FCvaXBzfC9YNeEChTBOUUkQfzzO5G4J40CU+Sji/N56UPY8EZ7JPFuLM7+q
4OmdlnwRiYKldXEPctDDxTxTgYccEQy7PjpueCLmnUF10+5qZwsRysbiWaGXkMeP
c5Utj5kPgFj7QQaHXh3ipmSYxZiqdjtNAIi0Pj8rg6r6/x8VQpaZ+m2GOUQaEfxs
JC1MsvF5WJ/AWEp1WBv2ynUdM7fJZu0yvCMZ76UiHWR6vHzyvpKjT1owu4+5/KwK
BCulVVqJrweQYanf7Bo6T7yEWltYNBtxdQa/kRCC0Ac57ajUjegn7p29fx51oWZU
SWeeYtmlI2ivB5e7qEFJ2wCEIVBAw4EK/VKoTRU3LfJUk4Cst27lacJKzHCfYiA3
/la82IkyhYoWDcK2l4f2ErvaBUYr02W4vpFQWdADu5Ygob0wQ6vL1VFmga2mbYb5
tI87ygDePvtjSqImPNAzbuVzeQpvBBLhWUyeq6sgZ2eV1MMsKrF5clSy8tnA5FAD
/6qdkJejci8lD6Hw3ttDrU4nDuDThS9OE7jIcHP2KBO2aaXrC2ptVztaDinncynR
kCYXL6E2s87bY/BMJULa8cyz5JxQS4TL4j5lDivlVLdlgkHyJrRSAlydwpN5ecbH
6Pi/xFGZlwBXOXMICWGQ5CA3eiVk//2V9nB4Mo6qCnR2kxEhvMlVwcELb+fbh5F4
PT/DzEWEoiiEXVNTnKhn6R+W6nNWDl+6VyARilr2XNNwXey2rWYHhxM6Qunmgmo9
dHGu8J9eroPmh+66RvBmHZJ9gj0MmdCwr3o/5J7oLbOpxUNGmIw+dRKGLsH6x++8
Dg0V3LbPgecSPUzCwhAvnCLLTXh9db/CQs8fhf+8Jcd4wk0RiVRkbetOFbXjBmBH
4UInRa46L48BWNO11ZcEulWiV3O0thgwao2X/88qQKRL3HCiX22FJPwcSaWyISiq
M3PlVcKH2aEFMAqbjJPfmqd2w42Bd/BUCnSueznjSanYJIDBgMfo7rS0ldg35oTy
FUVqcm9AexTCABKeWVGgS6Oe2p78nWcoc5C6cgYwShluFBezO7fGZhGr4SAnqhcz
96JdEDNse43oUySRw/adPPYXaryujYZZOfIWycGSxKT52ZTHu9S0QDer4zZaT2mw
AXoHcrVf+Af40FdYx2GH/fGbmrJp5yA6aX6A3KgQ95Qj/UJP4ti3VR7hdSzlxvN/
C8jg37psoH/k6kBRRchynBTIwCzzbDpZYkgKF4gpp0k+fCZ0gBeawycASP1BBg0Y
183rCwKIldelxR0b/PeXuRPoar1hs474vB4lfxQWyA9ycyKH6GKOJrBJS7Yv4Rj5
/SFOlvw3heyQeEIwbeSQCRNkAM7asc7YIfwzh8grrPqdEjIxlUgKfLOBitMqsQxN
LXO2C6NlU5LcVV7nKTNfGX/mRBTKtwm8sYNujvUMiCoos2VmvD+Jb8aYV1T+9Ig6
xzw9Zn84kZgjOar9klAEct62TtSz7AT4/7UvivL31ak24+UAB4MhTehzdhbkVFQz
f58U9wv8KiSOi1C1ErJhGvQ7w/piP3JpInUL7+FsTXSQrdNgt+3o5et9nz7fBdx6
GE8EBufIfB3xFF6OauPCV1sxNmmtqb58PQQnkQkrSXZpP48QwaO9m42ALPtQWR32
AY0mKRRDmth9VhuWgwG+Dm0fKe8Zti/S6QM43EmkNeihFf1oZMoHahOmMZcoJDKI
SQFAASVtqr1hFErYlCFLwXjyzRWDjf2jwAksOKTth7F/wA3v6rcy86pFiVBgTGOy
yWFV/WU7JC83xv/wso4yL09+ZaHA9enWNhYQHz7BIHg3JM37nVKNHif5iZD3vbL+
nNBat4piC60hmkedkJoqJ9UKUwya4u2TYAFKnKO62/oAHs1In/+pT82HPVsTae/5
EbGvAT364wVstHeMgZJDCeA1ix3yG7z4ZHC8eDwd0hTBhPHvE7PZ0XbzlhD7R6Bb
+dyYYhi/YsngL2e0WzAI0qrMaweYqQUlG0BfUSfDBHSZ536w2LNzJOP+wI40IG8a
gxnF5Z7TJCjSJJJftdyRz8EM2M4uXF/RMlaPd95TpNaFnDuewdR4VkHHVC6VX34R
M36sdaIngIGeOLDtyfpwXKpVZ9ojsZnpXB8wDKzqpGfh98NWUDOFFzpRVA9565Gr
0AsIXlfOu0XiRKRw8wBbKwPxOqfqDec0su3RFRrCnGh608qKhKzWenFhCm7x/o89
5QH5Qol0OJFwbUuZPMJIgsXtRUr+aIQo0ef50+oDLxtPUB0q6U3pEwKpf/ajcGsb
TYKAgre0WJAbibHz+a/WMU6L2mzxlT5myZz1Gi5bYKClgPc0AY0uFXTorFeXFMEf
1KmkU+STSXBxRAhvTNl9nWwadjkk/EOIMurfnjxrQlui6jZFL+WXmR6DZO6KNmJW
IowdbgRSyUo1R0abjgT9fUVf3QXg53ckkqDg5Cokrnxq+gB922+eyuv80bXeyULo
9ZaVxHTN9KIcGQNwbxegQyisMdIhRBm7zsDBDrGJOHmJLjNc4VMM/CsSs9MOz78R
AQ1S5dkESwp6RErpTHooAdiTMSmGeWB9eT64hWetCYUJwj37kmfPXWZyOLrUtp2f
IuhugxJAwIoekCu39aQWw7ACyYoxu65yiIRrDLm+0z8xdB/BZDvE8woiwHWzek1d
ZqmkpySbkVyePPImTf6E6cZ4B8NOLfsa93Q0qhIOd9s1O2DsKUJg7++CuEmi4gID
FJIq2ox1PB0UYx2KSMAwXExCpWgne+7oVLpWrwxWHiucuu2kHJ13FMvvg7uf9leB
iAoS23OzTaPA9Rg4jcuL2gCoSYurGJadYoGktAuqZhqJTvidmJEYnytmRjfpeCmM
AeN4IKzdyX+OFQNhGqkDcX6Kvo+un6UOOFBSPH85QRWN/4FFTMTxMWVXBnMcAh5f
l5Yz9/Y1pt+S9RrUwm5uaSMmm4qO6kCtpPS6XKfgC8jfekMB96wsXW3CYvuIl8qe
ALFTULWAMGpuHu3VryT7f9um2DtJ98qQEGUNDyq0KjAX70jLhTKN8ymD4sjxNncz
//ty0Nz6fsekzg7bbrYLvP0iW+BZUXHBbrgBdGVfYZ5qgrusPMG56Qkf6LFmBEDS
tUx8x60GpzO5iEpDFVDZ7nXuAhZDRDQhSyK/HljCYH0rYJBY65DaUd9qaMPZC1Md
F3Oma63p//7UyJ66qJP76vKazMMIGqFk/ljW9MFJU87zzYt7GE45eR3nF1ACPXNi
ulhVckAJKxL281LnsCt4EFrtEFatxV4zSx6dUTLCieFplAjE6hW1TVD8Xsk6Agn+
Yfuy5vKJJhqYTPusXTzaSSPIeDkIcMFUqbA0sPl8qXrvA/UBgn2kufrneDMqDka7
grlNDfj8HuD//5QmrURbYc86ByJcMbYNGXaa7lnBUQ5XtKtwqoTRTB2BH9cngnLI
7WVkhqNPbbHPLHqVfEyuR6Klrg5cV5zUO4mCm9Wt9GWwvjrQ32sOkS1NeM2bLwC8
WQaG7wm/N+f6YA+t9DKpRoIxJj9xSaARv1yddG5skAxzLLTLgvRVpUN+/Dhh5sEb
6LrcK+1aVjAAP4/kuwosui1j1lG2igDl2jOz1D6w7i0g3mhRcsszxjx0fZEGFF9q
cSwhIxm0dfHMRXxRC6es1a3S4iPtW8MzG45RLAkyJZ1I1BIVuJmWz9cLwdMYNPSP
BIuGcGN0gQQ+3Qd2gMJeQeQVnYjVrT6mBfsjU+7AvedkcEqlx6Yh05rts2cc1EEV
zmd4T/BVj98viP+iA/ztbeIZPueN9UxU8StFaTo5+rskkGVCVMV8JmUrl03VzeMj
6N7u9XxjKikwyZi52t0jMgd9wCq0mXp24AZxx+VmZLbg2qXiAGSTNYnOjwsjnhyn
pr2Um1zCMkpHbvq4TQhn3tLfTkUGqAD0bwQhEFwcpKWopIRpWYrfCnqR/doAIHHb
bq3sgAoVSipCNQKi2f0HS7LOOU3MWvuEj3+aEuRHjA3afga2/eSW+Wuz/wzs8raf
FdAH5Q1pbYB0PD8q2ZyCQ3F5MTwRM+5AQWvx8VMOBF7zpiFBf2mVQPZVImjQDsap
/wJFidPdcVCn6s/J+c2PSefWZRHohzx22Jhk55NIOzgwpXI5zt1kcDAbc46XRKnw
SAUO73J3eAjQebsOfnWuAXPAUevhvVbgHg3LywxEDsVyzEvdYeYQ4zALcGnTq/8y
Dj3KhkUGVqacPSn+gGvnqbWxBMTxvb2hbZ/5Qey7inC72mwFw6aoQaB4SMsFwS06
FUEiQ60DRNbUDI2eHcBpSBTae0J1TMmZvoebaDqbd95IBCsinhWGuczi+nzlPXtT
NRZkJdeRM9zSVs6kWXUIFgD+J/UxKzz9hZQI8awDX9tjGcMvNzy3v4DRIbJGFQcY
1IfSBHLlBUgUV/o7P2CEmZH6AQOiwJi3FUMRn0g2JTSN4MNKRhLsUIEmaTCXEh66
5sXdma+AoSI4BFysEwArzy7PkLPgUW1Tnmxf45nkvYd+PmUWFqTHSUlk6+Ym4hlh
BhYbN8hBRY+3MIfD2IPhQs2Dnb8nrqyOJHRet7MreoBjHoLzu1iqTXwKPoIFZJpo
63H7D8aFAg7ICOb+DhMUXZG0LE/S6cfIkWbHIrVFVWFI4+ivO5AzvB3kDHfkrqj3
tCY51eZQOomfH1VXvJjWm/7h4R/QX9MHRsKmnEwc98HSrLmloCWgRqcA5LCHNzZo
2QdKXUBSvE0aHC+vy/YCZB7KCtbqMyp2h7/oHHQaSzbdTwTDJc1n+7sKCGYF4Nx7
psMI3dBcB5hBUOqe4zteEf7TgGpm0RDmfMbu6G2UkwUOoPMHusX+AV3KNZP4WMEU
CfsENGBJ8IMVG6c+QhanSFLGsEdOZyNJRY7Xrq5482we82yIplyGzTSHEqdw79zY
iBAIRqmb7E+nF9iz+6oC2wnRAjgprIdWI9e6WMlRGYpBSSf7nPrBTcGrDyai29mV
wECDnD8rIIP3i+a6e9szjVtugGH0gMZTD6mW0jGWUn/EECqrmQA03vX8TbWUQ1LO
u2qe0263rWetEs2zfO4zM45DIkyRSsea8LnDDQyIu+HQ8QF88VyuPrC1wLz+3ZSa
MRRb+HYEwU7UlAVmZm71ikr7XAsW+0A2Z+jpUes/9dCkGBOj0WEWJnqT6IqMQzDZ
cur+c0B4Se89mxm8E4KoTOGdxRIrE8MZrJ6cFp+lCtYlZE54xg1i0gRKlNy43SDm
H2/sVO5xhpuUa1QgMXaIQi8jJDZVtdawfvTn9rzdoXurbgFvE3iOcrVNgLKgGv4n
cLbm0dnewzZU6DujjtxmxfyMjcv5RmHCcS9AugA+vpJItWe4ZL+4cIqMHxld+OLe
Bbdd+zw/rCtLtmuB1+PeGMO+s37DrDAMlcd7XZCrsAIZFkqZkyvz/W/1sL7EV8Fs
NsWFV4z3z8gJ3QuDcE5KIXL9hp/3213OCKPte0WApsbHE5FIhYhg7sPauvHuzuZS
d4K2XXyU27D53//AWYQhkcb9teSrnn17V3xY3Da5LWNGGeqFJUto3D5kg+rNq4NX
DjuLQfOslDMlUxz4CtRy/3m11uC0361MLMW0xWUYjKV8fcVDPea+ufDhRGOLSv/8
m23e34B+FOu53JrtiMIAEp6gitgKLnzhZwUgbObcb+W9iylDCPL0eS+EpBtH57HR
DO941wDxp+eHC7GodgbypbTkyt2fagL2Fy4LnZFHUBwawcH1cbl9YYtQnbNw9npK
4R8wDx5ud4VTx0U5wgZBP5FUah3arh9h1eovRPJHbKen7UiYn/EMS3PDuEJxQ0w1
orMtplgziCu9r4yS9BD39o0IkiFJZsVc/zO5tO6TH/rqqY2urfDw/R0yFqj2iZ9I
MI+FRFIi4+9rXOq4xwnNgd6c2ham9cWAdmg+U0COtTqCbG4Id56I25pgKCSC2c2C
Ok2ibL+DhCdu143yQkRWDHU1MtBIGNywakkEB8CaCYhHkvUiM0oRdnmkCdr0t/gS
fR6XPV0pikxcFxx+X7FFN8kl//VuwL7I5UUPsWLVqObrOyMwUIM362lg0BXUjf3T
K6A8On1Hc9JtOqGY2QcCGz4CMt5gM8nG9T+htYdBw3KOJV588vnzEtsTYHQQFLbF
NY4p1Ou6/+PcSLXr+sqkz85wQmmtIspUGCwPihAMKsRjCafXv3w27EOQxl6dkLFm
+Q8rDxM0U/HAa7BIU/Ln0GUAzYFgYpN+f15HXb9twT+n+Qrcw4Db1JGnCVMnwv9h
ucUuLSvFJF6MI6CxlhSasVFDI0M8J5+hjl2aOryifpMbg+WCcC3lItM5IZuuOK5Y
J26egatgHG8dEkWRSUp+Ki3ar4Dt0faWs5aXZAnM2D4zmvI/Kil9pAhcjFt0s7Oq
/NUcvEvkDuvigZ63fId8+qTaVXJx6TtKSOFNbs47hg8ub799n1Dx+bMdqlxzD2c9
phvyFw0th6Mkb2f/HyPCSCdR2aWGdPlvyZHZOQxcxuHbYwLqvCaXAL08GuyAVW9w
p+Ao3XWZyClXgVIM0dbyPf190CY0t1EAGno6ZVWcj2u52FJIiRfE575mSoCNPigz
3Tfmk38AAb2jVbjnix/iK5lJuEb9nMlwWyo24qHPIACXL+j1fYCCx+xTnhC6Shkl
shnl/IE7MdgrG0Fl0Ntt/DQKURkXBrx+d0BYx61Cyc3iS5hIOVuYejkBi5b4bkUC
6Y0RotT4NhAcESpaP+z5czUTp3FZJBdYLy8C9wDZE9USVEe0l6VJs7btsX8zhBEK
zN96eC6dV53Fz7XIZ34spMaz3t2iQL04/yi3VlR7j9qrv7LC7hZ/RcgqVXAvWLpI
QwZllqcb+OWqD5MJYyH5ZKcCk9cxcowrtEe8rsni973HN6bhfNQydU7qWQ7SY6Lz
DGlBXdNdNKcbCV6wpeI6bD675OCO3F1L5b2W/s8m5xGjPGZhiBYRFGyqdkF8MFyo
FA09NL/CPxOjr02czYMrEAZSVWjiphckejHJCV6uaOvww9z3PHj/6O/XoQtIBsjo
6eO38gO6kupT6S1mBmogpR+NfBbSO+q3s3IQMjNL4wXH/ttTjSxe5YpN2mxgS8oY
tb+4/xvYscu59s3oODvnzWxXSLvFMGEQTNDyPPtGo2Im9cGGb0O8b8NP0k72BP3X
3eNh0ackPCF/4kCYvxeSTn5I4ZZLlTJHveKC1M3/qBKQCm8teG4T4jAlTts4hA5B
F1AbsOHDCE5hDABOKCGrGXEsl4lf6x5FozvosJojHoUw3kQGaXx8XJiRFVloIhto
UYV851IAlIohM/jctIE2wa5wQf13Tis3A5khx+U+jnUgqx2hlBc1XftGNd3dk1rO
yIgkdwrEQWwDnj8YK7KTnXIREqWizNsUrEhkxCR9JDVBmalfF4+gknuBX8rSl0UJ
GITP0L3ZMszo2vNO4DIFftW+oKrBa2mHr2ONqThahqSbDu1lUtWdOeFa6QMJKVOw
bnnlR9IsyTWV1CshVB32zH3GaEPOhXgZA+yOnFGBU/Cjbge+hBrwcXZbx5ff70A7
rc8dzA8KhiSkaA6kqGF8uAvONOhQaV27VZt/UtuVw9aloOJv165FOrBr9FiHJKkm
THPFpVftWIpDbO9ruuegWHmmjEYBOKlIjsxXkoiPRwH+HEsqzyV+AgU41GocjMbn
Qwai/ThkAzcuxxYLA9j4JfUYKaHdiNwg/1CeKDGA/C+T4Z9wAQs+TtteoyW36tgo
VaKSNs6pALs/chIB43kP0JFxk73/OH9U+ZtThlRhvFG2JBddiYt1IAJ1TQDai7ee
S2Kkv8AIusZ2Ll+DhAqEk6KNGO5MUqTbP/5Rnlec17NqevxxcGVUEgLbQcl+eGDK
XMB22ZUme1mzLQRXS/vTWUJk7R+WFSqb/VM9C984k2PyJfyjF3yvf99YVt6wtA0d
3e9CoHhzhrT1E7CS1OuaReg6R+VIRJyQkp0dMKrFpnsbHY53cf4CCL6i9c6Lepnd
2qXKbXEmVzZWRdChYqmnQ3s4qfjxbeITnWakW33n7wEHvF0eNg5C3mIo9PY/y8Dk
SSTZbKiBQLl6xTQfcxlMRfUs2fWgYAR7XG/vwDh/kYui6bPr2fxCQmVD0OfUJRuA
CMbCnMp5ykStf8kWcBGfASrl5vj9/m5WfOXeigQI4Mq2lpkzZGG5zHulROqEYGWn
p+x1qoNeXjLgW+r6oauPwvDogy5u2SSbWtIY1gYxUvlsCxTITXJdesLYRuAP/e3w
PkzIvlymyFsmBSckfTnYoKGa6tFJQz+NOtLAyTjgiwFacY8DTTXezKJGRY9tvZBt
9IC1I2iTMXKAV53zR8exhIGLIZ68iw0fMWlBS2U9CrlY3G5o9SuJtWXPQ6ZBO9Vt
HRhkR0RCiLyIKhCGKhyvnZ4a7f1diKmPU4dRJAGsBuLTbd5bVDAJ7oehAwNUzLqy
SHmaxs4M3JFEEtsL1VmKx/xZk4V5y+45ChXfNjRxlTDwF9jIrUU4aaQyC7qpt9Ku
D7kEmMa7qk4GklKPxIOfVhK4bGFyk9MUTJ3vSQq7VCaX3GmhklPleUogvZto00/y
nw7rTT+b0q2P9B5dblK2SJRDJIN0EsQCcvqf7NQPnFLJrla4rQ2tnLUkC3UQJxYM
Rsl2kcwyQaBuKFK92p/X0Ai5voIHxZA1Mw8+VmV5fit819V803b3h68pZG/dKyzM
REfzZdkzIw6kbewEnOaxs6+6GwCegvrZsb4PzXxGbAU9XXw7ZXyRvHlFZPoWevGV
dgcEPIkb4EfJUnRMefbIoK27+zpZRrKeRRHHstSK0fhaBIOMElluoQNE531VsRSU
jHNEKDiPtcrNUnUj5ZJVQdmw8iWv133z25ZBlFRo1Sm7rGhvC7DbU1fRABzuAcDh
irCQ4SgHX2uxmEZtY6CAseR4klzVqgSWMrUXrTbCI+HDsE0CFjTdjDpq2h9N03Jn
8gHjRImGC3hzoMrCQqbROcOlb5Q1Qi+mB8VwUwbxaJpiSjNA/vZ72bx4TQq9Dv8B
j/siCncyVeGTJLj64IWOd5tiX1zIQto3hsdAG6IAbjtupbNn93H2VPArzD9V7c5O
F6PJ8UXpi7F+pSNTIBL0WschOpeGPTcM/swx+Hg+lHAjUGAw2fYy2G2xDiKczlz4
XEepE3G5TPevi63NG0wOllku/e0s21ILmjLWjEiDOOxKSscRMWkJ8aQJh3xPqYnf
jt4kxKmD05NnZOlxc9l1dxlwEbpgPVl7tk/MNqHKBMfhb+9uo2Ts+qLkCWdibKqj
oXz2juoiDtPFSkJs6cLAUvyoPQhCys5vQNtwu7g7oM8+KOWH66B+i02nV7lGvAoy
i4UY6NW3vygnrq1hd3NTFyOnLM/CXHrn76uoYq2K8iNye0yjBxwmmEOiARBIxIMK
GJZjF6jHIc42C8u/9NcQUF9S/O8EbQ5L/215m/HNsI97JOqiNHzuTdClJaoWOfCk
/zUqW5tEdUUf7ZZ3rFPC4QEzGuELFXZpUHRF1oYs0dIlvk8Itb+iB/wQn9WkczgU
bqbCNnu0jYRJg/o+VngINT61gyCbJzfMLT9GTbpmq5PmjdmHnt9qS4gl8VBEswoJ
h0s0+zHS3J9Vmum0Xxwmv1761DhC4QKZkaWV/sAtiswSYBAiAkdPndLWvflP3Ll6
0eQNsoebLlwjZN1rhJ2/b53cUoj59wCJgg28Su3fFDl8nQAUZw3YMO1hcrS8bd1P
/mvAFJM3El7Jilm9vmx1Mvsju3oy+9e5xirT4KRjZ/6GQarL2jZP/dtfp3/0SjSW
p3czzRm6udsyB1dQeGvWik/Le5sDhOtW/IL+7jgQ5v1blFEA65Gl58Eiu+C3rrbD
/RyksPwq0No4jxn+IT1SScGuWz68s2K9y7q+aaLOQya4mb/zSLk83TOgk8zz+SQK
YMxdPvRFzGUqKZodwe1oAL44BWiaRFW27QrznNZW4sLoRFAzSx7tKElRaGyegvFo
BiBEJQTcERFEln8wa4JyVpFmrff3vgoy57g19IlPE1ejTYf2o9y4PtJhWEJNUZ8U
H0OhKbjdmUbwf0kzXqKXGOTCEZ1wqp/+ExUE8eKGvuuTLj4JpT2uJvv6mKYu2A9b
AUMU1sEvVfDwSYvJYnb1L5D3ChjOy8kvFgyr8uA+dbMKFbFta3IyNLk/ShZ8uhnP
NLh7d0HuThVQ+rtdgzgZjTD4g3HzXw5bwbq/XSb5MMOqMpKwPfOHMAWRt7Abqi55
41gMT5DlGjJbmIZAIUZ0G322lDODpqt8k0lfA0RtEUA0VKqYrc3vzUh8axYRKm3f
//5IbWJWGWTjOABmiQtCrN9gNeDreJXVbuLRQBojpzbPDuCLbExAIbTS6rfs2zT0
RYR7TDuwtyEFTU3OyC8aLXvhf6jjvHF0Ulr8T+0i4fFR8RDwLVXAyBXz10WxxAwj
x8ThsvU12Fbw8zTPsG0Qgw1PAkccCJeUDcOgBKuEeVxkMvXYotCnNkSyVbGCIKTt
8nEcquksjdvYDGmHv3LGfySYK8O0NS9zTEWVnwITrtU3TpK6nZmzzVNpE6o/nlkz
e7yLhxp5JfmTaQvXBeL54Z4WlgaQbZTXp1FxB+/1iqVekgZGkipWJhNPow3X5Eyk
8GPqDF0p/bBBCByiLXj/G0qkYm1AC9vQ8mbhhvOu9kQh8GobpNYspuaSHW+xMtr9
jO6HGvMYiVhqbvuo5/idRKn2QyEKH+Fq3bkVSZMGAKqn8+0H4K3I78vjJsKgVzP0
2XpyzmN4Sn0no2LwasrffQK7YSmyEMrAoMcwNwDk42dbrRi15nnpTDfu7Y0gdFdf
OMSXMx8ZQcCLi/7ADprnf6ywTE08avgqY8OL8tx04I2fU6U/DH1n3MRODFUhfAXo
usEUDo2X+bfTTSy56oNXbaxEJb+zoWOKzHe2o35LPsGd0MaoZRAK0iQSJkKe+V2c
Ime8xbOPpF5DEeE8529hsf0DcqrcHNx5zd+9cXk9jxKWhcY7Ap7OeL3yADoo4xfm
u6BrGuVhJ4jt/PdyWqlSTKiMeXVOE9WLSWDWKd6rTPcHUMuyF3rfkbt8Xxnaner3
fbKg38ekq5fiW6Tzvh7zKEuGTI3DHeAweKhMkmVf2HcmO47JoxDp6Db2yvDIrtZr
tkJUnEj8rFMNXTIWR8I7WGHPodGDgOBQUn8ybLVq3TrDru3CStedJ4n5NAcpa3Ib
jqtDbVa0TyK2WIjIqisUisoxX/pdCHU6Y/Hesa84luL24MgksDAIdmqb9oYr04L3
y+Wr1XPNPqRvdAlVZdNDrhMEuGoZ7H/ixMTEuq8fdhp4NPYCgV0+45zoTElhetVn
/hn+HNKLWEmSq77Wl5HMA4BWXdjSRw8gm9DiRn9Y7jOLpN5WYmYlSUaPKS/t23yj
O0b8J9pfZqItNVSqGlUCpy2ATryBNuf0OZac2319oSBAhS6iV5J7Weiws5Is00gx
2gnQ44f8H867mLVyn8y6qRJZtpEscu2waltFUbihiNG61xujfjaRD1SbAVtUoHqO
11c1B9dP4LlNWD6I5H8brHVw+CusS0lsGo5XN0Vb3ymbOlZ9QOLRkZ2ENHrYgHQD
7fb975qBqhfNf/60SR/HFdTgGHZnkSKX/kWjvs/TsHK/nUK0jqlkMf2x2tJtaV3e
3mvwZec8Dim7yrtf+ttd2ZlvXTa+ZkJvqZdLj6eqmAFuZX8+n1oaaAU6ZrLVxWlK
vXocX4su11fB1v7LRlhd5Ed5kbjvJ6y1rNarfeq9iq0hq23Fdh9Sme/X9KW4V7O1
RfcYrgXE5F9VffzZESz7tIIHRTr0FIT0SJUo2Y5ahamw89F/WgiRlfYpvkZTghNe
0jpKDs7v0JkMGIMz+5eTi3ikmZ8Kq4HEPtvQ7yJYrcHZ2BEDoTEBxAQ8/qTmwBtQ
R+4xb2jB91N6TkOp4/peNZUlzu1MYeLy1YJj2XJSNM/t/Y6tFcq/DmgkpVFDxgCq
i+ZGKEVislrcapqMsfIkw3q/z3hkVtMlXSpw+NaC/LsoYOoNFFjpduQTGa5Bkd5J
Bpf2pLK31aAX9dOCE942f6YbQhct3piN9CNgkNB15HeG7ERfbH87bAILgP2uwceB
+RAsY3aME61k2xnevdzOg9OrrlHITdaqF0hjK44Qchd5lXqdv7OfogWJ1bsvFKlH
ilqNHMw93XAdoDMzqRRjSMRoX6KkebZ0ycgtR5HmSCvUuY8IEoFCb4mXP24jmVCJ
chiAYEawYrrunjvpyVHjYeXYAET/eSaBm9INMa/rpro1meWVhmHT8noWk/1lGHnJ
svT8qivEXdqhwdhBAZf+bsJCC3BdiVd9lDRSEC1RWeqxNf2tBeZd9gNWg3IB/Fuk
8UmuPcdabBZnrGNQHHTJ7LKsCj4UsZABYDGuvn7WRXGvTeqXL+VazGt2l7sQzQtr
G44teOyMVcG7wj98veVGoRdNF2oflLI4n56wSReN/NbOH+5jnNp8614ni3Z7lym+
qlolWw/KsE85/+JELw2oYYVUZtwff2vT3KI2PANvZr4Ey9Mb+eQFKRDsN2hI+QWd
agmV347A7CH6dGyYL42QO1q3c5WVbdR+MbV3DsZXgdDniqJoR/5ZiV0992Kd9AHN
ztRf2LJC3Q+B+j8en04q3EvkzRvRIg8d5aUzoxWFd/EUbnHXN3f90U9ohnkM2AVs
zSws3Bc3/ovOCVd6a0B5P1LZ4vhDmYL2ZBLvVVXv7MRyzTntRl1orjHVEkmD1TJE
2oAvYyGxQh39ezwtZM4ijlkNcQKTL9zZ9Wsa4OrXoiYaE6UBa1H5SC6YkIOwpEIT
89LxVNBZjwTxfGl9NsswR9dvW/ao51S8PFfCZh4wIUscNY+97vvCbEiY5E/BPMju
7IeRyjc5PWEOzpj8E8Wyz3nl10rlsIhTWVSrentDtPnvOuMhmqJx09BEbm4qnijL
wo4VcGCNCzCeMBjV+BjYBlol8HXx7z82hvXziMTU0CXrxnzQK94GfVhj3Rpet1XS
hCtDHhuiKEwbp3vZXIvnClcpleCxFX0QKtrIvZa5ULXk7BUdrMfmJ5ekjRm5BF2E
E49LIv9M24of1LW4e95H4GDNQG0tuHq6Bl15VPkL3Hc/8n1a0D8+tMXh9FdwZ95I
Jo7Pp+V88fuEPptoE1hw/7082ydFjn7IrXP6fkdFep3xAf5G1V3m8YlUU1JFpJYJ
NXz9nEpuk/tPFs2iJNBhiSGI0bBbEMOVLm60IH9icOWw6HslFr5MwMMTsAXpUMjw
ZMESYI6v5R0RYLBa9mOhgXzR+hhjZ3kaqvmckpUHNtS4tpvB1uwTixJZjRLZ/YRT
HU2X3HvW2SWgzs3R6bGWmqr0SsvA2AmlfpvsVkEuWTIxwMcPc2ZaSbiCIie3/P+6
bXr4Py0ANHcOxIHXSAF5SVkT6PGl4BQCrIUmg9/AUNTm8ZsI2N3+EPwKqSf9u0K5
E28ycwGK8BM3zytjCa8FmtOXHe3ktKHggXeINBJ3I9fXfSOSPT+vYW63YemzJ5vH
PGedzAuv5QvY5gG6z8jUOw2vhpXjufvZjuWJp8JK8qwIAT1VYDK6/rNxz/gLZV6M
v8cyvBuHS5Zsg0ltnNuA0giFgNxZ9d9MYNgXg/5qiATDvHxaR+Vs9t7LxdKlSXud
np/69n+GJtGTnoa/mNrMTDL3D3yYom6uG4uuCqHNfYxHSpAoD4LH0C43aqFMLHog
trriUYjBioa4B1xl1bVUCHk7nN6b/IfmKFo9RxfgmThRHwLFWzLARRymkIwIec7V
a4+UoTCVrIDaQIOf5v1xUHU04oKYMCCytU/Bl2JrTGmIOvhAcBzLs7ZhlZImg5bL
FsUmxqoZW5rX8C/yA2iwKXKvZyNGDYtO370AgxKtSjXBHlb8dSIss6tDK/b7ojKd
iMLMajt6eeGpbmdpHp8ezbq4d8tzXyhRq6pNxWZrRm9XKMe1KzaVYexzKW9h4AAT
WcNi4XmPSKunZOmpvBTFY7m7KDo2XhXUYLTnpezzSarSdsyHoyyvnD8zqu+f5YHM
w9jeVKFexPZcNRat+p9cTDuhZf5xO0G/VyFUsuVyb25/4yxaTkGi1duMK82kxEWR
kDXL8wL6QwCj27Ywnnx3UQtM/EesUxu8iwkif8qA29uZNigUqI+8FHPiY4IwpFLx
l5AkehTe8eorXWqSZ7Vsj+VQrsusnoRcJQzEJMm1qbHNYzk2mnmieCSdGa6FhOsu
A+VP83l3GF2cA9q6iXSi9F0UqcOapLkCXWoT3P+e8lZQrMD3nehjPMKyibxys6dN
fE/cskb23gE69a3ITo6kYGYFaV2X8ozt53pHbTo9HfAOS/SsrPBLU01JAmTFCjRy
+xqVbiX5lIJmkt0qSaEc6MfFWFQDDidgeL1CaSV9e+cfMO/reZ+MGxHXeqUozZt3
SaBEL1dFmdy0fgRGwuaTxul9YcULWdDEctebjmjNGHtbWlwCzvtvrxMn4eJjyONP
hNIZQk2Hm3zbrdloRt/iJt33hkSx0TDdYU2wEAxcGv7kzJ2FBJBgBtYtos9vFbaq
IW6eR/hhHvDl6xC1veNg/BodsDRXSDJmGUFKN6SubntnO8eXbyKFTcBGMGWgB5s7
mnni96/z4UxeqvewPG//KXOItv3laMa4+zxTn5CULLqiC7l8V6zvRvK85ok5JuGf
EXu1wAwbVBtph7JlHJvfCgSJNPYMlvDoZGzF/34L2253Cf0WGmLLtLCwh17XtGIa
yET7KEQ2d9znR9wasGNCcX0LA8Ur8cYQG6Cu2PiY6Wz2R9gJ254jNUnK/zSk4TKL
eWbfcqcscpej6fyMzRiLFK3AD6xHwEgEUYbLtM1O7kuZ8bBqvwa2TAFd5kLiVXvO
GcPo0HgrjFlr331qM/5dcWe3wtmyTOSaCREGjKF/4NrSWfoT2qKMEbiAYqCGN/Wf
cgIV1/Gcq6ER8bFAD4biksfCMpqaV+V93+72G2Q248yOA9Many639KjZuuSCg18N
wLmUxugB6kO7dJFixdepXU6t/z0k0eRuOCFExQSM6D1+Qz/q08xvh5o20P4nl4et
NR+OD23IEKMkRSh5TTI9U9iRchPMTBW3ainVWOlWKLx6IOwPfNDAvi9qsmFw/b0M
UA/YEprZeFWXjZO9VgS7KaOwVyN53z+avWLnaFEpRdhZ+tgXEGGOT9AT8LUkIL6x
qlpsugBMaMFRmNHJVa+e+7bAI8682rNCSldNkNTzSF9jK5ll+bMkQC++S/YuYr8g
aUAVWTXqO0GoNxGbDAH2ynrJEgONGWjn56Q7nQJHukb+sk87ry9gh3lj0NhIFtrx
UIdRiVuWF/EPO9Hja1Xugq1mxm0c5LKi2wX6382AH8E6G8RYNu5+QO4hHHNrRB8T
GEkFYGDD25DMJHHBOSggGLLYQK+2NEooPA51cLAmzcyW8O1TgxZLjw1vNrldDfrh
T8Y+dhX5G4/Erh7+fVtfPBjp0E3tfXkrT9ZaobN35BstoKPrz22lwWlLj2rkLy9/
yCGQQbG+mUu82iZMG/+K8NF+fyYzTW8lcYXkjxQQoekcmkYfDJjuoaaHVUxkUXOA
pvv2genGtgO5E5+em2rR0Ki2GQ0SXYCXe51RCDKSRnPNux8FtDLEkEaQLamn10sQ
rR3iowxf4RptDjoD0YR1qvaCDVmDPQIjOXcKep4y1wMciatVskERdTTTFqdfjaFr
o2VUbP1t1+hRVa5SgN28yM1uX0yj7QbYrmSFHRe7l8OI28ZcWSWM16myBLP9TKLD
Dyi0KK5m1sGpmYwAy2IpW/+D3hwuGSpadS+L0kHxgfToEXr6TEiBMQfMlWhULs6G
nK4MbD5pdnDz0+O7rgj2SL1xKzAw8Cd5l1H+y06TlGMnNauL8wYaPbMZmMulh8T7
uwzwrlprAGb14fWSVkR7orMTEF5odbzpigLBdwrpNfVa07MvRFFPUwtOdmh3pmnz
Yl0CtWecvBd1JjFxgaGyaHdm6GKgkjlfrcyRHywNxQLKkQ05G8qZR6o0VvCo8B9s
a9HMvqIF8Rh6Sa2hnXWygdEv2Y43yzx5633Cpc0Y8FylK+i/atAT0bBxeAVBGgKW
45RW6+Bpj+leudLD4ckM/aej0fGCU66dzQBy43R+bedszt1H7og1+koAWcOM+mNe
+gaOat0JvplR6BwmbWkxsqNYd4gDD8mOm7Bhlic7fmnig88ElUp1+cuYGrB70D0t
FpV/qQlUy1S3Yhc6/bnyDgTt9kFmvXEI5DmzXwvbVY7cZw7GdR+tov2h/o8470Ka
JU5pJia2Z2BTjxeNKCDmTkx3jotTj7LQOysc6WOVgIZ7IX5zDuIIFzGh8qm4cKuD
CjDK7xekoJfOCPTkYYULNsLyhOIXUSNkNwgSifOwsLFQ9JRDOSGqy1g8pnRHxhj8
btrXrPE4Yju4Zmc/vxMG/UrakkOqutTRlZhm38nC7IOSfwxXG+nlbadQF/NXMyKZ
uzO8AqxMlHdr3oyXauxR4h05hf/ue5A3fTuDPBokVvyMbgCi0A0aEuXM+0972i3A
uNDb7HOtGW2mGJlgaK7sD9Yh3uCuMacy9DLoFqNP0GTcSN/MxpB4aAxvA4ghDWeR
bWw+KZsZjwoxTYhH7rCnrJOPnNOXypI1swUVofStGauOQ+NT1T7Ji5XameScqM51
El2MoaB39gMRTUWds1H4MipOeUQm1i+dDS6AGfI4r59TsPJWlnYQCuwbR7DznvpC
KFTZmz1X0qbwxX05ZsI1fzZO0BsfqfSOb2t4u9OrSPxvji6+l6l488npM36alCUp
vhY+XXkmURSd2Fs3T0usWhATgV0HcH6cZcPdXESPb17Zxn0eDM2n7cAPd4Tf2oEE
JtLEDRHj4ejr+clzUnOCOuTtHbELyv1wfAqmJTehWJumwee9LUdo/cs9yEnrLIbr
gJqHEh2H8TmJf9lmYOh3WBeT+2I+km/Jyz22DmpITxFBqp+XGyxj1JcqPMysWGOu
D6azCfVo/dLm/DWs05wdDB9K1PdRUAaUVpJLlPYOZ1Wr+AR5mez2H5VeNRt832M1
GSld74mA2IgsdVExxSzNsRRS3f8rNo8aLw4DOpHCjVz7/qaK/hjbmmLYmdc3Birj
XLFbaYobqs3aiUsa+ft9t5KN6msutTddHictY+Mox+THsbnqNyBmwaZi3hREVQHX
fuQSRYQEEVb0GjNkykD9PCJ1rpuf5r1LLemPVqFEYZGM4XrHClLk/ZHczhU4Ct7p
/YShrnZ+hkS6b0mx+71GbAtw60NjMcmS2xmJo+0G+tbR3oHSEQVYc87LDiG4JTeV
kkzQXnpYLO615hOLbNv2Kv1htmD0GVJTOzmu7pzHZRnMeIvPPg+7X8YonwJy22lb
7yWD+X+pgYeIUg4g1gUaA92/FPGEx4+pCxR0vnGSt5DKSQDtXBXCOpjZ7y1Yx5d6
0s1kUrlTrPW/lti+medlXG4bpVMEjvHTIhV0HuAUDVTnasKOytSRKr7Tq0JL6DSa
Cpy67G7XwYHnMmGp0YE/nJmg5icHtQ4XgI3RDBmlG55msDzzd5OY+f/WKmiqJQj3
PyhY0GPCY6dzL3PQSHvuS5yBksxXuTFJ1XOD1Osym9m7IKgxooSqDSSqAYmgKNCl
mQnvjSqKeVI3kcIuGxiPswNis2MauEYa32/DY42mo0rekg8YC+SogV2L8gs6+ojL
XjZloMwwGVy5k6Kbg2ZTAtm59MQrk6KDNFnLedOhaPcjuXly5tPfRntYvccA6GGo
35jBf7M5bNDsM51DANNu//LovGIq3qbQG2S3ZRu8ZwmDTJWdrFATJokLDcmRKLKI
cDQVHRSZRwGgm+FZIdKbDxTcgrEr8MbacitVAN5eq/4R3uedEdxr9mQio3UdvKG7
SWmJVnyxolUaOSZErf7hDk1IT4rD03geOwVobNOt/gZzX9P+ciFwU8Gu/3LY8zLf
PdvyA9B4ibt0PnNYVjPjdyrkyylDmXqETdgc874UzgiSIroTE7dpWNmjApAdWfwM
zQKp3cWKYGz7KKYxHj319/0ONP4NDqxwRCR5+JfEWE4n4pv3BD4SYvj1DfKlxj7k
glHpf/6ZKfHYEdZ6bRv/snz5hFYxaSLgQmSnBOsnewq+iu8uF5vLBZzr5fMFP4Ia
Tk+cFZwtN4r+0HJ9QJ8HfrNE7QjAH8ICA8U/M+/neVk/h6t+Ca/GR9NDKyTUSC2r
obMHUykEh4YCn3UQPgpiFI7aTS3ZxQvrkxRucK/wFC2RhxZqrgC8mIq8pPvVk3Zo
4eROKkfC5d7e5+lWzBhHn9SjyqJBhmrpyYLcBCkrUyoK0K2ODUocCTnTTF01ucCE
s43HkYOm9+TI/v3BWMm925Y2CtpCHqh3hvFqMtt6TNA0nX3Fu7jQNta4sHlA2znm
ScvJCLJGMpJPDl1KE88SXikavQtP5tPUJldggD1tHD2kQCOE4M6Su5SdjEE8aswx
LDAN1NLCDWC5wz5NsZkBjDmO0YFqj5ctWpKhOcxueFx85eMbCCNhfV58OKIbExUa
eyos7B+gZui7tsmbTcn9BCe2f3rjZLpCU8AiLaVbu/sCcBuMh8KnmzNEsUKAe8Qt
JeXXPwvY19S+Lh32gRMrBRdhHruEQmCyvAMSpBN6Z5hlSUbIj67oBajRCgUbzriw
6AKxqPr0DBuB7TiKq2TuJ0SYYCehJlwmfIwB+5/Xg5jclrTqjMP/JbMAYqYp3rCo
DvLLa1zr8Yrl52XADyMVYR6RkpRc+N8RuO6CQFn80pByhGFQioKZ5Tw0zjK1Z1Xa
h6TFe2W++Yl/6d+k44582i93Uib2U3f9ovFCgLbjMyRQ44foGwBYZfNtJHJg45pW
hAH5BtRGj0V1MP25Rz+uVxIMF4f4CPkthIWKGvmQcUBrnLyFeQ46JLI4GE9KNAxA
Jvvn1Uv6trDP2M3jmdhV2uzlazFTo6Gc7McBfYkMabqDwxjyuPNYzFLgUwBmA8Ns
JPc3ayIE491338WtCQlI67pISjzss1NICAhGWH+nfc7UiOu7gr+dj8Vh7b57nh8Q
v5eXETx3tCM6zKoAv1xZmwUMTlBADc9bOI4pWBkphl8U/fDfC/+83Wm9c75WJ1S7
S7yX/QxzEJHU49fGEX96hbHJ5BQTu27HiEnWs15re46V03GJ+etobXhN72vasi4+
LiWCmGiHCk9pk3VDaC33Vt2hIN3DpMUNLwRUZsMnb7hx7G31qtFYZOnj4hy0TWtM
AB60ip8mscOPztVGpuW2xDdKQcQDHhFu/UuiiEL69Y1kJl+dTx+2FDrV4KJKUr/r
njb2kjxuGJu7ZdHn6YFeHUKznNJvojSbSvOrRSlpI+L5ISCsDmEPRq7HfYCxD59z
ydsR51sFcBjzk1X3fi7iet2NRufL9IC5AwSlOw16llZmvJ3/wclzUc6BWUS0qMT5
tvK2ev7fQKu1Y+I7Mcpj899UEQrUZ7QcLYfHTbHFS9y3kqxwvZculDuO4WiTjReq
3bbiEzxmx5ACKr1YwqbthTQJYK0oZGmmoxsbAScL4ti4UIinJWfW40PW/f922j+i
HAN5oTKp3EG+1dJynhoDDP3AGj8mfEPt+QuWsJRmL0FNwxObg1WNV6Jf3MU91C8B
VRRStEmps6X03qm3+iBl7uTwjz6v+s+/siutEFYNyx5tOP/X3YlvkXV8t+FoLEFp
Pnh+Prty1LnhKHycNd7IuUCOJ6xtu7Li/j9mQTFQHyEImb318mP068lOC61pSFhs
wqlhW1NyC0ODljippjaAUUgv73lqv16UfzYRUGCN1RTqoi2+4YmIpbbJY+sJF0DR
xRyT3wk6hzAl0Z+vZwgiMNNibVnGOnwxwVJx30U8Y4DWCMJxj8qEL3TUFMOpoqE4
JrrMdfmdNyDAg0XRmoxkd1yiJvkMhv5cSLmueqOiElO5EjiWhr2rnjjhmYRx4Mma
3O+E2JHGEjh5CJeFqJUVTc0ElTHGcHMt6wpeYDuzAkeXDNeZZ8u+UB4vOP4cr24s
loo3USmjqhExXapddyJ5yBLfxiONdagFghq8h/Ecb/P7yELmPuTAIXr5GYJnXpqe
HO/k4oHtRHNRLrtfulcCryL+8D73aoDgsMoc1q7wom5vL09tpi3c0REFN3ZbxroK
XjgODbJO5fN/XyfsZ3zFLbTLXwLExuWaCtEaTGVKT9jPzOHdnxzVQbzErgJX1ogG
j0DtXRCHKShHSlF3WIz2/YrJqtTwvj8O8SUWKgMNVpuzNTRQthfRWx2tdM02Ki8V
2F7yGkqDffHOcfvklBM4OFzMJIfEy15fkGTutk5bB9IUOnLSB2FfzpQrOjCVCLL1
Rm4VYFenmcJTeiMWgHH0rluoBbtwbkE8gdgghDXh/Wt7VrIeqOvtIODMed8xitpQ
gPV65o1zd4unToxeZ3Bv7sSyyZlv0BKQi5BDt5wQoGUhn2zARpWRl83QEcDyRTaj
MrRxTNtfINKLTwycVndYqJchGiK+t/oEZ4nwHQ+lbJDPPybef++PuT3fTp8QoRn0
q5SzNZ+onSorWI9m5H50//U4xe18VYBDSBlOcPDd2kQDTwEtfVVLP62J8h2CRE+v
eAoxErc5pPuSSZRA2YQJ1pGKpJ5MF8oKtFcjq0ryajvVkNO2a/64tHAlo31JBglT
42i4hMwgwv8yC16U9SEEuAIkcasWbzW2OsgpO2wOwHJ5miMIwOUGjtjtbXBQQYJh
iuh1Cdb2S/7S3klfqId1ty2IKJR0mwW4CKvJ0SiKIB1LxNKnhuK55OpFihZmw4ga
omyB8MfhCTO5Z8uQpS1/shYxIt+OQuileQ0zczAUtFbT4ec10dbmVyoLcvBasGeR
05R4HHw8Lzyc7bo9hdq88a9W5AiZknUsYvhT0hZkM+9j2fqbaespqARNW0e9CwES
Ms52qF97wbC+NitQNfmMHz+qv5Ao+lyoi7nawTATuDpH1SIjV1q8B8qtRWlF2FUX
n26QCRIvy+PiHt8hyr8a7REM/Hz6LBXjNO7Kjkn4VPy93NczMFy5HVWNKL3FZAsV
77XbKkkH67epcDdADSx6zJSzJ+fp+UuJBLv0Yx4lHCmywkSfdJruPeICGNj8V9uQ
EdLvMU/4g7CzeddB9dNl8TOyYEJduC05fvJy1dd94feBph6daWExYiiBTlLuCArl
iCi2p2TcTeWmkBl4SRf07fhIiDhaM2/5WQSD9lTK6DV6XL7M/NmEJjRfTryHOJPU
GUAVeAoztnIgxY6JZw7A6QVjGuCSqHxCchJ2zk1lezFdeKpikby2pkBqMdEghNBv
AswofUvz1e4xnZpul6vW+gkT9OSfLFGRjK4mhuwp5CcgxBe8nxceqGZ29GKLOH+J
Yp8aSjHKbrDPjfjRJ8TsVKa+weR25rr+ZvpwW3cOls5zLQcC/XH/9xBxUf56mNGg
utTmCYgDfOqQpccfnAR9LJHgBGZ3Fnc9rx0O+PJL6kg/fUEY2NMVxfbcnsL31aBG
dDSnM+B9r9qCm1SFrcIMZYcWutR6QIsfNQof6qJdDHTRNym9JtON8fOVKNhn6bQ6
gLSnxtGzmZ2vZ2wd7vjuIuA7+neFehlAogDsX6stnCRC5Nbo1G1O5uDA2HHZ6G/t
tZjtF8Jg9JT9YlsC1q4sTzfS5kJnhz0Y5RPPHbFgJf3+hthH8+392x4UC0TO4xmf
djF/GOrjR+zBahgKR4BZhKiZ6ebBxw2Z2sitVfdd2gBpjIvyxrTks35nbjPMaLug
2QEBeSff0NNrhDQpUp1m8IC7t95R4Lh4R4T0Qi33LUCMNURHOILPgT8+TazqOuW3
94z4Qc7cpVmJqhQBcPOdt/F4sbmVLawxDXdEgxk4ZljFtF0EBI9IUiRya6g+W2xB
7i9jLWLsrMX3M3/gmdQrO/+plFO4Y4F5M/NZDnbx2KEkITxM+GT7DHj3xOjZjI0A
Vs02kmRnCi0pXibpmMFJJ+u6pTP9EQxB2zIHnP3XDQ38enMrbFd5AUn4DIpDji7R
4WT0Zl0OoT05scPanxA4BQGHLuNnJPoqpTKN4C/QnOcyx7dbt1XI2JsLtzqt8fax
9oAIbDbCvRoPGRfo3cuGpHlDtARaTOOs8ztWcRBqfcLt44a2KMrZOiRZoe/SL+bP
I59DvQFRI1OO4lq3ch9JLn91SXFKmc0ngpJ1SvmWXQOJv81yfmhkwsxuayLtUV/7
qaBCXpG4XUK9UMBgbOy29OZuCdxIVGeiAdudolfELrSIRjQwUOoRZita0eHXQE3Y
THS3WtjSerFm7BcnhFMaFii5q8bdYxIjELRt4AiifK8AJEh6azCootN0ioxFnVJA
UoqzXkPuYPGq6h0Yydoy8xC3EvQkvWMGoj4i1rnXBeRx8FChga8cMBUcZEI4ZwGs
yxtMn0zRLmMKiwSCexZQb2+pQHqEQeYlrg7jAe0VyHvrSwqEdcl03PTTMvDuz+qs
YKvvVZ4HWO0Q1jYLzO8L5MQksvAChbi/Wzo8Eq2NmlDZPevoeLFvZjtrn+JhVmuj
L7YTaLLWcZ7+haelN3u94kEZ5/GM9syX7mjmG8xcu5B8ZPO2sZWluJ6Wh9QNr0y/
2KjOnd/AGNtVfAzcgCzLY10uhrmDYXSTJtcN1HjesvYrJ3IPu5Lsg3nOhavuneI9
T1TQfcrBnkl90XDWe70UVEPaZm8iWPGxXrjYXx5zeXeWteT0Uh6lx2bG4tPVqVcc
I5yMhp5FHzr/1b/bG7tIvRvNLbLhT6aKE7wMIAt+J2lXKcggMgOpH+A/47zUnRqy
wwGvrvTwEP0OObdbxsp9Zz5PTnAePsVFmXua7dJyZsp4J+NJfWWCEWOmMy+1Qd8O
b2CXLY+0kanec+7uzt7WwTKO1//G4ybytBYKq4/lkA69J6+mQvsh+BiSI9sgvJHS
ZTgwhSBp3fYOCVSLTZWcYfDZBKBqttwFwbNQvwcfXl50UFngyG1qh9e6vMjbwaJm
hSYay/WgJOwxVsq7t1VYfqTe9jgyFo4dIO0VTt+aqs1GHxI/QX8eEXoCUT/JyTNz
p8Iecxp6aJDP7uftBoTUM6xGDh/gPlySX1eztQiUWz/W4pj8n6/jvj7nj/iVP8qA
13027W8FAkIZuqXSuro+e0OIzisR/aJowrdGulZvf433L9C1kGW3IJxevA6Q40Gs
9Ullb7GmE1Y5S01jz+bWcxiwpcbbP3KbbyagcZochLVto+d/+FebxLsTTmNchNtB
g4Tja298EYFEmDMi7a+ZB4l5g627BliHuFHWDiluQ9vbwWrvS8ANL73od4UyiAat
m3frjmkarWdFnPu83/6JWU+7wJJfw0qtG/Wuo/MZbGlzH0P5dlmxeSIu5a+ZoKfT
fZYI5ElSRSboHetn6rjiNtWguxpcvYXXLQzhnS+TDelTCU0dvHQMk3/ZK7kD+hkL
TcaT/JMTpNJRXL6z+/5pGyg7oZz2yApIJZv4xPJ/WWigl09r9jF40KslvOKKXINN
afrwEbxjaunOykngAFvN2z7BbHlUeN40A7r5He1j7U6e0kNa1xF5WjoENt9eNjFE
jPsux2KRcPWTQmBG3GGwUg/FzMhtc1xLQa3qUiGcwPgLLJq7C/oD0VjiVLLV38Ql
KgWVbbg3LXlm9xn0o6besqS5g3YQkERbGCchRTMiCrNJh2ukIDx6eyRRb/7ADPPR
cRe4x2LHnVKWW2h37mbvXLO0Cv6YkU1Pdzmxnky8Uh4dhYe1ct1rZPURXvn4UxyN
goLEDMgMMQsLziceXaK1+h4bpkuWCygGhnWgIADHSuGMvM6pEwoeKiuO/bFGSqxZ
mDSB0GaiZSfoE/btolwb5qpSUmdkAzBW5qvy6uyVRPDMY2q0kUjp/zRFIVdDbzUr
7/AW7MdpdxcKZ5JIMh2SlslDTOQZkjYFhKnIJwPKtkzs/n1cGoZ/HZBbRqtSyQvn
HXzeI8rv9bZoX1Oefoss1SfsuZeYVXN/F8MFr4mWamIsgSUEnaw7J86jb/d++vlr
qD9IvFuZx2E2jZAWA55FCTyMVRWL+V/r3WI2kyAfACbxxZJ0F3jLx92fysPtE29A
8nazaHwWKpI3kyFMqX6aNpmINhW8kgUN2g8nEp8CoLoswGbUIGV9UmnOt+AU/CVW
CA0qq513dEVZpDh6dokInEZGGSpx0Obu82OYk4tlYtAdPjFwTCrExiSYqspfEi/D
z6pquczccdlKka9DQiRP9rp1jWgQUJuahh/M/6jcEqkRo/RoEh+XOzrIUJW8n70X
NQSiKa40l6FtMz9ml3DDSpafyo1WHoR6HYA5HyjHMDxcoUGtzYaZglz+kk09OGLV
3oLart4GXoGi2EBOyTISQRlF22Vekknb1G6RguNFQxAuUl8XZ+VmePYVCLoFQwog
U0VVoxEIdU8M6UVMNCq1H6+o/h2gKjiH27JmW2jauB/7Tjd3Hx7XYNXAdEhXUg++
AfeG8ciP/X/dJpCMOxN5DFPOSOg2Ek8IEsPHQB5z8aHEimSp/4JNv+jvsWGGcq7w
nUQwJeAaQZCe8TV/JfUfzPuhxeh+Q2PeAPRgiiwy523e/p2myaYtxWOiPVPav+kO
qWE3Q670K1vFcflSndxkOYBpgyT4IFxykuH7M/8IqQQRQF/Ch9dPcW86XbIJHAVg
tMAThatEjSf3WItZuwGH+8Teb8nsxUJEAq5fBhTLd6RKxt8jk4Ii3vyKldNAyARd
3cdyUUuD95YVY+Q9rd9eI9KeYIJsk9ygTYA/MHw+PBPKzlFgqsKCd3bUOUWzub7l
nmp/uFyzwQxVW0PdcdyG6uJPtHKIfjQaHLG09Pmaw5ew6VkeS5zbv+QBePNabjzo
1nsSRtkb1FGNRAN6JDp7XgfFOuSBpBri3H99y/Oa8PmLSBwiLX2gfrmKv/l7CNgE
LVurw1wYSt/7WkuFQIaXBEbWtLxwOTWye/GwiL3/0lHQxgND0l441ZzfjykhNlXs
tLFSLEYOa49uFfn1ZanN8Lg8B09AiMrNPZQmgxidXDz5y0LMvy4e5Vwi0bcL5FAA
HmbaRuIxZROLXT4SH7AJMPStiOxOYb1Yn83G8Mgd4m9C5fz/L8asScF5MsrINHK0
t1JzzPArVnB3IltAr75V7VI6xr7Cw5A3Gm1sHLos7RhsaRW5jzthEpQX26wAV/Nc
VDnPh57Dum8mQqdAKamdO0m4zfTcpgb3RE7Eq2bJeJiXt0adNCZ76ac18kGozlnK
SfAyWSPpfoo8v5IFonGvQw2yL0xPAAjeAUHyg1V/BGweahG8Q/AZzCMPhOQCo5vk
ya9QuFrnc4+SxlauXIUWmEhqjjl0SHRBNFpjQ93+s+86A5TOzIF9iMzgZ4XT/3oD
8QcpfBx6rkkdAY7eWPQaNBc3FI0ix7U0Mm6xMh11zfIC3D5ieBDsBVSKesi3Pz5p
dXA5R6m1B5h7Zl4xM7hdGkC9MYjk5sjm1hGJ/nAKDvZ9YqneyEmBR07DWJNogl4D
s7nzCPItPGINfFlqHrXevu/ICycc+ry9udaB2S2CWFXNrKo8QNXBVCQVm3rheKXW
ISGMc9N3JUqa21gpDry3WBmVUvD1syJij7YcOdpK5ZHQ/elMGmuwlPtsy4RynQt9
7RMzyh8i2umFXzigpzEK70Xq7apgxG3C54GDYXJyAJKKINufEuPOwkpj6bFFVPFE
giYloNIegB/Fo4IR7kXOrKrJNDx/NmwPrscN9L7vQfsCfR1riUF9aZ5uNpL2seWX
kqjOexNPdn4DsCnmt90/MM+vkNBUPJ0JzCOjoaURIUtoVPsAa7UAi+d3MaYgGs9Q
r8Kh5Icg2rmjd53AYU/G0ZOPEmq8ASYPmKWPe88b9INAv9peUglRXyMKf/2mR9EU
94KkLIfi4sXOwmI69Y2rsNb5U0GIzA0vA+Qy7LDAr30f0wg9WxCJBNOe5b8xhWjV
AGFgN+cD3HHf3ELgQGJGrAYnDHMSYrn/4cR9LBepUJD3kqaurnpqe6cT0rDjqQ7E
OXZdBilZGgy02khF/kgXmjaulz0UdRp/2YTE/9T/nbx35Cc854cpGK1bnFg8vUwe
vYVGkq4qSphOjaECSh9AnivhK3+6zTJ6VLvnohH35dNqtzwJracbDYJWQhsB47Da
bknzMAWZ9RXrBCb2FR4llWPYsVj/jfP8aAxutn5zwLeZa29d7bXsVqf9vcUtOXu0
yQeLMnOnm5uTlsIEJe/HooCUQ0vmlrbDwKdPpeDD2c0uzhRnd+tbvujXqKcsspIz
bEYWzIxzkzA9qr+V2XglCQTbNNOVjRlRBAjGbNzZTbchCub3cZXCwpIv9KhWX/xh
KaPjJIMZPGd7R2Ros7AEIK17289SSIRYzplzpUX5+kwyNOx9SdjZgZjZVfLNHCIe
Det150CGYEKL2/9GhoUd26D4U8UCMizJTLG7YyxzyfMSuySzC49q8OwFo8HOZWsH
RU/yzZPQPTwJ6YzPlPZmYI4zISPnV0+oPn82yu8akhI3deRUcL9rTXpw1UERZGVm
Xsq3CmfRL1aZASdQUT0d+XQuKcFDG7biDxAbUFTVhrKX8Q+lqWo+WehIjAkNt/5R
YsT/6rJta99QAmarTwZrLbFwgc8Fk1G7QV7yMqKFXpJiSQVjY0W0dmGSYBeR/xkA
+BSrYlf5mcehtitOi4DkxUGClCn5q2M7ybX+XddosGmMncliRaxtDj6Q70rH6V1V
9ObBN2SypHtyqvWSxE/w+EJbdwiS5vZo6cX5jwqP4aP/VHCijSeUJRPFw2Um0Upo
jGYiUlvJmksTug8UFD3wWy6rNnixer4VAZCUdayp24bmFs0FazxHCfcbixbC/iqT
ruL4CoJ8JM6/5c7XzuWsa0ECeylSei8gkm4sBW6JOZEIoLNd1GYihsjnVJLsXynT
WrqTSUyjwZwRUCqShEmekigQfukwvkv4BrN7lKTq7IAFiDV5EWL82CjGuWNPYsxG
7jTmQwRlL3HYBGeZE3sBQW/YwN4TKH1B/TjvGCKBSRZA+M0IgMWtO6aQYbz3oURt
bmOIkKAxFFpFLOzF7kyb5tc1Ey7to8Vy8BDD6i33ZSk8aZXzIL6RtvB4ig7uwZzD
kTDYojCc5KKFQXuHjupMjVYqlldl5jnuYlQHyjV3PS0V0+eoyYoy8JfqRAKZ2i2u
IGiWc0LY4b+/ZqG+ZuS+thlpPJpOYG7V7h+U/A4XpeeP1kS2gkCt3a1FMvu956bc
cxUaqnzeol+v2s2Zh3u3dfJNa+/7an/SsvtLp+e3qPi85DwvlvG2mdhjzBGblCEu
22DOtF+sBKCO/UwF5wa+OVLuzZ9oMJka5eGZgKE7lbRgXx1sHIdqlB/Iemn0SMJX
opyOMOexMOoHwMb9D5vcyvwUJOtYUUaTF9Ek7NqM/uPPVyIKbE+TxlGytAvYFNY4
Krsn5nSDTKHcJPjPsh+kF0ErgMs1VvwtRRMCkZAP62vjwLwghwMynofQZeDPb3fr
AfsIAfLTEE0mzuAHTEUkI49Ct9abaQ46X/fQuyehrFNe9gsBJWiyTL8ArOt+2h24
mbOCbihKT7rUHPQ+2020D+2bqd8ZXm8lNHlYbNKTQyyfw1IP0Ll2ezpJ9IRE5jzV
fPsrAfpnhJcBhbN3qXZu8WS0lKSH9B4VJwygUnyj4AOAd6vvXQVjc7jO5YyKr2pO
gi8vxROAHPqWI1wW0oRMDqY+vGfhL5cxNNSYgOVgo2AO68RpjBUa4+oRkuSLMFKn
gEjJfiM5Ql5ZhoCZCViIn4Yu/twytry8zTXa6Qx1MpMqCiFUKXIsrj0/bQQv2Poz
rxhLGlsu17Ay3nKEfPh3mbDnBYqU/YPSkZ1By6x1IItrO0ZLIGgTh6Mky5Pzey1E
lcX9KbXKtQq727L+9jCY/4QgoFbOhL6uRhaYWHxLWY3nJnYdrsu+IxMoHmlyr/8P
bg4peFU4dKg5QoeIDddaY8QlIXP0Wq1qOjxYHBYxh00Bwk9gYWRS4242GGQygP/b
bXteDuBnUJjvsry9pCcs81cPFnyyyWqla8oPybQs/Kj6Dm1CImVM6s41IqO/E3X0
Pv62Os6ExXB0NnsnH0Cw506JoUJU2fc5fshrwS1mGQPlvWwllTUG1ynHzVsiVaVE
ZsprTaibs4TC5GlGvQ/4o42LeG5GjooHNAnu05Pdaja5T/IDYLwDvO8cF2KQg1eq
5GNioc8/PxWBzStYfQnOIW6+nAUwIGXfjAs+Tyq1Wy56OToCBl90p0mJIUii855M
Yh6bL8MmKk1gufOTqInrhaihpY3MKlM63PibVUQ46awLZ64kY0O1T/SRdUF32gRx
TtqsU3k0A88wJZWc6da+lJJKXl0ronnynSqD7UhWDljSN1m2z9djA3z5F+G7z1+X
G+yPcvUcJcA1MaIjcv+rowYqSZenkvk2ldE2JWrhpwrIB6q3KnciVA3dPPj8ekur
2vP7Vcz6xC7a7IlL38q0ISuxsvCCu51nRsS7HpAy7AcTAXNLw1RbA4PYgWDwbRd8
SuTA2+sftEFZGQBCW+mrs+6ZUXpS6vMHGflIYj0qDL/eTuJ0GXrzrDDe1TdGfbK1
mO3VqkV5isl4zWGj5SFYGy2rM1qYC0iDDmlHlufUbXMIaCEeFbOpHbBtn+vyZeI0
LXZMaRo3dzp69e+9jxn+1nQl76EFjueHaJCzG30FTUFb/WdTb3ECoa8+QlA6+R28
ztXvt2lJZZy0QVbmF7SzZrnmOucTmIbiuQIioxsfNbTYKhbpBn/o0wsMRGyg+Q8h
s3TjpzLlIXtAWnj2oKB14QrGlYsMyiI2aj+qh0HYrkYpEWFlLYYzCHcD2x1263D5
VIMJvTTaOYNKzmvCJt5u5HqrdBAizmJLVDNSPwEWiybxVcPfy/hEtz291X5KT5dm
MXFy8cqU7/rMO7Xb44+8qHC3c3eO95URkmg5aTBCMo3hqUGtHj6Sw6Ik3KXYxXam
ADmULy1dT4eXPJTCdsYHayg5hmrYXEKeBY6Rwj7QmGKPpPtP+ZrVNu6GvFMQCE8l
TWecdTmnwUaH30Jn7g8vkQj57T3GuaBLQHBvcAuzqgO+zjQft9LDqwGiLQlxohYE
LOyRF1QWd57Jpu3ZkNvRNF3uoowJ4n3v/P2ZrPq5YPXcg/t3yDLRAawyYUjPTEYM
di2C4F8hJpM2mAKKV9ZYV8290XVNYX1GkHrWneUu2rStHbQoOjgPjLDnmC4+RDJb
4/4PYet3Gh4VkE7NPIQIz2CfxXGcIwiJwOnQ0/e+u011nnWHD7Kf3OG2U8cb6H0a
HZCY3rvQh8ScrC3OuPA+m5QrS1zwGwcYbJpMcbP9CCgmTJM/cVurDhtNDJafK9zX
9TaBOa9bvUrxMuO/MG6vab+yUmUjuT3/Ld4ibTN8xoeA6CpHo85qN9JD75slk1kE
zcWRn6TqABB3TErRwyKIUMQqHUb1uQvbvX74bMll9ky6AnhMJogVbsAC27GR8N1X
XbXL3XSFIQLttjkMfMTI4FrAhy/2jiWNuD+GFnFprEzVldffLZP0ydX4ZhM5Mdfl
J/cWJkPWdeb/QHNw3kXTacdXCMhAv/JmRnwwkg62j3f4q6pVLSLyTaHgH8HtSEEz
OrYaaXbjJ/IszQmzdBTi+fDALx38dbppgFyHQkrg+dV4uJcVR90836jq4u/LmBlr
9d85o/kdeRu6RHMmVFJ1hAh2zkGjiP3FE5U+YFK8k6/1V48kCepUt+D/aQrSOFxZ
w9vWobWQ4V4fcAsxDTOI9YiTlCxYbvLxZXINr29DG63mvroNC+p1fzlEZidjQer4
1Z08HGnpNGIEpd0uyms9QBNqvIqZsstKUsAJ/YDnu1hygDAoLzTjUt7klYpGIYwf
ef7hxinbFBoGpRiwoeafeDbKzZi7urqQvwP7wgmX7mPMO4zMPjEry/qalI/KNCYJ
MBEBLyZN/JPj37qkY0UwF5VusRdEOTu3OtDjAYUqR/cQfvTVL1Fj1BCoEfY58SO+
+gMa4yYf8Y5GhNcv938F4K8a3kU0ODtF02FI8djfzHnt1aKxSoGZUS7wFk3jqHFA
wBfQ7FTOr8LLPFcw3GqUgcYmJTv2tRbddiz1LEvZW3PKWizAcn4qUYzZvAq0gbhm
TTP1NsdKZWBMsworfkagRE6ja+jp4x1dNDvXGBzAWJ8FZ32yRRdLL/ipLvBvXg5Z
h6MeYvEpEjoKY12Hq3RsOti6oM7HC3QhBDPAAaKYGgYHtJtYjTOwZdAPDasqUPmg
HEjRDflp/KCbwwzFxvCeDR1ChTFEb8QaHVYHzZE+3s0TTicY+vY5WifN54UO8Skw
FdwVaULRTx7x+r10vXNWSJOjNshWrTJSx3MLrHsanATAI3e+UXuHDnrcgVXlzF00
4XOfZ1o+aDmu8EFzi3OmyInkiQiKSrEN4h9pkTy/yzTRvnUUWYwBB7+tkuqS2beG
yQrFtsJcL/B+rFhRI4LkP1P65SBTu1OZ/t1JpaKJF54Bp+wm+jdFDhJHwhYMPYtn
/3NhcxsnffF+Jxcfekczba5VleP2p7tWEa0SpAhd9TeOyderU/Jy4mMpNbPdiZeY
baSVzJpFhMM+xixcQexFakP68wx8M9lrDed95G7l+b0bcGDP67seBSlB+Ku8cQ2f
iwxQxYKT976jOsnicVyZ9EMPk/6OULEszdoKROUCSW9m66GdVbvx/PFy1miiM3CA
VbLldcw4bVjBGhBF5fto/1hRAk/mvtWCzhxnKLw9JcccBH364s2gPOaVCMgs69iH
nc0BGYU5WqkBOjj14/meESL7EOZhWnvoovquk0Ip1AhKtlXtDgLCb/KlthfvGN4U
Y7q41at5KAaMOIcmq4WRZ8bg7ksheNje6uhImG6lT9TPmI7dnK31VGnVtZHJ+Mej
mYeZW9wbSDC4ddjvnDO4lVczGDr32M+KqCiCYjh/WytPiQ/fyz78H3VsAyvgKR7+
uXDseM0LpMimn+gn1I9ZHG3tIUBbSMZfC4RIbHB5lNh27Tc68kFEQhFvUsI/JNOx
vR/qOx6PUOdBmamxI8mAgn9zJ1bUwx6pR821WNi60cqDaP0OvVPuXX1KcE2VsL8Y
tRAsHvskQ+9vjWFrEFlFrl/m74Vb4BHbCpUTiKMTipBYiVxAmxSwdXyG6XnOLvVq
DkTuGBG7siNw98JBD/mTz6BNijJpn9ec04gkCvVQgnY60M5Rfeuh+YaYu+N65r1C
jtkm4p3vgS5PjD927tDtYHMiy/1R/bMd00n5BTQtyGorFa+C9JG4GZc1KVpAwf1t
xDPmlKMXTsjoKnLVdFUVkSNWndWWnou+ZEym5l0VrXp4zMDU9hiMe5LF1Lros+qT
jVrsnDumV/CiorvY/6xv7SVxwCcg/lAvN/m9QXboNhz5eKDQqhMoodN/7r/Y+VDm
mH9/CyvymZat/q4iYpxeWyJ3tf1QDrznSvM70Thz4Puy5PhjuUjrWwb65+eWFFJm
cEiIMhoknLez6HPKn7B/oqVq1pijNtA7DmhScm4TzhmA+9Fm/WMCgyKlg6jROyuk
yfFiwGK1pgzHyhHThTCszdw2l6RbdFDJk4MR4MwcefPfJeXuDdkBX0Ds4w7NVqiP
i7A8mcJUwfkYrZy39A47okkLYtpgeF1V2f3ufq6sYOO2VxM2OY3w7QFAcQa0np2N
PxTwtvDP5EhXBISRnJfshbgjGiLIJjqwZaZtXs+ymSEqLGbGekWWQ5ZkwnnL+JJb
wtSc+62vwkwXSmQrfYOV9+sEqOChwjXhV3468ocf+/bslO9pidueDJ5+yEinhQ87
HIMQAEK0yCqrc6Q45g43g+ibd/smrbfiMSpEs/Mq1JYyGGagFvWy7eRJyM62qOiB
o9ol/BstpN+aMYRW4LEWdehGliMlY52F2feScoVl9WGK4N/elFhgam98HU4xad2K
TFisaS62ZRP401pWfZosmdjwGeOWzeVZbVGOZ2Q2EnUB31Ic5/kKdpV3SeooseS7
qY6yS1gxsZEsgOloCkecw38k6FVeZ2h1KKo7X6jKwsF7dYMPCKeRn92KPn+3H2xv
lbiXMDYtSYDl9iwalrlnCXHql2r6X5hC+fd+ggFH20RWMWpCori7j5iVXjBp6I3T
hJU5SdK55p9SDL5EwVPoHsdNozi8BNh5f2s8cssK9t3XklRtb978Yiw5+gtEVrXM
70Iv0yjl2uMc79i0LU6/yauKGZ7lXfC2U5WxVUfMLE4sWlPjMDo5BJC2YGnK+huu
JD6wiYZk+tNkBoawwB6MBP3fkE2z6swi2944WaDCWJ1E6pu0aOYczqGFiFZ2xvLX
xk6tcHkM67HSByneBDRYvPDanuhUHp+BbF1phrXIiQm7/geh/Il736aJXirriIie
MUZPubHjc2ho6oJgWpmiooTHzf905pLaMHFEc9VTRVHtyqiJxi5R4AZL7XsRPwbJ
tTEQSJ1Rwt40oBJh7YpglvdyrJMrgoxe5p1qlZ+b2cHmxcqeOUy1pNAMhg/bWQlW
JXK5h2D/VxFfZcsMmaJXAJaOM6fMUofjRSjEDYnYQfbQklADFX9s/bi5On/Noe97
Kovu6PfJE90co+kxy2WzVgO3TVPAd1ny6A/HH9dnRDYTbk1Mzq73YHfbmjtU73kh
5ETPWql/FHM0VgIas2DlJnjzeOyhlESokd2xiqnRDco8SR3Lol3dotLXh0HCH/sW
J+c4aTRdz5w3pOnEPLx5nUKgmTp3/+sanbQ8B62y2MF7YULuOGnURWhNmPn3fob+
1ICfGf6GWPLHkrgDnSq9msKqBC2+FkWyzSKSt27BbrJTdJXFZwkKlhNOyDPZAHQf
MqT8z/olic25xy1A5bM1y2qboQhY7/cjOJLbs9Dz9ciNGD8Su/WUKyvuVuocouUa
EeUnIBE1Huork+MI7nN9msx+IeoKHiZfydMjmyi2VFtKhQuC2zMs8eQgBKrQ2QQM
TM0S69A78VXag3clTAZri8BsRKP/gu2m42lbO2hR3918H59t8hZKlMaGLH6oKd7b
RXvnLgEpalE4jJyippp1sjWSU7XW0mZwdXUmns7uRcYGIWBzM/mHbsQT75OOYIFx
FuzrVR004cIt+niCkSC8NijY2ABOAl7px+CHSonxDKyyDgeDTp6N4iY39FFWX7Nd
uswtlyEh5IYJyv2qWF7+RAtsnjLj4qctlRyAut25v1ueEpIhQFeU3VUrNwZBra9B
hY1s184qbkMRrSjzkxmHikag7R8Neu+Nx2jETgwBaX2WrwJKKHx/3KQlSycg+2gC
vydrGG3vCQcaad7WAoiD6c3CjLknhroRvv2+31MAwUxkxT/919AHz3mrggoZKDin
IyAMJkmQyPiyA/ktrVF/VkVfuAi7YAOrezsTd0m5PIEd9/IEPY2YkQ5Ed5V0iWWj
t7U2gKz/LdgpZZTiJ6zCJe5i/9WChpcYMi8HcJQ8ZZfnwNrPOd1n99cb8trXvSvF
NYzGP1oMVe1GSNTo9ZOnJtsoz2KarcYQX0dc+0QyZ/0QDdv1FPlqgzpOdYZDA6MM
c2Zx6JIKeeOLQhpBcpFu6AFmr1BLfQFGN/pw16+5LtmE3DxZK25QKTFhGYnLWWGq
JciDwUtp2j4Vw4jEDlH0bjYmbBALk9rD+d0RDh/yP4rJG5zXIJBF12kDCSS5wMRS
KDnYjFOGcTKUC24z+HdKpszgbqWzlo2Yrv/cA8VXBZfTmKuYHibR6CyJFhgl7QxY
O8GfN30Du/NKf/5K2W8ruzl0GkY9ULBlteHusllRg+lohxSFby/f7I62kiToIt66
L2eKZ5+8MJxQINoWi0DvZg00BIh+s2e9rnjmwwumMAfUs4+bOAVsWcVerlG3hBCW
/qUsDksPqpu78zBur8VWrQU2P2uVorgfZ+SE0V9MjXX7FTrXXix22VJGfszZbkbG
OHdTqnNnUGKsBgIz+Wp2BeEvYRAbj6RoyVw0mSCLxmQyIlgy/+PU0wW36LL3SQts
gM+1p36jIzPdqn3xoNjGdFsy7k9gZ0USrX92awI7vot3NxJIbhmtRqjsL4XgSYzH
3r6buyukh18SHJrebRW9a0LDbUf26W9G+jlamcURv9wWYXOS2Yrf08v3tTGDBHq/
KT7wNyJYwLF+Guf3yTS0EoST5sCP7JpiYjmHMH7GjwcO9WXFQkRuzYTnytm9RwMd
W9iSxPjpVQdlagG07pIk6Z5e6Yl8pGBNlBZYOC18CV0m2Kpmf8LeRhLobJsH4pbP
U9USEbaGgkijupEcT0x4XVTtMPjZdJ+w0U9S98/yotIy8mnw/IXe7nenmS1ubvM/
xmFp5aCNMOTsL3DffqArsveEfd6OpFM13dPqmOKfnZ2QkrRq7y9UHifZ57b1A1EO
4wW3l77E563HWhJv/oedA4yJjTw5c0w4jLFlWwLhSAGb/L+HNBqszLZS1k6wAxrM
YSH8QeOmjpFqJys/6a8e6R+7eJnSeG8Pl8CPxvK1e1nqjR/fpXVyI4X2p6KnOez2
R/whncCPrm5iOl2CT3f8Lojtxs62kzhMpg28MNGj1QbRyPtbbi432t3vBEFP0Nhw
rlbM57batypRY5JIbsfu2f7njSPQB+WVUye3cYZqYUxLpZNAecLt7Nd9OrgF/nca
BbGUp0Le0dYAIjAJwpXf5OlSXhYKEaKhtOasxw8OHpBLZ39SIaNKSu4cbihpzUuX
NIEfjzq09qR/w353mBC33JxoSl2QHhciTtLMEwQ6fUpo3sficdW7vBrtzd+ooaV6
nSa20M4s26OqnAtMPTB1d0XqYXOhev9INcocZau8ViSpo1O2+sJvGMa+LCNJsPe5
VKBGjzVjiDUKLLDGe/x5nPM7ZPdCDeUtz2Vb9v3AbX0zrCMJAVf6j7+l5QZdGw3n
9H9wQOdOkWhIzWNtea+cfnMSXLDtMr2I2Ct51bAS/3rC0Kz6ePsROu7cIr/q8krn
/nt2VPjHGbm+13WZ5jwnrkOUCq4vxyxz1FZ+OhK0Xogae30qPN/X+mQxoVaAGjsy
t6Pdw/SpEDrNhNvTfErbyFkFPiMOtVb0NQNdcF6yxPgCBRMXReIGQuwkBwiESmIu
m2E/BcdsmLEcyNTLBlyK0ijMZwFeHAK8dq8nykZnNlsQ36JOef3FdUykFNMa+PR2
MxvKHffEj9NiT0qwcZxGq03f5s5VCs9MwZ2JkH2CyiMIV8DGf+LU9kAEL77LhJaE
V4or2fyAP/fe6GheYB8mcTRdQB+nlJnDT2VQ+pKwDY/ato//7BrZfCsL6aezOed8
Bos7PEDmBldy6ZObzFz5o9NTjAxFR4xzzmc04KKtwox3DD/fQ4+7mgJZ2HMMfFBa
VHncJ1dm1HMJDiLC/Bj3t4lYmzG0YzIZzMwt8eQRal1yc5VWiWRI2u4wHnY0zw3K
+Ety/Zsp0IKxO9DJ9GnrpFpQY2JkXsq4WkA9akAtCdxrn0MPtE0QBJBMqP/nMJF2
7ny+rRw+6EJ9e+f1Lg4b1kLl9Uy2KYDnpzctadH/ZrTnRKhEniCg6wasW4Dxc+55
uA8ljCEpt/Xfy4Rm39vg+shwUZYuTrOdSy3p0uBJrOEGg5DFw1WFqmcB8bxETFfl
5a2uk7vFYmoU1adkIEFN6AOkssCSEa3MAueFuM5WO2aaGTC1U4/3hOOhlBnHpmR0
uYp2+CfVyglm9DBGokM6kW4Tktlo2rMrohyzJAY2ab8YZ5Qh6j0DwUcXIqijyJCL
s5dTLosJtXFvhUNGmb5iRB0D2T+N/QDe8MxC4nAQGmCRVuthDeKp7qU8kpkVlgus
k5en2nNJQpGsSRXKkSDYZ1Xjqim3Pd8ZhLnLNcAM16ihaKPiUcTM7VtprQFzfC0L
CZhXvDbL+xSRisRFcUIn0eMOk0+AU1KWamEoXiLZFJCVIa8lHQsN4gRdUHujVCL7
1Bwq6ABlR/FDjzcMlKbvBMNwmaWiOG4M7DRDP5l0Tv5Et+xTsBzs+k3tnxKaz6hy
Wzv7pkxu5JvJmTJrKgReoU1Dc3ycemawatI9X1G5n2kMgqCVLFjpeNKIZYBayqXH
Y7fhsHBjOHjaDglw0iNbp2FRQs9x4fuFnZRquaf4Ik6aauVxFbmNFb8vrqmZ7bzZ
22MrDJsDBBnuVwVqpHpW0t3IyjBYo5todT/yb445SPUgpeR6t4HqNVUVlnw+f72O
R4mrtVE9oaG22X1fyWqfgJjbqWK67mrrtQnEHhUEn6Y8OghSNMMpGBO8dSvOP8kc
IHUXJqT0pbv0JQ2LpmZCu+XBuCK44Lx+cr4j1XVJ6QGZ2kOdZe6QdHCX3WEZRc+X
cVygykQvbqSMSpS60phKn6iCpTH9ymxhJv24/fHQ3Iydq8nYa7/hirbtSH/sADNu
9Wcjfnq719pP3vtcgnMjn77E6k6L9wNV9y+hfTEG93meTl37veSuCMeZd905KKTF
APuYLWKoS5u9GPHN46xLTcVoB6Ku0QviEQuZFWJ9eEqMwuYUcPJ2X8pdJ+URGowv
cISKyBaE7eDs7RkBDR4M05l9HTK/kCVDKx576RgsO7Fw7tnYo+GrieC5PBP3cXnT
FDmwDKOEYAsQ6mUzW1k6VUykQ/JGl8PZzaeQxwFvjxdXfCHAo966y9oL/znwuzPT
1ouraxMjdv95OeY5tgZNS47fiHiyGIDZmiADVKruUz2Ehs7PNZpLogS4k72/ARk7
K+7FaxRhvrBxlRw47/VtOtGXiKBk/0TsGrmwBzlaBuMuH/AHlxiB/HGrOqgJ7ZxJ
iVkKfKsmw+6mckT/bLYPpHsYBYbFSedn27Y2y1/VxMNkrUeuXUKheAfI6T7NY1+L
S6yQ1xqfNdprRbrukfQEN2g5l70Z8si5OG5hZ2FWOz2uR1OnnckywhtHL17kVY0D
X/3pWehxjq+eDyC2Nfla5ZeqyZlfwrR2gcBSoBYrhAfyksw2AGFKRD3kY40RBQnV
y7jpopRemjgDzoGafM92N+oU1Yiq2NX4htoG7iym/ezQhxNm7l2qIeshRVxv8JWA
daJO/Bk8hcUTzeBR97/0XNg5G0TVX0atzpciZQAQB3cSekg7kKiveYTd1bK1OLlw
SAuTmI55VYp9Pq3Q1z9MCkJFeKBE1JuEFqtun7WKeeL1Fz/wM3f1XTlir+r0n4ZR
PQyKcGfqeWodrr90ow1XGnSHxwDaYuErKn8xicSjpEEBPCPg9kWnSUfvH91vJDAd
9lCFSwe9I1bianSAi+BUCwPA0zdD8S+HQLd571dVFzSiV8bCVc+fjQKyhC/wAh5Y
LNyJKZeafqRVjpsF2JDdmHV5tUbvCd+rP7Mqr/EXHsJOcnWmlssvvwGocS2LsrhB
Z3D39VbTwG1NflBcDKpVN0fwjWT+Zv11Mtcub/Gs67+HYQRXOBUOlhkINoAx7xcx
V3NWK4xkVVW3agBQxhWkGdNaQW8Ogxs7XDtTu+7ONvP7lK4/FEQtDfknAxKw0D69
LoikGeI4+oxXVxCd0PFRTS/rAqTf2JO8dnHmwpWLpablHs1Ijr+dxuhibJnBFLRk
cMM/3wCBn07qmYLS47nZCycyE/QlF23d6Q56qm2Yab8XJn8hO3plKSpq25aYXJya
ziDpQ1eX6f8SrBqbapTUVbUmDt9SLQxi56Dj0hxzz+Sj9mP6rZhjDmq7Hr7TAX6q
XgxU/+sZq82rI14Ca1jgG2Xmjz+/hsP3uoJEWlE9Ek7bS8vkR4uHrtOszwmw+Mpj
Z535z5uYGQVzMYX7yO4TWSdssj/jdmbCHGnF6cGBtRMCD4ZjS1eJ7QNKMOqZm1aY
1dvIsu2n95JCMpZBaasA83EsW2M7hhmwN6RPfbyN3bLAm4rkOweh54gkojpsy2Lq
ElAlVBErz2oCKjacq2HhbXhdd7AMRTOf8KciXZL0ukoTWA7uXF9cC0f+iNAItESH
GVNoagar/a6greBIOKhd5cODJE1pY/FYH++BnIHgv+XEVac/klPytJjfFG5YoI2O
uybKQYgM2VwYuzWMAoo2IIXjzF05sYGIAV2jvsKW+5VixGMx3uudAN5gnMOEvl2m
jpWRsukgySk0+tQkHn8XV17LpyrGF8R5oI6hWUGCC99V+42OZScLCzvgUdB6xH23
PrKkBFjeYwiFyEwBTu8nCEgwK5ily5LiNKLDYmcOJvkFS9geQoOyoMF+IzQC6/TO
lTJEWoP79gPPoyF1qleJ6b1yx1xOxug4fUWsWfXnyhUsJIOlUns7XceymdjH6i5o
w9/Z7kIOZ4+wM8GnjyOAUBnRmVudnOybJ91aLQz00bySyi2Ahbox/WxMFXEZxycv
NH/dhBozMHT3vjQslL31QgLSlsLgVdsVtVcm5ig2PVvUBPLcSBRiY7oEuHLFbH/w
55xBvBZNt3xGlVFmFCMZjzWR7hzH0WdtivP1bnUJdy3LfUMebB40VhYNZ/EQSLEx
Jrw8U5e+9s/CnuahKv2rH8SAkCc3s315sj+JW3eoIsJkdF+uOVuvuBM04UdnQ3Ua
h6U1qjqBmwo4/hbAvbIFZfw/3W+nn6VhlGzdrssvJOZUH2ltOpLN0stpKHDGFwFZ
NaMrAT8Gw4o+vPQOjwsNd/ooNTcSPW13OvZPf//NrxRlhn+DvqJrIJgzEtp/lhtc
Wo/ly0cCA/ow16NR26ukF62SWhxIp5nDev43cBJaTJ28wJR7PfG7LWsNGCMGbHmr
AeAlhulHl+6j75JUusFWla9pOjlrR6FBGwgx0M6X2lIZH3M5EOV3mXWfHBJj0hbz
gHmIlWvLIO/a9xnVWTy3aS9mHDR4zmGr0wqGqxJ4rPevU6P5uXASWQwrRaloCPN/
Lw4AcN7Lir4KsWWLCbyBiI0+Jm3pyYmPf0e4zrWYCRPO/ksEHmcdNPW8L2VJ4LSO
JDsYmKIxIrrlZpM4FtNmzSpX8nIUNM96SAa9mO/sZemIKGGCbnFMRriT5C2BGMGk
LpG2CHdSUMI00xLzRY68sf4u95XCH1mB1Mv94B0TsRRObXJlQj9wZEJJN9V7rbKA
KCZzBHF8Gc8OomhyKkZ3en8K50/4NwzJTf3TGMwBwYt31hjKc3BzF+loNhmSNWtx
ld/sagRvEjq5XlMiKymV9uShSvr0YPFrYsLR9Nmp8okaFoqr17L11q9r7L4s7haT
E+V2cQ0yE1b2f/kqOHD/pry4E76MQ2zekpm36fDd9n9eMqWMoKVKubjZ7vE7axOW
qwOYW68KEchxly51hQxk0es8tBk+gjl9kTQJ39/wb/wadD26J/D2GRH3EBU3FGNR
Y7Uah2wLojYMTPOlBjE2oPfnAJQRcKaQaBcb0fgBF1tCcMssqCf6joHV9fVTcXgZ
qCqueP3pADcmC7NybSRdrE5FZjWbhSQ1XnCLO9wYHOzZ5LmMyI7pks0fYfD8kefn
PWvBAgX+PzSyU314zDeVPnRHzLM1qRTxHUVnB1/1T3b8g5QJgnVF48hWs/cLvSKi
6byrlVXinaznTcXK5JvG5xWCa4tGdpzFZ3MXHFvfINrlrFpGjGuNDoAnKopmZQIY
UIY2E4RhBYl/lL8qqpDQqDi9Q8qNhO/vI4KaiQAMgbrilvsk9rACEgMlaKT5Q6Ku
GVZCYjACeISREbltfgcPS1Yo32J6CaiTJ9iSobFvHiZ0pqy3KASYndAjg1iioUTy
fEeXGMNgrobwdhmT7WonLcGkylsE3XpyKFCpWB1KC1Vt8i6AQbikMTi+amt2IC5k
2pekgp4+baKEAc8WS5YS5B6ks1MszU1unfFUR4WBcrm6Tazcm/2He0nlae+yFTWS
PCI3629sIxkX/8D1aA6VWn+oEKRp6FaR1lh0mEqaVtrnKkz84bJhZhVPRRmQLf5g
LTxY9HJbaLtF97nDzX0f5ElWxByes/xsBUwVl2XDuTTdxADEPRmg77jPExazVHRT
9Wus3iJbF6b+of1VRkWTaQSlZXKMw67Dn1+bCoYuRU8Ph89BgllSlG24xILRUWgx
4khq0O+eycBQmKOlIrHwWdoEMTiqBTNNBGFrvfMu9zMFF5FeZcE9xx9Zbvi5D9Dz
XbJrW3WHedVjFbenzVEIY1EFvgs502b9GYfJ0eOIOjLjNrRJwGWShZ8k4VBjg7oM
KCqh0h+0KcA+yCqXQxRlMLKNlfbJwMUndK2MRyMnX8tP0NNPzHjxt9MzITcuVcXA
YEXgc1HIp8Tw+nsEtb+kUFWa7+KliYRI0I0mWEte6B7jdRr8MSMK9zd4pu7GvX2J
MpGsydB/ao8k8Evx97ltgoDZ8gFygYr/wMnxLySNO+AY0Y4MPMyjovW5vVjAe+A2
qclDPi6Z8zZ3ud5KIpSAPRYHwM7PnMjxpjkRJbj96ncyLQQTAlAqg+fjwfCS+IsA
C/AG82Z4SykLb2QmVoGrVD6uhovvIo0f3tlQsZuyhHePtpBPrV+altNEEd8gCnO7
kO4VrW33GM5ypfFFxmhMofthvr/Nwmpk48w3RtQF8NvJGXcXf3BjnynE92JMn7GL
Xph0VJT/dTtUaEkAEHob9Sh1v7PiHBZGcEwNgvi9kCn1mDZ6yhujAhwFrzANJQjN
HsXUQC8QL4xBWbuVF0pSiOrTHIfaz/zAE4P7La1vHQw5m+ODDWZOo89Du89BX4ki
q5cx3QZHLntESvq4LyIsZ41wNAe8Sa9ZzmGwg7p/HVP5/bCL/7iInp+BICJVerU2
/PRMsVNn9kHXD28XteR2k1k6HrTQTRB3P9oS4G3xofKJolx0AwX7EfuHVTH7uzkQ
UM6anu33aM95WmIdbxXHOxp6W1oX1DRss2TU/RquLwt4+9D05fXOM0UOSkyxSllu
Ab36lsHAMM/ZonRfKfiAyKGFXoARFZ8KHrUxttT7ERzh7WLRRY4iO+CDwjRzYNXp
flakZ0PpOSuFR9axQYh7zsZ/oVV5uBJNSdcm0tC61N24t9/H4HKkPCJqSEMpAoDB
TM3aTlPyw06XTt4nTPJQ7HYSmAisENOYd2tJ6aImoUuN4Pn3zUg1ntRTlcBseqMN
c+5JKoKa5VfO03HCpIDn6TprEk3HtBNAPhjWKDzSq83275K9bgsaDECOUm4Qisk9
xgkksojzZ28AbCnOxDqSJbZMNfuBpsXcZwrilrWJdEVc61WihleQLcQ6CucKRp5a
98uCi29gIhh7jW8L5LP5V+7wclTNEMPX8syuGaUlJnSVKnC1qlUygkXxGIxDxY79
ZnRJv7jY7MqjetVE7m7OVUuhHGBga57+LZ/wEPsB5hyB6OXoNGo++wTnPIHaUycl
hWjyBJlAVjysVf1FFwBQXyWHjCgD1it+lb7BOfjnC4iXx3DBYY6EEl1/H1eVqUC0
vG/VksoZa8exAEbj985yVEm5NKDbqtPpplqegfOle//wIEIDxP6c48W9XlWfCAMi
OCYq0q7qahfmodb35o4zSOLXU0rszGTAz1EFq6QcuzHpZorr45fGUl+Nv9FoJRCw
EQm+RE/eHmwYLJfjZMAbNYVtWFz7fF+NIUs5r69nHKWQcAsmqWlnk2cVtj3PvjWx
p9GMWRW5RpCOCKXkjwYT28HwINTtahE0b8riyDoFICpJTtY/xbDnviRHLUWDyGRc
9rZDx3phQdwC3/2kLF5MLl5rna7oE7bN8C992JtmA3ImKh2oUNdrD/gyfSMZ85Vh
Ojxh2tegLFq/KnrPKlybbk2Sif0od9WUaWtYKSDw1G92YbH5s7NAPgasO6MmFz/3
ZFvpLhEpZ1/k+1ezLqOCajmelu7cQ2+oECyrXeBrCz/tJCdvSXC2xM2WpxUYp99z
aDrY7x46k1nKBSA1XbNNkdZecdD+I26zNed+CF1nptLwRHDxc+gc/E2FOsZOLJ+m
K+nD1bB+uwekSzqCTEyxYmI7uPdegxFKqqsy4M4g9ywmsxzL2zDbOquSrwTEVPi4
SX/S7BLjCxFnjvew7BgZd7GC4N+HCcg9jxHQD28QxxepkcVw8DC3A6Lix5EO6gaK
T//OZG9KAHJjPx+8c/slIUiKEwT7ZIya8hAKE253FZGm9lnsbY5g4wH4oXPa4nZP
C6xsz6pjieKJKjkBYK0ZLDJBplHXNjfLHb7TwUUOc6qfcn7WJ54nqTIUGftjousb
/dm0Hc+Os+qUIvu/UczxaC6U/j7Y+fa770UrSUIz/nfseVb8GTOejqDvA2cLfdqh
AiYLRyXm1ssI4FALx0H+8GBLiBbrOaYudEFena6E5Nw9qdXrLyMiX7E0NjTzDa8+
rIV/TYmTXw2gKV34b3eJSJs2SbaV2tq6D7cZO6hPLFSg7DlV1S4dDCzwR11jMDlg
9wWi0j+QTDvrJAdSygfyVgtMPNaNax/Vc8W6JsTAYhz7MCUin4uuPUzEFdg2suaO
D//tJoS9sKWm4dTg+e3c7cYBRpm7IJBTPx6xb5opVSqO9DmuMrA7CaJGqGj0B/OZ
NUdWmc62cKKMvn5fiYCDJVWEfoUfZ/RvK4/AvVZMdUvmtSo+CUKdHNGY9GiZJ2Ts
oYSAw7nKO35ekWGqAhjJrwQT88x9TfIobxjq9WEp0HHuAUeCAHXJvxO/TBHTJOVw
2vPMuMuFkDA5aHBLyjvuxe9fWnG4i4CiJRjxm8xhPxFQ3xTgLrFCRCcEUCATkDwW
IYpyb/jle/Ofc7oFMsLbB09S/M2z7Nn4rFfvjRtFhD/aMo7mtiKYjyNUEvC84T33
b3VrI3FHX+aNfEGSICyEfAuzYSfiJYhdThnt48gvlLrOJnOIA7isaXgc3haa1kU+
wbvFsoObW7Uy159q3e0fK7YB6p763knC4W8yNLFZlSKF1R4PYWVkKdshEiY5Iyyv
j9VYUj8nCjOYI7s/GK6ENJaGsno3V5g6S+kpqPQcs4YcvyxLKm4lO2HCr5kfPAuo
VCwr97w9asi2Sq2XiDyB6mbmjb76EN7ELLP3w4c0eaoRxFgd4fPk4cXF31V0kThJ
bIeaPd1E0jYpm61F8w9fWisfzXuifj0rbZP3f592tCVu9YVodijaivGOZceOXzM7
xUAYCXH7HeRQyqMu8d5vinWNbq97r1BJGUu35mEb9TgngfUfxLRjUFS1K1pNq/uK
mhwEKiakMf+xbvlOM0jk0WGjhwyVpDWoIwy9q5z97LJiUy8k56huiDNase8kO+B2
npmcIa96Fh3uwp3SrBJp+StNX3rXJl5J18JtU5ZNzi0AnB7F+iE2f/BTZoyNCi3M
KUkdfvEZbfzm+Fkyt7lyb77HrDEpVuZQxOZMAKFFSpBqnyYNxc71ops012g8kDQJ
w2iBFTvEWWnsk/bw5ut9HvOmLBcnt+XUwOXXj0Vk4etqoZkC6k7mxQiZw9x3SEaQ
BR5mC2C0btkN24yU7mK1NPDO3HkPpVLm/48rgeooAKIzZjzOKNLgBrZJVNIT/n1h
J8Qg6HnRdHOzle6u54J0/It59u180mfOCwCHXiS74mhRXCYjuAkzvF16jseOOu0F
kau/kOd+WYcSucJBJF91VoJjSZ185fOzaix1bZ5zv+IBDeW7eAb0aoApWgqi6NkX
DSvqm5wZReGh5GrWaMK18oxU7QMZtnY5Z57MeTjfzDYnFlrXBcsvJ1B835r+p6Kx
bopEI9XOfyQKcbqLpd18GxvxsXGeOT2UMubPGZNTbezh3X2e7IRQymaMbpyTENLK
+oSsEtV1XBt99e+DGJTqe13TOb01LQR3Ki6I8NgNx2uXHDMOw3X3nh27fxOJJfo0
kt3bVpo1vsWLZ2BMCmQmLgikr+eoUz1e2IxsQ4u6FewHhXV+FjXWSKsDyeaL035n
03HrIzakb5WyI2SIWiObOmgAnIoj655WGfuQmXGdRpJcTIw0bAtPiBkItiQ3atYe
v47Q6sFW0Wph2qyIFeX/MSZpEt1Zf6A5pGU3URxtANKS1lKWgfi6JMfeispLgkze
gOUTTEGzsWnx/z57iRLOwv0Ndgy3+QmrPw3TWrtwnlqKLtUL9nA81r52vj4CJkuJ
7kd9x0pv8a5ohUxLuy/4XOXZNwXXSA76QujGwDbB97U2S5v7ZGwVgYrMwxstOL7r
CZTsnRVNMcAJlfyHFxao0T2UrlGfURlgC2Kgj3LJLTwXH8j3A4usYudBZFEPuPW2
fk6hwQeA12tkx2RRed7GccpOyuOKDXIi1NHKQLhQvD3AfTyXFWuDie9opk3diOXz
4IIwW1AJBNIZaZLi4lqOvZUrNoAaQtY2K921cUYHJHhnRSpUeNM2C8GP5ufscvRe
zb0OcKJ7EH2OpGTc5AsgMSfJjkCpreomTwdynUlg+OJBhqPVtDSP7A6Qma4YwJWN
l3kDLGlkGQlfGRUJ1DgLJtDE0bNmdD/nXhdkkONOg8GtojGdKLXiFR0euG6KedvU
r/a+rq5hIrETlDRuPUhwj7FSh3b3WA2hsHxGPdIaSLrGOY5GltJvHtxE67Gx2TDr
+BGgyxg/UzSwZuRVCFRfVgJUEcULOR6dCJp8Dxji9viYsAIvb3+2CNfSEsMnfLzD
Amv3eV3wBTiuYXXzpNoEnvBjqXZN/BGKFrK85M4cNZTOu45KmdK8tiUBRZC175JJ
Qkx6mdxVTqgYwLByNLhWXTIskcLO/zEgBffFqTu3THq9ENVGwIsECMLwqDqtVZ2R
NNyOtVYYntl1erwgEGI/IxtBAzQxa8Ew+wQPn2PEZLGyxPISconYBS0Wrghmo93n
4aVyo/yd3NOAxwONM62oBl3OC4TtK3OpxgUqY8jI//rThM3VZaztc/SQPG7DXocG
LJv/op9A8TRXklqaMi7ZOHhmz6qz9NjhP0/mOjvUcNPSGaSGKySAJMNech5sbrjz
yjnNdvBsBBivTO1xy3HxJvEBPwLdgFXMpatArA9838Hs8gh8mqPhjM3GBECrJCGu
XjQqqglQFrTA2MIdadFXmstOYp26xdB6hlixMhzOvwvG9BizsFMQkSAToH2hE8/D
lIJSDWfAlCJ54VT1z9KBUvxKcyf8ISAYOt5uGOKQpvMNdI16lM+xZ2WaTJdlOMdh
gLlOJ/v1ZS0J7aYHs9K4zCiQ4n6bWZlmZSVVzBAHFU8FQlr193bafd+Ot6mLdpeQ
6Y/ObJZ59+t4O8xxw0yGms5vGimGQdleAAEQstvPVtSX7ObKYkfJvBvXBWYbZPq5
rXivUIjKXyxmwpzCvOGWyD7uhrumOKhoovKABpP76HGAjN5leoED0prOBxddAgNo
zMP8TJNvqIM47P/C2K3IZUVfX8Agbb+OYblkxbEW7i/LuLHuYY7YJpA+ZxjyNajQ
0QRF42id1DHRU9FG41HNnebj8i/zq5xdesy8kDC/PZTCTXqg9cV1bSiBy9R88QC6
sWSGckQze7zcrT/1mL/7wG6kotf0pm5H73qPZ+c1zK6GZ9ThOmgHMIEIeXwNLJCQ
pQoskP8ODsCMX9X8QvqhwnIRONUWatW7bfHPo/KmPl6M9gSZ6v73R7OmPFzn/5EF
a2QWWaEdakQyQMi8+eN0esteRC6jVi1pVeIdX3/gSXwHgZeF2v3By5SLUXaBoXaz
31N0YNgdgH1l0+mT0eSuABnne0rYRFnhlF4ldemhR9RGfoSGqORhbR9WPptbin+4
91Jfwnm+cB5nn/UoaQNQs4ra5BPEpQOQcG6a2BZL5agIwpjIBoIy/QnekSiA9nBN
5TntEUiu36EzG6S/gRlbVj3dDgmsqx6Sueaqr9pcp+Qo5CuzTIWCUQBXS6Q94Yqt
AzwD66NlNKLH6XffLzfWr9YLKMoF6ZwsId7R/eXX8CULl4j+C+9VG6sz1rgzYb2H
5cKgXGheBZoqd5KxkL0kJR9D+t6aup9DGgScYudeW1PybWa8PlyHFJQmNk/ii8eN
N4rDlO4BaGpt8x9OuVd2ldML5Q/9ynxl9M/aYgfKnryc6G9AGhODeXXvi3kg9MlJ
Nv/UqslJpOpTI2VF/H5pKJtoA4ZQwq4/3N1/9ONFFwywIMoU45R21DRf8QNh/PTT
wBFQ3lzEueCpXAxMYaKdl6znrPe/GTaY+fdF1oOgkR3AHHx8E4rgTqQ0uuB6yFsi
mM1dkO2EGepIhluUJA8V2xEDMmKHKwaVaxfofOVolD7/TxP/+D3apmy3AJkdu35F
AjhA6p6ozpYXGFIBJIDG6PChgLUbyUXC/mgcsHW8n9uo3yLAK4Rs8haNs2KZnlMf
AXO2TuvLRd/fZmdHOZBZICqdZCVU0b8H/uAXZ9UEumOv1CItx4cRl18mIzQg7Ev4
P/0ooA8tabs4lDoHVQ+YJQDLn8l5OWCMyAW7qkDHERO51Ixg5qf5+myGA3r5ZEJ2
k4P9BKxrj2pyPQ6++c7d0DmBmyVrRavnAk1XUSp8uwApAM8yLaWNatWapYfCYNQi
BIJ1WuTSglzFsFBqrsGubv/DwiHaakyrH4Yhdb1gmwLg69/ovu+1ENQ+iN3v9dRg
H3TcXqvDgG27Z9+S6VQ2rZuLDp4TZbrHyny2n0Y11fbzdaDNMTyUtL/yeGjRLYRx
TMangoQmtbNrBqfzsHApOWRMzZf5NEcH2MZ6LH19nO19R1FRqwca0yMAwFl6mJXW
IDfJ/PXO9rWNgV/U4zRPx7IHMscQCd79+AiTqtBqY7SBRvI1V9BqeB8paP+huJcq
IVTbZWk8Vr/6/pfrmDw8yrwMPCf1J4yUpS680KNw4W2AIuLK933R+D5zV5O6jPvK
zebi400pA8qgbcmgLS8MdYpykJAvDlB5Y68jMEvEr9SNFnMrcFMXVnZth7xTrbTx
uoPJHuQJfnOHAO2cW/5Iy2l4dKu8DKXsSPASmLcik2svGWTmH3RWgD5JixlzzzNR
+j7TU3On2TcLTftIOO1E5pwqospVQcpgh3sOqt1UAhjiuKm8TRD7LKsfWoB5UxqL
hU99UUSCE8Yxe6wE271TEiGqNbL4gfxTW6SvMcLfSEtgXYOAxkh9eqyzUoZWuZn+
lk/vZQEGv5HaPMMHiXV9rOgnZcoA5eAzToLMhswsKOBA2USDNtaTUHNPXorxzTeb
YQtgAAceFS4MSJ/cucqqGLVorG0sdiTlTTegJGqoQW86+F627Rm+D2F2G6c/Qh6O
EoUHGefc+0va0wfQz3mEEjYaXoTFxCLpXFLZjWMHAOic+zayH44UlP9o6kb74TBr
QPohOxRl5fWXrkSwnq19FF/B1YNoqSHCSbmAeOXipkCkxiRWOclRsM67WUpLzDyE
J49ZECATqzc0CC4ttnoSCccRTyLPDyqgGiw1LhU2KjORz9jt6MLSA6X4ILAOTdTX
zG8YSH1Wy9RleJnbTrvUYknjgRTjZi+MyvQWyuUGUTU6R2qa+YVXIJqpgzP//qao
xYpy3va1AM9TEHarwn5iPc6vcryxZMlMaZiqIrERPr3Fhfw+BF7OVW247UjjZIBf
oYfMMZ9AwNQcDRkKuXIXnyDqZtdlzJm0/qNAWTjX+VH4HHOl4GFK0C2P09IBLIWp
CjWdzvzZWc0GDYS3X5DafzCGMLFLYN98mI+QMMdbPZitvzr3/hXE3J9jXR5zshme
jq5tgwQDl4H+7odmJCD5sWUCFKWvcf9a0jLn+NHo5in+ZeBnH8CoTkXM/5X5fzoe
4DDdgp19a2mFuCeFTNJ+o6Sdd5U8lcI7lgv42kfKvivEpFxiCjNclCyCyNTxyOqt
5hRKNpPN8Z4bBEFnw05eaZqopA+5jdRGoyIOuXpMOkrHbfa0x8Xt4NLV7VMR/DnH
B+OhVqFMz66WO5jHxg7lN3mVE/ruVaT71auXz17Vkz42ZY0GX0Uw6+TsJqRUE2Yy
imbmMsdGiVe1bmbYFkqoSvsUoJmh82ouFdayDXJUDBmW2/2Db0J1k7WdnZiD6DYA
gZ5U3vASm7hx5rSV/vEEoQO40NYT78HuuWXyZIJljIXBTx3bmZQ1/DCpotQmufpJ
Zp1mU0/1FnTUPpcsEmwPrWTb6eHxPrPzjpNel/ehAMytvHrJtTvkyQeq6wegTcNR
LQq8fEQhZmPHe5Jqf/WY5hlgkqaLzwgMM8mi07SeakEL1sJzGSOnyY14B09U3d7c
iw+MiRYoLvMegMsfifMmzbW/sXCeAJvqt0y+0roezUxEPNswLY8Fj4a55afCo9W2
D09+Xu98zkJucDgO8XNtfaUj+0gb3aFt9ac5AXVGFvRtC/nbtheqNRSb2kYTDb2F
nWgNCkICj4QwwKl8Z+cvdBrzk8zQRq0zxkMiuomCk7a3y012YhAIcAsP7Z2ZM13n
uF+hDjv0diaLMAy5dC/uoeASOlHeVdso1y/Td5DQjbf9KSQhFIhbpu9q4qxe0EGY
9F4xp5h2L7QeW+Yb2AAz2Z3IICk301ZtH1dh3Iwar+jBC0zuV6AnDK0i6xs3xNlV
cLwsDuzIf6b+Qnc9DnI/8E0BgC8CCh29mzao4yonhJgd/K7rFwOPx7yrQMo7WTM5
/8pBNbjKLjWZltG0XsGAMKl4ExYlWDfb93cFWRN2jDER3Qurv7G6K5lSw50LTkI2
YmpEW81oBZ8XB1x2BfvNKwKbLXPuTG4j6eBsXk7s98fSM8cwqtT5EU8RgNcud6+p
GxVHD/PHGFbcsHpnf0PSA1bgRG9ANBg4Jj2BPuZ8pQaPK5HAxgz89fm3doR2sZnI
Fes8Wh74kp9D2dM+V7nox+n0dnvsP8WgrLuGhmy2wZXcdcnVyucieAe9tB76CYWU
fT+XUK1/cYMfpX7Q8raVMXwtgdPp0npa6bBZKNjKmMy5txThvTYKsnr0qXVvIE30
xHTWCL7cVctkT8CWuGtUSrxl/b5Itu0rVTe0J2YWfwNgXIyKeU3xwJenFND3gA3I
n3Xyk7XMjT/Vxz7DJ0hxVAcC38X7/cB7OEb2t5m9+M8wK5f7fZpjt1JkepDA6kBB
pEWorfJB1w4Tq1BJ/mA6amvV5YtrBG2Pq8lOBbnrA/wnAHv3qusih7CfqCX0W5+M
oFXKuLcF0AZWI1d1Kg1sXlJY47INY0KRk4KVNyBYIPgQeYzXxodl7/wfC6Q5JWx5
VMhJU/wRgKzdDmjsWFQ57NwMGueeDslpOD+/gOvGZIq4vMqFDXGJCNQBrWE8OZEg
MnG3JXWbG9/H3+brJlhRZ0GgHTGQYYN0OZI08fbq+FEzFcFv7XxXfYKa1B0CZ+4U
ccprNBLDF2pPa2/CYVMVtr4eqerVJPW6OfJbM+4+wL5pSMhIQHExZw0xDXJq7Gaj
lemkQ+zVXprTjbvOoEEOOMtNz+gJ734ngVzj3JlxViVsStve1u6u3N/ZxeU0agq6
sEXSOtk7rTTtLKQ1b42FxWVv7eKbM50Ikd1sc30KKVcdZLFdqgUem7KgOSCPJm1c
rkRqr0KnoGsdB+cbtA9lD+XEaeypwbd03bnKE8JE3AoLisQ3/IgroqETl1hQ53vh
jNrLT9+9M6pd4qUnLGXPoWwexxazK7tKE+lPMen8t/PDfB6d4jK+EYOIhRmaK9o8
Jt5zntmbtsc1Xt5SK7PBhlvvE4FuJOQM8W5SBhDqf6NfsuZz0Rv4/FwqCDTzpc2q
8IneUeADnL2wXiTVSpnayKVYeXwWxkx8BSHf+rVbS2TAOvMC+SiLi8hdErgJg1fb
A4qY8u2Ynn4M8aqSSi8QYXatYcRYDqQ4z7+8g0r50HK8qZJEvZqexYO0ayiS4xw0
PMEoqgKp/9RzgDMut8EYxM3RYpZb/5tJl2u4YkRdAuvqLecnzK1+itsIUHdpEPVh
pZ6FHTZaKv2teBgTpeQPodYT/bJfbeO2rmLmS1kq7lmmyruiv1Eu/2NOi4hmim4l
Z+ygc9fIHo610NmbIE5of6/2xNDGQmwpm7QoM0lKaTff8RFsi3QpB8xumZFLhaVL
bAB05LJqXik+dkacmvv3EVYQ203KtmM+IMtLiYKlyQbxzVGqmHjNygEmSZVMUQY3
76UrDiFMgWJc3ccZRdCSusAakPdoizk/okk1hWUj3N7IIiGnjJQPwoZmZ8+HG4Ij
t3wSG3+omaDaPNMfr4LE5hSECPrHxJ8HscZMfova02A/61PP6EYA0VKhPk+y5TEN
Lhe+IeFr+WzFRrh/1V8BtY0KlGZ40Hdum43dTN8TuoCur7aPlafGrq7RZiQNFobG
E9XnZbZ6e2YWU7IK9HAM7kes2sDdqd7pc+ANf7vz/a2rgAMp14W3yzoj594+5ijd
f0OanVjX8uk3DVZoE8P78kd2kPHEYg4Qw5G80s4BnARxiXYd87347F2pi19fZva9
BkJWgH0J8e4r808u0wesQQmwavRmgH5JX/yvpscBK8tZHecwUcs6do80nOO8yxUH
15AepV2/ZWHGIF/W9iOjgZ6f/9+jYHo9G0+/vMxwZWllvzadBepnnF5peiyZ2nj1
dWSCrytR0QRSGp1M7KBG8iLWmCAx8+ch17MaNreZbN2E7uQK/Ya2RFi5OAVVhdTh
2nXyefwUk1YywncEpzc5CJD1eCDh/bNP/z4Fpsp7F0NEusG7fCpyB/rb1qN6a7wU
ENiid/2aSMpYhqxKPy4hdaZfAYSdRb3zzPTUVaJTuHSKUY8InsgyvKCsr0P7YwHK
tVVJHk6NB4gRMvIY1kPN099WpqTzzcH+Wbphdkr5k/oMZ0hNhstMGJ/Hq9iSG1ka
5C6/stEGAUR8nH02E1D3lOaF+Y4L2+JOF39K6Ks1m0vzagdCJSV9wzwqq3W+1tKn
CNuqGIoCi51s1N9SBZ3DNjTPEwJQvvhzaIHzx03sqf3TZdoI71Jd4SQmcEMOotOS
AWNNQ7lrTmpWqOXaVQraTDE4faTpRBW2mNYh7tq9Xs6QBi8af04kTDGD5SbidV5u
nm/2B+0kszN9AXmP+MDD1wnV/3jXUC9OAd6uLD/4mCJ7M7Eqq94fWsbJGN6AivLQ
JlDcY5jjAESxio/Nhr5QnOIwtmBEOtiz1uXy8u8PrPW4RdqDBbp1/uRubFWfYfY1
WyUNAy3klY2vCvi6MwAoeCEi9Z/q544BlEEW9XFJX+XCkRz3ljlKCwWGFXXXHjEs
y/hOX8eibRbgdoiqgNvl5eVdqNTnXBFYWZ/Qo3DL0eD4DgPp/W8jhlUtnclhVjYK
1ExymPq1rgMglNIof0He4YoHT+SwSgK2kSwoUtxbwueAs+zDzYQOihaPCFwkiUWF
LGY2izjpisHlq3dsVo4AEQoLs0CBCnCaD/MqJqOVJH5oTNOjv8e0vKeA+AMeRnsZ
S7+FGCitUeWSps5vyv4bSy6RKRx0dW0tsuKEchcplUDnY4NfouECyv/c5o1M6p+U
HQWwF32eEYp1J70nuWhRucbCLXMiLSfdgVXxv50eLo6DSj6eN904h8FQj73Gn+wM
Mp6c3BGqtNmRQZ23Pjr7o5uRp5C9mch8B/Ep3Aqxpz1hbuiJhOu+Kohh6mW8gpYL
pHT/ger9dKUrjHRv3tQfhe08LYg5Pk8Ex2ASqPauJkCQaQooWr+9w95P2rmo+Q9U
xAjX7s4t/nNpoB6W+vqRfUELjgnCMwi39kGceGgUiEoChZvuxBjNTgliD+5NdH5T
D2cOWwlnPVngf6nV4Zzdis9e+da81me8o9O3QoQ3XPFwzr/+dpbmpJ1j9bdS/vha
8QHNg2uAOJGNgsuZYIVCmjpiwZxD1o2iE9tmBlolO/Xzn8UvcX3ahyEGF60wpIj4
FZDnz+hLLa3ZlZHzOLHPcdstEBMNltLvd2iFoMOO38NLxxmmFiSuSGQ3M+cx1TIC
HxfCgcjOplrUiIc4gfzpmiC9+QQAxZwJbzUf5e1a64ov4B9sppfzzndS1Lf3q4rS
0hGKwn9Y8szSnwAGm1tzKBsifyz/wgZJ4cSooKSepZeamAwc7moORpJO9jzNvJdc
ma5Resw0HpQNUvbE7CSBcn69lCTR4+YwDJdMmSeBWMtbtnErxXAiO6iIv4Ee+Agz
49DRFv4MBJf5kEZ95UiH6TXVj7Zj1dt4qdWBPV1uCLeIlOi1C1Uak2baD0MrWoJy
mp6641fZQArRqXyizOygZObP2apcLnGWm9fAuolEbRgEk/QMEYKo4Lj+PYwEpVA8
ayy0SssZxgkliKLGP4rqF2cHcJibGxXvkl7IM7koeGQJ0Fow65VGF983YqhyoBfy
ICp9srxjJSwPVWvoAvE7EdbPO89GW/41UTxhsQnruhufOgz5UsNSy4NJTnw9EjPn
fnwxu8K0JbrnLEf412/g3pJL70N3Y0qYIqOx0YXuGFkOZmB7tfxd30XuGRX+gV8e
BU4fVO+udeRD3PptmH6Hm98sFBelEKjwjzGTt2FIgdrv1DrBWOR+VmZTvA8zdz0b
SaLQQig9ltDp8PHnhNmumi8R5cJplyfs0Z269zUarfvPFFiiTww3NWHdcpaczDOL
9bqylZ2wSweoG+jmB9paz6KeoRObrTYO92JTW8BhqLUzmZMgqv6HrEHjyrkS7H/F
amy60ha/98qZBEMVWcVQkhiDVVKKi78MQzeKLHMOTqSIDqN5GsJR0IBgdAhS51Ne
hdyzQa2NOkZbfEev+tBM6VTMygwwlSfhn9G/zWLbJx7HMJDc/waMHYUuoBS3WcNZ
o4PoKNvao8Edqwoz10GEz9Jiyx7vTal0jY//El2FS7cBoUThIQQmzzH67FIqRUQt
DlBqmlTezck8nZN9prUAXthtN7LVfeSpzz8TgzAPXOM/dZCtrVCvtbzmkeHk+L4m
FJ7QWd2gQWRi/fCh3XB+xg7l9FyyJJ+tvtXfzpDqYPgxATVsIBBra982p9fEmzog
6bTbkXHD/bd9A5fuN3G/vKPkUIf/JKpR3U1A/2Gn1mkp6Rl90azzy6Y20mnLfwiE
Beti0uMOiCKhDFffNxokhXAGnBFKgfCXQN1G+TYoDlZrHoD4fsylfbfUczwkdVt8
piZT77TwwD/3aBtf40aEf59k5pJh8iPTomiEwfuSDXgoZ9kER+zZRPl3p5+qmMjO
2XiiCH5gFxrpRHz0OcRaVgbmB2MtTHkwJx+JtIzFlc4adf80oQBrPV33GxMpx+uT
QM2uTg6nD+z0yFuQkdDeNwdUA3Z4zKs0CnDlh5om3G5K0e13EX2NEhDhCcge18jn
ULj4cD7KeIO0slWhnY4eBlWp5ZyXpGtlz2mOC/xR/3sSgVyXePeqB8+nj34tMQD+
l7MSMk359SMGDOF+8zAFABjKWotEOKBUMgQoAZGFXmfISuLA0U+ew5odIShAlRj0
YmDtK1SF4V9X4VhsjxC5MsMHHX2C3IpIGD4MVnC3QvvfzwFY2EKQE3j6cJtS1SFS
VJfBHwEQPAm6cgVKyTYFzFSD1Aa/30i5hyw8dFd6FXVmINXEG6G4tRz3/f+0Mhr0
1umvswH6ct5ANmD+w6vShxnQdzS5OdkNVJxKTqXHW+uBEkk90ayySzC+cC45DOk+
1nNjAIGyWrhiDpevP5gMu6Y3Za8MR+kBPndMbrI6RZoYM3hKS1SDrybPEV0kA7hA
eY5QAMQjEbYWupFqBK+nrwQKiEJACda5ZPy8rdDLmu2/2Q6cYdPhWN34VGABHnzl
+ow8PYndmzcwKMAw8ZFCgkcA1Vmr4u4uakUxll0/6o9T0P65/xs56qeVWU7e+BUJ
YvuTBQwjWhRaANpqBXz9c1bNldgbJ+XawXAYgeQUIxp9Xu4rm5GfRfqq+OKtmiKs
3fhtfWOKrHg89pi+D0egCV3s+FIepyhECx8gDbBKwbOAfVc0Sbrqhc6+ZFi37CQ5
I4n0IH9dNFpUxyzDzJKcflWKMf3xYQRgbuIcRSsmqA++EyPe/n6/bEFEesUwEYQE
ccg7b7CvXyH7V1aFXmCto26bUl42eEG9hI5+nSnLeHEdOJ9Dx5w5Ox3HnkRpXRnS
oViyLB9Y5H4V+5wkqtn3UHCveWyEW+xsvAGa1GyHfn4X1eVJYrBhObUfPMgvMQtF
ODZrIwU4LS4NdMmN7u5IsFgJOHl5OKqRB3r5I6T9XtJs2DOT4MfDZpCCXZH8sa6X
egPgF6GfTl4Mdioy8L8dQbFjMOd1ErMtvZ+cdkPayRMc1wVDh97rXFzU8ifxfhJ1
bOV4/3xBm5pqkIY7a5peq2mO8UxtLGy1fUZclVe4aTzJv13/ZP+PsTwE6nYYDtKb
b8rRuQ6R02Dn4pr9Im96NXsAKvWr56q2yv9SIGa0/7+o5nlZH5X/8PKm+uw806Gw
2t09li4NCiGvF/13eXylhc/BwtWFMKatk9rOyFWA6Ub0x98py4NoGmCtz+DzORbO
AVZmaolkrPEKf5qXe0zAPCfcRBo4t6z0RPX+usocLRfIrfVNuOZYCMWZJdzFk7mD
fH/Y6qMQHUB7sFAd++m3nTxMHv+0OnQlsailnfR5sM7VGwQMqMxOFGVF0ak66mZY
cZ5HEDL8kUOqaqqHruXUm+HqhhffE2Kimk8vCvJTurhq/2XT/pfejny2b0glg0J/
AMU0kDGEDgAfBr+QRuD5dVZ10+GLSscxC8lzqvfGixj8QdsMge7fbktnAgWEE93T
KO47ndvXSt+iro+zVZ75pWtIdLp0wBlu1gdF2b21kR+P8HvtABvUWcjYuPjbSqem
ZHBQJ0gJ3AZghCwjwXajSynbWdIuqesaplhhezTEqJRD6UCDsbwuaIQa/xyf34a+
BfYl7FdPyUNtcV3RUc8+hke19H1EIqVl2VWQtr/IWba085IWH1f9U3Je/KN/VbtH
IA9vrN/CmOjBhyoonMlrjtqWfTUck4fd5eKelCphMlTFfsg800cSY3AhRDgprS+M
g/Xie4QUdsHmxnHC4KgcsekwRvN6jYtZEUX4FYPnnUO6X+IhixRE9wNzs7oLVW85
cmK28EIB/3xdgXy58S/5ZyykamMTh9TIkl337Q5GpHLk15IGA6BO112zgytNOXg4
mlNyFw4+Yb6rRg9ukz5IeukARDRwllk03DTEyhQahfkcXtqxL55li0ytVtL+WdAZ
A0ppGaEDPpz6S2kisEYzS/QQP0wezCfbvIKZBJVJ58m2pJAmOkgUg4mvQmqjbgU+
7rhEVhLf0mThT6oxR7UnshvcaguOBdO56jtLkVMoAItfO0r7TgefyVsZCuhvImVg
DJWt6PwvhYB0Ke1IweY7S4IGS/2Qb1A1tddJHOoSN44HH0Zo7WBg3zb6CN/KFJxt
B/UmhPUjnkbTlrsGm7X3AUXQG3d6SgJ/s/2AS/Fm+PtbotH0Oo0Fl1nRCmMPxbmE
cbbpsuYQFtYs2PJM7Q74Ut4VzG57uxITLnH3giCaHebcGrfyEo+meZVDvXJqPXN7
QY0C/j/15q2nT56w6VJELEFgeXTWTU4HhhH5sV+tl5iB6sVp+1Lb5CUHpMNj5xBa
OtdWCiV4PZn9GI5TUMfEajeEiCVu6g7gPmjZpbysi6k8Pgx8m6CTfWTngsHrC8om
fZ42m/lwRG1udgLwgi3xenpmKBH1r9WSn/upaC825KkbU2Dc2dnH5zhiMqiPgm0G
ChLRKii0tVVbW12CASggERUysscANUOPYP663+zur3irR8QWfiYKryJ46iZOI+Qj
CpRGm6DJvXVOm/fHABZSJZkuX3vjL138fwnLQEIvzlAePZ+z4lUQqG+diT4Ipyxy
l9fmXvQN3/vX4Boa4Esya86v3J7OPKNZ8wjKI3adoTbeN7/ErhaS1+cjOY8cH0XC
Og/JhiB5zic93fGiGCHWzh+Mj2KIwNxQT4UZsCP6JG/t0NS82kv4XyrZSUidAn9B
BRhCZq6EZSVKgSQSovDG3Bio/pYLz/GR4uEZnnPOrwXL4GafoCa4x8jQUHHr4IpX
d4jqrL3GqxECCSw9TlKT4LjGrTzR51WFlt33aAwZCvr/9LNXtI4IBc1sVS1S30XF
0dKNSh2wBhKmkVzRifeP6QYlXcnHr2aw57a+uE4nJccYohGhamAi54p2AFvRIhM5
sVAZAFVYuoGbUKzljf7CpLaKmhCeDKVWW9bVenpMweDpjwBlTLMQIN/Dv0dWoBCL
gPmGyJep0HP2cro3wv0NfzJRfTdWxYxnJLL7ENWO8bmwzUMNYALyAkoSTpmBIHB2
yHdUe5BqRC9GTmHsRzpW2++8eBLuzW/FoRq1T4N/DgqXJFiuxaRUiqkGFrSoKKeu
gLnIKtRnO+3qj6nVVP8bmCtNKQ+8eh9luVhY3IOgFjJeznyYtDJAp5EDzdWaxKQm
s/Yh6rjt2ZK5T0jFZXUWqygv3VrFY+/d9c/ygSYmFO3aLZIQwYXoxQhYnEJgRyuN
8ZWfcYavyMoyaubyWkNz+FwBB4cTv+W2dQ6uOyLNREuY9lC0SR5alc5NWlMHbog9
w3FwDh7GeVLyLc5ZSQ5DX/0FbJqLF6VOUSw8G130EubjOVIAaKyQz5I6t4vbS2Bj
OeTrABQ5c3U0LhpxROlMOm02dwhE3lcKp8AgaNmFgve2/ozlY/vVD/2oKV0xZdP1
FzppdWcMTEvHpmVce97X22kRHmXsq5UqsTztfR72M2lpu1tCgofyoyISivry8Xby
wlnd1jbt7dltYVjA+E98qOI69nknEdMScF+rG8QVNR6i/Nmh5tySnc2QhkHsuc2n
U1EO1z2BMG8GZor1KEh/1hN37uh1eFAWQCb4SU5/uDeSzAr2IvQifaYipk6cMNLp
k+/KotU+hVYlAPQGAK2ph56bHDhilCIUrN8Zfp9bCJtJq/oOWzETMKkfM+HdvzaF
suhwNNjEQ9EqcpP2HLAOfDbTCOC7iID5SmvuIl6c7leS7OLB9LuzfFUDzZXHdlk/
62f9NXS+9vulpu7TSdY14nuwSHMnxSUTs7M2S/77FV7nlUK+PaeOLKpmniQNVVFd
uyoExrulIKEksw+uBMWlPfqZ1aajkMku6++8JdDDgAkE3GEbOCxywHdvHJ5deGXV
jc2BxBGwHJh1FywcBHRNO9YHFemoQIXySTqEC9jhRAE3HDffST/DHy6SUjt1P2aD
4P4gMTCH7a2wu7BnQ5uNrYZ1f/iJyDLyB8oca54j6dGNR7BBhgwvx4XueQ6PXBZr
3Qk7GPvqgPObn0p9XjAIfRNc9ZcD9P3TTT8TB2kQLL5oCOYMSyArcfU4hqxRPdTn
WVRGPdFgin65KGJ8aJiyhxcOTgcs27v1nJyxFvc0+SIuQZ9nYkfemlONmbm7ans8
LFL1dln5iUBX6xeJE+dO1L/fttWx2Ti8eABbj/tnM7QVA20sh+2O1/y5tfbs/fm0
fj8e7LNbkWhpvJWlx7VhO6gYyMz054KOQ1Pt2dHZmZnTZsDoIBIOtOn+V+RLVAYU
qnxC5su/wLMMlHiiBq3uzpa8WMqPyBp21Pd24/O56flGICHn19csi9NBJ1VVns+J
aYrckcwCXFSLSxYgtR66LDe7GXvIe++nFJiuYi5SQr1Qw00ev9mUE21TbZnRBz7i
scQclV3Vuj5wdF9fJEaM1lqtpP0yQmIPEkiz+cb+3jlbqhpyv6gQq5VldDr7n3A8
W2fbvuDAcZklXrBz2X5D9AGxOm0Q7OEaNWprWqI+skPwqjJFogpK6qCmQIhNKaPb
DefaffDv14tZddrd+uILxM3vYKsskUnaokBikw6hPlhQJELk6vXr5rO2hf07zWjm
d3ij1FzVPtB4PzrQD5/K7yXifxjFY2I0EMa8XdITO9HTY4gUyuazzqdgw5X2bv1h
lkwQZuyg1HFCyjx0Hil6i24pU+4D9H1flxAb/xU/QK6ha3TaW/XnErGoq6TqF6b9
BKJmUKgpwQRNQLVmkULIYAKnlPnrAwEdSygFRxX7VLW7xhhZXazySdJeGTRoFcYb
zOMFNXWHWN4SJmE33xr0mvXShuQVIAXzpCDDHmRZEwRD8idEEWtqnhX0vpRRAxfd
BKCJm7gZEr4XPr/RFrfL8iegBhNz+I+1YFF8RoCiQg/yYHDVDM9xrxjxdKLywPLj
q7YrDe6MpltGvbGh5D1RUHdQ7XfiwATzqE9dBo16kBWsIZq9TvQDnfe/RbPiUPp+
03ZwTzp9xmbA7Zzh5VMLyM8yKh/ssH4Gy3zHBLEemaaYmCVLGqy6u2Iv85IWEeO1
9cHpRhqAfZ2VdE2BkcitFI0Dqz2W8o9qtgezzxuVN8yzKgWlJ06Vt/rnSi4bY1FC
v5XS5F0EgVsSiFCLJcrD4HbFjkqFy/c0InZ17Ejk1IAJcw0T0pnEbw238N+8/xwe
dMPLtjGed1JQvDBWoGS7Rlt3goaHX71FmB+Hz077DOWv94eJWNKedSCj6j+d4aWT
pq8S91nu2dZL9maurCW4mId/qmOmLPx9ulMvzYUFn6/V8HS2HEPPIQJZj4rMPvqf
Kvq3Y5iO0gLlWzSMLyIDApIoHH5jXJtrFmhsNY/PQEtjUfy3/BAFCi4e1SGpEjWh
WYZDV3jOfzLLVATRfI8yDmZCBYQBEFuWgHboyCz1S00hiBFSHwdfl+RkY/K3f2xK
aTQGzqeE9fyZHxa14e4b3Z17JLWRXFq9C4fJZPt2unpmzb1WjRDKo1/96d87qau2
4LTLpVygCJyqKzfueE/y1MUOL2oZTzqjJPO0GKo8Mwiu1fGRa99MX1Z4cugIhtgU
kE9bS1WUPm+1CU3oGMU1jqwTYBPgNdKAJ6AtjHGOgjLBPLOb34C13YN4gvJrKp/o
kb3cDUIKYJ48c72mHlQUtaLf6Y5btplioWkuhlB8fKGrFw0OnCvrwOnY2JDyGcWz
zO+MKxtIqXJt2FKddWYf/YKTRFlNXFxY9HvIthwr6HVFWVcWPr04xMFObyXUGDoz
xKMoqU8gcQXRQNl9Qk4ibfLSWianKEnEkKexTDrVN/4HS50+AEbIt8rrZjzD7s4u
73xdfNMoNmPx3Q3sMQiwG+/NV2MWYkDxDskZgKMpGo0e6WrooPyt1As12ItkulXy
3Ma5+8tby7RxOmcro8ZeE9CJhbiQ3G0We3No+9U8+waL+nRHCfZiz8riExJWexPa
o6TkSBqvG7g8104cRAtY0caBZw7sXj1xSxb0sU2WMXTeKqd7PaFvbjAWrOsbLEWw
uanJwS4LIHRrVYjNwPShdH70205Z9XBoYEAxsFBJqyr8sNNDz02PVJJblMdHQMVI
lsjUH2IS+R8hONtha/tlNn0dGCDzTw4MUz2sUcl85NmwL5sgvMvAZEOGjgc1xiUP
dC0q4R6WojNOSJnE8zNwwjF4UQKAJR5sws5SzAIUIXNpNllqdOT40ynwzg+WhFTS
7CXz8dKVyfF811UoOk/0yKtsSB2mHnpaLx5qYqpPOgx7zL9i0QyVxAiag+i+iMMj
+rpKHPkCOZf1qdIHq8JM1+G8E3NInEFhJpWq2VfriYhOnML9rDrTEWZZ47qX6XTC
2qPKIeza4RnIsMdtLCx+pwvdPlVuHTU6lsbZiUGWRwSZhW1AxCEWBe9rpUzF1yUQ
RDqfI8yby1FKWURI+dZsz+JcGCDkJHGJsEYIC5WP9ivQbPRTzqx0bqS877qeyWdU
GYnwyW5Z2AEh+3isEVmkWgJtPizM2npays4YGM7G7hJwO7dkI5Pwt2V+dAmwZpX6
59iBNmVFIPpvp4GP6U/2W3oHfiUAVpWvoXLtUZ7MQ9XZOkOYrFLbygnIf6idjwxx
i6TuLR9iWv6WtHs7wrVgm//9kIqMtDpOagfhi6BNoLRLkX10jGB7LGahk/qb4KlD
Q2xYAaQnsOLDIP9R0xbS6kHwE21ahFFSkgKI3FeusYghFKmKakfg+zaErYiqalsK
Ltckvq47LUYgeCC7JWc/HkZTH3uRSrRECi+6ZVB3pMf6wZVW7o1eV/cbwLCloFmn
zaDUE8qb3TjuPQIiN2NZIDy5R8RyUukm5Ty8g8LjOtB0wDdfWy+NJQU5zhhMkd1Y
Nq1+P8M1smve//RDfng/VDVJdqZXxsZGRmHweBxKbm7F7PwrJ4ZCUYDlMggZKuLK
d7nqtRbBfkDtPcozympQVwKLSmz1QHjJu4GZB2t5P+q46tIa9ptfkjJPmBDDytTh
GiJ0PvTkyUeQYU01LW1Ua92sy4kCFebKak3wxoKV4M1PEQIJbLBnJnwQ3laqsEl3
eaD5WNlGwK2TDTXCv/lrEBNjbmNA+dsFWH1PrfMgSG/WAz+xABSvp1LlxbXyK2KL
fjvUqFs5U7LKeIs2BLyrCbBljdQIscusDDFsqlTmLPJryqxMxaD/vbpAFa8l5jzC
RxYQ20a5tvH+x1Aoj+bD8UMRNdt0XhNSTIDnL4HodrDeLX0+6jqitYtNSLEFhlEz
PdaprHIYPvejMuoF2qlu4GQM9ghO0l1LNkNDLEUHpcWqSXi6EcOtv0w/oC3zwX/u
mUg2lnnFTCPF01oo0Iov2y2gzE01sV6Ii1dvsuiWiujAMZNGolj8d0/lAhmPdRgQ
+3zPn4XjjDq33pynSnFYO/boYVwGZrEAyZpE/fhpOom6jKSSUc6l7DEehUmdiOyO
Aj8AI5BtfIur2NCEIMnFY+a6CVQzn6cZWq90bb7xo0N2/iH5u6zFRxaLdSX0pCQO
Xlhji9PB68YMkwDR5owskWmzGDcFJqsTplRS1uBmy7m7UAfqVWEwtA+9h+Ad4rRx
4zEki22GPW6Qhi9JLrwoHL4jVSAhN+EkgwT9g7e8RLhSn+sKvqCTcLMXrmPYP+0D
ucy2HfsWJJ14WQTdyffN/vgxn7Jox3l0Y9i0W1Z5S2ss/2zwV0OYMF5lJdyRobst
bvAAJwS7mSGClrj0Q0iLk1DJEfHVKAgh2458+4asFM/v4PXk7gApHHOu0hsd6ggk
OyXkjwxuzajCv5oI9bqVLMjuMUDOGN/sK/+a26OEF8HGX5lvANjKjr4qqM1T9Tfj
AMPxlq5+lF/U2s74bA4G4w8qHvPwf8nLDUM604feNVgKQhwpt4hmQVhonvnMnVgd
61QSYHiUAIQk1oN74WPtQrTRihHlAFepCNeanaYSJhJFthf/m4FBOiW2op6HDvpJ
WUGFVve8cNnh6xic0pTkBeFU9XAANy2kTAaitdz7E89gNPr1f+Xy5osXvWypVQtu
j7gI+jp01GsTMsEt2HGqSMfvfHe98dacTC4AjEFhw3te5Ypp1CWNWDKNCVnqXjI9
V2XPt/LFl+A5TuOgSWBchR0u7YpPTJRxaPtbkVyXvDEwc7do9h/YTgchGY0Fc8hz
ElqTTZM9BzdRyy3zrcMg9SvPi1dKKzfNBn8sNB+w0wDIxI/AnJviLKBcLIR51KWJ
VE2a/2GOUrAa+CvGdk5EYOKtV+n/Wv4dvqG0XfJbsDCnmhR4nshk1TrgMn6PfEH4
4qFGAUDct68j3XDPa980l+MtQdKPwRae7oVHUNe0nh+is7m9e55WGZWc4J7Y2TV8
tntmQfB0F5Gw/hFyzv5Nq6b5L9lYhQh5u3VsqMcgqQ2JFyCtddWc3Xvx1GXb8+Lt
dFdw9K+yF7IIjcR43Yc2vA8sb/Ds1EUafhOEzxXoi+3dklNPEYshnL0BWG7/Awe0
8kVLrgbG2DRG41IVycKj0+bnzbfAuPYwfQcuYtbjtTo1tFEn5bpkKBpRwksQbCXp
ysA+pCIOuksUrjhHkEVDc1DIrLHaMeR9vazAmWRtpmX/gfh6dmuyt68S+GcX2jFM
Wh6hQI5+EegpjR3sZ6pKpu5bKDJ2E20JJ6u0CiO/M/WRC8EJfxYnxaIH33r2W/Sk
kQD6F4SorVnI1hxzYjbBr/NufodlR5thoemFIVS6rBgBy42lfff0b5MjzS4FKzlA
f6UrPlxTB7NjSNB9IrqtWMBAfSWfdqdDr68Asx0itXh1J48aC3FZM9sBZYqtfzd6
IZEeOdqDxy5nI3c0NXpbSARTK2PFAWl8bYiOhxd0ASPe/I0UJTn8UpEbQEV/i58t
pI/QOdxPcsJIQGXAsPszyxr5P/Db0Gswlo2492+GFX5ABqfY6kJsItVHBHqzyRqy
IoDS/N6pqbXGnn9RtY76Y6xgz1cnuHfVGH16b8F4YF5TWFErqkYFSF3AcVX6aj8M
lPgWad7n3YZZm+OvRuvy5TgN90eeENgAyrxccoeB284QZcYz0sIFGYKDeYWUKb1N
Xm7H0S+x2bkOcPX4RHsSi0MaAhaV8cY/3ve/hJkY+Qd4GUwsBN91RIqVCQ7lLII+
U15liTcboWirffCyGXJsLmx/kmYaq1lsPK65HWPNzHCexz9k3+6mLYy7115ewWon
5bBgeCXlR8WhgR3vBIDT9aC7aJDG61gyIDq7jGC6WCKTgNA0lSXMWeVq1M/qrszr
F41RDg87vbTeuu17QDKr2SpIlWTJ0QZsIwYJp34wvzAmGPrH+NxwewlXfF7An77X
XC/21Zyq0DSOFxsuhOP/dTkS2wQ7qwhNH0aYhvbxbWP973dL2Aw/OaE3wl9uNk5D
O5mB7NopNq68whvDdE0EpdeHiWfuhu/K8NKM1hGo0yLhwwjPYEJA81PXPcyS8+3G
Z1lth3CqopMIx5H7F4xHsPXD+MtaL7+884fGNvs33gXbv4/yn8g4RoEuVY5ndSjn
C8qC0Sn/tYRJL3L8vRpXfdSyt7MJGO/CHf0w9eUfTVbjw4PGfGBYbAwW8XpSrHpY
+H3gmMa5Jbq7146t9HUYm9bI1zMeBFClHNI11Yf6CfFq5W4ZCRhUgx3chk01uqCY
V6Zmmh4jKFUcfBpHzg48BACW2L3I6yfEHmEjCV1NJ6lYKCIz6y9aDyOFFcTs9ZWQ
m3rWqcoL1R4DUO4dNxkCCYrvIW0/wFVfo9Vl+3GuJqJj9vYycAuQHDBxgywNZJWP
9keFKty0/Ge5UzdEJhtkuNldvSW0tSbPL/aCF7p8X6nravZMB5w0/4n7Dd8mKPAo
utIWnb6HPOLT/zv9WgM9RgtMansykfNJnWgqWZ3hQxpuqx9MLBgQ1NXmoJmQ66hb
kUKKyiN/9acXDiAfhEH4KAu+iS0OqnXfGz4blAgbTXZ19Uuiu+kCjE80PzLgNwq6
lVozvpFsg1StViaZOCYtI/BtO/jG4PBHJYN4dTwPLOG0VQR4DtykeIkaQ5EbzSsy
p52U23qnlnujWoLleotWCjFoN6h+M4PSWqib8WSNOjhXwXFyTklpb+rmbtoP31th
vbZFnY71H+TS/RaDL+N6ZykvaUilcNqfqXKvT0V8cxg/3NkjiZHEC3wyq4T5DkZB
+1ZCMzRYiVJ74cxfkVkDP9swKmxJlzOEj+P+dT5JnYzom4ho9+b0vUEK2Z7/fDB/
kodKBLKUQ4LU+X6En2uRCkO9XqbwglIdpsdrS1Ny2z8SzzkIDd8j5MO3klzKMlhe
Ew+jbzHprPuBA7xjI6n6vy0bgIxVn4CabtfeMNRelqSNu0ai6S7s0fKffHHQGLs6
AZYgqmkjkp0GVjvbK4PvJwSf7gd2CAl660ti+VwN1+Ks/Jc2tlO7IFrfLPJNwDsy
3gXfWhXAwEHCPU7xZFhb2OHyZEVAfWSiXQE+ki6FKoa3zSBBkpEaq+LKNhPlVkC3
5GSQO+0ZbA40M2NpvGf2w2v22VmbnH/u3tG0pY93V1v6egikzWjCkP/GSVw6jG0b
8fp0v6sYLtpMiPmVLMUEr5VhmyAbdkK06qAh+PRc7cALa8IjHTWRsAKIPtUXyxHJ
DPixFc9FOAcKl7CIP9ZCDVaUy7QgUZvRDmVt5eVMgY7pjIWAs+D9mPPkRfzJ4xgB
ROxubmzsklHyksIvdTKwM3FJUToY2OGL4PjwxqGe3dSKqdeI2UEH9n7bNsl9p+Tt
Hr53Q6E48gJbD5SjLD6X08KcgJVMQtii2DHppIAKSlILtn6KgYMXkVfkWGSolar/
hGhH2TCROM6U6TS0B4rG5J3ZjUqGUSTDiiHp/1m50DbpgawD92rEtUMp0ZcvFxBb
aVH+xWXYMtZluhkXeN/ghF1rN1AWM/1oct10N1gSzvJPoEPSzpU/1av3M2JQLwVK
PdZeV4LK7NkBUqzsZvewV5oPxo+S+Y/Qqzm/EZEe8GpsZQ9hqSNK+85hiNNjpfgn
8D6JBYdJ12Kc7VROUCdLBwnkXZft8WilH6p3hazSuU6zvBCumXlfPoXkobCuAWES
xUl35pFDcYejB+QsPPjWrNQmFFR+fqHueKIlMo3Apx0QOXW2ZlZy9Ijx1gwjh756
ReFkvu4PZ3PFZeaxoQ/55QK8Q3j9X2LcmCz5SVOT2gYcvRYEJkv7wenq1/Cx7+rE
+hWti3LRFeHlrQBZdWC/ez7AyHtavsoCxkf+joy1vE3LQe48ckmgoeI5EdbytYEy
n5jfjn85yFMZ1NWwoUQ7QCVx1vuOnh4v1skEQvqHp9frLzrpwLp800izQyJtyWN2
zk+57DVfx01hy2tpCNeBakDnwSCIG2oB6TP7U4rN5wGt8BIXZwR0HY7payZgubbB
sh3JDcG8Lb5hWF235hIbu+hF2vOSB5HSmRIe7Aii/IxaxlXJ429565MnoiqUVot/
5moTj3H9ondLWQdhEc+qrydyze/dyig2FzUyKKrGc51WhKgRXy1jJuNaxmtFbwRF
Lel48HR3DjNvEi7HaYRmmNlCvl3yUfpW5U83KXfKuaGyIoFhg+R7DzRqybUj0xKZ
Iq3JVBmeqaBs2+Jqy0hV7Udy33u3Y/3KgN7vOto3p9rqeVHAVQvGXxqn/0KWsQMa
tFkz4vm/JtxjYW8hSiMnVr6EN5n5ZXr77OySZv3psw1me2P8yee7N1y4Y0cl37B0
BhGbytSc+YJvnJ7hiuGfucY1S3LIKZZSfLPDqioJykdDkGzJDLxBKXm1ZGkHrmF7
2MV8Kys+x459ME60dogGoGOBJ2RSaIGv1L7Ig5gPuxZx0bzs5rW9xId9EcFVLHki
A+MiZ3EAELxUHuIXzaDcfoNuKyJCUWRS0Q7Q+cmv84Pj5NXh8W2p5j4bauwikex+
EEdmZRwlMNjSbIKZCUguuQn467tf/qiTqRLjqs2RIGuKQkC98QLwZehyzTCSPbIw
OsrgFsSagSZcc8RPiSzxoH5H3zSaVAZpFkEXaMg+sCvzOUM1ARBGTySynYwcoRNG
+fD8Rj04W9NxsM5HLgpsZ9IHbO7tj3J2TJp32zlFivskpfwMr/0JvYjrBJ7sC6HQ
SUUAepyF2nHfy7CMz17ZfZaVJ4k120/3DJ0zF4snoGRYFHHHJPTsHmmP50w9/2xZ
zykmjCqV/pOFzln8emuHKY2t2EAzoc6c2diiCndzVUKlV4LHGrMXjNi1jcvrVVcz
q7UyglpwARdiI6pGtEXbV3gsbEgmHAd+i/O1beRyX7g6St01AXY8hPrnk5ZCa6uY
ZlEbtSUKfRw/ZV6fbeI5ZnYIRJ5RUaBb/fV3dQuO/7oP9TfHLgAQcZZhqMj2ywwK
q+oNIV4d1sKe/NPfXOBThRMBJcjlLvpw5xo0z5ZVCSvRRseYZnE3VRdlNCeSGvzw
9kLHV1s6PGB97FahsMr55lFRUMTGbpBe1TBTsBdCNCqBkMn+OQTcyeeiNI05AAnN
uxlEfxcapkHal9QGcqicTOyXUBZ6yFDT3K5f+xsJykdfSx1duJwnqIkcc92k6SuR
JYLGl2VYvXdyXA6XKN6AaleHlCXx7Ew8fq8n0lVHcY/UlISItw0NUX7g+Nl9bZgJ
hFEWlrDL6vShgMcGcU/JRAqlqVM2nXs1EmjsCoBdPO4qARq0s80Jr+z1Y8EuOmoJ
V84JQo7WhigXzC/LH5xtGuCmd38iwCrK3AU9+HZvP9LVIeFJ2Cx0uvNROK1nOg8l
TqnkjIb9b0Vj/m5tszAxYHdINIilCZG2OPcfLRx4d1f8nQGjckss+hgW5ezN80o4
VocHEhcO46lsAUw8GlpzLwlO6XLQvFDAdbHxtzu20HLL0EyXt5jDk8Q48zhQZR8+
FRzbBCYYg95EDp9L2k0DYeIv6TPDGRwJNFLg998mWgwsR6ZHCc4T3BjJ/zssojCX
W2s4npF9h6yjVV6fD3Y26qcVMpIf6apQF9SC+JI5TxufX6ti5gK6UHdki/aEXDvf
O3j17ik1Wn7/TsR22Vc+oBYAK9tZDnBOUAtDE/cULSi++Wm1JPnx355idF1LrRmK
saUK5fR4RK1ISt8SM1vN+72zyCB8Aux5/tGPuPtGd1/G4sk/6Aswr9gA5kHPdA7C
V4eUTulW3jLM4PT/6bMa+KjmND7wo5EV7+F5x16FF92ef/5KjS+b+LcvVo5NAFkh
RVzg8Eipj/aETqu1yGmzP2t3c3vdfk8X6APh+k2mXkWjKDXYs93yRuqzsWEaUZdv
4tIodJw5Q0ZvCAeCWksHF+fGkV5nlEQ5SmVd9W2v47DYkJH5rzJE0OwGNWRukt2d
uUAA/uoJ/vM7xzsFvd1hqaJB9rgm/n4EndNcPrc1IMJPiy1xzaWueEG1HgNaNGAA
GUfPyA1NIBwzDHXF0sql3m9/gkOhVuR+TPS4nFLruttgT+NgVYSzJFQcVdI8i0q8
HyvkIPzCwFNZ1XZoVyo4J7TYdSv1PfDRnN+pC4cJn0GMuFOmHVzauocw6r+BYBXC
M6AATQvRgknTY2P+rpjSUXET/l7MaZ8FLf7HBhQLSZNPTny4bkKGrW8U/rdVBAfo
rX9K796cH4j03tCuMiYoQ/qEKxDW4VqdUClnZ5t1uF+Dldu6SQvovoPZO+Ld6psw
QiYee1pYl3Cu7zUsLV4fbhAqyQgheZHyW806hg4uohvrj/0g3g/h5TWr+Fz+qafA
w9PBsHGPeejkhTE14UVV6sfj40wi3dsCYnUO+NaTHVN5V4MLMLfDpa4wNMf5py5l
xPRJtUGqN1bkQRBC7wrgQlIMEeVU9vrcu7S8tJ6FuJv42dg3e/0LM7erqdkqhxY0
sjHilqaE3pCJtQLiY864dbUdfFfzY9QJvCxdHUJzp+X76zrXES1U+nBgFdq8MRBp
H7JiJ63FqQmHeHcLscfmtCUj6JgWfg63UnmUyaj8ZNry2Sh+DMylYY9mOfCXz4AI
jTHMx1NAIrt/Vbbo19DCHOzsPGhVLgI+26EF7AtN7kKjBZLIK/2umlFD2vYVCDjb
ygvQl7Qd+f5YoEwC42p5vweRe5eSkG/kZRqz/3U1TArGGn1Vvrb2bwvHOqR6GHXr
92I1Ry3le7sFm5kD+STJoxDg8N7LqMzJOIduORqoTfVfszqs5DiWWVSDsgavyuS7
pFfhUYQOXf0LVnReUjzOmtdikj0DsMuUEECXjpmGFz5DmvJvs274euRn3lIjhx1V
yS4MoeB4GbynKPgt1c3xqVMfWlYo5tg75qjQ/DmclXixPVGLChN6Ez3+loyUzybj
0249vkViRV1SBeq6JFwsnZptPQ/kwfE+syI9+XD3P2bHnqPLefA+hPxNI7j8H3i2
KQi/aaOk82EzyEfN9h6548X+3xlmJPHuV9Qsqzs+Bb++2hNylwevnb1CEpbPYHU2
tCkqaanZR0tgo37slgNg4YGeisxas7pUlMbGzisiVcdBzTdvLVSUsA0UGDoxYaIz
X1rAY1Pohc0kdP112YGITU4roQqYDlVZb9bR0F9WMq8BnXCkEZtmYHr6NSNr2vO0
WjCP5DGYHitD64xivsAlE/dtn/hkB8c/kX48z27gVJaDeXZLeFMvQ+brsI0lc3WA
SuBAiS/uVOnn/TWaZEchvbijB1EYtlHj1aMMNia1xjtQnCDer542cI5f/h7OJwGN
hQd5t/IQu55wc7ZoudKt70nBJOIQ8WTogXnCw4UWqSz6+T/e+YRbDQYpDfr9K2tG
DW1f5PqMTrU93+GDHiJh0fOLX5esnp1VYBpwwpCsAkZaeBtHNVs7iAgOHddt1t3J
1k4OHAQjVta8kIC6Df7Zm5H/VkAuz66T2M5ZhOxqfevv1GUcrdHobw1rI7+eNkDO
0OB2GCC8RuoR3G6MqI0n+ESpQHmjc6oxPEbZVLqcds9oG0tLHO99mUJxNmEjqzP4
S4lwNwFMZfoIQcIe9CfqBb/6wBdIqV1vX0f9xNIlGnMaSOdlNWFbSLZAVN5noYzy
UiQEt9wg0TK0GKs8g2kiCZ4yhNG1qYD+rL6PL73Vcdb+dLrF+RaRdIJhkZrPSA8T
LOpw148O1zXJYv45dxMj2tOHn1lFg49yMEn+ykmZzDSblKNHKIIc5p9bQU8Rm/Qs
tuObpKbtF5ZDp4Cm03O20VH3McATUZ9Ww3/Ekcdacm5pBoNBs9Z3dK4v6wLoTNtb
NKK7j/DWoPgLzQH1Ykf5i6/luAp12Ueok8dUldYi1n34N3rXxcx1a+jkFjJZuL7/
dcx/V0aAFXVjScraWl/bxlgKe5lpr9EJSfMReDNMKiMyv5ahAKkrqzx164yGVe80
866hjW7104tXPcbb8NIzhIGgs3BksDaZR7qMbx7ss31iQA1eo45Jn4dFexdKdXtO
pRsBOK+Q/Xcwy6NSj1w30/u/AmXnAZiPF1fIionpTDQ9GH4VVSbBxSBq+rPD3k+m
+6L3pNyiClyXuHmzDFrP8Bx1RvRh5YsDZEzT9/mIb+WwKQUADjf7o/rRa0j21a9l
BhHjLWBKQMCa0EqSo2sGrTJ7TVag7XcaGBFrGW2q9DdduVBTeAtmcNuA7rZ/LObI
VXprlb1N7h5e3nZwvl7EXO27qoyfpxCIgJQj/WIzsFD+usgpsAPVa8LUsTK/ELNF
Zc1LTzH0dC73IEQuwQXZw2Du6+RobC9lqyT1C6NzjC62DfUak4ptR+IbEMa3TIG6
OJ3XqCipji7af1hOWZo2G0T99WUsAfOVdxy5i6aubM2MEWm2DJT+PBxpxlNuIW47
UpiRVXblqbHgZ9NsKGShQbXrsEhnzGIgo2BiMwNvYiG3I3Hztf230v6etVuzhMDz
7vFX7mAtPV+0O30sWST88t4wXZIBubDoWFVNCfNh1dYHyeq6OBO1wummQGjM9OiC
4VHiRrxYGNFGHJFWXkKKI8nYkpopYwJ+LKtobXU3IFgnLDl1MQBO2lxXu3GEEYw0
ZeWMcTWYvm8MRvT07LWALJ6dOo2PekUicq2v86wEj1VgDzSa/IWbrKKP3MvLvzGR
5KHR6IscbTPpH0IDNMbfOUpV+6zFgb+xLdeq5YJ4mlsb/6HiJJorfuDYhpKmUEuy
yETbec8RvGF4kv28wDR4UuRKhBXXJ2IC8a7JEgCPIOzDULh4tmbs7foT5VX2MKv3
DJ8JpL1oUWbuaEOGNN1wsE7gDUmd7e6/BrCLNIks3+HYL2aALbstzt9NliBubXFz
TBNifr+AXQabF8sKoXnd1bqCQOQ07qt+XQMbAdKOTvtNGvUD0Xwerpdg3rgwHUqS
Wu3wDoWiFLvVv1/kBrhJgNTJ4XMrxJMsigJiaI3yA9hQPuDohWY1R2dBeZCT6lkl
KVhtF3HSme1AA/oY4LdYFmbMg/WyfNBajDcjsoNu+jbVRv3qQ2HeeB0wcNZcQwVd
WYxSyHKY0jfSE1FHBVr/yW5JKjeMCbH8u0gOPQomSOD5fmDs+n3KDvFXZWFyyff+
CEgIXzNF/NW273r1tyjLebSWXndKFX/8BpCWPPCt9D1fFw3R6e12rCaR0lUpCgy4
vZPzqG/J2kDN6Pe86RBdKZsk8SVvVnIpl0HwE2n+1upUuXnljgo73T4u9oBqC8J3
lgKpxL0NHNdBguQ3Lh0Oec7LWaaMeG8dKmQvyt/nXwCaQhUrfAP+vCJsHAHZl7NQ
0QLEcsannVryAEwWYKyo1KQ3lJ7bAIyTh9TYi4pw7IpLyKZxKyaMAMF8ctKUXJsM
PFNSCx6ETuAoFd1fJ4SNGwtNesa8qlu2w7+0JcByws07Ysb0aEbR6EI5JKd628UG
cmWnmO/jjSy1aQP5f66VAhDJN9mfECeSZnms58HhT6qZhBi0rxIv9xCGtDV5wr7v
optQm1z+9q1NVPchkOzqGqrHROUnbIJ3+MFgYUPycuV6GoC8IkdcBEewFcBBwyCX
015IwLAlBNxzNUzGxZ8K3KgRYDpCyw0VJDkjanYElwpnR87W3bPyHMz45ptvWTIW
Hx+PY4ZxmOIZ7Xpw5H60X4XbNF6okx0/OzFEQo81tk4MVxNTJSTNm0UXESi8vUqV
7VnM2fyxi9d6rh4lIMHcpVc2pHj/T+ljfeQxmtE7qARIMf8xlO6rvhEHFkAH/KLU
sr95ebSzirCqHkOw6bGn1iQS9tyb6xXbgRXcHAftYV/JUsbWF6huFnvj81ES18Bu
YVMpsP0lobTyB6gYSyiHRUj80qxSfl9XIjjYN1M7UxE1Z4tzgJxBPAxJX2YOMJu5
CT6ibG1nrOMJNnWd0rAyfH6W/n+Lh3BF0SBSSYs6DMlEI1HgBqMRfbt0KBQQt5OY
JyQlhTrYY/PSyQkMp0haQOS2XIk2VkozhKbjoeAvTRJD01qPXI1UqIWP38ZGmLJb
p32U95uU9MPCfBO1j0s27ASSewUVh/+WQxRCtR6Yk/Yczlci62daAcfM8mn4xJpM
trbZm0087Hpj8nF6eYYABDygbeNFRUU3d3kbuUkQva3Wx0IK1HDk/71fN6JF/+wF
LO+lfU0u4qBs2Ri5tTA2hwZuQgA5e/6SbkF6jxb5zUQOzOI5BA3Y+He89f+rihK4
hdOpmmo6aIWZVFJuosg8G6Cy04XIylMk0O1iRW1qvQNr5FeJEQGR29JIl464882j
PMzEArWjY6JnEdUx3LXD2LRCCrllrMcYxeufKEIEBJ+1CmU4NR9sqNqMwncVDobD
4+WSu/YbRSNms8oO9vStWFftMLbVh1ZO6RGyXRDCgcc89H3IOnl5S5W80oXgnDKB
UIAEoG7iGRZY6KXpxXShrIGwkgzqGXCFAWbKfMv6clasBRzjtL1SaAMjWArKjQoG
YEvgVTuyYSZenSjg8zNVCn0A/1jPQTfDrsk8y8rNdKwaJwX8Ycbe4/TG257yaVTj
ghMC5zM3+NfFEeXzxd2E00LhjlVZDrhr/R8gO4TDKeKz1Bilq2gXm1RnXt/eOxJ8
Vktbu6leH0x+3mXuBtd9LT+dgUwHcJK06mrttSuxsGfAl8eHFVoeySBvDW73y1os
5Cd03Om9RVdvfVcIOVlTUgkjVs/4PX9KLgldD8YJCQyc6jX61QbvMHOKF9z9JE/g
OB/9v/+jgI8oCRtB+qurbH7PFPkDOmPGqvD7dIDhNXiNrfqJ5p2GAzRPxw9kyJEC
nrukU/dVw0dpLR1ssAw9eRg5AcARZiFoReyJoKCJOIk9uwx9tPfMKEa4kCRdecTq
G9zGUhSvL0qAhIUg0WT5Z3Mpoo5i2TVmdlQLgin7O0vcpil7Op3f+JcfSvvwHvSq
IKiXNTgrl3s6+fldsbDS7phqoX4mY03ta5DXy5HYyvY/InHOaTfAOOQV3GYRF0Pi
0sh+3qXfk72AUd7drqFdc4WYPoi7NEO8kMqlFceibkA8SMptUd4VpRoyd6r/N1av
XsWy1pd5iJCDqA5M6TQiaXM/nRuYiVhcLRKGbjUeOZJ5P2DrrMzZXoO5/XQ/lHDN
7KB3S8uyJzAepQg2zWbQi7tjG4gIuSfs4m+NPmhhI0YTMXRygaeuojaeC6tvYWxG
grms0ng34RGIg+75GHLPo1TOByt34ZPT69/j2j9tfmT0kymq3rjt4x1wUwuY6QuV
gqI6rKiqDPm5t9x+KoxiMDgn8vmJncYsAPZZn3CrMdfIlZPSA1tM0FA2zfx8vlYZ
0g1fdGxziyQxyE9o0ghy9w0un1Cu4mNDR2ABX5NcfckTCtUNvBu3tUQENiIw5Ehc
RJFAjD9UboG0ECil7dc5nqBWgozw39P/mNjs8/azoDM07OaGzZJ8rqGsfaUZdp8Y
jcBiz8zTizsPcETfiUvBo8q52XC7eBBxCMaMdbUI/jpkGU0iuxOCTwptsfGGS1cv
6O46GNgU3Ub5GIWyq+q+EPUCDj2N+HL6AXA0SeM6YPobEQVYCbk5eYHlxGGBkFrN
PoAkba3QS01eR1JngLjbZib+wxu2NtJAOdb7zo2SDcfb6fQIT96fSCP4Tkb/nS6o
MMfoOmNpN5HbOnca9JcHhuQdQUjC/seEncMI8z9d2HBWSSBMsdSYngO7D1R0AAnk
zTZgTqqwzl/Ib+8M0SnTxkuvB8y92959Zcyd/a7eG0w/hSZcZsTvnpNRovVwsd1i
mhnVPQGmctfFpEjvkmlLIZijfNyJQpQQGTTKzYjLX1/jFKm4M+1EFMPBjyLmuikb
FqphibXxNxqMKEMiRDxI5y5u8sbMDNyfkGVb36RwwqDQfh+t29g0mY1iCprc/0F4
wgzacfy8WFKAoOMJk50TEKgomp8riOUeb9EkVZuAcjUVTgYSs2XezfTKqz35Z9M4
fgLBkRsUVkUJX8v4WMDEDGgvy5lrD+pkKAJlp5Zxd7qhoxnFKMV1D54E6/t4BKGN
5X8zC73LYnD9IfoaTT3EmWXsqh6U0C367QwyGKOavB7whyEkY/w+kpwObPC8/iax
H0tix9SLxSLfT3DRCUWAyX+Kuh1sHQMQY7CpwFsJKyiMHdAAIS0sknQojsV9i47A
3xns+SubvegpJfCuXVVGE1WdjA+Kj+yfXZao69a1RhhOcaKPpHsV6xsdIxilWh5W
6Kcea+T6n3AssfLQKD5DRTyCQT5HxOi5YlKKUM84Ire0RKJjdKHrnd77bHGC66Bg
a7jUhprissD/xQSJsV9hlSbjT9njmQc2sKbj2RrusR81nm14gknQka36NU6/RAWu
w7cWeaVmAAQxdV5ZhD0FnqyLl73YyP4wc7z1Nn9ySRCLqpoCBY1FVMpJaggB6bcw
rMYZpfz9EbEdKOE6q1ka3HKujyx1d1J9oqFNGTH/pO1dY6xpJ+eHFjHUhR4hGHuq
RLz0EeQsku63bZFqaVfZFSaGtcp1kbF9aI3wtjd0ASdKzAk35s21efgs6GoEsWdn
MdHW0rGnE9s9A5ffsa8xfA47UI3T5iQh7kK92C8XBdjKN5QxgpsgXdd+nG1/n3Pu
5lTOP/K0RWS6f9DqF5DlWsqt67+LQ5i8bN6UVdIGOyxQAUQVQTOy6dXD1DEr9Axu
sKVqt56aOBMtq4zvsBHMrXOcnwbylJ4u3F0S1Oiz2p/T6K0GWXx6TUehMVQWTMxJ
xcW9QiMDeNhW8zJeXTFvX0ClvKB7GCET8RpTcHxeY85SV7w4JXdCGZN2zzvFRkCq
uChivPlMAWkJfWIEtyaNit+h76qMPBHXpC0YNFjHJkOElL2ZFvq/GgrDluhZX37m
3end2fdWWhUPM1yNORWicdcuMvTahEIjQS9jMawNNo+v6LnkjvjVb7WnI+bjZ62f
jfvsMsTTVaMVJEil2aWPg9S7S+yLJdHdwsRFqjyn8m5yu5Htp2IuazxsUrIf3TdM
XB7f/lJYNtpO5BqzgIpgruc2SE0JOUDrq/I+KebcTDKjnnnoHoGPV3+3IvYONsTa
/zODSy2NZhqXv9LpZkkiNwZbuuwpzKy5V5Tg22JNeWJUnSv2m/uGDJFybT8JKRsG
dPAVqHG0Fcfg1rGRusgoMXM6n2yef+REOdTbfu1QZSHSIVCol6bcdMG+DltdhiHy
cFOGhk5spZXyyI18QP28nPvVMdNp1mRzVvgCvv/cfbhZxVxWYMCwrs5sErwazu1U
xfv68BCCGXsCL7fspdAD3Kvdjxf7slKym2imbmGwXhoT+uLdPOGOZg15zO4t4Jqv
IUpLDDeEgdns9rSVtcHLRpem4k+2nssigNKRFAvg9pypBJvsa7u3wZ9yencDf7cZ
zkYhgy7PKNa6JzC9wIUt4larGfXA0AsSFOEhBCDdnjkYKljQla+6+bbuBGD1xVRp
+ncyCYaFKaMAiD9dY5AOQf4dbriP1Irtn02V6XsOD/6sz17U0njIiz4mRbb48BXq
40OZBD8MYG72pjCd1E9GiAqgNu0qPE8HlOSKja/5GGyzbfaTmOI7mJzHLCwvV29I
lWHe8C7usMC2abKSNhimLamDt4LukSqZJIDmwtZ4yyjAfMcGeEwAQIxhU59JUxAs
zkdZUFGKouFUpAZvvyIs041EL9PdN+PnYMfwZbvH288YFqr9+zm2Xd5r8AxbiWv3
K/izYT2Bi1AisjxQuM7sTRq5lNrmvyL7Vbb1F7TGaNt21fDGuZaKwa7csgaT21hp
qSXtrvaUgQu/FRxp/OQI9tCzmqSn36A9DiMdL+GGdNlJ2fTsZueJ7/HGZvs6KsA1
kq6n7jy4DXL+kt99KJBHZHo1TEo2zO+EBuKp5ajGsZOsB29qIRB+zfM76ZpT/crL
JpNOufsfO+vXztXes/de4rx+FmvoMWIdHxedGuet4nyh1ZL+ddwe3Ek0ykymo7oM
M4IYwYvVuyY9K4OHMqh0wMYC/KgKgWDr15rmSwFBeazvFXx5aK7pMviftlidw0Ad
3EeEdlmrb4WurhWZCiK5p9N2KaLyTbx/1uwOugKThPIR9w8x94z8Dddf6U289Z+S
1v9L1Gn4QcsGx7T7gG9SsgTPQUvJDty0+o5FxBwvspUAPHsm8Sfwx2m9dC4j4/3F
Z0vQ+b1Jfl0R6lkLR+8j3igRSAMxYAAXmTN9sLI8KgGaxLLLEQcCa5cdYkcftR5g
HeEBQHY6uSQvyfUEFDkvdFYQdtcALt+53sdZBpGgxwhzbVXrMVWKMarkgRKX9B1G
49o8owoPnBtMRx4zd/Q1ol4IpbJjHL0vT99MagmdtluDFYHkOpeshICcDSP3RBp4
9sj0vcj4Kuo+Cpj+/It1vH9GGfjx7xKGGLD0bBKUkYMr7uXM1cOIYMoDdwrOOhb9
fMTudlBtsVEj1G4i0eY6wkLaMSgqO3CdG3kPsSw7XuZWlsNmc1BUbaRcwwJp5pdG
5AsSnmjVQCDbzpg7L2kz+bK6QRmNhXa2MFB02B1sRvPBt37BWSZg+WPpSRYSurQG
PiJKsccbcYDTjh4RgVoUzc/OdveZ+0QMGVUSl5kMFB9tfo7aofuOWkD09eJ9pdWL
RQWF27TCeuZZYLRjbklMV1Tgc6a9JQlYnGATNZrT++Of+zTB1qw3FGphpubGRpiD
G+QxT3dagyov+yT6Vfhyc/7jSMQMpnpP51wD0hyqCeIgBpV4gROCTiULD2IImhRM
10KCAnyW1QDUeUy/Pbh+SNRJV5jCDaW+aNryyez8v5pnGslctgYv3PwkEtipZGJn
WtXyz/FJ47KS8dfjHypnJ0vpeRp4zBU2HpNB0MhUxHwUToXzDYDv2WZEkqT75uVV
v/oRCNPpPwkp2kQfUoqMCmzAp1Uy2ilLHqUqQToFGffRVdhiZbn90E7E5QXogoSw
pa1bz2b2bPp/aSv36xD7Y7N3tyXvqPjNt6IGveV+002A6nWhwDoEuVGjPmqIhtdL
yjZWWBYH3mJtZKlz+1IswL2OOMu1KpDL2Rk2i3yfvOfSAEMSXcqa9NMxfrJs7riz
8fbkyREG2spoQ8J9aWE/ykesG9CsO3FwCnq3DDxBilP0uY+sc3tdQwesvcIB0WbG
Hdjy+3UI3JtEYXD5jQsPQvqKrOgl9hHlaOxWme+Q3ueiEwO3sWiCzpCbVtJAqiBJ
fbIZrEPNPHDGlXodcSQxK+nbA3HPX4uhcjsBxH8uuXnYF+L5y6cPAzyzkX+EbuHd
73/L2XfMVM7czS9fzocKV2xiBK/DRV0UMA10Us/t62+3zjdlQHi1jhYF6NQC4uWb
ybfHb1gMacKxFDIv6HIuarJTewY0fcxjwrv4Gn7iifWLFUHtjrtubhfkplrTKl9v
4ro7sikd2Ro8iRPSzKGLS7xVDvN+r1/M7bLhMM88nVRfJqQq+N8G4cn06Uz5y/Qj
puhcl7qw4awdW9n9RTPl4v3UhgvSH4RjnTLz+WNExPembJ6yyFwfyWOHd4E7hl6t
NMU8I0g3NJIwvfcWcY31KeJ9KtlPBIlSX8cqOePA9j54klax+wVsRpFxkTMYAW1z
tBpjfDT9zg9oVNWI4m6ZXMFucSpB4QNP/dwDhLe4Fok3/ul1gb+i3yRmpmSj825A
l4OumP6MrBarfoQxZh43nlbYSYdm2e+5wiRzjbRAwqQW0X7xu5l6THMxq9taqOD8
v6hvE6bUWVzsvpj8XXG1SeaCyvBb4UJBD+QMEbhYcz6exrTtaq47YIZDp/LKszO6
ZIYWI1PFAHKMsVVoinygmvVPXrF4isF8b/q2u6aFvWSaoLuYbyExjH3RjcuskUae
IDMxvCRU1j+8VRXrbHt5bjKVnhB378au6BJsxdZNR4P17vatm2vO41PivXHue4my
aZMpoUG4oXHsRaGA2nz2K1TqtWIny7V3z5Ep6e7fef5X/0ENgqbCfYBPYcSHnqjl
PExooSjArsoUAmP4e3n64fgIDoum+ZiFZDKFc/C69NL/fKfnnjFnFOiqDkZB8Dxk
jvqtvvJ5FH1Ts86lGq2rcQfuntVmgDAUjV9HE2+sG0yZ2aHDO/0u/u+T0z40wgV3
dzl/tYW4sSgPwGskLFF9cKz/YJ1z32lEweL1Y+KbHoNfOQ6TyzO1RTAX7ZvNJvAs
qSZgxcZxXHG/dDjqZEX981+b9NaYNEw4JsCpNoBM9S/dbxo3LAb5pLoNz/+Q9qhk
506plrNoUICHH9sarwpJxqjRjEUjAFMAJ9RokgNCAjTM5dfhA91NHl0SHPeCcUXd
NqTr2AMBuPgEpWGJzp7dml7RNcVFsB4lljAQan3Exw+/UeDobFtFcEhgVgMOs6dr
kWCzxrTPYYMmK52VR5x6XAPfVfoud36snhBrpcsabu8k5TjUu8/VtQpSmp8FTh/B
4QqQhk9lrxkRl2crVA6Rq6RcuyNGQ55otStU5tPQ63z9jfss/4SAybCz5jTZ7ULZ
oTVYzZOoOw3e+8BDPNm1BlTkIUXdvw94ecysN5Uj3bSxbsxsa/p/czpeDUXoP/SA
9YRlLyNPiee2Z+Y0r9ft1jHdD5RllfJRR/xUSwmGfQvqNvaBxNK4TDLAy9isQaOt
CPb+2bb8Qz9u4O9wxw0iqXLdBBamEe0Yf0KWGk684iqGIGUFODbz3yfwu1spdIuI
+zw1UyBwH4HM8uMiqk2BJ6gnB1lPkbc9JiMcvQUuoyYWZEfiEow5NAnm4kLhUnF5
WaX1/fu2CT5vylMh/jNSxU6Wl+ZTsPHvb83cbYIIoBAM2fcGA2qfDaNW0tu//RxC
g64n3Ql6H6bJz3Twm3GxL1oyewpy0iZzPgtNQCoXZGLAR8F6SjXPexwN6Wo6fHO/
QzxXPDF+CcMjevwbsngtKMA0cN7aa06+Ieml6557yGVgaxeZpygDuj0nan3B9Xye
qlO9Y4NAi04krKKCmk1xRVJO/33+f96sfOHRlipYjDSpZvQTMSY0TETpDXn7xy2P
NtRy6InQDyO3mHt6MAiKzXS0JBK0noYu8I1lEuIU6uUcQ4ZGhoJWE3QqCFmpBzyV
LvIEjljaytSss2JA4soMvDXlIPEEtDd1a7+ZpWWWHprL/8LMDSaqTOWgTGe1+HeX
OPiSAb+FbrDtyTShzspY0lZgKVv9skVl1AyOWlAaI8vLsRm5QOC6mBHcOrQW4QTU
+7jbOH04zuh1BdTf1UV4Ay8Nw8TRcN395nHOvxaOWLv/LdYM76ZDm5xJA61HuM5G
iuyBa36zDAkGlOhfPCHI9G6BgZ9DusVf9w697/kJPVjZNIDjAjVLi8pSyuvmf3mJ
/2rMXGAFvvkVRtmUeLO8r1Z9J6Gad+A3qCESH0YuO3l/ETQOwfxXyhfBviHRJ8Tb
eI/0dt4tPKiTO2OKBz4dOoBHfr/teaKZw8rUyEbGEzOgVYrBEO+yeLKnErM2XZB3
YdNa/mw4b/0m89Kl6igJiEqLFykKfuGlGgInRIhrq3LunTfBMoW33qrHYdoSVMHF
1Ug5frwH1+0QmFQMbSiqzD6TQAc+0cqH5QxM/tZ/tCew7BT4WtiMURu7mQJ5IyEY
klJIIbnS0imXsBdgcGgDbZAYT+MVUCCbZXPU+SE29At0FvLi8rKQ/vZFkJLJC7w4
Xikp3p/FqNhcSRHlTXhhZe+aotA0NPQEMUdStGlt0YGEBJ9PNERrqmlAkcT27OmF
whkps/Xj/vXGkn4HzZ6SaeSoBoobP2NX1fr3MqjpJLQ4Ch3T4OcXyiAi9B/A/Q2q
Xoyepq2Ie+rlk8Ht+G3w3vRkk062Cgx+RLgZCmi8ekaFYYK+v/4TiHb/5FvlzMvD
He0yTA4E8zrvttY8q71Y++jltO/CeNpiPmOGVrYpczQBlXTmbptRUsq+WPkGw/xe
8Ed9OAJVznvbLW5lZE1LuuVDJhe2BAIzFy5Hwtg8Bqy5c39hxIwwBhJII2S63ijq
5IG2QNuwNbbpk4pNKVDfnOU7IiaiTYOuHcMqIdXg4KBbdcggMb9ILpmDRrGzeOOq
S5uq1dUI/itJKyEb3lZk3y5YllauVVBr3b1FFlLTAB8TV5jC14f20RuztN47z19P
3Co9CYkidMsbUH/ZPoolds0Bd14GeC4NTld0NG1105LDA2TEslyw5Gfu7vUqz53T
LoF/PoBZkCHSB3RjGOHPu6zNuT/tCuSEFThueo+iBNbcuQqMk3a69BAQK6JamoAC
N2BpaIuSMq3WVrVKpyMy6sEts0X5n2evixwiOGEk3peSeo4pDBs5XG0UFeP/fohG
Bx5ow96sMbN3vJN9qWNCgxzwDG2/DuGlIkgnoQFkeSuXpk29yUkUX5HnYo2vBbSs
rMcx+t1FVty1lfmBOBm56TrIXqjgo2jinsHlQVoC9oD59Oa0JuHIALNdrKHl+hvl
orOk1HJULU2slipTJVyxA8jWfcV/aBw1VSc7pwizvEnL0VNa94tF5E1mLUc5Awnp
+eN1XMJaFx+pu07pmus5dThIQiR6tkDxoaCn01BdxqS7I0ryTNgm86HpDqxpo/kR
35patFtmyfdcGASC7mn4o9be1s+1hCAoDOonJtUCJTzx6Cc/6TG5Ct35e531X3ja
sg/0NV9UZxv0SidQK/+2H5tk9Pb6UDKBsGMJvj9kNM+kO9W7Ipmn5rQaQTXFP5pJ
xLfFwVYZhMjoO8Pi9FJz2LfU0EByEhZvCl0ASpF6KZNFCk9ZB1TwkXmdHZ3xXQ3B
kfK0JxUXvs5NF6OQuEAQkIR5vfxoO3q3wZkykR0is339UwCaAOA8bmPWkECb1pIv
EqqcHGABPu+qkGoN2ZogaQ+T+uGrxLvIBSqptelG9MKuX/KIImAE9QJmqCf2y+tl
hC42vk5qIvHrJRWTFwvf+4nG2HG4hip0QnNRfUjB+9Bo25kq3YFk6zVcRieBVBEA
dHRThJig1GKSniNG7PwWtFXF8TAW4fOeljxdIsd91u7JBn9Gw6uwK8jV4aGTfJkL
N/o+ixACR4YZ1k6yKHTBAJVQiOvnFcPnpc4mFupNiEclEUOsXYQAJlahzX41yPVr
8RiBjozRKSFn2+0l+HZ8wvO1fpFxsC/vSSXFIai2330y9rcg44r9wRwuXeVdbaMc
Sthzxakh6NIvijTW7mrEZVUoSsN+2/91/BM8DHmHs3f7qBLns9TkqMu0vogUYX44
7n67AX93YAQfWj5fy9KwRtAFyfOnyR0YGPJmhqR5GpWWGMQyp0cCR1pD3Pwc7Fz2
ekXdGYKbdsGjVTWcRNvamtFi9djjvqO6hqkIJtWOmxzw9ZVhopsjescDN5s6jhId
/ZuqkQkTGUJ7Mhaq6RpESS645lZ5g/pDSw4vTmVyHNJs8oeYssBroia5TUiWW/lm
21RJ46TmFFqweyO21K4kbMtIPePjplZposN3OsvjNFXZQVnddaPXqElHqHiJFpUj
s2HM4L8lF3L8oGjWcC6FxjNOPSy4OFzps+uSN17ItrfLPjItzJb7yYD5AkIoNU2q
ojSAHuQuoQKNy0WIpjxjSvr2x0ZWz7/zIWpE+6p3nSdf+u+7Bi1T438ZIIFY/FsX
KN1DldF8+/dJ+QkM0eBxxr7QHCKGhRUhJwQuuLhIYZeaM8PS0YKYLgXhJqemZGNZ
6zLicYZQki73TUNjw4/h45HyS4fr97JT1P7yltKXappz0hgeREUgB7b7qcjDtX8C
o7o2+3ZKFhnTVBoBBGSJNQSLF2G2HB+8vvECpFwZuHMfNqMzakTxDTTWXjpkB8PU
dCfCi9k7YJ28M94rRBc/otL5OA5HnPJlVwKJwE6WYNYEir20Tdw6SvKfqHsT/5xz
nbRiZTj1N1VEFwYH3DplYN2ZjM98B+r9fwEFc5oQVRZJrYX8GBUNc94WFbkw/Whv
LBv7gu5IPfEyb080I8H2l0HOPT3htHQCMKh5UWqAl/KIzxCtPTpNLtBejAXojQS+
7ex1YjsKVBfzrAZ55nGZYiVnpVEgh6WxpUsKn4O9YefLA8dsLnIHZ0Pvlz0J/q/9
5pkITbVYOv4QoHSY0tu0zTif+pcuxJWiNCmEWBapRahTTYiF/YiN4Ivu+Uk3sgU7
Fza4y8Q74KK7jIqC5rz110vpWz/hE7yZaQ5NY0TCUbUdhWFBrf/4b/IhaAcaciJc
Yyp5ONwX3u9ukufWGs6LivwDJo/Y/B66SAlYpxVZEpkA4Y1RfkvOFO8ok4UgJgcK
Y1AEyHPU+jqZqF1ze2xR/+R4d+57Ju5ZTZsRo5zWQIh9yrFUHTKhKfqEyiS8myJ4
ipJ/YagIKHQZs8H6tTqd7VOS7TywL/EJeKgW8URdD4fUW7sHVdEJ7IXZma/WkNXs
hILP/5D5RQmqOstTPVL90Ey02DODzTTfmcJW3ssJfiGJFJ7S9PhJ1zqTaa3+FXio
WfbsTyF7/uL6tb4uHIwfC4IDauWHdiXX9XdjJtNUuLglIZXVC2XjfVSZRctcck+k
vLrOQUOBz3ZUDmfOgUTHwrRWf4CUiDWThtybaAxJkTfoZHAKaK8ekdIqDD3IPuLF
PC+x0jPkAedMMf6PoDav2kOErMZazrV7tCn4pMeeiZIQIkq90IW+h0GmU4KWEI4/
xYNwf46BKJ1nE1t8aiw5RtSqj5aF4YdRQlbp501DTS4WyvN7XeKuVui1+dVZAN9a
bDzv8NIh+NLsBpanDoTILfdQua1a+mrb1Cy5R1Lc0Kj70dHxZwc4Rtebpgav/1da
gqRmzEbg3MGtKSiMiHXwOtZXcnZ2Z9DvKCjmaRUm+lErDcykwDxvLyvAQsqnOy75
BQ8uD3SSLnSTfVW6IkzOJtDZ9O99w1gDtzf+rEd8+e9iWkFYHSP9etxmvCHDHaF2
OutJekdBaMT2QCuZ724hux4hbYHZczaCQLU9fbHHWytLFoh09DOMTIacQ4mfkt/d
2fZWshws98ajYmmcc+MMqw9NLIwgnl4OnlgJ0xoHnMhCbsIAfx+MbhsK+REctbky
5a1zVw7PoXeGh6XguUVAtzdLMwNd7cUDK6qF5lJ1KqhkcIrzno/nYt7GgcWE7An5
tvikutmJgkR9iTCEQYpS9cZvYSnMlHk5krmlsc7bswqcJK8sn4HQq23MRNJAJkaW
N8ne2AU4fyu5wmXoPZuunOyRKby709eGlch4PGarYLER/i4JVLXRppfxuj7G6a+F
Rrd5AfyWe/RArfvxfHD3yGx+1yAtsOfpEIBaOigqYGHlrRbuwxFEqjqQf2TPQabS
fylPj8g0v6BK5gl6UV6HlXJjI7xSllV2w6yxgh2TIofRQb2+w/aJk5S35BrFu9lF
KUqSggfj5+H73m81x7GgkmVlnHxGXJeLO4nbDKSG2vNZNLTEPerb3vqrbp0MjnGi
G8+zmvgUgv7WvZdkrhOrlpzuYoFyRuCPOipFhD8WdaDgFCMjQHHlHQQCpn+LDfRq
gbI7i5mr3V5naYPktuYjELESrFFf9oqMsiTx37qosMLN6DZjcsxndMj27fcsYaIt
JVPQuyqq6yyN514LdINLr2ewVEeyI9qqWbJ3CoOOKNZbRyaXLCYscUD0AfpFsV63
mwRhZlrDwUbtU91ZciOjg+2VcDcOf1zQtL+5dCNXD/UrqVZlyxojBWjYH3XP9KII
AxkJp8lVdKKzAzu4ciCAho/JetJyOrVIpIa3f0LB23BMemgpfi9nbrnsa1TwJ0fj
1lnKqDnjR21Ra4IO+bHL2mOrXTyIGbymaOiIVY9UxJDYz5BP8kAqgAZ6VtKtDYG1
uprFfM2Y9i1vqnor9XQ5wpthWOwbBgRbRfrgVbFjdkUmAPRoBJwUTxaNOJumS4vi
wfbY2PVfzXjX7EKyAGMVL63pbMQfu2Wyi98uxxB1s+z3rEchsVzC2F8zVrNWuRBV
LhK7FPtfeVB1O7KQad68DdusYwIpcjSCAxnM91kfumXBbSa+iBubCnPI2cGfxSvm
HThdk3v3St8dk/Y8CccKXk1SJDUbQZsSLwHd/xw/D2MYYXQhqHAjnW2WKdniXN3d
aiJzKKUbmdovfk7Td7Xzhuhp5zLFHdOcHGsPG4XgXh0lSaGnUgwNv+4SqWFzPwq5
x5/TOfqxujzv+vC74Ahstm3TFEBTH0Sn/vKcezNPRDZ8rFMjJgpqyJLihyqVFuqo
hJBv26Wq3TMTEoTM4I/13g/otY0GKgmfu2HLx2k/3e42yw1u+IsLfT87NgXdDeN2
GDnCZEE+LkP9wo6pNJV77PcnfwSY0vYVmpZJWCRQSzOIixX+7U4lOyh/kcrxJHBW
424cdzr+LYinAWEhaHbPltvENTMujlcJ0PciYVObbYyThIcsu/XJNeNX6tSxI10P
Lsa3Lp3aH/xUlgxC/wPAePxUL2cuW8hyPvxeIhDZeMSLnDe7aYoFULmbk1JtfZEc
XGyZSyETj3byCehcZkUnUF7EXm7t/mgMUAIK7JpQMnmzcPaa3a6QIUGbAlyG9lhV
8jz7+xCy3VtI1c5MhRgg0imWVU/GCBS4xiLETKtiZUbwXnUrO1SyrJJndrY3WG9B
gILac3/m/10kk9R7KWtpGj3JYSYxWdlhYiFYOPeEB8JWdfj7tmZtp8AyK10WXqQL
V1DHmhvMKxnB/Gtwy4GHfxFj87ShySrirYuiOlxnTJYI1V2xxyUUX98+Ve//TZLw
y1LFr1bP9O2v/VO4euOSChQWISudpQcDBdjBV/isgl6b+pRjK3d3O7xK0m/K+G/2
xFro9NX3ufL8XkQ/NR04jpkWXpOQOTLlNDXHoRNtLCpuUAEnnyZ/OYE+1eDoAHwh
jViyvlq2o+tBkwEVbSY/n2ebtnQd2CwKiftlxSf3ou5dVbrjS+fjbzPBdIiPrFJZ
b9wNW8L3uGIWbz3Iex4TDZgminCW+8BAL8YeF4T9MIML9wnrXyRDokueZ7dZq42E
wslhGa700nej/Wgj1Snye/bBuxztFjATs9dA6RoXGOZ5+J2FjarXp1DM/ynhLlZa
XhAyQduMVoB+W8PkwqaTMzPAtQ9AW4KQlE/oD50iNLk+LUCubK5yXzSBNQ/wMuY+
QGXiVfxge6s+p0L+byPVUOnBcNtnzjrhgaZey0qggx21Q1Vxn23/1OLieQEx2Jb3
L1lqLj42xvDIZhMdvi0zkYa9mEkXM0gvmxxPt6UjdnLwzymc43LdHZuhWRQwXJDa
kwSXVxQfBKL0+hyaEA0C0Q7AVLuXrYvgBP7QB3oJmHVOy4BuwG0r9R2aa+mhlzeg
MrM3KAsek41pY7sXPWS2vR0S5iyhrP9GMwEPnecUnLezTslvFyA2bksSaQv0/vyl
bHZU8eZ5WIiXhILbmSP39x8kYkHLVS2GTka45+OUX5iHqE1dylVYoGhH5Ocm2Rjt
aVVRX2o+AFGNLop9tQX74wCQy9FGySYeY3lqRoH+uNVn1BeivEnc/JoYEnfnkTlY
Uu/PtYYhypZrcfnBbFbKJu3msqUe90lZaH8CBzvAgYHfh1212e7RaXwfO/0uMaxX
NPg/0Gw5YshZzNh4HGbhStDcJx4o+kpgsqTNJrPGTVSeZ9TtmUV1tXwfy2Oxw8Wz
ITZeAblM0GL1xdDyZwz2MIS6v+NrsS+pZ3jn4efnga6OR+VKb6xKAdW9+AOW/COR
FGwLSWSaPhQqKd9KhRL1Va+AoEfzTaJedq6TUtCesj3A6p5kEIlccGtUz0Svxwe7
kNO/O0KcRQJRUyioW+UQtWcMkzZZaiqcDixUuY66b+FDH9miRrMOR0eZOioPRe7F
Ts9fxAT0bFUV5kjxlYg3Aj9hzDOctW7cl2opr3D3HeV3wH1suj98e7bpFYyWj9Nb
vRnMF3jtSXQnbLY+ZtMtz/M3amh3oLHqpxaWR9dtOyInCRSzCnRrDd1ST44wvZsp
9GpUUsEtis+QQ0L0yjV/mtyM+RDb3naDLpzLeZUJfc7dblTKSPKTWtRKnh3Y4a0D
ftIYLu+Wp/pOLrP498DbtFxmiXFolw5VA+e4CWabGiHTJuLTwMUWnVRnSwAKGHoG
Je5cKJQpFpaBSTiAbNjfJQY8uFQyLJwyu4fwsktRTWEdKMgwb/AMkb4i5vVOfJtx
p/ngCUghGM4Zeq8+1ASZkBzL9wNt4f83Av36KjMOOeT+hgC3Hb9W5D70+FlgNcEi
HeWsLrGSOVoGG2CyyUOp5ElF3G2vqnzhkwjlm01RmaF/LyycVSG8HfLuQKeMhC4X
pwnQHpU5L5s7HOKnP/Qn5rZqe3YYe452unpUtG5WpbSku9mt+aDjBeqgUGe0yBtU
R8Mm2qKUmeW8JEX0tJuY5FnxzjdpEkauETHLcdnTfVyKsA1xB0pXrPDp7W3c0P+h
gl5KE4hcPMReK1xcyeVagxv2upOJvqed3Gjjt5J/Bug89NaGNeaE0G/bPXLeggZo
O2WeQ+umHXnGswped060A7GUrCImtuKiE3tawpB3tAotoekBXVLRU3hcGWdV3pys
8fK5TZzTF2CM3BQNxJPSejsCDoT4n8mvzC6LsdTPCDlGFqx7HXmZ8EpOdnYtLPi0
9R3GShb0OdXqHwLC10yh7Zr0ayb5uQq0XK++VBGTdpdV3wJFxgFaAG9mxzFPWPpJ
AOLZbGZZA1sX9r7lSXN2G+Azc9K7kVG96U3qbpWPXKl3WFFzqJ2x2WbE8ULTfoAB
UAnF8irLvg/ZQvPys2ZtObkMMhtoqQApogPtNOkJji4mcUPlPqUBZN6Ln1hQJ5w+
Gkrw+7MvSiu1TwcNbnEcoFA58EZ8ZykMkfxKOBn7dPgdVwXFNwux6jjcAI/Fpck9
IwHTlJHxw7ZSpEao9TJD+8fiP4LsuPTORyGqfiCxVrM3l4+fCZQ972vn2O+jlkfu
5mIG7ni8t+/ahOYyoiY3DfueXXM3pfrC9WcDZ118o6zQPz7hOxgK3htaP0xs3g3G
89QlJZE7MPpqe9f4TUjdvtguR2f5aw+WW28et2ERUhVdOBOUPb3B0zd3HpXRyKQG
BoRHEprjcp2ZTa9kVZwVOhCWFWdonkAQV0XT65MI6CmySnTOwdsWTiTYACAZmqN4
QyQQAUS8olcAkZNmTLnVYskxC0ahYIhnHyaQD611X4LIwA6XiQ/y7R4rIjK4EUA7
q8yOdu948CPd3efxgTIYspYyUUiYySc8YHx2taVq+RRV7FaI+9lp5ssMHZEvybZ3
QLnCOpex/Vlvuwt3M6NpEudLHiP7UVZjJSU60nIJf1QcigBdWphrhKDPuA22oSMT
RnA36R/89Fh/UY65JDZKM/FkRoNdcgWhSniJnWIo7ZoEJNBaEAUy1D+tWsvE7LyC
3tGUsiJc+2yFYHRmYrB0kq3H+S0fvn70A7rb5YmVB6CBxC3OFYX9zpC03EJ0vb/n
rQz72UB8b9mNcFoMLxritbUdVAD/sdjOU84LNwiXFsXLtJec0xMkQgzIOrGR5Q+s
qfQXXjZWiaTne3pC1DrMzeJ0M5pzYPC36maapmdGT+YXCzVk7Q8iu+vRhGAMB3sF
G7MLCsvPT+EqUZWn+dlKvRtRYnKEO6eWw3IlkJnuyIWdQtJTdeiABoSMmMmrl97X
W3K3+VpUYk1LSQtagCQyzJoQCzs/lrULTwH1+i93Kxwq/E7GwN1t6bi1bQNrI2EG
3RJ+zxC9UlROYY3vN97SkohQjKOjRF04dDkC7rqW4gdYsPcBaPYABwVStaREK4Cz
vl28fvkm4yGHaKB20EHIYp1yqx4W/7vsaqbmTWx5w20apKqqeq4PkSjI5udzUlXu
QNGAi7L2ba2OQJv7ieQaWzebi2jbX1AsAXMW/KKOD2hiIpiFvbNwpXRd8CCq9uat
MzUmGAP6vubfv6SJp6769GiFrxM4j8QUZ9rxBe6JaFmpGRKs/7p3tn37q4xhAs5k
MmuaIN5gcdV7U0DYggDso3cXSEtwLZduWBsf3ZFbRkTMh9+IdfB265vCMsZI+I6d
7gBksmo8iMJIZVto8sqVGzcalJEupegnohBg/yCP5ANK+RCov5XRdHQUhGdAEmjs
mmePEZ/+khbnUICSmAuRIMom/MMd9OcVyvUX1TGHnmeWMRIl10Jn7DvWm+tmpxae
bGPQbXHBIROwK3EwiJW5oLcaHjq7foALLZEhmKdgfeniZkSQf7iffCAm62QpwYho
spVXRLUGa1g1IRm/X3v3zI9lcSiiZOiMOCojcgvbFmR3qF0GeWjlnwRrCFB/cVTY
KtIm2QYv6kRD9MD2760qBIWCXEBaKiIbC97ab72lKyd3x9Dh3vxpwiUGKCv4JtKj
OVJX3MUFt3irknxpGOERdCz8Ml/kHhkxBfUOS6+nZf6oBD71ip2YTKuvxW8I6th4
QnCS53NF6Q7HOB8fITwRyTTsk6SB10unkTARLcFI3GR2v6EycIQUFrt+W4jK8vWr
0IY3Rij5sRklnafyHG+Uv7NAcb8TRTyZTAROohja48Z0NmR1T++D/Ka6RRponCgm
u9Zp0gchVf42Pebd3fUTeufzrD5xXig1BE7Kr6YwKOSWf0BAYlW6siCiVwG8IB8H
9dLz1fh4sutiiDZDDpk2Oht56Yo/W1OIXecgQj0oJg336wEAhFdph1T3F0teGVjp
Dqox680iQato+539xfnzACLLZI0AietO3ZP0wVR3jXq3bemMxDD5vhZ9UDLVYUwa
rwZ9IqkZhTJpCJkVt/H0eeWJkMDY3Lgkvrp1+rDct/87aWaRJz6pcYITEBcMyrFW
CL2YNlR0pPLnFlszmdHtML2tkfOHRHBPoy1x9tUatN3V3ZFH38TvfiJxXYv2u93A
uoiozxw9VlfgiFs3cF1/PB+a4JOSLqAPwwA5AhCiEkz9vQfpviZzL51tmjPG6vGO
2l4YZatSjIMDE5PY/oCfsS28PfvLv4YfcO1j/5aMLr18V6xS6B/76FP8qdQBCp3t
Sk2OdNRlfr52K4T70dFiI7ablGN7pJIPMBweN/mugMCfRdEJL8uOP1oVDHsz5MAI
3iE5nkg9IBD3FF+eifYXFAkFqr6C7hX4h2/LEUxL6pAU2sawFkkdfLIq+ja6udh/
nqY7mYo2WafWbhRN7RVhe1bN8vxNFyELdd6WTENZjCSlJ47xHrj48qm5miLVMxkN
510VNQbu5Qjre1Hn2ILfnqx0Czb+3jvJomW15iC7U8j91yS/xqEeLDGy4dRtt4oA
MDSOtv8TV0O+F1oRhPNkDlVVW3Uud0rqx3RwOMA5Cq8r3tT6YNvQqKDAjVl23D5g
qRc5EcSyCekMsVCvDvb38f6hIomQ1yeVjSukerwtNAnsXRIWDiZOvi5pIp8DnzjX
a/KEYjuY5CR3M3iQq1KAyAw0/DmuGR6Fsc+X9tdM3Oecp+cG6Yohzesomst/thNa
kPb+iunCYXiX/xAnKQCk1+SZU7McI66F9R3vqWfCUIBp8/hUhxxZ5YFLK1iSGiYO
GgoNvGBY/CYMAiAy30xcD4NbK7tSo1PE2YTT3mdFd7VMVI7ncyXtUZeU7la4qmBa
nx58PCnkAapurwuhuOZLXaPDPCI6VBby8gqXZADaOFendYNZ1l5DqL1bBoKlVXFO
CaABYqkp/DLh81FjhZtnazIyjuPthNrZNOgTmupaFZZz3bBO6G3fR84gkYGAJLt0
7TDT85872f4RXDYjIvAfkxeZIYcF0ZN3nDUdcFMjEV51ypsonvmnLSgVqUDytD95
zaYNC8oPWnbEIiLEPBIgkn11OXhIKgjh0uDj5Fo21HM/hv2eN7FRlW4bC12NyQgW
dFn6uSQ4aJWYnLic/6LbcUNe14YCwvmIRhzximlvhlG7uUQJnB4pImua1REwkI7i
YvabrhODkDiIitmhtTwbT/gZ2II3qHXEpJlhxQZJCLoGrtgFR/5ArwOy9ioFvooY
bypTIsTLgSiwESJV7A7bBPpwXWo1af+NcYK2Pja/BweMtj//32dVh+VaYciLtLRj
jRO7kC0yA8wDqdemyQDViv8jQiY3HR1ODL60oum0XJW9Rbxz+HnN5LzsK/ChX8k9
/IQGUoEmaRAi5mbx4Nq5vgFYv6GKfWMZmbmDktkUp+3+R1kN8cf8300exnYn5JSl
ct7Ol7NqS6dv+KJjjHXAsej05tqZDnUVc4oaMZHv0gd7Omf1BR0TUZV7fOZC2M4x
eSCtS5hDit0M5SaVdfWJlXveMLJOOX5qikRYnEhGZMUJP0uDgGM+2Bjj5wA/H0an
xBM8gtZtlblNjvXJ5xzZO8ShHFsznfiHi5vN1QVkuCXH1ZaSROunP6o0flV1NJdi
5aaG0ccljmZ0kfybFYbzRSOS+yWkGxppuErn1CInUceWKilxMIDswl9K4sUhux6q
VHCoEgoWfLy2TT3ls+kf1GacIdN1Eehcr3rVSFax4S/LLDrLBRM5VKeoqWnOjejb
+UQcp0Mq9hstHAaAMsxj3/qBu5bk/Htgyq644/yP4T23Uv3G9W2McUA5TObY21bf
Wizai1LZ6y+THRhfZcCRvolS51R/Zq5P7Bq8+RBXUcChB/RUfgwy5yxDC69PBBmS
mC5ACsNlLKZzV9DaDtCf62yHTK9Y16/ZhtngWWwB+smuEGR6geOhYIaxKnZAvEaS
Hjd3cXO8v9h5zqaTMUuS7as1EcgUBJT7DSaF4cHT0VMnXYucDSJl60j6T7u6F2g8
F6tuOvtNVjuEtFuiWD1lZ0zHwSDrtCxUnoH+/4/CRjWw0uyfMFVLjY0iUviyFeIC
LqnF2c9uiw5zAnRSYWIM3IknBS57bpLaN2jq2PF5KsKiNVVk7G46elRuGKY/8NZr
Yz9GxDCZw5hJmF9v8TlmeV1lkjZ0xKhV9eENVeNWDu4wxiI0NW1EumUAyG+CL4no
khZ17P53WKJhbmweVFGxL34HQvbROcQEkdGsxvQvbGHnSTbijpKa0NfkN+SkDXLU
O9MTDU1LyyhYqmLmTcxA7PRRT+rjs+9Scpwqr9cxbUPxf7y12qJNHkdKdSHfj1uA
9ijN1gBm4aS0gHoh++Gxv8M1OkESBhREFK6s1JhgWV+/Wx2NN04JAVVryLjwgKow
tOH/2c67Hz2+GLYr1fFlo0Mxccjfr+KJr0FTuIf4HU/JfQ7APuO9vtSrEo29BOFo
4E8SWsDPG+cCpCs8H+MfGscM5r0B+9vGHGwutTHwhfxqBfIpUBupczxGW/7Xm4pP
UibgrNx3XW10McO5sMyAc+Fm/0F1NBANgXu+3mM84xjkxmIfdVt970i/+7TB1RwP
2YQ6JcFSsoFqYxDV0bciUWLv1+UNrURaaHOHxi7OL7mBFdRnBYTXuZhJ2tnrLYtJ
OqMXuic1HL8DzJDJYIdmilyRNnYum05thitfh2x3wOMj/pwCNl3Fa/0q5ZDQYi4c
dLlNNw7zbYSgMWj6SZzcqsTacoTeDx7A5fchKxaIY2cRx6Jtb/fFk9j77o/Zd43j
8o5kw0v8+M5hBo+oJieKkqRj+U0hNCSrGt04P/K10PmfWXhyZU8rantCtlQNVCzE
RNNVv9YbWwLL0//EX080FvJ1iTKr+dFvNXfIdIq+yxD0HxwHVlx2uygM1Txv25G6
b98SFjRwSS9tr2u7R+XkvNZXu2rHjgUa7/F9O30UMsAJnDRkZNVQOGjRECsXXTgd
OysRYhY1kuApi3d+ChLev3nsu5YrjCuZ7Nfa1aBQRuiS1xlSQ8lepZ9zlzMS+be2
R265SIS1lYcfwCjZbfCKfFsWl+5Ijv+BAhLntVWK9TbQIq+EpCJGqI/gxsxNlgom
Nykze69dH96JeIsHKENRn716/Tv1LWf8TZWpA0lDcilt5JTsVrzYe+meX/3dL2lk
dxH9WtUaR7NerOov20IJ0gYvtVvAHrZ9vPdp/oFYBkSyH8LzScmNm4AEwgf18rBu
PW2Ua3IFc2qn2Xz7hRK702oJ4NbIdobmjBWQm53BMCMfB+XepmoNAMSTrf3S2H+D
j9aQvtO6JRrujTBp19HeXO07cEJUP+umqTp0os/9gp21a/VGXnFrzdQ+x/S087JI
OSk5/Agh+wULZMhZT5HI7nPx1ym0mkf932/kVpSPH5RZLTibGOUXzlifncIY0hYx
9dfJKFNgsP1RnWDI5KTTQ2EBrK8WO0rUprk3cfju8Os7YOYmX6qm6t9HbWmauXxK
26+hG6VO/KsQCtPC6xJaOv7zFI7vbvzjK03fZnYlCrc9uEIPb/2ZmQIsrliwqQ4Q
sJC4IT59hVs+SERJ6GOAxS9AUB+PoIhUrKNeodI+6NsZJKFn1AVawjTC8vRozpMP
RHt2WPtP30oclUL/oIk2rEN2QmFk9Kct3O+ge2xvFkSmaM38b6kRhJMvnxrldaB7
kd2l0VsXE1vxnM/RbviMhktjwt6m2KQXlhBY5DX2pEc9pilkVroNm437U+DsVdIp
QP4T6smm2RW/FgpYculndiue9/FIvlCJgnadP9aVhE3LZDoIqV5VOwVLVn61BTUY
W1mNX2LKQU9hKwtOWrCu5F6+TnnMFgMQvAyxJIWLtZoiumKCC9vw3eqvb635W2kX
kEFjmPaJLP8AAZdeWrpktYlIIhNqU1SQEohWz1n52Hd7qHNdAGLYl+fl9FQZLqsb
AmrqEhwsf3Ge+iPUpcNFII0f5b2GwKgooC4X8a9aqdnsn+v1OdThapRH/Q5WTC/3
qyCyarLnWzdFDM0RTEWGqitmBrJEDByDCe3tllp1lDvj/L0AoZ145DoDczcGhmyq
XI3V2OucOJt72pjgsBPTfgt2amJCO00fRNFB96szYikj3KkXyZsKnc/5xK8y09NC
YGwBwbPNFR+ZEz2C+lRaFCA0M+M7juae+zQ7Bde8Yuynx0BnKU5/A0S+y87XClE1
zvKysqqZ5qZXvwpLBsPQznAYlg20S326mHpE6lhdgW0m0FIbd8kG1n56sQcteOvy
jJIBhChGEulo0ZTQON5wIcKkRd/kN0jxUVMPRjrP0mhS2PVbJLPEDnBwmnkYKH/r
IKiVBAwbt+qnoKmVR/HKBEoCXCv4N4A+eMd62B/WDyzBYCjYjd0vv+X+9jADyJVV
0vtAdvG25qduwSf4xn3BWGU/x/aEO/KsfPjxnyqERYcUBGVBwBfH0Kw2DkQJVgK+
Nn2wToYdKJ1XV8u8G973//tJxODIIs+6gpORHVZFjhF5E9U+IYH2iPW1V9ELzLrh
BP4rC4dKWHP6woI+Q0AoO4+1gEBdKFmZ3IYVbgjjevq5P/UvTIAG5EvgVF7mHRHi
Y90fdFLcoB/13S6p73OIwDz9l82CnAeYT/GpfvqYnzD99Md2QLkEYJ66Wh1wZOIY
z2BIpFOs4Dv3Ce8EzGAj9k3G85b0gs/Q1Dvyx5jEHljfEeQZqiZEz90SoBT3S1H8
fVCjwZFv25luklZbYU8Xiug8Z8/9eEjpFKdvoa+HZBRjXFJh6gkuyBrV3EVjbrak
LZ6BA4z1XWDPCIq1TeY2elgXv0tHJXH6IsFbERNXqliPWQaLdDD0E3fww6FGuGW4
FPIMX14N8Bho/41ScbFgh9IO6XV0JmQLZPcp+x3C7gUAvDp/tRtwaEIsk+0tuO2Z
T/L7/4wsG/DPI0Vwz3LTsxNaL+YTEwYJS9h61vRW0VuZaEDRU4nf+HOFmHZA73uI
NYSWu66yN7kzsRGHVZbbA9tegAfz4soqgcLdgni407FEEQEe0iceGtTBVm5g7149
gFae7jUtDIzsTvIkeFujSoirq8itgoe+O3xVI5NTrWc5lAxQCIu4x1hA5/lQ9ool
1oXprfTciHS9WDJWbz3xv96E5+vyAHADKyIZKn7j+VAU7JkhEBWamVLKy1YH/UNR
EtqBsphpXeak5m5N2aS9xXOEKAlO3elg0eLAiqffI1rdiCDeBY1J58P+L8qjnLeT
ZIiPwalBpHHkXuIwkQV3yBEHBKifdHczwC8j8fl8eK9ilFbW+GR6VR+o5c9CRKQR
Mj7p2763ZMNiMYQK2ZbqL+LDkVaiC36ksZ4dznbyxgQB1A8IG/8iEA0W518tx8VP
QcovCG7xFS+zJC8iqtaSEAFEs6kI1pw8vsQQ3y2mUIrDV8UH4Ng1E79u3B0HAFKn
UxjnmIkXfbGNGchcIKwL7135IM1P1pn2QJLewk1Bnu3EAWTgUZjtVVl/uO3wvMFX
kp3vYO/KW+kx1v17XRnLKqGwYWhjN0FUC+D8K6L8OMqCYrmvhUnnq60jCEJS9uFL
2nxFl5LkWlXFXYzCakegXOPBOP9r4K0BuaqLnjA9WaL5GRqaGs+roAjBrtSRbnj0
x/smuM+lYYwrWr9TaFPvGw0zkdc6J/GKrrdI8Z3b8lrWwW5MOZhxYo64wVoHyvYu
B2prbnwlasHndSk8MZb+JJ0/FMm6wggetO7AVOAJHss1L9vNpHS9FaEmh7jBsJpL
Za9w0ADOZtYJOsaGCZgDaBvypbd1P9He5+1QT7QB5UEpb9S2BaH9BdZt9XtBfAYF
dr2P4z3d5eHbTyWOsVqs22HXKMXqc7dcYzyjDxV1BJHuH4oImttLQ5j+kdqXg+OK
H10q6NmEfCv/5OXWG0k2bg/vknRWtSOZ1MXC0p5BdRljHvKvIM6SDGWXmr19MHFe
CQwXBsXk+ad//BtLhvjzNHMJPuz1tMLM8JJOFAFwgR84cKr9jIrGAmw17YBFW4BF
ea3Z3zgI1rrXkqc9g6TO1tAX1qjvb1Y4k0CsDeFJZdIvlxQADiFYemLc/5kTmiNb
mKoFjETZ0xAdnn+Fy0XcFeRs97ri+4SeJyUuJFVpFSLxLfupk6opnz66kxPgv9Qo
wW/2mIOk4eVHGHcgOZNf/BhM+JQOe2Drz04bVIqD9zfqXQoM0CW6okrF+zj+rf1K
++pVLVOHH+35DAn4qwplNF50pbbwZhXGdIsLZflCQayH634WOQcsRkVKxxBrNKg9
KVKwnbHmulAp++Nj7yb4at6kaN1mpQwdC/HXVWZdWLgKmFE1qI5Er+n/5BI1oVi0
KBQ8v9UafYVyzZde/uNovbj5n4ClEaVIJvhRYk9u13Lkcfuo/g8GbcUez9sVx0y/
HaAosdk6Q4xPqWPDex1GxAac+DZXRQpui05kF7k3qzPT6s0lt3eUiGdS7tCe8/mg
5RGg4t54ykEK3kh8U1IcOtET6hhL55X/KJSUOdHm02hNBl4xCzxY4aSJtvg5z6qK
5FhQO96D3eYbDwMdUN6895n/m1Z9guQPsmoTBj9pXsy5r+7jufUqmmKxR+ZrXxbj
JUkrPaW/5iZ/+oBm65Rl0pRqlG7wj+vxYdGTTmoQa31owVO/1YUbhHUB5LTMNc1f
ED5eSDqB3pJi6yqgCVI05BOPkKrAPmkXDIAzUPWRspfax1JIu5ztlKz+bWjIYGP0
6syLERAhQacJbjmU88mlwIQVQjNIfbQUoQnDni8KChFyXSvZId1aTzOWZftGzGyu
6scifVebW22EE7JcgrnCsSrJ02SLzGp8C5Km6YS30MuO3Fd7m6Aq1YmWK+56oGPB
H4JnGI3nysPmiVKMiiG8HiM044O9v7kiZf5AxfnmZ/y0I+vZXtNfHVPHYFgzTokI
BiQnMtsnal5gUtu51mOqeihO/fLS+nksEY0ZYj23y5vNP7aDS9Fm4giytXCvpWNq
u/2/pVmrOX7b2IxKm92f0xzBQQ8ftHYDAKIAWkXLumDdzym5YdKoCVYcn5GNwlYb
VDjjA0uFF9PXMhOmxHdN/JHIClIEHGgSWne+eT6pF7b9IqCjBDNB3mZp80Xt3ifF
Q8MX2DEO+45svNN6FhYZG0TGFojTN8lamDNkJR+6oMMzq9E/3qy6P5hIyV00F4lS
q2rQhVf58enz7nGd52mbaddhsFAH06q5KRg53IBULPSK7l957q6Dju5rQV08rabj
4UUdyDw5J33ZtqcfRPd7hz98NTfvv6bS8apwBL3bHXKISyn2X79LFvN1JcPB3uld
JQ5TmESmd3Re3X1RUJBHN+xrptNj5/nxb8ktRORBkACvJQ3tNJ8vjGOJv4vKgAMI
QOyaRXwbq5NVrT6srsS4xo29bC3HeJ9Pi8emUbv9vbW2bj9+pXZ6ikG8YUb1Rtz5
n6IAyMfHz+QSz8SDWjDMx2mXOEe9JaMDeWE73YJt7jVmVrdKm+Cx3fJ2G3UtvwTP
1oZzFsVsYatL9+aMTbLwlMpS0Y5bDBtTccTWCrSfgAGwL/fcHJnsoTCANNyqwfGx
a7ybvASGf+0t6WsO5j/SST+ifc27QZEKjBdISiG/I5mcOy87HUKGGXdRMspbXvnJ
yg1nqJ+tlLYLMICBamVg/EJ43NvN3Z1h4UXUWdb4JCx654sG9WWhOq53AA7DnfNH
09xH3+9WalC/ayW7V8cPChEgM21OPtJGoSyGyTVbsp4e0McGYgI6Kbamt4k7t9CU
mTYRYibT0azdJXN8IDZFfWN21HoJ0q5Hd3RBJNdEoCCa7StxwF9Vu0XM11fVn4b1
wl/pz7prvBnkV6IhL3rBgcyJp2UFqeJGy4M73Pn41WqB7+IzqJA85R9HjcHp1RPo
wIaNLoAsKlyI3FsgCzgyQNPzvNa+Gq5yEN0MMs96q7Y4QpfOFsLXF0Y1DV4wFRqM
ifYQ7dngrSrqb4bJUZ6sauq1ThRNNDTUocmqKS4plPdZz/J+QZbFziuWgfYcGkMq
2TWIUsSe/zKvzMcd3NPCCEoywWwi5tsvBJpFQW49pMI5pQuxxLlSSczTFFsAHADP
zpVgWmR1DDgqg2bjOmt8sWtKQo8y7hlGq2cZ2Y1KhUThr2Z7wKQy3B9mWZur4JeS
rNqlnaLjuAzeMFOEcj4KnWbg+O79HPTqMY1U1/zMauZwbSSxfapGbcB6v/Xr8bzv
vGgWc6lw5u26klBVBEipRp1XUSqRZmOnw8LdtNYh89yFcgjqbQxZMxybWjSEXHt7
xbcJsKlF3NbHBvi24tonvHDaOcKDtFjqDh+9UDCNOeW5zUcUcI04TvzwMDJ3af3w
QxRQZWqFl2pDzPHEZ4Tdl+yHl1exjX1uXE/qRixunEVxrwyNRIdT00lsiCgVGxLY
/aiyvmgPv6EqG3VDZTf+MTVqj8qCRTo+M2k9sOInfXaUy0ZbdGHCd2iizT/hdqyU
oLlJNdAzglhanEjPKG7psfLNr/R74zmPuRZqX30s53c78OE/Z5RcWNy/LtOssn//
Nnwhb6kbI0dMv2kHDlkvLiDAn7hoCHqlq9wLfcvlgMxCfNl19+rVENo9WSPRU21M
AOm9iromxgvp0doUJz+8HUYA0Kj7Daxp466o2C45rdS6WgjcCGMXH+a+4EiCXCyA
olFCuEPLSVAPzsDUQmu/7W8ZUBGsT0yMvNA41Vx3pId/d66G6tbekZEHlKj6zydV
w2WGdu6BbGH3+JH5TNQHrJSfECRaoZmR7BhRLbSH3Xm2tQc7gFhNXq+dNYX1KzIJ
Rwoq3OQRACqO7RaqyYGSd6A9djw1tSLA3kiS1VHbUYUSgmnO8PJFFYCDL2+YShc9
n0nl57CXHza5mBB0kl11IxdTxJoL/yvnUwHlEhrD4Jbi/AQj5893/kQw4ssM7jLv
pkckP15iCkrCW97tUNrfZi//ZrSJYACuN2gJ6bH1fC9V9QGPVwpcefKCDeuI2RgF
ZJN24OtjKgaYy9pFOZQfWRzde9qMy/CaQvZMTWlP6Efdekti6h4F0QGhov+yuNPm
LA61EeotQsi2Z30eovYXsxR8eg8Za1EJHQgnnrVr99wDTweRP9KcOZpWMN/PJ6iE
e0TDDKGLpTNHKIc0pqiNINEqyNH7gUGTon0zV/jaz6hX1LOkIZmb1WMXcPIw7V7u
wHp0SyBqGl6uJwT6DQ2fbrIOA7HxJBf3yHk/D4IcJ9pSSeiIg6Pwz0SkTcSe+LPM
yHDr/GCMV/+W+b9DbqZ+elayYi/O7iUap7vlAUy30+jU6wU2JfURmwnjyBoERM/W
ChHhNhcffaYykGqfO0oXTDg1Qufx+03XhBIbh6BXDaeFgbFQAqCFXAj0AjI1umWS
n4H49qFDRvQEi+rp8+ZwaZ/QVhyHUWNKxQWcVmxATnB+FaP0ZtM5+JUXLcqxDkuR
yKFr8b8w5OtU9/De/qHq/uI7ZCmES2TweWsmTbX0dACzlQL6L4P3Smh9thrbVbPE
6vf5zccQiaYm8T3queGZD4vCRtsOrT9GxPsTnfdwH5i5ZhKL4E2zuEVeun+NxUv3
jrV+o0PAA/TgP/X5XZiL45hmbBYOio3P8OvpY0fxVVYj4sVIMByYBD5G1OUNIRvR
L9vSZwiDYy9c6ChNXycsbjUaI9MXQbC73I6AbdqaqaVA74aEcyvomeeml5D35KiZ
JF9j4PqsJ85fLWOSS8h7cdd+FIsg+eNzg6M7xDSdeyLLjpBG81j2O+eV3ZhrcIW9
7gHoNe1N3WJtsdPwUX4sW0HtX8mCBdeTd4WYHkksKs5GDejEdDcSKnip+VeOQUSa
bRAiP+D2YCLLQnN0Qz3o1V7geRiW/UTCIyz9cQ+MzFCRjPitQhv7ojlf/bvAFFiE
G0wn06VUq0S7Mp0Fh7c56M/KzwHAwXxRgyOfq694NM1SHobyaaK20l887G+LdkNi
TJ5NNXuZ/YBy26RnBXupxD3K7zNba+avxrJeDzOT1/AkwHjMmPnk7ICWIcnz0Maw
H7SwlN7r/sPJUSm0kQbM3capwOF5BeduK5SOEO/xJk2wNRJ67YMzGIZisHh0yUXi
ngz+CCk3WYRSQu2F1P78mnqJH6jGuIRCX8wQzHT9/ngwjbR2ebUfQQlohIP7UTXK
CdoYrtdV/J/zwzKTMgx2MkaQWbJssT0lPww/B9uxaDd+3jWGr03Rvue0vrKowYZD
915G9fAHoEveL3Z7og6cp5Km77SSlERP6g/uNOcrKCpWm5elmlK/r9lVPO+G8p27
RTqMzCtZ8MAe6ke8BzD6jA0E+I0neIMD4VK+srK3DN6pA4pCV3d2xNg7zsDRSNKa
luR4daRxd69/U7ta9IPsXvPq9B/a4hfLJSSydyx9n3fDhwVeynCqUTi5SywiWwWG
Jh/OiTxU1cT4JpnfZcWCMouSyDJw8noNpuW5yM1ohu2zqu0dF/NQZbOQflK0YRRP
iPpTlzyRAYDi3ey8ErRH/20SGH4lb2c9a4fm77I2rH7RsYJN81CbYKWeZkbTTZFC
Sv4kIfZcGocG+poi3ynDBo0m4P/U3LShv7c3dXsbxZeBmp/95Zi9bjBAHUs9NTuM
lFWWvUVJAmeIFRv2f6HOmnWuEPNylucIkKXu1lji1brhBe1QtjBEtANEmR9ZanBB
5RG9Xi2vdcWTJDpVhOI1CBrifI7PTH7mFK4uIrvQvGl89vlyaAgefNSDG/Q8eFyz
GKEb57i3DyKFJZyJkjSSJyHCl1UyINajfWAX6n7bWDWorAz+/R79RTnAdw9H//mY
4OLRi0F3UXc3IXx3oKYbPfBfP3UB2Cglns+uXT8xr4YsLXXvTfRXWITWEYA1Ruc4
uc0/hNx9S9+NKVE6aRbJE1iiRrk/WQ+P/qOnfyaYKr14Fbj0oRyksI9smhBnsJYK
jJxpN9IDgHRbNzD9Qm3rVJEwTqoe2twXty4zHnNIjafMcfI+PCK8ZhKTaAhbIh7H
jPaNdxmhuvYBk3f+4WGHNI2YwxC2p/Hn+krPPrKjjauibGf8wju0HfYUcnGo+6Ob
w8PHAVDIROHLD+FJ+giDPgUH3in2Z2G3LvtWgVXSjdZI/Rid/J6alNOQviqOFAcv
R9bVtoJS/ekb+YPjn1Mf89RGr4L950ejKt+BmAnDkLjVcaWZSx616aUoQF1kpsov
pFeZNKXoLZ+cHV7vZHAHWhI3fdYlfmE6CmRmdAO0KNByh8b6YT5mhMGZ0FGDC8P1
/A0qSxX3PO/NQkQaW56PxmgBrbi9VZQoVIO+WkynVqcaxz4dcHCv0jOMUmgsj2/+
a/2bIE1/pj1FaR7+Hip5Sd/PdzK5t9DPO3OquPGRl/te2bnOHmkK00DTYPdX4yMu
VFeqSMnthsVT6eOvK7XsnF5b41x4p/V+iSFAYcaLKN4AB/Kq3H66+0JkNuE7hNNe
gQL65bwl7x4nN+t9WhCUptq5rK/gmeKrLDNHaPUx+jjy1A6VUQODpazfz777wy9P
YuxxH/Na+Fwtq7xTOgTLSmeS+E7JdWIa/eD/4tNqCdxsllgc2QB5KU9+RZwZp5br
TwnGZBuRle2F7FNa3xpjtfTPapXiAgM9B76IBmrNHLNNjHvyjToBeITyDaAjcOem
qmhsuc5MIsZM2VcZubHyqhHx726++aBnzwyJkXfzX/MiaeOGEeWqTWzpYgsaaVwH
5DO611tAZwPoXmZcFpzgb00J7sKZLPULhlP4tbmlwzGraA7MfWQqKSR7vW9RqJ3r
F1fvum6t4Xr9Zl+T7+sYOSTLksuzn1/s35KwG3AiVbdnS0f1LRETulsmmriUZRTx
sVu/kwQgDgAxbf1pTEgctRH5WCDFo7uZ3ASlAJEqGcOW33YxhU07YZL6LiHmB1TM
Hi/+9NU3/D1wyZiLTfL/vw3u8jTqwQbuHhwGI3ph8mBUgVDcbhNB5HUsnBn469pj
Dkvf3eUpQL4SOkraXjMo29b2ZEFgA1F0werqZ3vRVtIuU1+eywOXNC3GDnzKcvSh
9KiFkHbsfJIQllc3GXkxWEJFg2ZaShGQ5lq5AMOuc1pRWqu35ccJYztvauNYwA0X
zWMOZMLtQXgVF0SJQa/Gs41iE8+kTFcJncwQ7dtD+1vAVRaGQ3e6I0OBielW1gS0
zxQyWKNwiNCJkbFLjsQg4/dR0aQYw9nq3ilUN7MGvH2ltNiV0NBRJKMWexcZ0rtt
sJFyaufNtFBSDLb3BR2sIgIww+2Tn0bqU7P3csb4R3nhjaJ20Ts8HRgkaw3NOzCS
4OI6Os7FNF2kd6f6CfXLk2/QzsYP0Uo0M0Hn6BhnMOSSgMzfL9soLoYlAR7QzfpD
s1IqYr3RBInY/bHDGP4YUpPT+jyxyBKgGltEozQF9zgGwYIENQNffBKfGlWYjQRW
0KcUokRxt4EmEc/sPEm5JcLYMop264XI8o1GBc3IZJbkYSS7p9QjV2gvXJC364GZ
i9eXFKVnBh0JydXun+h0IVB1pZUddZgFPqIUIHlh/Da45imViDH1V+QjRe0wXaq8
GH1EGpEElK6lvLYNdjm1s9h+Ir2Xikco32TN19hxMG3d2h/JMivOMud6wJruwOPB
V7E2eU4BQLuwjwwR7kM55510FlY9QsmIWPGwC4IE4z35RxrpwgQkq1xdFId6oRbq
b6CFMqWuGn7Ij7QdJohoIMpSTNWYbLG0P4Kj1Y3w4MG8zcbfZ6PY3QN3yMj+WGrB
qotLqbmdnlY0guyc7wjF/txSZ4+czCrUjWExslx/LsfP4WOY80+ebyWZfjtlsmOC
+sMVubg7TWGKInLGuQhGhTzi3UsoRNDo5r1bPoDRHyClhcO+TJX9H1MSo/DMCRwa
18odi1vtJSyvhS8DN8Ht6IfRZ6h4OlU/VSbhw8kHNODELazl/aqMumaoWjqQfpF5
mNl6USzUDRdk5bZw9UrV0Q4s7haUS3lN6+6KfMBTsRMmlS9g27PoLbDy2XQSQq3f
8YaLuZDyXomoCoFUGNAgUTFdKx1U4ke6l4NvNixHzoVUZTZkDEsWMZin+K8jlpuj
EJ/o3fPdFOYkzOL1ANqjOsfbJEFeyq3/s2iYs67C//Xe8ewubkc7zIZk1bQ6Fow9
gFM5mbr1Nt1svBDPz9319XT9njGDITvZ5qqgWyufOIJb4an1clpQexiihkcU4wxW
tY61IMumNuxl79htq/hRwmkgZ3kzk9dIIkEK4dgYb+96d0jhmXRnr2T2F6DBwImb
5g0E7dSZVtArakPBcJjV2YktExWzdaRMd9w3A6NIMYmnUtF3rpQxe8/NnB6FtFRP
eOUzan25/wH9XaGRlBxaO01gReOAI+xZirvyosoFVSuEXjVoE/fFwT5yFqh9NuOg
ob49TVaXTL8NhdwxMy0UOiAAKoYVfsozshWnjFPsAV3ZMInEySUghimIsTaY+936
8ah8y314hICeF9LM3vmbGBoSk0SEckNAhniRHPsRDzvlpk70+d3ryZ+8N7ODSklx
qYChaXalx22ggIv1JykJfe458rUZvSaSDhgtQKwvxVVDcOiQCS+SLGQzkV+D2WkS
15uQ9+B+tKGLedbK+vJc5Dq7lOkeh6wbycGJBOWzGgvZF4/Iaa6/o88ZloPOEHPT
Qiuev8xk8IngxB2Ppdf3hIO4ViXvzq+CmhsqrEwzAW9y8sA+I6FZH6LwhO65z8fR
GNuLtWsHiBfL2n6I4xN88F8zX6GX3JKIOZc/thV7cHcgOyu+2GhO4s6lUzmz7THs
St5qehE347WoAYn+JvgHkO//DLvbzImGXUO9KgeKPGc6XPkQ/M9iSZ56o3Ymtl7U
O9DzKvKWU6IPDm9HayQ/sOffJ+RaWWUujvcrb4x5w70vetb55Sh3YiFCf28YTzNZ
E1jI8+vQuSPoaGzrOBiXdHWvdcGnOElr+bwYCgXPwhTJ1QBwRUsb29cxtwbWH6Sx
XOuUm4dMdpzVMLXsxcmAJ9laYfQmEZlZ32bOnYidHW07a2isXmqPUXmNfRp82JC7
eqt5kQy5ubJIQBSlNOKZniygDzJ868TVEoIFaJoFWf4XlW8razz1IQSrQOkCUVQo
VLXT6VKfLfNIOxq/KsmzkdDQKA83cYB5OyPItluYA/rP2w9M7pEIx3K+1+7V+aUl
u2L/WRyuykBV/bl09tl4yRdNrgBTMfKhs9PwdvHkkPui6qwrFQ5Rj/o6tDgQXvXA
Zz6p43xEFlnWQlJc7V8ag8syFp1qHCKxnfIOC3awCocFXr6DMtZuZOZSR8ZD9uGM
8eZeTRZC9S7ggDIYEH98y18tVhR7fsA7YgZ8WcQhOUe4Zv8tLlF1LwAL/GACxPaB
yF6N8/rUJhb19uYTpc72RwBk5gcH48F6ev+YnHjTc3YtaZ5/e9l/X1quD8gJj0FA
XvoW39SPlSTzOJDuli2mKXpV4VWYlkuR54LM5F+vhez+v+E5n4XZadbvbscYjcin
lq12B+9yS5af465lR6ZbEPZdIfnJwBeGRERgErwLhBsU6fWqqYiEcjmyNRvlDytd
+bZC3kbwwS53tlkg5A+OWceax6MCf9SPTnOp4BESgHJb4NgkfROOV5FaNLF+0FLj
5xEjWwelCgsl4V2tXBTWSEJYVB7xaPq2ow0O58HZdjiHtTaKJRQLxc3cKZsck4jZ
dhuYb2naJHcSqJVAt2svl95XwTwgxPeIeYEyH+/xCqut7pQvuU8yWCqmU4x8nN19
4MvGXsYy4F0cmAUtxSncdE4yn9GZmjPy7Uc6rYY4iZsDhYf2UX9OM1zxvZDVLely
DA73I3zulQj3cVgXUEQXr33NHUL7l/bX+e6y7t4g4enCrJKUe/5Kky9EWt4IEhCG
fkqPu6wplwhEEi0Qx6EHd8ZZBi7TNgotPEEcO1mhaYUkMD0YUcHQOlVuUWeMUx3R
qg4GjUECg2gh78iepxEMLY3qw/xNwy9oZrxkPplASxvHsdb9P0mOruJMEfiDwx/1
aG232PeYBAt/FRDP6+EyU/HrkRU10f8DktGwcE7qO/YTf91paw5obGDsW0nDAlCO
RfADaIiv3+BBYh5TJb/uPbJFY1D1Woyr0U9vNva2SD9eDDbImR2t3/4gvcCHWaaP
FHmoZvh1JFG4E8uZID3yI6WOdKB7ptOfDC/UZg2DowmLDGHGaItqHtXd47Z5SfW1
MfQceiuEWZqN5iPsJybTOFJJ0LzX98qAg8VQcP2OTVdlWcd3kPu9ACplLMyZ8jVp
xVHJ61P5rN9Ync/t/0m9ixp2AyLi1IcBFjvCWZ4Q0Rd9dlNpzkhyOhXQAMnTwV9h
H9wQrHWq7WdhlJu6kQmZl3MB+21bqy1e6S0gt8c5D3AbpkstIsUDord9w7wRHwNi
spQQrCKe+CMb+fmunrX7FpPNArmn3F+LYoXKYvtj7RbxUTRRAjf+nf5QGLowhcvP
bz29OREGxVQ20NJmzsq3D2B546+4dsE0NgWPV+qjA60wIFGtf2mWUmiR+3thxMWh
IvCgWY1O8VUG4woZd4l/X/aVBXYdOTjI3JAubRSzkAvldmWE4BoM+U86L9VLbgbx
xzsyV+UKNEeRz01SAN4CwH/UCT31l/TFKbFFEs0K8GoyX0pdLuy4qxf7OMGNnw8u
BMUhZb79lBtnojtTy4zt7x9STEVvygqRPPv2hTuMe/p8aItElxrW9p9E1DVg3syt
KUCerLpgVLg52aOA2QkVfKp3Jo88Y98Br8/v+PqWFSATrWnOSIc4IJQaXeZAcAZX
Hyi4l3NKVtVP8SY1m6KPQMeHl6aoY2Kzt+uubGNhMldQFuyiiD4H39fX7ZdpBN0j
Lw/xoVH0KOPyQAyOsBhRCa3srYbndGY29osYcPpo7xDCzaHye5HgeUhN3UUz6xgz
KpwI5g/R/8gsVVqarrhfy1ROnfYfLoW7buDdk+d2DECKY3GL2F079OiG6J5UkslF
WV/tqdbOPle7KU4psC9WhSo+yTJf8iuOuIzYdPQZHU4wlMz/oXFUvNJ/yiKkNhVL
w2zZY7JqmJX4uHWRlOd45eTina6DrqEm3U9Rin2nFl1GZJmKS+/QJo1FZIfSahmw
JeX1iz0Vy2b0wz/mlFvo80M/IYVPYR0+QDZmZXdVKzovbJaJKsPdxb8eiGc0ElhA
WF4wXdoHMw3DVgXtNLS4IdGTRiSkcIRZv3miv2kQQIYCH3RRYq17vo+8NMHx9ZeY
IB0pK27X7Ef7SH6QGY50nQwkCVt8ju/mcZU+8dkwm5/dWgLPywzIGCw2ilpD9ZVt
Rns+mXcynw0kG/WrqnF3Twa+Ua09nhmOWEBzXz+XCrfQIhhIxfvIAW67uZjL1ISd
oUe47FVTVWjaXtTJMVjoApQ9H9hCt9R0Kc8LE1hhDf06HrZm+JBG13WwWkb/K6DO
G10sYrjFoTkjyWqr5CNQg47xivPExT/mMMkTP+WwpZz5HT+GFiLxXFFkVfW9vwAl
d9amqdu6U9U/mDriOJ6HAxCEX5yyBcAO83TLnbiwheGU0yUNHDihf6aw//j5vbXU
8/9fQ6gkkGOOlft798dyKooskifpXvhe3x+TX5Kfb+ne4EPJo/nRsBk6DGWoMb27
ZCdSxLzlTkRV38G5MCbjOW2h2Rw16qi0zWLa9mFBLLF5U7dLGMogjKNWvhFNFPUr
a2tD+27L1/Cfb+k4gQJOBBHMSDEsXXxISm1M5Tz97ROYfJGTmUhdSKsI1MsaHR5d
O5KBJs1QsEqgGFRbhYCy+00vpSE/PhMtFi++l73/wsQV3I50HwIay9+HTtvc5YKi
+/uKahfw/v6DP/m0625XgbA8yii4JmAHJWUHKx6hMjv5P+rfv8H7eWPTBgAuxmwi
yX7x6LsCECGlv3s8yAORoWGa5pSWmteM9ZlOUfOGmOONKfvztxR1cSz1S/ZS0BxF
LjgZsPsg5g5SPqD3oR9qh+3SY2OajXM0Mgfj71JiBOWfAFZEaHK1E1Dm2sbhuo3G
kPZMbMCPC77VC2FFbdE3V0SHewHMaNd3mcJ3Qfo4FpvToL1PGKmuB3cptIACZWsT
46KSvABoVhR0jcXibd6z2p4zstAFSgC+++Yh/AuBca0ZzuKohtdoG4UgqU6qd1nw
yqahL44hUiDWuZuRe9LNp08A7DD4CTz8tOM7cu9+GroBIXtBRPBH/8bKtz34ug+y
S0LxjM8lFzgL4Bi6i6Oh/Iq91iRU9BvL9ACeI4pBkrnsIKufe70YxqHNm+fbN2c/
JVn86nAszUvIPX7PdezRhjxCEMLu4WKdyfJMVtnrxw06mg3cbwu8RfFvxvVfavPJ
anwhNlchEPGYtXi6Lu7oorU+btzThh1MlbWCrPUWs+MIuWHLilt8vwaRWjYJZMMN
d7al1W7GzGUbjFypFpPRH4Pa0c5SzSxtxpawoMdpiW0kZ9cT7xq1gnwffDJabzAG
yvZMlMbG4VjOJ5QTiYoXPIa3899lAIKaFqUWwHFb4A2BaKIJfRAPj5pJQQMjULsR
n6qIicjt0rkqnkHAaG+HmmXjEtl5mOHGJkLx11X3K7ppl1tF7Mu9SYruMYNhBUYV
OaGRxTf5MGIwUVqwHgu1LZq+VLgpDdEdG0FwW7yrCEiVOtQ1g7eIOeh+IarGTZvB
5iLCLtoAO/r60xb4UEG+MfQos9dpBfdw4uRGXXiluBl6DAY2yJb6RSCGEFMFwWuC
AQfyGCj8bneNkjZpnFoExdqC0GPxrkNJkiAi1yLYoQyUHtYzeoFSl4Toc4sZDdLy
Rx43Dm9hHxJe1xyqA9k9LHOetfv6ZvkB0nwqTEB6q6bqS5JL3GLhcg89SqcUMkJw
WhAQdLYK/VKYOAp2gmzbGDRKM4nk/bI+UZRH+aeG4IYVykA3/qXiFOzqqcRThC6C
9FuDB48AScVcwmUJd76EUQZWRLYcCgmDxEhQeuTNcPAGg83QBN9BqO/w+cGG95EO
MTtI4tpzb+zNCnx7W3qXnLsOdVysaaamxBt4lxCWdoRY6xK4V6T/1JmrGiD3g2aZ
WCfhHoIP/NkTf4qM7eB1yAiqWq4oABpbBOt0Ht6ZvKFoDoRWU5m/GaHrSBn0GEp0
/JDWv1rRH7H58BtZQNVvdN0Dd7IRqzMNi7fwtKd/g0XORD6pOpQ9o0fzOPsUBLla
w6l4vji5YJo8mqGd1MSMbvGWWLJZD3mT8ec/VZbOD74OQiW2qFs5LHSrGFwReJGv
/Pk2+4+vHJN6nRgoQ4EqHS+raY52dKgja/rFzaTfGMeo86a7c/q2MB2UUSBD1stj
oO1S+ZE7NZjxTECBbi8dMV28TeSMToigHJbn5zqUCKQuu8a/PIuN0CbElclxwX8T
GMIx1GQaEZfqj7g9zqAP90ZBGrsDw4vpf/LDbe3hnnqY1iK0GEISTK2AflV8tmjL
7ULgNKkPvJhLTzBsznXnKmJJ98FJbsSKYgiXX5BYDBOcIzjks6KDOfr0GHAK3Xmv
9n7v/j9kmGL4aDtOeWLtu9QKPMzmh/4NKIKS9KkoZe6AdCfrmmLdfINl2M+dEbk6
8Ive1acVbaG1a3DyA5Bc9QuVp2JUo8H2P02tKwBLBxE479EsySC5Iufym9bnq0hU
KvFDBhDmrZnoK0tau8UCYMvVc4luVTVRkfyS5SNdW1aQuETm0HAM6P8F2Qhk2/5h
7v52cEczGwHhz+Fc2qTv6d/lv6B1k8yApHY5FmHtA+MuoWoD8F765bgDdtCv5h3C
B3eu9L5yLdIMMJWPV8VzsQpSXpSMKK3UWIamqYQEWbc2t/ezNzbWg+OfTqT1Cnlc
GeQHKWTM//PRzpsAoTanTrymP4z+KlDLsNvD+Gz/wO2N/T8upaLLqcpVTyJHgCup
ET/HgBZUAtnrJW+UL4ThcSJSvdLoqnhopAw3nlLR8zn2Oh9jawLxsjCVyafEs4f3
N/z6l8vQfkUZmAT5OZEH/N0D+3ClIyl6R44Wl3J7iEUPdgChyFU/DtRgHsEaOJyW
B+jx5dLMx1R3DD7leeOIf7piedLhTrjkv0YQQxFDeWiEXnP9Ug84zLRPdIiRnZA2
RWdX/GDWKGX4jh1bv2UEJEBuvTw8lm9jw2akCtLsYJDbRYyzM9PewA5HBqsamI7n
CURp16XKNukGSp5Ue3Hmqh9TZJXMexQfKRiZ8vsYchk68cHms09p4HEHwsgamr8k
q+6Tzd1rPJi6Ebig9yfC1nrfQRmZWk8BnaYedj7nzk9zzqiWEcmiWDfUtqJXfX0c
lmyO9gjTnX9bpcG8ftHiCL3JXHXrS3J+qXdIc4Nc7lBHLoK6g/Wa56tYTgixIE0V
VdZkBg6csqe6CLrt3+pooNPS6ayjDxoumdom0gBlsNGUCmYh0TLb84F0Ra3Dn3Nk
Mh9S9FrQfoiAv8KB6UjpkIf8sl5D+ZDnBnPtWy3Iqw2qNgXY887uiE9rDsN1dpGW
GXnm0H+q0GswsWDeOvVDctsWd3X0fHvA5gQVbQyMTh559T5l8MOSRLMNDcJHb+qn
jXxB6mB1Hh20JVMfT0Tl6o3LDuqLETi057xX0i+F6DBwD1xIDl9MmylLS2R3KXoX
hDab5snheSH4onbdoCtardSFNHh7XgJE1QlNw2H25TAWfTBzgK79MGkedQxJZbsL
eC03F9A8JyywG+sFcsZhdlLKQPYAeSZwk0pdiRob+50d/sxdaKpMfGd8fVJVF2a6
Gm4ieGDJeMLm4LMZ+1gCTi2U+WBzTsQMUmaJBv3XjZ5ml3gpCGlZcK+s/T1dzhRr
vvgZLUeu8Tki9ISyxNBJMqsgOzlncFjkzHF8QSAIQWFCnUT1PHK+JSozYVrM5rhY
UwxexKMFDkloD4qFD66JuwpoGDb1KBPNlEbXTbUDcmfka5OAtG2Of2nbdN9+XS28
jDDlwbmVbxS4dNwPnpQDq0x7qmljUbsWY0v+9fG14rFZHQ16QtZrP5v4KKIggm05
WxyMdp5dIc+ESqEYUiPd8EXirNMR3+rt25uIOcgcGjeQW69vogDoQodo2I2CzT+B
bi+bGVkWpmcJfOqNQL/I1bVjN7TQsTF/3hpiutQGO1TyMLoOk913rX6rEjn0pdtr
rGqcrDlnz5DBWLvtPuA63nVaVTyfQMv82FFB6fKOpUPUVBrpOVzuHN43l8pAR6Sb
lNnQ0szzLR2eD6C0aRavSdCjEr7V2n4e8sEkQcXygtDuvRLGJ9TpwKzyDILvp07O
gpqojrPu+NFKETgWlLHbL3PtVl0thKl95oShusVQLQRUA1Y36CHDeNCHN2vcnR8k
MDajv7beG5SN4mzDGAT0tJ6WCzL/LM4iTV/I6/yaT4sElajDzxHbVJbfxSJl9cBr
KOAb+iOWZOcArWCXUPtxYa/KNXPx2cXSgZJgKOc8jwYZkWIawYyABGEyS3u8/D+F
gtYNjQ9jDG97BoeEOuxvfoTwpERWeCaVQvXDBv+GD8WJMtyqP5bLwdY5WOcdDqFm
e7usXmU87XfiDB2tZHZ4h7hDKqwS0XINRS/XHJxWk+MDEMKx3AGsERBPD/ue+Dsz
RPueYBIJb0sI0rpLNE0MUtCvwBRjsqDvSDzrwqhmdg0sW/AYQMQ/VFEI3XS27/iB
7znH/OxpxefH0LSyk3c/Q3zWmJB6JC8kQEUXrt5+MoJ76uGdParYV9NZZ3TT0bIp
xG3LXHgOygEk7D+xVcC8GzwIKdJ6U4ZNhuZx1eznxGN+CS4fyJaIb8LoTDrfSMOE
yfssR1i7w6j6aPkGTapeKOI+bw49A6uXOm0RTKkYeVNjcoL9az+0qw5q+j93sxi0
lCcSASEXGR2htiN66Xkr1OvRaDcKMZVU+++Qj2lMIncfYnhOV7nWUkhhSBKj1MO8
AwAN7lbugbu16LOLpVfhlOqgxXsaj+Elh3UbvxrmtBCjpeJRcGjSTkQotZUSbf0I
y4d7j+ZeDDO2U/8kUFqQznG0QdbHGHcXtLTNNaHpnmqLVS/4gCRlUlhX2mfjfUfC
RKDtM9dhjdVcbXZSzTkCNyFAYBdXn9T2Hxptyn4L9DYKnMH2H0x13Z0YhqLzdGDe
y1OObapbnhnPnCLEjCbIaCuKEp7gYUu+W/xq5UZeoAB2wJkdW8fUSwvTwQqBdUZV
g9yidfTFZXsm0emePp+52hOW3I733tfd1TU9kTEvyTf5k+Qf7fhNBLUl76zrCC0c
uN1XOCg6MjLPjj03VMEO1Ta+TIt6M20goJ8SL1z2tIoPlNXfQMuIS6JS0DmGjlTU
BGC4M9PyfaO7aeNCDOAgAy3gvIf4t1lCMlMqMrE7w7ZE2Q9fSGdir1hqIRQb2JVZ
VLYYjwlDgzRwnBHIabiETwdh4NUm/m1lNP+F95BlnX+VFTOeWa/4f4lQLt/Q5BVm
VGSWB57YCZoiAsM6tSE4S0GYMCJ7hagRCFXRMUIaRfDm+MbGV9ovoveoSFj/KN2v
OImuB+XznIGmnDXTvTpBtksUaN1o7kaeqvBYgsGu2H4TMm3T7s/sKqrgQ8q7IJ1i
vZeMriJAho2ekrX75koYxhkp5RUwDnmNDnydHAx8vnHaJ3QAqJKs4BRBtbiOnBG2
4yEoLiyz8HMeCygHQUzviUpeIwrUpZNi2vdTupXKNyveVgCRXmIJ1wtFPg01qyvu
uTpeinmwzOGiRYn66LOoiVfacXXk5lioYXuuh+TRZMfdP5ScCa8Jl8jaqCt8FJpE
puZL6dNlNRD9fnyqzGEhRoaX8Wp8CVsCNAqRBBrTT9RXnCA5DU6mG3nrIztEBjm0
4DE6qAF+fZEfaUSjCPX9nexkRzsoyftlceQHvaACyH+LH2FsWWof1ggzVtDOHs6E
pR9vVBSqjDTX/fH/4omGBO4Sr64ldZ/fMiJedry1QrgktyrM6/bbfTOicHDvCJZ9
fWlPxwGpQ+0WE/s1fUkCfOwYJog4Bm2xfCcDuUUf5WUmnp+6jBTphQfwo9p7LdFp
rhQ+JmlbJG0D/i20Q14B5lotaPN6SWVTH5JYTyTW4aHRiLLdmdAOvOGiAn1F+5ms
fFbf76TOoPznxq2Lc9iVI0LBfK00GOfcLGo5rvIiZ0gLCWhtnfIuixBEDrJeUmPi
x0g/pIAlXZB2RB9Ogi7kCcmj20PCreyFHRL5ok2y7M/JW7lL+SKsCZ4nMQURvwZ9
EP0RvHUuW91sq9uLpqCplXx4pFZX+zVBPD0Qzv/JUNHy0tD8ZDkCsrMXn+k3TfwT
OpiNLI3nBiNGsxJQbLHRB42kcPRM4rJHkk0ojYdTWjnya5XpXQ8BwLm2aGOBHwrc
aK3ckDt0GS9XENOg4PEISDcUs5lLyZhglYsgWEAXXosUnlQqq7Ij8hEp8Y8ey8Ms
CvFaNZtcIBlQSg4CtM75ryvjzt5GfzyioM6x9x6xAeufprEkLxe2XfKgM56oUbea
oh3lbTUAmR4KzFDjgtRnaAEJyIhYPNd202+4kIdOyoUZxSictikF5Gdawhd3/0iA
Il45NKNekxXka5IpqLS3IhBKoj+VUYVVHAaQuL1ZQXSZV32zHvrDxmRwIvM2GDcH
2GZb1jEZ4VIGN5jq5K/4erBgXDzc5qTvHYrLR+/x0zPyYum6elqlsJIE+yHyUO+y
YeWP4kEv+9yNmobDDsvfZljjKjiN9OYSm6LT/Yv3iPCPQXy9N2cYON9IsQ99LhGK
+C7aE9y/LpI9WgmaAW/5xI0e3icvM3SBZe549/5uxe/GFpmvLg+OGN+Gnt8LWS7Z
1RCg/l/rjX44Yf4rTo3KqMGR7i1aWFFR+j+gtJXbDvM9oyEOsBI0gndD5Ri2cxUw
1UcSuztRtFsyu67wdZtp5QVEdUJWweaX3tlfvr8e4AVzbWJoog1MTXaQg+RnRofs
XrZgC2EdWgVySxAy7KxMwuUvF5OnW6Bl+n8tz5Xj369ugdqywGUJrS4A8YqQ0Ue9
g2uY+kCvH8sJCczLoKS7JehNtWuKtYcEhWo/yYSgNJAeh5f5poYWGFN8iqynHaBP
JGi/8I8LeJZbgE0H4rr6YAUfx9yWA0udwBV2kQEN+zqoxUOmE1pxYAD/5s+oof1l
8zXyJ7pkXaLwg/uX0BvMnalgMJTBh16lYKXB+xxGVK9evQ6wIbRo7L7MgVtmLSvm
SCU2kEk05ZnRsSvBx1J8MQML7Y7Tj00iki/NfsylffVJykpMNokwVwAXv+7VVEhG
kWWshThc7K2WSukoEJtb5nARLcLpN1ObRdP5RTflZ8ZtygDskWnnZUXNqb1zkAWn
8w45/byntZm7dxssRQUf71zzYuHN9Kiaw2cBxUsJyyg8x/2m9ZivthTkfDVH1ALu
e0hAe5beInqwW7yKLfUV+REpZxXe9b56J0UgJAXVyfEpDbYyopO3YDZiyBDWOKdb
FLK6oyZaImvpZjWICy/GdQ30IHpO8l48eJjvWzgAbjBh7o7TKcWmippimxqBEbgn
6QEOwNN0u58sRvFrnQAJSZyokuff1/Kr5AxB/7Ona2R1BHMJaneF0r4fVSHlEC9X
2wIDG3tmMhUg8Q88lS5B5BAHqy7ZnhgNc4TEmJAlMluj4ArEx7i+raz236fTUUM5
xi93hIVneliKI0bxNR6Eshtl5+7YYC76ekXAeuYqM++YH3J6rTSa7kWxMxjUspqL
Xu4KerbnSY4nrpE0nRHBkJfmoBqZ+FDaMOQC0pe7IwcDAKu6HKmgPYXpLkAbY3qH
3SCJhc1cDzz5XtGLxKSBdX9TG8umDRI2IhSb4yAyx/34kgEXK1duqzpyBXKhk5y5
ZTUbunDBz7hnvGlflxe0FoE+UtGUOEDOb83B0Ua8oc80QsgE1/prbgTTlV0MlC+r
IpXzMQJHtwRWNYAiSGfZqTvHBk6tGYqZjv28Cygw/mxgf53kV4/ITefN5Mph52f+
Pr9jD1vypnCjg1ZZpHSr4/RzkoDybxmEWf4/s0t+ul5P00zFLiLrLJLtPkIj/ntZ
86Oddx2LjcIOsTDm/px1XdSYhgNOkjCXUtmLz+ex8e5S2WyNrbAgrfjchpA+85Q4
2SbT4twgl5nVwVxq192Fvm72W1HkKRTZuYnvdDzzD3duPBix5c7FKiT1XVW85Vva
MhkTZEcaTR5G2y6uq+MPrVvEP0kgQOJBXkL5kG3wCyWQayzBIV7jEyhgXJckZJk7
oDS3trsxJsD5KSGimmYk+CgIwT5s0fan2P9WkX0Rx0ygkRJ+aIzySk2zJDl9LEnF
oqYfbEHk8w9xKXPYvsci+R+uOF0fiqJFMaG/Aw6NT8RJowuxLkQ9AuZQQwo6unnZ
4zdIKSypl3fQXOQrJ/4nu8lC/p061EZCBQsfDm9NaBuRJMNMXTqigE9sXJF3yabc
j4vnZlVH/H8qS+GblnkiGe1G8gHVbASEVOv00Z06pnriDN5t0KObLFygWncREvJN
vd/IkAPIewzQ3i2UjPNq47AlHG6491MkDAiJWsSPjVi2vGN3p8MgIAJyF/7hQA32
tK8oX8lO8USh0eLS+EPZrMgQl4GkN+gF6d/h7nD5BQTqJl9cwMNhQeBrexaAXKE0
NAEGK1zc4EsW51FQ1PfxNA2Ll6vB8S4hlZTSSX4Anec1+F5R635Pzxfosvu/+DGh
PpBtwzc7YGAjHEEu1Hehf5Lo3yDOcN9nBP7/c5Kw6XInSYR70wTWIeBa8gqbm+hg
JnyPD8Dg0MTodlNdUUZPRGMk42YxppKHE0eoJkCxG2hlYJ2U8mB38Sxw99gD/ZcK
q2FUBIk/qzevBF4nm2LctMMJcqjeANqVc6HdPV/N/ABdvcxgNijrXMMeH+AP0xSY
hqG4AAeIUekyVvZ4pqUSIIQ/rY2xIL5SbIfEKHuZdJOlXgREIFMVcBg5LIMalOCI
ZMXG0TmSgZaHF/af2HvV86PUxmlWZhAGU5eVYFL3kFrrEgQZwXHBUuGOeQR7O7Xd
TcMwvM/Fo97ocBx2vZ7mQTZMThaFmd6QXUkj9RnlHcqZ4LvHld509FNgS4pYMLme
RcXSTXfwVU6j8ei7LkleU8u/SrYBfzGT62VxeVLBpT14rpxnunT43B1S8ZRdBT/M
m/ZsBIXygU7RN7fWsELCvq7V2M8r1Z1uqJyOI9MM+krIYgjeFHDi9sY1vZnV+Qq3
33dEt+jIcoudIB+RmW8PaZJ2SG6EyxWZczBVJs+cUMX7xhhVGl3Hg6bczf9sgiVX
548l40l8KsmbB6dlNmg7lHNLl6xwRe9IUTCq6M21bROX0iwP/gcESHMNv52BczK9
o1HSEqAkbXib5vLsEuJwFCgM0EzChTmemxPQ3VeWRTn+YUmorKD3+FXDZT2LZbCj
AqfWXM/sQbHCXXluDCZdqrKi+R6fynD1FJNeQH392tAqaIjJqZPSJUGRe3i2y9K8
kT4TVfybN1czygUT3Jn3JcltGftQgP/cHLYP+DB+NVvnfcPjwHSi/+WEDIy80Pyj
CQbM89r49K0LMe+oN1Dx73k57Owrt5FzFq21g+x+yXPWVSB2qWLf1+sAKIRsb6/G
X/RAV6jZJmBoKXUisTNkmyZO9Kv5FjgoppotkG+4kPexaZgXl8KRIWEVRRXju4bS
uM3imXF7WNAsT9lvc3XJVucyiJn5LIj8JztiQVgbrNnjvMMI2RcpdAzt9ksKSuzg
Wez6D027XrAXgFbKt8aINyn1A/5zWaW3U0LkfLPNJLTUEuVw0zyoW9eDswfnau8c
CIG5FmiAFqtD6aRdcrWzdGdkd8RhmHU+6bO/QaqrGTils3Kws5c5qMdUik8edED/
ptX3Y+aTY4VJu6i8LC8OyZGjcHEyyzQbBwnysCRcBcxsVq219ILW/vHQd6UXY5WO
oY7nOzm8k72eD5siQjvQr5G4O8oxYtEumE6gfBEC+vNYmWYsbr6KIuIzN5hjHxHb
Vbo8xfMVCBKI6Q18ct9IckMmJ0+J9V5lgRb/NW2+fcT8qprJBEkL2+zWbTUesB3Z
G/IkawnQWmbDlIU6W3dvRJCqBBIHpbwlW0nDKn64zDffCBxEdxs+12fre19OYIGm
OnvlfOHke8f20dqpU3HiGVlvcpJ+t6eg/D0uprUTb/OYmmoWhmHIUwKZjDSMCB91
MIYgrEsUvrcMqUcOctD1lU3q/l1Isd5cOtBaJlUmt3srOuNtjhtIb07UvJLnDKlP
SpMmF6FhWIkjUzOP+sG3YNslOuq7kL2rbkw9Pm94fXkKoe530Ex+4Xyt20VE9oGT
SBKES+aIIBkZbTBdpz6R9T039UJqV0hQSdWGRM6eM8GkTtRze0e7r4OGYhmCtf1l
1EgNHFEDrE4G9qsOUpABUl2Wi8by+0Zq5nxE3RsTcdNYu3iKWH37P77XsDuQkPBB
q04xwSVAeo9bPNJReHX7z7eNgl06/hly5R5ALuDOVP4NFt/sjibPy523e51DnG/B
4I1pBrBZPPIYt0DIqApbfBbj7qpV7OifGZOuuxfV+3LyzGJ8zeHwiYPDij34PyIW
TH1F0YwfCR3FV7inIt4K1iDm0QepoVpIs7Ks83EvMf1Ga967wzaXBEP44lHwPkWz
6+2YXHzRjey5+SCleAAFGbx1L2Z9nu9CCEtIZKi+hA5u09jS4lXwwG6imvKinRu+
v/EHHwwTiKBrTXAriX58XFwjXttwJs/vIFudQc6MQ/NjSd9mgkFqOkM6t9qYUwD/
74NcxEkD2rliZ2Hi0DjGMw/VAoXb6zpzklC8FGKNtAw/s6WkSgegiPmgdHwA9VnF
ED54N41YI9mURk/JOzbDf9i40XTfbR9VnEpRoFQmjuMVcJI2e0LbSnXKhamOafTS
yJ3V7QZcbdnyfCcTEjCPEWmsNRpXVaERv/ygXqLAidLQvwIZTff4OmQ5tdK26AuP
71o11lyTnsHXyv0dAWOZVK4wHom9VDQw1GfHDhadQDiCOpSdZdST3/suaVLUufpx
XthExV32ROEnjhatbregmEc7q3X6JvauhPWU0pfDC/90dSvDuLmA8n81cnHDCWID
Nap4p9HZqVODdNh8zGJ4Svvho8mAoBYrVFbZIxk8TBdEl/FCHeRliCuXWeRUJsnR
dCrCfk1Z7XCjD6xObLrwNxxVc/koZo04tIXaC6/D/krWdWAq49T3YIISFK5h/l66
DJcH+INYCcWC+ami2N5QlsJO2fkAFd5RmQDNtDiP8B6DLd9nLdujPqaSkF4gYi16
DtiIsSlE9mgZXGQxRfMncP6g6hY+xGHTCbANYFp+RaY19q/pR3q6mMnEv5Y/xYy8
MbCVzzrmP507GcarN6lzR1bwRpysY259rsdVMBfs0tF9LKreU9aFiegfOYIdy57j
FanlWfvsHmKRsRztqtxndLqJoWj2WbtlW3qXtrwK81b6/43sJqfW2juJjiVVdaLp
pPevipVZXBzAs8H2aYwxEEL2LUUBImoVdJByDWdi/FwqNglOwIrCSGcM9JVMWj3s
nhwMe98iGnxQb86gmoZkMYqBGI47d/YD1A7OwArilHJ9XB8756LLKji9xiRuXGAw
EjZz6puOcbPCmNYA+a6rOxYTrnsB5S56enCAaVnoZm5ghlIyx24zBkfm3mTn42ND
HxOMX/gSX6IHNWcdXx/dp0A98ULTxg9RMXPdebi//u4bUjGpq/I00r2UNotSlaYE
WhsAzfk4WGJr6P+WM63CLGUvEXL+OMMFI+VIKcJn7xwHIvKUBXKY3S/FiEC6llKW
edcJix0Pez3X1MmdjEZZDHHWwfWRLcqwIZqhc2YQST+OvD+tCyYlewVwWaz9R2FI
tR0NZznsVvZyjB2eDygKm9czrFPUBX+tiBnovMQRpCanTXn13UH6R4lJ5kta6gQ5
zB1yH+a3vr+rjVFW6Ef+BnRtyMMh+KltYEZfIpPT7KpZmcv9Plv4EvRvv+4KuCS5
GSim5mnD4RRGBTlwG/h047PCElB+G/6OQazZTCQiqOUr7RU6nzLfpBHw6qfKMDv6
xJImY1Lf+hTU4vYuDpz3V5PKyDLRsBqULi6d/i9Y7bOFgeUiztAwyTmK2XGnR5mI
WT3L2f5K86zV2hNdV/VDLhMIXXfvVuISayeW3sU2pBcl7u31z+TVmitGvW477nVR
rzJZs+yuPIiKOOZDxhU3sskCX6AeXRc99TpaBjJGqoqYNE5akrBpTL1D28js2yPT
KCvzm70q3BtAeNZugC1OoG5NPMxuWRP1gBt+L9QTCbYQAw/QJBDfEju49ILqEZSa
Xv9oIyJqq2l4zrC2h1sHt8X+wX2ExJ5geGLAi7vtMDO8RFJ1jAcwk1AzomuNe0aM
ew5xi7KfcQF+f7CoWSaeTnPlt0N8f4HGhGnCvpZdPGKkQAgimPmMvktar/Ru3FyN
OzbNku8hH/xiw5ik/2Hq7pKzTQMbTmjCbFekoY50YooPMZF0RKYxFN3KNdYLRgkY
j/choy9/w1xBRwlIOnqqIbzUHEv7jjrOUFPsLcaZMZd7WGIec2MOizKEtQKMk0w5
/72sGQrDf2YVqbni8NbmpkmYTSmdAvkN/+efSQOovV4zFbrPThFyMrC1p+Xq2xkv
2WWMArT5aVl8PGgh6dRm5LhgK7ecM53ju40gBotNpugonTt4JV7GwnWZm8zvp8id
R6jVeqQMd7O92VoeHQHrWT35AoVPiCC1fTRxzUe5SCWawMbDA0yZEc3OhorwLGHn
x3MTKN8wdr8jROOiQPZa1OU2pPOszb9q6bbTadqc0gRYRik1cfWtTGFko5iQ+mVa
9HuPV2vdAt1M5wLzhdkcfTMxBCBpKhEGn+YJeL0TX4mAoORGfx8C8BllmguPu1d1
nFxpWBz3+p+UFo9Zwh6S9J8y3VmMGPdGvh5AkqshnFd+6Sjn1KSx59mGgckQzbtR
iGJN1xe+xP68q5ZqwSBFsm/2U+3Vh6qHARV64jCg4AncBS1X3pVvKVq4VU3yYD8u
VeiToz1BBQyYbKFgvmuQvyCt0jmwX2ba0FYV9deA1eVy0sWBldSelbp/QbndiPs1
SObqWrlg48gq7rTIQUrLls15gQLYWK42sE8BKefUxONVF8LKz61YUct7ZXOBuAmj
DIsgBfGF/4sJ1IvWcClptxgZS1QXG46P1HZYlktUOht7zqlHVBG8t2VbUADX6gF8
r4Z0M+2PjOPSvQgEeZ6JrDkOShG6rT672/9p78QdWgLQ5QGSqVlmtpL/609Z3BXS
Yv93qcdLtSKf+DKgNyCfOEM5EhSVNWEilUY8IH21uZlL2wNbIcuUPLLXRqKVSHqk
nkJ2FQo7XXK6H0wdUWnCUVyIvyznqCErY1cwczuAWwSJP0hKdVniiKauTbao9r+C
on5+FhGPOZV/I/QH59ySVcpUS4ZJpUNUzfNfCIXD04ljs7YEcOd44VdbalLIvt6L
GatGN5O+pIIW5fX14kFUyIbpU5xaHkODMcDW4f0T2EUvtGQ/YTha+TBkAkNjs5K4
+BQoiX3ueVfeW3mvsr9BGnil1ZzYB0bJDvgLyBeQ1y2m/1H/3gd/x6ETVNWklafT
M0f0FNuaA6TFiM56+u+p6YYKSAKi4o0xT4UFbla1JMk3clxCJlXK7gGvrt5Fuh/A
r7sBfbVP+TMe1wM11qRa5lkhUQ9uc4x+ejJg1BMwvB32KGEMVS87dOp49ZHV0+y3
+ErPFyjdmarI0ZnIPWxXs8tTapyrUHFamD0ScrvFzv7lBwO6Q0jh4o3fkAPjKwhu
C0skQwePfdSo76b2buUV4DYpvvf2sGZ5ZvxsG4pdaGH9FbNvDA8qs/MuNJgXfVNq
6KoPussGEoHt0AYubg3m5jJgbfThbAD00FtkqUdkf5z+aQsnegiFf2XR8XkvIVKK
j/ZK0yGNmhbQsKrLINoS1Q96BmDZLih9JcAF/M8T+dlJGEGFqC71Erbd1I58KgVi
JWYNURq/AGdf0lXO+dewjbLm1Y7hOTiNekvUqnXIWyA0JtcgOVdtG8Zxet5vZ/gR
9ZanPJg4IPjzuCT6JJqyKW68pi/oLR8e85g2u1ilnmM9qgnpqF2r2wGq1JoT1PmX
3bjxtYX0T+UWzQjECTB1tXZBaBaI4pkw3N4DndNmLNu2SPtdEXxXhw6QQqP/BgsE
5OrwmnXZT9BjMY4VOIoCX2yNCQKT23rjm0XwWXshN82Vb/AQbwuLvlDTuA9KMFZM
uvfVO0p26Fm7lFgyIFIZ+S/wi92G6F69H7rdLSf2AFXPvN+zbx5uPOAY/quRxGgn
5COwxvO69Yh1/uXkf89nHq7IfijSgj3sVKf9Vqu3etsxAK6o9chw9FBxsEXoL0O/
DsWvaOTbQV2/eYMVrDfSMJfCkWmSlPVJ4Uy5KArGtzU5JWRJ+rNtxWpdUqjYI7k8
GsNCJNj8HIygtTqWT2G43tJ7+jeQQFTHFZWC4BXVtqCbFYdxjyKcrFTQAtWd6nR7
6+6SgVFb7n7L3MAeM7zqsAXlxAWzf/RRhzucaaey0EPdg9MyeJG48x1n19S7eGH0
fzoDQ2Akre1Vlo9PHHB9dtaHqNGKoVZlbuaFMn2Qx5XwmXvyAry7lpJCcipaPpUI
koJnl3BSFuTarXorUTqvrGeygPN6zFV5gOzUV/hWOWUSe+Xz8rbrd+K3+3wgb3mz
0Yoqm5ZEXZwnUBN4dhGcDIs0oR9zwCZCplYB0P/nnGWHQ4MLMTK8R+9btmn0LA79
UXFwNZ6LUDvQRrBl5MwsGv1C4MHkOjc8iYYQCBU0Iolo0cLzP74gYK1qRIfGWPde
DhGP7j0sFJIEaGVR/cW20+RaoVNE8rD6YVzihMy/wOCf5xq1B5NJRYoAiArvTLLB
Dq303E9kOHy+GECJhMN10WBDHl0gxh1Mgyd4nvg+MULR7/9pRFyuhYJnhUPTPW0Y
iIA6cuveeLxyhfn+xzmgCYlSZabagvBubaYvVGWPk/MJeePjvDweijinMgilulJa
x0mfLiTtyP2ZR+pT1stSU86vUrrqcdvgyVc5slc69QJzLBIAzWnCJRsLEJ8RDLG1
O6Tmycoep0sUhe5PCiDePrDNWLJdsZut5Vr36OzPAOiVlsExCHcnIMw8MXUSRVMq
k+oj7lMBii91zw/XJjh5DvZCy5DBUNlYyljAdmCW900MP5R03GNtZMWye3Wq1Lii
NA/TGk1x2I12oi3oltZLeu8rJCjfMFYsmvIMnKVToV3rmERtwTkrKRZK+liAdeEd
NGVKpCP7xc1TP7z/rspO/4uZ3Jh8/UbYTf6NcEYds8DqBUCsO+shxy7J+OJJ+xPX
48VWNJ04ZUylGQlLIN9QkeOIdd2MXYPWH67NT5YryltKbO+SbLa2YSzvmlZs0Rbl
icqVZx1fe7SYbYetX8+kdDtym6zzkm+0W3u7v5SDMLyhmaDhSLGIR0QGMeLWJhKK
sFZw0ro2ZnXBTPcTGtGRB3K2svQHfx/Uh2mp0sgKVgwH8T92af3ctfE9Z/dBxyJk
el6ux3zxE1H+Vw2ywTuk1LDreXZBjZX6gGL4APlgISIi1OclE0wi5hROUdXv39Hk
kA4594cyXSHRMfj9qYL/eYLd79Ee9FxuHlb4amiEswRlelLnpi8AYA3kqX/Mu+GZ
29i9Vdv5eGlNtllA8nClhamvctlcjBdJGGrpt5adnTd2qeKV5chxWiq69jxidV1y
oLm/XlpZusALS7D5NderlYfrkoO86oie/Ba4+ARp1b7ppvZ2qZb9MS5hBOlUy/Ua
njwcxgfbEcPZT7IITKE80c6ZHxQwWHU8fykrrAeIfI/tAX3itQBu49kEiymKGKwQ
+jW9AKyXnDvkfQWNObNgNuc1XgyJtFt27dxjHXC/P2DrRyif0vnRLRC21Ow4Q88X
2yrqPQyvHTU3r1fbLEfGuW6czfV6qEw1bYqCBWk/zyC15NqI+mXeRki7qacdsMQ5
5QzYEUzXDAA4naFg7dznWdeXnb9lpvOM0Q+q2c89fOgcPvkH1d+Eg4P4EFzpOigA
bGH/yB/W3mYiaNBQPBoHMYqL6jomsPZNkVmfV0Pw/Dw8GGI59t6vYuC3aJS9zoSs
kBBu3JR5aLAgLs72VlY+ygvhtJbBdxzjmVUnpODxJ7PLPAilYRlN/pxf/Nt+Jj4c
mL2K8laJ57rn4Ujl3/BvhJwAVfH4572JArHttRfUgbvIK89tiX2cGFFR51NBqPdR
VL0QRvcdsCF/kn1Ee2bTZWHS+nN92hxYdOCTH8MilP+UQk9TRVbqHaJi1uHYkvey
snylTxE/1dnB6eJu9QLl8Hn5xPfv2fhUpZjhJ5e3J6f5iCz5VIgkItCRqMXmKYwz
mVr6F6AiTqWJjmtQGRyFemJjpXSMAS0Z6hn5/S4iOy1ov/d7Z0E/YT6h+yfBBOM9
E7Vd2dmTwgwXzDln1OTQGXXloheRCBIhsr+HeK4wk1gYhZ8uwtaXJkf2MEKfaS2P
BhPCeGFBObbYqbdQ0S3ljiJbCX3meVw2gzht5G8o59kpfGDLBuv7T/ZXGZMieFTi
hKhtKatXdCIBoixTdjOwiGgIP6RIgveoj/4b+bofBBD1XEhg+YiHSEptVsZuKcPD
F4sRav8hL00qDUynDufXNZ7uan2wvELSQAhB00toZYLfim9KnifWvB88qvPGw5Os
TrKVLohx13XPf+3o9ly/RDp2jbNR72o3ZNyoStUArNDtOk+XyL/rPztoCmAHbZT+
a1fmvUsrlotQ2+vLYlv/PeEyIdIaXJpjij/YyhAUdoURS1leMBQXvjG5mRfTdeq0
Kt1+cZIu4ArW5wriX9Xe9CxrRKxEZjBfsAY2xszPCLXiHHSN97JYI5inrAF8MDFS
3SqgIjzopnmkIQuSCOvM7+SenKpL2Eb5Lji8Sql8VVWKCSGgPKZFnQqOdlU5NJon
9gFWKyeUwXaqubSeZeuLD9DJ7S8khUpmj2Kgkl/rMgKNbCmPOrxsxN8FQhGCcivt
RYa+DrJqNpL82CYrmsZbPF2SjA5LEE2oRhSDDIA+Q6nHrOdP/7vmv6U9OSUn5iot
+1BLPknMaGKRCAPwGFbWTCxzsiOrTEuIjwPW/rTqC4Ymb1Mj8/S2pB3/6sD5Es30
49ePXU41DFwvG7lqy2nep+YzcC7B2uAaaqgNX1KUZM35Ql8vF9E35YYj7x8JfpgD
0eRrZP1RX1ok2nZm0Uv8Pzj9xohl85MoPJoZh6K36/jNtm9SLK2u9ov/HeZ8/rLQ
aBLYekQIW6x8Z6rOzHWIzUuIBwl5pVyCzNC9VMvY4Lm69LJX+sbbY2PRIbndFB3r
4oE+LkB5km7lghQbPsfbKYKgRQ1kUhzJ/YynDYtPNAtBDFLsat92UgZu4JanRbkn
HjtkHxr7E2tA789aRkpTR9zgbAv5URz5nUS1mOCt67W6f0uO5uxQQ2n/1e+D56rj
A4dOMEa1gO3qY9GDF+HFrk2l9YqE7DKcg9NJmcM+gnRsNLFmnYtJ8eIR2Kt1/WcU
z1hzGHMJ3KFPE3ReLXVt6jqq728e/tYqV+XO+vX+P6ICx+83oRxfWwa8w6UNcAQ6
7LlA3CR4usI2pPqNaHm4u4ss0C0gNHMBxUwcv4hL3OKyLm2ZonfJQMGETjv4Nq8P
1S+/O1ev8SCjRZAMIU28Ma/UFavbflFTOTIsks5o+ccT0gwKbd1Uk+fhFHUTEtlG
Nz+be5HvKcg0aRp1wZDBQklDLxlwTxDAblIELxg+H3avMseZABC3sZqdLXb78zsK
AJKbfK4cG6X9T9G1Y/yRYOlNzrtcY1dyY0/vvVwqDTbVcFbSV8dnaPzDo4VT8qNv
FRgxpZD6FwaXI+fJ3+HoPztNO7E4vQw1W0njQTDAI+5Rnxuo0SVHfnsN9zQo9rhe
ga6dh3rVrGOnr3/NWN5TeLIm5alWxWF+0ywS4XiHWpVv4YnQD8lowoHz5uwHG9Xt
uJ4S1KfDGRrONJG/v7m508ttG1YBmCv0DyNMhGZr1f9k6LbHEmRRWk40Rjj22MDU
v65IEEVLGQuORtzldo5yM0aQu7eOhkqrbkjiS1BXC2hKT8r7NxUKEGVqTK2zfKLe
8yyBKnPQ8xdm4RU/3gi2by65r4eHUjeVG0N8KHZG0g3nWWpaBzli4bVGbWrwd7xl
qOwumaT3k7xIu/Eziyxzyguz/A62qzeEgpLUGZ1BUxxPQqtIeqspdZEfqvm7CB5+
yTgZtZ47toQlv2rMVZVuBJn5KXol+iqO5iUgXhXkLhIUsmP/2WjtJhxN4L4q27IO
TuAhcfch6phOu1gvUd17UNiI2QC51O/ZIrr6Azm5ovuROscsXtTS+todGwAZQdxV
KKyQxyO5tglLXyo65QX8epVL3NQwsrJwukNgFPnmeGirFKn6jLKijodNhxEThNqg
B8vOMbGWucXnWkC6hq77V5zljmgsfCdng8Lvroe0Mwyjg6Qj4bbAAJUiV0/v2ZKA
TpvXbi32U9BJGIDb8FgWvodaCRfntJjHqDZN5ZrzmDyCQtGV1pjWB6WXGwo1ZCn/
eLs4jkGK0q74Ig1RVonLwaq+PxTi1Z2hDZDVJwOm29PQO+ItwJrk1322rM18QzOm
X+da/RFSORHX94bm8aTLYx4+WtVVPiaI5PTTlXuAQVAlZmRWhp6WjXadUpgftkOM
M3kAeMtvfRkmOM0zqFIkaJm9uuzkTHl4xe6gVolRHNfY0Q5EgVQStCiubJwcksLI
Vxsnge9hzf7g9FQn61LFN3MJ1EJOCdaJrBfsnpD0SpyqrYYkOAihQ4ukaIEROpRr
+T9B+Lgfofkyn/p3qoObhdbGQUVcCnZE2BvePyqFhREgCjNR5KK9Fw8Tzvc+t8J2
mgLwR+G9caI4IN4xq51ahzSnP1nqd+3prgayShwcJtDq6gGNcH/6OZXv7Ytr1u7H
A43YpqQmBUI4csBo8GzMytk2BLK4I7KmrYuQnLlkyM5ZsInAtWSYzKGHDQ1701Ge
jvJTsNXlFKEi7XBruOCSd8gCsOoXafKuV+t9it9GoPd9HYe0/BEpozulgvRB7a0G
9jgbbt2eIC8WQ9I0mLJbTin44/aDqiV+9QxLODeZeT55hjF4f8CWVaag6K6/sOMJ
oKrrUj7DNYOuNkQk/iBjhH8hk6Afd3MZNztkbmt8X8w92WS4Jw53vrDupbB2/FVB
UGejZKU7KhWOvaNjzFnVTx4fpKPjfdD76ClBAw9Sz+Z+aTNmEzG5Pn5YzVnWFt3f
M+6ydyzKkATLBbp0lRkmhg5k2S7jFGqXGdk/Iw7xi+ahFksZuhHuu/f9uB8jemm4
XSQ+0eAHd204FGic58PyXfuAZJ8557Dx03NtaVpX5qVyTCReOC+sc/CMtA1VP6mV
nuivUDBP8vaJMpI2LBycoc3rt/2c/vaubgKhRp4yu1eKRqCQPQRRwz+vhldaOJ/E
OXyHlpEPzayoI8IW53Xji4n93i2ZlLK49S5tRrMswfjO6UEw7xmdq9R2vArqnOdT
sZwii5a+0tce+tcklWiZww0YDq+Wot19UDfJvwqL4jUZxbptMDgTzZ7kVZhRpgTL
af3eFFWVai9gd7LXB4cVHgDPJCHguddUyPRQ1dHvEaUvrTQBwDVi2xAFb6b4yhLF
81KirrT8fszJ0fJcBOJipllRFCpO6my65XUb6VSCOUVCFv4m9/6e+ygZhMyYe9nT
Zrmheljouuhrliz/QMIuqAbgnYkQBY0+dUCI+Qf2idedC7I5ZSiVnoDepv8PEjbK
Up0ThVMHJYi19CsG/S+ZQ1U5nopbpsLsnCoqm/29Q3TJ+IveGka5BRFlP7WJMI1k
eFHUEyRyfzBt9WJjx8obRAxN2hAGeu8jVU16fRdO0EfFFczHITAbtowWPF4ys3I1
amP6jFl6nT5PxClpS4lWkgNaDFUNKBqG32RJlsar81Ri+t7T72p/WzCiOic2l9nj
jBMP3/0N6qS8RYZqh1LKaI2iSrjNYD1qDDmoeXa4w3HC4+u1MK1qLOJn9DL+AcBK
rVxAt7GhbU96IAxR3ixeZh9ldqKMz+5lg8289YaTdRr5iwIcByZDqfuspHVePtyj
YtT+a+87H0ZViOKktIp6fRsmPKQZEmWvjd2MF6Td7y2/DrRNbARE2S5Tzw9Os8Es
0pevXdTEEZ9hq4Nz9vrt0ZRVLnRdA/46gSuNaWuSwYZJBbfhufd2nBOh2zWZ/KrF
rYLoy9opNv/LVt4dczk96cH/NAxUJWJXDoiNs7KwM9m6OBGEOandrO5DYrDLIcrH
FuQ/Jp7RtfDbCxMvricdsNqRsMM6lvucoLz5EIhuwHiHGofBG0DiqnbiB1YNRtAb
bdE/ppPb3tsT5TA65Jo6JGztLeKqCitrnULk/1fCxbwBDJQyivD2or/cOmQN6jDO
0yXAMjefmI8NngilxcZt/FQmMD6bNNS+ThnDxXxjnXEuf79UXhNWUV8IzdsSreYr
rO54CyzI828sMdQiqV/unJ+ZrjlXXqRk5g0+8nhxdg4TZR4wxOJsc+6unz2tc5Sf
/I3kFyJJuLVy8GNh20PD7IKjda98kZt5JGlGfzn0+GxcEWTXXUaprrcQGwt0fwve
gx8Fi3k6+4uFLS+iwLDzWaqh/yMoPL4xb5kYOs8BC+XbR5KHwKBJLXVs2bx1KMpH
sWiRwYHpD6ExqsDEWErtAuBhXFmbY2MMYBm9GqIIZUNVBx91RUC6nlZnP+PSn2lf
M1gzNWSjwfD4FNZi+FM10jNgszTu2sXx+f3CL2A/crut+SNaEVf37WWJcBKTHCZc
HBVqcVx+kDpoSvpn0X1WggMTvGmIBCNxl9BlBc2RCJyxOCxF3e6Bf2we/vZvdM18
zhBFaKJ3n4K8cy1hHsdCTKgeXVxgiu2UsflRMKdrUDm4LOWIgFKeoOwm5YLm3o0o
2MoZuqL4aWuyMLyRYHGf+2T/Llq7PHd8wrfYltP/l7HkH8yuZNjtYkHzDbvovpuT
wjh6Mcv+ayWx4lGGitk17i4kQReIgNzXBXGGweGwPm9Wr1ATTE40WtKz+1jNnMR8
oXdT/VEC6xoNdURjIKP/8sAWDNu1Vj3P6XDwHDWOFT6F0xqk0iGVaX+AbbMIYeao
W7PfkebSTtMeOFaB2TzU5//I+SYOo8glANNaBpzoBAphUTvRt55a2+t0eBL/0yUd
VyRd2hl8qTqga+djy+Fmx3x7KClp3RJ679tn+O97rUqujsUVWWEDqQcMwcXZfNN+
mv9zhnWSmQN/46D8/ovAScnUZWgcXJtzD+fYah6A+lq5A4gGhaTDery2X/JSUFP3
oGVUsiTij+tbtaePQh9SMEpMX8b2Y5L+/tx1fjUPdSsWu/2YIxNPZE1jK/WnP4ho
DaombZl5AuzID3YuiEViujyT/E5ZwUIaNDEvPacWcWqHHcCRDCBJc6qa65th9a/w
VllWKpUOzoQeIaP1zI2avrBojG/VA320lfXc9sH2/uLcDqlPv7xAJ1hhH8VZ1IOz
mqA8bHyw/Lty4JJ4PHJomFYuxr3tVsB4s0fb+ePV6hY+kOaz7rn5qn9tTgjPfBvv
g08WLw28z1RAEjSU6D1vIBUyJ2UFehICQ2qdDBLZzvO9gIYh3t8tdVz5/37f+SFk
Ib81laZA0LRXg3vOOiA9npFFzYYGEWITEIAs0vh5ZkR3mJSwdStG1e0EvADBnKR/
HrjoINXrWNH4gTEklVd9lqfMHvkcv8vPQopoSqtpTMKon2axpJMN/dUmLFixLsid
hAh2ppWAfOrHsylVyL0Cd5526gLEEYLNuDPH8o/zfvckXeMwD/XPmczwqzxLmzOi
A7I1yIBp9tg9T87TeIT4CBS/Ng2lNWT2jzqDywp3K0BtMgG5xJaFsjdIgmUEUuyO
PStiDibafgoxEInPpriu5oLv8klk72wJGaO/fd+S27Zhe27df9nWIJrkILmgyt4Z
mSY1LKr09kFKGxrOF+7UYMk7Rgp37Y1qAYSgz0gqb9tS8TMoVSSewwj5xmOs7e6Z
WU14ZVtrq7z3TRbA5e7MqEa/TbIZU7YTdTQ2I0bUBr/OHMfjYXUz3ibrXdzudnmu
9KWppH3oYSfwX+7EtGiB5l/2ODK/b2o2rO2CU913l4yMdrFy5Bs9jBBBtLCuTo5A
vwZWhDv3g9z4yWLieWtbSWne13mxcIiCddBbA6WEpyMyerrDKWs5bZOJy/QlJQHD
qhTxKdG//FdduQC+U46VreV0Ra3go1qm0rrHfUrNDtB/b4aLCf80P+WLMbEKU21L
8w6/jWV6ipBfBjx9LmxwbUlOxrgm+8IIIHW1G+FxhhnrLQCgheoUfuCy9KdJZEBg
oHYsBmiBXLfWixYFKcsA/HjTKfGUt/x6G7c2vfrxgWFz+k05YhtVQJvGVH19ru6C
SDr1zkk0rgjgW2SLRKanhQuzXT+LPHa9Nds5xUX7B2yUamTyCKYSfGBS3BDfr+n5
hI+wVLObOA4kpUQi6A/GMYiDkvDTfA1yebzBFMK/mQMEAqR4++o496V+be+d6dpY
yp6oDt/L2tXgQspfNkzTGSs5OiOUKhKKeqtI6Vs/XR2HtATwZfG/KrvEeg0cHZfh
lCiXrDTFHqY/N+5kE6xIMlVrpNBRitmsbSZ+Hu4iCsyeVGj2n6LiSjxRhFVohuO0
ep3zZRZwzuUqNhk8kO0y1BVV4jKIPsTmdEf4gr8t+E8B03k/V0YpRYs5f1cj4bXH
q1+RGMbGilk9WSUMBox/w8Vb7zyG3TgKcbENCKbQf4GexncB3zpcWODY0sHOtkQe
kzmpOLwdXyHrVSlE2+1vf2lsj1eiQu7GV4WS9y+QYyf3SVvkrlkWFU/ICWuWi3gP
5Fmi6R/kPKJUBXGOACxnan+u7Qz5BrKsg1wjnyxO5kr4A1SPOmyKfIrX3Vhu45OD
RrhvTtwNg0jMDck1mPAjbZ/63BOJOJXOiTYDTNEgyMrUzwxTCZGUl7CaTvj4cf5+
gjR28A1i1w3VTXfj9kLz1JPpaWbdjkZbjYrAkIeKVf01PlYji2K/Bu1J4fHD+cJj
cTPa2BNkq5mKG0VuNCPm8XkEASZvNo8UlhHH5GZBNhrVspVVAyqsdPxYamIdkBt9
E785UBgslKaCC5Lwr750AyuKAbPO7cKx/dCy2dtxw25gEHaUSixTrUO5TWHIiRqN
3k08uP6LJCKFUqcy3gu8Sm5C9usmcf+dL9//22V9lViODMM6hfDmoW8GmG0Nax/U
xD4i3ayOjuskYoYSBOdHsDWSViME7aHjHyMvUNEIZktyUl/8eo2GQj74VHEk8C12
W/QNV4lEMJ6B0BHr7AYvY5qjPx2N3zU5l3yG5zu5nIWVk5oVbwHKyB32wAJ/U4yn
kJzaw12QTM9SLgVKQpJybu+GcpL50PISifiifW3oE1DiKzvEUdrnBeCvuoelbNpt
BVUAmgjXxj3CLnN2T4/vvsjGepZYOS02GlZC2m4NfeQ8mxnQjz7ZKfIsPgK3SfpA
z9MMIg379YCCootR4hbF/8K4kE8J4sMoANL1X2TS/6lawRI10ZGEmVfN8JAzUa2f
TWFA9IWsH7pZAGDMLHebo5JcVyaWGwUtC1gnady0BYbHKJMJlPYh8RZ+4m8kMakC
MNvzcUqiGea+pem+qXj1girhVq54gR2D0xW/E5kbxDSi/53RtQz4mRdX8fmSmLPn
H0sBlCQM4PtVb45SnEQunYQT7G43S1jsXtM3D7FhM8Yk8938C/A0OXkL0RHZBWXx
UmiuKru3Gok0m4FF4ZGUITz76TmmUYD73wi1xMVUV7/wep8VVTi2qNdj4QkrUdSK
hVG7UsRxPjR8FJ80kvCBzQWCnn4FsJ1FDtYwU2X39N/Ql71KhofNA3GCs4trORvV
0Cdj4HcK0w+meeArGFG/M1M24KwBxr+vzTObUi9G+zZLCdC3YfxegBLZmzOhceLR
fUgfqHXNAaKG/05pOVQYWDzmFVHQZ00/s21HXzd32bY4Rxvn2Dno/Z/cVSV4NlHE
vn7UOqU0b6C3kI4211wTSpLO4tFAoDc3Hq9JTRf8d0ptlYOmwCygXsfuyv45TRI2
7gpL3x/qs2SQ+XJ2CbAR3UUeMeAXBauz+MoLhot7pDrMNhmwvPHk1m9hX0MUZlrs
b+L298ikf1la5uabeMCKkLkcJMZZhEPW0ITb8mvvUpJbyq4ThowIYHQj37tFUx6F
5WaXGT8RMKKk+fYkwMOVPlBuYowGMuuE333t5Bf/FoXntYLkjTZ6WEGxoKE2jL0s
DEOmCfJ7r7K3aox8QqTg34paMuO4BxNbKVITdzhJZVrA6mF0MDYiJOjSmWsodMMY
YXcBgxEQBokUIEuQeMPTIaJU07hDYMnXTH+OH0APKAsA6WcvhFAus8YjiNVxFi5k
ZKHtLCLh9BpRl+2eoxPUSR5ApLuyFv4LUxIoIOFUbzgIT0hDf1eHnofyNKMSfJLI
/tQyGbPk9EvuEeMvMpy3OITvW2hoBnhr/hk4S+rgKbFXJMGm3P1GFZraXGWxI4wB
xm9TIY9uJnDuXgMvjvcIkRFmzy1DlxasEmm6tWEacoJEYhTUdiHeDLU2z9wHwKOW
nJcJnhqM7u+8eKt/kjEjatuua/vkOiFBKgANAMp6i1myc2N/9LwBWOyf/goQbLsN
n2idrT6P7G4yhRlldrVi9a5T1XkawBARvdjnTa4lKcUSp5NncTOzYBPT/OzUkzOC
n/w9uctmRoheNPNKfKKozcJTRcwmd29qNlARO85bRaFBuIX0WaSO2gfAU9hVQwxT
C7ORxJoYzuZUTg9AmVT0/DgFhhQVhOcHdSUSrsPJyEaim8kU1NeI4a1q9xoRS9gl
WsHgAXkbhb3xHO0rbipfg6bIGEtbwy5v477c/mv1u/39qA3Zz7raY1gOd7yTdysY
qaS8bHEADYQCRqa8Jd7mglhsBSHCyGLOdU/EEvjAOXauUQRb5faqSDkdGl8P35Nf
glWzuwzKdIfooMGV33du7mFsOvzG5u4uao63PJPc8jE+ZifpUAhh+3pt8hQop3Hz
AEALOzix0iN8Ro+d+PbmDxaF8N5Y5GYYd5guJoys9E0q6U9p+wV67avIeKmwQoGl
7t2mkHD8C1zWenvVfbyaruPSC661Rw6FiL89IZMLvdpC0DW3j9yRfwbPBXQg2aAT
8eXFnRGRW8a6c8Rg09lpdpH9augcQkoJY/ABD9lAnrEyRdxzyFxzG2mvSawE5UCK
AGeNS6frthb/4NrHPSt2MID+2SPt+//gUxMy+oU7jSipaN5cTO+Al6jwKQhSNJ9l
xTsRtMuwjL0so6MW2LXAGWInmPnga3G2rpz/d5Ubsg21edZPJKNUqKN8fuJLAAuP
/6rbmDGVYrs7OsOf3z9kp9VvmrpuK/mdKB7FbPSHpH8ypC4O4C9giw6IMoGp/8Tt
17jdCKZRufS38ap3gCedZyrh84Lfk9cJOqGzV7zbVDVtRi2ijFF+rLVw5BnuW3TN
WGC79nW2x6E1OEAn/TmgA0AvwB9Ksu8UQMrpeom2sXLHv7jrsl0oixOjJ6hbtfTN
jRBZs6Wa7rX09hOZcnjZqJNsO8jYGWs166B2txAQbdd5G4lbzJ9K52ENZA8FH86x
GZsZM5Zx04QIhT9m3y3FAn6bnDMxU17oEez84gZkERMRWhf5XHQovDRlZsF/WzdI
4KGmYPLgeh+CZiFyBFcZpRhzuU13ozAmkatS0248915fKmgf4Q9Qu3yHt2X2VuLg
DH7csdoTojqPWi187wekrEbzLWndq+tN6LNL+/Oo6TxdOyZQ9mbwfm5huRh+kk01
s8qddoZeSA6S7UWaox46fE2hKiREHdG3c2Mz2HDx9ab9vgQXTJ1yEpGjh6riRMZe
+n5Ju5da1Z4tjdm1MDx5jBUkABPFMdlm+WRSPvdpp24E6Z3Okh4Yt+N+gvKsXueV
kKv7rMaRfN5TK5NctPy+OS3h/dZ1h2KhPZdM+keoxVISP65GhoBpkkQArBCtwUP2
eYG5r9TE5y5YuBCbDcUp5H7kIWAHTh5IM49V4l7ncQhM536vNDXAA1nwjMusQHir
m0ZhMpJiPaO7jrPWQByE3BfVfPtDtMQWzuijksjmqR99BU1eB2VB6Xrp7u2ms4aH
7UA/mwdCZJjQRU58r4Hnq8YeuEJL8QXS/dfWs/Wk7n8z+0ZWvgJA2rzjfXf2Hbbe
YXQDoW/TxIngujcfiiRKxTxr/V6CQDCHCqNtj7UymM/9F88Iqr3zpy9FDF9FNaUE
6YUYAOYlFoCKbExXuPjca4+vPDj3GtAKzmZO5XeFhgJg1rBIzSXn/CJ3eQJXPfnI
FH3DaCHjNkb12GEKfTFSA49A7doxBQcpxPsM6o8jKCyi0eYx2sIcUflbSC/LjsW2
wcxYDf1uxo1JUZ8je2VN1ayy1VT23kDOd6zYv+4ifhgVrF53CH4rnTKoAE35PdFh
5V2ACcfLFNE3Zt5GGaJUxHQh7Ghb5CnqL63mLiOsz856w4zRvoKXgH3yL0WC8JR4
wNlsVdx3C/hJ4jvZqkW7MeuJpG3/qyW0MwK5lmZbB85Bpx4vzfHEFxqqoWTapGtT
yyyV0Z5RXMdxpKKECAQHgY0gxxgZ7/lkjV3111ZmvIEBY3AvynswWDKnxzsjaVWY
czN6uKOa/MRNPlJ1Y6xTMNJ4vkk3VTdf/uHuZUGAStFJjxrb5bceJ1atb+wqNY7/
yNnojXRrNw8nLb9I10gFbUwaMAIv4XzVujEzRAyrCaYa8U4kgh23Ev1QDMFw1han
P4zQArCnUSGc/l0Oj59DG9/TfWA4+mukDZB+q5elvj5XESB5bsiRfR9QgCj6VRxu
3lVV0YOFAdl8uTWHZio4ctMUHs4as/Z6VtV+rzvhZIOSSpbAdH9msUZaYsH14QHJ
hV09ryWrzO7RyMGRzkZ6vIdEYsGuSDudoISfl6tkzYE1jZAw29GjinJMtquYlpmT
3CQ6iC2mlXP6hWR8NJXf5ThAeldGnJbnY0ZlTWHd6N+tqPVtAUHmZcl/MbOSGuB7
bM8YAATpTLdguI0PlEm6WeOM5UKbMfE5gSdokcSHoWx/sI2VnGotsal+7y90xlI1
DsDiIwxGuWZcMsdaZ95pbzk2/m3VwXEbQOO0pk6N+K3/Gph8MLqXrBIukPnAp5oY
mmOIElvSbR9FOaMHLFp9xrNTw7lRny5X+f52zXZ99srgfCJXnzChHYL2m46hp5rD
I4HAc5mkQGg3GHjUgY26iFE5tDLJv4MAvVLL8gF5QCbUxudrjqyY4KB9UC3PM8TG
0feuAZjuE1GNEg/qSKAo1VxR343I1YfLgRCJz6qhIMxaInYL1stchL1+YfyDYqm+
UkycVWUK2WqUL2SAysDjraAX1eq2awNHTGppSLHtRYmUrX8HkXyJffY7o8tLMHFm
g0oyU+fmjse7DAvnxpSVgBohbN+Jp80FDYtIimPAp1dox0EFuohwF7f6I/dKDPEP
21tinbDw34s2ioTlZd6NpY2TUCM0cYX+5ZVRSxVXrbYtNo57uyQg7LsqSwiZrERN
jr6qoX5FL0eKHwsFmTkDUPyDA/bVvB0DAooKeLq+pAvAeCabFlZvDC0BCCHgWt1R
gg+MhjfMrXWh2jsAau1Kuc6xghV/b3dHv7OTsh8MFcLPGR8yqfeJQrID3SJg3QsT
ZP0uB1lLRCGThaEd5tH23iym2MErWvRJVP2vz46BwnpT7gjEO13Dt2mbUNuFjvak
5AFZBn81cHpcEyAegEaR9g5/TGRtZ1NO8naunz8pRyBbI/Hr//u0wtyGO7uP2Z2b
/KomDQE2fWkJnZ873PrZd62GdSDjVzeelGXcunUzT8+DVkocLZz5sTVWpLfb6gho
HMNHAWoJm3PCh7zKQazeolkaBdkITm6DqEl4DQcoZ7L1W3Wpfx0+SZ6c7FwkHjY3
Lz66Kq+b+39aRgaB/qlIvEL9pA59R8HfFxenGWcBsyVN/rbUnee5UPqntqxYbuKd
kmqyDvx/utuQxaVp5O1s9607F657Xeuw6kud0+ygudZM3gsvMUIN0bWCQFOn2ZUV
9aOikKrdYKnrIOQXTfLaEfh6j08egsPkTGvuAnALJUgNxR7Rd+ueF0CJfTGGQez3
ZWbOm5rSXhyFaPadHAO99Kt17AFnYSydRUooYG5fiZMw8Ac6gUx/t/LI/FgpBBCC
AN52Tcp70lJxWYaEiLpGs6Tx22XSUx3rHBIhJwQX4TcJOsAjbjuLwKrUGKpNdBuA
sb7OvpriF/zE+8c+9PtjSaCdqWxa8LxF3JArZ2v9wlaOrJ/aqkPiNG8Ye6kfhh2X
Bu/GgXSt4lSdopwSjaA+Wwe9IcnXaTmCrh2l91EtzNwYlnYal98ZKcrNUvuCOB/8
YUXMYuTQnmbQ0nfAaFmpQUNVnRQZ/9YxSlyu7jPFPbS9WiHxjbuvIeYVOOPdTnMW
Uiwz7g5naW1CeIQNkZiZ6LXRXkR65eq9XJezz94FHVCOdjBllhktvHWfimP7HaFc
lmW27iNQIkyNT6UXraJ4o8smRh5O2X0RyC2VonounK1itEqL6lOrFnAn/IN7Q6V+
FNbkGUlD1lYIOEUc5WE+9fi4yARLSkBC6RLdE84J4vYcIiXlw17ivGwIQEdRzlZT
h/WyYcHqpoLxSbCS9nkn0Mmp6944QzXoxj/cR6msY1oRqBXkDgFUbkXTG0XcyZQh
2q7AI9zzHGeXq0D+3QPn7AZvZ7tUby5AgxanS2YCfZg7jD4AS/UKevCcXWCzyaKP
+NLj/CFDr93v81m3JkrERxI5yqyYMFYTobtvuMRpHl+m8FNOVacF8If91+QE3Uzr
okB4lNKZQ2i0QWEDBUvrN0UtqH/Zt2FPsqpjYr0PQRX06xau/sNZqLS2LsqhGldZ
kdwOl6mWhkEgv8b4RfQRREnA3ID9BEFk1GFyfuOGBsWYSfv5nfcHckhdk1EEmSSo
kVr6buMRaA4X3xjRJ/mjBJeZ3mSSNgL5RGIpCjvR2+k26fgjubwLbQpcwC01A5bD
59R3b0aNlaXkI2D9PsaQZTRrS6MZJi3Yd7r0X0AKXKSnhDyKk83waIEw0p1sYI/I
/u2QjlZVdMHUbs40To7DAdSdHnXfuZTEvt6guiUkEr9eLCJ8aI4zQj75YPS2/ESH
aESXg2Gh5sv9J170elOD6vwccjxYoNjrj69uI/56qsBk+WQg7z2Hj9SLLg1HAhhi
WJD39TN3Q4E2rOX/GYWiZ6sfT8/pWUGXNTgT06yBHTepLEYjGqAlVntN5eFYHXJh
aGkg2h10j2d4wDxI36B2LZk9AXnZwMqUC8nqhW//qnSk/9gB6ut1C7EIh8SDd/8L
LcQZI/HflXNZWzkdJy19NdlYg8A8edYSCnpUDs6NawEeskpcCj4zvieEOQ9+/j+e
fpVc56bGns86JLjIia/nHxGmlcZq+Wu/XI2NFRpWTxKaAQ5fvq0JGDzLXd+PMAQL
2B6w2k+ACHKxsAxAmAjCc6pF46NF/FVyyjfgYJBKUwqN7HIAFooBpqPe5CSy8y1n
zXgdD9jtk9jWvHhM32M2cIfLCVNqCJT9JAYiKBZNjIiVZgFtV9fEFA1rLkM/9578
hgwguqtTnoZE9D2BHdPB5K/ynArNh+U5c52L0kA6zr6cQqKupTsjQ7Rwac7zQ8sZ
pBs2kpIE4kKRm6RFQj9p5ZJDxW34QSp00V00xoJbgddK7BnCn09qfgGmUX/M5GjX
ZeNQXXfhEfwx/ctiMcm+0Nd7pac9lbFeV12bIRmIX+rphlfj1gA2tR+0hP6emOlH
529ytxmx7/i/49ZX7nhOYeWYHMrrzZXK7815rMhct6nLLhzX+nAMaCy+/NYdwz+j
Fiw8Tm7S52AjUVXPMQBknswLEGdkB7QVZ5yS+P/81TYidRslQrF2tJK+xC2TBVhv
a8nPJEdaCXk66uj/xJ7ADlbb0rFbBV2Q7jQnUxj1cUa7r6hZoKWrRkbCfZ7uSJlM
wYaaI2tzYJHWXq0BBNRioL2Y7oH+kM4/O+h1G9jEid3ap/DiqJyhWjYmjGnCe1F5
hgVQqzz33IRV3TJLyDy6YRtAa9jtaybNS0rewVTQhkDEaR9LVPs2suHCXESF6g39
y26GXohmcvkUDy/D1/9Ml4g/m+LqD5dhZe8ADVU5VDJ1Z5pDH3+Z6OtjP2CGbZ3U
uLFOKDWO59U6qrMJII5ypFXaj9zFPzOZZrygQWNT15VvjYaRUh4OBXezJSBA+1Yk
hIFiXWijgONke9jZ8n6AZRSq0N0261bWJAYO8eHP89GFdXJe+Z5Hy0488K+5iHD3
q2RcT2xAJ0eoJCFdqqAdZOUJKVWrPgLBHypqIQnkI1vOC3wamuYN/AbPQNZbhOXP
lGFrF8E/yWOh5db7F01Oxzh4RqBan8K23wIPL1PWsnZ/bhQ3oNz3/Q6vpLMsUWmc
Twyvr93tGBj0JcEdol/cUF1ZD73ixxUADQDJLSdJBUtG5VxgjBZ4gLtW2lE1oLdH
o3ZWO8rm22BRBEsWRxpjw7hp4CRJh2N1q+jC7YCi47AqzW/5rWUTl9ItwLcpwbPk
1UvBEF5X8cZfNVqFiJk2ynE7kZ4jqJGoEA8t467vRAaQLNeJ0/Bw3G2xow1TPjlm
RgnZEyGGGZUBbKTA2f6HMHB+uzrOZqxTIEp0lgM3yW2HpzU24xZNbj0hX8dAPq6T
wlRAXAcgnwn0Lu/8oPMS5Qwqzu7qAHtj5UNvD2t18+nUaCUUA341d0Y042o6Dwq9
pgW/xaXl8sC6RIlCkqRU0MLrnpxCXP0uGCKCGxndJq2+eackPaYlfv+tu1XyFxPw
xZUzEgEDC7qECTro369s3NWs4327h4LlGQ/FsbnLWStDxieL8NqcOVDdzJlCgzO4
0QgoxvESuxNyDAIohnjMKHQPKMm8TjaDYVWTZPle022Q14CXcChIUbEkuzWxot64
pWF5a1NEFpo7KJPPlCme4ETx5OKOyz6JBSAPp1IClN4AM0+iQUoc6fhsYoKnB92D
+jxQJhzNary8ebIzyuepWGEjLcuNoCZxgSzc+VfFFtEZPQeQ6DnAteCscDXXwHGo
jJq9n3kgX4Jk/8A7gm8TqwtCulcwoII6+1qSjfN5oem4pNBb9C0q/QomMgWm8MzN
EZySKDiXHZRiGVjFg5ijm95J7sFk7MQnaAlOxCWDvnKINzBN2k+agsjC4ZefV6X/
pfha2Fd845AzZtJvHuaKq/UvAR5QQvhpqgK6EiowjZJR58QWd4+4Et4RnBQ6Vh95
9lL0Wm4Gl2yZKOmGDF7LImsQENTpQKO45uUOfo/34Beqzfonf0siw8WK2mI+iRty
a43lzDUMOlwrn2K8owvBTknb+4Eur1ncuVOaLM5i24EI46Osf1Qo5UAgYV61WQCq
UYUIv3tr/VHIs/66hCV+SPQJWer/b7LpBNt1TIWhFxUXjoBX+5siRsAQctBmEBOX
W//3Da4GFEILVkRSwLO672nB1Vw6a8mG7J11v9bqJ6Q6uJvASHn3XOQPQy6Ymr9y
JJMsMm88H7pyQhEzhsEO4UGLHrs0lVh4w8a17Y5G8+XF+JeSdRtndsXFDjYsUaqA
1VoP1mv2GNEFiAxurprm+rMtxk8dwQCIG0Arh6/2hyiw2FVIMc5X+DuqTLCikKA5
GH6qhdO88VyqpBWcu8v+UqL+DkEPV19BJF6ktZgX1SUiBiRAJt88Lu+Hg3jJB9F0
sObrZJD8PoSl3wkL6cBpr7Mo6q64J1b5mQMENe5ni9sUzRDmUYz8J2WV7oUH/lnP
HXaylqv248FtdnBryyXJh20gOzQFVZWK3ONtbByFtpTLWubdHjTZ2J50RpuQqWQM
GpIuUVJqnYnMt4/2jcl+ND2KAWjcU+q1fF8xrVcgRToayOy73Wi+lQDQfRB6sTtg
rDd4rbpRsVlGrqoUSl4bCkDqkFdH6H2hlymdu2Ky+3uuBmWTdGQFWr934bo/7clV
i3nWFEbCPZ/r3Al9u3CUvZtYcQfUJ1ywKjhj1PxI8h3RPA1hhzUBMPkgU+T2Duzz
30LNpKQzT1eotuURPOLXMrKIT18k29pDqXzWJrBDFkDVbhjqhMPaVnumpmz9bY0U
MrQDkPUwR3GcCgb3rFsO0jMu3b5QyI7+SYeNvsKll5uH3Uwf3VevAUQ6iesMepYp
KPUJf7TxustRlG9qO7dHfR9lysEIezvKAnPIJ5epbZRcCBZZ5PQ4o+jyGCdKg4KC
W/mEkumYpr/V6cSg/DMr3mubRKS1LAY1G3DlzgoW7Lb549xsMRvvewS8XIXXc1rU
5GMRqnrlGwkYUDgPmt4lP2IYl3inEkr+oq0e1oohlCSTBtM2d54KTRUNbvXuUgiw
UQDwwfO9FDa2pbKFLXhb8cRrHqxI/AnLRTapzAde8QFLyvx7YPBmC632TZ91ITns
BJO37/mwC85AUTmG1mGONYBs+yIzn/nVGZegzzsEWBxWs0/pbdvQQ1l3eAXuGRUa
E+9XocICwp9fLDFEbd9PjkwHaMq1l4JldbkrtoWPRBg5FUqYIr1z47TqM0a+Pjm1
ndundBX6T6OqyCOTIsi/yqhO4YGqg9v+qjM6PdmYvZmKwlCcqFwIJhlPkrSU5+vQ
m0sdW3jmZRcZzT7yRdIEGCZPRYRH3dTpDHWPYVoPyUIbZF1X5DwCcwN3MiTm680U
QU/zJgPpuYXEoUjPkNe3cqdjhTjjgQlqV/ptWd9cYejWJzZS3eWSh3TJC2UrUPcQ
41coRJzbMzalL5nmvOHZZj8Jw4s8nfq+xPwczvt0jJvW5LrvMjyIE+WdgskQEqA/
MO//TJ5vxzPY6hvCyqYdkHF8lpKjaYDYZkksZr3I4PMxVuAgWqVChACtnv0R8Qsl
YNqfUUUPIAhNLPxcmQzdHFN/u5B2tKwVbNfUNhg9PlOCMd6aUWu98i8/vSA91Vk3
vev0uQ9kLCwfBYsPOL5khMF5UVT/j3i/bZdYWqtjQ7pKEmE7aQVakL/LFcDOkr8K
xejM5W6ilugM7avrTAYfKIQe3PtQvdSdIS04v+bDyPM1ulXFv/j63wlmOU3KnoNC
Et9e2hefFrINT59U8OVe4IIe4n7NeMQCuVMSCgad5VaXbrevluGi/L2UB4Tr7fVN
C+zj88GxfSB/N/7Bzt8h5SuZY62qyILiXsylbljrsia3M35FwhoRhGFta8v4hFrK
Yc8aglbgJQbM/tblnTjN+FEaRhfXmtT/JKOCtqWDpQZdkQx8EOGMSq7RpkpSAe4e
zNIlH0vZCQXXqLLUp556QIbJxtxnAgQWDfgT2eEkRSicBGf1lWGwwbH3rXWD7b6j
s71YkN/wWo9P5dsdoBvZcQtbWt8U0fIFBw5MlXMoyXo8nfJYlHatCCTxrYfr0IOy
28Gis/JB3bQKO2UqH8JORDmIPXV+Dw8lFSwpT6eFijUykVQnfTkrJ4WwqgeZ9tXb
WCjp8vEJsmXP8eBx8mvY2aH4nanHTDfYajevRwvZMmy5kXfp6c/wiaNKu8cbWQxO
XWc4lzw1Pug1VeKfIiNwwsgim8fWiXcdPU3blsNEZHaylGxSeywB1s4FAnuOCLEu
JvY2dUBMZ9/TuXGiUUqnGUQtQ4WNAUJOodsLU0KauZbJOYD0l/0/j3GglyZ8Zmbs
E6zkWX3OghfXdiqTTy78MfxRQ3TgxkP8YVH9lKOpiJWsUIZgEYnQX54CuwWvqj6h
tSh7HbSKpEhZowhc2mCaFebIcrKKHIo7xW7FyZsSIBLYBvjEpNIowrgST0r1bb45
DfwZKrFRFU2LTX1WlRWLbIwO5wCMfVwlgbJ9WajFRr86w/pwQyUiA/W8Kd1ZV0Sj
Ge7VHsPaI9pwyDfVpbI9MWiaSqm/PucnkbVZdLk+J1qOhIMZNnVt5m7d2qZo/lWd
VXidlkYF2Ga6PXElkdOcSQfaYrBF+mBRJNmB7JfL0gntM1cq7yw3rY7slMIuMAAA
p2FyYdVX4ZyK69Dw3AwlcFGGFyHDbXRRHi2TPRnbAQvkQokEeo17y3IMmWV91m6Q
fT1W0OP+PxOmsRLpI6kWhMhext6nmnTfu1LVIj2iPCX5AJQLEnkiPIWFik1J37+z
bnhJmRPMvBEqMVzzVsDqKrukCGoTX/+IvW0hT4hyhAbXYHFsLPi9SwmRyDGGY7z5
RRlmvugsccS4YNPQu/8Q0xRL+U0qSQSi/JdwfaVtbbSXS7KvorrQp1tjrS1gvxRe
ZldoC0h6IsJ1Vh3ANdpMKujDbnMNbfukjfnWDoKgpNrIrTDmWySznd46mBRQwL9U
yhA1cC0wuRDZk5/3hXAESQ72ywEpt64fRtREBIULXY1fW6lxt8rMIuXZ+UjOm4au
/iSfZnIsdsltb0It4R28zs//6od8o7iElXa0TAmOaa+Yw/4L9fr2WznLCX5bRFd4
EU6zDIuXd94NMnvdOcSxhzff98OUJpi2VDnTCuR4GdRYmCZbGVGZeTlmApEPzmOn
mcFT+RLmcVsepWVFueIs+ItVRHS/XKhCTcIiI9bCtNwmoxJnja0TmujqwKvEEl9P
hU4b3GwZnMY1tiOxSR9sRkxG65Mdp6pFiVIXdAmTe6kJ9pVvwAlehNl1SUbF4Xi9
ArBA4U7CcrJhGDgzIjVARsvUrPaYMe+BklnfIjXiLVG8GXNDdwjeSqewLRhphUw+
9Bp6QsRPLWw3LxafSji/GbtBvo5pd1HWe14Cp8Aehtza5224iu6XyBoKJP65PWr8
T491AMBfDVeyoeFNvAF7t2CNQJk5QnEmAoLpLmhp6BplIooKppsw8fOhS43Nh8gg
BhttzVxZdFsamb/e0EdubYKXv8i/ViXcsogXht7mO9eyrOl6lJwW7VCtUIcTjpog
ZnBqksUMibMfAkPMI//UBQP6YdPOsCS6R8/pSKqVLBSquO1E0uqUrYIwRCyC6W54
nkXtWcrcsWJ3RuFEn4UbmQbRKDeT6IIQ1u1SwdqucvowN/rDB1ILmXWoyZFscyJU
UqcKH9jpdSfYukgWDOqfBgxsN2p4axvr4Te04wjtgiaaXSq26dEF+IXXJgUzvpRe
LnoCXVTkj16qx0acOO45VDtKJ3sBEPK1tBnturDMQjZi1/SLf4keFfb04AUepaHB
RbKzoASz2ZhWk4KWsQKGGdDog5f6/TKPEwImqBGLcqPgHygn3PjThuIGW9GSPRYN
o2O7M7Flmg0bVHr+mkMQbA/iXtjwnFdgpcwI0BMUZx0YO25j82Vuf/GtTHTlUg9Z
S5fiavgh3u6d6uIdbZOZVDwT7sbUboiRConKU6uwn1ZpABWE7Dj0ra7x3Jwj+zti
NojgtXscirRL0GgK6RdSitDwiUb0ZC+QOA7OBG4crP4nlCa+bH1uHqQyrxScGX1r
jhdzUNufECpxjzQYFNxnpqvVwr5M4OcqRwSi1AS+E/aMUeNW9hJXk3Q/qvT/tj9H
l5u5PJQt6s4kWg2acqG9onPPTUwsoQCPGylPHigmbWPcjr8BvgQKEZj72W9d0SIj
Y7M3bx/W2e2NoT7lFCu5hDZPJk9UVYWxW7OrOxu5YdvMyjAfPpiO/MLqaFvqdW7u
5HUCajU53YfcCFIuUZDXdS2SaSZFQtbnKOu6W0uIOhBBcKJplGA/34f7w55qN+aw
lQX0e6cXA7Ru74ITofQi+iUQpVsjxk5txMOpMXXMte0zp6UlMrCtOKWnN15yagzA
HqLc8f9+XGrzfuh2aReqnTIC8s+xKzK8FPOaMNfQT8JKKlI6GBhm0H0ViPwlHkWh
JBISIH77C0HlnxaFmcidbV6lP8BJzfFMLp+NRvcUEL/633AIQqFwhocO26l1awZe
gS7UanrrFNe+Q5+932G8i13XsTs+GLZgs7q2KrbB8iUdWDtn0u0UMrRRil/pRQwS
BKdlKAeDqGz0m9l+gPFDL7PszypUhDr7WVGaS3i3igMwnVk0CTtwvbewVdaKRZaA
ghKrgAWakk7tyreSO5os/vbmEDtVlaSB7eduDdTwZ6SGqAw8JvWHXcnmofbL+6YE
qUGHO2opc8JlLyfriFW+q36TxlY7C9glCFRNUGtJ1UTP8gPIxdyqYFaxg5tQO0Ps
o1WHk+cEydIXjK4bCVxg9iilQE6jX2gVvZhGzR3UkSS3zvszRYAtG1GhgEik7Axx
3HBpN3AZDWUBqLFMQzqRwCFnJXspxMgHCgSDhDDa4/OkXz5vae5DhX6nK5Y1fiIu
M7cSLpEcQfnPUVdYave+OwpCBGHrWRNT0CtgSCcVSEVxXbB9l8dIpn51dORTfBDF
EeVnlBCds+r2mnV0R7XZIdA8ExS7jFbFhvzT/09pRV66BT0BvqCk4velAbtLyK9r
rZcN881zN2/J/kFNl/DNT3qySQtMIFbUo0HQF33pvS5ZRxvXc/+DEJMxXLJWnnUC
QUD9LaMGKzul1wgok7NB+9pFSvF1FmfXzgFWKNGydKdH+hQf59wgr6Ph3/ZjGBnv
B+a6w1P5QsKyxD2/ENTYpPipSoixhUTOecly93erar931W51OFSZVJlto5a0Ayn7
zdW8Vrqg4cjI2xwtYZDQfgXFoDvstE+wBU5XoOpYIB3OvD+oM3zzjzfH/49LTSes
dRrUlG1VHmDF3MYiG5NNULFGCpmaIUY/agy0t2ByFeJ6E3FG9Q06VyZyk8MmeBIf
gAxpKbKvT99KFxEAc7nc21ihhYIrHUU/hyU7Bhuh9kGUn+Lc7Lb4wyAMEuSeNTR2
loRXEfJKy2rs2ALOdb22VU/gbNuwt9IUThxJFHv733djmgta452baujSA2MPejHy
WVidg6BaSfnRxWYwZXmkVopce7Q7XjO6rjZHR2kJa7shY0177KvhlC1Nn75wKuvu
AzKATg8MTmVRI2U3MR8eZl1dpnD/7Cxm7SYmmQfXUpBS+WPAvWW6P/lWWc+uzfh1
wf2KSp650x+r25RWhKfnmVqZid/W3v2HXukBZJywe69m9MIj8G1T/J3P2IYIIz9Z
aE00++4HHB5r14vIKsSjWi5eJRbBMQACkOYO0Aw2N8aCWZ9z7tFC4YVMd5zWBO6e
xG4bXpyHVDC8ztHYTZKCP9hrbUKR3ogVkmpzdl1oGim7lp6GqYASPDjM3kf3Jj5W
4blRP/K8ZpGpD5phIOun9npXvbE2vBZxldU2xGCDz/g2ROS+0yYWxucGoS9QpyOL
7A2pOx8ycMLelUyKAD8hHEzkpwJL9KIi3/+jDuJ2c/MfNEfpA1A0oLG/rINtcWNp
He/mNovSNgcIauNZ1Ssaqok28RoWxCUrsXfIpmsiA1XRBXJQ7A8NH1Gi57f2w6af
e31z/NwhbL/2L5uY37P8XiBIfc2xNChhL3SKJmUc8hm7T7QcoPWSsO9iI8XGvz9b
cooc7E30EOJrE6KoYUGQdRYmHr4lkSHmIWIvvi+hB8zX6yNfcGaSqVerKtvCyk2O
2BG6B0dkMSMfYfHvveyPevB8p4mjqQG5CMteDVh78PI/a4E4G5uwyprluIAHroAe
7ERA1DBU+sHqU+9svjjLu+T146X9j5TohhmVEjKrjFEnc2lmFX85R4fs2xPG7wHX
cMDI6m/chBIpH1O53SYDpd6NaObFX8jVvry8sD6//IfbkiYSYCuVt5KiycdayBJl
cf9XEPCHZFPB8Wf0AIU2dCztWf9j9CjLGMBykBldNg7SXQAXkJBxJkZUkGfZoN9X
yi63lsxiZodKaCL3xSk2MJ0cpO8SJrt/TiA6Xo9MvfKo5RzGT5FnZD3QW8Id8osg
JLFD4t5UNB/5msRe9pNcrttkQhO1HjNGiOKR0s9j5laS0u4TEkAyuoHTnWSR8EnN
mGhMeTCTbhuo14XAJBRVn8cEHtjiQeBFaq/1saYMxx4pd3cWCrwg7uEpv001PeCW
giR6I6BmL+j18mAtMZDSrdSe0iOfx/+KCWL0f6srn1/E8T1bktBoQdduLPVx15jc
jSglwDNVRDKIDL7aw62m7Pge2vtK1V+O8bIzwF9xTDQtI4GsUh/R+LTq2DLZOqyq
QJqy1TJYJCtYH9/qxKBDWncu6UHzTUF70wctj1KCMCHqtP9Y8/6kSymUeazGAH8r
izPpW7TUJ3/Iu94B1LJ7WcJvr+iZ48QI20Ryee4qvbq8Q/b+Z7FTZS2cuV1MUpvI
VVb2fEWx+k4e+6jpS711qXAKw45mKmpp9C3BbetnEX5NEpM9EGCDgtMvW4uNDMlY
vhXhYD3IoHbZkalXraKU2sbiUI+jVZw+0L+FG5vLgezTlmKpn81IGZJ/WP3tQVPC
rR3mnUUQ33Q4RjIJcdVdYQKZUxRCmiQ6y41wrLORJK4fux4g1opVeynZCs9RrQnZ
/DDm+B29nNzAs9Wz/FEyZhDskZzp0772G75zLJiQ0eZKqVrVNviy+JbekG1q09gv
WVateBmcF92W+sed8oG+Fq6QQAim/HDikfT23yCVrIehRKmwiB5efWKjMwSXzCT4
Hsm0UsKnr/w1E0OgNWChEvTN1+dn11HoMpnafc+Pod6N09gFfcl3HecoP+ab8X9t
xD8lWfs7o1Wrbe1jT9/6NKc8Di/uDPRr14IlpaNf3VTXDWwjX2IjCIEKWBJkMpma
3CfuobB6U1ScBHVhkXNThAiYK8fjhWoNjZraAIf0nkw9/3f7r/O5lvgt2UnrqRU/
HPMyFKaEC1WSl0/UM88lYud+f24JOrJ9unRy6vOjM8D320apGuzwlQQLbkG+lN9q
wktkEjAhdYTu7KfwI4kwDZ00UfbxHwZaT0h230D8ZJUbZYnvlrLM3u1H7iiEbT9Y
tNwh6FZ+JPpVkP+JGjPXg0vSPJfQOeD9GddpDhzKXECBhpSjZgXB4hCD4k1sEe2c
9YyzKyldnHLtsLoE58klSqgqPVPKYcNEAeKS5OxQakRY3I0GLNp4T2Gb710osEzx
m5B9ZDFfsDiyUnoTNOQmR5TMdSllpBUsVQ4hHTT+zGXDBioyOBM5K9cKOQivyAWU
UKwyEsUNqqt+aUs9m4eQj4h49aOVNw/ANAKMe18P4NgS0z0lhcfhDKYhdq9xlLx8
EEMDw91VwMMggvNQ2rJxMMSHE+CkXwdU0h4n57U6YXndGi+U44S5umB5vduBHBUm
SDyOU7RMoXW1MM5rafbl/9/komyPklyiOwd4zv5uHMkoGoR2HihcKefhf+kUXTH5
k6XAsQKdP7YIZQppOsoeyQcYfGYjifiEJoo4oVjRk2Bur61pMhOuArQGkhPZHYO1
yVtV0DQs3MggV4kxAKdbNmI1EWBJnWgdsqLaJFY9JIs6JclaRmOcKGoIoevJsBeI
ARaog38/0cqpUGMKctFkNUoZdGuMwxOPHOgC38PaT1xtJEaKAH+DQLF0+v4gPoxF
EcLQj8r7Ndvc9cplzY00pPC04ml6C8drf+sDU3xVv5KAVSTjqzEmtbO3J/EvgVEA
HRh9WHh75L6ccBaKEjaxn8qHzQZKT4vXAV8AjKdjFzcrSzUVWn7UQwBM5dPii4M2
ym8OMQUVAYoLLM7xrdIgz5gnDh5B5nkwzGkkc1hS8KN5HQIxbs1fRfipyTxsutGQ
HrFAThxB//NdvvLKCVIZrOLvTFH2dGG2iNl+tsHTk1RBJrS1Pr5PT8kt9ZbqWUSr
Zb3XjctAW4WZ9Wo0shDB2ZiGNCi0naIlJyphZEoumk7aci4aNZ0SkabGxuE/5cpw
24YZ2hMsxNiNazlM6GsAxF4UvFQcCi0tdPGMYFvcf3DpWHGY9mCY8UKKzQ+Mmvlj
MbuQPsMM5RDsgeKlLEN01fCWCU01panxNx98a7qg0iAbb3ne4Y0CMmnZ1DfzklHy
IZ/pTTD3QS/B2MLPYZmOYgX4Gn2gtlW2xX+VgLDpxSjrhntXeG8Kgdk9+QnvGZ/6
uMKYvH+1XVHvO11sfFrzdhp55PSJBVYjQDD4GRFS7xgTyAZ0k+43qCr/Jv1ALvsZ
OJWheZhkx0BgOjy66EWNCLQ6UKzJ7eKmyqMZnngVvUiz1IQFjA1cFh/VKKQ9FXt7
PHk3rm3tfPm0++RihnuHbrDMuFoV6WaNDqzoUxDhgBIPcmK+PQkV56o9P2nxIEeY
hqqx/BZOIRqMDkGe424wp7DoWlmO1+xDqie0M+O8Ehkkrrj52s8qJYPNC82d+e5R
VYFBPH4fUlW4kk7p5vCFh+Iry92LgTzDUUlo3EaQEDHzO3SapFonwteenPNTHYsZ
vBDu/wZPIhxGDCM9YRFifjTTQH1r/VZqt/nypnNgen4VPimrUsrwDa3h03XNrnN5
ZCgnyo4j0zq8jxIJmQbJAhUaObkQCFmmEiHKry1ZvL8XJXIAV3BYs+d0MCZ1Hbjw
QuG51SUbgeFoAWYSmmFm8hkUvv/hAoIlrZyVH2XUEmBglJ+wPYCq5XJi6kFAox8c
afbaxxq12mSVeuyarrKpfkkv5n2I2zrLLi+c22IOTm9HMko8+Bt4ZN+U3SHdFacW
udxQ8HmccRwRVH/TCZtrHUdye97p1xrdCBGTsaYYPF3aEz/O30RLRuzYlZT22Xn9
+ZYk+t9hZ6WnNShsO1FpH3gBLPuQAVinfjycI9F4KOYXsoEzYfplX74qZ8eWMwpm
19nQBrrWOK+5u8MZ8X78DUDNgogw918JtNdgT3IS9Nwnl3df0tztX+CPzpEbMr2o
3cwqvRiDK3tYU826J7EKsILv18yAjO+12SjSR9SXLTfb+GXkNmcwDsugGgdxQqMU
kf+aQpekUnKULJq5kg2ZLlSxGQonfugNCVxYNbdmxUfsi0pK/vkDtPwmYu/9BSQ+
1VuozTQ9yZHGYU2yW9BzugIBJbSNbzM/q9TMGlXJHBRtkTH4gDD6xx7KE0/82MQy
kSGLP8LAzun623UNEv8l0ZHGL26t+POYCMZec9ySGKhZzkjswlTGMG/CX8VEbHuM
Qbc3RctFa/6uynmbBTN2cGoennYMK7rq/gqxGrYmK6jRIlSkOwW9dAA4e+cwuSJp
ZzcPjCxQe02c+KKgpbk7oIJNOnOaYwR54pEbEyNQp3BW/XsGiOFLISZBnRGIdZd1
nMqV0but6SwVR8W7I/uY+CSfJIMrj651FsPcIaWDOSuUfneGpzyRRXUeVjmZh6Qs
dyGjdyNOrR9rBfEuZXt3cUEQbuuzWztV9v8AhUkeVJuHeBOfsenfTpsg7hBtkrWO
wSxcJt+ohDkZw/9EnLCn3GModftzXIzLSIxF9VtVorZa5FmZqMcTU+Ng1GygfNk0
duV1vnK7q20goEWG7SjQovjhVdak8qePBqnZIE9bmcQaAzuuWOZGukr21yXg8+LT
rvFXFEPLuXKYvcO6h+4uDUNEUK1KkunE7FSiF218OR9OJevxkbz4wP46k+sUQEIK
sPj3AlqF7t5grmLLyI07QcXwNfanqi4AbCosuxvs+du7zrucCEK0pDBiEOfhR5Dh
jO5dMwdqOY7IYUkoSu8slTQUvEJT6YSdC/NWNZtSxDlAlVl651vFtK6IYOMbLQ/t
iIDBve2PnWdWPr/KifWB4+f8HbXv7A94dubayqegHUPWJ0kBOo8+59ver/7BzzWY
b6Y4qF+7990YFQjD1jaVJ91C2YOj0LUSBdGglkIp1dU22+gDrgmVsCeO8XyhHM1L
d3ZWUyrRvmPvzr/OroBAK+bEa2VRBFDzqswqsIh80m+biffY4iAe1nYUxbU5LlNy
W4QIQk8eOfdjD48PhVMCnDylbPWSZ33Yh4Rv8hEPVAYk/DJoP6UXQ7Sv8vbAm2su
aufDNNf1irPbFoArVk9MfwS20QrDGrJGfgf2boucgbe4b2K4SZUa9rwFBaqVVxxk
FCw/nchI3j8zmygL2/4Ni5jZjl563i8MuRL4HXQVrovf3UXTeIBKeP388bCrX7ou
/fJOg7aez560n906sEZP6ip2dszv8rMkTgSTG0FKFmBt0s/siR00h4EsAs6J3Ajb
gnvSOV8nkfa3a9kKkuf59TP3q6zGga5HXUYhxntN77C/7SSg05P+oWOvSnXld8u1
bq1K2EPWIKFh4LdFHtqxrSCBrWYcazhml3kkh/eC3TvBO+F/3x1kPttBkMMpFFIV
seiaIQYnKJdWeWonPbDck3P83MkM0OyKMGs0v0BGUnWm3LULo/2aFAzg+xQQU5TC
cuIybdQuXZHcDJHOHZuGoF3D9L26ymRYj0wK/kSZOwWqBMWXamVNWhoXX9M4kab6
Pm7t6O6V4X/5rG5KY5Q8jxxRoknX08KI5r6GTRM7GNS0XUcz9yEpo5AT5JMJInLC
TlA7ilTkqXrqK3mCXeVy4WaLB98NfOYjhWb+haANrSymTpqsP+9aQE/W2QiKLklh
axB3Qghqj13Q5Np3Sk45AedETurtJ90zO2pFCRzzP9QU28/0xw9k8DmqPBiJwM1h
RW3XTmbO/vIS4PdSxfO/2rdHfKQ6koTRpr1ssYNA4d0j1KNpHbrtPj6LXSDAK2Aj
VaMsSE92zp6+evJSCcTURx64sYXNj5Bxiw5JvMW9XyI2ASdzbJ9NsF4Ta2WbNWhc
WnrlJ3ecIhQ82nxmnNPVOwoZPiEiprxjNruu6dgwO8nK0mExicivlxxgu2ImJmG3
X9cxCuf99c0ewW62iVulK2/SIjIHfhvhZrvTWzThIOuXtx9PPzSPr+Nn2+Z4HS3i
lO7V9j7VQhXT7SiE+D1d9qrUX+pv8srWSjYgQrufSkamIw5Ct8h0Lgr7JBoh203b
ksK3FEy1kx2XpwYsXh/Bj9ez+kAHJLrULZgtZOU15Xg9tuou2CQZ9b/jHuF1o+sn
cPN45xI4ZXVamOdSAoiMgJWWnPzxvbqcCAuAyxSlBa/EL69JZoeo8CJlCSUDZpO2
WbtSWGqkoOAtF71CNDIVGl0DLbMKnUdLMMyjy7DOUl7u54y/VlOKvKV7Aik2Cv0C
7D5SmkMzvJiA8G358NS1iTSkklYnLwN655Sa3szehWNpKp0OSC6IyoKhN97HdOu8
Y22AjyW3apoOH6h20RcV4GErpa99ZtnGazXm7Y19cKQUiapAjMQjCzsN4Ti1uV56
y/gfve2EACKCuHyIY/Q4rxas242D6sovE8C41i+gMgSeReFicvWr5La18iOn+0Vm
vfzwqyn93QEXg3/DCeHXk7RR9Pb3aH6gwbtcLUDhn5hE+5EdJtdqL61lAllayeFu
jDS6uwvKJt/XHBYoJAQcwTSh8ytD+m/vnQxlFwsL2XOjb6UcGl/fQXcY+QF5Pq6X
zaF2DWe8ZFNWWTtgKZ7Nbfi/6J/to7r0v2Abdu527cB+WJE0s9VAHrKC5AijnAJp
zEV1beuPs0esdPxU5QB4Y4z80IGYN1w14xvREi0pxPnOI5MbGzvjhR9WA37bc16A
QU/pWecHxM5bZeL4zs3ojaf6dnMY5VgPtUJBjU9811mIcT0NOam1+U493Fzmrwal
a/daLBSFoeCzayr+0T4ISw3F3QxrywGhp/KWI0k4QE3PWlqPQxi0lpU3Bxnxs2an
McP6JncjGk5uhLrn8pPStnZLzLiP3KR8bv07GQF5xSqpXj808qxIUZjYQipdcRYM
UG8iWIc/t6cdF/xPj1kUqWZs+WIHiMaltjgIj4cCZN7qsg4eTJRY1oCkyNuQBgjr
ytmHEQOKfH1eAWouul86/85piwwYTpcb/sr2GD46r7MSlEav0//FDztL9NmhSy7M
ZTzicWknuYiipYMQHaobAU7EWEdiD4jbbL+jfQWFEfxX7ehwWjbxVLOFNRsqtMQ2
8UE4nHDl8NltKtn+4jqHOa7Q6g8inkosQmUxhEAGd0Sl64o69m1VvrfsSOx9NFkR
DhnYsVlhgc5Lrf7Y91v5iV1cHJUvc7vQxnZMmIQkONrFYluhoMV0PJdrHWoJX616
NL2vEl+DguwBl75keMwCmAZSpY0MpChwnP21k+z0VfnLqiO9IvIBKGLl2l2XdEQ3
LWVgKeggZ1oXcZPF38SLpGqLqz29mI2de6YyoMDyE5529s+TxKK5+wm2B8fhLt+6
Q1+eaUVamNNc0t0TTSf0HAHwnqn/3YlIPbbmsbO+/Cx2WOR9P6dn5QmHi/gRTas2
4HN+sfhgdR6+sVn38d1Yx8G6Ih+MKGZgs5jeBY0pO2ROjP6vEHIusCG/ctj2GpJT
7O25zyGqChoiQfPpTA6meT1c4tdR28erBFRNnf+YS0JCF5wRk5+eCec4y6xpyIze
WQcNOYKkc3yaVBo6BONp2zK7nhPIUGoRn723N1kRuuy+729hZul63eU1frpwhdJR
/OAyOEBuw4tgrs4QurvUQwzLBq3a7JIylEgdp13rtYN7wb17L9MOJBigaaBoyByT
MZ6JKSiUwjPAI4qAKG5WUdwud2JBCJNeCM07hwnWckEhiMVItzv3eZ4GjBJ835Gu
+iAh9lbxfWJU/KA0A8tZtr4xN+5YGW8VkI79kK02Fyc9hrT/cDcij9q8zAWWS15U
jOLTgEwIJYEMYgd0V+9UUxkcZSn1KxRGHeMfnwRQlis223fIvkqGTsxNykM+cjWv
Zd3sRmuDl611oBnMg6LZy4XBseVi9HLUDRk08qoEjtYBt5cvamB+Xc1s/OaelguH
NBRc64Vpdhy+3f9cMBKnQXQAkPYNv7wrPr3+YMEOcy/65xJ/ZQFsivvb73FcglsH
t+dujBjDglPmZkX6injTojEMoEAPx8jr4zqf16eKuHueLPHh+pVqXWnQaslFB6uv
c+bRj8A/QVOXxY0N2xajAwERB5SUHcCv3Vl3tZPz6fAei4D82BJcfLkNc9XsfId5
M2/uL5wn2GPw41l7kkr6pFfaPMfqOdLPGBRuC7aFh/FvVuVi+EdXNXb2j5cCV+LV
AAoa368REVP30H+dcRVWiE6kw3elkqjFGdxEoWJQZPUWjlMP2l7vfo6kvk/bZrfR
uE8FaO9dEXVnaJbgqUMoMCmBPf0LwSmk/OoJn5riMYB3QnES5rDpnRQSX3HSU8Qp
QFgxHuTWGBNzDs3vrBa96SsDOxehim9wjMRgxK9c+x+fV3UV9AHdr178xv4h9AmT
2kEdUmqpYqbArdL820hwbV/eud+uAYrAlu2B+ImoHsUvgCwJzqME8d8uKJQoZla3
otWM7gaigONdexgmDKmPOIO0DhJFiNPo622ShAcQcKVTo2v5opRZXkwOh8BHRkXc
x0uOWVSEzpAgKqyJl6zTtHqL4hrA/ACV4T3HxCNY43pTzWAKYerFl169i5VxppjF
BWSpZZIiznISgbzv5LbiS3jon7H7qlzp8Wpfh0WpdDQexcz6jvGYflBQhS0dG2Wm
v/fcTyl1W6IeSCIoHyb89yLw9SwN0L3kEEzEbci5S4RylseGd398PUh402dMvK0/
AtC/kHdCw5/6GCpDIokIH5+5pJ/k2SQkJSuC513pmZ0tbNrSbLhu1lVnXvD+TtMh
tiwcO6ViJaTG5opHHN8ESgzww5GKhQF/Ppxk7cowNyrfShx0KBAqAvveZnuHXERZ
9yHRfCciTATRowcBxK5ZAuJZpcMNApDD+W5CzXZdYzD1JYLv6zgMz5JtBzg6POYK
MyvhkaiEQFgnkL9T7d0vCsz663vefjOajHFd6WIcazT6GiypHSZG5peZR+LH6sXg
H9al5t7JIanRadsXzWM521R3xVtEG9Gm2DIvhrUYFmrHyemF9pasfOQjUdJp54BV
9s3jCzPRZ6Y47JRbi5HBYgDBPo8OUzMpKS8Oouy+MHuxQgQMaG7Lmk5XyvYo/ctx
o9BP/UFKyMzWnJWPhB8vWpLMlzTICYrW4u+R3O9cvOIsIklzvs48V8QsWYjinIlw
Yb5anTT42yT7iHNVd/XR6FQ7xSX99uSGhQwnWWuVUKQXvUbu9raXW0qwkvz3KXX4
lDKV9K/H+BcQLl8WON99HpopUCOhlV1uVWLzMw341gOVomoKM5lrn3jG7hL70b1Y
S9aItG/OY2HjWT2ZcjhvmFetHItqZOIZmgOY//7/anY3cx3jHoMkQ3Zxa3vfNyBT
pjED2H0BR9QhoPDtUajjJqSrwbteeTuzRyh9SiOGe4B0sboajPbT/cDibjqVQzIr
gkjIyHqTp4c2OnUBBoJ0EMQw8+32SX5WBkRuEqugT20rETibB72QddD8vHPB+edH
f63yFingqF/pDRbP9iVKqDTa7rEI3vEAFi9BNmd7jnynvaPSSKa5K1Olc7i936Jg
ksERlMYvMK/sw55DaRJEbbex6ZN0q4uFZF3XbVov0A9qD/hSUlC+rF8Ac4y9W4JR
ZMTlMectlAHgsdH6RzHzIz/QJ9N7fggiyN5MKLOzXxI2rsz4BTsXhls3cxrg4R1x
sHtx+LnIAm1LqX1TQhUXnr+2ST0aZyOCcyNE5qZ6sFiVNNFUne/P5NxFmPBLQxwF
0ssHPhT5s64cdoNRxcMajll555NK8P3YvjiajzpDqy7bDwoAtlH6CG4aEzSDGks0
QrHjmnZKBjbsdhhLuuk7LEIhdfIyfJDH13NnHE75QSl9JiXFQyv7ecMrYXjmRw7e
FEzeN8FY2rSam9E3oko4kaa1wdRpsTjQGBwhOjbAIRKB4QbhlKX/qCbTGVOQGHK2
XLk4akXTUMjSIzRESbAN7KLPpG+7JvifDBc5eckPKczSXeFBna1gUBKembLr6DFt
FF3CVMIgqZugq+Wt/owaDN4fUd06Rcclg+uI1iYZZ8FGOrWhK/DeTFeqIQ2cKV2k
BVNn/3SrKu28rZaDuUTBDYOna3Vo1Q1urdCv2eFLyGdgSkhysizPss3ZP3acB+rz
BMbm3az8XBEXggQES2k0R8g02m+KMeHDmfQDH8o4JQxGrzUOc7Vmi6r5us0/8Xth
cJxPudBBvfonlsgFaZkQTmigLcmQD7/Tw6W58u2nq2yc3spb/d/McNku7Mt7SvaD
5KSKEH8+saaiC0Kryr0OBn8PYqC+xUOLIOk2wtD3nBJ0DflfYLVQgaYuXKwPdAOO
Ahwf07NgDWsG7sO/UFAhfdTpZ+vWfRmvuJaA2HqrPNSdM4ctVRNcHTG+9NoR3CsP
ts/NY+y+irxhIsSjAnyXWBejV9wAbrE7kg8ZgomnlqyIvqhve7TrjTKPnN9EPaU7
+Id8mA1lL3N/C23eh3WfuDRf89lemoVwxIK1nrx7/ynD6D3BK3RRS0lUDoEziRXQ
u/2payUzFV0CRc92wurIO2+vxsCwJqMEjycvIw39kZmVuIerXjN56vgBQdvqEm4x
HiHpJohkt8NBBIbBgtDoRWsHfc0Swc52MaljvlTGnjZhsEgcMqLwJiVWPbnW7s5A
kJQOySc04VzrrDKx4zWx2GXQQIuD8wxuBpKT03KB1tBuJBRNKQ0qnpRZXvQNVRDp
7/31JwLSjkevVySAhvTIX76BOkJ62w76aSngqBbTaYPAycQ/l/c/VxEjgyKig6b1
YazEq44n/d+KJKO/gD0Lt1dVcN/5NQRESc2WbQfbU/bbo1xasP7MeqaCify40gMt
x3ZPUpzL3hTIhsTH0pWCr7ha+yOaytAulheJNid0e9+Feu4K+CMfP3kdTQsaNKpb
T7CcYUSiJP5OCrfZX1m457r0Gzv2w3iju4ravd60WjQkCshnFp6yZ45b6DbSEn4s
m+bbkWIEFgjd0Bt8VqMnt7eldkBihO0Hr9BBcadGI3XEs42x78k+kViU62QCFFga
6V2YMwffdXeBn6WGJrfKY1FqnDXTy/zErFnkxzK2lruR4R5tCmew9v1wvZGL8uzt
EADdIWwLDycX3TeaCVbNRlREzNGZpOOpqYscKFAhhO182YmN+2LrTgO0158zdpqM
Ws6RAXKVorK/kgxUZHOwERLx6GxIqs8FoF1SQYBQI1LZgBhxfTDPabcgSsWRxP/3
hWpaTy7XyWc6gD0HKt68bu+TerA9rnP7Oj6aoLNF947Qefwlipfl8QOeMJUDfEMY
XKoCTiCl5NsjSkpOY5Kb90hWsnHuVQlPk/WzgPHi2Fj5ecjqABxYvPfRZoZ9n97z
Jp2Zm8KbX/zcZtZ+sWNZj+M30I9pNbx54ui6SEcocIGxFXpIjW8Oc5buUMZrDuO/
H8QuqPJjEdjdL+rAqdrJebnrIBr8P4hNNclv+k1EwB1LG/PDZLK5Ev7PRDYMDzfW
go6JbC0NbuNgJf+alIQyYVBVg+8/HxXzYGQPv4WJ2cO4iNi+AUqqoWizMCKeMgiP
8Y5UfIRV6PUVwiVJ8QNuxRlK38WfnlGphc/H6EGfACpcHTPH8KxAtHOOYwurMrN7
RTRc5tqfkMTq7HerJlSWvaB9p07nfrBjv89YDa8IELjUt6LNEzTqSH9SY581jpps
E3WnN0gQtfQ/evIsczL7hJe3CzRqARDrMHRdn/j5w9OfE1Iu0WMZqvnOsrwObaBI
K5D1kUXrNMdAAb2hAIISOIr5rLzNKN9Zbk+Desy/gi8wOE7yVljd/7g9S39q5UcD
evArgYeUPg4g3jGe2Iwn+9IFIQc5lcIRhUE5e6CfKcTtWrBJqiE0Vr1C7JDC4GM9
CN2BQwZpp5SXUodYXwT1+j+bUTM38ca39DBVPbjhPP70P5/f/CTZu/wAYUlVL8We
XYjiCpXgYaK2Icm49Pae/jszvjDVqnCz6k7N5tpHXyA3LthxHPE4yaRxmufjuigJ
9IYP89ZlCefbo22cwKNo199Kf2RR80pY8gCpVlskdLL0TN6lYBwsyZI3BS7kcl8/
yWQasM8XPBj3JtAPmuOTsI169THYvlnpMO3SquBi6hB6wRtdmA4Lm4eQMAariZ4d
YyNWoFVtcyb88bDHBX51dcwpLgLYwAEe6RgeBqSrEQyKVQOhgyzuwM/lYmmeTW2G
jYN5crOdO/jVfMoTwD63n71btliG0VHqm6+FIBD8wzJ/BKSrh8Scxak7HjBvj4LU
zM8VGOUHPfTuN1PGhhPTKW6OuZ5TaJHaJ/NczHyfvlpUZVah4c6RuCE03wZXz2yh
OskLc9cVn/3hiit1dsa6FQZOW7i+nFZmVkACeVRzyq+n+rHk1sLM9yjwKC5tGVfe
BApPaQccxXyBmGHABvaRvZsOmDNVEHaQuHvuuSS6AGVFXTu9lNeDEM0ElRz7c80W
ba0Lu7LQM4jZREERvuYYYJlMiKAGi+4XAeTxlqsI7EKy+jHlsAIiqR4Dp6ee9UBR
7Up9y/VtdKH4Xzzvn1/HvvZwD7iC56A0xeG5vC2t1qA9uUn8ynjdXuBFOKRU/Tf8
LeoTJ6Dy2ulkF73JxE2Pgj8JwXd+GxB0PSP/Girq44DCQ2Oc9k1m+/3rXc04R9g0
2BTLhFiXmpYzFnQDDYKC529M80GewcLf+cu4GKV+nBAE5t1lBGolB7aP6wunDyXf
FObeCVF7SIXgXgGK7aXqFIVWuEBED4w/+Nyih6nx/6YYk0f76m0nUqy08rAm/M1v
cmQHf1Eb3Ykc44Rs/3nUYLfJ5o5Jvi2bjQtUfWwAXkBde0ln4fM1GZltR3/NwV69
p8mXBZPRyMMLQxOJSqKR2nRgpfKTLomL6KFOM0KQbE8d6jTcqHj+JkfCZpBl5dGv
xHMGTcTgigkcRumnXseV4Fr1NE/36jLmbllQ+wM6gpopONfLxgYKN8BgDXvyDHlq
YJLuUxxP1I/ucKCGVwDTHFc+KuJ0NnlNqPhFu7viP4x5a3pnS5Lt83PQ6xnrbhru
UI2DG3EYO+YYo9sKXj7u0ZsmgToRTbi1wUyhaFWcchdaTTJsnKonBiDfSlWH2gLN
OqJWQ5nflmFGLNvB4hIN2UVDUcFnHJLnw3DDueU/LHYkRQgL1heIUviqxNd3ZiJw
vs8PaxP6pnd2QZxRH3BnC3aPtHj1fQSpvlAMy6Z7PZAbiQZ7mxxcjXGwO0yTVPZn
RbvZ6yQISTgFf8eA+XPElfwJwRpHiaSS13qrYWe4/xllmh3X0bffju15C32pSMIv
F4HqQRoYfLXnjLICiyOn4PpszkQzN12Z+rq8FbIuC8wnbqfQGzNYSvYeQgdySKt0
GP690zIqwmX4ZBFuuSeDYOAzCQsnM1gzS+iDvDmrmqQ9IRu9Rhwzv3cK0XoKfCzU
THx6MKK3lxdtKUxWf8QgSj8erYrN8EpwtdljOkhE1wKDcpIj2T3ou27/0nYoPga4
mC5qPBulWZhFSJmoqLRg0jlBdpSFsTvW9IHevMtH8yqCMVlNwfG4Xndf9E7l/IRO
4kJWEj14Mu5VYn1ZHFJ+26qYTl9U7XO5AQR3/t5vbzsd/NBSjXeUhcA4ha74ixR5
67+4pToeB0IUfss7fz8S7dzQg9Ze1ABNANzXpDx0Ju9UkWjin8JFVif6td9rcK+p
QI3PK1kQ9HOEMQukwsY0DYj+4BOLMep5NRvWU2mHkTMIL6eT2GoyVMaCgDoihlpX
HcuYZ13ptMY/wFchC7mpWX4v8hbPjC/xYhlnUKR16Y8cJGIgdgLdO0x+OICsSRqC
bGlgO7QbQdfDBa5FhgPbmz0+iG1D6fz41hMS1hCTmXtfW0uhezD2FbBw5iVlLEry
qkSVBDGtCDT5bahKHXYUCQ1XtRgq/XsBfy0y4pKA/Umrgp/N0j8I5Y4cVKmZLzyp
H1vEt4n6jer0AcsMalFKBokNh1tyPIM3f7dgOYC0uwjflQ611TBYjYt5OBgDsD7d
xXcnpf/QzhTka9DcfYRdpq5AvhNYCjare9+O4dEMr44kRsVCBFPS4rnumQUWuc1H
ldhSQxtZuojm/QemyXhF1bEsXjxnIzrGc5Y7RustAS+Wigjt6Y2mWq0OlvDqlVM6
f+9/nu2bl3vbnnLdtt7ltFTyete8unWvbHvOOdEQHdIooti6Q5polOs5PvzJBTob
EVuXLGKBRUKUf9qZzHpnEnWzOlStIyC1xx0K7oCyaIF7O9BLr5aOmqLRz9wfRNlI
Ce5/2GasnTn3/9omX1DRlE52hWZofC3YYVQknzQgb3RSFsVULu77mD/TVVyeRKVw
OOTaWkD9RaOAYF4dYxdk2HRpLuRp1KvT5mnXtd4qEElUfPHjp4EfDApxWjqDefyi
UOnCPnEW7F+ljLjWoYkSWPorG7Vv8Em+CH9Bd8exgqFUnsUhF3Yu0j6BHnDQT8Xo
DxnJ0rHVLLDqiD5wbM1IfcZdQOR4UgqDZh/ddz0RnRARD7cNlGpa6VolIG90vE3d
qBmec4xuLIHg4ONfSSsFEzAQqww+g78MYj8L4ewIOY3eYt25MOUfGoIvfLDVH33C
q2BPaMciBhfYGhRP9ceyxfparuhTEqLA3vdK4fCiVFaB8K1hFqNo99FVL7tUOkwF
fmn2YzvkuFLGqfe7JkCnM5LB+/w6sRsitxLpxJmd4bKmE2fSjNeDrnZEjw3RQZcL
k5yAMTW40mF0hNzjbbA75SlELJ7ErW/0LaI15wXAzbZ3Ya842p269p0p9piwhQyJ
B9cYt0fqaPqQvmFbU0cs3IqWeUZztt6etAQgJz0njhW0jvzq0UcWjEGnzoEp/xl3
kSHEkapCl/nRr9wCdafakgY1J80LE07+t3ig8v+UwpC+G7/nwUaR6spkL+VuLwkF
t2Q0uMvhB6xZU6sSijx5Kwhq5eVkVaYts3lDmnR7mWO1IZkKRgiypVaM3eTa99y4
hupNtmj8SEjZajuW/jksTx6LOfRu3foGrESK0GBNSzfosz5BoG4gIT0t7ZSmGL2Z
U/p3pyE6bp2ENsWQyO27qY1EP9vap4BY9VAF94XB1ZCIbdE6SNXuXMhnSn0QPZgb
O8a/3AeMH7eCapVzpTyNo+FQB5M9DMmiR5czENfoZ6qED11bvF4aOXw1kR8KDSov
lU2NXfncLy28RLDiVdwXr/Ox+geL8EydnZNgpVTXXJi/VPfwiRFq8LsHUe7eV/oX
m6SGGcywB40a1uY4iTwJrKNSUeHLQPJjlPm4M5g/w0Y7t6vz3Q6ynPWss6l/mZb+
p9TZRimkkHVxeb0qUl6x6Zn33sb2aTFIsCO/tkBOb3GPi/OD7Fd+LbkPDYv7uMCP
3HdXYKZL5D5KHxnqswwbsGbr9CNVP1e6dMYXdsAkDkWqolqXTHi6MYetN478CYWq
w2IrIMkeX/wLVXdz+V8eJm87QrjZHMRdKFTgV2fOq7JP/rMOL8qHvT92c2XCaQpr
9JSmmBKDooGI16BeO+r0geZ2muTKp+RMR6G2aXfCcuxH32W8AojDAbS4dH0bnwcY
EkF6hb3EvFhFlzV6MtFfRCQ33Tv5smOiWA8Wn63zyLlawN409gO6i8acQ9TjTSX7
5Zw4hFoiDp06fUZlV0fCNspLzUKjxuRdgKaj5V3m22FJ+HGkhD5RAkthn6Y5FbMQ
zIUv8853BQ1QPZJlo3ZEI+XGu1tKLqOKygmATn8gFuR4FE/bGIWmBn/S7GvUv1a3
qpjqL/4L4kp7qXqaBeKi6+9QzRz9kG8RLdXJbRikU1mjkjzCy3fs+rdxYdhJpkwE
3HeJ4VCx1vFoe3356AjI8uP0U64I01096cDi4AiATiw/cj0WAqSu4WE1YF0NXI39
20TARgezwoAM7ruQts5bRliEv/4bQfaDGYHY1lFl52zbnyfxA6oAcM78wc+P1hxP
quDXu++z0Y7pvcTWJnwswqzghPZHheuFWiF9nQRH3UfT+rRv1rRYZB6m5Es43eiY
LjDFQ3SZYQqpJrepafMtJZpurGrxTr71L6Z9qR7kYBpe4ZkROOXgkYK9juMqbsvU
BLllLTl0NHE89xTVWruoJdiMcIw6kaSiWZEOD1gzAxudWcCeBJyjQzn9arQW/yyS
fwUV1vdc5J18vZPhC+bmpPx2x2A8uOsnQx8RzCTIMqbFo0Vv2cMm7hnLrqj7zKaF
4KJCZIJ2Al3Fm6gboaBfyiRlXFExtTZGhYvfPwBP+ZWLjRTyy8RiOYzCepVKbFHd
eufQtWZo3kPt8p+OSmo9SHw9GpqJu3rYO9AvEokjKBTdVZ6umxxR9Tj8J6h96tiZ
8Jaaj1AlGbNuJbPabm78yGZ98MIvtds/S4FyR8EOsRfvmRLfee/tEVS7gXnGhW02
nExZzjS0rOhLZozsmbQqikQEVGWktuARUNV/LREV72iuPVhNOlsT+nkojj9XR/S8
RVIavNAPftrcPGAdQGnpt0JfNNTHCN2XRRRhxGr5LknB+RXwHUyrL6TRQo0F5Rgn
Q6mQg5Xh84+bJhLDsGGY6RiM7bGBy6Z/MEId1q904rUfcsBXeiNNcX28ByV67S7A
oQ1pAQ3k3JeSqUSIPimQVh6pZqnVJg+rAqMIOF41M0PgY/EEqQanVZnF77BWQgAU
X6j/di2Mp8vUA0duCWmQw3eGCCXlW7F9z2Uu7EQBjwc8ItePXxxDVYZ1QXGfxo4p
CeMG2keU3ummxx2SsNKrpi0iAOhiJPKIpjU7oiajaG5QSFMYHAxqTm39yXb/xo4n
hQysaoRnBuU2ZywqpcLz1KpDuX/ganL6FJpYeoqYj8tY4a2s9as85aXWyLP0h2zj
q0NY92H54ltRrM57QGwUPbPZnyQoM4u87rFE6nnh+FHH/ZjNSNWs27n2KcesRXVD
Sg/Hc8NVPGVEGmxd2kkXnVsF8R1+gm52WBjBYqpoNVd9z55tu1CpuDBcufcgNzOt
LYSM3SBDhHaHv/adRPmPBbF1dIaxvw/S3NP8D6LDSvDaewSlDZLrSlbsV7S/iWlN
NLK4ikx19d//aPEnrmAuSXeKfyaeczLRLwLjlqa0Wo23l84Zot46qtKikfHlNyPf
Q2YRDKfHC+Z+cCSUrTZzA1Pe1a4hTrR9V4+3j9HVfwOH/xgfgoAeT2UoCn7hi+4s
BrISCjALR3CO0cRZwVXgEvQDiU9Us7zlGWlZrESFnycESp1d22XXfNrkTTpVgmwv
6DfKne6iLpGBA+PUfDo7+QER/xKWkY1GEiQuUPg9fdarnjIHGESss9cM4XdYJ1/X
rdsd0rvLHyBwnbUPWAhjp88iHjqrmwI6men5/hvsdihRcZ/sycQkB8/tdp3huY+M
59X3Wkr1dKI5WwSqqHjDaq9Z0MLFTFROupM4LWZJHeJqmADGjTbcGgK9oUCcaRmj
bIcvJlWP+wkHTXN7L2uBsSuM3ZQc8D81B2z5SvlUU98JtzNrKm7zROXO35pfJNuF
CLaJpFBvT3u7EZtfgqOhQMojNyEs2SIt9UHyx+yh3KZadEkTzkkU/Q1onvcCj5Xz
s2AdFW22ejl53pWF2NscRyxYkkHxrmq4AuSkRMX0iBh+G3rh2SHrmmpEXjDW9K1e
fex092Zzfhe+MGV9y8xWYC4mtplDF8H62/1HHQmPOMnWtmcxdfxPaLoKnEMWsOrR
LXLuAae/BYlgxvMq5TCvvmggpPbC2pNVlKHmX2pfysMqE6/3VoTtyxJfJeUt/bil
bd+DsAOVYd1qEPrEsdN7YNCTrCCvurc0pdIKxBBOh72jmQ+07o9UKCVOMuC71Rbs
UmBgX6nAK0LcaVDSTG0em+BLHpJkwCpv3sD0+RyxQsReUsP9mwehIoAWZIJT3p7E
IfuVC81ee1/KyTP2fLmc6VrItCfocgHTTfqUuwijXZSErINF8ai4Gdie7fmPSrLM
5R9oaSRx5nkq0vCk7tZ3EJza/6uUToWV93rNS6PZWIPeqlLdADROighYcxORn9A4
w5REnOioE9w7Oy6/DQ6hjceFCuhtuds1Hx1Vq1cHn5NbjIN7JQ3Vv5SM8C0z6ytG
1BiyPVbjTgGsJapJzE46gkn72gxWvRHQIOzrAvMLRH48wNZpDJux6rtGucPKeer4
2f/bq2a99hMhNA6EUDHVYCqV9UEB8OrRJcyNo2XZ53La3Ep3SN8kSBgzLyMvbPCL
ZnkCjIaZEgDlboWAKDuqFcAVnS0aCQ2uiPAs/2ZEcQwRgfIOIAAF85PN8pghLuEw
kSujQivlbPWtaHpNgSD/D4dPp/aHIa644iOjzfuudAB7Iyb0JY8jFJ9OQukyTRP1
mkSV+ywQCPADl80dF6uEwtNTLw/cnOoeknx3jhuQ0ymlxgM1SKLqSv9fezG10A0q
iblCb9E8AxWa4Ie0KwDX8+kfCFA6IVIkxAo5lfXKho0xNgWRpLtRJX92F7D/KjAI
syVFznGAxaqMbVd3F9n1nmSc6NXiotjgW+mBeHkz5tCzW12iT0Ew0zVVPDEDDQTu
7SNeCVBwvag2YwYS+Cp01oHPmhMJajuZx8vG5Q+9FDWqAEmRR0Le0lMElDuvdg37
w7xPl0D9hctmTOuk5xqnvCPEetLN9eL9bLIjwLHz5gfSSFGKWYduWh5HKdlv8kjv
++SsEEqaysdi5MZ2xveM75YsXZ85Dx4iLyVtisNYox95tC/8ntoePJyTW79mJHTH
dpB8KXF3CsCEb0do6XwXoZYf2nTElF8uJ76koah9Jn7JD0zWXTtCx1TnjTq8spB/
VF/DnYwKHGv/XHOysnem9CJ/DHTOlYwcoRfnL0WHiO5QlgR8zSwo+Wksiw8liqJy
Ye/kfW575nabKrvW/JM3TMyrbEVGhqKhojVq6F2KOc7RSwodL5rrtFkD4QsMrbcw
IEcgegWXIiY6DM7U6iW9i8GsLFmDa75rgJNl0l9FvsDy+Ko7aecGbNu9OzJSXLKV
K+7U0Kh+pDNw+4074/DAdTJHyxJn3sA5mbw0GryVbdQxutuF6THQl+rhvRJJyG4b
G/JzWmXjtwjS+Pt7lmJkAGG+xDMOr3FJmVObyqNYq4UyZN5aOuqvx0jZtjgMQp8p
Rn4WsFzuiDeOiCJUlQ8KrliVMrzReaNDakSVOWF/BZ9wA0giG3fxEM3Y9/FQ+ta5
3geAvMu0EbBzx4VeWESgKiP1pFA+B/N3981z7k0xvlvep/fBKyViRygDRHdG2YBl
9mOqOZ1MkaD9oDhVMCy4GpE5Ejea4fNOJXWADQh+f70pBTjM8YwsIjrqVBnrtc/q
0cojzWvB+wIeFgwTQ86SKDwSzV+ckARq1cD5nQPhfbHqFW6RdNdvUH7St5rJWolZ
oVGqLawZAZKR3R8spZ0zuwnQmvcWv3Is82S4zHrdtWjEP/tp80WtFvVbARMgabP6
PjhVAQ5+WPifXuCkEvgg0hta8HD4QWKmB220RCANigJZnHEt07u2YSv2c4IaO6bE
oIgH++Zi8h6iAHYB9KhPtFPLYFtulCphgUv0AtsgMdtQRRJGrsSMOQPh0HODwkt3
DsesCemSa1M5Oj5RrV/pItIN0obOgr57uepXb2tezR9FERgkeFseCjNl3YNOpH0x
SCdRZa1gg4WdZhH2fCmC4KefnFRii7sGW3XvbCnPmwG4GyOLHAB/nlhTLWeei4PF
reysOVD+Nsxrkz1ADaJ49CYOq0D6O7QZRSWhKD/Pf9g2Pv9/19ECgn9LlIcsFUXO
C+jfPXSSs0lp08jo+Q0+jFKY34JMImFB8MUsW6P5YDOlh3cVBL2c9Pkl88sToHbB
Kmp8KEUprYJKcpVehVD77pcu7CI0FxPfDRNBETeuZ6G7KMg02sSFOfO34HL3/lOr
UGZX1z/6A/39JGWIwl2b4AofJdYOKNzmFHIYwH2K2dqwDN7cGbrwjGKtXRn5+X3x
gROy9pz5SZeIITy946fhZ9Zgrqj9S6Z2lFrr08oZkn2UePo6Mh3JD+hmfSoQiBFj
jgTbrxMR5pX6JqM+dPNGLYO2pM5tGiVQIvHo1TCMKbN6kn7wiKk7mufFwYH92qR9
DHDOrZFlTjjFDN7x4zpWbizOfB8b6R4M27Zr7AME2ay3xWzI35Zb3p6WdVV1NMnw
R9cHmeSmdrYZSKlBaejb4Uh93dlmviU68p1XC1IFmWEurueqZdegiC7qcxkQqnjB
vHGujqY/axlNurD7Nl7NUIuPsfAweUq/bkvnMOtKrGSnNc7YcWe939cDKn8qNv5p
Euj3Va3hrkIXI5zkslRxdt2YrZD31GSWP27YzeJtfpa4cE/RrPxSJTkeXTplwVrp
ZTYDv5s7tQmlCimATiqyFs/Ov568JsFN/U0kPZw/Kk2QCIO0t85o5DvusrOfRVKc
2SuYuJJBNED6uGsbVYMrI4IBw5NTjzIxwd12Fc1N/YNfb3t2TYyPQZ+0Ll0BuHFQ
fPVVZSgk56WxVjq/reb0B7QSpMy83LKlrHSzrzJHS7N711ayW6cnbJkYZh91UREw
sr4E45Iy08TsMbOFigx44L96k+ZteXSdNbWMSXp8r2xpQTwLqX4hTmzoDtogQ9cC
zkSIv2CEnLCC6BTRmKkVh5YvN4TPjlSCPCJ/XBfjUlHbWCKqrZ5wkbpyyt/3/Ujy
8Idwi5OWlL74FEh1JDysh/8Rq8Z49t69YbQr7t/TJkyqKo88Jzjti+RD27GDJs6c
yXlvnIvyRa6+dE+u0sVbStzjRQTzZLQ3FTQrTEoTL3mFL8/Ab363DVUGq6FxiZYY
ZoTKK+Cvh+zO+KYEWAUXQtdCzcMcryUYepiesKHynbjPHP9WslkP20Fr8X+jGkXK
X2ZXDMGxwYv1Mgm0vGvpRF5vUIHnrBo3twz6tOC6HaS+9K9H4HkpJgg1issgYYUy
xBlKq4ynU9aw8BcBdis1l7M4TUGDLQ0zW2mVotgi0rR6FkJ4RWzodA0KOk0MKNLm
HMWQdexVmVPr3U+CmwyQSKCoC+Hmo2rdFvNQwEskPiunptzol0MSJZD4WX/FOjRU
uBlVXD8EhvAhcZ3Cvg8/SZ6TnTAGzVW5/FZp2oN73H0d7PzS3ApMq+BHsvJlIGDk
IvDbY2J+8Y04M502nwoR24Vi6Rk5dateMiJFAa34NHnKnRDKX2oBbFyy3QoecwQo
Hbw123EWbK7NjMhi1sA8MDR4AfcNe5DHSnWwa6D3W3fkmb0WxybWc+hU9NtnYVbY
CxWQpvTeA761pAFucQxGlQRiBFQcgdk6SN2d0Jr4tfV3xjAPO24KDlCD9k9d2lxF
dMYqTgIgzxEP0zf/tx3rL4ha+P0vi9gCCWm5MJoAmhjkbK1dkm9alBUdynWcYfWp
X7oNy7RbtbHt29LXLSTT/Pz9y8jdw2RykY8v9W3nf4lQQO9lk2afl/Ja5tqLB32Q
QOW91Sg9P9pZIqJyLLVhA2/KMfPM20d+X+4uphpQMuQLIOky56hs+OxvblC4FeQW
H4vshcb/CQl+4sp/JRVhckHCANoed4j2z08VsBflD7KEOYDPTRxFN4iK4n3LZs4S
qxe1g7lBFEppy78p4zw3ms8A/ZULLd2iwDelBvqPfaKqmlnkKz746cCPnSq00yKe
De2UqZtMenN2Z2R2DDPswEsRzwtyKjWNPvVA92vsy0t/lqNmad+SLTwQVzKZ51dh
tJno0YWdCTcqAEFnz3buf+LLZkenowfYBrmpL4ftAT4bDqQxnnrMWq+u8bHwQkFg
cZUKY20ScG5suAIGCZDtMOI+Zdmb0u/Nngk9qkasARDYzIKR7xOUSgxZ8zgLMu6+
AowBfomO8rgJiSReRG+5sjiVmPqDt50GWdI1fyehnjpPwQ3/A/eWv9Gi17GGcjxA
dgleSOJYuVovWivcMCUhs0llGyXJmC34Qyzv4I28TXV3hUxX+EgHsAM5x+4RiYap
4BYjM++3sYgsN76QcSFgp2kd2SjOILqsU8BMIdB8b1Xh2aGVW1DJ26y0AzWEBEMH
dRbAhRCvu5lcLFhnegFQJLL7qwS1iMSJ3Y6mXnI2jEpaOO3SbSVDmGhhYvRPiZeJ
eaxnwkBwMWR/cvBXVqwnocGYNs3hkHPiLqlKh7BhCh9RDy6pbr2q7jEjh/pYo9+i
Ad7ZscMRQ7qVGMZWyZxMsIrthSlOsvXSSknKq2+xeWjeXXWngpqdSAom8H3RkXtZ
0siq1x9q9eAOYjbwb3r+NevshdBBSb/qvkptEAe0BGWOf/u5xuBQ49hc7/0iijAt
GyRo3S7rwG6jrERXZiujEx49B5t8VfckCAr7Co2BCGi8WcLcRVtzJIObgZXhzIPr
mGSSsvwKg9NWOM1tjE3B0NSgfPn28Y1ceER9DA67anIM+TMY+3aPhiHpW9M2j/nX
kxwOMaWAtFBCNGuJXly2FpPLtJ0Pa7dWTqkFCb8Ni1OtDvIrPzyLYgPTGADDOFJP
W+9qnKTRjmlL61UULemG5R4Q574To8mBEPp9vvPbfLsgGw+/jU2hOB/KymmgpJWv
XL312QyCKgYYuK5sv9izppyU4PeO97/twbmzQkWqwJgbZogEknGWMRtCvVcNxi8e
aj+RGeml9AkBFohM50MPrRNf+cz0VGBeF83rRYj+SxNsKayAAjt8h4q+KpY+w/JB
7Pxaok4nUKCYLCZmYEn5L+DFf+bBGKxCH12H9Vbobq9XB4F3j6lrpmhMG4Kht00j
bPsVcY0KXGJP/FOdxkihhGcKnHeIIxa+VlwPFItZdTxOms22mvReDEihop5Z0VlD
0+byyjEMvTIZFTXfhWFfeGaw8G8Rb+0w0lMKBZCMw9GpAzPeNGm4xj183z0Z2stF
2J9ufjn5grF/Rir7ItoWl2UPECMInxG/glNvm+8CydkRw6/5wNAvhKRgdKEgx6lP
RbbJj0+1XddkaE5s3s/N16TITfnOXGmlImxDr/FWIzbNyfEl84VBVKF2c1Zridrv
vjxVzfUe7fNcYC4yOzVMbtazD6WpnTs/0NNCN9MZdICaJsPfIUwZhVb5BrZsUxOQ
AfbM3tjX9FCxhOeYRBCvZLwVzuOyfkvVo5q0ShylceB6zdD4PrxV6BznNZoNpdM4
UkjqjT4aTv3Tm/jYLh3Xy9I5iaHS8lpaNd0pdQIiiF5/tkwGgN/AQ0iabWtCcYb8
KCgM9UEg0ofkLjLwgDrPbhztpoIhP1YlVNIsevrrECQte7jq+oduyyWLv+VTPAmm
fyuq2Q0kK8Rq1cSTEqSNbEzkVqW/RtCsksD/Yuu7cO1KlCH+W11V8L0ao8z+l0O+
o+opUMwo0AfMDSFAJmNWMNHnBrcJEhfmxQRj3fmlYnLcaFN+lpC45ScTnkGkkR39
g7eYP9cbyEr88w++lmlF6nPFtwmRHq1+NlWFjsi5HgL1fnFvGl331EN6KqXt2u7g
KmkRTR8f97T1y8lBqQ7IlftllMuHjezcjhkFyNS207NSVgTwVsEzgDZZaxQrkQka
tXygoPaamsW8onSL/E+CqVPda2dyaX8m/0z5qWIDm9FzEpvG+hkxN1G2BKvRWAhU
kdZSHK16Ha6o+Sisd+4vgVS34G49eJn7HGyNfCheUWXdeNGS7uQnhw/7jeHjI5XD
ORFJ24TlLxXmX+6DK4G5jpJZpkCbXuMzBb3d18M3l2sXCGNr42f0gETYEtys8nWP
ocPNkSFcRwQFcplFhDczA/5fUS5qDbtgOVeHff4UOALVZ90KwWhPRMVQ0eaJazG2
dClAqUPMxd9lv5qok/SYQC/FutPxBdXmsdlT/rYWfm/nJIrRm9jS92mvEukqQfob
kPRrxtAI1u/iWiAlm6XDZfmBQKqOcs1XaR3X5KwkWyLuIw+TDoR6tB0k2Qaqv9Ol
LIT50IMtIgcslMMJxkCXzw9dKGLMv+MO/eVQKq77vtQFMNtT0ZGWIEE7G+CEXyFN
oI2JN6N7rUbqZBmcB1QPCZx3l8XXdNXenANRzxejfUXqAKG4r1D2llImC5uGaJwJ
kjFildo3bGbhBrnLi5GKct2TnN2p+03NAHjczy2V8YPkHj2gp4QLE7aM5o/cv+H5
cJhtJQFHau6JvNGl7Qf4Kp/9/27/cHOCAc89vxe/D55BFZ39G4+tz+RmalX3LwFT
iFq44zQnN2AtNKTI1YuvAbEYRSGarncH/ZwoirkBIgSVEumu9yVnBsRo8VA2Iw2q
cCva4a6bQf11JHjNKvbPRGXpBEmcd6gs7Eu5jiXHiOOk9UtChLXOuVeH2SCYtB2O
NQ+vgYSMlVkEoT58mIhLRWbizvfcAtr17B2yWX+JEZ7uVEa6mCtfOKuZNwMJkP5S
7cHKffq9xfa0TbtSVU1GA7714TKYSmUAPSMY6AH3P+VSYbYq1dKyANl6Ry+nUIaH
Ha5iozSOkAY3zVm7p7IvR+NyHbFSXslEHkqGSxu+2Nnn9TgBEbTRTQ6IBoykAoLh
KOOYfbzu5iMSX/mtyMOdutUl82Ha87/kw93zD++wHhxkEPOUbWtLD56zRqqnO7xV
ipD/KFDIcEHo+TUUEvPKqmuhFrtDou1F3Z0wD+FuFllrSqDfZe+iOdbvH/Npne76
WFxyNAQ7wa93wogcPd769IMvXXgW3e9MKizWY8nwcrhrttWROZHNziC2cs0QXz+2
nnfgeh+ZEVmuR2dYInKe2Kybim8PzH2Wdt2C52VC2u5dGl8BahLvuOLI2q/rl4th
6tauq7Qr+yzi0c35z60bwTitvASVuoi7dXP93iWsvLQkeyxOQxvHzx4PImoRGTeX
B+CKhp24yKy0W31Tzj4ESfqeF8iVliHRmkpSWPKTvKSsEc7wMW/n6+GgaxhqlOGv
tU7YC02gccsmMeFC8sEYEgYfVfjQsDtSh3aw2TRwGTrfoC6oRSiat8YvVd0RUC8x
gajGNlQm81en72s7sxMpB/o+EsjxiGPeNe2DdLtyw/sR5HfSbi20AeBECClGqnRF
Zw9VxvA0tMv4NOTc2YhIs9BhRcGuw3NAfdHRrtpEAcraUp+98uSg+M/tsALxQL02
kYGCRyYoIf0g5+7DzPO69MK4EG3vfQnUopfgZesOWCP8r7sVXPXYBdi+f6ESBdU0
n/jN/k9kzN5JZrzQc5K5/e3iTINoGPfKDqLq2++k0rq8NgQlpYG3UfaLioNSgiXF
Ka8M2kXw6GAtjzGFwP+uZgF7pWeekRmYRToZ4Jms6ZIMK2t9tq3UwhvGNsln2MN5
0H7lOjWAIx9LWZUgxj7kcXPVv6ETe8f714l7AiPrOmtA6detIrErsmiEopREMV5x
4KPT54+/IYgDl7OK1ZziZRFB7fZrM3AzakzNO1mf3fAuyS1cMJofjRzpcRgLpblz
P3JoWYQ4V1IvTrMnXeJ93Q7NPG/kI/htxDsMrTB7D8fNW/sEsPkGYpoMYF4HnksY
KCWxJSvQeA0k8JwKTY3lQPX4TyxRXwp4xZ1vTojzxKl9twYdAYdYLdTgnDu6SPxN
/wtnHYicpEZeHUAx+KoK2rWEPQPVVae+wL+wCykHwH7asrT01BaeJNZBlN7T6Ua8
iUu41Vy7BSc/5V94bONIPrLbSarX5M0pYmxjvA+46EDl1ur4BcB/yfk3JE6Sia2C
8VM2bvYSSwE4AspABPP3zKFJe3IROCzvmRHVnk0EMIhvRmrrWQFyDhrO4SUOuZ52
nQKdJjeUNT3TecYBPiYmVDNXjJkjdyx2de3sPbukE40/bQjEMgG1p8IlUVHsij6+
6Zzbck1MHNFVJMm1O+/wwduHwC9QnGkgJB3RiDLDNcEMZubsg2t/9HScArkXdQvl
ui6IcLndINqmbJ3Mw/qjZkhNUZuyScWUr6u+T+lPNjQ6WyRdPe9PTC2CH/oTLYgn
ZeFu5qW0l9MbL5qpB0wzgBrz3FSZP5dt0m9Fj5aHrSs4bTooGXfcXWt1mjkz8MHh
OnlcWeG0vYK1W15PlebCWDyMpLdkf1YrDZdeRLtWYpZsaD7DZJXkNciRUPZrZkta
qbDyQ7xmThEQmCDGSagFlPXweAE591UEZ4ao1M6pMIUhrJHfXj5Ym8+Nc8lRjWME
z9PixD7/Frnk9mUC+b69JIuo7QBNG6hgyCf3iRxY6VAtr0eZYgfuBi3rPbWQfthW
w5PaRWuyXuFRtS2elakzIC2I0RtTcfRFUBPA1jcoUFF7/xVU045LNroEQyCSzyVE
PWn63Ny6BjM6q91D7Q+r/C/35fkngg/Ahb3KN+AyccDcc6PD5h4u1EkqReFgJfX9
KgVrChMnLERsl3rJ9CvHDVh27K/O/Z6/NuQcLDX9mDCKjiVsLw1kzTsMO20fvqt+
In8+O+YeIBnL9RxSDJqC/xhQoE/f4mJWCv0fcm+qxrVHEd8i5HixTLlT1jzfXbWI
oVx5SRi7IujiHLyvqjp5ubie/0TW3j01BpPCUOGzWmAthNP01mWuEVvZR3cEsuGD
YRsWpA1Qh9tO+yLKJDHbjwn2vQdJv6P0fyWGlhIpdKD25AjvHnK61vgVIZ8S+yRe
FYDh72MNrnDnIUnuDeKIKX69PN0xXDw0pCCHJ2Dnzw9HqtLERxy42TznFagSTTiv
aH0qCI/znJJatvutBmxYeTrf9gLIjvySd4LV6IYP/9WGtJI/6eTuVFEI8hSzXGRP
5VdeIlPAU8mRGqlE0YCZc5rbgkTqOIkQhDwgbEEwraPpKMiR98HdK48KU50YGIyW
qcPF5Hhk0aZStBXbvzw3Ih6vE0xeoi1GuLMb9LSBn9mx8J81Ts19Fg8WKh/jdvdU
6BDsYqZJ18070EKlMI2uXtBUQm/MfE6E7KChACyzNUWUZ7wVHoWl4/0VqfrAXlHc
sKZx+Vrxj6lks1SHNvtaWLelDW+8UybKDgpCy42WKp4x7siuK/PMQoxxDUe5Hbtg
N4TMEDQHdxQVxrfyZ303Kkmomqo1uvM4OWnXfYfcj2xhPWGXUHpeL+XnpclldzFB
zqOHwFR6ukw6MxjXI76HW7DvON8010Bl31iZOKBbXASc6W2uKmrYk49zlSZ9Gm3i
Vt2OuHXJlGEw5IJ5wl3ObbGFvbIxEVm6OkT7NXXS7FEoxXCwDrj0Y0zN6LtCbsXq
jSa65ZVCjuscxB0VN8FC2v5U5qmFpnKXfElq7U4omyZWVnU8n3ExfdkylV7dNOk+
E0PnUct9UxttmgG88uqs9IMiwLq40lGNLoexXNeR64a2eYT3ZVqPV9MuULAZwx8Q
+HHjk14x50NFyvzOc9V6D+66zjLdmDXPdYGJDiGur7T+kQHYUB1HVwfndZ7Ys3wF
6H13StRugBMuYlON4ppE30THck4h+gSFgTsO/m5zrleuQl1vpxvDMpCkBDrCtfUD
Hnitf6Pw+oLL0BL9vVCKa/7ZdFOdQdXIjXs+iJpKKCLNQtwi6tAnWkvI58VRvYZo
ngyJwKzQ9C4+f5o1yUJrWlqDXWF5kcicQdETO2D73MOHojePl65ouM+Wv9It8D9B
fXvoNpzQ3SGOf5US8adx2KwpmggfpccGFOJ9eH0nbJ8xqxPhol8ExAZNRkeiRlr3
+/abPJskYenOrfSfk3gAIizXLUt0CN4wmW4jdegM/1PDS9ThOhK+LXU8tOvK2apF
qrm0cwBbey5k9sh1sc03he2BR+AUe/iyxNJXBsBxb8ZJEjejQ7gnakdzqrFVm9C+
z17/KmojDjR6S7wcaNE98aKV8LlJQASiWzOR6wS5FX9AmZ6iEIHQSVjzqpDsQINt
hKlHs8WjdOwK7LzRMwtM/ITcmptyytqtcZeaiacN0oUwGKY5RtEqvsTOjNN9bEDO
9r8pJe3nbz3g5gOt5GFl5EeH71d3vSrzz9u70DNT6MArQTcM6TJ/hKY5D7gyahe2
NmKPUwBhVBQZ+xlUL6d8MywyBto7RA7w3uOVjQLZ6R8WE8mt+w9tuQM8+CQ8tZFJ
AaAqQzbOEhMeG0bfEM+L/zbYpsnKjzjq2/0WiOBxYwPZfiAD7jr3bTO2N8LbQC3j
5Q3xLisLZsps1H0VdR7yT3USJKcP/XK9jbR4Mqpw9hs9EOurQsfs1xm9hy6gmx7H
R9jJMdH8z659XOTJGXtr0523OBN2BdeYrDpTfH1CMP3FxmRZtTTSSmzsYI2s5xm3
tb8Na436rj3KSYowl4fecVXHI6BvSV4nrzuDLkHMXkzeoHMxruI/cazbhNTtFDi0
SGH3FriTxW4wsmNwyn/DuTeC6Lwvexd7qexLGCxRrhM2FoXYulTtfHuDUbVNIvlr
s89Pe8hcNSU0v1K4+S8D/S2c69I137nJmQ9vWHbMVQutxHqKeGd8llMEbk5Gae/O
eUrNnW8wUAE9Mn828sIYAKKzH81lc/sVMfFVNShLw0bDqULVPcKmxfBu+auwxc79
lRxrx4yStAFXbltRQeEgjf0uFSu8PfO5AYID4rMkHmLVWJ9pVZJ6FBgYvQawYBJf
yun8ChDymzUpOoruEf8m9YCtBHiqh8lSah5fyU71POaXKnb4ux+hQUF1gQR4fcnT
MXRlITz+j+C3L81bt0nCKlhu/0Xjd4eYTvMyBjp7yfrF2b8/6GYKexFU3fKz4otg
HWsMr6cDwMLapc4zgeluR+MumxLLzPZA+737V6KG0tYp3uFQ9Q4fFGRJx9ibvpBE
deBv029+iNn5AYSo2tKdiS9jhnoy9jZae0OA0kzVdtemcDA+TAMzDBMDJea81UXd
sORg8vAhG/SHs485RLebDGeWQvDNIPx3qsSaEoeLFBjX57tnZfvBSMzcOk0QR9Mk
Rrp9RHKJNVlV1SC4q1oC6Wb6JzqmooMSIjjsnPWyw97Nw4yJ+LjIa2AbjXynY3Ty
/jeiYp/q43eE/ngTy0pXTVSjZgUWi9TdHKuaEj9Xvo0wfhS/JAbUtdZNepUAGQMu
CtBbah1XjwxR2swUmB0Uf//+x5VXnVVDglRQGtUUd4wm9z/DU1IY1Ea6nD3AnJX/
6VFDmB2jofzWrpyav+lEKfubDZDJXYJgCwsJIELyGvwqAp3mAA6IwxwVqIrvGl21
iDHxBzXo3AWyRe3oEHdEQwdbH82glD/0aKyhyOMGoHowOvXeXtaBsv3RqwIAC6nO
7P+9DKa4lZp18i/LqmJDdh8MFqNxDbtYf9qj9wjVuTmRW2OYm0fqlw93jyQZuVi+
Y38zaNuU4dVvh17ML+ktP7ku01P184MX6bEj6Ustnwp6tCQQPMJ58up4AxT78LXU
l3YtWxGOSBei6NP4n0lZm0IUWKLLHmrWh9o2Oomw+1776xliQRiATXCbTV43bDlm
UqYk1PLB31w7RCtELoQ/wevW7/3lF3YDXVw4d8XnDVFu/U7dw7Jg090c1Aju1klr
uYINSlOvWjk9YFg9COBuVdclbEJu0on+TY41b3Hg5b9FQYt8irqQOgDU8saDKK/l
LRjL5X/w1DrrEhLP1sLsBmMiEaq5JkuWZO4T3QN+RKCPpi1VIP19XcMXBBVcHUGw
e/ivy0zlEE/2Q38RGiqjc0ymQb+y1JuTmXgsEwKWYWIdidTev17ffG9J/jwFjEu6
yhHEhvpb6U1FGy6+dc8UpiqjlHl7UFsejQz3bOwtsnEKEERdRScwNXH1qAnhC/sY
8OI689XhNT2nAeJGrDBccFFbPm3adhcvMZNnKpe6oP2ZJ1ydA16GvVforBMxYAKp
LhSM/w7USrrWXLRANNhskMTrm3HBf5ooA8fzFh8MZYGxFzjPGyWRwtTJw6XwLNGW
87h2z54pJC8oUFatEnug+anB1i4wbzQlb3zzXr6aBq4yziordPnx6HSlII6F1wJr
pQxw8gA8Gm6rdnPBtMNZCzW+ughzTdermIGXPze3mEzWCdFIH5MdsIQDl5vFM5AG
uaDRfZ9dUXKOfou9Ay0sVzjZ3706GAoXHcftAVpdDpeUP//LqLTbZAV2uRL0xEme
Lf6b0GLXB0+viA7ZntIPnBxvUcy8XHTYUoqCJJ/u/kTobsraoqAkc3BbWeoCkzUE
sujKYlXjPivykNW2aaFl8BQNrkepYxUS/u5B2U4URhM9Dnv8uLYuauF7t6BaU7Zt
raCz4FupIY2JZyDSgkMFGAQWC326dhfFd5cjKKtRnUHlMpGM9brGBTdqrQv9AqNP
8mTm3bfaCSpSneJSqXls2MjrJurPwJQoQ8wBmlfFbwbh1qfd/XyqfRF0wXl54+/+
DgwVYgJg4ye2nlJUyzZVvFL7FXJlyANs32H9usEsmSJdHI+e5hxnbxfIsTvdLHou
E2Ci5fBIM+14wEzBHEWrVrEAknSfVc+iR3rF7Q2zY7zmju7Cohh+ZBoRitGT5Jvc
Hv6WI0shmuqJdZ3Ba0E0klvKgA+hVcQMJKBLh3MsH5uGSchem65ahzMNWWGTXcf3
A9raifILOYVvXgZk0DyekOfIkRYYBqqVh8P9FCAbFJ4NntPd6Ax/Gwcyt+rVrPJK
XN9TRyRdN1EiD/L04/GQ4CnbKALDS+eKHwQhcM7ejRh7sVqGu9K2Dqc4QakbjQHX
ehPnvKFsvzNod1b+Gd1QVPGilzyFKIzje4CT+SkRChDVKZGiNYgar1drM1iYrYIY
lY5rIR5FD9AEHsSbIWtgiGAbVjEgAa2v9/5xqopAQEMjv4IeRs/ymzy9+GVMrLfE
OV5g6FRNfiEfLQqaqhiHvOjkqjxulIUeDnaN4x49qCmkLKg+wVZwofbSO2EiZZ9r
rp/YFEFEXhWJqeTHQ+PK9MBS++QWrMirhgLq8d8KnqZ83fjliJnH8cByb7UXz1Ln
G4lm+/m0fZ75YRQqGtaRxmBG9Rq7igKxQ7LsKREuf70igWdBTduezJblhqvRDTsn
0BH1AK88lM0aFERH0dqWfr1vO9V1WsgzoMynGZ+fpZJHJwm/ldvo0rUMWP8r9hfd
PhfVUgNWOivolbV4uWsLi1EaQoh5rljXSvjR5YnuD0qjUw4EaMgW/Dm15rd9Z4eS
Tm5417O9CXah4lI+rGCz0VskXZ4/reMMT8zfwm7qulzaECZ5OQBMBevGKGkfsqld
F+R9sMxcQXXO6TEIwWpbttjiUhWSd+1WMVaGkzYiJSjd1ZTrX0scnQtZohFZqkvB
qukFYWEygvn2KQPU2F2ZOQ/IWoAvIGNUPXMC4wAePJ35GXWXSmWuyeUrKJEP+9z1
9dDOX42oPYZv8gt2ERSJz6LrRqB5cFUjT5uR7PFjsz0hiUX07Qmi6DGM3PC7HS0A
gl7uiZS0P6qvDmeYqJbwk6zHB+7FQ4taCUc7MWmSfTZB14pjAr1YK8XdkkPogiGY
cXz1nhYE3HOPij3UJjs03XTqOXMPeP2tLgb9hrupxnEsN/jDS5NBSrSMveE0VJfE
0+Xyl7IZb2rfw7N1t7m1cHfLLyWsUpIDyLTm5jRvuCgAVAY1z9mXJfkBaX2yDqx1
bWl5xy7vAQ/HEpcyGTWRUAENGRZShEVDwjgNqPGeXqMixP4MxI5g4p20wL7vwRjp
53Vnz0NLHs8XNRuREwE4PSYJKgrZV0vTQppBeXOu5QIt2F1nzqdstmksXm9wE+yq
rJBujYcafKo4utcOcXFxoAms4W3aOHlqixLc46nd0ZxetRnzjnyKqsTTtWL9/WXd
/lgsD72aAXWSfy/AVXS6K92bqVQCbjSxYzh/ehK5XS9bugXxUVzZAeeKBmxkghc2
tLZCraq9CCHHpaVoX14btCxgi247qAgDhnZpAz9COOC+008QTHgwCMyVr12rtCTm
R9gHk8p6y9fk9ZElskBaHMfr1VKELfhRqUuKuXadrMPFcNV2fJDrkIOtRuqg5BCi
2X+W3aFGKDFZJncl2p33v1qJcpeauWuB0dlvgNzMd510g/6akxfXUcHznuuFN8YO
b1byORR+fx+Nu8X4hbQ1wqKYiIPGRxkCRIMOSkqx2EnWS8l1YFu9yZnjOvP5sic+
SWMuMTP1pfOxg6icwfgdieIGCFLbmDekQRyVP1h0LA3WVkoLYfDEDh+/fBYnRoRz
ya+Nkcnk1CGw+SRhyWSR+462Tr6yT5SrVoaq97iYRXMOFP8BQfJABUEoDmErdo/M
JssmGiwMzTg/saQumZfigp35U6W/UV8BuzGiXyc4qWxWZzqIW7rIlZ3GFVqrLvqX
k8YKN9yb+E8kfbCz4j03CnMxpm2dx97SMoTclgxUWSg7zy01PZui57fNItbycGLo
yvMuGMEfXZq3F7uU1NcIFRDAM7/3TYqSx7+TOoqXb2N79wCN/eKOv6glg9uvI7uj
fN4FjmxyV9g2cC8SGDczlx8XZr5daRBUBUMSI4Rp5YS08lDOsvyRkiAmR003mFW1
Nf9BUTZ2eRlMqKbZKWp241rdr4bHSlmv4R/60d5VSO2JjWG+1hSyHjg1IaNqXGhR
Qp8l1y/Qbf2KhP4xfsvQCav2uZCmrdodGvBrks5SWOFhL4RT5ZJSWQFOzlqkZQ4c
5N7sfPwHSumOjPnQpIebied1lpCSxV65qfkAYl5YAiz7Xj7LfrfAWYpJXYH7/BYd
7/UmD/L1+1hwK2eOO/Kig3ir5iLoSTwiu5iatk14YMjhMAepn+yPHbOLTbDxDgTE
72iM0A0BJR5XoKsekzGuRWfeR1BkMAUxoEbmwBBKll7+F4sr7JQVe7UOgA97V38k
urciKu1PPPwPF656Lc6OKn6hRp7w2r1Q4YvDYRwHiKEWqPnOGP2mE5s47W0SKNAV
Nnht4mi2C2LjTEtP+7myG2pOI7V0/G19bmNY4y+4Dgp5x1pKtuTtIA2e5sM8qm+a
acoxzNE0gt6W3dN5Y9bWVCzJQ1QcfSj0uaAc3MubinaPZC8UfEFHkdfAIxk0m1nG
cl6PGBB9tBmlG9RKKvks9Woi5yBcTWmCFh3BVynVArdUbcyGBDpH9zssr92bGDPu
/KTL6gPHoT4EDMt47nUzIJuWT2CGkfmj4ERnFATqvHl7rM77xRTYhzvzu8uzglmQ
khATEh7u3MSeayW06NmniRDyL7b6MbfKloFV8oqJY8jDjvgqeAAol8fVPcJwg5Co
9lJ9pSnXhRYjtCygAsFDzhy90AqS0Fy1ucfxB/odQ2O1kUpof+niPujY6mPDnWOm
k1CUWX9gTuONskDNMezPJ17DtyFRFsjguoifFaBkDtAuVG9jJWsGJ5ZdNtr+2JML
UidRYz7xAo0j+KzBWES5Kvj7gv3q/6Ai0ntRGJBvNFZqy1xs1KvX4xJE7ICPBB5j
6aqeT2DzvkUQ7bfIzX6pcZGqTtyYvzOatTSlV9jhvQHHVQnvSXmn2haxVvoh7XuU
LQ0eDndztN1R9uNR9NnHbrHBulY1dl2MSfMWFze4UnZl2163FP+P24BXXehFKwyL
/1FznkVkr3swBNPxOe06tt/Xp22JcVomxIaWXashLKLDEhc38ENZYJV59GYywQ6/
IBl/PWJCPV7la5fl4wftBtC3VHWKfjjPf4qOwJEBFBHxiQVtE3jUCRtiB4qEfIx4
FMlwoTKGruSd8TE3WmGxUJW2gWzwozGnQWnvccQuunf9ULJ6lr0d54hNV0oR2EXT
AoTnvTezjfgjyxtX5InHS/E/uJKIqSpr44Bg2mwwAT1KCySrLE7rT52O74FpZUin
LrZqqhdeg8YHvBuBRXhMF2AaUluUY4dXPMbt21Z6i/hpRZBkLxEbX1QFnsVQ2wmS
aLdp7qeCLlvAb3yetNJi5jfUonHS085Y7GiY337CAjrkJlIpigCuUHcPosuH+8Xm
qnnNZNj9mwuymX8QUz6E4N67B0Wrn9ucIltIopeeewo1J6A3LwO3gefPZbMwXFa/
lwCUxTO0YzhNibRsplYLHSmsXl4VIojLs2WW616izxf8rvtRFMlHhyOsNcVJpfW0
HAT8i8haxqcM+MG7Il6bFHnLwOi/US+f3cLG7mc1TWH0Bh6Hw4nXuepui4BaPJqX
mdYItHJ4RjYvdEIS/qXeRZh5VEgcNERlMRaBhlRVdhH+2vLbgZISpT/MPyTfCpeQ
cxuVlMjbNaLMR4QDKjtgJ3wXrOT7wOQAfSQRnnUNV8xl/DEywgu68AdRoIRTO77k
zceeDNzSbQISIizJG0YRuWSgG2prRwLMbd3oj3WlarFaeCVyDOplzBLkNyz/vZbT
Fx1XHy8Dzm95uM3AGnCT+KpOyhV3A4uZJ3krttIVzoVkXTZwqtDORaC9H+gB4cb8
RaQLASBrgi2KmaNyQHzCMrKSghfKQOgpyschZdz4cqaYN9Lk/VN+1Lj7L5bm7d4Y
fYOiXbdV9kx9UbmtNeS8d0QuQXnNchmZHS04JWXCCFMGU3h5dhnaG0eOaT8+/tFZ
7VmPkcfflwIYb35z/iDg+RbeJxZUNMXMC7imMbcSooGKK+nSgEM897gfDqUMp2lA
74LJtwWOuRhCEatxg783lOMi0RjHbjzJr970qYvruq2PVBWWZoT/N05sdy+oitjd
/06wE6793mxJboHCnbXKN2aAABY+xuq4KZOCC04bEa68JTiGKj2qFFc5CbDjno0l
kJ8FR08nGy7T5/UVbbZDM58U/7ZUneMLfEUv1ODzYcPou3UPMh5PkJCqVkeFxt09
H5zf/4nv2N9BTCqdlZlFabjhTR11ygmhGYzjNx7OWn70uiXj49bm+pDjlNP08zTt
oHgYcubQeYe5UhUa6Seboz2vW9N8XIcamDCB0uw6Xw0BJ92cKT3HCvo+y+GFTWn5
NO0BHGuwY/oBfX8Yg3DS5NkdzyZehHKvgw+21NrA1QUNlkiRNyUVMjRCynrBfh2A
Wtml7cTNlIgWmP/Cu/Q8s0MLvbx7wgwvZENxiZvKuVCm3gOtxrIRAHU0LmdJT3+s
XWT14p6uSZsMtBpKJwHhZ9IIonQHaPwAyKhNU8nxEVvy8MTLBX6/Rl8EGGHuNs6M
9wUcychqBahfUig3M04TlqTxi+q+ySxTO8RK5amlxT2Jq4LUm2MgiqmH4iZsfel1
RjbeKc0eg6rn94tLC4jLEEzayX3yOFL92uNDtQSNoSh90si9i8dgB1V56dta0zrK
4znOPOYLKYK0cKpvpPu4hOpXjzLk4zqcmqZsesDpYYb9kSpxKwD0r1eDCcw5elr1
C3OU3LCY7iZMXHm37jspltOqk7VMpYN5Qz+btbARI3nFGQJyhtP7Jw7U/kgnbjza
BiRsMEGt7x4tZ5+4gzLLoMi2hNDfzw0vzVIz/NEGoHTmO90vjiXch/mn1DlQvb5N
uYlgDS6z3QVyWziOW+H7CeCyVtPEW4EctpH/hocjwhgWElmXcm6oSrJomgOdiDtz
CHV2ZYP9mB5Vjk7ZKWVrohhF5xib+QyttvRdJRlgFGv41DTqJg8+UryVVhklKYcP
ZjkRj03KEPCIxBvzYRfdfS0fa22ei/1nvsj87jnqVELnJb1TmJ4Pu1y0bzoZPVOn
DOmytLpzX5My7pERy5OciQbSpMdtOErionRwxz5zijV1bvcbjClsIv73TBc1XyMm
/Pe6ySve8Gyh+CafLK85yuRuc5x0QalollxC8I4YcP8w/fXBx4YhCMZwLAK3OOIQ
Q9FqT1FHsiulGGAJt0Ykan2VzXbkiGy8zwMhNCUYGfHyadDzKnbFIVNkUJmdb6wN
ye85hXQ0vZQyY/U386M/SC92JpRwD905mKlVJIJPNrnxSRIAl0HLpZ1W3IcLrqI8
HqGfKsRd6H3z3wGzgO39ebrvgfgfu1o5WvWzGjmt+vHRfiQOAkaqXN0FiR1IezIJ
dbEHJeAh6nO3SUeC9qaaEmZ5dIosC0JhMjqnANa4NSfb56iYwRW8kGh4qdYT2yx0
LI0BALhYRIKeOaYTAThG/5PUo4p/fPWQNJ8/A/YfR6KhJVxeZ/wUqrLgU+NI5zYk
1QAgy+gP+dbwXiVX8RvZ6S1+eQKT/Qpl1jMufl2I1QtR6Y7gaaZARKXqRNsnxciZ
OZhN4Hzw8q7D92S4sKnVLHQTbI1cRvPCXnKXpGX589hg8GsfxKXcHmkeJZwqv6Ds
QFf0PUG3WmL5W/dHBZVdtWFHg4BYHkdLC2xORJZDovwdRZjc61KQtAjTvFv9AsPg
S0Si8mzzYv9qCMr8Cn+z4fPidLwN6ZeQzmVXLeOPRhrBsNbWKSfz1oD0e4Dmevu4
Qt+fJRQycJqKX0MNeWiQ6gPcRfj1xcPOSarCnOJMsecrFOCmhEu24PfhSx5Xd78Q
pH75qSFSK1i3/VE8KKBru87t1DmnezudpwkgchlxU4yAPluYfDwdcsu6O8YnhIzm
kmirfgsISzW3bhZZA73dVFm7FbojAXz9T0t8pCHf0VshdNycEpvz/i1GPhOaI8+C
V8/IUO+xjCJY9zBxM2OsIN+so+34R8LT0Nc9Gj5j3nLQ1rOp0bTR09XANPUpRqHG
Ao6rIEnj5P93fR0muqLbNIhD9Zqz21PcdXuA03oVoLy2ucyivC2VnC4CLLNe/zi8
KHhY7T3dfrO8EXdfPABhnF29MoVqdPOcWGijcrF+VBhhy5tfjSGJhqB4YwRaHacM
MuWfBja3+8sjWerbfo9C3f6WYo7DlizFDkTa+UShP+SfVVjIpg1bt4123ifEB0+r
hpXS/Q51K/UITdxcb5IVxLapF58Hij+zFX1nm0rvnw9acF654LccYCR1ydOQB4NH
/Pzsvqhb/+6t6pI27ZiA67N9WFrmiqCiVus6Q9jNYZfGHJvhS2LccbaXrbXJyK1f
erGLCOjPk1i27OeHZ8bWB+OfEVEFHExFVqhHHb0+AsZjc60IJT9vpEIh0AxerTO6
gWD8V453QxNc0bByVOpOeZKyqwGn8r1/CYnI82LleLkXMwT6bNer/sUYt15PmDuo
aARAn8URb7pryS0F2kmU8F8T6Dxau1K5Osg+jTurULRWRkimNmNJLRRngmRMB6Y2
qt7QiD5tdRbArcY2zCytps/BDBJnlWKyzbGRuWDl8xdXh+2KndHztK8dyMY+iDoc
q6MIMM9LvCJhwdlYIa/9olL1CnZH6QbN7iNorHBkth3ksRYSbmmTjST31NV7AXGQ
G7y9w3JH7zBJ+rOoNhDYNPJNXqgncfT3fxHPfui3aF9t2b/L2vuYIKz1QPVLqXDp
JGd4ZQAgfEjdKAIhG+861ePV6MUMJl7A11p9UpJaM/HSZx7fo33y7vkwSRItyT/S
OnAt1g9R6Vebq7ydOwbf4XQASUGHPtBN/BdFg9ThGIJn19huF5ymzfvSIPUzbTp9
embruuxOJnscjczU9iQ/H1SeDKkDWHc7yc6XtitWbxoiF0AOcCwNa70xF+TFlEG+
pqQggS3UqgBVIeLdbGyl5qG3xj7C1/hN73rw3804XYDZbNEr2xR1+r+oi37vTV/t
RUAwch/RiI7NYHwhavC9ZHH386LTj2cJ1CslGE+ZjgDvVvMnjg+eAnqwBm2Kl4ur
vH5yUN0uJjxxYN3ZevD60ktvDO3tp7/YAvdnbeL3tQiUQypO/OTV5WDj4CLdY3eJ
407q7qZ0EM5xWrOLCyPeUaQpmOIoRSid6bTbZ2biiD2Su1p0q0VK7VQWWm3km4iV
H0Vdv6jP5Z1ZI6RRVN2uupYiydIXYk9vs4S5fF7r09OTs4+b57WB0mRyr0kp0F3s
2Eg7I64CpRbDNru3/7TG99nqLb5t06G5WBxE/g1SuyTb4n4NvDbV0NGVkfKBvFrT
BxqktBHdcAQrcf/UlRnQ6xLUFt1hToo+mvWCV9SdkO8oGWOmtUYjpYU5xNk84Td1
W4FfdOFG2RxjYqsQFiSMzXoJJK63sZp+rEsVNk5mO/pfk8Wiv/hLHutp6JMhJ/g1
rkwB+j1Mf76G40/sby7ieQ07v23Zav+ZBIRCbE/fbE9ezBk3wqrsQ9XUAMiDS5vf
CtJCpDjZ0GSx7jSmx22zzJhzBWbYjrlq+aaoNJxHcnFjMajCWPZcVBIWJahcb0Uy
KURxX/xt8U7DIckfvyhiPgNe7zUqNfHnq6vRrdn1COvMsUrezCXfuXPfd1Vqrns+
Hw8hgyRqDGa+m/VacmoN21Q2UMJ3ATI0jbGtPsjzxSKSUZ58W65sbEcKOrUZdS8j
WaypRpEApH1CS+xYfrG5nZeSweA7ZsTbhgGs4YL82WZHPn8RDs/zPU7Q9EaDYn/4
oNH+UOIuKfZ+UaCdJOrl+hliqB60+RJD/pkLb34aMuC8f25xGFonHKUP2LkvvAAi
gAwraY6ENwh5hlLIXNtQOp+p2npwDOvUwHWdXq0uhdF2FeU8Gf5P3zTtkvdeSi0k
Em5fXNYgaQVCLbkPlHu+QchuGepk8ZaS5H7/SWk9KBgU/cxsch+yIwNxgPmX9ldY
PCTvbAD9/K/couu17WtNv2CqQu4UMYTTzXgYXgoplhrj71GvvVxAVznZeZD1G5L1
crAZw+TH58q2yIocdrh0XC+EOfwI/Fxpo1OVn/i05G/fryT0Xq1nUetFE0QQ/k8r
s+ANxBScaQ3pSLSFoAUzQKk1fxMTR3hhoOVxXgoHLiPn5oU6i8dePN284VWxPg26
B/dClnd7a2gsKlNC70Mit3v0KQQxGqoMtUw81gQ/9xjw19Ba5Sg/RRedP2WhyBT8
zPmD3HbUqMkGEI0UZZeVv+/puQ8ML+ENyO0N1+vacog8waOyemaNFe4qjruSe8oW
9hahNUQWdxFarptvifUIzqJwBVYkvHlMNDTpJZ94np8Hf+qRf2wJlzxnfh5xJpob
oT15CqFouy0QN/D+w9w9NW+lVyGXm3mA41Uqw2aK+1TIgjzol2uN2DyyMp6bEDE2
MVfvcEiTKrbkeE7d44uX2zLgIy6tYwXACkC4YhLLrWfocvTy7hyZwEGriV5dXs8O
Dnqos2hOVBoIFgMQZv5LTPBKs3R6JcmY2c3yMwtE4g1/fZitbVP6LJ9PYSB+YGnZ
N5dpWR9bUY0TIqSR4Wjg1o2YLR5/ZMyBY6ectMPzYLgcf3bwXDVxPLVWpnFW3Dvq
Q6hneq1mb8OQgXANQ05iov+3HRXnv+xUzEW8nf+563Lpm8urYKqWAdZgdSUsFayq
7LyCP79bVaBwTxNKB4xtGt5qcS5O6Wtmtqo08fi/U4VXesEI5/EPWv8I4b+q27u3
ZnD5mArusQBWnpf61DZLJVjCTN5WXzryCRVRKQ/2bFPbzdGaEIlU9dsCnYkbfH7c
6rLUzhWmu/N7RKrKXkid7URottQ62y52Sa+d+Fz4ZSAehbGKg9vj+0ufQxoLRJjk
OBnWeThuuV2PWnFXAHNzQqiS+WugWyjN8e4fLtlQm2ZKL5zcTU21PRsNCEkprt7W
8ZZ/eMHuS5UYKMqkZAp7Z8NdPM+cRhQJEIFMOGV8SF5Ijj6o3LG6BDm9sssj1IZ/
dU8GURh8y/YiB4978MgZ6kBx7RUE1PvTiJLFVDI30r0pWGNdPoW2QX9tQLCzsUSx
pqeYCXKmuvRXpgcXd+V9ZPQUjY9e0XZompAx0Xaa3V5M7+HXXJWj3vIdLnri5kgf
B0e1oF5meF0aIFxd5KFuKnrJCB9K6YEIYqrEJfDOyZyFzSvRerJ+xWVzODlMIEMj
slT6cxSbbXJOdCH1z6Yg6hxW5V7RN5k/MUXcZdP6upVNHELpbUZz0990JS9UeL4i
VHdlXXL0+ZHD7QmEV6CfjXRpoPFBXA/bZ9yWnG6WAVRgwhbvfKMZsVpEb7fx8xZ+
NwjlMXGZ9+vBIx7ubKuL9I5A888o66hAkAkL7PES/q6LM+dB0va+OwU93mc4djOX
8y8wJtUAqxJ/Vep+j4SIKDN3rHjxETq6NsbY5vTpk4KhfpzfQHPSWskTcj0bMF2I
3o+t15KJMmPbtK+zsXvyzh1VXEdIiRUCi9DgyVLojj8aVTbFog/gGKPqGZwADCKc
VQ4b5tY8nvuvuamAanmZA+UVUkC8xEAmJZAl0AX3aql6qFSoLhkpJiWVrYKNOJeA
CTgtY8YBhg2Kmfc3EdrRibfWD1C5LpDS8JLa3wv+G4RJ3WKWCJKiLcQb9SwCCTfd
gSVQcbMkB/3AHH8L29hQRk8tYpbXoneKzFs+PBh3UeDVE2nZdIhLRmSY+HEQHQz6
GWvN37cRJffXj7NUsFpQGEwU6nZEB9u2pZ1Tsrv/uGh37S6wNsEeQ+F1etLbYa1j
p7wyZTU1Q5SNpC4MvlmcKR7V7i1RkQwUnCX7jtE3tJGmom0IVwc8e+0vfZXwfS7O
Y34tmTxhhjk1y1Btmtwzuyra+QLHefaZ8Lby4eGT5AwCoMPmTHNZRJLw1sFsSeCY
Lcwx0CyIYnT8koYGRIW/ts4Ffljf0kEg1YR42nnkdtm2c90zkiw95AuU4UJY+7hx
5YEy0NGfYWXh/A/U1l1t7Le0RQ4oEDdC11vBVf7gUQEKw3V2TeTDsRWiALijOSgR
gexUuXTCbfe3EemBBPUqcumR1Noug/dlPUrqkxYe0gdVrCF4KrAM1ojLLNyT2X30
j8xeexjrbtv0hNRz65r241he6yifFum/9WPZpDaxXJoQ92OZPJxAcSV6pzgx4990
6ftUxu0Ft+MNkYca4xMkfSDv6MfF8HH4JDZaqVrrLv8DlNDDugjdHpHk0NGo2nue
/xgPAjGA9d1pTAO6vDdZcFUDsIQVIHEZUt4IQvLoRacXGi9+r9GeYozS9cMNl8x9
mL2wYyS08hRHrXVGcxfMLswcQwvPn6Ncq00L7azItags/9y+uzhogziPcvympUQI
kHaFCQ7E/NIXC8DWwY3Tp/DZ7C6cyDArYVRso5E96Ia+xl9Eu+bEfmzOdLWg6eLS
anvTMSIBozqjt43/4K4WzH80SC9CXjAEC3SkkczjRNoqmMoIM7nKigYz7tuOpSkA
4CqSqqsA3gi5fBglccxUd0ZPtjP/2zROTyhauJHAuvI0ZOu5fmzPIa9oNJgVBud0
6Wxhc/wEM5sXopDr/uy4y7sYUST93O05IepzPl+YVaFcqxBOYzjbjbq3vGyINqmU
hglHrq1lGnFKc4WA+ntQ44J/ZIsw8lEhFWYeSnF3P7TewTovtDsp4s2C3LsIi/7N
6Lc3XI/276peu4W/tJRBNpSjXsB84OGPrpy9rjf775QpFVVwmwfBT81kxWocqNpi
NWUuHw+Y4fCDFlrBgfqUSRTbWlYj2G/jeOknlJTTqorheRuOoSMJRaMWWiA4QKAR
VFqF2v1fHCMR2uhiK2eyQZngTSP08Xzo0xMZYcZwGfdzvbto8xLo51fMlxGGncKy
ot8mgKHZkRjnKWZQgr6TMZHaO1Keax4Gfl4qN6n1vT63dmviS04OT6isbiwpJE9v
z0lnofMVvJIb8nLXpy9iQxt3Q/ldGPrYwz6TNVTT7mElEWzgxzjuGpNftrKd8T8m
446u/kObaWpG8mECleigWzMe++3sZ3EXjZGwPu9Nml/nvdDc2/OM1enkXR2e5FVT
10cLbVGcmO2yq0iXiuPHeZTdIBUpkNOOc8DVDbrfKrf9LsS66Bi84o7n8D8tJjbm
uPqQv5zg9jd4+YwIRlAzib4+d+X5iY58XfZVSoW4UHWxnSy4tys7Bpkd1wJ6vbmL
xwP9+yQBnW3ybLsDKIZhLifCjVe6I+TyaoxRVkIKyCHCGe8Ay+/sZ9qmAfzqq5dG
WpFAt1uuAnN+kHaFD+FCrfp+KXd/l7BKLJllpwm1Kh4oSuPsbOKQ+praG27b8JIv
Y9gi0/2O3chAYg9aDs7GsfYxcgGt6RJODWTNpRva4gu5TRKwJ1lGK760ZzL40SY1
knuqCim6DqXkJNVSS1iQEjLy+KJA7s23hchnkNEYqG5zjxmK6jsJFFtNdfq7QvkH
/lYgjsXJK9zaKidsSji3xdp4OHgmarSgWjhSQaVGcKrheheG6CKHsDBT4vM4/LiF
Tnq202HzhlD4UdiNvhvLA+als+4Ivq91QlgIqaGAgfCq05jq6DPNmXDP1dGY4LdK
XzCN/HfoPnQC+wBjpgAb4d/F/57Mrg+irXJh11TRg/VsOiszMsHW8i3zBM/jmSby
SCSKCkZ7aZYNbjZRg2paeSUv3Pr6iVNejVRfOL4xEOtzqriXBzl8u5wpDFvslyvl
rY7jvvaJMTZLgcwLWfR18IN/8wf1q+KolG9fFeBW2d4kcgVrbNtLKGMEcH88/XiJ
javAgKDrCENzd8Y3bbUWCp1zM+RuAVx2BspknZRr2UI8ntgd9ZSd2Jl3Ent0kyt2
llm3SfO9R7e4a+P3IFicz/i6U3hDHPBgX1cx4sbBnSPzj4CdjYvmVTNF3cQ0joiq
IFJ9SsxISlAtdcRaTfojeuXuFKZ4JcCgVSfTUrFuEsGfhSHM2NgdNvPN2mFFIiUS
QgSdLR69cLeaIc1EAKF4RSjXAPp3M2nHxynO+RlcAbd322ZXuj1DYE5TIzoe5Uq0
S45Sdk9i64xHodTkjtInIzzFTCPxQzMuGj40e7oIAEBFe5JOXEOtc0ZG6dDAnL8J
+7F3vn/LG04qn5Xx2TLXHkuJO+qbxwhyX7O574XNICBh7VAtCgHY3QMmJEUp0Dm5
CHx/mNGjaMKw4y/6Eh6NN0X0roX5hI/DBytCeVaLWmqQuwHlgYpb9Z8zxHmjQ5SP
3tkblOtDsfub7DOajkgnwy6VOiDkIWbak2Nr6PMLanJ4P7+yQ61Z3G7p3dF0mYMG
HrVO2hkzXhcJxKDIuu7Y+gRO2DdcANiU1pGCwrFaBr3xBHDdPTRExhvNb/gwO9s+
4xeJU4A7Iau68JDX2QUXEkizWN4lhN0AZ1wXSNJ8hJ9A1iFsqDsSciQls2LZAQCU
N5F8La9j+LJXNHkQqAnRJxcwhaIIGzF/+mbmwnStKFnr5AKaiuvgXKcQi4sUpx3M
cGtxhVswUfh/KBOsU+yGsCFdx2ACq/QjEgb2qb9Fiam/J0fPlaOMEJFjwhEbbfa9
9G2kLZmjRQ1CFRtHkJ3fpWNiross2AON8P6lUve2OnfbbP5we1qiY6vm+A3IAubv
d4y50CX5EuXw7htu7PMTj9nQ46en81PJ+WVM25hnCYD5HDtDEn6eCBLyB0VryHBx
8aGwikj6giJQ+ADvCC5Ev2OD0sd1XG+n599myYv4XHyNjhT3e7Hh4UEns3m6OABD
UViYjBnE2ziYt6vV1q9NTc4kiOk8c1gqcVYMB/sg43LXJplExycCHGqYya3QC0zE
i3Q4Y12DnkFE1E4xczFJDwHM/R6AWHLAvoGn2NKsjAhP+s1f7u2RYBO8e/MXv4FV
T1bb7mL8Dz8XeRyecp/qxFLBR3HTUrQva2enW+yfqvXQ8gnfMeMTlZvSBR9OPhU5
J0liVoyVMyO7UnczMaP/Z6Mnp0BFOsRxop3Y5y6jhl3PfaXRHo9fmuMagks2PCay
f9VQM9r2FAWdwk7QoY4cDz4t67C9G1MpZSls/Zyfy8R8rvzkoFU87Sr4/2+63Txa
aKG9kUIMIZlcFJ/ine5M7XcyUsG/h1YF8UJ0ts8l4pC4aq7xvYaUn7iAf4ONQWLO
BoOQzvMCnFv8NZJRFeO3FRl1f5/Oq3Qye5ynpZ2MvhzatBjWqYeJpb+fdHvVF1ea
V3YJ3xwgGeWAJ2nO0SGfodOly5GJ9+uhA8sj57oyelOdcwVar8VUX0GLqv/aPLOh
gZOc79SmiUFXMByElFd/MfNx4eFWm5//z09Y6S1k41SsW8UMYnjt4WoZNlZeZUDS
JRaYmSfGewwru7W7opvzKl0gPqn8SQdhl7frjkvXydzbUxpOICo1dMcyPEMwO/zI
ACF1t4Jm7ZzqpjnpU/WpQKQevDaobbFQYGWNV63fIkOZ2S8EG6VIboGpyVGT/5XV
x2d9mpDtQP4TlMgrT+aBtWhBRYq9A102brokpFyCm0lH8wCXEEy7FrJUBiyuaru8
ayltJcAPXI/TwSR1Jue1SJxR5H23J9wvox3xOGyFnhjNZS9LjIFQ3NcTEnt3HoZO
rcZbx/zuOK3djdK44jB/StnID8DVbfyj74vLrt7YrQtD5xAzRhqRN8xHs5y3+eVZ
uu4PbVcNrZS5SP4WzWEmZFCYKydrrS+UCBdRx1erTHCJcH+Xb95tOJopf7lBHR/p
TJVJVGScecqQ8AEGPADJLmutqZAPnJunTFIaFudTsteOEAQjnz7Oi/0JER3mmIUx
zq9VbeQyGmsI5vRoyBvK3Wvvf8sU/WonVKupWP0JQ+adLFqqh53fHr4HNy+1iPqR
G16ctOTAStO4TYkFjhP0GeF4eXkcdWhMuHVci2mwRm40jGAYpICelnO/8wPaEiRG
UAYGFTKI8s2gAW1kmKdg4zizMvZs9VKXFbbxPqrcj+mXatIrRenq4+b02bqzoGP1
adcT0fD3Dee/CsnIS6zD+inexujxhW6QC5NtHWvLP3Br6n5mc25vKDI7ABc3Vm0D
B7EuUkwAaNOjb7Oy3fXgXpne01v/DvzGYNgfoTzDWZJ7nc4iUBByJisNFoN4xT3R
X3f7Grdkkjyi77t0D5z3m24hituoJl4MrJlXepLFakeu3zcGYgt+iVZ7noQB3grC
h05IDIuKrqhg7EGax00bKP4SKQvtkKhyqstpRBRCYFOc3bP4BDThhR3uzSMexEGA
60YEGy05L97BQ8oVjGkKlnuC7oHvRmnpypTYll6BV3NeUIKzUon3CxNPtZbq3qqF
l6oaoTbZ0bww/f2v+21x7pGwQcn9mxehDekcAUztaBQZX2ieLyG9XmaKjSGn61Ud
iYOR6inVTADKY35bkcPYwuJh4Z7Ep5etdD6BtqYUfowaSilM6gDotPUNONeSfSz6
gEI531JS150FaQrWGbHs9W865FRpFj0y+Xx1EayEMslKtcZGDSMRTdAFpmHkCkvN
tg10AQHmJO2Ezq1xppUX2cBzryNAHZYb7AdrS8egLpKDGgxSvWyAxf7g4EyrNmtZ
3yVGMiE4hHELY5a3EgZkqnD+tRoUqtTT9pfV0zQ00CImuysTR50oT18yWg0M53qu
59/L8IKruDMh/f3/NTlUC5VN5tg4y4bbLhuSS1WrPK5tZjrWOAGvlAbf5DKjdgYX
HjWR85LsL/XfLs7ot00foV9tXSrivOMcJ+gI8JMJoXFZnc3H9IgEWlWYqmR4eNqH
jQGNn1+oK6vnKmByBq6IOuU1gvdwdth77qzm5ZqgGwGDroUEVFG3dZ/D0p9AFk81
pLPGgJJUAhUGQKRQ7RAyc3KghwIOr7UfTy48ZFv6tM+2JHiArvp+/rkPxXvmTbUe
aZ9sWTjiHWUkYCt8K5QxSicVmac32lSHH9uF02OeZ3wlROhL5VpCPRQA34MDBoLR
ZFaLoKnS0qGd+Z95L3miOPAuSUEXRPjkaW+vjj2f1l910/dvxWT0tvxWfaGuz/jG
kqBr+XAbScI+mvhV3VzGIDHl1LVDdAl+/u4k/tNyFKo2ZCaHMNomAPkdB0onVNbN
1YbnxSzfNnF6SjZnnjiPbss8HOiqbwIX+gC/Gv61bVayia/K0Fv5btvMdQ7dJ4PN
Ta9W3gUBENpoT0aZYJ1OvowarzSxzU2x9Jfva+dl4XkJcj1C17d28yhcKeJE5BIC
J6lcSdHrUuA4Sfd/IAtvRUTmiHfj8IOvXZPBFZOSOtSwWiy8y4ZdkeS11dC811vG
LiEXHFAbMSrlu5oVi2hRZcXt42SxoiN4kzQnC0aXa7d5/zqcT8qcOm48DBPN51UB
iTLAimHTJ2iRbJ1OqZJsyO9K7YF+JVsU+3/oqbuvEfOH9ieB2Ijc+J23GIggAIcM
114kLBp7u2OlI1Hg0lA54/Kg3wOGdZgJr29Nq87hXFqLj31qpfaaBKN06Vu2rMh4
GNp27Pm5uKhwhmk3imKdexF8n7jPj4FaSdJdLRTdD/AnLjHwDMkKh6UoWUNJYy37
tVs9ZKPsWnPvU1ul6F4PxgBTnjr5vXUqhbRStWQMMnvoBo+lT3D9XTDc0rc/YfLf
lvlSiT7zjXLDVBsdEVoAvsYEo/HdyRF9fPMZp2ESDztGoaIuYlyjv7tngfUzcF5B
nLYxn8joPyce097meA7r7AFXUYSlDkSbifJm8QVfM7U8ACvONf0daWZuNnHDh9Ab
i6HV2AaVNMUSlxFXMjYxS+zJtpwlPwc3+k9fYjabtX6ItTeC03uAUwRx6UHDfPm9
9gaBYw1P0yZrKF3mSQSuylqGgpLCZN5Tt7KQ0j+qYU+lAHP/clHSBs8aYQGvxe4+
ruKf/5LP9m47vt1AMTPTEslojxNRtrAsxEEvA4aITMeVWT4DmFUpHAM6yRWVKtQp
8Ejf7VnJ3hXujNnMXUiMr0eQHAksUIt9FhOtQKPRnTB00dUlsPOTUmhRA/Z9Mb7j
FLIi68hXhgtHSVNLEVDxZtZWdjHlqkXD0EJAm6ql8zvJLrtVGDUE/tnf5z70unZq
vnchPyllWVcEWoC9rWy0hDKBcSG/iHexTo4HuD8/0s9QCQb2v5eM86M6Yo4HV73d
WXhAU+NKt/5v09Uv2EOTjhD9UB20JoQo7eg3PbhmxCSl1fg0E9WGL+efn4fW/VPB
+PnX7JdlDSHCJZJjIf/XbW+IwTLqZsoh831YRm39ZWPltp2n8ze4npDmtS4yNlDq
62PYeKqvsg5hxvChrwHAoNkulNFxH14RzaAPmkpZdX7c5y+qE2NlfF8Xiw3Q2IPG
G0hsRqCPUgJR9fWz2yLluOO0hFvNuOOAIoDFVbpp4ypx1RfgBzEScCjNTooPd/vl
0V2PXmxZ/kdRJM/ixnDpqz92lgqwEDQUNiwpoXN2uh4bw/4KwD3Ug4meWm3ywSMP
0rIjeEf9nc1HRBD2go+YKCPYweOWobhlDzVqhwSFQ8eEl+5YPtys4gMYaVM/pgDb
XqgHTH5RJmFftQND6UsWBZ5Tjs7rwrctM8Sz3ryJ0SXjcb/igJ18x5vX7lbO53lo
xM7veTv/qtqIOYzrOG0SiQyiuX/Vez8y09yinXfFD+Blej8werQRmda3VhTnPsIx
bcXqpOHU7NeF5SnLuYR1AhsCpyVcrfBAsGERWzwJZIODl8IjYTtdBz710Dia05zj
BMOmE1ms3ZFTcNLkVnzvlg/756gaWURN/Ma0KUneYTerW55FWBQ/LAFRL9hKjXGW
xFxzmOlSgL2acLvOv8lCenORqMly33mRtxPlivLymvd5FbhUXPf4TCybYK+B9BxH
hovbbicn97f/vm+1NAL4T2OADZjoOTdh6ZvyOOryqsmbrfXUgYW7fmfnqB9d/jOS
hqNOEPHvP8R9Y1K/Rk2hq3TVWm732W7qLXmMu1Z58INQ2KW6b7C/HfWJ7vi9M4BS
3YxoiyfCjpmIKjPut8TPNo+vPR88rw2jK6w7nnKLEGBWk7nmLjyEHoV/rUVsiRn2
aUmY1wKndk5wexSNAErvlWFVN2YCcEFHBBMKwHOjP1GiAp/2ytWEst8yVd14kNfv
/NbiSryRsV32q33/jDwFkycrjgcPG0x6Mf4MfjvC9V/XMEd3y98dJ/61EvagzCwu
dMxu41To6lDiDXR6qA+HxIpqQ9DxQRYh9/gKDW74Ci65AV7QiOCfp4TGLLirUkHr
NiaqsjT1QRZ93aO2tGAaLWTkGn2ecsx6Kv47j2Gw6mkyNoY1XRBBuOQ1LIe6UEsT
jam6LvXd325bPIlVoKFQe8QBVo0GdSUtb3K26Y4UfmagZa2CEqrTm93fsi4+uHmP
dhjMawkZW2fqZW2KyXUcA3UN3tVew+Y6GhrHpe4007qSDVNecVyMehLTuuFRBO+h
ZagWJB55w9TXqtN4w8unP7t/3VvnS3PmVjJqOoAYx9ubyR1UsVscz/aCDLQqH6kG
3dXHY+nKDfUu2oj95k/tzpS84ZujQU4A0G8g8Mfp+yq5lBJU+PeemOXcaD7usSCS
AzmJ/Ua2E16JoiYi2x9NhVjNfWhrzl6Ku7ofsKA9CxLyu4gtAixkVz0J3BRgPNH9
LwbM/XkNzGoBGOMe2PyXVPgjRfJuV/5JAYI7MmEiXhDIPxrdwmivNCKmGzin8RdO
TjBonjknjf5e+L1MTzYUe2QJhftaPM6iq3WKpg3e457cbeHF5gZqMRPIR5/Ob7+p
Js9XhaSKCQv+iN2WUmcsNacz4hVFaaYXOSeY++Gi2agxLBT0w/j8ljxTP2UgWkEh
Om2QIhuI8CkseM1v4UPgwOIQa0WxkDF6CDM5erch7BCNUrSZRZIE2kw/S6ys0qfV
uvzIH/AAtNNDRocVWWNyGlKzSxcU2x7wyHkW2bJGzjofECdeOUb+rbB9jyAn5eKo
P41t3oEl0LaJpolX7LGyJm+1qJeqHhQgINQUFu7cBmZPy1LS3MJFugmhzI6WmPbl
eMXTRl0//DjBb0UF5/c+jR0mtmP+1JnxhlDwBRkzjiazhikO+f/rLhYMICmDNzX7
WL+QBJhoHTlNtX0s8xUs1F10bT4eCqyM/J5mKtbZchB0f/gF4sBTxzeHJ6fEnMCv
zDCPdYf3TBsShNmRO9iHc+CTAdoF2441jADPCZQu1q4rtAupX5+d/4xgCItrRGp9
ZkkcLWWS4l+OSXtTy93brYu52HjA+Hk7N5Xl5Y+SKfqIZv6Bc7WDrLYpW1AF+Sg3
rMlZnXhU5T8EQE5gk2NBgzNvdR4YxVMq3CTN7pFkl/0VxEG4dxttUSRavgBSyPGG
fFXs9mTFgeZJxHymoAygw7Fj0vJORf219Wiok4LrXuc86PvMtgjhApr5DwzmXNsu
H1Eq64Ku8SEA+mWIJsdQ6a8DuJKf7/fKGsXbrJZd0t94YzQ15kaiFrLZ/uUuIQ0G
N50bKdlxkB5U/3IjCR6IVRwqe3fs++1FSkSu9E/HuR/Uh3FasHbztQ0Po11zB35G
k9T9lrYDxhaJoYwBcobj1q5eO217XQRxjB+IqjOH93bnpNGFdUCYXP4L0Q73M2zY
ipLROewQ1d5PUxPh1mBaCIHVapaXeKB1dS1WJxYBbKfkBXanqA5AG+BpiT1YQi0a
bIx2ryEFdO/edfwQtBwuME2qfR+t0ld6j9WUYRxNX/s/apLhJGMRkBRAi5xVChiF
31eO7dEw1jxXwuJmfNqUe4ehs6dyABjFIPkLyuxBE0u6vtZ9bwI3VGudr9v3mOcK
XPURQcgIvEQWAVX4AFFYlRDGQgSNX9ov5MKR9b/e1m1fubVrzGM2yZOJvsEszfwG
7kJLQcmnIG3GvD2q5CCTPKuu+/s1/+3RHlTZY/dH1HgiyaE24dO11hrF7w3x6ZHV
sI+oZM6Aln2lbL+DXB2Y4iGfzdto7NcGgwVQdLxpJaRAsoxrMLEAtwaqC59AfzGP
lGNbdMoDuf2JlIoJzVG0IqIBEQB/cKIDuNqr8Ouq0F2mi1kMFUI5SVXF4sj31PaD
58RviW8eavmNqoGIeqqLzHpD20SOABu3J14oQ43oCQ353H2XLsRCVfJl5p5xK2tO
CKamamoQaGoF9vpdhSxIrRBTWJEzhzN94fwvYxgFCxeDq95x49dDX0lxP5Ypwzwj
hMhN2cGxfs1K0299A/NU0lmTk/aiwXvocG9ViCwaLwnuzQBN4fTKDkQV+jRvIi70
mCYUvk2eXdbRM7mtIggzzh8uVtu/xKCto9bNSFdmfGk0AGgwoWeujTVH35CpdznZ
rhsbg6vvWhtdIM5okDxm8vUjBevsFgmTcQavWIFPQZiA+lb/K1Ivf7bXGnL/mlH5
sHm1WK88YAcrkbeUvuEriVJiozOrbfA+NdIEctoGSBgfGnD91T6fxZkxXx8qZrmP
1w7iwnMwKkWNvtCdRiLltuQY8seU8w1tINWUkI39P6pWJS0l7kEFcAtlLUJOdOEX
etZxJvg4mx1TyteH9frzbQJLF5EzEhwojNgo0M1djpe/Y/eyTM8UuqHUeb8JYYZX
PbFZoXsUqps6Z6n7YMZR5kWcTcpijgsFNY4yeHK66ZN22iJFb1KRV3sDWRTOIFhT
0IYeKQPCQLjjvs805u0jWQwIxwidhGt7Nx54XrypCN7m8i5Pg+aWgltgFQtaHgsH
6exd2vXijZG/IadIAi2D7KOsixhgGuLOSOD4hMKm29phGuoYbaakCkK33gwLr+Da
IumWKpCDAkl8hZL6dErQmHD6RLQsuyzL9ExQoGSqqQw+0uatn/Uk7qal3ZJd+rXQ
j1rcQjhOwHIwtcawrYGiJMPpGdXWNXERD4N0VQ2W5T1t1BBaTHYrIQhEPpgE4U2e
B+ako8hGSk8FcpjP6sF9whwfR3VXIour7hpb0seGZVul1iAERoInXt3cSgz3KwkH
NnT1QRLol9GcQZPZ/61UoCswbNHlQUHfoFdKzWWpwRvJLhI/BmQtGEQpJMMRSaj5
kMya/k1JkyzeGtTCvG/3ohwenr+ZCZj6fDYPLoB08yf5E1QSwNKRPlxKkgxKYfNf
Yc4MSQMeLKkb+nm/LaFKW28bk5S4XGz1Ajb31HBUk1tcin6KOzQqFOYTj56fIT8o
bOg7cGZ6c3MYbf1qnC1/EJz5ycuqvE9tASysqLhNhOPjs8hvnMqOVqJbZW1RNxHm
vKmM0e9jjdGWfSvaKRVfHlhe0DIJ4BmdvE0M4DE7u2Q7H4kr9EKjE1dcf49NA7mK
r50wUuW9+dCequf2l2wnsOK2K/Ejq4sKY1dTx46yzUHNBKD7Iq16QPh0WWFW+N+1
+uzudSerKGJoy/0yhsCEtEhW402CLTsPTRk2/EbA8No/o63PbiKuw9FB8/wOLKV2
+ptPrW4zczAg4xZIP9GWfeMZAzQeEw3PiRuZkIoV36rVIULtNEBDEYItBYU3t/fH
YXDMIxKykIbxgpB/nFx56Ho/tsXtmzMDFL6sphKqfTJBvoF1WsRIivbCGLLcjPrG
V+NhoW6XL6Hzd77FMHi+4Jo05wcdbUas4xvcgcWJUJ3yrktGqtPQgwK0KtZWjIvs
cYT/RELI1hDJ8/Rr3/Iw4szjodjRIhb9UgOAo4+mOgxHUrMDUaPEQANGSFD3Cdkf
GPc0GscwnY48Y1iKRwNUudRruLEqZt9SQ8Vor0ytNPFX/dVQqg4XrPpjuhA0IQoQ
0lLOxr2+9z5qivnQK1W+Pww4yoFVP3zKxFRumqEXYU8n4WztejTQgaN3EouvGx/g
E1NUOAnWnH30o6BvBuXvZw69DDde/t5Ua2/wYb3BJwuR5FeUXxbxG3pWd+l6vH1Z
Lbh7FfkqQyhrSJIzCFqtMFfgqD+y4dfTR8LAyk3WERLijStCVPy76KSCmDszy1I3
uoyb+Rd3oFlo9vgnYUdUtUJu3wbhBsha+EUsoSJ3GR2qpwsfnqNjGTnsiNf7aFR7
ZcEJI3ADycHRFNsWTb0UM2CPOLZSGEssFQaK02tcpjs6PnatbaAmBP+ErjKdZcJf
o1RyL/DvgglGsQHA97rRGHN+w5MJBknhlPz9PPpOBxBwDB3lrVM8m43x62sIDtFi
oEoh5bU8VWODze2rYYXWJmSMOLXKxnDboSnsE32VYQi+i8BG6cQl+TE42Ph0fBVj
Md60gkl+J3oCClAKS2zbm4ori+lYoT9KagBB12eDiPmKgnH2CIf6Emi3zFpIbgmH
uMqgNWL8HWa2P4//lD+2fVdRfXkbvFURZ4iwG+92HWMLqmC7O+cXkVKGS88Pgcvl
eins08Ov1LsuSkR1HzzueIcHqIqgPQVckOMkc1IV9rYHbmm8o75sxBsRcgbM+/rJ
WEMXs/Cbg1CMYr9hkb7c91DvSj04Jh2IG1U8oyUUKs43WJdGyebQQjUSHLZhddTM
6MQJ/BZzraEQ5VUtngcCbvd7wgQEKcboBtP8WS0n8aWS5OUjOuNZqj7puYLRbSyI
GNpwN4LA2yfPhrlJ32gVk6ntloj66Ab6JN8++7lKx7nHNRCrU+6+J3rA5Vv3qeWR
RQBsqL8SrY92YMDTrUzACglovs1OqDQ9Zh/A5OlV9hvLPKKh/dE2VN/4/weU4LP/
ctU4wcIzCEYr7ROE8QfKb4Jh6Cv4SkpJZoUvgvdVFiNlHVZbsBXfFV7VUlnwctZU
igSPiZmibiS0Ch37wlikGW+JuwgLoGntBHgMwl1LWXjkzJL66E3BjSGvvXjN9K0N
Hy5ck5KlnLJhMyNhxTqI/rFEWBe/ocnhrF3Xlkccb2J0SQ1GShSW90h1av+upilS
YLrOQmv29TmOSyeA0AmCajrR+3xdX5TBTtvrMDHX27j2qyPfL4MU3aZZ5JT9DEWL
2xJRR50dn8M9EgxQE2puRcx0XJn0z6bj7jfeXMOY6TR11Z6wxd3b9seVj5eQzn6w
snBOGFkQbOdSE1ERgwtnSToJHDUezcfywr0TmlbVfu/f53xMwFeFSxSO5EZ8G9IN
KICjJ7Ws5jgznEmbNaQHezlUnatD5oDM8RIYrHeI/5n7m75SPo9rB9kGrbJ6m40J
9uy/aFptK35IScf6bhBgikcoiE6a0g4Wi3rC+zUzUHUzEh1UAD94+P9BZUm3Ix4W
Vk37H+HUSXqiOR6m0SHhIhuilm+pqAkuqwuDjiRqpNHNbZqhC9Sz/lTKNuvIgAuj
BzuuWf7XogX3zROQQtE+BEbjIgtpRu/fSVqtm0bS9MKKbx5a7HLvaLywfKm4tz2G
bGvQnsjSYqnemw8v2HqzqS37IM5oCy2t1gRNGgZ5bmgLJWpUNkX791s9FM9N68Mp
Pp0AoFw8S3kKcIZpbAGEjwFGxjJ0oqMruw/SaJtiUygCp1waXsm7VSNnsIpqnWOI
yZG5WeAOo92eKhXL6rx4VHkn6tJ3/Qe7ixLJRuLwi0Bzb4C17JVsEtdWiAb5FNIH
BeXNnj5qnQJBAt26I+pTJFGflQEvOWdU3NAnn3dEYFJJICuKb3uiJujIDikxn5QV
euiA6TAYrrENyJrUQoY3NUd8QyiYIEkFJUpMRlgVA+j9PTZ9090lwppwRn9HqJmZ
BvnEs27KlPjJUBTVv4OJP2M+jvPTo9KVzdp7cF53ET33Ekf7LbPp7+QKZabxxONz
4+nVNUwo/NgwtC0zp2+9jAFkoxZjZnVn5+DyyTNMbvj837fteyU+8lNY/j0yN0gi
L3EWdCbQ/vLsXboQf3+iWr+3vET1wqcae2P1C7gsTZzDVMvjNv6m+3HBGg/vWWmV
GOdkyfX/nlgFhd+zblZgVnG3sAHTDPasazNcBt7Z1PhWBnPgn2gE85/ok8QBTdYu
kroYr73MTICaKKa08hLVDKQbWL3UV8ZGsDZ+C2jQOeWd3xzhy+SBkocq6lGMpGmK
TDGl2yi6tgGuIbREAYHqblT/GKBOAwU6ic+1kx05E5R4A3WmXJYFkHeNIEH1o+Td
9yIglHo8FOpiDv8qHwIMk0W+IACYuth/pTuCB+Rz7u1Fin0PpttPSkxSujTFKdH3
oz+qzOWlc3iUvoC7oka4eF8n4bqI8Kd5CuUWnrfV8xY3QsU68qhA7wQulzhxS5b+
PjVKnliPqFGul24hNHw550pWzqDwTNWpuyRx1NPmJp5CMSBAjbHlrzcp69KiaASb
1znVDTRBrElf37gF15Fags1vEzcwsl2Tss88oyDiocpr9813vVKtwsWDkNMP3WpP
46kOlGNLdofYfJ6lo4OMsIanqa2gOgKO4RYcdAX2gkAnNJirY/yvtWfzeO91RsMh
pxDLzLlp7eZxfN5SUIubct9G12ykG+iCcn4OIDRaMIexRzKEeC2hCwulaMXjSMc2
XeuQg7txh0s3XMQ5gQkCpM8uLbsutWEM/MJyx8yvx/syPS5vP9qvvIOmhfO6DgML
hmWoYORDf5zphnam/iy329/P6QKTA/LTYEEKojRwAYCUxt4lqeMIJSlyRWdqiy7L
LMirBG7VFwXng+SCwmVMmGzMDtX69dLUZ1DdQtksuGdaFu3RPUakdJGlSfHDhe6Q
YcFi8+bA5bx+lXM6LNeKobP3vgowqsdHQtX+NIj5DoIzkEjnLIesRVXiHmf0G5yO
88PWRq4t5fhDq5Pp2TlfzqmMOabM4BnXiA1xfUjze5kFhDemEX+56V4M2PeIF5Nq
rDvPiQ5XiXzTMVIWtC22b69gaPgZQlTn+9AUIk4ETnDSksEkv8160/fcBg5N6Zi2
KeBzwqnMEPJiyB0FcsrY+iaoO/PhW4lXWMeR2UOlz9qY3lLguOPFV6eMl+70n1j9
Y751D1a81vfLZZzgjfEC1msNyp0fwi7ycgYNgSSoDgXXZnXaljU5E3suqGOZXnCB
COhQMh7Nu6rWPBvsUtb8APi5UnJs3zEzrBjY5DmX2v7dXmaVIiXFzAxPGGsHeGPe
67S6s8h2c7ObYl44+oAd+QaOquN15dBdLwLHycgtnjCyR2aYPagw2PjK0vz99faM
QCsPFUpwlJdHHxeHMJbKBvY21ELjlWfKRmOc4oekXuhwKftq882KId1zjo8eHNc/
51vOH6WdxBUfaEwdXQQZlERlXSWBR8lj+34ClLY8IGnGqq5EM3oR3neLo5xlZHsR
SsRjAwcCje4BgxfBCJE5p00QatfmQYknXWu1sSp7v+80Ymru0f6SzVCu9TIBgcGv
eUaUXAo5+T95Gkxyz15jfgzN4EyPPcqno4QfngL9k7ojxpICMJtI/Ao5M3cNcqP4
YN1usR7ji9PQjHgHDRxmeFjqGi6WllQuDwZmUep0SrpKVIl7VVq4dxz3PuvNFZ06
flTKkA5vkYwsd5fEgs0UzXNyLgwLqrBt3gPCO68kizYHd2KUWV7fMbyy30UvClET
3ePFANpFmy4SfLFdXp9Y1rxnp6C+Upww9rWMMg9c0wQ1XXFtO4auCagNp1Q/7ds/
A9Y4lPiJHPvASEOX/BBTcGtoFvbyhbhToAJ0e/8S4Oi/Skftwbz/iUOpsaj6UY3w
ZlE3S+wNF3a/mbkG2u0X0enPDGLK4HVOT7MjyzhlwrUR85i7OMg3R2gjo5qJpKek
Nz6rk/cvyfP9Jev5pWN3u7XVqocX6tX0IVVaY5yL80icRB+Mgp5934DdzjRsSV/m
012B9F4l1Xsl2fMAvD9+jYInJCl2yedalSzSJag2JIbxuoIJgeQS3A9hoT4nGpRG
fU3ot61R1fa31t/BOgwCA5ga50AJD75RNvmJoRWvFcKb1rsQyrQohSlNQIcLXi3B
HTgIuqo74YsIkEn9yaQk4wvfnrAmGrNG/jNVoudDTDfw241B5I4GrHtxWZ8QNpEe
1x4rm+lksvtLw9wXMlVm1ngG7KuYKkFhTgLEtVwgYNXYH2pElVT5qylQ9tlKwnay
jtKKjtMhMZ1fIVqvn6rShxNj+CCmcrx5NpGyZc0kmoKEelsBoixFhO8Q3utJDEOB
rgGFpCVvRc4kApX8z7SJ6c9BmOa1s0CmSuLyPnZB8czKMvVOccRg6DmgvP6qr2PS
tKsBsyoHUIP10NoP9lh88BU+CfdBmWPLGfx+yIiL5LfjFhAPwuO2CeMwMKvPAD8W
7KtbPaVOJuvf3XMCXF7IwJOvsViDrCNL4kMJLV5hUZiIYglwrog5slQD3RJmHVS3
oFAuDyJ5LA+O1mKp89GmfdGBDQC2IluuwFvCM0RQjS+HDtDwrUlP6ShyQcH4vSMY
74zTlhODeMakAykV2bPfD9esNwYBcefkfHejFnJ7dGfju74JgNVs4ZN+6OxIwuXI
9mr2bhSV2T9u6DMLQYEcYhoMq+t8o6BO02yhaxXG/RO/k/xAdVgtuPb4WVO+oj6i
OZzHR8P9ky7PkgnlkprvsJL8Qn/s5E6sEUoAuGlNB4emCA+hKH/GlA6LmRH5xL1x
syy5/zPA46Bulky8bhId+XpsO9FPSjO00grv1M4wI56egSo6Fz6VGTmVsRhj4zBv
FrJO+FnrLoZBRRpHTczWUtTKviGrEaZfyrsuYZAk0Di3wNKbZ0qAFkFzW2gHicpi
Tt0serP8mguVNPf+BFbgLksAbMw/lec2ZgYZkD4g4HvT6+zPW0JpBrE6RyHdF7o2
CK3j1hhWypyRFShvD/1dMe6urE+TpJNPx3CKHGHrSt5QCV6dKtDwYdcENasAowz1
GtXBHZrOGJWq3OnZDXZUzO92uwpkZRGKfXc//W5XnWMiylkZa2m0tQo254NsbOPF
aH40hyQVOwZAduefgWA4U/f66HdI9TWDe6mUCWfU8fcHhGb8J5E+obUfirdtdDU+
fNIPrkDkbfP97yw4I/zzodksg3xsv8UB1wTQNCwUbNkfHlKO/rf2alniZdWprSiD
gW7UZKX//XujQEPxJqMJxSq0gK699wGMqNxIKunE3MCESxzUl7muDxH8C3AIh1Ss
cQNyjhQLYGoZwYwrlm1Mb/4UhsqAswrSsZyxrxBSIIyLW+qOCS+oNnJgln6Wb0su
YaOwquZGm2HNBosH7mwksXEyvBs0u7c712o7wsoZAfzjLJK592lBy8EacvhK9v/n
A1ajg8zMcT6QwR7PdqFooHuZg3Ao+O5kg8L6hh3PpDQhNm1gUWLgQJnt1yGDEECZ
4mm7XvnPIfS1Gcr0Js2Zoec6/fXmP9PTVcGmBApAxISlGvjPZltouY6a/JThm/ef
GkGh1bw0yciEzPmNOt3pQ00mvFJsKvLsnSQuCWt8PDwx6xs3PFbTQ2wgYQCZwmTZ
YwTZBiL4tEemvV1TVBWgvIVzOspSNaQ/LAhTuZECFNgt0sQyOHCm5wceyWbYohl0
lb0OLeypK4TM4XOikoqps677xG1HVBAYbX6uS9Bhsyo70qcI0kzRkwKIakokFI6P
In6e58nNnVWRcNVvG2qMSwPJHQXZTVlXyfwCUaScUhk5LRChtImiVJZMO7RldVEf
rqXrU9PCpHEF1p1IWIpue/5Qoh4CiwCvvlDb0ZdD2ypdmuMZq5BrdzfRX2aS5c19
5wsC29t6RjFvR6QOVYw3HCUJpZfu9ueeZ0sqMgsTMyTJtTbOkmCgJAPm64I5jiRX
0HntXZm4cmkaLhDrQKmsylIRe8jEiMxrQefzFRJBwQxM7lY9Tldq7G7nAAfyLjrQ
XQkeEgAbBGYlq92bulsD78PizXloEX+Oyh4R9oYZXHbrtCc0XUxheCXx/lpvE/aQ
Lx1TJ6xvZZu0oUa/WR8plFbl6D2Kk3ncTFS7x3MokYrdIFPVEcjpyfSwzXJ42tNx
SLElorfoI3vBAeWNRkBsS9nMymM+EMc9l5w0KdQzes4fM6aWlUwtMyWb4JJ0MYP5
rgsarSW3QgwR2hSsBRV2r97Utwp7TbGN1fTRERYX/69DBrueacxLbuYqeceLXQYu
x4X+r6Nbv6ht+ipOwypIaxSEw6ghu3vk5BjJGllysbQQlRlAoWZFfEnHwbF1ZFi+
h6lNgGZq6mpdNAXL1oWNW4njfmfN6jux3Cq4hn+c1PeXy/hbD74BfHO7MG1lspJv
/YGdhutLZ30bRaMn8+KPxky2h5pgjtk+nms8IOjlordERVTreHFLCV7FJIfn1AdX
vxHV16VZQjehEdMJzZS9Q+AXtI9kDrivyCFI20qOxKHoVyLJN7dBSnqKpWnYWE3c
KTO6BSgPfqynQncxObEuynxjcP3U0uPtgIPSrR/uUgS19FQrGRGcXnLYnqd7BHvp
ngyWVbbPXd1aVtU69Igzw47Vq/yY2Ns2iyYr8fKAvP4ClxTudbIN5A4SfOArw1sI
lwSNHd/z8/Hf7a89OJynFcFvIFYQmYTIffVOdoyatbF2PKqWrv6rutdCEPAKrNPT
VTl034XYlfL5mFWCJTwfxShYmg0DQLDi17iOOYMo9eZjXwIxZ/UCBnlLRIrb3ZA9
WwtyKd/07SJ5SVGBEgWjuN46QjYcumlBmD8ML0BIYglwkKnwkuQi9mJAjbdHFaQw
Xdd/wj2WYoO9lnmE+V7MKw2uAirxqdPXmI34lb04sZGMeKixSu+B4bKSt7pmJN4u
mxzjTmn92ZUkgsgrVAipEB9Iglnsu8pZgvs6WU450sX9duS38mPQWFoitRexNPH6
tZPKHDimoU7IuQYYsUp4PY+4GjyzYSy4DWeisUS1reSaLWOaRVI5tHST6Dx/pNfZ
gKtjwCaWlCp5Icu0H3tu3EepfNgcf2vKdCeZC653g/EOekFFkdOEMFDnDhnxcbgN
b4vMM6rbp4vl2vgP5JO3QaRgf73HXzOMLDeLiuxlA/lEQl5bb6+Gh+CM7mTHUSiG
SHQ6druPwMQbZ7jem5pJTKJgAXTyeMc+28PSM31n0SOO18MzJkLXWskZXCEuZYas
6R7qJxRkJTBLAG6MBU/k4n4hA7FW8aCEYHFkwlBd2xojgOtNs0Bsjp6OYoTmOIEl
fOPzsod4OtWysPm8A3Dc+HfU3+2h4D6pXvk+4u1aWd0c66iTgE3t8cCoeEzj3wU2
YJJDdWpS9t/U9B8fgLKo90esgcm3OpoAePM6Z/a1Bd5SKe2lp2m/updCE5HNI2I4
Q/AXHGmeamk97woHbwPG40i/I+KrD5f0f2OtGE7ZCsQGndMo6GtCe6ObdIk0+n/l
uSeBAbC7G3WemTaI/itSb/1Po7F2y6HrrMWJ4eBimPKjSw94dS/9IwMieANGBRAh
1zVOfx8Pezloj6ZSIzByDQOjTu20fk4GbCzsHzxjxGunraBPW4cAZ0ENiINynkL3
vSFEAFW01dUbBCnqrgBr3wg8QcnokkcX/CyJEtkTbCEJVyD/ey+KGIyrIra5EiHE
iCSXCl8v6J1gF+G3JU9aGzwzhc3+6Ut0yVoAJ9me83Kc0FskrxTKH4pRLEz///Wr
fdElPyvraYgkNamg/41UQputOhIM4ZYIdp2nTzqLHo69Iw/erQqMD40lEzfCIviq
qDPzkmUncCRIelsEr6ke6lsCXzawl1Hmg3liEiblMM38HtWPEUHH/orOzmnxicEs
xCDHl1Dwkitl3FKoaITB6DdZYtIjN0SKB4MJmzWyoKgGc9XQ8bcprfBaJWyQsgzk
z4EknHjskroD95fJs/1iE4at+aSumYe0KbChQJuZiX/o3yYxhE7Jwk1/uqHYeQKR
s/FhnKI/INIb8kSThiQHEvz76nYM7OUGOz8d8oTytbVj9mSCh3ASSZroGf5siJyh
yxA8yTIx1HnKZyghmc1KnF7UaclYGCXQ312pqjlw/QoArR4/IAmvwy4nwZGbeBlL
hDgqDttN7TzfrwGmKBjstovL0dBwQkKguEXfza++7tz/0DHBY2JJO79q/WVVXLc/
7MoGVzeQzkhOlQ8QC7EC7BEjylYf6WxiHXeBoKL7D32ZLny7PUiz65EzOFwgQI1b
ZqjnOm17cFOwhHtIaAb8RqYVpBp5IugER5DwzY3x3b9Hp5gFldbMSw54jDmN5lAE
LuY59wrMXiMCkd9DbU3+qLzOrkTZJeUSvTc4TWHdFjugJW1NEm1i9RwMDCbyu+ET
m4zmzVyOKnj/xvgFBCeEQB08Fw812AiEKNLpN6SbAEVgYzA2fN+WSR0WxwCUsb1H
HjluNI2vtCGOVLRVfBZE5CyFh7Fd0xwxsJDC2lH9YQK0CQghD50w/whI06U3YlQU
SfUOOldUcbOAz0tleFDsgc2JfITPEkpvBgHW3KYOv8cBPhw1TgzKuqd3GKa/JhQW
6mKq3zosodP6ixI3o18uH9c+q8HQTbuMLX1VFlc9dAiils8EHmVViwf9Zn5jM23b
h4ePCvgfB+wR/RnPuv2V3ypdzaZ6uegGvHfXu4qGK2pXWKbtKilmHrOr7Rl0SoSN
lU2/JS0qBdsevOV/GUUTtjpDPxxuJuZ9mWKsO6xFE0UTZs73IVtbJHKXpJWtvW8Z
DBSZqq4cgFsKsXQDv+2EykesM2HftP4gO8eRoMobBUm9Q233ZY70S1xpyZOoAbYM
QtiGUhgZgtpCXzpQpW+bOKNmPtEyiz96gkMSVdg659GO3NRZzFHMNQQ0pG6VdklC
BOf1+FST+GL4mi1V2xe8libg3gTM/2EQ6sDj0wauzIWGdwD4wyBdijJBhGhG1Eg6
5cRVYWd3bc/Q+L2/SLmYlrzcuMiAkYuUzCug6+esvb/KC7Stl8QBCIvZUZSH54Ln
jEzwniCcUi31YK+TPCxZA2D0NAcZNZVCId4uO2ZudUGOFudMJP+QuDWeDOiOSKMl
lMj3QrBqXARBrLDpZ8bOSld7shHlOdwO43vWJc31TeMC2A3l9Lb10mrgOeLZliuw
ydy8wX4O1quQl7GTiPTE+hGTDrwihkNKu2NZGE2mwewqzqC+xjapvHSJ+uxfRVEm
yz/uOUOTbJ+lJb6q+r1KC8DDT03yszP3ZmcjJyPo7NqEBLx7wmJQAw+EAhhCG/c0
CXU0Nkpkk2oSFveMdPg7dtGxdEY3fT2MthuK+qPFlm2j/CKF5Tz4+utwPs7OyAFi
iA4w8esm+L9f0aPfb3RvCuHB4tpkgO1Qg+f7upF3Oh+XYjcPOdA+0k3HZMMdVaZi
/lLS4fqFzW8wjgHzNBEi+KtCtsdTs/hJ6oh+pyi1Ry14kiKCdYoV0xGt5YsJhuW+
odcGvWe9Ibw55BxtEWhmwM+XIvVeFLL36TFhc3fGn+Bo3qQY1xjU9YtOuCX7hJFc
yPU3ur3Wagw/gjqOHM8jWgfxUZXbR4iR0dUxJAf7BePqH9usUMb1XS+RvDFe1qik
jxKq0ope5uPfqH7guhCCw38U2Bo2ZpYnYANbw1jXfV1elS8OzvJQGIB4TjAmOKPt
Lj77S+/vmSagJJKdc+box7v0oMoxZoZeU8BflKiu/iQNAYYMJzkZzxmABm+Rs9qu
/P0g4x7rT/5uBKWY/vwN+3pJuD3XNXrsj9o7h9Yee/wn9QWLTvGBqAVqiAXGJjp8
NW5wVkkOwIM+mF44NTBmaFTLUmVkccVJEW1IzNGEtgRg9PjtpPDW0H+V0rD665pD
65czDHmxOO2VcPn6UUgpI9dW0H+kP2jajC7adNmc3DeUnnSZs6XAzm1j2Ufz5UJo
sHvbxP8xYd85Fve0rrvK9Kdx4Bb6Nx0lrRY9uttjnWXnltBttVhik2kgSLYcAw90
D+XMHnNGhN7Rf7PcKnqVrbO2sk+2G502IlbqyzpT37xxBqdZNFGuxs86zbxJoh+j
LSVt69SGq+wK7qXPCJyEyvUZvkoZyw80Wuyv1NVB/WyZdQNv7SZPvD/gn4uiheDM
pzTk7f1ypu7sE9FoG/u2LeGpJF2fjbvSXXXlgi/1TCuxCP4tkzIjJFRZykZEz7NX
uH33ebvIzCFR1EmSxDwPYtXoCzsa27pC/4d82mlS8xowHcAqqkONoI+AGSQZrPvm
0oBsz3C4c4ijc1HffE2YfH8c0UsWoQMcTtsIY5G083ECJDeF2cT9n83qYTCkI5TE
ofQzE+IaEWb29uE1HOKGimBALGWRd8prj/7BGu9J2aQjjtFsyddW/1m4+5gCyh9U
cJX+/5CK+idr1A53fH7Zxe5PDcF4aeKNoMTqq08SFTd0snDqj7aSDwpvqKrzj4Yy
h50rniRnQO49+i7srN608437AqzPugi2ixfzgBG0l+yOLk5VMTnCs7GDVM/pUIoC
exoTeBa7SoO15aQDt154Ggu62a/Aa2p6M9c0HgoN8v1/HPdIgDSGnEJzHmJvEuMl
klwS0/kxs84ywc9dKVmdEe6dIgyRThH8JndV5U+HyqfLyxP4UCfDNUTOMoa4DKau
ji5VUehRs9ztQ1m2iH0cBF3NutoZ2hjYAy2SHpe7nMzbQWjNMFrYQuzpLkxm00FY
gQggntki4/pdjo4m0qxg798l2ibFlreacKiRj8rE2iT7Z3CYvp1fZJgCFXf+ptwa
BI+PO2NxzzPjIQ6JzxfK/2Tdcu1JIFt3iI7sTn2uH15FT3bU0BRCGK7aR0eHb4iz
OcWdFzkjhtwntX/6WX7BIvUI94dhlI02shDamFGECvzUEHNa2IfHYakgVnXkEzyM
Q8tngoEzgg7v3XinquSAcsdp3vX7fS/Ml2K70CB7bgH+I+WQC05VIQnADSAjUj3A
zgEuzYq3IiRSkHxt+qQw8QmbqG3pvhxZRa2Kitvt7C4ET+PEyLC2/aobtvszubxs
M+uwi2kjkYGEObyvgD751rRg+ljc67Er/h89aWfQg+JC+/3dcItXuVmHatgNrLlq
oIHjLINdtxfVvlO+CBu2C3tICMTtcifNErUuHKDdvQCVpsJpmEylFBBGSzf1YfPZ
dOnu27w8mMtNu62iIocd1CBnDRqqB8I+Wnkb8aY7fo1hSU0SnLmgcMKeTVvmO5md
Xw2+gF1mNT0mEP2wH0pN9KZ8isu0HuLz/OBkuwuMPiYHSCwZbRGVN7GdfTAo84VL
b3gsxN8NeTUep8F0yeDjob4PQOvxi8z1bcdhOZYmrKO7cZrKBUAVcJ/aCeEOjMHW
GobyG/gnzipih9RNEE4EQyy16UZfHWy85juWpuwRiTTjfKz/VnB7UPzgnqYU4W3A
3GYRNnTBpV2CpZHck6jKa3eddBXJIiyPJ8ZQBblTphsTQWy3LmcKC4FnTJYbEpEM
LRRp4TynpckLWupestHMaKFO6SXJSXMWtX04MjDXBxSmarcjtYoFOAV0sz2/gaEc
OS4j/otahUWcXwBDcnMJpF0ace0XFglpe5JZDNUI+AlkLRf+v7PMYSMw9GUHvn/p
3xJ0u1mXad2GPBHQAxNTioWM//pQDP4flF82UlPEQWBob1WYF5nRR5C6zd7P3h5q
3DZfWIV7kJDdNJH5mfZQgN0AjgCfMqMD5xv07ia1kLdmV5JqIFX402d2S/2aO15w
TO98w/IUixWSi1FJOXV9czO1wcCFX2hzCTQNClrj+H6lZ0SGezU/tkV65CC+l/kv
2/sD6pWjfAwM4yVgV8TxLuTMnRJyON5C6HZjmzJ9n3t1JAcERm6EM+e394Mgm4tO
O+McLhG0CrqenSvIWDzKoWK9wALv+Kw9aa0f+Fh1r5Z7t9R8IcUneVBfC01jc1od
WV82osxAuuc675k9yRhia9FWepHG+hJxqX8HMJzjAAoWLUG7qCgMVEMf5qOAzgXI
MdxJnPLXGyOSXReJ7iamWmCxp/4yPzsCAzIo94i0IHTHqkNGEaJgBZXnzgUGkpL7
V3MKb2BALVgLIMaNwlxXroynnLA4Uc+BVXe77BU5WR2L1p4J97O0lfwC6YRLjwm/
HPz7SeXYtTuBwjS9ifC//6crjMiO9V4tKTzqhueonfvChB2vkm5um2RTZgwvYXDY
KTRW4zBwjSJOOj3eohK1ONLeVBseKISQVBJ8cPnRP9mXQxwajtPDu+XfkJ79uEbp
iNDbLOQgVWVxQDDmd+CO0EEhSLHO8CwZ2p7GWr11pVfpgJoKSIyp+Akd1HFw+vF2
cQOBxHwjWDTw3hK+UUGLeyLyDpvi4GPI6sBo5HOkyrDsy6h6WJNqkLfC3RFaoH/W
h/Z94qEZgmZaXOPwdyIih59B16o7k0I3MWynazZkUa87I2tFX5iIv0vfwJZD9Em1
Ed8ReTy6wYrlGm3cDiio0VD+PVwtE9DMbV5xCIKUc22m0IrMCyTEb9QYsirJBilU
L5XQZNyA90cglwKIjrbzMtEcmvwTvrHZzySgxaZQ2jUYRuyEuALcbKVEqAfe71Kn
abQdqWK09PRiA759aDlyTUs+gMecRnA/22FBYMQ3Lpw/a340+7kRk2GJMeZLZ4+T
C7BO0g6ETADX0D5wbHIODBkC3+C88CmrWadEC+Y0lI9WBXuQEdGtJ7xDrJrzfaJu
n3VyjYb300vqlLhyeUMNxMJ7cZPcDQ7Qj+F5Wk8hOiKJ0wMNKaNCwZlUpey6GDv3
T3H/vCXszUmA2wZovvCIa9ZbxYOv28z5CKGXEhBZNTfR++qOQA+ffH0bl3lAbc7i
spLwkoBMk6mRtTFSP+cfKh9P5siyr18UMtu9hCSmGOpd8UruhINJny5WoE3CpxBx
vpnmXo+RK2FLrWoulOGbgogCU4B/V5P2lIglPonCgB75aQvqKlaGIpLYe82fhr+p
u9lKlmQ/0/A5EMoO1vn7YRwpgjYWO68+8Ij4zYW2b+puQ7mDdplpXXsaOuMsTdd7
dr792+MklQh+QsqehcxGBb456gPJmPbDI+QOb+lk8Iit+Eu8ov0lxzWtrNCHVtc9
WJxldiOexLZyXs7h4SbNHDK3P04QKsl+vBXqXwVO5vaa8WF00QfRHEcK9Mt4j5t5
F/oLdIwP0xTNEDzGTZtNYnv7WvILL+bmwrL1bPaw+b8bDd9gYyC9sRwKP9wWi4DR
4OSu2kk7MNvlRVFQpzu97BgKuDNOMRveBP2n7MREP3dRHcCFxTnHCMKyyn0yqJ4x
/yOdhl3OrSBHK9GZoAlrii5muAcs18MQMASrcvzbOiPcyEinbLRpat6AJpGf3Plz
DTlAVpWw13VUrvFs18Smj8nIqr2R7TVE9nlhWlRAGf5OOrp9GYiAo+KRu3rHILpR
igu5BZOFymHaJTASL5TtEZzJpCTlJyw+lqF3/9sbNsjQphWNJU74MYcqYXn68TAp
Nsw/QBgwcAx1e9M4WDTyIw4sopfKT4z0QNsMh+5uckF+OM88ObRD+tZ1m3l/hmzw
gJ0hX0Q/ky02VDTcJd2+dUwRlBAL6NjrFIJkxnx4Hc9K9T4qbme57QbNPCw1KMsn
BYOAw8Wj5W6PDOlXxOh+9PuZc4rT4TBhnNE4YcvCDTr6WRxGynkMinVoKW3Vu+Hg
EyQGtO4ZFQmmd+py3WUjzC0FQ4fWzMQ+eYdDW7dldsh9KscXT/fXWhnEJToBOCro
MBX0UKMmMl+P4QamZEIT8FAUE4AfTkzMsbFy+0FAsXZ5FRG+BJQM0dtuSSBSIetW
J/dgQtRoJryUKX4w/1PIC7heUZS6wKSeEDJ6KOkH0koWRzOCYa4G8LAkiKU3b/i5
nxj2+PrY9gCPVXVHyYC29jRs0kX6SNcuPsH0zzYGVLxprZ5QnIe2qp1bwz2l9c7P
O1MvDS1VbBD8g1e66kSjwWkseANVdjBroUEEf/+dvBO9vFYFlMBbecgaFDqMsDX4
pxTDJONalLrPfJlRbyutVc0/8C5JNWhIihfJK4VtFmbjPZqyM1+skFd5Y+UZosLq
uIYJP0tU1SMh7/Iqhx4cl4malLkNCsY4e4qY8lSErabEW93aABFT0nRRO3TBPxAZ
Ej0sodg+pYXZ42daISZW52XCSU/A5i5TwlsQLzamMHG2R2K7+Cm/0c/QOWWr5pZC
sZlA7rFlml6tbYe09Vvuj9ccDpgTTZ2BMashQ7BQWYyf7csaEYD16u1OkxX4Qs/g
nxMC3+aeqhqKSBrvLJhD1AcOX5Y7UK8PDGstvpXEcpjqkwD3GixwwnFiSTbOBtzK
JkVF9wDejSsRxnyVDG+6yDQO3Cgy87VUqmcb7cd9TccfKccr9QoiU53PfqNLeqGm
MIksT9h5aoszcRDEzWPgrSmbtfhNLlCdYb8CId7mi8rkRMY8DcCCfiZ64BS2EKD9
DM5yO0DypfsMtceD2Vndvr8lrNMTVpcgsPbC7VO2+mBQG8sfCPs0c4hjSLMReIrw
buGOlTe0nSXDRrzO+skpBrR6FHQo4dzxIYfTMlqSbMDIecJmK944KwklIyJt1z/6
oS6kpoXwPZIfS5KuM9AM1lixlQSy85SpVKla2wj8p4F7Ukr1oDs9yDiAf1UdBDbO
C+ojg1woJXts1uE2hmasmqC7xex3CMkmSJwa4i4bTtGc3bNh6w9SR3f69jVZYODB
Ql/euALI2tTBbDvI5m1MEFoB2AYdwKCc701hAxvNET5OudMFjhf9TtykjOEOVs/w
Czi0z8bl9tbzy3FO+76z9wzn9Mmi/x7+4w7Cp6ihZ37Y2oCJbtE8SYssPBQjNN9R
3cLaCkiwkCg7S49XZQ3u3FA4W74hhOL0nhVQrYSRFVQh9zALq7OPdojMfywxZzzd
xG3aFsu7TMJE3tYzSZdhTcrpMAVkcsBgqRU97ofECvT2dSg3gwkMXklx2ajYDaj7
XX10Nu6vHKNHFQ/CA/SBW5eSXGAMYA+2hH/22n2yfMK0Wcucd6GHrnR9/9MNq/3y
J5wGWbVNe+OFqnLJHQjb3O0JfsN39+Hgcckc1NjPw5chL7p+TEAayjhU1vMhrKG4
a4Zeke3QZUZ5B0eSasaoeoahhOv+IXPgy+vtSQCkK6XfqUITMQMSK9DfmsX6VWNz
9KR+swLZroyW79gxvcR5VEbpf1pwcVc4Za5O1vhJXDUCjX80fs5gXUTs55kT7Um2
bl/lfejkr9Z9yrzNwFaKWxJHF+3M6Kl84/9H1EwEE3JdwPdaZQZJIfISWtxLzloN
zlCWReBNFdazUoYWOz1gYL8rgbpjAtWdYNu/wPKj0OX5IRc6ErKdHPBygMQtfD03
NXeIIw3XrngyTcaJA2leROKe1zRr8WzhosKvwIGAHrPednnCcYS9hr+0q86dbrwj
7/qaCAOb/wWU4HHflPmDuZ+C9lySTLFzP0TXaAbiGOnA3V/Su+0gq/pMizDK/MOq
bHOfvYwRafggxa7feTMgDQLjCudcCJN8c5lsL3Dp4rwDZn/0fe0O3jTUYxJThfhj
4pS8/ptEIj/kfN+a/8Al8UBHCl+6wEV92tl24ku9KgLn9c/tbqLy14c6gAv58QB5
ZGsnX60JrHOyXUzsUibrWbuXIHBqoZhF7xSJ5qQeclz+adulXBtjFzEGa90uwAFV
3zBopnuN07bkWcJcX+Ipp1PmbZ7rEPvBq7TeQ87yxbWRqrNqms0kvngb3eJCiatN
YZ2V2OMvpwj+7pojLHKsUrPwOx+xD1kupVfpq5dqGWspTaH+K2vv5XhwdRayxXPF
7Pl5g0RSw/0QJJlC7PLUVWB+L3m2UdCU3udnlO9ftFEpjY9BihTBM65EW4a/1qUm
DmhZgzLRB1uQDkHjvzB5kME2Bfvjq7hY/8n8fHclRl4C4P+Lmd7XzJCupwTCddT6
+zXmkBhFvux5vao5CfVXX+vjyQsSaU4qKidIhRxKQ+JfljRQksWDEAuUQH18Vtmu
DwIab76B9ZUFyKIgKmSzY/JSJlfne789MJCEojjIrabxoDfh0Cp5+iGaobAy678f
KRkRkgKY3E5HZXo4pPsatjsrRZoG/7Qj4crcolJuWV0jU1D7lUpZt0N+5TPMPbTJ
Q5M1i3Yr6UR6dnOCNSzrsZbxWIrDOFyOrk1C/26y0suWYoFG9BoazOwbS9Ur8eIX
8QHLHOTGOToDrbLSQ4RuPFnfIiWk/vwZmBjgjTRlRRK+wPjE/rOEd32PYAJkMkd2
ReyOxCyZ6La9PuA7PbQwsI00CqyLL7gxO7+uQXRP0zke1DCAWwUFSlZLsV/of5Fd
9FNF8TLAXsYH8glQlMtIoe1RruVyAbRDkhVFbtKhrMJ4LvssXQnWx2Db55zonNa+
EfucSP3liSAtFN6i6OLz0Rf6dnKcvduWTutqfyfXa9SPq/RYVG7NJWRcghEU+6wl
vIs+Ucaqa/Uh6/ntEqnKBVEy1rth+gKVX29Am3WHhoiCPAYQkRqQM4tt4XU7KYwb
9WmtBKjpeQUu/rFxrwB/7yLVMO9Pvxutseq4LnGqrNLA9rHW4/y+lmTvmHxSWAkd
3ZzOjUzyl2KqzkoCGrqFbAMgeZCvPsdTJsg6eAC+jcnJ0Uayk8lZlRLd4qoTSb+z
odUFwr9Cf2rkjGXbvIgMxdBUmPwzxt/KvqI8HLgeMBkgDu1Ek5jDXgSyYhBhxR0l
o8K49Lz7/fS1TyrQQh0FR97hxjHHztAeLouav3ZFPVNUDDuG5CLer9Ilz7z5KaIS
EAKdB8uC/pw6iTpr8OTtHBvEpuM/x/KzItnGSoUiJmikrXy/OUgX0wTHbEunJMUH
FTNequnCCmBVnFgo9XBZDYnuS0hmgWxrIAS0OD96uBxLPgdthXE5PLbcWjX4RKjZ
oiqqEGDOpNYxNjoMqAATslnHdxBZAIitc+7OExCVGGkOrAtt1/yYkAZtakJIngzN
WaksEi6NMjxbU6xU1bffd5w4QgSH/eQsemDuohrFuY4UoUhNDuFsSX9r5nWtaqDM
H1s9q+ycj6zY47zH8GlOZOe0C8walPUErBGYqxZ2ljLP655R98eErweRFdfAXD2K
rkeeo8uoSfiVOGu96G/ACVh1STMLGf2qCgGZyG/mZO9O5doWZ9zzNjQswS7YpQyw
qKlQ0suf5AatEdHW3rvd7SXtwErrvJrUIeKNaWSHVkVHcH+ehYpyDh4y+3GtOBai
R5jciHVtw0ag+g2QYRVIcMJSbELOf7bSTP6y7wpM9biZSsvBH2f4xGZbzfYnIepb
DoIVgj/gGWohLMsUcfi8kmXpMOqIt0JelLYLvkyT1qDMGZW+//3KrN81jxlYKgwq
v0BNL4ZzwBFrxvP2BD3HkTAsk+cf9Nw7RyDLyjm/M7vQetBenb09Q9Riux6UNjX/
FITRBViU84oxKnR18PCc/8yFxx8t3wdH91ckPUvIpIx17OmpoL96WLuj1c+zwu8W
CqV9y6a5E6VbKdpY9hmV2Rs/XrUfrH1lYaenzd+zKwavyVw9It2KVWiZiaonKPAE
2TttS46nHIAgrMOMxYcP+UP/0kKg9emSzBApTmwDuhy2uXYqwHu8sHFybiO1uub3
m2vq9ZCMpTWQmWRlTBbW7HfsFeyuHEgeBD17oSYmee+43WZWehtpLaEpolOIrJpp
ZaQDEFmWTN1mvruVjZxBzz6J0lVqa0/bfT5tGNAPZ5UqUufqCGPmIJO58SUCZfgu
fGSUmPAnqvDPpzYUYv1vM5FHjPR+p2LeO09diWCe0m84OTb76ii929CPnN1XH1V4
U3Y5yltzJMUna4XJq2C8WNAqUq2fsPg6UySI7ZAffQw3ZrcpydWfOmpwT3ZrMi8Q
wJgJdJvaD2k4IO95kQ9YK9Z2xCEpzFNWrcXJ/lJWdIBFk4Gqvzh8GE3lFV0hI9Yq
aIkJEy66EbD8ckuhqGvpvEL2p6dQP+/Imjh2Qs3Uh1EMlFF+3+aGjSU0jBPQYbIN
/Nz+ffdLX42mATtNh/i8gikFZ9pUTmcVBxDfGbijmESuh8wKxDQwfmQ+Vmv/rJI+
GKbCB0hLgO2FFAqwhtNqvyK5w3LwxLNrTnt+daePR5pL7//AFfGRfx8mHa3RguzS
cVRW7WwJwSH2v6CkFaQG1RInyACokMUCPNc7mpN4pu9/yYfXw69xGoB0aF67A/rS
jMPjWc4jNC4F+wkFW0fdj12/3J4cssqf4S0aOEk3s8LSa5+cssMxb/xc3z6x3+Aa
HLMGG1LuVZaI5+UivCbuxTO5S7sXwnuRDih1xRfJgyNnkk7zhR6xyhlf+LF+Sd2L
W2WC1SxBbKkWIfcuQE02bhi+wXx6YZlQUhEv5MTIdwt4eqLziJ16HlmgFYdaAo4t
0Y2CkHntv80X+Z5EYLdg6oAQT3XAnfMv81ECHv1gCkDXWkOkDJmitZOaqnmSV+FJ
SIpuPngDQQTcobMons0UYhLcianx53TLWqZDYbhUi/oaEL0Dk8pkXAPh7f4aTT/e
kuR23x1OVR0CcMMx8zTqmXM9KUewU5gpmjFdsBDOrZaAzVR4e+pYxcalKb2Xmc2a
B+ETAu6EZpdH9FXB/rSvm0Ud+KwHCLWHXhFIMsSFiy1XyppcP6o14XLxkbvKPgDs
hKsi5MPwxJ/DX0sTFI61eDZBu8hhS3/4JLBAWzn7nca1UE4wXCv0LXlxYvB4b0HQ
lfNKQ9H4AhHajl0fxzCn+lKHGe4afumPIz8lA786RyyTw0+Ub6j7IbgRpuzVqYtN
Jvsxyvnwf6z0zWUqUZBt34/gmoSjYkAXeNY+rodkZSyp91FjcTsZmq6kElvC9yyi
CdSChANPvE2AgJb2rXxIuidN0d8fW4z1r1BaQ8fVGHpwjyTbdiClxeYQazvXPUQL
1lRdMun4B6JxoP4b5f4f4c6Ms1Ov+BcDaSc7L3M9e2GMAp6WlH2zZDwbV//u+Izm
cdkI3TWov4A5YLNEc+d8fx7DINSzcG5YPMPtrKOPhHuhkGAsF953WCLw/zs0NzrI
oPKYQ38TuD0I8xyDuZBfaL0U+QFtSGpYcwHxii7vux5gncPywLDvgpF/rB1c+3Ke
e3tZiM29YynP7FhoTK5vvLCNWmJZHLdgIF2IBgzYbv2JpkFP4GvZJH1AB/HxS4TQ
/SHtAGPOTg2JX21Ko75l+BPOqByvwkXnJT3ygGFRNbx1spkW2poWNia3/bNTXc6b
7JtC0DlZ9fS4k0g7HmEsRIHMcuYxscQsSudEU0OQJgDvNzmRAfE674ACPVScrPVN
JX/YFOTKNE0ufR8dTrMxzD0hsPcpwhKZAz+minz4SJ38Hg2HeQWZLGmRQiVi2J0i
7J4Czxqj9MqdzK0XMUvuWlzMdoq83hKMJi344aTc6AyQ/rArqfGRqottDMF2hjOK
RDUKTdPk0UaVJyz0ROfhd1argroMT7Hqvy33nuhEYmLdaZxbZEyts/8d2XzUUyfT
He7rwaeKMTEbJyrrTLcNQcFuzCnNqbrJmjUmRUPuxxSvKxntJbg7yf1rOetDk5dO
BYadC8cIeT7G5iCJhOfp9qwEG0iktFPrNoNFRk7zqXWdJKawN33dmAtzBsaIgkbJ
4Zsbjxg154Ttm/9/G3MvckO506CB7qouU08f2s2q+tmHabbJb7GZWQTdg6V8H6zY
gN1E+is/JiznRHY/XRwRSiaZqFkf8gUt2zBV8uZR/y/sZYwSMXcRJuydwgiq80Oz
B6WrGv0pk+6uWj0s+INcZfggVDUXV/2B+5XghSEeRQicjaNSQviLUH2nnCTgj1at
SPk9ws2fzAyduJ2a3TSMki4UXYo+2Qpx13QmlHHUQipKO1ge+0B4l26Mp4443xYy
GK51xCflQPNeRSk3Ud8J8zt2v2zVebjWk4c7dnp2DbEwbet/nprWw53ZOCPVDO7d
gf8VIOgQU6OZP8xu+y3IZxe12uDeKtnko00opDAiOga3Fuk5K/dcDOc4gRsng0Kg
qjr5MuBEECyQZz7GcOfT3Dwy6ZZD59cKCyqY51l9CBnbWftoZ9o+SUfxcwJshcaQ
3xk32hs9WGMycDp9+gHvTXaXvAF4/cv2t8utmy/YlM0Ajw29pcJQt6xAHwCm2up/
JxiekPDdofzzjeCszl/pvu+0/XSkionr1nwA/SSYOwNe/Yp0pGwwwb70QqLVfeUE
8OO+kML5I6fBwVSarp+UqFtOTTDs9OMbl+OJueZz+5ykoGwTik30/ZrBDs2H35+y
Y8Gkdw/UkRO+1SpRuZoCwv4ucvkAjeyMmh5jqfQqxKA8jIh4znCW/HdY15DgW/qx
srkqai/4qWHvfjTPcdbMwoLL3kONMecbLJ68Nlsx+N1HLWvL5xHqqHPIOjLBofDS
CznDu0dQtq3K2Hb959A4eXjdsFqU7eECn7+XEFxVpc2v0DXmqRLIWjdhsA/Qnn42
5wYC9fgXZr11RBFd+8Kjl+IGkxPW6hx9pny4uCrBwJ/2sPP3zsu9lzYxCJtVGVCn
I/GQXud/AARctmUwmwhK51QFf+ib41rDHWB1gJqdoM2+GrEx8pkPyPCWIEaXBUQQ
ovgBsoGwVsFWssCMs/UR/hAvLsuFR+zDdXHwhi6Fzc4oIxoysC2S9H5XPuriH107
2RM9+/PsIoRA30SoR2h1UmH2bUSbJtXi1EaAgb0H4jiw2DrB+fOY/4w8mxr/ruxK
fo/Qia/NrPmlY0bVTaLh6EjsU2h6z/rrIz+jHFP6LfDi+KAUH8bp8XC07/99Ijm1
MBx0lhwKCJR3Yh3kH1wuChAMqYtUlBrFidy7cq6aGDcQF+YDmebx09XbwF+HQysn
1IEJ5iUewIPRGTunqPzKOcklr8klI2FFxJwZaPN1pnNLmZwsN3jipCzgqmU+Ofi+
dh9RQgMvs2HzjgPX1I+gHrlfiT+Ef9P2JTA6mfmzdDba4VaKJf4GExJUX4Zx+8ys
zhgEwxtO5AoZclRACmAeEE/G4H5g4RY6vfRsyFd5rCnOMUUlLelTwDcolH+3cJpK
/L06n2MzFEtiq4nbMvJmselg/NI29WCRjj+YmDzVBHT0N3fUUcRqf12qJjRIOHgb
1Zx4ZdhhujVumddI9VW2HnDmmc081ob/KGb5zG+OtzaaD+eKUaVEi4So1x8MC4Px
9+URf4o8KiugF+i/AXMJipyabcgTTswLbEkRaPRbPhS3wSUugwRrAPTy7Rl2AMVd
yYAR3fvHOdA5lvvcoBHvPvbRadcMczixNLO3k7yELZMKesMlqHP21QlaWmLtB/Am
Tnv1xwLwguLFTVW2hv5oeS7aKeTUeDkTCASATl952hfjb2SxfDV3hweeGL9X+L0r
9Z9whr37r5AqPnMQm0aNpn2iajtM7qrunb/ap/qxNMO/A76hreUFPUO5TvhRSdtF
X52w/ifm2QZqjwTU57SYxR0eH+jjjpjZfYZDjGcY595h5dvWVpKDdlU05FyIwlGE
fllNWwDi2Qe9jSy0+gDBeFVBfuc0bZhc08vZq1CAUm4HG0F/KztIc0b7QKmNQQbu
DzEUPxxtfOzDVOtwwrQdyKHSRQpGVD0DOV9tn2ebND6ogv26bhupVl25Cv5ZCf7N
sfu9EP99MgaK9Q8h/1Nv3W2kEBiOZFT25L454KA/5RnzqHq5Jn3ZP1m6lO5Rz1j3
VqXwRMubW6TwkrhfPfVF4WeTgy8mA8KrS3QAXon31f7h9gFdeJQONT1kQVTiFBBw
lNXH5s6CPvLxyLrG3N/fxQQYexBE+/mouzjfsoDWWCUnQGpm+tPo2jlpdjwveDR3
BcMwY+WG2O7q08z6YAfYPkjrSyHCt4sHnhxJFZaxWHhlA/BiURlSYafkAafc+rD7
G29SUR2NUBSNkHu54r4T20JpbppfqpYLuIpoKQKHmu5SsC4AXrCa3nCFuE4puhgq
kIac/6fH9KwLgaCt0o7/294xlf8g/8D/smggb3dQTpWOPZrxsH1m5/oNrbclvoJ4
b1EcbEZAHvly0n/07ygwqts2ef+iR/6sGHE+SM/kTlA8R07qgDiimuFQermGOvOB
7et1Xk0EL888ODD3aHOJkgDuH5uAoTBg/5HROFT/Di1qzYEUe80Pnn7d6WgaAohE
rHeDqpO6lQ7YcOUxHpT75TRqkZkv4zpW38hHOcbAQPyGJkyx+EbVcaXB2Ucwj8eJ
4DIx0tKYCT/tkJUnTwgIpZrcQEZoSkYSuuRPkFyUq9ziJ2m1DrWAfrNqhANeMPjo
xJnVlQxy//FuhIdwDfYv48oyZqWynCGAd7URYDCwBstcHxjUFJ7C3coxsmnWamyz
ERZbLHfFM03JGHE4Z9binIf6YIEDl1ECxEYjlwOQudOOIrNsJP/CjsiRf/M/6tfe
HjBgGq9XebYvcCe8Z9+Uc8KWl4vXBR/wmg6YwU1gA4lJxwu1Tefar80UzU0didwh
27gX6twfhUMj2/199b7YgCRNZxtVAJ6ctAPnTibsaIZ/+Jq5j4Xsabei3e+kCwHt
Q/rrJD04D9FYD+2mKCITeFkILyi+KcmavZq0PcvxakCHkmOrXon5r5YjIsGO6YmG
Hgi8N9B20Hd3MQY1gYr+uUnTOgbb41ns7Gd765cslAbstI8lJL+xydoFxjV/IovT
D5p/O4OqE9oW002iGVWc3UIBeXqLDTywY3Q9N/3YbgywlafhmiLG00g71KG5uyN/
loB8MMbiiI7OdAFjG8WfRt876RbA5MM7HlaWQBZyZCtQCKpJdeAOkqsvHF8vPZQL
Sspvn9zoW8EfGOWr6kkr9xgu8E7omB0qTMAzolJe4QgSpwsRLXd4YVBoIrGk2lRS
4/EqSIY+M7a4nvRgKXkmxEdtD6b4iMWejHlzy6rt55m1DPJOj1CkXv4vLM3TqhW/
hHqVMm0TgoZmYobnZa86eKaV7XYVi1/b2QH2xAb8OP/mnGcBY/OFe1iuefXkTcBy
b09yeNY/PaFz7EJJFFZHnBS6PW9Ig2OguSJZkfkqmQqxvZ7ftxRygUiWF1h/CtV6
okjrDsg3flnyQ4+EYQDg5JGRiz9UPgrbDVBlqV5ph8kYZMmJdg9FDN6I4kVPe4vW
M2AlpEg9kF1KWDG500HRMpfhGwQqeX5vljLwc30f1jnHIsqaqsdspndEHL0auv/e
Fq2p1F6HwL6hL6h0UqYNwZy30XVkdvQsjGjjEdEqI+Ma5u8ldmMAXvJVvk/9JvMn
zMwRixNV2pNzjvYSFQT6tz6eq+xShjFUvQ/rZXX3pfB62zl2T5LJGdY0zPvOO4QB
F4hVmQYBcdNFOw6o6gKU3Dh07QRdMnvOI1BPGciZe25V+HnLdpxshtAaxw03fG6+
S4PYWQ3J9JuQs16qhsOS1mbafH4VCUnmF42j4vBCo7xZBSBb451XIRBa0K0wGRiE
Hqw7g6YjpEw6KZYqhmR3c2Hr5wdkCyGmKd6eYBNsziuNI3IBeQVjwb/OBlBj82sI
cvNQOYbxK9MylkT59D3Cxrl/Fh8u2cotM5enELmCiYOZDYcEe32Mrn5J+RFAOAlJ
KqkBN/wZBdoisKGMuopD28qW1UBzTKGA2CADAXEOHlgvvq1idLHxDI1qNHDTp5DH
yQuv7tXJ/0k9P1ROKsdK8Cur8aE5wuamFB9D2qcwGGs0KR4tdJozLa8EaUUpnowG
8XvidMuHegMnQ7ZyKS9z4R+yh3VEsVj3z3/aHbZ83B9VQAva4L6NtdZhoZm9PIEl
9P0cP0F/AdJhhWSmDVHV+h77WNtaOh3Gj6ERURG+PTIfbByQ67KZ0aI5k+6Pn8sq
jDCQICkHDxuNFdUIYqyO78FLHRbV9WcUERftXbW8pO7F+XIzAJwxHvDkSrv6GvZR
/XZnoJjday9IE5VSuj4DODgqnBLBIiijeQ75iK4tKnP0NSEwBYzK576y8osc7jzf
zgziF9SfR3LEf8q7ixBHOQvz857OM9WzhGAkMgWagPhE4Lzne97fKBz8I2y+XTHW
TcN2wxrcDvz4RPLkC9UnP8REVsneIn1EID2YYxWYeXumvVR/ds11XLMDvPaePWIo
vA0goCI3ZeP+Jez6OrwRPv3cY+IICU9F8BJ+zMGLm5nkWOC3bcA0LPXUZFo93Gri
e3F0btELlp6yFD7BJsaH43KXdbRNXZrT8xNtTsqO3/f9ZlTcUBtOL1ZuDt/yHuqr
eXwC6A/K60O158eR6OaiMYickGp3a/EpdMvkPA49HVTf73AdzndfoHjO6OnKRmtG
ndzMAAsktIQK5FVIq2LrmtdY8SWjnosztBsA5CySGrJyKEsTbkkNTzcUJ/nmEfuT
CLCB4+HZqW8v6Vjt4+PNVV3Pn5MHFJ52ArlaAclKVxYcH9PNjtacxrj7TUb/GXOV
FL3DRHlbkpZGCsglHz1x483emnuP3G7hPcq/2w0ZWH5V/+QppLOobTln2N9bQD6P
dcJHbhG2IrqpF16dIBiz2GNtxEDiuQCGF9tMlS+Te78f2PvNJ7lWnBsE8H4Aca0K
0QNu+QVKZPuKUr2VJ+KvTz0xCaJw4x5wYt402t6OtuY61o6ipLelNrWkvNGyesj2
kq51ZjHOaoNIPC2go5JUYbma+zyWBo/ba8FhgVCitREzsIVAK/9PI46d46YikGWG
v9YdaeTfttgKWW5cuFcj/QLH4NNMlcBTlRUCDMeMvNilXttzcvc9/uiPxtXTVgNc
88ik+2QinzVePex9waUcJQWNoi/nNLfjYj+KH1F70LbgYpt+GzEATu69FrhBOII6
7sFKEp2FYNTAl8Op14ZuKq6dEvBQqSmxvakwg6ClF/1JEEopdcjvNm9lYcTBEn7b
ZZhxGZzaJ5ywZShtbP2yXHca6oCx1tMYun4B1+6wdmG+eu1Xv/yEUD+T8PrCoFsY
QALhHbIdevBfwb9If1b807G8OC+KIf5uY6iiOqtTeTIIZIdLq+dfSLvdyvIX8w08
K+9IMxoFPcBDmp3m7TsRnktCvdbee0kWT/FIbGwgmprqAq2H1kif3KZOLBmMxn+h
OhaNUUxS8VuDCg5WpWudq8TOg18Toovo5FU8687wiOqpFvNXXEewrHFUwjiVPIe5
ncDYhoGHgwdssaJaScfWYERWSe7S4SGf2Saxl1UzSW5Alz58aCJYZoiGXSs6XTUn
6SWhb/NVZwZanLbT/pWgG+VfPj54nA94Sp0yt0WyfS62rmriW1ebTsG593jBVMlV
TLosGuBgdY8Ikt7WCJp/f3tc2cxeDwixXKLQu7hAQqLDUba7PPYstcOdbHHPJ+/L
Cad568+KhLE+1xw14ESBsRmnDCWNGgsWLjaMxb4MN1zsYEEoY5b9/f3ZKP1Firxt
W46VHGOcSglbH8EZ5xHnv74RRX3C4jpQ83E7tB3JU3K7YoxJqimmgyg98Yks25e6
V9YZqF+o+jNlSBC3jPtq3ClYWW/ub8NLoMkH38YGYCi6NWsoUBqh5GGAlsLGrsac
nWSFeNbdG+jVefVsfuiHHhxrH0OtjIppooRBM+eamQzIuFG7oWKzqUF7fAAbXgLM
d6EuD1af9nYrUHYBVAbNiptIMIBfQ1gIJwAkZnZw+heXX067YaPvrPXIuml83du3
eJcVEvk9hWK5h7WlnlaHpTNEGumu+xu45TT2BcY4yjccFZzUCfcQrqwAaDuPEX8Y
6Iz7/ro/MTlr02g3KpzUQz6Y9t7o54Fol/Rz7MEEy/ESMy3NineY0gap9ppPLUif
jG4/UF9bkIKuEVVYEtD2194/6jOdrgMwLoZ1V5FbjrsPSjlxmZ0tPlvaxeTG5BL9
NRubUXLoyWOykWr6TVpQ1B0ObLK1sgpAJ1fSGZKgDbYPznY7ZwLqEzI3+bRTQIU+
H7746dSeRFKo4waOzy5WqkZlHd64ilkNzwcPWePMpCoD8lb99uTiJ+F8w6N+4Egw
LcMW1o9f19LvZSG5sD+cRi3/GqsCTvU4aKPf/s+8xY6Ma7rTlIHrdUeQWdp7SX7B
Kpx/va0HnoXh7zvd5zg6TrHnO0GcOY4sP5ZCH3iYpA/7YnRMnBpQv3RvKiyQX1wE
9riQ3u5Fkz4FEnI42dqZ5i+/vhE9lRH8erc3yEGioRWI6zTeulhzcAc5Ds9eHQQE
RuTm/9/Xr0lUtX2FxBV20+jwphIZCYYyoA39YN7X2OuL+SWDBksZ6wofQAW7jDRk
O7cpJH4WKjHDk67Wc2L4r948iFY8GuI7a6k272sOUkOwOROElX2o7ZCiOFDRj1AW
wpZ5HUptfKxF+G2Z0udM12ULwEO0/+s+Y0s+adm8LKEzmSpyKyDIO7HUIgxL1fC1
K+u5t5hCgcoGrlg561rBQJgMImybLdIbr/iAFe267GN+XgQS8pufN52HFcEVzgtO
AJwaJjMZTHP1ljKdbTML3TtXLm6ckaeXs9uL9l4RKsH0NJm/KJJt6a7Y1vK0SOxV
pM8HU8G3gV1XgkRBaf218ZeoI6uu/Pq2DJBo76MaNuUBi3nnoqze/4/g4DMLAhUi
QLdksJMeaztzuz+cnjAMXWXBqh2NR0XojdWlqP2nXaPNjn4hs7gw7NmWrXCUEOLy
No/sBWrmpZnNbJ8AoNxgMBvVgKLBrmDOxaQw/82GMbzsnrkGiQ00ICPIH/VJsRs1
NHLLF+GmI0pwdpqBRCJd/88u1mfG8WZPf8iX/qyK18ORau3IjK/yN6wdbPDQWNoc
/FqGSD+U2GOofq72i2scbQNC4cvEC53QCJYLVVrmsDllQXVmIvHsZbzj7yC18ndN
N6oAUO9FKSOd0jLa28Zwcco3Sr//zW28DXHtP00I02nGscmw+gXQKPT0aYmfh9Kt
//9zngrFGpLXHSVppfapG8ajJgluWtP9RyX5lV1jFU2zBazUPS4QxRTMrfCSCbnN
j8+HdQFOdGO+zl2gBbr9iXcvEo9RdcJi0kQh1u8WW0w7JFSpqBKPZ4lFg7wrDkxT
czi3yIwe927XHreczTnt3Vk6Kd9t7d14wrWJGzVXYKh5YHbIoi+1NgZks34X71mq
FwiyqeOWcWI+6J2GD2DipKZnqye/T2HF/++xX+yR67j6xtg0QG3Dm6ztl0BlqKag
8INVbjc9V2sH4l4vzPuMiNwnfQnXRFvvapA8/xvYOTNyZIR3kIR5GqO77b6s6kzx
ZTa2sDBg1WGOewEUScKAWJwJENfhhQ5ej511hjWk1soVCzH9HXNnSHpxAlEgroQl
VbpUAvgOGrmFlkHOUm2CYcwxUHP7rVvu//ZeeFsRw/qxzRek0fvq5twEVMjssFcu
3lx0bt7xrUgCCrpU3wWxVTE3kkoHduhLfexzckfyHBZ9ZT0uqG3/xawkwzLFtjcO
2Sz7h7ycKn6DYzmjzf1Cx9HTAJX2A0r+fV5KJ2odUXHAl/dT0kniVQun5As4vt5w
w7HEuMgQN5YWqyaVbZlQfx3J7GCFkMBhLKSGfq7LbXD/bA/iTgp+gqAwHf1UJlHS
SfNYyETf5OpWTo7PAEWtfvFUXrMdMAHUhdxUcRG/bLi9J16ZJ4Ongw1Zqz+qgGvA
WudlpXOd6Yc/M+Axa0Xn58Rp6vJXo4vcVh5XueWvvLabRNm9JoQAjpBd9sd8kwQ/
S766tGQTjpmz5VwSWMtiiMTiJaHQasx5GtbjeWzjHxa7iK3wnSrL6+HKQvlnFsI9
dmhNAuhh9hYUZLG+WHD4Q55eWisLRV70RBAXHMLxjjmTML/pQZg73Wh1AuhZcSZy
Efqwav+Qxp3QgVxpy7nPNMfDXZ+GshQOc0f5iyKUS8ZBgmRJGZnktGY6r6nPRT2P
0t8zdfy56ffg4gpmWjVKHYNkIMWHgGfNxVg0Ryr5BnEj5pMWS7AvsGAl8CP0rgXz
klj5/uD8n6h/zdw3xsCo3dUWjWoSI2RzD1DvyWYdLZZ23JIehDrT+z2ns5hruImK
y5FEGASLhc+q229/SlKyD352HcKsU0AHjmcKMJB9iJsXNSQUww6rLX0js1lgNsry
6qlHy30B1i1FpDFkwBZmHdwMqRpOCCwjGcwJh3Mbnf+vVrH7xe0CziMgiyvNJ51F
/u3Jz5fr+OE7lF2AEArF7uF8NLr3qPR38XxtzIBof6kVhMy/aZFzVbq4enF8KVq0
HFCodwarBfKxZxWOcGwMFMDqjF0MYB28opRDO7Pr+xO2THhPnOEKWUFqpH0ul9lk
InyfYZWw7MgxEZF4F3yORDEbwnTKFeMlzgIj6FrBIL2lotKyVD0o0467z+OqK7Ju
kycoplh6lasaljwgcO3Um8kVhL6KD9FkRVlAichjwjC6tQjnRvclORxYvXX1W63T
hGboXYC3w8gGW99p/vUmJcbw3FTvB5qqDqteqjAPuGayBDWO2+CXnm18kou5XMFZ
OBOKgkxnfQ0VpVCiwu2MH859dUEEDxDYZ/ogauYn2bVJQc5t6q0StbhB3kU2Docz
2fKSNwEKU/YpnQ1cCSd4Oa3tFBc8xxnmBMe2ty1jySp4UPIAqnxQxtcT4q4S00bh
63f/8fPaNcXPSzqcwMtSYKJxKvv+aT2N6uYVkvEul71Uj06jBF/ZZbbYYBFdCxjb
9DeAr2mEw0xqKaoI1OkoXR32h2NhGe1EzdURvRO/nIjvuRD791niB7Lju5cVVqsu
pxIjZ8rV/1NB4uDPVBHNn/akfsyeQJyD8MFgW+cdd2d5HBsKy+dYHswgMTGl+EDu
P266Ndqp9pfNa35UTK5hXIds1rM5gvVqLT6alsvma1GjPcljBac04y8sy2Fbkhow
oeZHxQSezhLgFPJz3Kmswmxfc2wLivvX5zWKovYBxxyuaFwvS3qHRX5TQdPdxFhP
8eYFF60OmjBehBQNQqh8nSBzmRoILtaaD3n6v4rOjjVLZE0Q6Hpd0t1PHnCvskXn
FhvKwaW57l7UatcBb3ngQHaO9ssHGH2cjMOZ7rf04JzpNwEZNWtw+xaVX/Aj8bsx
Q2+RkTGiwkHbvjzI6k8OPfmibhMwL7Mp4uzeenpyx3+LYf5/ZPM8B0X21jD8XKGy
tlEnxSbuIGBDtI1m6H8z2FQXB1kSAnKp0fPkcczfSytlwVjYlCNIVpV7rNdErOhB
HTlQnNAjFO9RS6cmmG6Az9T7Oigp7I37J3M6TXOqwWTDvzLmGe41xEDDQmjLAhwZ
HSd6KgSbmXK8yDi5ZcjJWkNuz3qZzohxytlaHBa1C7Z5ank9EXbQLcden9h4bifC
y5gmvg1aoFOf8jEpW+l+Upes8ophwTEPGalgQLCM/NgcuPWIx5WCwQVfGDl8p4Q7
q36neAYtHrZ1XL0mht5mX1N94aRc/ydRr7c8zBlc/ixtEc1sUD5axJrKMlpGjQBO
FsrDB+yRhwiS8bWA0RbGwqjXuHZoymBShTJvM7CJh+MSWf7bfSGWZOSTDKOQGdrE
9JQXe5T1uXslY58Ht0YShvVvUWxaF/rqfdjcwsTEw331NUkJh/gmyOhk+ODom8D9
7qAsCtZFHCSUhuGpLD191pGg0fHsUt8iv+aFXiRdkITwcwJBMDYyKOsblc4y2/L4
vToXyQhVbkxNhc6+yfjUiPkGZBtvzQGWVv0rP2VPGU0AuUvXU9HaG/Vs8rzzwWur
m+UYdI58pl7XRKvGEHUGzCdgJSknqJ9VVuDTVozRjk9HZO6O0bzBevBecBazTHxd
yEUdjpPIEH6bAQBao6WxrOrSruHtyZzuXS1ZYkU387ukRhHnBnXaQ1kzv1804oH+
EbtjMZ2H9v9XM3kR20u/bxbGdQiIFKWxdYaHnXlfeHyVHONkXYN18XxP6Tbnw24D
RWZVWJ3zoE1gsx14bOzk6B8foTrGtVXjcA5+WaFYsZUzyst2Uu/fF82/0Gd0/IWo
Vh7wtMcwjfy2vyV3Pe9RzPEwrWGVENv5OY4DhvkysHeyUhbzfmsgDUnLA9sHdJKn
sndsgtfpB2twQD9Vu4RV0J1VHekOvvyyVHns2Fk7wzJ6O08c4yaQeH+I4lOMEiol
a6pqXgjF47oBuFFCMFyrhcGZqyM9e19wtSe6jpFNReGKs7luYqv7Uxwqk2InPm3r
aZfll84xBgJc9KGir3L0YnfnSTV0uIbjLOcKpcWpka4TiruA2sBmMHAp13vUBPHC
57etO9PoBuOKl06OD54Mt6vukmcWaLLmjffpvaCYHJObEN9kIj4ZtifgIW9i1BQk
RSRp8Cafzaw09WBD8HqoND+VwC653MnErPzoXfQNgE8mFOxKKBf0nZYd7bLHVl0q
e12cQmMlFsLtv8uaT56r2g0d8INY3nV04IMXu0bqI7cwXrKqFf+03LiyAwOJveGx
otuT9MEuI4TqIe8Ha97UFz1q+dADYEUFWSvn6C5im9PI/Lmv3b0XqLYAAsZxfRLM
7RvvF5yEZeo7psHfzfnOJaJO8d8jSGhYT/uG4T9BZ858RMxkn9JTRm0uKAh1QyNM
4w2ZqJJnyEPTpSj/EQ+nfKWK9rk0XIAymI4cq3R2ui61C8LNaTLLQneZkckmmCxp
4tQkgm1wtON6YlkXh9+166aPOzD+mVayM/HLvaRrXs+3J9OlkMsaquR6kWzvs9W1
9a46w5G2RsLWSOvNVG7VvZLIg3bzEcH95SmipzjXe/ewHaXsQJpPvMJRRFumpssL
/vT6AYTEr66EfKl28HKCGWw5OsUhCpNqObWtGlDIaa+mhyh2tiuOnWbLlM/2nD8c
9vViEKPfWD40DhgV7Z36YYfFDHR1cSgw71JVMH3wvF9JzkR3j3KPD11/+jRJ4hmI
upaMzLRP6OKpcNCLr1UhLDMHGxtcUW94vPravyNc2xyQDDJr/E9BzLh6wQ7DYkza
J0qcfcaqV0K7yqD61hPTNBuZGMlpO3rW9p7LzAbb029o4Ni7xFIrEXf1lsZG1TNU
LqNZaFhC8m2cao4IHFUNpvqFJ7iPI7oDvvbLq0dKmdmK+Fmnna2CvJDEwHbW5Oiy
ihcxPGhHn0qeszNvSSupENoC2DZOo4HYI8awSjGGrCJp5+h6fjjUMMx+M03s7ZZu
kzOlIegtS5G/ZD7SOloscJAwx6D8PyA928lvpoVlaNtbdu0bwsdOxKc522YXTPrC
V0GUAtxrzb6R9V3rP2KUrGHY/5bz7DOEPdEXfSz/dTszPuSC0diJ0PUGWMh1Itlg
60imUdXvMqKeyludumpffVaorAUt2lSw2zX+J1/vRp58xUoW/tDPu7+Cg8ebSBee
hPTM3xWtc2NlKevq/G299bMvIsBlsWxgb16J+G5H1K7VvZCJX7tMbymLVWaeNCzw
4vGo6CBelBlhewi7y6ZRz8axWRA4OQUBsbq2Oi0DCP3nnDzLGLF21uA3TuH3JebS
LZjJbgw74xdWkmOp2G4z3WBPk3Vzoixcrsqpq5blx15XhNVOZME3ZEuCr1iyUmST
r/wCIGWKtUeRmeBEY588XV2U/ldMSEJqsEyzvbuHWV8cP9QNrrP/hbY0fLw4V16l
eqItxjkHvMxkdr/Gtz52FVizRbWDZq8fctyCQXg6wAysQc2pKO1/UY3nBMSkQyQG
eW7/R1hxtOaG5aoMcein9B2qQmcXZngF1ueK0z8Xl1ysjhVr+wEJ++bssKcRHRHE
2SecZSn9U+2BErOw0+qwP12SoCOLOSN16Vts/7KbJs8jO2MWqpiEL5LysNVfJdAI
ee/CVXwRIDPPSAbWmpbGi7O/PcX4t3+/ainBWHMyKdypQMSV6HhXNfJiAkzQG56q
k0IzZBjS3RjetE9or2e8UXLusQdk53tasjJIBDSJwPRK8WukSQeKWLPpVP8dkpId
XOtz9ta7d9pAWGG7TLrgB235BnuADRmTEErt2UoW13210Rf41e2th1P5ETE2w+0o
WMG4pycIdxFeOViOP8UWsl1TXVwwP/YSQzyTSjYfvuOhdGLtDmbrM2qqACcnf8Qf
dmGJ/A/HC+MNyVWSTfONArtYoIZG2hSF6TQKsNzgxVn97N2tJGxYm0E3/Ixkt9FO
jHg53NidSG9LBsdc+Ywt84/YUjNRvGtE07gNTbsEwgQB70Vn25Mb8GUzMULo973a
ZLL8f+Sq0dbaSWosJkJp4/tDwP9r78JyzU9uiP2E1wLHVOGqvlmNagawYlAvkIxj
+0NCrARbvTMMzTjOIav31vSIYx0i3v2CpS53shNapsqpBK900OryEol/tXgU2Yic
r8uFIBmoDcnOv6zuXI1Q9nKoWClBzQAFps4Kk8oBuT4mcVNzuWcqgglA6UpooDS5
5TYqCWtXC8FdINheKLTChPrPdBbO2oHuiDrbLFDh9SxmAm62gUrE6mYQxWTQEpim
rPl3jqdorcfPCdItgKoYfUPf9cPzPXKNGHK3jEuSzZ7SACpPOzH/h0SzFSIzFpTt
uHUqgDip91pwXqf2VpkY74cM7eCuDXUmUnjApoZoyL2LnEgJXeFHUYb+v33znkQY
UxetsgwcpkNSheT76t5RwiM0MO9HxW6+McGcQIQoWMvrTNsiIAw4QC5Kd0/hexqA
Nv71n3zdHTGOZ570XRSrMexE6k4z2TdRAosveheb6mRAr6vkkW0yAY41sCbAlXQp
xbJ21p32dC3X4wGtTpf48xmGAcPow34+CdksNrpLi5RfvxYDgDn9fwx/UyULko2a
rmSK3obJUNowb0X5yNjU8G8QYDt+6hhRfcY2UQc10IYZRNnkXjIVL8dDETb9iDqa
nvtZg4jV1p+tnMf4CunbsWsJEOJCnv5fsotW1J6ISPDDgjXNrML7XZmG2B1GfTcq
SLjvPuSiF0M81B2J/A5zLwZnESz3cSTUlGU9XN2ffQs7eyNSR0EISAhF7yM0jr+I
YhwEkOngZFCXR/n3Z9IkgegfV7aJQchjfAf/nXa4vqRVA84W3YZ0YMbak6uRlbrR
vjAemIw8kR9eQrYhTo8xv4Tb1XqrQNk72JhrNSuqx7JmnKPEmvXfiRwR+KMeQxQ3
WfH2c129gWR7yAeP7qgUS5181OrLphFUkIBqcIYc7yJVOcPMujjA+296V/8oxb78
cFCu/rTki78VFnkuzwvQXptLiSnd/rksN7XGjKkEuP+Kbr9UuWlOcAWMN9QTXBOM
wNKbxEbpCEyaGhOEpMzPeVEl5ZeedLRT3S8SmnBpo2IwASnuNgl/4XpeZP9B4/tX
feanbrR+FVL1b2Ep9+i5ehrTDNDG6pwdkYFbzNCn2G7cN1GgzntZtLJGhZOXO+3m
/iF2tRbFTXvNB4ekmAt3fHxMTTsLZn1rfEn7v4ubJ2fS+T9ChtkI8qfuAdlV/oOP
/JMIQoR/BgjcR43nnjuheaNhwGj2Xal6u6N4VX5BkosKK7oXA7eGlJz5MdFovrmf
PPDXQdkEITOEDx+tkYTw/bWzz9xVakVVPQfzXcRJcVIYf+dJ2oTcZSdfjyQ1Y9KV
eEef8nBcREVNcVnJc6BYBlPSU1MBgarUxZr5bXv/itWAb8HRYvsI/hrvIEOyNYjm
zA5vLPbTvvHXT5Nn2dOeMFqeLxvcbtUnwSaDbAJt/0gVsHUkH1XDDhjmetq11FwX
c0kZoiy/dHnfrFTNpZumRs4YRKEgMUdPoaQ9AM0qFW8qhdw6gWh/OaJwk1r/Zz1K
C1/pTaEeyI9iHW8bqYtQcaobWqqmPIOab57823q3SW5B3oHh9Tt75ypZiscg1wHL
m3L2vnnUymSrR5af9C5sheRyEFgFxBnkWDa21wDNvvdT62bpRun/Oc6gXqA3YHXi
jN57NrHTF1BUJ25d727lzdFcu50FJpRgF6DQPu4UmI20YHrhsDFO/RAN4i3YnaxL
eb7MIhCtbIRt+0AGOp80VuitE6pkZHtQhiG3oAuMoh0tqePKcrkPuS1SlsWbtScO
FeNAd4PMbKfa/qiU0CScWVt1BAemo3vexU+iYGKwit67bKC8Pk7Bqcpkm7p+sc/b
9PV0BY2znbD9SnN//T9q0xVhaZW6AslsHXcPgD0YlyAtgcgoxZSN2fJC4uZEDfFi
I9LI0jreZ6XTlDUqO3vXGAZspqb710n49q0yvEOUUmzcaCcTWMEDZTIUr+4iDD6a
l474KY13UpGTVl+cxE8JUDKy2RuO7elAM9xo9wHRqLsBn1Mq2gUDNGMrKgYYn11I
e+M7bFgAQcbi0oKFSzRuRjd0DSFrXRKYOKM3tk58bKqfEnQ/TkHBqE5GZurfqV2r
WuqLpmFK8/17kjOy89gim/UAvdBrY7VaNx9BDIz/xKb0SrCfXQA237dbWwkVlzmZ
i2PwuByiiBJbwBYLLm1Qyo2Qq9RzDMNBPJYxM+WVnI7MXSnwwncodE3ndHcJGCR3
aUlREIuEGjvlRYP11AyceQqStY1JaKWLuO8Y1+6eovsq4pu25qmelHjrM/PAnt08
KpIgWx6Rnhjx0Uj/DOJ1/zNKDWfhX2b7ZEJcWWDcgrFAqQq71SApCSW08Sl6OMt3
HwMYf12ZVYIG5U2Ezel8U8vT9VWXK8P3qqKcRHCMUSuDbf96dCHGLWtS/lZCeSN6
3+ID/I84ip6RSR211PNIR0ZAvYNQvwkfgKv2lVmKZwIMlszIqxK1x5uO1HZmrMCa
HwwyhCHTdUDIvw8KuA52FTPvrjPBaJKlx5pfeIJE6yXVvAbpGUCM/yYy6DEB+j3/
146b3e5mGnfrg6rDlU7RvnBDTzuBVcU0UNXREed03nJa/FDU8vmrP8KSUqLdO1BQ
FF+FzsJjQe5pCpM/3xZArnzCG8XITFEdUPNsgEeWri5fdQg7b2a2hazYdBkcPC/M
0iKoPmdEcbf1PBmUUxKDu3H86f8V9xReVaiQC6x995+68FUJ0cInSt791MaDqXnW
3QLxHIAAmH0aQK4ZYxhCm/4HHCCbP5s2181VO9c3/mi0rHzUZGrGdxzkRSQIFl2k
Ia0L2RucqaNsqQNj82Ug2i5i+hcwp7z92rSE5whYeQTMyE80iKoDjef9d8jiinIO
ktPC2aUtQj9bbeK72qCwW9dUUaJqp+QqoquFCSCqBsqBJNFlv4EvAe6lyOa+IGzh
zQYJuB+53wcZd0T6p1El/oOHMzY/JM3jziv3Eo3O3tJmx7x+zaC6y4Ss4zaxqN9Y
KuCiI2J3mH1DC8cUcXMwiYohoqEsRPv4W4JtmhilKYNjVDv6Ssl2iwJW00yfVmD3
XsOeRMbR3FzU7S/XDpsMrmMcKEFBIHOIQ3WdE2Rgn1dFk4UQF4qAi8eiJL2eKQWL
A/FyeEMgSHeRqg5pN77caZJtjEZ9um6qNg3QrkWKn0RqxzCVVtb+qPCFd5fShyYT
1i+klZiKnv+L71hikU1LosWgbTz7tb26fVlmt3r+PaaOOx1rc9s8hW+eatjlzTf4
hqzGm8OV3IfOo4axkqUgXPihRuLRL87rD6SIoolnQHYvPBFhdF0IXsAtQxDHJ6iz
ASW/Puk/NNC0L2bsrVdKUzP08A6fMNmT9F4Rs8tpfrk6t3AlM/Qwpi0+jK5HNysi
GOjvSnL56UI+jv8+cZ4O0STLJ3UtxfDoLGiI7auUPbN3oYYLCRiDDL7A1+iUcVBS
KgOy7ws6VM1/O4JB3VD8K4yObgvtmE3V6fPIztKvnJJcbVXdygqp9qV/bJoliThC
RmSm2Gyx7ocdIF6GxznpblXefzd1nH9k17uw2Cn87OheVuNoAMV3Hs8JMYIbdfm8
dXkD92p41tDtZOaG33W1D6l1gDSqmhigfPCZ9wtCj5VTHLrZt6H9HyhaetYDxj6P
Op7unaHzm6jqDKBtfWK5ckedBVZ10ZFyiQM2mfvL3WEbAp3qvd63WFT66ybb5TY+
Sws3R6C118//LNivdnZFQWUoSF0KFEGvwgxRf+VqB1YvrwOzaLg/QHwyW63E3+2j
YrB6rQI0lWzlRLs/6wcXhz562exUE+e42jmfwgg1RnYzG53auFKJH0RE/otVMVG/
+wZmPc99mejzEERVU5vnBJHMFbE9vo8qS1/jSeJmi79MfHzMR05wh3sGD5c2msJE
31eNUdoofN79C1L5wtJaALGq/MCezbi/SncixhrPpd2lo8AgbfapRFD9JM4Slmkp
ZsaoRK8/TxYD3R5LEDpEwPar0x2hGOJ4MfT2x8uaUqUz1oSENGXq2Qg6bRZVRVQ5
WIOpfVUDsdpDRpetBX30zKChqQZINrTpfNLMKO7ZEEEpPaf7ltaQ9QRsHNBN2fGg
v9K9JUCeKRA1noXfolqn7gRbI0SHDHaKkdlt3otABF+fMWUEuneYc5oQe5vCmIqz
64h8VGRjO4hN3auGixVvdmtNvZHyQqnJ9VDtLQExOYyyS+5xvoufnEEsdQwLRjaV
octWQu9yBOm2jfq4WFiPJaC0tM5DExkZszBba+TtnB6IygmlTDtfG2A7N9ukv+Ro
NEyKUfjdcYokxcsULr4vCBbmgEncgzMEsDaDMAveTrkavSE+QB6FH6hckz4amz5A
der7OTMdlpMgjrK0/I5Mj++tbzQ+5kLve3kDvgXOaFYG8S5pTol/bNPai49JTbq5
kerhMC7iOXqHmyGwUZ7uCBa+opccy9kLhYqItJL+q16WmmGr6Caia5gDfhQitzjV
WWF4r42ElzT5lP4Gl2zhwYzbtyjLIXoW3Vo7PPMTU9b55vs3AIO9dRYPW4Zh83h8
GAkQ50DajdPtxnxns7dMsRfUHxY1+dwCZdEZeY5mM8HIs7hsWSxU9j0r7oF6J/+M
qGrN7dZmKWUuqcK8O3WySkpJDFjj7DyF/dcXTxRP27Ft4GeTJp3V2lsLb5hZ/Ter
XXiePX3Ubbw48uTEL9vZEx0/BaOHRHv4nlqu3xab0RqIRmTIdTLJ+5sTheRbB3hs
Ory3wFdtMy7Ein4Cm5EPhBPe+vfue63u8NLcxHH9QOFrKrhajq0YB6aRNsBDNvR1
BVgRCWvEFCZIDavfq2nW//9rsXpxJqoykAvtXbJtz+n6mzPDZKPcVFWqzhBSpUW5
wUkl8Dsf4Nlb/hzPmJ6ny5w/PDA298bjh6Jzkz/byC8ecIvznKIdMhFf/lpTUevQ
WmysYRDySphmoIc7lH2Kod3qyVOnZWt15QAER9nnodzbe0Nvw9u8ux7CJv5arf2n
kYOI/n5yRe4li0F5Ch5dUPrn/rtrDItBUXyncC9gMq23pBd9CbALkOl3TfnU3Pmf
qmx3WNOu40fRyIp23EskYALDPyTTeL04i6r0Yd5v42mRmPQvp0G7OkQrjccDX1ah
Ty7+qmoOSDuCYpZBTZJyCRFbbRsumeWIwfsKTBe9CV3mHOdmkCZ2wDH/BYkd8zqH
lYnh2yOT6RPtylhzpLme9BQBGAoGppsk21Qbm0NprwoadlquvuReI9vEO/pcf+dy
3xVbKfYUotckkO9pEqDH1GpeUiJVCcTX+eV/iBaV3khI77z23PGcdJUVIbegpRHo
YKhu/C+hzy2OJ1OU8o7CmY1JbEzkaa6pesg1REE7ePEJ6OCCqhipvLyRtb1uWcuu
R9uCzylF015OQlbtg3cUjyo0jvVi4A0joMvi6BpV1yyrV8Go2oMgxKD+XVcGxcM1
MSpO4k5UXhsFBubce93ysenUQMhNWzMX0fV2U+nV5DSWuQHw5Ctbfu37mDna1oIg
QENQvitnDA+Q9xfote6ViTZKFdKBWvWomW9nIgjRdtHo9roQZyhpT+rQOjIzsg+n
nJovCkwlret+EvxTGHTIl4cZV2WZ/4LnjDAaw5UxnB5Lgx410E3+9nTvfX51BsrD
aBEpPSpgLFaJHsZOirjDPoSepOiUevKTSTVMeToJAJCJeJdgz+2A8VInSMOKuFWu
aNmKMEbkPSGlawAPyqW2ravSuS0SQU7SwcSFRXdnvUY81g5M5Q0/pekEftz8h5rh
VG3oJTzRWQvEXfvK+3kUm1Af068CCzTPKfS1TOFd6cKqg3yILvpdIZoItGo3X6DZ
7y6iaACFBONbOdxyanHohk0JC4IBSAWyWgamN+vXdhS/XuegmO4XQu3tmxxuHacw
MUF3rfzmFW7VYNqPXVPmLtKqcwajx9DUr1Va33SfVX3R8viiBk55BMZ75ym8MePN
sBgwFPB44XvfLKoNau7Z3Er8WDjfXrb0tlj54NnArgJjJCZY6Tr6gO2i9GVF4UjP
pjashyf6dX9MfqidNXlosjqiqWQFt/DQSeohqxg8XdRWuDa5/DZbU7MkCFzlzNET
JbYhiVG9faoUDc5a22GYd5B2ipbbT0SlSWiwQm4xOT6VkGxhnVKRhdxIrlJFYiFu
NnHCC11ajxk/0D9dQGJZn3siAkYy3bj2LBqzOCDJHsCsT12muTuWSNe+QZhCk8iH
3ivjHzkATq44xKUunFkMmz3cFfYgVNwbw2SwoyM5ydHAzOfSl5rMaoO3LW1AI/G6
eIerbTdJ6ndzoIHG+l+xbm4KFRmyohCbR4HwJjeU0o32/lD15+Xn1GcjpnQXuBZh
1Tnu8POwJD91Wg+xs2ShfpM2QmAQWRTqIWRU5iFb95ZGdMpoxhxTDjpYKHT/MLQb
wVgPKb63xcDYzFtl3uauPmapWWLdQyNoIa5vpar2KPVnNojkEhy85ZLOC9cLpPwL
p3qNmrB9w9dFJhziyZ9lEJasunMwavEGZOqjnpb2rfrhpLZGJowMFGoGmw7XNrVx
5eIDDA3KRAzmp2yIgfbzEMLQ41l9PolpAP71/vyNsKJc+6LThAhTMZX2JLUMQz1N
BF6uancZ/S9aOjN3QATIfV2CyoArSueygjhrm2HXOJRo4zzLW2xd/DxLhebBvMtI
qYP6L45G6/xPqs79gK8Zd04eXIKUzvQP7SwY0c0v8hti2DiR52csmYHQosj6Wxti
iCF8xiQEIL+jThn0gt2cpdqZA4BF8MmfN4lYWEzVif81hnJoZ6LHlaT9tPkJLMqb
pv1UqSrJzRNN9X3/loXoX3THqwLG0h6+kZCwREiUpgpzG66spx/eaEvay5WYbxmc
9IxiSMpYdfF7WbfL6Qlo3fEWaDw7TP7slh6xTTgw2ViMUsp60L0Xmu5L/7mKaGC5
Gh/mwM5QZFDbLOHW2y0ZaXXXq4BmncSSLRwdYQJnCjUAXQHnIm1jdmAvtdKPzGgs
xQirpPbvvzcjfwIvKssVFJ5h5JdLTaoqF+SNbwaNAjfoS7+22iHYGVRkpER0kPuO
vWDpFx3V+Iq6O7zqJAVCKpJWXWHwWG60UZr9BQbTW7By+QW8nWsvIeGQSgDzqdf2
RO6tBUkG8hSIrFRiPvEGNSPy+YUnB/LyVggfaxzDjBXKnHYGEmdSTl2gSldtrpEz
ecAuwdFJJVn79bF57plPxP3FlN7fHqxnvKoyZRzBqJZsjjYz9V80Fe7j/0Poomq4
mHAEvsXxPv/238oeFOUAW2VO73Oj+j+Lf0bI+xxtw9cOMI2Z0YmQ3P1Nkj50UKp8
qzktNZyIRMIqCQB5/SH+D3zmvVJgoNK6tpl0T7sthtGLBUwZwDu8zihSgwV0q53h
2bDRdeUpj9z/vDckQ3v46Y8PnP3E0RCoHhpHD6tp9NxWSmltp7Wgd2DfC66QkAOr
G6VqsKo0MP2f3Wx+cNw1BNfLxRINXUv3hGLVxhJqL+Rt2c9lFe93lx868+jCYTZy
dT9+rhlca0tScfwz+Z2P8jTsIc5rp1/NSzRFUbhmcnffoEYVz0erlCoY139e52Wx
D0VP6c0wUeQzTtO7FGFDHWDTxTvxMiu52zVuYwQOEzEt72zqA0ZSUsN3nLsS15Ep
6xWx2aKKErSu5FNyuSsBt1VRbpiiVvTY/+qM0Gymps78ATIYD2jJG0+8c9qNrn+e
jTRwiHXmP/JTbKPbjl5qF1Q6W7yvvyCQsoeHfG/T9HFHnQ27FrlqtpY1QFXsjQ7i
nR8fLmhRULFqY3LJcMV0UFdIx/dL0BttLA02jfumUGsY/1jyTFlFuzW8me2+NuLJ
fWyURFjLl20ax7cnBL7OQOE18IDetDHgUz4Y2FA2xpqMJIgTA9hroO021z4MsJyZ
ZVCYa+L81qXZCJG3FUWEhoZOFExCB9M1uoc4+TrwQ5akbTTq6EIjR8mOigqfDUeY
KG2A/6ZI992igd2BXJ894/taSaxxpOR7EGU560uFQl0U/E+TeWwY9v0bcWON7d3W
8+GJB5+UiVEWjh/b2+gxPPoY3m3C54i+wmjI/bETc4JIgToKvJQ8mv+4jPDio+Rs
2TX3WEpA605csR8quULLy508S//ka7wq22NHxOcL9lpWfVYldp7p4vpang2aPsti
w+EQppM4gkIEs20lDxWcv6iEbB8Ws/+O3OSCgIvx0zI1T+NssnSBjENODhQNgTko
DyvWkV4UQGu52yV9ISuCrZsYDVeTF8OMLpisNdM9OwAoElBpW/kdCBIMpnNDurZh
+uPWGSRInYC4uOLPlcOYcWqitnUyBTATvO45S+5ussblixxCvsxzdyB8CVNB8mNt
iJzLCkHptP2HXfF76OektIPJuAXMCJaCV0QUn8OOy4PnUyQWY6UjiMqJTUSxGC1k
ekoC/aRvmyCDMmhZfSi6VLnUKekVS/PywbfZfvDm+3jbvqrYCma26llOzcozpZY5
Jtfcwu3OA2tbzux/gg9wGbuEaFwdxAlvcZASrg0BZ20187Kce0yVTVeOr4RUTL1L
B2pQOHZXQYV7uZwK9uDXWqIXXF31PiztkJCUPBOoc65ySczV/h1ltaIxQMwynUmx
5hRvOHpdLdJWROiTIue6c2Z+MrLoY++UFeBrLu16gPh8+PtS2atgH1juekzIuEkb
g2wzqaqaYc3iPOBWBo/8mXk6NhKxA9/FhjmKSTts4rPpL9+6149WPbijhCWufvhQ
Sy2RhdM5WhJrpAufOCi5TZLpuQ8NZ4ZFtu5LbTjRpjJAiyXmP4O+wKyEj4Fhv9kE
qOYEL8DMMnd2V3P7FBZQrgApkg9IH0+gPpPD1/glFbWBWIvVkXAW/pZVV/N+1tA7
1W5XsXIzaU3fA6ho55SFxIrNE8rL4Fs94Nckauin5h2qzA4I5g5VUfZfV2ekLFgo
GqcB0FooXldLa+keacHaYsiOth661QEJA6MgjAacRj//N/sXDmiCjORRhMXsUBT7
x29GCUk3WXwlgJJkAMTgmjOuDqxB1rh7JzQ8HlfpIXQnZ86FGeDwoZEEaD6Gw8j4
XdG/ZaGBh1/gi4z0e7uNEP7MI5XqrzbxTZp7kJQCGrCbU9dOMZs9EgAmqFpMxs0o
gG2q1XHlh+AbpbAJO8ieHvDssyGxQEZtlOziqZB+12GAiZBlS9FtvGxn30uZlY+6
uj/C9xJMflK1b+YJMMR3U8l2Po/8OF47Nvly8ziwe084x+2rgxPbturcQm7Vgb3q
ypOW3c6SiBmIWcTm4GZxGT3HLyEvQYg/Gm3DVO+nodyponTL9+URUxED/0oeTL2F
jPTK1kak9mxSzcnQf0tEyE77f6RvuapUQvesxtKIoGmp2Xgi6svbNOfqMEAkTpcC
k6vfcjBx/Xt1MiZGqBoJOfVa6024G+Ii73LOBJhCTOqKFL+8/WgQxZa9jWmajFnE
EhaWHs/iE043fUdmUVn8MQ73LPz4bcCRtvWCvK6ZT70qr9OLRtxzneJRozLApKPx
nbFKOrdFlBsQs4vgzMNKAhBcQOSbBYk5GeKdKcc0WYYH3oS3KeS0vPnDANWgjH4G
J9xh8ibHFkGFBX7TB7sHIKJk+ETLnOS5SNW7GpqgnYkZhVoTuu/UKh5Q6CN3ZyJ+
PxrRwDHzR4MMtKf7xDRaFuab9uk7sIukC5V3lfxpbqSWPr8150O3qj34LxedDk+a
uac4lfljQYEVGBiqrSqZbE7H06e4iy+/Wo+NDpb84M9aGXiKvgK2mH9NwEwz8ilw
G28FowtM+29SIE6xCT0IV/ppxJ4YdYEnhPlM4XZCrnslBDAM5YSN46E0YuCsXJ5X
OMXO3ZvUUFd2sNXMjzLJV7TKjAC29xWuMyzerqv+4n4Ql+/xYaPZ7REP8lDCDXkx
/OiwIlMrlwsZKx9setTJ8krTHoFRU8d2mFK81qFpKdmmxoRSMjIaxVfQr5FTVO3G
9yi1XqgQZ2TIP8sWE7CgUYzSZcpzO1MA2rq5RzFDbYGmO9gCVQIowA2eFraphUll
86yKStXT2fy5k47DdlVWqMhWNYekPzKGAzRTkYSPee5h46tAaRoHX31wHUwPQct5
usL5bmP8vAj4Coog/iYsQkcWnuYcRaBRVP2JP6o+SkwrHUj2jniupMA8p2h43DHt
rrrGg5ZcPRFK1L2xSnTQLXfPjl/gaxUs61f/udgRsWAnWMMrtKbRadK36ZZqmvMf
kPqRA5B9N/omnY6XhcsZHd89H1diULD74LgGCTbJW2LcmddEjGr6HXZt35OKCkMw
amv39JE2M7DASv8cLpUxzeaU2i6oBON50EwGTY9ZO2OhNp/JrCoV9DXB/DtfRnoh
6lJRLAuR9xhQ0inxMSRQOnQU3x/z9/lzTIzUDqMRtGS2fKKfCsQ8GEeMb6+g4+WG
Jr7PnPyArwHU7aH1AgoO903AAVVkuPrVdmef3z/ibZXy9NdVWYJFjeEJ2jRXhXPv
IlRvPPu8KikN1yzE/Sh05jdOV5nx5fZ3OeKqXnEcXFH2Hn82CY9j7DTxoKgQK1eu
UlQgpHLLZS10gihjAtMsJ5VfKlQkRuoMQfN6gMt53ptMwT9NI0Zstylo+GPu8YRO
xW0Eu4DmPeR92h1Ehj+1rZZbD4frwV7UkR8t5RevtHFqUt7QK9gEhzip23ZmgwLH
esRIF4Ulx5ZcHJPMm0tpS6PuwNbVE5FUmFCedG/1rUmewz3FR2JmXjzTJ/1egoog
y4FMyurJK+vjK0wG2cqgmgXr13TqcYZxJnIR+B3Xo7/aFHDvZnlZ8GpcHimaZ+Hd
KOchi/KxJLLOhLHiCbloS4Mq6duu6l/nvnFEocPxZOvq0TgzvF8g4E9uj4tu4gsV
zSIZtBCmzr74rq7CpHhXpeWTIyaMfCscjsq8F+UHI/tggeGEod19ouelgzP9VecA
laQvtt329jslHS2UjEUBG1woiNffWgiJ5zcI6KcN8PmmjGR5TKzVbTHzoZFKDkGi
QPNoDSvekxTp5UoxBthZqWOXv31P752hkEW1gwgJSY+eNx/ha2sZ+CQNp22lhAhC
flbnIh+6LzaPbVeaIkocFpyq4v+UQFPH8tJf9luDFd5cy/VMZU9tWjJwbHAqcS9m
Hk4cKvYYlAy7vz0mM1ubjAAGbBT0CfXKc6lWuP3Uo8+zL/HAgStlzoobMPWQe/eC
hapwCuwA/voDTp/sV8kqSmDzbRVedm2OnLUrsIoJMLdnCeBza18kUEtd51xAU/eO
McRdOHnsTtuBp18QterwmGvph8mTPgmzHKnc4E6wbQl97hSdNyXRsru40jplaJa8
Nn0d9p5YE5LRnYb4UwQkHgvR8djSUtt10kea8P70RMsG0Z6Hg/iRMNoREAHLEmxV
dNeLMhEjKVXVsBmR7rdIM4NF4AXmh9SwoKN0l0WnltOm+kKuTXJN47jh8Rck+53F
XPO+N+mYMhUY5V3lKlFxN0fh1A4NNrHifr9QjonQ0s8SIuK7Ta22SnD6SFd6DRp0
OK3ZKwK0awCNh2u3g3OQfri9I2jxNdj4t8Ro40mUyzpcy5xuTgBBrTqfJqZsnLmH
jzE4rSl9cXRvHQWIZ9JIm5GppOzzV3QHM5xYcKn8CMisWj//blnFtdGdvWVFDGSQ
NFdLqMGgVp7Gt8l39V6k/tNRteVG/zz5LHxDWnZBuDBP+eL/Eo9abOYNvvTqpg7P
aB/3Xz46zaM5DIv5qs7NhpnrQw7GR6YSO4UvKu5sH+0jPFKIPtd80TYcBz67+VEG
9VUaVcizS8A+5plvkdGiayVghIxKiFy/nCOp1vvz25X3koZOQjqykFSTIYGANnfg
dcWAACVWWy4k3v8IHx/4q+iXzBnddzo6eyKzzL9kLXoT+DUzgVyvcXHtqOc8Wni+
qL+iIsQ1/cTjzNfCocTVqCbyIfP/9xmBa5Xjlk7chzvb+0QkP6mTiWLI6NKCQdfa
ntT68+OiHGeHbrEtlN9mVPSrSB2LBHzDFH+Ap6mfnpb5eOGYy+D3dPTKIkUnuKRU
NI4j40OHJyReXymQGs/GQt9qU+qt8rIetHjXUDVhxoyUbJIMagdpPGDiiZb11b7m
HSGtYTLLgjXMFk7DO8wtS98PJ8fNx4J0lkkIvjJgH0MElh2GFfi3sPFYMLKdNaji
0M3M2/6vBS1Zg/3C5FbYISy479aYrQ9DPuY8FhtB8tyFXfFoR3uHmFwEg3CyEGKn
E5oEOit8WIg6No1c+mtFmwOeqha3qwMrRU95UCjboUHiBMI5C93goAXt8SA0xw60
aH4g7wUV1tkC5S1yV1eJCyhVakUhFkHvr+zqyokUOocwwbA2wakXVoqWKNcbsw6n
vqTkt71fSQx+Ir+qmdzcQEsuTnUw4Q56BN8V5hkO+TKVn2IE290qZYNK+HplWK9p
ej7ovoodlR/tyuVkCXHwL8IHGmhwyJM0Eve+UrVybsebrj8M1sjEZttv203ElO6l
q40uL0YEbunvNZWlAvrbtI9kBAW9csvoA08Sf8Nbhu2r8L6vfkDYwn1XEgv/SzxK
lW1OlnHWMFxSP4xbbLelFgFwX9FhBv/iKQjSHm5aWi4KcxU1/7YHmMxmy2BclrlD
zJ6RFRTsMSR2kUgomMuJIS7ZLWGRo6QM//F2hRoTUV25rNDSGA0njZV9+XzMetxi
LJp5Pap4ik1fOYVO0VbPYazG2FlPzHNUAfF5CHOU45jvAjEb7VVKfl/R24aQqFBY
3hxySIGUPiUo7RnOd/grScomkYvKa8+v+QIxUHzMrDi4s4zwLxH3V8Wk78+Ih22S
/p5G8+F7HPKK2XrSHLBu85goGZ86GloDVr2u1kKyr6IATGXsAlv4tZ/MtZlEFuKc
oCff3+vRKrkfR6zhIvMzqkABPLgI+c9fryzhtKv/2Md454ZJf7Od7JqdFxP6lfSC
2xLF5zCo92LRy0udA2CEfeU8fmEW1viWHTe5bDeo02hRT9I5vtO/CYvESTyY42LP
VbUQf95YoITNnrLxIfi+pMc4dKNpWjwY9STNwHjPBa1/JqxAHPGzFPtJQbOF7GJl
iy8Efu1k0t9Tx4NTgEIqxl0xqHsx5rkvO/XNBviqAD0lfZFwslSOCGk9JeBv5UrI
GED2E8SBU99JW7M173q5M4qOS9BceqTIp5uz8GqzXDUx14ToTErljvs0mVjrnpNG
lmXusgecid8h94U63BLe7/CyKRqpNt5dByfnu6ZS4+B81hTQEDXEu9dypHBWtCE9
JuJBsHYr+45z7XeMQ1/oLDcz62+qYLP9K4DBjC13wTnptgdRk4VFu7EAWR3md8Lc
byc+bXjnjbn0tC5wqvUJ1jA+s+lCIw0fqr7rAe0jFp5ZJxDScL31dY49PaJTqabs
sbd5cK29kK7JCn97GT20apKqQBteIS2gRpVesa1uIb9E1Uh+BOv8MofCB9Raj29v
U+WQjg1ubdP/+fUCfkPbpHgeMqL1aTX95sycQMO6vpQ2A4aWQVrTY0yek5fTrIdb
4GDswZgr9TaisqmVXuJDZjJWyqjAH04AHFopI0z2yR+8zOw2Bf41mbeM+OECz6JM
WYzkC91Jy1NhNWSBjUt/1Q4cAvQFwscbsGxFbP7TC9RiDzhO3BsgtzvL24/6g2OC
WwlPE33yd3xBrdT4vp5MKnyY+7tUAIjFlvI3K7+xO7sx3GxksXhgCP/u8hMX4VuV
hGiXmu2Xd6AZX0EGerwIR6izPNLy4LF8GphjitZT2GhjC+Sqi2LBQ5StR8RMovsG
ECPV/7Zl5BpVC2tVXBodTNrqro/onratJZVENK5xXT8dvhB4MYoJaRI8xnHYgspn
fIrqM5qyHWxz5awa4LRo+FoAC0CGKHj3SjSfNihH2nlKC2wh9PUFCUFRc3OuqGev
u6A+lovyXjYL+42Y0FM6LJnyD8g9m9OL/yrVoDN/SndApzXy6YIKJjiNN3qoz6mn
xzAKtLkXkiNkodUJ3rD/QUaIBxXv87eeJB5n5HeShcYQFWQ5s8y7hQuQjAMlxbS7
eQ5iWKoi5HNcXsFklgop7cv3xqoh4qoeakgJfyu6+oLVJXxFaElECj7friG7qbiR
TnqbX+mxBhn5aRss+6pJ++FZMPkbt2+ZR2RNbqyuIB7y25YP7cI0FNQVu426/4qU
d8kkgdkuRJ7hLqz9XNgzcXSNRY69pfAGm3/iJqorGmwqI1R+u9XIBUdFIrZcCV9s
LWwHBaz0H7TCvVT7YEIgiwlDV7VuxPwVaXyF54IsTvus3ujHHUk/eiI3HJtkSDA+
S5r7jdcUly3O4B4JRELlxoU5Dm/0KNd35jo24Y45n4OONO5Z2G9BOwrnCgyCsVTC
eVmJxZBovMIO1whJ0cNhRGALgka5xWZLeqGcmd1tcUDjr9R30to1kbHDfGc7CH7h
NllkqTGJ0W9+2STsDlArQVP8WuoFUZUqagLihc3zM5kzTLSkqroAJ6ucHfc7wT1Q
yoKPf5QLwMlWV/j3XjWOmnLaMYN9+pZj19xcQJjMzoz16KymXj4T4sSVGZZ/rESO
TL4kN5SKHRfKe1kzyWvGIcV5ThWThYRzXjDBFutlqmo8L0v5MjEGq9IrvR4dS/h8
8HBSMoIeD9g9wDKcBlUphDjseKA5SwbN4e7Z3mrdkW57fuc2jm3mApziL8j09qLR
cEj9mFyzeyuf+ujtcm8Dkn+e5W1qBXg+BHsH9mZBKfZsQF+JBuESLRN0cwLYgi9F
xojFMfYAV4pRw9sa4TqF5WOm+JkqvZH5c2kyf//u0T9btJ5ZP93ex3NXudbSsU6e
lYkcgFJjmWqHGWmWMaluZytW6N9968mzhqRgGrMg6B3IjeeH1mHLyTdSIC6V4PGL
XA1Hv+kXopQQ62lpMQoRJHwfY7L+W4bBpnuHoB543sp737HBbDBKjOIptZxCgQsk
rsb0pu1FiOPXtuyl2DutWUQu8KKPBCKgO2dMdAVfVDK6K31DaU+QADgo/9+ptoal
V4MgYTN8PctnYKacMrEM0mjVWiR+tTCrIQnSFH7BDGTrBEVTXTIxCMEJuVnICh6L
im6pKHMKxU3lE28xrEsZFGjGj43/HrBNKLmh6cky1PpO1AVkPEm//uLmptqiLgIF
CrqE7ftVB/JnpxpcjyJCTcLZfWj1TVfol6g7UrzONRVMO5+1tn6R1xlSbl0tii02
NEQznK4wWtoDV+HYivPl1Dc+2EX6PW4vFgTVs2oGITKm2b/hBEz3karbH1MYs9Mi
kpM5swL9UT3SY3JOJrZJse8x9s6yGiociN8laWaz7a3BkEhn9QKWwdgrKNFxkTqC
DfVpVwRICpBf1ydaTLpMR6kwlzxCf5/Wiugl3LWiluV3UkgiYLwe5hB/U2CwdHa8
Kfeev2tgH2RpoXeW3MEZ2IwP27JQ76umwvaYe6HX9faKZCtjimeF/5SnG2g9pRDl
QZAl/c52dxol5we5G4wvYuyltxL25tCMhlwkVn1gihNTE+knYAlybPo3iPBlzZqE
xQe1gvUBwzbOnB7ZaTklrtoYRtxj1Znc1k3rGeUuMRqAgm3FudD+DZj+0npUVjjU
DwSQzdsnoJ3OD2wlsiw2/qhMMtYq4bh9L9xaxyLV0I3bxWBTxHxrWGiF0OjyC+bJ
SGnTHDXEFAHHY2aQOXNHlTyOxr8CFuOZcv8rf8t21NVLbAFX9WrGTXzLgtgfS3md
rAMwwG+uKJvDiEhx8iTY4yPQuILKXE8g2N2nL5uP/LKy+NeijFFz90t+e1ckox1V
s57J/UxiHHPuYEJBmcT94FfIvoYChLoF0HKwsHJdK2lbDorGPDYwUVcoffAY1eho
ibX8HQzyowh4749wt9n40cSiuEW0OV6xqLKXviqI2gYCw6cEB9ADPav9CemnVgdg
dsGudCD/Hh5AlWq/+YvJPkX7iNiJlppmjzPKyegnzji0UxGDG974fKbHyWg0MLtG
MA7ROZAR+OcQcvjlzlET2Gc7o0FFZubMd5WtSNhnyquuYWTqVzhwSbvviMK08J+G
w4VzSR49GL1SPXB4Ui4XXcOVP58MgVYkEvdlbpEdOaSpSplJEs1r9EzgA4bxBqYj
XOCMqjwFbwnpFcUdnxwNyd62IXEfTrzV33qzJ2+72L/g9CYMk0NSNRzsArkGezyR
NrrEhc4GjUoGCRB8LnZiAsPfSOWpTPS8VgmRhRDNNf7bvZ988+VjghhzT6M+VpqQ
YWDx2Re1lv6t2eEk+ZY4PdK7qEJ+WZTHpI7zXCV3mTvtvSDmrs4kfbuFIM4PPJv9
Y08fj45hZslX1b63IE/v7B/7Ja3IYLNp6u/e7trG2drkZTffvGLLQsH1Ajj9DMEt
Y4rIG/ULWFbA4OgCfr0myyGGb8XcdlNcmLgiSXphTwLPrv5dC6+6T1AOjnKf42iH
svLecPfjYOdSMo7Rl82DxeJJ61MAiYW2PrwrwiDzJqNupXufYq2FyeX1wq3uLFYt
olwAXCBTKuVovK63nKGIipYubjPpRzAy3VqD4KAACpnTNCj7s+Njr4yMgWhGTRuX
6ewQ5U/O71EHRnG0AXJyZYHnoFdcjjWqL7JJZDmm+0GicJyya7kEXniz9pE2Uwwv
TNuw7eG5PnO3WpDBffZ+BsWTgmiKaGHMH+gTuVpEyxIO4Mha2wE1qx9kTzNJXoVL
nC/3lD3WiFMv138clc94kcnUaCZ98h4r7SGDrv+p96vUWPYug++eb6kgN+AV+Ntj
BliAzp0LUVarHDYk4b0hf8i/95ISHpokQC2cD9gwK7gxyUW9PGa7dqYiu966cw4x
gtkL/A9KpIWPQ4wiIr42fpSIOs7moIvNpzkvDZT85lVpn8sVY9rvaZebUg53si2N
fu2+39Ej9fbeWooWEyCRSQfwqutxkzYK0ZyKi3qpxJlxsQ/wLNv5vKZ+BpXUitgw
pt7V/0EkJuVB7fpRrHWkDhd1/3JLapv1WNKYirJkzQSfDBai1nf9D8WtGy5DB/aV
670JK1NQfrPqLHHH5Xv9WVzBzF9lHYOhcPyESn06fEApBsFUVoBw0knApUYiAZGX
x3uYrwamBnVJHdHpoEszaEjVaQ7uTIpCEhrsu7ciZT4+9y6FNOrlw0MGEPbgcsUJ
4Q/6iWyccUtcgUrqsSJUgEsfN+PiPpd/+6+Uz0I981+bYM2OloxlT3ghf57g7rdU
RjGjLCwJ4npmOOZ7dQ0i5EE4KhDB4xxzKKR/UTjTJQ9nwjyBWO0aFIXorve4/AV/
/FK2TCAJrQeSvprRj7UZJna3ul0Y+ppz3JtDfSfnZBJGlBBzaGOyGYhmgoJcAlMS
GiCF9B02QpXRnhNLzf+N/wjBXWiyT39D0CH/YifYowjVPcXi2lfSdFrpauI9ghhc
XtFyVOL5fB+AW5fFyWfDYAbeGYEqNVgxDbUxDGZBYqvsIZgivtFdeZkhqfr7EWdy
UiTRf02Tjq6b6x2qwYOdd02ad324XMk//hpt6MUmU3MxVBKFGO5sX4nYALcxmgKg
DgTPrIUbPgmQCm8pJ/B8iP3HmuJvNuoI3m3d2b3qpYIlTWHUyqxdG/G0j1iAtU87
N8QZPFaCLb6owdddtabvhClRfpqNJy1xXvbPL1xuED6YMiX5XEbp0L7WKJBczZmx
Q3y8geDTf5gvucrwORlHwBveP99363YS9smKlm+7Jn01P+WS0uSaC4IlLnVw6Sfi
vI8v+0eVhjd73hXQhj0h0StoC+DGZWBiV9OBh6bAaftRg67yYLKx3FGvXuyESnwX
tQbbuY+EAKIsB5G0IeMeZ7iAWL8Te+7m78tip3cgT7D2IwSyhWKzOkbFBOkHG8rK
ZbkiX2h/OzDOdKyc+gvzoJKKeaso9CcVM/Sq3FMs41ttq8NPVgE4Acv3sR6JdbSM
e9/XE3Nq7xCdEEYBhZZhFJG4Gm+yAAHrSJwiEZfe+/Uhq51oNcGpilqfCGD6bzQW
ZNeuy/2Ht6MD9k7XwaJiQgPg/uuNwhz1qvxevX9nGVR+SVoC27q6xC/xhZl+GAUJ
AnCVq9qs101PuwiybarhUrT869okgb/5yn/aT8KvOA557rpE+lNNdpO/CYfxUK4h
d7Gukg/BCPrif4Y2rim4GsOmqYllaQE5lDYAGm3EudxceRjb9k7bBXUQsQseyR1z
JSJ0oTDQa7+AWePgCvPUaDq6QuTee90MvBtePY5rJS6OjZNZYQg6J1+XsJy7J3Y1
8rSV8hHEJFaym5HAVoP5fUG+fsoRMIxq2ic7SCZHw/2kA6HjlKib7WUGotaP0FPH
Q5no5dnFMT7jFydESDzf1yp3OolvmkYtgTFKNakxlVrIOJr9zF6Ldt7myjUnm5Mm
75HYN86isMqGSV5kt0lsaFZ0Jotq319CS8lTf9cd2D6fziruAzg3LYIJws2nMYLZ
tsI+QPISgrNzBiouGe9LUEkhFYmc6dwkOoFZ5jsB+SuNoVQTmh0FNp9iz40VlAkc
VEPFCigAc1hKVHLP9NW8CD5/yVqAIqf5BvZO8ZtMTAl/cG6u3WPov/n06xIcHrE+
qC7F0pynTECfiQA7nbREsBNfsebHE3DTFJa6gqK1VoEO921Dvw5aUbuX6ecgX/Yw
1Tn2AZq/Nh63XGcTvB2cYurGhdT8+hoEv3uzEYMpS2HLoZdywJaVrrSwQqYmPyf2
tOkBSiYaM4E8AraMyWoNMVIpC/TfuFk1sDlBvoMog8PkXDwL13kjjpS5OrrlR2II
9yhOU8Xi9t9Bxn3c0N1tZs4PhMxcQs62OWrRyFQfCnrLGUP1y4H5jP/oFATBdWw6
MhWQ9M2guZypW1ewaqo9EX0cy4ONnFwyiC4Qv8JZEMGRb+jJXF++fvb8TMvDsHGS
j+ET6lyxroKXu6ch3QvAtHyqQzel3wLHoMUErEJyQJ8wyveppgv4Wge+xMjRQ/S7
rZwfuKlyhRLusCKbMp36uApRd1rW1vHs52JP816+gC8n14wduyFCtpZLVtWSVFEG
n4XXAig90pxfJynDlqH1XZsohNP1NLartsEosbMe6eNFX69Cf2fpN112asv8fE5m
S1CWc2HGVqYAXGNoqjAkqkbqU28/HIh9VAd0ta783cuHADtkUAx8EoESGqAfXKRm
TRpLeTrjPRadHe7e9ZqH0ahZDDcOvWoOhHkvOcZXIzXO0KMVMXWNM24FUMK7Uvre
w9dzqCxv/8ORA5V6ZB5CqBSH5F69Dt0EmKwHTd5AsMRjoIzxkC9qLd2qnMZSJDx2
2iV8uZLB3cZNKw3ntdiUOuAeVBxVdSJTM2PjW5waU1bSew52Ju2STyGM1Lx3IDet
/0mgJdFGVAT7mRZzHmjzITS85zGIjEOAtSwKG+Z64p6FqNBpukr4bWElzt5N025f
PtA/b4wtKsg16w33WEojQbXKFxzI5qkN7BPrS99M8fqolJE9ctpHmv/N5pdb7OGe
KiGa7U+KylzI9FHwwqqP3QxmhXAuqJ86zyLiEcG1pqTSBs1EPIR8m8KbLV3iO3Kn
XJzV0BL5oNSV63CnSPlLjF05hUGByfZcIvCtAmPw5UwYVmdSeYM6vOlOksaZz1ZJ
BmN9QArzx6Ss9hx3kxXfJlY8fIMhkgeu0kfY21MJk1nDeQKlRWd3a7Efbe4rRpXd
VSplJxhmSCj8ycRH/oZ+JWEOZrlG2JhMQ3AZdxZjw7JSJP2At7Cdn2BvxhJLSZz1
1TM7EMvtWW6q6e8txm1FAuUBztDhtrhvLfmazcrulHpqUkFzttxsW9mrIf0Uaykc
h5lYCkdAUVGmnlLV+clT85jDFVl19RqWryeCSMUH6gxJUScerJCQLYiMg0Jo8W/6
ZZnVOLMMityhrti/DCiFD/nc1diu8n9inrNT9cT2qG5UUriKwRUiV3wVwihiV3om
26QJENILByWTxxaNOvBXHvz8tqID1SlRqEROP/Wf+EdTxH1SWwMkM8+MQtCP3H80
ObSHbF+P2ACNnwMOohot4bttmP+yA07kr2DTJZAkB4meBsO06P2eG+UaPRD/czcD
/dMzxxkNRaL/DivS14OICiAT+Z6F9lgLRjsLo+Xcf0DMQzHqQfqRO2VTaxDdOgLd
ObuKXO9vCeve/0V3H10EVHJfAvRsug6bJxcbjRcMxujqGyQEs0/BPVXdKxcOHM3+
f4soaMhE9hSCPIFjeb1qDaJaOp+VTjC3aH0GOhFUoY/N68ATQcgskEDwsdm5lJ/7
JACKnISOguPRYWxeJUyvDXdJp/y7TOphB3xf9krDTWRaih23U6zzNZILTsibofoc
/Uw9vtu2EaSjO5XZd+J1//un/+XXOn3N6DMbKFjvwQ+igTv0Quh6gk2MfpxHPYES
xgAo59lTttNvGf0JjjLCaI+GjI7WPm2whxBdscV/x4LRAVc5e3px2FVs88DQwDcE
A8mqG5Pn9nDgZu1g5o7NdZkofSqZq40rrnqmozWloXHax2pVKZf4LqCPffO2+xJO
PXlLiNWQxq02F5KYoCHCkl/oZyjEvGxG3kSauRlq/2Gchqu9vJeFzbJabJ+HaM5o
mInHtnLWjs2PqyEck9Q1OL2ibwG3URVRdawyD+nqPDKlC+Mce+xBWeDqJioHJ8es
DK0spLDcsXZIRPX6tqJB+QSnjBbF9w+xdQ64TpBbQYphDYTcVzWu/MIxrX0yQMN3
ky4Lxz0xO6xoxKCGxYFMcC1fZfusHvLeHxM5cFZQP+5s48HeAe9BxVGb3yr78PNl
yR4M7oZeh/7iT9lNL6hjbdkzLIOvanwXn9YONmqF0EDREsLP9gFChEVMN2GT5zK4
Vn6D0f3zW8JaKHrJ7nZVYVs3tkJT9jb196Hu+Gbh3GmRRN2PHdIyCmO9EkpgftFg
B5uf2NATcYK3UT1TmPWEA46gEl2LakEnOYmMeoH/XrCuOR1HJmf5jPHTE5hC27wj
1t4vYSs5MSFb+aOaeGUHf1qzxMs9JQQSieq7ySKd6ceHPnViOTuy/+m7O4KCokEj
2SLJsrtiLVbgEywn/qSIB+ZG2dMmAhKb3XRWeUFEk72mM1Lx0UMuxZUc4BDLo3h/
9NBjw7xz84IuRdro0XHRQpRfzywHCZUpG0c6GzTwBXTdRakc0V42ed9E77rjm/J2
P1eNpfg5ccmw66EfHcr/B81G5tQZQ6c2IvH7CSbWVnC0QXKNKMOX51MHvtLnQwa8
SaFmfgqTXwETKe+il365YUUYp6a55ZgOTAjKIkYfQBf+zQ9f12IeqMQvevOHGBu4
FJTb76U8gqHQIFXDGeeVKZABGwlaB8SrImxf6YMjYk2fcvIQ82ZSr87bxB4u71kH
b2FfPnZ583V+KBvRHMIFfbnLy1exIrZiTNFO2sLQFzLYEkaY+QT9GXbhUobc7oxL
6GjYoM7qkIR0X/+F7vfLK09dEUGlF0NN1n2fMSwRz0d1EQCIQxdxr00FLIxj0La5
G/wiq0dhgTcOQW8cjRtUe4h4bTR/idYon0qynzowFh/E67wy1ht8w+GU7Rlqtd2T
lZhAdC6vJIAH1AEMMYH8cSsJi+lTmfzy0/YjZsXnabjj0Oh6Mwp7EPegqkZypZ6p
xKpcKs89F0rODJPvxYyQwiTUW74Vnhod7+XRA2UFiF9s7dmfTfPOwpVkRRvOZgES
lbmyKTsMCST4kc+AcB+0aU7moQtsnD4IOrr+AS0+ayz98I8MpUfaV8twSbMQGr8G
t94/EE7MCG/5rnilmW2NGIx74R9lYS6UuBHEM2v4ncGOQU7urK7fyxspSApY61g8
UJr7eIVHIe32nFvqXZ3/EkIytEKuTyvrsasKkUEYG69M8/9vsEC8iJJ5VCFzF4ZX
euBKEHNe66rhAzGQNM/z1QFRi4C6euh2L2FVZMWAeQ2IhAc1uBQrWbGJao2da62n
p6J3sU+K1v2OQFhiZmnRpQ3TW88dvRPcRusuB6DS6dCqXmU0jHc08TSO1fMODahk
8iknmya255u/obe3AErLDR6FscH8ObZbmDomfTTA6NIsiK04eap1MvzcusKAhej5
4OVf7aY0urmnhHbXynXHyrGpxTfUnqWaWxgL276ZrDA5wrfaTvKtOB9H0r6JL8Gz
niCKmBtuSDNCFWuK/TnLV2Z2feXis/SJ0w2d8c0U8phV8Z5mhz7jRGzZpbYEWDfZ
S6932e0GegpPWMk88e/cE/XaW1gMYbngqvTU4peUbSiZ65Q7IIGldeyS+2oYJvEQ
mjYzxmYoAqGT8eLCcjzLm70IXPrPTaEnRWMJzVbdCrbMwt0e0/Ua+7QENp343aMm
cQIgHgs0HNgDV19nq6QICnB/PQWKPYnzWOEiy7aA2i3yCDk+LlNUpJ2LRPmg9MvZ
jcGJ6ZvigPqxkywWN/aKBVl6uEj0MZxy4A+7wUWBbFOH8JtJBfpso/J6qnE2L7eD
UX85DuYW9uLSJF3Q1q6bFHgqY4Tlvu9w3YkHvn/BIvD+WQ1Tzi9cHkUgVeEMaNv/
vfqT1PSshXiK36pGi63y/A6nQZKkf8369F104PdWJjhI/KmoFOiBaMngZoiFIeNv
e5PZ5HZZaXY2n2kPVw1qoehMu6X4J7K4Tb8/Yy+Delmt9UrTyLKxfz4VePXsKAuJ
0fXkOAvyrMOkW8KOClbgfArgH5ZYfzVckPWnPnxUPHoS9h9Cb54metlcAk9EPP6Z
4Te7Xe09ylK1PlcMmHL/zi+lnRTNiC1nnv9YwjZi03UHjGkd25cy/Y7FmODYcWLV
YPXiz3OHnJuxjCngdjVMsq4UmFVcq7Aa48sYc3ccNTn+3hdHoFrstcRZ7MxzT95D
1JRmxPJfsIFQrchYePItpIpfVnIkHKklBzb5UQRVVPItmVkWVLX/JJsskNCJsj2I
2KoeL0R/Sl6Xl4T8IaahvxgnXm6USvWAyndJCbP8n1wxn6C99QhGw1UcFtze6Agr
h3+iXn548+MhaDi4l0C9xtTys1NKiOddBU1lbp/cECE7CwlpiCWH6tAJgMmpjXeP
HW+2vy2gqPD0JFb7PkKOau6T1q9JAG4UkUsobwrgBTeqia4QWIfvPPW7c/A66IZJ
7dFsvqjHWU8NrmWdWyaNYUjAILCHD/5LNx+HEVTIoia+eQUYfCE59W8+MHFivd7s
oVwGuS7fMqNL5YL+4ziJtdc/7l5y6zD5cjvNbtFrZxx/pmrwaZXjjFw01gK9U+Ic
d1Ps0wK2/+wxXP2u5L0S35WL3bPMU22E23djzebn5PYftjvI74HqpLKUo+8YHyoo
9Vl0+6c9zVvdbcu/boLabBBmqGxdQNieU0IJ9YZ9HMFjO3awvUy4aS7GK2myfiCf
vOBHDKBdK/6GlcTQ7cZAvgMqarS7JobUsKaQ7F009ILG4wkllvGuqfOfmdXekiaQ
k9K74ybOEETXoRYI/xYNYXeEOzNkg3kMyCMg9A+S8556/hBGpQthw5pJZjP3fIRO
SC5NweSAYa8QQVotLGyAPCNVFUCh3eFJDeiTu2jEbZ0B7os4/UX662TNUrEDoCE7
JejX99x+kxf4oWn2GHZ+8yUsaCf8emsWckxO2SGAO+iUXzDt8z4nDlIap00au+n1
+NukW1vb2AZ8m8v14SJpCV4LTo5v7awjvpejVSWFeDWW7a5ttQWq7REhQgxOGmmQ
8JrrJVM+aAUvGkeW+NUG0jOgG6m8ju29gchZC2ZHoXXPZ8GAKp1DHnaEJ06S3OrP
gQRiAmqYo4kS0+Z1R7be52WN+1uQXtIqrz8/we12O8fY9pgWcROrZgVO8QajBhCU
xqUOov/I9wnSB4ySY9nlmpuiyAGzqO9MwTXdunFyk0vfIhbLXHzB7Yfatm5YKvWO
mj3D397xkICtoINstuwf6ui4x+5vkAriactcA17+F9+cc9UZNj70G1UToooSrN20
U0Pe8YaFrT1pt/oGntFqqi9utM+0Ze6uf03rqnbu2osbRkxzgLGpQm8Ca3sDZ9Jj
rTwIUehZ8uYs8nE/4/p09Py6DaLg6OX+jd2e//U7vH1FTzTo7prBeokQzX2SDI7b
FX1Gs7hZiTrmEbgqbGKY6OnFa6mVVxxdMDgLrPqAloFaoqYH5IS6hOGsL8CY+9dd
jSRs3+9fG6pk8b7HtnohanwMKoxsX4b3siLueklW13EsRMlpLj68TJRyZC3QLgqO
mZekN9bso1D1WjtRKnWFLq9gQsxPOAUxfPcFS1bB4obrECj9PdJMdGHerfXwJZMV
/ca/24Nl89brHOQ9Mh7nsCpAggBsQYOSuMvt7mTmstbce/VEyWgU0GIUXJcwSXMY
pyya9UE1i/L+aXt73rx0XIIGLKrhxescgbxXdKhWqB06fH33iM24KL6D+UjpZ54l
iU8wMKkHxx60CcxwGULilLAJFLs/jyQ4Fl4i9DadGHsKw9FTUrZMJe9SxgWYeXLw
dQXl0T/ZocSHxPnHct/EOx8umkHtu/brpXYzUfbqdHWZXPS7kF5b/ZxFF10EiKML
BWGOuJH+qjXkLxmK0tI3zgzvisaTRXZbyljJmZXO/1/sWD3Nb3r+v+Hqgn8hH9EE
04zjT5N2J63i7OB/2H/uAW9QgBehcLYusMlj8KUfsOiF2srqwCXZJ6w/QEVLeYKr
h2ZJeUSjXPcY1uzYobrpB/93mzWh90g3LQU/3SCO519Esng+AIlUqWI4eU/z47pO
R54JdJVFlumbhDed2WLkLFZ0vORIA+zwB2Tu7mjatQFAt/lRDh8wYpxlhaKd3DtM
eckKYtBCytR961kR3m/mU9Gf0Ir29H1HSrb3jW8LgFvAjNa0LB6rLvg4al5Ekx1r
BjCpcMCIzMJI78wIap1vUm214cvics/98P8NRkF2NjHyfaAOZ/bhfKF47X7xEuG7
WGeLPcuDgkgRFrtCcyLg0bMBN8CVdGPMiwNSiwOhsJex2YkGL5NA+mDqeeKCW4Nk
HhAg6CbVe/zlDHCNOa2To0cgsS+doloN+aCIRVj9UMdkTY5Fm8g6xsFahFh1G8bF
VgqclYhuJPiz5ZXIj9SItP7hjAFl6acFD253zERwCa3DvCG9GLx27hLBJUlIM9hf
GiR7EXaPL27pNXCL56O/+ezsgL5eWMNqHf6owWeS1bbYlSYuR1NIHltjmsgsKgQr
5RIV7iP0kGeB1L+gwp+SG4wSNuVv43voGEwlbagSGtWT8Xfgq4TlBfHWcOZ9qQCc
j/zCiBVzX5wkVISfVdhZl5F4t6fPFCyTcerfqk2bAe+Kf7P7kwB0pbp+KkBGrabP
AaGmc3Zbh4LTFgG8CzYZTUuP3i1pZhJ+TeA4g4ZCEnoaean+KWF/z4sWHvxBuUF9
2COAzRDWyY8IQEA7PyrChnrV0XxboXMMwwUaaGffFE8YpQzzrxMYqP8lJ3P15SHd
F+p6lIOVgu4Hpcpl49tsGzYVUqnqxuc4ChOeCQ4OGhhKXJqldvBv3485W+DGw0v5
EZ0eTGe+56h4nzQPkKnq39ExQdp5vEj2JrM/PHrUvEBxQ6Ju6pIwRQbO7DhTXAM8
P04tc7K66VuBkRRS39V6r17/KtJBAmHXxLGaQHbu5wbf3TsjRG6+k3Gx13DGIEVg
T8LZP/r3EyN4vmrEinVPPRv9tbvF6J5mqxikOKzOTV+eSspv8nIQcVAxwrmnIHfm
+NJiWIoGtak82k1grH4AC/aEHbaNqX6QShI5bAfNSkqTFgC00Dd5SJrdx8bXGmPE
P1Bw5Er6zJbUkRlWCm3uwTpjm8rvJ21Q0aGoU2nyL7Wh71oWOt6GrN1gTVqrePQy
aMRhMMA3/ABcMZksGqIS3bEFuJmYn2fN4NT9P2MbqK80oayiafL2I1Zd/Rkfo3fq
BH4Ob4sCq/COJT8QTsz4Jmu/606QPSob+SeO2uF7CEjsFU5/xl5KA06vABR2pRGr
wNsRkg1DnKzrw/iKjP1D80O2NZUG797vHI/ZLFxutxN4UPlhSo+8WYeoKr5mxHbm
HkF1mPO8S84iEQ7Wn3dlGLlxo4Y8L9biG6SUB1FN5LK3Yo8yvu3P4rJg9PNl/3ku
o/WeXykQhYY64Rm1GiNBwW8nRELFZHbqYB2pcM11THkdz5j7SpMZzLk4UBjHx+G+
/yhTnYcVK+w6Zpx+sXdSYg4Tfjq/mHX/HAe/7xltpHoVl9gv4xtDSL2B1n1yUr/u
zmHjg7seTI87QmEzmnP+2D8FuV44FGbp5sPMwifb/nTX6k7gBqch6lVSdTAvR9Qd
Y3fOi/SIf8bU37eNvyrdZN278qcdBX2J1cw3KuTo0kZ/YjiFFfXkblnrA7QbNEW1
yhjIWJFUuZ5PnaAGmBZhMJZyG/C6tU0pwH45xDg/k5Drr/6r3Pm4UZHhQZR4kr5R
fgwrFwMx8VF1kAoXPh5AD386aqEUPwm5fyvV5V9KIk/e/hcqyvH4UJ1nwfKN+m+1
z72wgODJxCxeF8FdklvNqXie4cXKT0TudvBehH7iK/vzfJodb85NXU+uvqZnUnpc
oluA4CXDbR1pz5reE2OFbaFBXA/sOxYLSUlmSTZfr+BiABjBil3feQY5XTUhyt48
pWvCKB1Ut/l7iI2wh4/QZISdNSrcAc33m80HYWLIPAh3eXqpoSNstm8+HO9vzyH3
NC/R0Zaaa/eoS9we+CGrHlHB53cDKiKa/TOGwUXrMBuMH8w/xWucPVD0MWLLgVjj
JvyqQcF9pvtQbrBTlbKw+tKRSFFwANwKrYBGZI6k0Z+YM6WswPbnaxJ0CKSwgLM8
ED+jpDHs2MR/dmhoiXksB9UsX0iWOqohgXbbTWaPKX1PnUbhzXAe3oFp1VbQN3+y
6365VgKHzlxyUFvXY2uPX/J3zK3j0BL0XtAXZl0FBM24kpr36oZOD1AiDESmPKcl
SnyrW2lGe09Dd48y0eTSy18W21qg9muFhB0VwuxLl9Qk6DeHUAsiPyDIXXQOpU3C
QNSXsNyHANPv8MztMYzNkWJ02AzQYL66o01CWw8Taow9YkWoLxCFonVDmnFewRYc
5cVRAafte44g1ERDfaMNDFhdlkmCQvA4AEifnMKbmmv66a79F274h8s9Iahcm75k
5jPZSJmtLDDciPzsLO6CsNo5Se3C9a659V3ir5+1Mi4vGyNdzqsfPa8DZ8G/iGVe
QlRIp6/MFrLgChPGe1vv0lnhKRi6MebQaezLXk6Zh9oR+f4ALoxWaP8NBz1rtB8p
SIzjvpGis1XM3H7rCRbgif93hOXSr2fV3s0mDjljzZEu3HD8GmLJkPOyG1Eq1k8w
XZ2jF5I2//BAiLj4R82u2cOE3tcEvakNd7i/2CEVX7YRPUln4l8vSMtFqJ/kf5SC
trTNslp5Cnuub4pn1wBge70Rr10lpHsBxjXZYYr2MncSB4ueiqb8aXmYhsj2qHWG
STjfJBUVwYdxWe5cOvMbf3vbrOe/jrc5ZVCz3CbFn6W58IX7FNttJS6m6CWumwDA
59HXC/fHUEjfaPxxI19yVs8fxRjRXeF8FRk4rv5mpuEEzXg2ioHzN4hNPC5swk9Y
KC4Ul5f4usWq11Zh2WzYVgU+k019Ox3nkCMhpuSKWf6nhB3rabpeszJbar9aCmJo
yQ1Wcge5tmapPf7x6rJbF05j6w9cYfbgnqgQwGVmIOiXNFKaMEJL/MmucpAXUCI0
Xlu6LqkUe98w5mhLotT+AuWg9HGQKt0TE3aPhZdYTq99+YBiJLjJIhay3DuUDi3o
EyftCkbfjFf9Zo4vYRSXBryb1TgUD4OQtlFK0DKz2y3GcE2Apoz3hZnQv/VEF97r
BjEILHE6fLSoYekMPIQlelYaZPRyh+kotvV2F/zjugNGwgW1YmSveO+jLjSSaA6C
zlAku6PzATpGKsnB5IFron3CVog1Nu3gwXIGI1jN7UxMN4IFFv6jec/pBFmBk3gJ
2553gUQ+MLktvYB8qxMnVvipEaJvkcjlH0WQIZF3/2EmMl18mi0yVfTxxD/2KR1s
JkVQaTbYiKowI244PeKBH4lJDI31g/DdrskGrrQbgD+xaDCRB5WgA+DpEI6s98zl
B6QmwzLY5hx82phN2FAy9J0kUDrKeIXkh+rlW0X573QvWhu+7/zYGGtGeBcIdgv9
tk5zQGoEfFEtQBfZ2z7VA+/5DFRAywwrDcvqJE9jQmacFF4n/lC37+L3pTxeZEm1
Rvtf3LJIA7Dzf4tPPubest9KDXBmdVSzxLuj3cQLcjDDvANdG9qiWMCUE9ZFChFF
kO7/Mu0e9ugDhVW0SV5dF0lDtWTiREG0hdAxR26RX45Dy24HLGCRUW0831sA0I/S
M6MQlyTDv5fsl57/5NuWwGvlsBodGX4vHjnRz1YVzA8U4UqUpqAFiQNZuo0FpqVr
u++atLej0copmc3Ri6/SF5UEDV2OVVE3HQLwFUNl5qHJclaUfluLRrRHUJ6lbKtF
n8YsolRsqUw+uw3IT0+aIPbdRDVMFYT/cKc+COOb7FwktRFyFxqlAyMskgU0uXXI
FG3YfoEMlyPRP3gVY7NNBw8lwgQq90a7MyCKRI0hrLnCGxrhCJpcI/7dAGOPoyIL
1h+iDlTBJEqkJZ5V4/jC4fi5CfSM2SL3ttzalBMCiZsTS1/7XiF2autgV/Rb6PKh
vGn6n1mff1PuaZH+r5M6Xp+TkzzlKPvQOMckF8OUf+ASNdCKrIZ/zGhblTcspqD2
xApUICR53a8DfJtCUlr3i4GhyhcBR5GOBITYA222kTB4u91MdDBGfPCc5laCJ0i5
NqM+dTHgP/h1jnVhCLtwxBW8FW14E1dHSow6+in6MnooRPAE/b5aElnHG4/T33KS
I+XpcIwBBfH2jvvRx0gg2Ii+bfhw6bPFQ4yJSqXlIqR5lSiJ2ePwRG2pheJr+2qp
5UjKA7jxxIJzqndXgRgMs+axLiq9lRgrmfg2Wh3MdJPEGFifWmTA9wd4Zjjf7TOw
DWAX2G3+rpAdNXP1qHmgsc14L1VUYCyFQbz4J4Q6fCTXmRlB3wmmNxWzXXjSAdt/
wTw8QpYnxy0jIzckpWZ7BC3xcPqfz9+ZZtv+VU/Gs9LqXCpsaxaJoM3FPl/xp9tr
SdOTWfQdFImbaCQNs++FQTl4SPUWeKNOnqkQlxUOIr/BBE+mAa39ntgQPvLpFIFU
Py/u4z4t8DNWhhIepPvW34284jZwT0gsZg0NDdkSGKoYj7HLm3iJ5LIMJBP39lml
rXV9Ou1S2uWf3bHTe0qYroCcpxg3/nJ8XCFpDe5nhlzsJsoLHTM3f8pcK6DzmUJz
J5nqhq03xh1DZSxnJ1ztPo4FAkKT+IY63IdD0tT7TGVK6cUe2b+s1EMuuNOVA3bq
jimFvWu+87f89gz6UApMjCvuIqIpIlXkXov/NEx7a0CGOsbyHpb78O8q+iFU8sTL
Uf8Vpfve2e2BsjhPTaM1JnpXHyk1NijxjY2u2OI1GaJi1x4/dTDSdmktcSiRJb6J
RJZRB0XRTRqcA0EE8vqsZwRmBM5JUgTRVkDNFNTxqAxbnY/C+ON8M0nH558MG8Qw
kuxQc9wBdzYsClTYfBqpn1E7y8lJ9DVRva5GzlNzup0KVB+WvmddkC7RYovBIGbi
pLLIfR2X4aBGtIJy8iHgebTEbnX5eVyjj4db0yw6GtcC7LS50rtK18K2vYJ6oG6v
ompNIhc2+80e7g/9J4evB9p2u8k124KD69/fweNzL4iE9T3RvTHpoCxTsDhnTMh3
3vNMNWc7QbYrJ93yvHquLzwFMSCbtBJdGKPNvDwfDCVxxBoE3VilJ1PsTvcVq+pe
uuaDSIBdeEgSGmR2iZNeDpMZY1LgYVavG85V/7TfwI2mhHHgInCq55X4EwW0SAH7
4RKUO8F8U9U2TNckyeuFkqO2897iobjEBRnuc8bdgwIRLXQO2baxZu1KmAyEjAM6
LAEOQ+nhNIpHSxMGllckkkmpCDm874sdlk4aXKUKaw/TCesuYOE+aS/6ElZfGZsC
pkICBDLxnLZV92d0Q/WZyc7bouYP7l/zUjC5i+HHLHtYkcTbDd0N0WSuNTZEiyI2
uTLPPHzDMBTFzrBTUReRzvyjBNP/xis2xzAhDOnygIoDzX4iaXU1cMlykpkZWoYU
I+PaCNvWhw0Gnt02Xr68mLmEN1YHwPaNRcPO3DZRcTyHdcZ3yt1WWva62FJgLcxD
ocbNgHHZ2CU364k+ua7+HBPXo6hzuamT8V1fgt8QLxZGp1vRSqJnfu69SdwO5HPr
H4i2+WzgNuUItc8/d2CcZEnbAkZi/hrw82Qi0NIcCGGJAkpTr0P77Id41/3QsodM
3EJPzsIaILkVN82W+a78Bjamz/6cF/Azp/p/tvlhK5hiuoxnVp6M/6F8crskQgIN
YWURX6yTuJgHX0wb+dlkYeoyxojd40mB5MvNQs7pqaAJZTeI/qOBWI3fYvhnRBo9
gMNvUoamBSAmIsNkJTDf5DwQM9oLwe6okGNDPc9Mx+/HQH2LQ/GYrXWQQmJndq9R
qXfCaR4OcQzcUoMIp7jy621NwoeFTYBZ6/vKy2xyeTClVVoMFXjYhvZ8sO8w2Ezq
wUQVYr3FmEerbPLGiZNVLe4QywHk9nADH33R5S7RFDhI6cP25hVkkskYuht6MKS/
cSgqdllYlpmkYgqVt8FTpCustl0pVNInGAQx/C/4kGYpDXJTdHUXx9ZDppqnk3gr
K0esoVK+YiyEOR4tA/3g3h3vUT96puOa3E3/QLcRRfHWYLQvsAxUfV9vhOpysVRy
42B5VyDx6VdxdchuNg1d/sMfjb/bx8TahkQVB2KUk9jfk9NRl/0GVOiepmq9/SOb
5tYovwIbYZl11DwO1p2TJSifuVdx0HMJWsEZeWXKJTpaAiFtjbsFERMceL3FEj0y
C33rR/mfXfd7C3oNQ8daGhWByR07//uqBq1A9ncIKRMytMPg26xICYnTF84ujaXd
sUJvuvxyKgXdBSAI8Ug+fBy32IJ8KSHDKA58z0j4HsgjtUuHj5NICsS56ery4QSx
iM2rjmPKe4Hyu/Smrl/nrmns3Z2uTaqjuIx8LThK1FOSxRhHka8JeVHb5gheC+Od
JeoOY9bQb70CftoFGcyJjAsL2KzjNT4CAuI/Bj6lCyTJ2IMXjVwk0EB8qLnYgLAf
Q0SvTXAxdpWeIiRZ/sYlkODJL6g6atdVko566yIANJsoCWN/GAd+6WeMo28ffOEk
6/9qRvx3O4HtnbUQUIY5ZZKTt+kUtgYvCL2iSX3pRqNrzMFS6/GSsMb4aFyefp0U
yuEW1rjQaL6FEB5SfuTJNlkFIkktnLAENX7D5o45S/8F7qouX9we4COkKk4NuqqV
f7DZSDhG3mfdToVizvf7gtCTVsIyQCOsldo4IqXYUN1TMNn0ozk1yZHD9pp44JYz
qoZRSDQJdFRMUwze8gjPAVXp4WLflTCJlxk1kKX7CG6vakAdvuZa39tRQyV4t941
UEzM21aXh7rl4clmdAqEafg5EQyMY+qbV9M4Awnjhty3Xl1xtL012pWXNimlccpQ
dTAmJkDRALGES/Kz1FAAbuKDYoBD46yRB4gxbbemsC1dS3/NDOqxgizK1RO//XmL
h2Y7ZwusawLa23UVZIhAd6WGhrLneA0PKGLkqStaRCtl5GpS7cwqtb2TbroS8BSs
XtLaBKS+tjauiC9zh2eTTJ4R5LBYeW5+8S0FjU0sYegbB8YznZ0SbPIBAXl2Bktg
MxKVNVhg3HXpYlIHABaAlg12zvfZJDOFTMcoKlWM6JEtpMyAi/rXPqMhmAVBSZOx
trd4DtDG4Tu60O19tbX/4ez7rTVBaC1cc1f2K4RgLV3cpGsyb3cS//S1lOKzdBQT
IOoWIulJDd4dO3HaNoL9re9KGjyaA06x1ruYbuGENCO34mRSMus3v0S1tM1FgRz4
IGe8B3ON5yXUlIYFPBM0quz87KBG4VPUowYCds5TtJsEeyco+c5TuH6TEkGXTNDE
pA6PmI0ZDH324mTrR+p5zFI6OhhH3rpJnLe5pm8nPH4qeEBrzH14atv4tmKq+PLo
B7IoSUUPsIKAgKqodsUcmXDzBZbpavs1rwCZ63cLERQuYUH85IzTl3WZhxbmsrgj
Fqeyut8d1T8Q0CW96/0kIYXf8by+ZxMDtzqn8SmjuT0EBcJJI7oNkZmSHmxF6ggV
MTWk3+UNQrUPUxAjFvHqCWDAbTWSVOuwVXFlqb76NrPLawXJ7GE6nlsJ8rVIZA8n
toq93wozpZU3zydAbmvEVWZG5Qb3NthJQwtuxh5UB92j7S+/N6rFDvXo3gSGmro5
a3E0hRJNh+vQz+7y29XJJ7NJ8ZBinMTxx5PaFET9DQRJWGpfR3dJR6fddH0fZ8RH
27vvxGKEOo6YYZ+IiKZOnAWw3OJTteu0om/J2zWf+DLdlV+MODtHJTJ0YcxXsyIR
zUHYLAHHo8leVcQSYYtzYhkN7NajllVRJ7Pi5Y6a7wAkg+DOcCv/W7rrX5N48AtN
0y/ahJ1WOA6qTxlduWvpxgchUz1XAi1x4lRftRUm5I3SaJufsNW5PFvndGnP9303
WY7S9ctzC0lwbKqBULsK/utrNwpVo6/srBh1ZEn7qckz2tRDeddbH0qXXOUKPiq6
PZAPmFjhickUuNU1gT9HoaRNofMy1GHxiqkkE3UbVGI78ShPV95MzR7acOl0kw+T
Sevv5S+qKzO1Fi24Lw+l9vBrs8N4oGTn3LxDiWz/u8JUGIwZIxxUWM9jKCviuMPA
rg3cekf2VNSr0nradUCejlCMV29wfRHyccBYUE06UqAGOpdNe5LKG7pPnVqdJbBM
CQJEi9XdpSm6QWlAtWTwUBm8J+DgwVNkZxB1Rww+7w8uZ/eClsXyF7a+HtVE7Vi9
+dnZBjFPpqEP4xhu94Jln5/AE/jXZMzxqj1ImNob/h7Ok/ye2FgDFD5tU3GjWon5
r9/kXcUa6TEqMWA0dUIz7M1mh4+stGqZqtWea9Ba5Pt2/MhkbMkj5kgEJ4bFCIzn
6uArNu9oVOjg6ZKrHtpOJ+XAoot6/49rs0dTEDVs6ctnM59du9G96RTnlvCf13dp
t0qJkQi/ycA2p3aOZ68CsuxCdsotM8rZ3OmzwNZrCvwz+5R33Mok2E/OGs5eOQz/
Nygbc6MQYrVoR3Nipno9nElsmM6yALBNKxc4viFXQHRUU4dcmoWdb0V5uVP4vyRp
njA/C4RPSfzZWv2/p9ulktrklCpWyjxGXuj2N4bgDEYA+14MS1ARyOfrLllXr81r
Y2L6g/HaCgEMWHNPet+lFzkjpfohUcoY2THvoMJrp33Z9d2Qkp9DhaUjVUmIZnS5
IE3Rl2IrAe0FfeWQIenMeIDr9aQ4LkBSqFIMq3fnT5yryf16OgzBjyoq9k5WZ4Rt
9MwNgpwUOKiS2sAVQ0pSIslhj51MlVTzoDnOatM/64aDanZSLPUDpE7zGKTT2hOi
4JBdnIebFwtibxY7MJ/eZN9WE4M3S/vJwHxbXcJK8h7IqV7oj8E3TcjFrz8nv6Ty
eMz5X6aYR3cC13gb4Qz20YBTylrOt011VuASSHAgjG+elLzJGM3Nj78w0tCGrggr
vMP9nl/A5LBEesqN3CYybvI8ec6YLgSVMHS2qdhMWVfZegQHW5/WVCzMEfWaT4Yt
AAODIa0rlF+BA/3xO/jJE+P+19XANzJoGCCeV44TCf+qROFpBlITlVEtWf8f7tj4
SKc05sB6IawT4N4u90R8Mj6bLtALqnZtCGpksObWeUF1nDfDpaCz6G8JvAY+tTuL
7wXY6jeMmKAP/Qo347oMW2uXiuO9rfwp/hIWx4LsrZUQB1vkvwWugKJxrXgeBRyW
MzuR0XBmrJ8spjDJoaSKTG9TAu/N+7gqCAI7Ea06GSBvipxmg0nGBWDprpVRf6CF
WKHtKu04NNTVcAtHTTDmSTqZtMa0/gk8lWCsjxitr5gc0sfCLo0qIITL31BBootr
5R+k4MzyecO4gMkNF+ABo9XOaNV7d7tL2tO4nhizBUyPApGPE1D+LAhrUQG7EgGi
3yLTLptFwRJMFTuzWluEvmg99qOpOKYNkp8vFXL7jiyKqCJghxUhw6Dc+7N8x7en
NRQMfsXcXBjhfAbjyEpfZAzTnoPMLVp++Lm8WzIL4zN88KmQqnODqyIsOagO3V8M
lpd0PokhaZWLnc53sin788ZI0BHd5wThilH/NpZO2Gd27Xa6aaCDGg1Qbk/Yhq6B
Q6uAWenftt20VWNBHLmQpYRkFQ4kI/s/K7XNyo2dlw/GGwotQ6bp8Lsu+v3O/+aS
sP9TQyW9D0/2TGJDkUm5zsxxrG7eorVJObQ7tqLc+VnrK524TFZVOeADQdp0X73G
UBBVDE5KFl3X3SXmOUDfcLddtf2n9U92psHZbJEIbrLcbt1uqRL+4XDMdodVMYXA
DVuT7Mx7K3eeT1DOUoHTwjkAlGAq1SEqnifRPKpm/EV0vuyz8Ly/P+oc1XfKM9/g
1u8FikxWFNW7ZZoPFYpbnXuPDvudFE4Oxv8bwsgoDNilqYqTRyiwdzEOrUzOglOg
0PXouPDLMkyCe2+EWhn81eLz553PL7gc1JM84G7WHyM9vKEvVrDaT633yp3e9S4Y
8NkFOeKI0GoTv4jn+pguwG7orWPCvBUzNvPPxXEID8+XiR4qiM0XC/I6+FKYCObJ
qyWDDidcQEjazZVtSCbDlMlqMk19NTFvUd+yqMF0AiYK4f4OFvitl0s5K46zRFrc
D0yCdIvonQYMkcVJn035VwpPulvN2L4A/dtzhprMgph3+oa95xS8kweifGk7w7QD
ij7/4Hma7o4MZpVk53UXPH5+kQMRAMiCRS7aMPSMoclqtJuR4gZthrKi/MEPBe94
TN8gRHNwsZ9POUAAsJedViDvk2/vqv/P3zj2MeuGKNlD7iDs67QLGH4KMVRnItHM
D0/QlYGZYz6S/OyyMt45l45DS8tn2yMN45y+Qfbe6lI0r9Vle7+3M0wqdBEhjIgq
+IxG3TKDbsA2mKXyqoXsUNYTyYH8kCH6eTpl7BzkIvDElFwGuY4LV3/n876jjsZp
usgbaZSv3t0RfCyIPMvuvKTgl3rLp/UDvFBuB2gPTOnfwPPmm31fSJbXUgOEppCU
KByYO1mpK047UHdizKN33hApRga/OYQL3bnXfy6DnymHDQREYQaP5NbODMgrWrSt
rrdFmLCDn5aJ9nFtVUOdbTc5ympVej9hRD87yW8Ax9W6WbxEr4UoMhGZFFntS4hk
nok6GF21Dp0qIlVuh25WmFxO0zzMtH+p0IaBeeHztRLexFF+WC8lKMZd8dTcOssb
PJLq6QwXBs+p96v2qhXRAMk9WVXNzt8zog34/SZh0C4vxHu9biLvTlreuWZsdQ0e
3da9x43asuwQOZtxcGcxFJ8Ig91CCsWZtQS5lZZoCXv2xTw8TYOfJ+RUfdD5w0UW
iPKVNaN6rXoWfTroVSc0zC/HnYPXTpCZTOrmKPXkLQpTAnAgnv69HuUBs4CPe/7R
qpB5ywmVOzvKLUPtHGKQSy30Fu6L0nwgJMROMa0ibJLZ+GMgsG6xNlicPOzK5w46
pNJCNJDxLFJ7H9m9Ru/1CP3yyNgd/jdPcxQcjFSjKhC4xsowhkvy3XPy/mUvoIaQ
2PaY5rCn0DF/6bzPpYDJOncuQRrfS+jfXAZgGJjXUt+TqrvI1xlQ+3Yy53sseIvt
5w0J3QkoMCy2ToYwoLd6D6rz0OrgrCuzC+seIeY/Dnp3qX7tMm/tkHZ2ZS49k4hl
LDWCt/dgW9J7FBqNCDDyEumgVN6PHv6tb5czle+RPMr78XbBWmGqN3K2OonIgB/Q
/KcGnTTrgrlPJUecj+TwV3dwzaKoFil4eTKIZtxGRa/6ND3oomeiGax3/Y9beRY+
snaO/WhXP5pSUg0l4yC8oySNp4O8VRh1/3WYlAqk0S0QXwUEMcxFG6gTWnDoqFUg
rNofE2WKndazapa8uEVnGKdUROQzQeNcFsQRU1sNWTdhnJG96Rp2I6L50Kz561ZI
MKXJPCsYwqhciaENGeuC6iU7aK+zxrvE3Y7xS8HnUZeWt41jLXvoJZ2Krkh1a28x
pbwj+rC2JCGswG6AkkFUbU5TlIGLhOW0tsDLNZtnYHmWRox5ZKo9GBEdDRbWrVJq
1gVPlc/yWGMT4qjPpcZx71dTsJgGLGdzIkT2Yc8SOobPvRPQMhWBnfdoDRBberlZ
qwftHBBZ6PYzB7vlCDKrqxLhpqV80YquYXeT39VhDGkk2W0VXwZPJr/b1dqG2+tA
mjTUi5eB718BKetqWflz/h31zDwZ6v1H7bD1g5Hdn/7k6NyC7D5CpirFYDtd5zrG
wVL+7s1fTvVLQfRsM4sh3+nNXBQ0EVCu9cE4XkrrMh2AZ7zp71MkzdtO+nnvydIZ
Xx1wGoCgrcfuRLu9Dhq4atUKtZyyfVYhULi9CD/oywRxn1mSV/rsA1ygxKH/Xp6u
+wxcArgTTbUdhv9AH8nFYqmr6bbhFCYpj0BXkIXNqMdSMhjvQbb5J+9/dTHPhxsn
+5RKo2uaY7kT4BXP+ScFPwXLNuQodrFDFh9pOGjFwQKDTXySG60RX556B0trlR5W
dIEO3whl4UlCvJxD/yh8MAydN8q2cut+oNR2wNd5eU/woknN4T1cQLJiqH9MWBIs
TXO0JYGacyK8AwScYSpvn0cxz9TOcgq7rzS230uaLtT6Pnuv7hHq7UWaLtiwapWe
Q45l5QP93cCp1Cn+YB0q/2dmB5pgWiBkmgrqE383G9X6nL/4xq8PEACEw2QraRUa
dqimNPp2YkkukX+6jweWrbKM4OElJ6x2gxHRE4YozwrOhGfEMrEoU/vVOlpusaTW
/WZRGLJ9FDDHhEJ3jSaghYrGyw8uPTJj4OuyMF/Yu/4ZJRiV3amsf65rbawh6kTB
mKOzIg9ezlEQo9iTB76NaF593rjXqTQo7HoD26K/oD8xkfucIoCo8Umk9nFnf5SY
2I5d938daYCAD3DsryfwJ02OAxLfEfJHAlpYFUK4LfiCvf1/SA8QgvmZ0CSMzbEo
9AuoLgbEKX4iT3n6jacUrmzIgVtN3vKBuhIcYiMtibgR3SqxdfPYhcjXFZZh+mtz
rn1XwWkuGNepNTd9Eo/0FEhe9FJWdV47VPrCAm0WAd5eISoXyoASxKnOvVAcMb1q
8+v/4SWmH8maAMhGga3Ab5Bi+/GfCL/ff+6IqltPOme6UZRXTvF9oqXbUJMU8KSz
E0CVRZt9ON4IBYAViLXLa7ziOFZ39whu1Vf3aD0WDOf/CuQT65aLpqqaRL4gaAOH
h3M/H+vxot22uMnCKxTf18AWhgCoCK+0U/Oekmp7cqcf/UHDodMdkARFIenVrvUu
dw4J6xPpqaZ4AuIKjipyCxD/ABXYdLXtnRoQNpACM3RfedAemA66eE6WuofjlvOC
sy3e+XGe++i1+Pdu25qTLrqJfRmJsqAcOe4KhVlRuPsEQnQiQtJf3DE5LCdSYyi6
TfFxysVEd3Q/oRMYqWAo6w0k2s4vOEkyXydDuaMuT6jkuHor6tfyMIO89mXQY5XV
YABgK/PfEBufJL5uRpSE5ZBaZpG5uT+UVPonjAzlmgz9TsSKVuU/WBvKMi6Ewszk
KroWdIewZiO5Ul2uv2i3QsN80RkIFhXSto+4NMpkaapVjBja0o1JOYuoUtdClDie
TQ24xTRGeuG0RzefCBvpv2ZdRcfKKx6tz+4RUUIE9SrlbYjdBU/6lpPkWIbh8iK2
s8JWIqV1bDh+vIuTI3DEzLtRhIMRRuT9I7WfbcaAq6q+8LQsXtoucgjrxwMz5eLe
0/9U6aVUVmVTzcUbzNxTNegi1fQX4JVDgTJBA8vbuf6KALsNZ7GijjwP9O+D42cd
BxtImtch0Kg2kK4b59fkjJvsflKPjz4w8xif/s/0Qtz59dU6ic3gC4mdXRvLdVLl
Nl5bRqvExLHF8pdLjn8LHsXbBEH7WqRgGWrWL78sVs0NnjkaO6G2OR9zU4070YFH
DYTHuTBWshE1ndHq92obqzRm8JQLjniJcR89k1a/1tJULDHwQPtsRCC1TBGBz3YQ
8Er06idzIEUkv68tE91C6daxXnKwCbT8JBvv8eWJwwAU4fs1Cfye+e9Dw92SHdtM
d2GUMa0hzRd8dIUwfpUjerMS+cJAkf7QcjurghUwaihbIsQ51G4Mq/hSBwAw8+af
TOrijiSex4mmlyAd0pG36DyMhsGR8RIvA2fpp/bucStizKCZ70YJ2FTl2aQFWRg+
YF2VW6WBqds68LQd8uGevBk9S6Il+BRTlTj+ZQsADF6JyQTL8ju6nZsC1aCaySl9
ctphHNqHhPLCAzE09PHea9NvFdFQ8BRmjbmA6voRJq34hA4fWA8L8ZA0dNVMPxiC
OSck4ONcLE6ZoLHzafdbMs9T98f2fezdf7Ip5IBEe+PQvK0aOgC7DT20zsH8BEsG
2Re59Srof+C0I8K/PT3hkjJcAswzmv0rvndFQxiSlIZF+ZwPP+EXSg+YT1MDqjiV
5TwZZf5mVRkqui7cHBJWuOKze7LRAMnBnx/ssGdZ6lGosx9bRTKjsxPpb2pWlJan
pJxxkFJRY/iiK1Kqo9fdatq4oanuRS3/eAKd4m3wF7bwKdzPvbcDnWjmrytvt3yZ
UWU1Ee5uy1zgctQ9gQZYiYfacxXTtkVMRqTbtjS9nfK82L0d5jZPLG/YNYGu/YjG
N4qwYlUV+2ZyRILEhytIl3quSnUGfqbfbAWMQ30yJr+d7D7pgCY0CW2W3rJrClxK
DVhiMrKpkwlNW4bnl8AE7YUW9BuXlxRU7M3hzN7bk+aPCqasyQwV+h+wbf4KpJkH
mnCJ2jVNvqt9vOOJ4ZtJ7K41Q5JRcAYgn1YbF8jo06rLbouD5Cr7lgbfALHS7Try
+9l1/D4atKIyRFhfXKT8VHNiQWAncqt3mZCH95ySTSB1Xd0dJfKVM90V8AFUlOtg
2mkRjngkjIDeK2uGFtvQok/TWBUqIYTsfYz6HWZQ6GJtfNRsvoSjMAkMKb39i8Fn
oCo6PXOnYE6Ez5WInDE3Ew7HxQNhv5k3CGvBuXXRWbejYUcLiUqPQUAPcSuisK3S
wv+PgjWzW1pSWY+oVtoGupxDrLspkQlDThIvonCia3gwYdm2WhnX9DMAVb1VoZk1
8YN/qYZOMp2yAOpq3V/6emEKhjkl9/0oJaLuzjLhk7Okm3Y71jGmRGi3aaTDd+zz
KI9otXcrIR5GdUPYripTYo3p7slaMa9BAMPvgY1NzqkVhM2/HjjFlujRalu66qR2
4OTqYtKG16KzpYILhvaM1YgKYWD/ikzRYon0Jk9+BDRcRpJyjSJgrQhd+LLzn7/s
y8sTrfKf5HI/mwh2Q2fQVvSSaGAh1XctSvIr6PtPhbvzlqMnnudAzkjN/Anbg/q/
uw7lE7Pwb6goJwOindMJEywhnjasJPNvwHrGRxsJAoxq/sNvne0hwdG1s0D0fx6X
rNqcGoEfdTkmKrhaqTTm/lCQzB3OndrXmPAWcRlzxPp3qKxK3iyUjjEpRbALTfzF
oHxRtKan58Yg3xmma3TOeZVrnx6fZujYpAjWQDosRNcBX9p/otuhaoMf91ToZZzr
RUcNRZmAcQEEnmQIAGibsVGLQHr4J7El/w9AHm6TCONOWP8apeYSZUE5z2mGGSfj
NI/rLzvGFo3+lKnvYriwZmjuPqIKDF4j4x6pG0wKMv7XwyuR30hE+HkR8YDb3aDl
QsB0+FemRfD1pmUHMilkLaTBHcSElzKHQyLg/nxooBG2LggVlisNonL2OoJAIsjw
FtVW8q71BzJ0x5qL2wkjechBkVcs8FT/Dw9dj2+3VQWTpjJSJbqTULWpBd7yvGqH
8i/t0cjLUzXv9pFWMPKZfSggpBaMT6hhk7/sDrmTYpeY69F34p3NaAW25AHH6P00
gZ1D6unTz2AmSc0woPJaW1cDAlHfae8pv9SHlpHxVqECPdC+wHYwF2OZ1+iRXsUg
h0FPfWOIz55wTj/8iHtd5n2x+OPrLUzvln8yqLUpN+HZWbCN23kqMUnut4+UxfXU
Mh/aAnOLcHBRdVip3DpUI/WPIKBAcIb9VSDKQ0slkE9DF/hSgZI7szEHQikjoU+W
HJ3lEBHurMaoTitF8IiCuZf/mdTSmgHjPG02/QGGyNGMjgoTxd3a7GULSWcJbbz/
3CoGYLOs9aQUuBV7wmZkmnBC00MYQjrgdcvJcBensX0hsGoUC4lqwjnx1NloCqfW
dIL1x5ciOPqt7cYjadFaY9yUWmOrOxY6K7XmiJQFicwlCi20zfMespgQIkxnivtT
7ToNAORrsqurR2eOvXxj6fumF8H3O4G0Fye8fIzml+C2w4pkPqY5s0D/4avuTZ0e
MwzQlyLI5eqOYZdlKpx/LpzBbTc/8HIjhIeka7pR6Pt+StSgyxeSQWO4Buz5JTp1
RJn6ZiI1Ircq7MFpZeaelv7g3zNoP4e0e5wFYuQjwRdS418hXfX0ZV+tUR+YMDRQ
p0NXpvYLulIau6RW6L/l7cxPbzfArNDi2QBbhEznCg+ZJCdqu0ANmTrWtci8OE9k
6pGuKUy7D1C9Xwc8euVs8gjZFKJHfQkSD9nuBJB2Vc+V5pckjTrXMnVS/lmT2iRZ
CE8N5hmqJnzoAH+efX9+IGtyybG8u6HX7oxOZW8l081UQ38Ibdx4GZDKmgCyIQ/4
ZiaQrqoHtwyNLw3NjQlj5+Lc3PMYb3/A6FxkbL2c9Grzp3st/QEEkHQq/fQ01Fur
TO/KyySldHQtT/NBLFs9SEoUd8yUSON36f5fziMtEdfoY9infLNbPDd3oQfXPnR/
aWAAJ2DfIh4xp3uPWhqjy3i74qpUfQLQDF79olxhj6t0It936A4O39ke9d+tdCN5
5xISvbyUPj4BB9DUhOdPgRtZA3Qs1FO/RaI4rKDjLko8TQTEV56G/P540sGTD2PX
DCis3NQyJ/qBdiBHV9rNMStqlmwgNyjVqsWmwEX0hGac9A9RqebkFvjo/J/zJFVV
bNPyh8ZdN1/moP5TTnabKnxkMhvMgL++dtbHfCcUF+QMa0W7BMeFOPM1+AHLTlFt
2SRBqpIPzvz7vOZVf/36LR/ajDv5w38JRFgUauw5op4ZcVJ29CyAh58aKWSlb1Rz
gKbmxa43qcrINg+WoGlUMFRlcXHySRHUE4vVuWtv8swC6HFvhJ8nUn7Rrm8qAz37
Z2DKXoDv5CsRer5ZRa3bT/KTx9i//sv6pXtDnbxkzWQjQcKXt8BOwWtms2/ZD7Yu
YmtsaE8nq1SIknBiRbo+NvsV58G+2OZmtfJmynfCxqZgxOYfujEGWV2BWkTIzWub
H85PzEN4a4DGVvpy6YnnmFr8IU+mMz3E30zC64kSV7nBqZ0DaLQcmjwg3SrsUgaY
y/D85sdQzaObwzEKg60gRVx7ItPF6ybffmc5r0J4TlrZrpm01iWltkgMziU71lhf
kyymbiu1vByTV8OKhFKd41pftgHS2kbNccMdyM81KadGVxUH3VK5PsE65RoJxRc8
8OKsWjdoprdx2k/k5C63tzG3KBmzlRT7SNLI50qs4b5LsJ2O9YUjFPDiaqrBOe6k
AkaM8Gt0FyBBKvuXkngN/xH6JiseQ/S3xFrFPPer9xC2b87ZcgM5kTdzG9K2Cbth
BY9BmSGnvNA3L2SN1oUcEPAO8XEFnvk8+ezuP3UUceOIOmF+qTXLpg44D/6foRRR
rCMC6opMThwGvtrUyjiMTtJXFn4HNkKDp7Y9/M/WCCcLf2C7ql60GfyMNpf3X8st
m7oL9VpdQa3w5GTfmAnlcG47F5x1H3L81sjae2MbQfvsFUvauc6PSX72ScZ7UlWB
q69YGfqyz/TxZEIyUxHqslqxBPmLtoah9yOzFxBBiKBOuuHFefkKwcNx3S60EdWN
Vhnzj0sJ85U67QXeslAar2pLRktFXyvyOScSgry53B6UWP0KDTvRdxx5W3T7HV0s
Clus+FONRmhHwvHUBC1A++pWS2j3pW7l0N7XdhPM0O41OIdlKFOEuVtYQvXMrkM4
8ckrPvBTLm+N5NRjcTg5P2YlqsG+jljzjbBte28bg30Kzyjh8iHnd97YFVlu27pY
Bnwttyu3J8OwgsbrocF/N+m+mTIhC+ixYwOzMyOIFlnqGhZhyRm7QogS0y1HF3iV
pJC2kWmBgcxXUh0h9j46n4W50IGHI04iGFn/uBgwM6AU9cOTvAovFpHpASTcXTP/
fV1L22j4gxs3lScKp6ow4PmzKpaH9thVO8IVUuwmbw2/nmecEo+j/Mqxjst+E58a
9qfzpB+a5gZDd2g+AUGzeYEqSQhTW6HuenPByCHPmOlVBlLMOF3Ztf371fcWAWou
wNiieYF2AKNTLok5IGrz58APfvkBgV9CyV3ApVqhDYVs2pjg0oAHsn+qBwjhkTjd
kHr09DrE+tQKq6ZnD34B7OS/o4YBM2T9zZuYHI1wI+K1DE2MnAf9CUqR8OiLCC4+
G1zA+i7WF4KjA6w8UKUkgIfzmK5lrnV/hPgjxej5ZsSKZVhqs1gM6RoosweGXNbH
/l/lxv5kyTyDHvH28NS4Hy7yk0ahF2jKSlAx5N5BBJRBQEmp98FzjjRegfaneMC1
zAgQC19rvm78bf7tONOe7bjxgc+GKoAuVBPeEH1gTKW2anLSZIX3pMnF7CQFr/sM
ucfkgajOeuSaus1N038h/VrI6/qfCXNa7XEcMiXhL52OYCztR4Z2/cAD4/yDnVak
BfTnMF0qIdXL8sZlyrG77LVmZOzOyepKznlb45SjyTyGVAbmpV/IWavcdAO4S7x7
rNh7DOZf3oBejhBEVlBoUKvVkMuEIz6ItshDdlMgIov4Q2QO2/9HAnDuFGS6AXDE
HQ2gtLJ1Yh4n9IBWdKnkE0yQKPmLpxUlrg+OZ5iCshiKYhLJPjDg76bSa6tRRGE5
tWd15OB3Au2gDMcmw3cnUW32J207nuQcWhkmr/+34N9CNrlb6HZox4zMsngKCZXW
BKystgimUWG6WbnxRdwlqDrAu+SN655HnK31eH+MfTVAwSCDvpx4TQKnHdBYCKQ3
l7yU8uml5X58QqAN7wn57TI695zqxctrPOJSTjISeEgEdkx4KcwrqL5Zq4zz0wM5
/q4mpz1cHQrqzmDozOhBz0W6T0JM7VGSjtGAkwJ0gI19TNvKtGHOV2lW5XSLwm9E
qJYR8oNN1WNBZijJoYprQlvQxGfKBWdR3iSCD8DcBlySxWNfP2zOCSDK2aFEtTEW
V0CDdsW6BMXufXx6dYFrPsimF+yzT4TMKlzHD/QeXMrrhIe0cK1oRTOd01MS74DE
LM9BL3s/Zcdq/uQ3xAAPXw26uEhmU7CU0euzstxN/DVH8mMWJq2J47ENUtmWR9+p
T7qpCpy0IL7L05Oo8XmpP/GYCWfXtW/eW+7guOc12Kfez9elq8PpRaBHJb8xSpcu
r5hXhVd9H+w9uHNuPPc+Sov9kN2DFKG2xziycR/oCPRktO/NGobGpSrYRV1I6EM2
KSmWbjL3H6P4Exx/5iNzmnJp4bLEEoGiA2DteJVaGwhmyacM25f7WZtmgjSDoB9n
kXW8aJMxgOKSPZtaGTXDRJm0TDSXpgGf8U44YL0B+fWj0EF6Ru/YcOKmMrtHTpHd
YOeG09UpojYBiiKlYp1Fm3cBZD+tP2BkcYI9ndYoq+8jYF6kZIYnNMLqWdOkENzb
cb0E3Gvr3v4Fkh4tjKUqYelox2w1pyvV3AYXX5mpkadmsWdNQZSfytvCrhfNTtNf
HCA1RM3mMirHHg61uqUICHyTNqCLQdWOzevoyGp3msFHEhTFEyhE5mP8EnL3SDwu
1OEQO6M6RAEZiuq6qgX0+y4oWDnqKuY2cGneHfg+P96KYOmwBiyJwpDcYbu7jFx+
DKgnrGl4xs3Om7EJWwNK6sP8Y7kd219/HNwlZyZ7lihmcW1r1nyxINVa6yit+ArH
p3ia3//IVVM9rKBdbHy99P52v2AwNNPxKbXa5wGzGZ7Kt+6MKDfbrASWYACBaQn+
PTErQp1NVQOOgK2fZ53yzsoCYs/hzbRZH65uElR+rZAXkPy+Avq7AIn5SMdZaEjO
914RF8ouVg+23tecDIPKRD9FLFUtsDfu6qFJiKE76LKWS1Js3vfYKEWPxkoR4Rfi
6Nbcx9bM23eSTX1lWPE1OZKrh3h4PhFGY5yx+O96pK0MirIQ8FLRVbN270N5hRWm
NRMRNNnEUwdVHJrUNR3KlSSpFBLiCjP5FFafzfyFMPHct5YUxBVH7UgSyJnypP57
iwDg9k7NtNT4FI2L09Gkk3YHcrmMOeox3AqEkccGzxypO5vNOA8WKvzJPE7WYfG1
Bw7zHw7dnE4vN6ZJ2xHuc6pz+1O9zK+4UvYgu6NZXh5LEliMkFUtyn89AinEsNr9
Yy7fOEr3q/Nk333UzpRZKisTDYDLfhSbH22GaacEGhhIhHEQ+uH3Uv/F+q4PO9sO
cAUhXNVBdrktJ5QZiS1/B7Se8kB3faVJS9dcRNGz34cTwAV3QPRW7I57W25+3cYW
kiXZryiepDVlnWJrjgX4xodEpuub+RvlUbO+0e+bdxZxSjGjIgoTNS49TYGWoTll
vJuX/psP2XxdEO5lTQUaIQq83LaG1Ws9l8QN7g/mmdCvbdrgGzEgo+GCN1D7zLiw
Y3KAtguzl34IzUbLCINC4VZk9V2FWQR/CA++gE9AVVx1/Qq6M6hLBlXxGeSdj2q9
KctIVuFAxsr0+mI5BYFhDwnwB4pTI2PAf56nxWxW3SEUqYD159QDFTtAD1Bj56BC
F48s50zBhDOHbqJrP2tw7PbmezyG98h63aEtEyf/Chd+33LmfdoAKezQGJFHKr/Z
Uea4isLYvOgxJf93TngMHwKt0B5LPgWJyjzpCOlRxJRJYcPd3dR28DMgsvzS4I5Y
aVXv5M1vB5A3yAcq+H4+KqBL6i3uJWRThKvo816lyvX4TwoW0gKp6YrYTn6ZV7qa
fWqHHpYAexu7mcjj2eIkC8KdlR0NSX8I05b9idbo/Sgr2CpVAgHbre0IpwQsWP1w
5Xi8h4cYeRQbD815ar/44OXsLVIUT295XsCiddxrZfbAIiM+P6eaTfwd2zxo+vAS
EBrt8KojyuRbSPolNb1AdkAvHrsMFNaXJo1rEuNUQpwtxZLjDNu0W4NPpNquwh/Q
2qPvYU0sc7n1kWGvR/5yF8AKIDpsDh+jVxzp/0MDA/ga2ULuyQDNmRPPLBWnkNFl
pghYB+nzXYZ+SofiCdQiBwklE0XI+IXbJsjnJ//JWhZiqglYXTYwpI36jZF2n+G+
e1aN5wS4LgXcsAhwGCYA7K/yaQii9N11j4RbLiN9HOVOy19tMFCIH7jtCalqmcRF
R7/7fDvPsdDYx/MBJY4EAsBO+q4Ce1cPBXoz8aN1aPA3IgQLvh5LnC5+cKfRMwEn
t0Hzp1B+Vx2Sg5BhaD1zoptmxNOFfia4LCR/cItzzgFSg9nLYnYP6bqcYLmsoaPx
zS2hNI53otHdXOSTM9gplntzi+Gz/hIcEQOdBCRVtMs1nssVqk7ZUTiOJ09ioxg8
4++nX6xRAOxAsGzDSAw0PugaK6oNG0BWRLKlPSSSXS4tu+Jk5dV2ZIDYMUHCS9VS
3NSwxWsD/3oCMj99Pv0tOYasMOtBkybyepY6IyHHdUZxEQBI0kJQ/C6TBOZVqa8q
V9F8dj9FUwatMjCCv2E6G1fIRgvVrocHln3/p4aZ6HAyr8tN7EgY6odHlK1KlNDd
I/nL2bfQyhYI/FKl0i+W6N1EPIJ6eTEGD+bW4M+v4Fb2aZfQJRGDuSzQypKg0QhF
fuusJI2sxWN8P8E5Kn6h3FbJgv3zoTT1VCQUXwOsU6f+RdseT3S14HqOBIf3gSqD
KbXOfKNHxYau5AelThWaEhJ1u1nC6TtXT0np4pJTNU/5O7izonVoS5s0DaGfmh3t
xVPuOD/mf6XDdO+IKgYwMiyjaNr6PS+1aXgoYSIh9eNoM1V4YZmGpTj6YwQ9tjgo
1AzuPW6f4i6ROoHg/HoqnGsa9W3ZGbcVWSTiVrYs6IO257D8qBicnlHcQA/O8c5G
UTHmWYi/3H7tevQts5SVNhkyDV0x4so6bYVCotKYhBXGepON6f4MZt817dq3NWsy
aQS6usQ5VNN+1HhwBiqfuz0SLu2LG5pY2Q1IF9N4ehVRwwEw+NRXYJ0H7JWuqnNI
lAD6cLMHl+CqymqunxFJgfN2M8n0J4o494K6VLnR/g79LVUqKpmwBfJA3ARvQfCK
TiPcGPVXxwQI66nVridKppG8HnoMSrUUozIYaDC18I0/ZFnBrJhzd6HqPE4AQa/y
++B/L0VZs6a768escpfhTpI64jo67aCTkjkZOSvdt+3wehOKFPasxLF9c2pPfb0Z
I2UcWBvafCl/Xmp52tYVTpwk689hRvGro7Z5IGp4tyRw3HyduxaP9On1OdyjTsyC
f8JbB4d76nTYRTgBPX0ICkcTRlW7SGH8qLqxfbV3hSAbgRk8x34sD2EQ8HajpaLR
i8powzQBiqMas+S4Ci30d96IZEwOZAf1/2bw1bGikkHgkVBLg0DX9iMQ4VP7ywUb
NfLce2N5bqzV+QIM7DPther1C5sylVLfMOrzK2hN3jq7IaLhdNOEJ9g2AnXFEl7G
+E35f6criyUqCF5nQYnycxDhxCcIE+MspCb7PlF6WKFnjmtuA5uq5ODrcpSjvHfC
umw5CpiQ9dURdhJDcGAOg1rM5fawX8nIX51ajyY9KLfVWF68y3gSY9OLAoHT3JPq
LzaUNCw5suiUBeM794f1N2TtUDcGr8QsbVDREf9s7sW8JGgWEG/oHWEkSfj7HrQV
qCDTV6g6avjzNyp3dfNXtEGAWRA9xedML4yyAFXnFxdSCFP9AtM4fDqpZn8kmcX5
vJRQ0awRHbgEtuwklKYPSf2fd95IuhkAk64zN/mC9K+jSEKFRALImmeT8B3KSvAK
/5c91FrCYugbtDr+iLxjh9DayC0jhJdzpgtLrIhnpiwF7CEawcDNbRDUbp0Vni2A
nZKhwLW8Qto/0TeJ0r3Az36QaWJdKV/+vfMFf9ab46gSSAiznyCBs8HvLI+h8Qoc
zHqL+kietVWpEdZJRfC3tHfDAs4i3uYtXy99+5QRzDiGq906bVdC5cFIoS8Te+65
9iPryhVmWET5TpWoHag1bKLbxyq+BrBBh+OiqBIGGH9I7bHxUcp6ZRcnUbAXZKC+
EF9uYx+uCJX1OjM+w/R94AWAZHR7WA35QoQ049DSlAxS4Je0DGfQWEpmJrjJf1l6
syjOcF+y/70vSngXb84LU2wGtVVFAnkUAjvDziiHKV3S9/hIiEADFXVMhLS8p962
zCIAp+NOQL/KeWzLKVU8RyiIJiUBBLZXM5jhH526az1kGcfHYbmpsNg66/NBo7KR
GEfWiiAof6132IMFGDmpBsLXhzExwKIdyJuQHjTiywHbmPu8GBEMmHCIoeB2O1nf
EYkUkH8LY2+z0F2sY4EYEI/sxaVUyskVc3/4oz10nYP0VdQQh7IwBeSoniqXEa28
QD09pzI/z05ATDwsyJqqe+9JMP7ZdrN+WE1RDz5aUHXlCKqhODByNewKFWNkbJHo
F2Irqkw+NCPicqEhMxx7gNsfdxNxKiy37X4GD3zex+IFYQ/+ZhjnKsBYY2kdqoBt
xyU4oqCmPn/FaG2RA1w/tgR2pihbbn0zfYM9qutKULYrXw4oyhJd3dmJpCT4Agin
k8uJriv0neaVT0j6UXro/h29jPHmxN0DTuHFb5NnFrFPQf4BUGXhcM5gk4VBv81q
EFDj7xPgiUnqWZsrOUoYNJoZNPIF0X9WJkAwF1CfoEW2tJTPuHi6tDSnar21BokR
1OOxHl6ya7uXjDfSvApDMw2ylyLheJQsM79LU+WGl0qAzBJqeoKja9K22ZqTGcX0
L0K+B06XE+g8LL71dyenxpzfQ+pX6VL5V3sNdpAhlZo1pg4D4m5JTSnzyVAi2KOn
iKOe8Yx27kMAWCK5F+UVnqUKECfJYLtdFU1CjoRgqNcNYENLQ0XCxPy2cAizYeX/
+/tnql6VJf7ZLKPksXnQYSzp2TGC2SF2IqDQT0SzYRN5bENeSTHf6fLa4cRXCdNW
lrNVgZjocBY3X73wbsx3qjjInXAwDCyY64HdcPy7DSGS/ZEUZ/l1NrSsuEls8KMC
Xv4MOC/NGWielXQHJJmIXHcReRDB7AmrLMyDZWab4IQsL2Nydyt59gAigb3JzkuU
uM4Urpggjt4yZFZXQKVIzLIb6FOPxts8G+brAk9XmS45hEUqJd8wcMnBVhR4qch0
3Q4sQRKDFVIKzjYAtUDx7fGTKoY0HxFZLmEz82vj5TUmZC4xldVSUd35c+4gkAQx
QoMLuqh07Tw01WWYkfZe6DMqCSOPPgvQtyLDie28NUnQL5gFjuCAwWkWCPqwlK4q
vlPDVWYqKKw2XwjHTh8dq/95NdpEsHAbL8AQ6X0H4xa9u5HhgL3rwkIQGWbQVBsS
Bok1K+A9xp1XQgt38+EEmCws+cEAmzLzeD4uT57i7WdVyCTt3OCjm3KAvdnphAgW
s0ZYAvtHXymKmdJ7n1FTeOFIbsryp/bjUQZzaDoq+OfP3fBRbEql6t0uhQxepSSx
3pO2vUUx0Zng6vX6z0TUOfZiwsjHzpZerv8x2i+ihEAF+GGp2JAbC0yBZ3qmWGsL
hsoM3eye8K14Lb1KU5lrxOcJ2hQDHevgMQLuylKll1o9zENx83Ku8yftH8RPrwig
UKArzYE05qLF5Jpq8REDck+KPZJDHYLnwqZmsCtsiMw7c3BbPAQKwOXMGArkWHry
ZBPfwq/pHhWD742uiHQJM/fPt8MkNupKBwWPrJ+nhCA8KJs8N0F1H4SFfcOrajbs
YywdteHLnFdz3kN9uCm/z1CTSot7rrIKRhl3EWhOTA4WHjo/AmQIq9VRydunueg4
fHL5WT1zCkGW1X9kbd5bgNB7VjNiquD+tlVMBcXs5P/lmTZ8tdzI0mPc7wNm5uqt
PRZYUUrPcRCWg4Yo5RqV/WZiqQw80lmsrPYPchriPU4ZLtPbc+KgEwdsfwBEC+bK
MrUvp42Mkud21aumCJPrntSJG+pnVUi9FsYRpD7EgPpz/16/4sk8MxZkqoLUF5hP
ZStfm24nbYVPDKpwf2sVLsxAWW2uOwMT9AjRIpPo8NBrrChqtgwI2Gt7+7Q5wDOL
nXiqzVYu7kFpvmSGOH1Dm/VvG/3iLJJNG6V+JnPpaXqKmImMkrjqIuA/WAt9JUC+
XidPoNVTrqfMsxJxT8SRgTkpAgnDbZTNA1WBAxhtd33KTQxx86Bf8SakJ+Ri3qQv
NhDa/zyZVwYg1pNvJHWVMvVAhFDIoD/xFcatR2eClWwPQPPJjCC6SzGlxksZ+0G7
a2LVjQnR1ND2X4EqJk6Xa0pag4g5SRv1kVp6/OJRB5l5JI/bSyVwh48yf5NuikwZ
9XlBUktP1z6vRWZY0SKqCajyyPf9y9QWYqxeSUgj0qD7yqQL0t90ecy0lhPR3I+3
kvQ2DmfmvIwJ+wOn7miM3qMMQ6m0bhCLwWCsPfSks0TfjeqQH2lSYda3Gc75UB12
RQ4Y90+msYkaUgg1HnBc3B5a2vfeM/c2BiouixQkhL21x+IZT4J4CyHPS1xhkGrn
0CC6X26cImjL0VaKIlly351uqAmwYZcSouhufvHwZzZH8lbEVRRKTTnaAyLtOJEg
OW6R2/D3FUsXWb5+7yteGHWxp2CqF2suEYNjZWTY+ESdkQZ5qpi1ge+biOpzLqiW
vnC9x05SPoLpLLWL2Ig7j/200Hd33tbl/uqIOVgbS++DPkmhMYrD8jYULjAPAyF/
Tcjye6RRBAcdEVmNyerTQqZyJ7iHlFZgbmRfBqDUoppBbs7RLewcyxNLBDtmLlFG
ZJTsUBMtF67j7yRqlkuDWIbUlu7WJ5Dwk4r7oQCRtNdvJGpmadVOU84blriIYsa3
B1AbP7HphtPY720tw4a5APxTikR8NXy0eWTVhiRsodJcMaZCmOGqcg/ma3dyRdCI
JwlvvOJth1w5sscIQ89ALIft3Nqm06dzNGXvzgfsswaN4yQAkQKPMvj08PgwgEdZ
jGrgjP5oyQaV/hTMsVM7XbJxSJT21/1P2sVlPRFwkLkpSEBmSEOzvxQFglX4nL8C
m/DMVpi4jfNPtai0enoP7NA3QYsIo9HM8xtAeKh8D21eud2RBfBYLfo8Lr+0sMTc
lgufarLOxdoaJzu15vOZ3ZoK3Y9/jokytmXZIfkwDZhkMpJZoZmsRUZJp2KV635G
c5SIYLpekIovhSuuye23Ri1HJqrrrvfIPf7U88PoDPx2k1LLavkPQVcBWbdINrG5
+t8UrxMRM9VxTBEOsBWb+wCRIwVVosmlQjXALg2j8s6kB72tCAlakltP3jyyNH3K
yks+lBHjhCo5DKn3bktrSzG0gNRC5tiF5NSKRhIFqNeAN1q0Fzo1UK8fwe0dRCIa
fHjzznSY+7e8GDvX9mjCCh0j6NLLjw+c8ySe+LBkVxP6XdJg8MrK0sAeIJiu+MnL
q0T0U9pB7bTlRl+ic/UFeVb2NOMmBxpjP/ie+Y+gXWl2qQvVPJ3tuLH2fewKfGEA
1Ie2swp7ZU3IxZt4SslvSE0/kkz7tja+xxI+W58bFCLUWtxnVzvgaTRyl8VgW9OA
PgpPAa8sUOl4GduYC0cEGONefoIQ30Ld0FnuSgHtlHtyHDU3yZJU7svCB3xOMZN+
XrJw1cXhuX7/aAVpsF15vFyuoS6QqCz3Jdd9yhjaWkTcNN12HkyIE6EGIFT5zPAz
6qgFXRxJr4Sx0z2rKReZTEX++YtiwHjGNDbgwlfpxFeEXW25ebA9PaLH8HrIBcrw
0EZMG2s4KKtoVevJ8KTZod3JauDlrauZvkBt4+4+JXhNa6x3EklB1xIfWe6DzLbR
/ujVuxQYrhDMPtjX3fL2w6tpdygIZ4e1ET7dbv8W+xh0U/uqF7UkDo8pa/R1p1Wq
iPGxkGOlARitCq0zmoc6DvWqpCTFbUa2r6SRdgadeOCrZm69A1szxS/3b0QVqYVr
2KODLdGAsBde8RmdT49ydnbk8pPwoDx7tVVJHuJT2e+M+dKkoYSgoqzsjI93nD0H
9W7vqEXL/QdOmgtWtSh72tvNz4ZlixXJfxbDDAMz6ppu3YthrW1cG6KxuznP45DZ
ksnTvU+WRkf2udVSGSZHJ/VIMnqqT2S5cbz579aBduAHC7XuBRpwqYwDqH5B6Nc4
w+s40C6fhBX90YTYpXvnkr5orTPJKBR9/DOfaVItN3MSxSFPTCp4uxLu/a3UeiYv
5iihgk8Hq61VnPJDZAMYn0Peb/QvZbBJrpM7IuWXfYZYJKKvgsZqwHjZp+PmkqYl
2bqc269n0D++3e2iE8BxrRiCqD+WRghS34BU2wIfliUGRlK2NjbNccj8WXRMG50+
CoDUEXxp4Ojvwm8r5pYXPgYB5AKO65k5Imv7Y7+XvKvzcPePnZiR4KPOSrw2VmCP
H4eqtJwbqmCbunqiGd3Totm72PI9N6qnb57kOSsLohSZyzjEf6P6Kkh/veTXaQNK
e/FacnC6AB41JTpCSXVndpfTHIdbiWgH0juTaAGMsRONdwOgfJfH02Qu6QgcAv8l
DlGprplqGdrNanSSowlPTrWXHGtt1U5mXKuDpX/EADyIhj0DxQ0fGP9EVgw6lxxW
60/0swcG1IwHTtERYZ8kLuszuxc+QaO+jUy7PjJpE05bh4RRUoniX70JXw1NBISd
q34+RKPbTu5yRK0jF+vn/Ojce6/xy02969yRhWjUfHtanOmgXNwAYS3z8B0GpDHg
7FLSoH0m4oQiu5+12T14vV/JZaMEF/IUW1SlwI6iRtU3diZfRu0Axx05NerQ2Yaa
ZciyxIoD1rTvUp49Vxt5xZCofvER3YZA+3Sihp6+/IoVghs6vD9c6Y/OR2LALjUs
g3ZvTVVqkgltCHmicCRxdT+gk4ma4pxiDLBSV0G/0W073JFNq7GVyxrk58m3WT7t
cLNUj0lU6oH9vqm0g6X1l0VBF8hYOMYEk2BmROtjYXxQZsb6eux+SmNyG4q3YCQr
sHfFmbhm+OBlJyz2to0IqIl+H0Oa016NVGdKPWuC6B1sYtyzOcLAupyBfmpZVAgd
USyOrdeeRyYJgVcjQ1+PHje2xIzSUk9ZDam6U6q/IuDvJ55PkRT52hpYsrStxWNB
hFBd0ckknKadE4SNSNJnvhIJ9m90wcf0mBmsAcgT8FMbDbae13GfgAmDoNlwOCiL
+naK2FRNc8pcuqSzZUqEFheAqNNYVU0yHh7n0X1ZYABgeMm52h9dUSIiG1MrDEVZ
Bd2Ih1JplKGjFsXvIbJ6JEOqJ+15TKRiI2h0aFHFiXwzj4/g2KReQTesTiEIAJFs
I1Y2Jx5uFVj9GPFSmmL0784IO3O27lhIF4xWFYoGuVEJPTTaM6TrZ08zRO4xDj3m
RQSK2WpPZGRcNf0qMAvXcDY/9A2Zp90OBXV8OgiWGso/PDY78lg9QV/jOaLpg3dJ
XEdO7QczA8zReDD/tNIHE8vAmE7x47m0kwGYaCGLn9ulP7c0wqeaa1taIi4pUaCK
PkcxqplRPNa0MH2KCbnS2L/Yp2b9iwPDk0gHbiosxzgleFKGmOc7zKf8UGq6MEzb
c4XXNJfobT7xHoSavnqcv8ab+PKQeetKx7FSoux8WkvFYtxiXn+U7z04WW9NfhdE
eTNjUdj8pCBl0DE48nBbf+jP2U2Pzh3tnLlsxk5s/sruUp9EqdgAqbE+Pvdo5wiV
x3f+F6IelSewiNJhIlyZ0Ptae+Kzw/oew2jpQXBhxFVEGem8FUHVr5EFl/MpmiSV
lvS72lG9pKAC1watlv9GOsDnt52q5TvyKDNyHIjH6ZO1kfbKh5s4XZu1XJCZPFjA
ICKvVYo0Pek/qSZaeDjVEUsbOP/C57Ao9m4zb3BG4Qf4GDYWclB1RB84OEvlhdno
Si4b8H2Lyw5Qyxnak5U+dcDctpMBJcYSPSOqDYo7RUxpFfX4Lt9rRREBxAxj0E2q
TYq0iu53Va0bS0SHi7pNm4aqFm6oaZsQERoo/jBWDs2kysw+pg4bG+ECexMqrWFw
jkNOI3ghhRaKepzNwjp5JLFPfKot5P5tMRJpFzKHgUWvTCsOzCCzatC9k2UCxkZw
eZiYqIg0hoNVC8WEG+CtUOYAaxNrzXM2wiWPaiDOjg54wQ3tY7zFb0klh8ivBxC5
XzDo0IclLGM1mqBs+2F4Wqc97G6jeRtLmeBTe/5AFsoUnTpQ2AelsxHoVNx2Q8NL
6VJrW5P797FXAE74WL3fDoOnhSTndxnfaaAsn6zyvXLHNONFT1trDP9lRDgZ/ZFk
+UUPGoYAs5Tv5fufdnuwLleArted9eKBnR86oIAjAsa3mJLV4B+LBPNeNPScWtWU
sOe4Ky7beAmgb3rk30rcOxxjIN/K+FF+5zh7/z4DhG8F4y7SD4wtDr2p7xni8hmx
WpVNZncRTQyJAz7nsz4f7y5DViIoDQIEhkU1gEDz/zKQuzyUCgXCC1RAnJqq/Dir
88LiAx9UKNm8+dpZ4C10mKaS5f9zBVt2O0Ib1WY4TPf7Vp5jpB8rIYf7xY+JI/6+
E/fAVsMXMB8qgUnLkIIx+yywvsC9T+14RxhjSXPCOqn2wR/qLJ/giBnEk208EuOw
0e2PE79iwL2Ek5Qz/0XCjmIfhXByynLNkDnioHpVt5IUEujx5XVRebphZy35/02K
evJjNNFQq39GPLTybKyJZEZtwEi105+wYh+s5TkPUDrTrdPRmirG9M010yrRQ6Ft
70Cd+jlBnOweSHBAzZRdrSP2RT9ZwBmUCzScvRyw2YEsO7a0y/CgvVK2y9kQmJ2R
4Krkq9MiHw5Tb79iDrcTf9dC2lfB6O7/+ONLI1dFKHkv4UI0Dn/mSx8eA5qng8V4
KAKHDOxQnVT3ENMrs4KaxK83WAcy5lKSY7mEFLWhWgB7jFUlix9ZZse6zgIy11vO
f5aHf/V2XmyGJIrH3V7yKZVCkWNpOhthnSdOdJ/BR+4CAtlqba9F6OYOWhQtptsn
hVBSug8qIBQTIZXDSYW0GEjOXpLF5vn4TIMGFuol+5BvOYu3kKB1fMuHdje01O/U
/8WcfSxmAZMwD+MV6bEIZDpL3Ihe9kbV+jwBWD6ZJgXEIQpnm+HTaoc+eGO2/vEu
vr2ibbKOh46FRsvwZxokbq1diK7wTmsUSEeGBHjJ9BX1XPcRWgRtBiDJqXFgLjBi
biIjt+nWOh8ORKChxe+FvR533iISBw+nzxkfiKDxOWYEt8s/MkxwziRWz4xfUkNn
+Gl9g+hAUpUfzmr+JUhUR4PCus1BPxn2W+LxrIgoZeTjzqExqwvex97anRDBMY0x
knz2wVnOJiVSE9/KmUxDNCJXLfXQ9W+y3IxtDZuo7UXEoSbCiuI/7ja0l4jbfKN0
lFFyhdX3N++cCta6Y13hcIlYk21KcGQeKL6Z1CBe/MAj4G+rIbY4NiHK3VFYbldA
LanbOGtr4GitCLLAZdyoYVhtGCoQyyTUt5KLgkj3LoSB66wPNQay9ttIhNa6gW2T
/QJVHU/xXTKaN2wSv8HyH5ngKIYQR0JRZuVcvvRq1QZNX5CN12JnkS7Lp2WZ1Xfe
fXOZmDZTgImKC+OgRfKDWB1mvq/d0BgjG1FRuJbgevqPy6i82cIPGw98lBGhckGX
12aJniF1/hw6Z8w6bsXE/AgqLQqMx5ug+Bdodkilz3Ixu+sg+rPurAmG8sUO5MbY
3PYrt/PPF4SQ0NMZoKpbjt5sq6Pr4S8WEm7JnB9jDz2V0kisvX2X83VuE+KEd/p8
Qso2dYwHBNRSa0ZWFtxNQNQjqiLJ6q1IeGuO47bwVOQQ5NonzwTxcPZU+N8svSkt
2uzuXZm72XZ70FvQq0D8XPgBiS16940Bf5KVUpNzoULU94YzpBAxho5mqZnDdORc
n/XzGmQv6kZEWWU4dQX00gksTEXRAflP8zDrt89HlsU3tkZ5vOx0rr+S4AMlp+kY
dT09btYTMk9hp7q2boGW4z7hDWG5Jb62Zi7dPX6Ao+viBOjqwklW1EZw8aiCClEV
Z5JPBx2YIVXnqskjsURX2tsbKsmpX4/Nycpz7R5JQnKk0bwtNEqFWOdq+0wVgc8p
Hfl0xJ+nio1xgAzFJ/+GHeBNiaIwrqCrwcHc7lNu6r6+Y1KN9/dFGhzDeMXGE7DB
+IiWZO36nRyi6KEtr8Ly0T56qfmcDzrEdbY9efaRCO4CthLYXBzlhYL8tIa6u78n
Qiiq5StULSoc3nyWypYI4sa/RQk9c1yHEhWzAeilDFMasMzQFAb/brLaCq0XT+Yq
YdEq+p6KkdgD3wdP7w8G7MLeplpzK7G6mCzcFXZ7sFKMmXuPre0pjh5tQHRSjPyp
IafmXPVsBJDEQ6E8IMvmnCYos3pChOICf6GVzj4/rOfURi5FQzyppw7oItt/9484
UMztx/ZbJcyCuMdmb4sgbyyyPi6Bdlwsya0axfR5d/k12Hw20HEvQLellA3imu60
CzY3OA6ADLB0HR7L738ww3VD7mQlmv/jmJp3IaGczyGPCDcZLBSaiVTPVAZa4JYk
Nlh1mzRRAIdAXaCjHQnWUoUmN/fiJxxd9Cl0XZptrWq0pNS/UmM9xK+2WXCXk2Iy
E/9uHZDug5pntQez/5bCE2UT5LGcgJHX3eL0ly7ZSKGILOLFa833g4dTxu6QvAPw
sRKpfL9aqFTBJJtrsOV7lzSPZONABvavv5rG6t7IJ1VVxCKnKwokvL1luM7fZKkM
LJWmjtX2aNJQaI5pRVlA3gSNAMsXgVs0+tET8qaymrDDaqUfdSsmNiaq1WRQQu8x
J7wUe37Naxxty8SiuPl8z4CJT8LYbkkrO5C76zpeUzwdVImY/L9QMjiUSJO4IGO5
W9N6iwQKbjq3ieN4q7UzxHbnwNPGY/ik/AM4b4GbC0tRXLWWQSriF/gGNdNz/c2T
XjeUg0i/tfQieWEwpY1PLIDIr3Sjp0NFqhdYxKAxoUg4FYRZqJkBwIvgb2pDdtv3
vRQZ0XtvX/6p+g2LQBheVFyTRXZVCiQIzQv0GVg0qbYP7Jy+JqOlO0gaotiZntFC
WVhUdchvUcAfLtYeRFVIzTrPT/Wv1ibt7FWYk9ERmBbvBjINGD1ROu8AOkX/7dj3
pRUMCH+C2rLdEfSj2YKct8+QXm4JIshrEhEu/Q9Wb4flw7YM10OAKdiWv+k1hWuV
MrIT8eFj5LhwLdUOUTpjxFwXiLuf3Q7uYr00ITgYjfvjUtGD58vIOLsZM9NjUm/s
nNPhtm3ThnYWW/iGBZLkX+Kl69fIGTw5R35XGEGBLwWtQqxR9AdLn7bzGGUAhx1R
sZZaJuifnU2dLDchny0pv0O3YI86feXWs0gz0vhNu1WhgSlg6k0XMHh3RQO6h49L
s24AvsbjHPHHS/x63L7IGAfRMtx9IdyCE26oNtBGi9nw26kyrXLSzA8ddMtLEKzP
nvakTkcyHraI+jvBwjx5VYCXopyEGEBgcWJBgqUhseY3zJoxdeWJPK4kUd3bWb1X
2KNZetoHmFWGvYWs1RKAfoNdleS7mWqE49qcr7uT9N7wfQYF2TD3enb+VH+FaElU
LfxXaW+Zk1cusFcua/UILRDCyJxU9Ofi4dXumuDwu/vXIddTXWq9ZPIjTDmkxZlI
Rp2ffckStJ/RydOrT2jDuRn34Tpwso2MfKdUaeGgmEwwt0UFUjwaIRZHiiH05OWZ
fVFJulL7kK1nfeB4TXZdY0cTC/JKwN4Ej3QCLwebNhZsPgwlVNamHzUNf7h+z/LK
UiUBXE8Vp44Y6gJwy0lM9/xcGPaNrYT80ncTkw4XA2rCww5HE2peSWSBs50HiobH
z7ImrC5m0EeGKjNty/S2NheNw7sGHMCncUVXmMc0w/jjC+t1b/wr71yHRYE/mCvi
XjzGV8SqxVTM+WTqOs+ttBeqEsI604I92nNYagjvUmACMBzE6jwW2BhWgwXr+gFT
p73rBJ1Z5XnwPPl46G5mHPut32eglEGjTlTQ7B8Wm1/y5eEHJP1hsCreBc16djgC
8u5STKJJ8MUsDaJ/0xiuDjXX1XLbdTXsmNparBVdlAsMIJ8Bsb7b6gPa9xpzYnup
g1Uf26cQgXgmtC5YcAG0uJpfWfDZrf8VAC1Th9EXcZgHp8+xOz/1p5kSle1hS5qx
C4F24nTi6eYQ7xn2SkwiBCnA1qFxahVwWlo0PxjPC5zz10ERjd9XZOXl8lLwaM7t
IAmLKstu63q3qPYU0Za32fmD9T46Pr6yGTOEEss9n4hD/UaWbUIWAku2ZAk9DEKd
63zKbXqcbM0fsCXqzfB82Oy3sAEfnT7jRTChO20GIPkNHe5JMZlbYTcDkvGoC8ME
3E73OODO2hwjnxGPH2ANrfpdAG8AAm3YKwHxEDOGUXOEcVIkqpQcDk7ByZVynB2R
pRJdXwOaKPnJfWqfGavjEVx9CF0qG3mRTxAzK9c1OB3+YSY99KBZbdW+VDHbxodU
/yyvjsQi/mK/D6mAzYcfdBiNq3ln+w9QCwtSZa695QeeFtPjunKNkrWEP+H2aDZd
No1VqP34+Bl2HYci9Mf4Y80E2kvlf1Hoy2HtLNrl+UliYQZs4tqfywWl0T2CeK/L
acHcABfiLCqCCtRsvy+ZcgDygSkjvI/LaaxPjzWbTmfegDYtXri76DRU0bRjqmwz
lEoAogka/v4C0Q3zoEHI1QP6Io2LMd4upmw5p7KZd6hreaq+Mp98Nhne7CT756JC
7ESKNs6VfkpbqTxtLwA8BRFt2/EDzKQCjNQK/ZzZw7ya9U8jheT5MHSj7E0ZFFAX
WnYJccLdOqaaMkbNvPFskfaqcgHWBEyi5QMn6/daWHhs20LJABY4iW1SBrOwkK88
ZIjN5tA8nvxioAGCtrgRoxawM/44942yTwx9aUGNQdwcquP1QdW4Pf6bJ2FlXLF6
Ie2gUQ7Zqk+RSqc0somZk0oJCOR8G25x8Kc8uNVQHC7xJ6ARh+0Tz8dlJnaxx1u9
17dJIO3z5um4XrzqH4YPkIIZ2PMCdRVQisLhynhGVnj/sf9WgMU72yu5HFXlSrox
758GyEgyw2VQJO7Z2lAA/H1smli3SEIBYPaMh8oPSMJ63iFi3T4PPPQonB2ziQPe
OENVlne5ChfVnZM4MKdGYv4XFOzzxTMhw/vM+96bnNb2ejb7EXatBGVZ8xn4QVSo
9d6lXCESLACMKuRL8Tey1Wc5CTvGZPL4DLAh8kNxIPfEpVlZZAjSXo4MD/4TCcBp
xbA6pOjx1R51IqGLbIDRv+EO0M9t5hD+wqITaztmS0BJUzzLVxAkeoOFqwu8ksS/
EIt3p/mAyGrnn8gjf3Gpyv4Q58GbesjFZMrZuqjADFQEwbOQv829AhfcmPRxhrNo
D4jTDWytG3EEHJq96sqJN7S7ucKxANl5SNZmWYk3ehC/QnQA49rCu1XOhZTDl9G2
XpqKI/U5lQSFUZSUtDOJCKSIfJ2ZJA7sR4Wq8iCcw/KYawCCTs/QHsL21fc4hwfV
TPvz3HMuxEjfTl2yTKVdWw36nUs/8qeJ2P0eYy8PdWgQb8lsiHhjlRqMDQo9Tus+
Ndj/+9Dg3W6uiQJZFnX2IgMbdnN3winIpUUfc3vkrw6nPAwsHefR5P9Wr7sBL5hA
SqY1cq94Ltx0/bNnzzIOZ5U9jy3JaiIpOg/PKVj4LWhsHUz0H/PyT8SVhnrAcT5j
AnIlobGE375hPyzohG3pQa3AHvCK5yqDXuWPl95RMey4iQDMlLg4kCqP0pcu4qsZ
/et3K5cUMewt98uJ0gLGorHbxV4ON0VVa++Si1JprWBfhoLF1RQJs6BsIU6taunG
uo/NLy2/xMFXDadiBlstqt+PBVNASI5tKK/vo09vqfrmYVodhIZDhf1xujfYPEnd
FwYnKTC9ASf6K3LcJKMgFLNTcRK1mwd+TslUNw/wfOS3Ni7ChsAFvAp+rDUDKEWp
9Q2FLlvGHIkLljZ4r/u2hJrE0kdmBTpnSdQoAsPoFlFb4r6l+XF43uxu/v6JtQil
S2fl7lSXF69XG72du0zQXslrSuoxbOnvJORa2mpl7i1EzQ+TY6xWrk8UUcWA5rWX
bpCxNhDKN8qohJD69nmDddYsVmFJcZpBy/s3pfMFVu/atDbfKVECRbSq+FaPo+EB
d4MO5AnHkaMHRcpxPLI3YTEY2Cr2YuMTbVWX8Sq+1tOjGglUnUwpExUQe5ADLgLz
uKdX/SluZDf8iZJkMPBABwzTvqu+ldFcW5gUbxGxa/jWT4TH2SfOL/lC+fwdauqI
oLt3zb+XNow5dnNRzck2SaSnSZzgtGlVbqLGNMXTsw8xJewXEhK/rdML9HmYNVLi
WqcygQtwRjXaZbmRAq6KfGESLbxZ+pS8FweywrDqHCOxnYBoqiu9l8nlpZf5Ms6z
AuQC/6RW1mVDdK4bxKAs9N8CTRplCYfZPtSL1j73zybymDBgy1+rT2xV4Us8F5BH
fTZg39orbFP8jBH/0x+4AeRgPRg/n61be3trlSCo8nuF1PkfrmICE0K4vzCWjcoo
Xdhw87zJhuwgSRfr7fmJeNHZVD88Zz0cPNuF2yqJATHHqkew4pEun3j7rppeBNN1
YCC7F6wef9+PX1V0KS/XFsPA1RCOQZV/PfloW0CXbl108bT4Ow4cuaSkqTL7y6mb
8pvUkPjad11m0lcd1EjIiCxFjoIozu0GCOhb0/RxkMd2KvcWChANBX4JyWb7AK0O
us1s9N7KfV1R97JWOPsE+mA5ePCbGFZbdbTnHK06vsWkHWr6BRjqjtpxPLXkndWA
cVXvP4otPZrd4X1VEKxh6QujZpo4k4BOuSYTkFnPZayGNOW96Gdm2x6mHcgoYD9Z
OCAF5iYkrmGn+4+36NMMgyUZc+41tGBi4ogNkYlJUzIXiFnvd7oztWdcl4G2IRNZ
hj4gYH/CiDJT8g+w0IJ/CaNQ/I+sQsAX80p38KXjZ2AVUbp9y54KsE7ozeM308Kb
76wVbcg5Nv/y018F697B6VE5/S/iT5i/I1C5hctDTd1FGMFTvnjVvPykz1CVT3fB
gsNYx7dXJ4z0rPZg7t5IhnE/K6U2/4GXg8d+Aszku4e9ceVPQkDs+QU8ywrH6ZHJ
qbRDPiLqZzmyeUFokKRLYcYF6ZofvaK3KS4Y8e1W/r65yPWYZdjyTNBhqmtz6ya3
U4xgfXnThGe2g2gdp1yNRWnOl2nN/+km/qtaLdkr3vf48Wg1beW3SAIPTOdUutDW
sLb/xwbtn0MeYpRsHOcHZQX8CKe5iek6lpQsivdgj9GJTNlH+34VMqhS739Ln6qS
+DFxPB35g38aOE9W69J7D46ra7+tP+6DkeWSrqP3/nOOJ8E9/saJp6NZC8FCpdgQ
a6HpxOABT1qS5lXZPTHgzgjSiobf4rmC+XOdKa+1SfnLYl4a/+MsFxkWfSCpA3Kj
3BI9tgl0XWH9A/MNYCf9giOglXZcUhd/07VxuO7yW5hThqZj546Te56cbfSKdCRM
Zfb7Qpz+yXrpm7Ctg3YlN/5y/bQuItOkqJ9SvOmd/UcKYBUlvmGRT0q4zdNWn1v0
WzL9+ORDB4MnmWt2vPnOJeE5Fz+OkOwRLkI8nbGbfoBKq8AsP5dwal6hid3VR4Y6
QG+9b2t1Gypq5dQCToireTs7bIGO7+WjfEvcbbg9+oEcl2vYAbJWX8/w+Q57aOPF
AH8j08wOopIQ2y2W5bc+dtadRQmvJwlOp6EHvu4JMK3a3q/Al82ld3qe660UldDe
4leQfe2zdHrkT/EqinlFcNUQ9sMP/sQQTPRFKb9oatuJRVWNmihEhFpxvPBtLfgf
7x9e+h+3FJQI+03b5XaHBml7RJlen7WP3kZPHRV5yQauX7HghOREZedLPEZ7Wecz
byxw3HTnN3nbL4KCYQ7GHJ5R0aqPg5sPlaJ5iMzsB7wyP4xN2FN/R2+WiyaVj36O
Ul9ybmKRllLZefhzeLhNvi0austwxvvRr2cYEHsYsUz2Ps8/6mdfiH1cQx0K69kI
pSnmMGQ3xzHH+c+IxrtccCfZ7DYV46PbsL1tsMbbtKHkrnQLDzG/oJ7AZufMnTHw
X6MuuFJxaz23alECMaeZ9MpPPGolssR51jX3qwvoo4GY3k3W9PCgasl5unV69D0q
+YHFKexvZ/Cl8I1O/jQ3c9gCGWMEftGaa6O/1fBlS59hgAZlazpIhIlkZFvMmCHM
2tEGI8VHn9svBEYghZ3y+jlHEp5cH3BhUGgB9LXAI99LzQsQb+xHVD2n4ZeuWcjg
hJI0s4b6Q56ZEimvMI4ikYd7RwfLy1G8+O7aUX66SAil5A8uhbgxwRWayumXILK2
8o/jeXZS6SxkUJ7yyV0QbH0fhxNlu5TJ4hrC5cycoDyOYCqVezeJkJcw0oGfJyu4
FY7SPbcRYRZhdFsGOvETr2nikC3yA3GX7dIGzOTaDYxQ6Dv9iaFkAq5EnY744xDj
gtM6/0gDhZESBaTJo/p/u5HQ7Qc79b3s+WvhLNEvBvTQCdtwpP8+Ik/G5AFuSG7B
/RxzYLZPSrG4OdM9FqkS6vp8JtkGlEbUsLnGIuB+pJlww/4M6BKh2BJadTV96wY7
z4AeC3ufHQExHlG7OlP7qIkpQb51qibMkFb40UVc1OSVvwVIBbGyKhOrB+Y0e3Yw
YjOSPBalwzHJ2UPSj1fdyztcbksFs5RPkyK94Pa51AcmgZl8zfuer/jdKI0jA0sx
4i/p2kg+/vIbap5bZJR31OQxxMNTPZWs9xOaI/6N6uad5BXE63mmZhf24Vv51Nao
iT9W9FhALjZa1KbeJlqia6SziVLsNgkOdzU2OlCbgBPapF+qfhYYY8NEGx+8vFgk
n0GHCOcd/3PCIqZZR3toVh6qjGcU523ZqWpLK11EIu6aUJ8AYYRLVeWmJv5i/jxd
9TprpdKkxaY42s15F/zqMYyTcOPXvO7X7TktZEXLy6+A99XViqRSYZQLeydO4jtB
RxsRvEWoht9gvv3tzDM0JcLjbkbULnGKmSC7ARVGrHQLNr+HvmArejhxEkannxn2
QMM4kR4188GdUjkHW4RnClP5E9R8QeIdOLSns0RPL+0VbfiPUOGu0FLSuF/DZ5BU
7ghjBu7WLdVCZSo1/QsVeBXgJb/Njy6ir8GqugfOpZotndLFPrroDV+h8K0ORt8b
nRIGk5du1Vt1XiCCmnHH5rN5UR2xVbgNLHYrLqr5SEW1LuiQdEF5qKyixOEETFwN
WK6+cl2C3yQtSAZ+g+Rs+1mw/rOJ2holQj0dZeSDEmMPeFYC4ZsngIKvm+wlZsUi
cRaH4M7beKMpBopnBQWvqkMbu8ywj9Xi1i4seLHzxTRC+Tk+mw38U/gt16RR0e74
iE0WcgbI5o8fMEYtVf9vEQZwKfXax7+ZDsBrA2WJ1g5/n63oYF8HwWRv0IoBHU4R
u+ZGag9GSuz1GfFxnlr3oy3ggj3nX1X6zC/cN7hOL9DrMw3+BHgeyFbTHq8px1ty
N3YqLKZlQ8dn+cNOzlJDjoYFR9CZgN0DUKvXibBxyQHoWhMQUcipcx6xVUDeMcyG
J8b7SREOAZ3X6bajz+DNBc/bgeWSwVxxcyHJaAUk0pj4bcx0yQEN8onHYPBSDANr
egxsWYYOaKS4rTigKMPhUACZI+y+3jBrQ1kOE2gW4jRm0U3nukxPHlhDMgm03fJ3
7Ld80AjTVBdeBdtawCMBipXox1ln+qB6uF1KFs9it0gw/pqAodMHb4sMJi9bn4is
zkza6PR5WAZW105GxgcjLPh9wyT04+XuApw2hOn+m409lJ25f53TD87Gs+EcGgTG
DBN2F1WLhhEHvAQv/J8pAbecwf6V7CnnrsbquttGEf0Ow3HuEQNYCHH8+md6uN4G
YdQBUQuba7Y/D67mHPs4DR+DE7r/gBWGHE6DIU3vQW6OCVWqsZgd6C2uxJcFT/ES
r8MdwGzgnkQjeX8G5EQjbjJ2Wm3e1hWBwwpMuoszfA0e3f6IVn9KCc/DpZB8zPK7
JWCLaNJD3SdzraRx+o4XWyxPkh9eTCEo2re+tiwN4XYwf+ivg0Bb/qPL2I0vgxnu
Wg6aAQEe6rUZTTMGgRahzqJNGnRjnrXQkCzxEptH0COr96OAV8MqJCi5vWkvX66D
2B+U5OVMWWg8b8DdFzcZRuCrvZV3v0hTgifBEAOkSso5+bKxoKSgGn7rMtOJ6uxX
U8hiUogX92dOTxAVah/6K2A4pcJRM+oA4jDeIBPJivzZ1nSEWZzCzvmyp41FoibO
0Tz0RItS1IqJNPz4oPkWHc2gmBpRexQhV4SpXxNpzUrHLUydDNMAsWEXqMky4vb2
SAkUIH1e15DCtCzgLGyeERn4rlaj9j+++WjLtai6inAXhcg8AhMek/gFmnScZ+n0
zGe9xxHZN705otCA7oEirGIxRUvF1Mw4X092tfE3KGG1wCEwTLn2U9XKZIoivLTG
TkjYhWLMOx4q6yITA/svknifIVMLP+Rr6DpHTrvSRp6g+NiuzssFacYmUifjgtVE
yI578JGLx3I7+L+Zn1vvTtwUgkGEQvLuElc9F/uOLRSFO0vAqjafG9Edp87/mApj
0fxnHUFRhLSzZy5i0oqG/kOauW7etqm6zP8blcoFh772AIdW+/1qZ1MeI//c9ckZ
NHokB0D4TKy4UvppbqcDua+ar44sOkBuzRLOgqoCdZSRue6L7XUeTsykW62P2Xlm
/oP4Xq3Hqg4q+GwQUDpAbK0oudKH5AuyWWtlVGQ2Peu+rCkM6tPrnBYm28SrAuD6
lACK4NZ0+n0sE5qdWRKPuPT0BoLbp+4lxeGtgEbq5Vw3ixBxaMukyN3FF4Ja3TDd
qwEgpK1vSQc5VrJrC+aW8Q6lpiuyQ+fAN4PkQIdpFL/ucWSjiIs/rOzqe9AI8JH/
oGooXrll8PzrvuzoiNPpiCGZSmxxIl+esyXBnP8npKMLVRMaY1l3joyZwyt6lJyH
mTJItpIhzZZ57T2S2kHoOeqZfqx2T44Oq66fzUuv04Cnu9H2hQSc6vyyxP/2DDyd
1WFajkXkNycSdyhS/oqgoLA3F4hDlYXY/eGDYr777P0E6IovjdvonpeFnKzrpygq
DE0Fq4EVEEBrUtwjGoVXAgQPsBVDAGD5+YYoRNjpnUYSH0OZOSFsC90+/xJsxEp3
sTxprRNqVJqzkmKrbUVCQI6PK9EnZdXq3+1XQYRy1gYrDkToUVmB2gfXA/j0e3Go
hLUHBXMc1K6J0nCE3BuBqYjDh3ZyBWAO+hRjs7JdrOKyneoC6D2fwdbX7sUef6ru
1iXwG3m0AxV2HS2gsk3AczTaq7QZJ5OFJrGXzw6SUizbOufc3cttSyJIo1uJeBJ/
hrwXPfOJE94SQilTWbJv4m/Y2hESCBr5VLxuREvM9kAV55WouNFHI9K6kcr5wsDs
QxmQgQukBh5nhNgAh5oMdr1KH5gbCD1+bDmdbwiiLZGofu6/W0IvPGzKDjF2HmXe
odUpnZI5nBbXNr3FDrEs1o/oKxbONo3hmJEi0LhP8oQaOq6lEXLtgKKYv1vv2o3c
z2OUnlzNw8JiMEUJrq4SB40V3yA43+IMs5ywwhTc5popA4X+F+zmEbnbDmB1A+PL
HwVqPCcdHd61trC89L7Eob4bKZhst/iBClgIMs6g/wX31gXqOejn/SUNKVMA4cP8
mdzq3ajRJQn/yMPxYRH7eJxRq2IhHhwftuMOLY73g1gvjgvBTVEsQItRfu+NefBt
KfyzSuLFE3R6s2QsyHWAhlx3H2EZrFhGE2mj+zYG24HCQvujkpzb5abMik7XmGGG
GTScWtgoP119tzSxbWaQqYobHWrqkmqijzSZunReoEdfhk78CCwmYnb4PHJSI9h8
qjyUYpOxYiFVTWqxqvSNZE5u/QZCfd8+jM+1AhQaNwPPWsEXqhPEznycTF4H9HJh
dbHg4ySk6FV5qjVK2oFjnrhXjOZdleYehI30MHrHNIHFsfXhmrrk4wyBCEVOxNos
BxV/dF4Zu2nkSDukDBT1WXckdfuYYdDrUffdHrZNIg/BcUdKzUFqDXftQSedOJIR
0JH7TBoA5DSlwc8pM/4XeD8LB9oXiQbF76XQQ9yV81tBUsD5TmCyJDQiUcavUUHD
n5x1wezeFvqa6NV1gScJn8zQVRWOYNBf/XNM8KP02FlKFD17WhmuEnYkQLO2iL9L
w7CH3LtDT5IEQe+Xo3UAqZRXz/H2uCCk7v9j56CluogrEKijRkerXGsRSncnHfW6
QN7/qJMFh0tmNrFw0xqxrS4xR5Fi/9SJyiC/bdWKhfyL2Z8AJa0Aao8N7zVArffJ
Bp9Ok54sulWwRCC8QnnAjN/AJXK+6qAz5cxd4HmKj6vJfm8AaQq4CU8pvVoXy4sL
sZ5L005IxQZH2rjxfc72DXERCfledu4ibPkMyLBCkFip9Wd+iX60OZO9LyFeZfD6
yNfMiL/0aG/EgcqDTQ/wfPUsl1D91LECfdfxkR9vYvEViWWdIV5R/CTLIU7drDKM
jkawDTiPQUyFzxwPCZihZG0cSQZXKvj5wjYDyuM/aqmz/hnuKt5GbqxkrM0GbRxP
E8+YxkqcbBlJbagTw/iGnzR3xO889q9unmOZ3VuL/VwhNiOakr5/w8rChd/4bFv1
4rr/YvtL5vyJfKZLSgIwp3c+6F0Kbk8ibTgono3aDP9YzhES93yUbedlFHWbAvwS
6l+bDCByqK/v/fCglWL3eIW9jtnRc7GgBufw+OeF2R+BQ0i/ea02f47nwQCYG9o9
EySW3lCDf3yx8U3oLpYD+SCmO3dUAfdVXKbhIkDgAXKAZEdz8H2BT48etVKSugL0
YF3ET2On8jH7GqqoiR8umLOTlWXoQXKV9C2+4HVJebUDEdbbUdDo4VcUNfyYGZSR
9pF+BCqa4D2RckBSNkC2CZ9TeX2J+7bs/d1QoFp44ej05qW8B/v9Y9XBJX6VO9Vx
xIEsXwZReoqRQKylgIEQms2yAzkOFNGuSw/NTf6wOxM5O0l5RrZCkUgY7ayAdqhw
9CVn8HfGDHTakqdl9xWHH2JE9bfK4urkkf0eL3TjWYVYbd3ekXRpAwVKS3UE9pXF
A4j+pPhoCJeazACVQ0zwGpC226mxgMPvCwzLwrBpV01FFgzADj78Q3tRSFqAaXMC
7F5LUM43TW+YA5sAXrc7z9YEsOTeumuS8HIZc3pkIq3F/PE+UP3MCH92LhMiaXdi
MUWyy4bFIKw2iHrZ98K+tHKZbRlpz7c1fGB7WLlSwHilhrTJlYmMBmS66WhQiLUA
IAP6opZA/abbUvHZ6LOLvi3vGupg85cRfKiDZC6oNuBnTz7K15bS/+y+zfKzI/bP
+cITuR03ylTNcBYpDB3DjPsuIj9N+qqGk8Yf94f1JknwvdQQhwH/7b4tLQT26PO+
mesxQ6TFcdxCN+bFhnW76mt0Co1ZtSUcZHTteZkVuohFhJeFv3nXmE4uqfDXPd/C
fae0iDOmX1qiafw/Umu7wEHqikz72kRqXRbGbD4VxfkILXqFK9/I/gVqNPnAi8oO
n9xCLq3nt/ZG+fROKPTfEX5TVRjFpzcIRJrtgY+7/zUbd9xOhpoKGHe5Wsfm8urX
jrDcB/nBE75rFane3bSrtfxCeiGAFnFT1j8SjZ1XLoIn1s3G76DgTU/kvKaT+SZ7
G1TJ0w2WwwH+dhWKTUso2dXsDgj2fVvRBy2UgR0uLLj3VZgH6mkKWiheICwYArDm
/Miual7If1u2+dK2gaQafUvWGwYbd0UjKPac5vCHYulS4Up/yrOYNN/UE1gMic6y
rmIKNO1yiOncO8WP8b4NfMi225+G5DRVurQqoLBAmXdGB1XIPqwpMTTOgeVmPXQb
xZIQeNUBOoXxaOcgmtvLU5uNVXaRZOWPWWCgruIngU3VA1SwoFJdMq01E1CM28SO
WgJr/5j91zhnHd/o0vvYDrXAeZSb3TzPYNOrRvyj5hlyNqz3Vy1Seiz9thBekiX1
20KiMfMyMI4qtuxemTZdMU7YT6YgQPYn7kJfTco/XlRdXH9L6w8+/qPWbkN8ugr3
t10Tjbc6CNKf1+xrU/9gIOdTXLTlagp5C3AwjnSmQl/EX8CredYz488uhlTSZ9sM
YRYTzBCHrnwKEwnAU18MfqFA146sMCTv62VLnuePbSJigVANlnCCIGzhIDhaYLx0
+G+Qi/1TKj2L9doFmYCaqSt7NTo9id2TC6J62uGRPn44czr1cSwe/CX5s7AalA77
huPsK6MNb/xfB9z7v/EYpQWW7dXGo2+6yenDp6Nel6zplA1TPezZqfUcBBWUNrvf
AkVfmUnwqxzVzdVH9racOqzBKODYW6hNTLu7IlEtVkQsuKstl3axR59G3bWlWQ6M
0EyXng/NgIrUMWLZgsayZ6FQGbSLgL0R6IwJbLP2tDMhFsVL3UksiOSqTK5ydpXX
A7UYuYQVAZelev3EeVSfL5CXNoiUBEcuF3Qri804bfAmgS6dSX5WTeDW7dKPRpXV
d10YkLEPO+u37HT54EbphwaKPt1gRKtuYs7XYSIZQwNnwjLF/8HvONu+9M+1rDmb
pLu6IOpHcv7SKvffCgoc7VF0TJrqcPQwwIiTYjUjLQv9Ogar7eSsKsPtuxcXqex/
U/70cmLFwj3h/RMOQHjVCGpbQi86EKzoJmLvLV1OgrsgsQd+lVLrhr5L0cB7Lmi5
Ngl3InP1h4q6cLzVqMVB3rwBxm+HGPGTuYrUKMX2Qu/Dih9+/zEW7DJRr/Iotmig
GwF9om7VK1EIvcd6ZFY/9QHehS1z2StvsXlEB6u7LXwoaqdOYITqp51vNVy/hlUi
y33R2gjCsbdxVYXuYwxdTdGiGX/k/vXwyahlp9JHt8bIOBHU8kRMzCR3xlrlj+/2
P+GVnjoAEOyCcTg8uFW+TMywvrBaZAOjoDdmNQ3f33Olqr4fZhTaPw7p7cSFlrLc
24V5sy/cADFVpfJ+mHAm76Du5KVVkAyM3i/SzNGc+frDhscf35DJACKYrnvra87K
He6DwRls96MIRknqCVfrVGBGcq1tg2qyFQOyUyYOewE6okbwnEpmLtGBHYurgUbv
BHyevwCvIhuif6tB0lMBmDtLDL6jo2DKN7SVlek3ZOrTi913fTOeDC4KRdHAMq5b
YQbUi7n2I+gTJA++VP0n2CInADXOS1I6UCzvcI67P82VEwWCiuqPEtGyLB5mOV7f
KnHGlDVml88bxzV357V1moJe/DvDaCgRpAWXsOIqt19OdjUCSEHnJuDaSU3aILtV
VjuwXAS8xYIzy46gA5L2xKjhlJ0Kr1jt0Q6SbzKiPGaTzD2GDaSpOIUeDjp9kAaa
ZDusYJoKO0/rVIVeL+JuEm4FrtLjK2vFVPmHhOXHU0rNnTDH0LC4RAgSingmQjW1
ROix1jXp5DPw7IwzR65jUOP8thkEA6yGKRKhlWIW/+I0uVl7fUaj9gqGHNwSYhEC
F7OeBiwF2fs4onNJbiJoCczwRwnDeTS2R3PSUMk2zCDr/cEWMkqNxwMNFsG7voEv
QRT3FsZuksvZyWPsqDf8uBe6C3pK8YW2QH8wV+SAnttG37xqpuK/5i0VbDpb+aeY
JnnToTEywYP+IeIYJCC6E7Dih4ecg+dvIksbaYyfbEJUHmQ7mHepOCRFzQsBxgfW
EicRMJP2XjlaN63pykf6CluuhmKfA8qgE6hb4H4GqXs/XB/qHld+WUEb2DlrQWK6
XA4+GZuFhcsZcfCRyiPwNNZWJPervrgoqOGXDM+KMab2OLZ5oW8MhOX8QZveP6rS
hbVDXIks+oRvY+CrZqtpsyAjFYYQluynJF5MdPIpUN9rOpEYEIvFNEYrhta0IiTN
IOz+N2cvWWlX/45p+0lXzFy5TpaLy9demT6Jbsj1Y38meE5uE/k399oxXyZv7nYh
w2BB96W+/N/BZLYAY6yyuZgtS5fA26boNHmfL9l3jWzN6dpohQXG1N0UV065UGK0
qthni3x58AFTA+ywNqbkzUeAFAZYTNGj1L3NfzKwKPTUZ6rDJ7jEhi9SoBQSmrwD
uWyvy3YtGiHbyyh1v0+0EPNylFHbceTTAZXOmO2d3kaxWbSs9Qiu7c9K/Eeud0F0
B6oWqsXplrOCpYfb/kVJzj9QNliAujVNJLNij0CJBQtBemN0nmIQMglu+/wr7bb4
nzTfW3OCKwbdiUSAuMcN2s+wUsNwx5lIcNusKTsZwqikb+ro0bO052l98SOYWqcc
PI3lrnORR+gWrk1exLEViPgXeAUIf6MTkZuoO4N5ZgSaiVS1qUR8tRHe7i5UkPRi
a5GGSBW5EqKqgXVW4VI9lGQLvzDIbpSS0w+lyPN6RT/hqzpYIU5xvUTKXyyE/+f7
05luAo0HsWFT+b1ckJxNEKapZQjnihpogs6dILWFBtbf2Y27a8xr8/FWrrOTO+Mi
5rQFa+1pC/b0dFJUEfzuBMea1ODi3+Y9oSC0067JZ7BCzsm5W6G3jHvMzwK/SXFP
NAodhJh0pxvBCZT/f6JmfloHZK8jZCxzN2DRA23IENVLw2FxoF4CkyUqvlM/L+N+
i8QF57eamgAdLRGc/1u+B4j3CcLNtlLRqPyj1K5iR++o51wdI2ClkfmyhuYZo6fH
CEEARIJmX0oS7l/YtUBBB+dGexPoIBkxZNSILlMghbYotw/mDBT69BIKWDMqrDXs
AM+g+MxR6O3G5C8+kgp1s0gxb4aCV6yba1u9ZT/iVdp2nndEun/3yQp9MbMqlVlv
BpW7QgeKu7Xj5fi/buKp0yupvVusZaIIcNtoEMjfcE9qw8q2BXFpPPA/J4RPKOU7
DWFZCoDXJXVlZZxmTs3cMz5N6UeSIFv2B/IEWbWpIjyH4Txnw5l3nk22YmyoIP9R
VqWzc4We0JOztbOfrKg/6VEa6tvzOvEfIPMMejYI6c1SxSqpmYS2uzYNN0cmDXQX
RWrx7y4xa6HdfgXuSlP4I0Jx33M86/H4RXGgryYDmcCKdWC6nVOm19+PLiQnRDt7
oDRFqs3cSbb31EAszbpmTHe55T4/zLKS+gB/HiSzL+DTdSlhZFMI6UY23Bdg7p7f
mRfYQllsbUUGdvGphUyZscUkG8Du5gsDh6FW8c6xRWhVmZfuSZ1ITcKEw02smPWZ
9uOLqtWXOuwLvKc+Xy/qTYBUGSnk6mFL6Grjg9WWASvIKUlMZmuymb6HOUIq+8WF
vGmz4WRi7duME4VpgTPn1LVN6uF9SIGqiVcEEHYUJZ+64S6E+glIa9Q5f6xmsp01
a0hcaeLwuCbGj0IPyYEdlb7vd17j8wD2xZTqWVSSj4p/+NBDBC7mJKuhvGo3zNGC
5DTR0rCbmLSCdNnRumUf42Ezky0Qt1nHCvMkfDEE/UT6OzphgpX7OeZ2lJwR/5l2
MRX12YtEnQsei9teMmKdFbvNy6z2Za26RPcLpUQhr+VyuhZEHgsooMdLn/8VrW5k
OBUDGHQgbtd5gotgueAe43owzA9n236nISmxLr68U6Lqo6VTLS8ycaW2mYUMro6E
X52vTqw0+bKacPhNFZEHJ0nN34GU/g05OynvQSHsJVyfn8KY7aJt8Bk8+5omrbpJ
cpUrjkZKHuDuekAfD89UB6HrJg65zdOnBvrG1/UGkY5rxA3lkmN3SjT8oDO0zK9s
/jaky7J6FqGYYx38PjyEY9sKOMtqa7P1s+TtkU19tD3F9LsZq5W4YJq8ic+1T0hh
0kAdFxdZv2AJSOWE0twVDi03BZSCbclBxgfuH3cKptuEmizjUqePcwMBA8RpuysA
bf+CvmdfiT1jcpRdyuloPPmtn5DZhBlTdZ7u6osHaQP/xzmRxgHDHHjhWDLEDmIw
1yXz3UtsvI4JmHvvYcBamLfJsaGM1APwJU/5HxGTSJSEYeTjF2l3jY/i7JCeGiI9
V3GfbyMuvoe12JVvI17KSyTqYOqREKJCpE/yiP76mic1Xc/YQ6HQixJ8jjjrFpNj
naPEYG9U61QuTOPyUPQRAnY6I9ImMxUJYPPKDesneWGhUzcgLq6C8woptqF1UCaC
2r5kmikZqOZ1OXHXHNvUBZ+T4xpucTlmraCcuMyxfDiotf2WEUfS2563R+qM3qBS
NfOJi8V17wKuGvsnHD1fLI/no4ORvI5TE7mP1niEtGi6QTBDd/Uu6jhtLow0SgFb
lj2uXrPdmN8CdsqZDklTvjn2d+mKwb1TnxQ1wcbwmCk7edPOZ4zwwdKt6sTXfAvQ
z0r3Dd61hjcYFI7tztL7Ynos0o10KsDKXu9/HaZhy0TQItpz60EH4BtsJqSKBmBA
pCs3EYxHtGLfL5uWVVcvMW/NVM/bWS0pJWI/l9KRMMrX/HcMD6vMh8xWFHd1fkru
dkSKSRGmt0zoLaGtzqPrgpxaoHQzf4W0nrMHHdkk5mqM18t7ax3WI0ZzJXuGN85a
3/9H1lm1ns86xbSVpiqD3YIkcNw6V177DgoAToNA9tpJ4x5dgIfi+PZxV9KdIXEF
yHusm2IXjdSuctggQRaKqtC/cdVpGntHFMlsHhtYZkOvCTJxyFQLItNHcx5SQNaL
tHpaq6DjP+PUi+vt1OixNOkkCth331+0385/+tktb2JGV1N+Y7EvoF1Iwgrxs2zo
UTr7yfP8ZldEsogl1kPTA6csgr5+EeRF9zCsWn+eQs7jdA41A9P3iEOndmKHG3PX
xABKLcB6uwWyakuwa3iLQTbps44IZaPROCO7OxrQf4kYs8h0ltvoS2OcjvZmepRD
aO6WyHO5Jtzq+RA1/KIlmd+A/vZv/cYU3czTDd+yK2kTTSu+ipajlZH4gHytamUy
E9fUlMT3E5PS1n0nHDyO+gw/3zRqrKbzaRakWHCl4BIb3ZynO/bs6QL5VfOa1EdK
9KiHNLxGff3SMOxCWpcIlCLG1mAu5ZS9vpJxFL0iFT/mW6gXvdgdMd24bAZtau5T
vw64ljKDM3a00zKeXd8CJzhhFka89HRkS8m60OLgWqqm3zZuNhMHEvgFOaxblWKY
+vGPapNuDLwEaWdIG+eRSwVRopiwdze+fRvZePHr4HpcwUoLVJzLAPUdxly6vgLC
C9axwHqNWm6mj8pWl5R16WlBL01HGpRcVuXgcXkzz4gCA/WAeUnfx57d6E90DMvQ
/rgqvhihNbYxx1+2rm0dgQ3Mm3NnPmGTjYlfGoEhy0sOIklswMiYO64/x+Pg3/5c
X39z1aixcHAPbn8ttMJarGztJLhB5qil6R+lhgZSLGPlM+6gVwz8NDCqwuO4tCRe
CugaRwXCX8c+8WP5d70oe6tRH9s76CYgXrH1bCQclRTSuUs3nSHgFuQbeIxNkWYr
Y9phg/hSHKNmkfoVJFTxVpT/8gaIMDvp1mt9zK4j4KAchzw+TjaAPvffE8Cle1ZC
2Ar9cfS3uEF3LU0dPSxTBb6m1kV14RqOY71SgRFov5s305zPIP7kyKAymf05j/TP
iuvstJ4yLGSdbRE1oUHVsgBjF64caU+6AsaDp7CGaLY34yOCrpPSJOZUiqfv4Hvs
OMru4vqvb6efiiSIxcbsWRw+2/CxVOfG366UrCwVW4Cb02Mz61Ae0PoH8b03U6LY
NmaJFE/MfFAOrJFvEcm2MmBgot34L4ZFt4oYRBVIb2JPUVngnxSLlb+bKI7pZGAN
63xGcB9lK94V1i1ighqd9RkmAvfg4hHuQoh7TSKehH82hbmL76VF7a9rNpBKFuvR
0Bt8Y4Mr2qqTb51T/NjQ4YLtpdwMTzGkxZAyR1OEIWc/p0WeUhhSFpl0QnXNzXDz
YZ4y2NHDvjC51bLDCbVnDp60RWP0OUbdV3Srro/mQfuJ1wIWK6A6W7N9Jw0q3iqR
JPlkvKYTv24JHxjOInWuNnmbfmQMhIjN5hB0LYexW40zXcQvrK9zJm9/MI1C1+WC
h5QQyRmlVAvlja/mz96khp/9Qtm29K28qqEsATXtRTP4amXCagICq9E0vlnqC3HO
eY5KUNS7o+vhClZixgLtxgOMZMcd3h7YB1JARN8EY1+asEcAcNotNlOqpNYEY5dp
/CtEStbuDr02IwKsPTVUMja6vpyAVWwhzs8xcrX8BofSF/3YrQtWYP02QJtJ6UXg
Xx1uUSPGYquV1qUmesIis4lM0X9TNjn53IInzctBQNkIYnrb63NqhAlwkpgjwt5H
nIyGbqZSPIs0LlsJAYhwuHCn4bvbsfiYSfcy5DOH1Klz/j2ETUyUIs65K1wY+H7V
wTot9Gmh811JJiAT14YEg8a0KyYCq4Ob0m9+ux1G/qPrGnIokwrgOIOSvKyDS4a5
BH5/EqFqgT3SHBNjIYJM6cknbgN41cfU+cZQO7oO6xonmrdzt9u9/FG1AF9f7HMX
gVjk2cy1Gu2IcYVVTKyCHL+lMce0YRiaJq3rucJYyB39YnsKGs1G42Zfpz4LJwNY
DZCgODSQOTzoYj4bQR9NDQjAVdMhJCVbcScDK6XNmZwSeg2GWshUGd4y/sj1aP3+
oGdzpvPqTy5SXLnqDZgUVqEVlFPLj03Pp8E8YrjnDHpieOj/SDZySbuhHj0CCYpI
TAntr06HZMkSz9iq/B7+UDr8Z8qAuU7O3snTNn3/xrcX/WDmIVc99VGCw3tfmp58
HqCKFhfk4tma9fIaXt8kGROwMPk/ntptgME96AvlWDQW+eOLs7kr4k2/ZWEV5PZH
zUoRNU0H2svrHvaTMxu74EzcYwvjfXDhbMJfO8Wiq02wJI/T7n3jYhDi0eE2ZIL2
0uKCP+Yd1ynbsE0Tuw75YM9tdS2jwRcZUWvZb7jNKPP69d5S+tbSfYh+kTo3JDYk
SPTaCWC0amDr38Tg5/fMJg1nD1bI6OwGnAfEqfFk1aIJ8I4K/U/l1Wegu26Pvi9x
eS2jYZ6yXGZX/2v1pAXJRCroCBXKjao0QGOGpZXiqfIyTkUSmSm98nBpPqSPgH0X
g6Z4yxtpivnQcx4KxHNePhwDLI0PrwRlXRbVnhVLEaZOTi7D1batxiZ0I1Mk3JgP
hZZyqup32fQJ62qFdRyp0Rnn4XMGsCcOTAkZQaDnv3B3B9+/E8913KwUL/OdocAv
nShrQvE5EXMkRo/ozBAwkZuyyVvm3GIx1+5XqaWiRFeX2JGYsGV7JSwAO0lhKeAq
0BDA1J6/xThEiQFfAn/Vgb2qwy+CksfHEebZvE+ig30X/emcH+2IGg7/5FzzirNC
PRXFuKK2A4JiLWvtJ9CwWKc3M/nCu2lNriuIg2HO4J3F4jAzhZv57ocLjNog8vao
PCnaKSzzrWFLSi0wiJrInxRfWfHCjultCwbJlA/NIucAIj4RoXDZeh3SRp5LGfHk
PW6LAxBTCya+ki3IVanxJnsN0W9E42S/0Cut9fbHvyKvpBxv8Mdq3KFulfWa0XAz
mvM7LtnNK/Gwc2sckXhuyKAlHaqJOoncOUdg+8ymKSkoPt8SU7C2cFBuOJT1bm0w
vxdxFtnbGiHaew/Z5A9c+GYVq3G3h7WTPsSL4FktR1l09pxWVW7aBmAs0Rev71R7
VHrLTjrWHOpkaHhsP6Np2WgrjJajIYaJuAyFNFuQkyJJrd/0LFw2VQMN//2RbeM9
ThZgluZmXl3NxUGgz9mAsVtZAiwbw6Qka+m6sOmdGfQs/oEVA5/mQFxZPTMgOLvj
sHj9FoHtQ4Q0C7X/SvUqcHb9iXQgDe0UKzaJeSo+84MHCW7/ywmS2CkZejQHFguk
knn9txQC9vC7FO4tC6PLxZ8YiUPh2eg8DlJsvMuLl0ugxqJzjGCrJZTHfchtinzo
W9iusqAUEwCUo92bCUM+W2kkHdwiXikl9zdNtBScDMj8OmKQAPX7PkZ0hJJaD49W
jomVDpDBWVUvmzJ82yTcs2Vn96zbRyrvnHbTf069kVRW87QwzbckbjPv8yKbZYKC
A10TNbL4CZfh7NaKvDyK0KvjY0nViIQ5rhoJhCuOKbBbwdiRKSjZeAuzSuLrRQPB
mRuvagES2qeEb5/luA4NrfEJAajf1RvSr86ZzQTI0JJIMXWjVB8PjlWpPULJtnTy
5+sGAvdwtDPJoCX6Cf0zTxsJ8aV4w0bKhOtLAKaoCr355Y5OMU76h3pTdjy9Y4dP
LSD+mDMgwyBv4nQ9cJCBa9n82lGGRgEtv2yDYusDM5uIjIQvqodxKWStSigj6PTB
zhjR9H3mtAxyMYcqtvisJXrQym/a1dtcbhy4B/ZDz6Z6RT22asFwnVmS5UEzvUtD
/bcQTfDdTEsugknfyNGGq+dYSbQQ6/f9rI5ZIrKqalMN30+v17d9eVWXt4PT3lXd
HupOuDpu9Gb0TnbZYbYz5ZPayzeRCa/GeMzzJ6S4gSdCFLHLeJlaaN6dprnpChY/
Gkz5aHoFtmYeJZu4KSG4GMdG3PfjeXhMapyAKKDeV0jYwM+/fjSKATlC1Q5ki8CH
louxvU7siRpAJXM9O8Y+Evxg0n1Ba1Pb17fkLcnXIbIs2Smn5F8jlZu9Dfg3z3hp
jP8yoeXD41UXyIvdRiqDwPTHMNb+hp5ywIICUXuypIpDR2T0mzEXvd4ilb07ZGzb
45A/8ZKM+S1uZ2YaeY+O+SRVSl57o4Ym4o7buOOcAGPVgLIlqH9/sTZ35vXghfmj
qsfSBaFIvzzm3MBBSR7RH5939GGB/B4TdfWZa9tbO0HFkGzUjKwiBmEoI0wf064o
m0DLrPwTJmKGZe9LT8L2Fkd9vy9LZfuWTkRBleNN9fM6aTBrU75d0/P9sEZQ7pQd
J3QHDiWwsx4nOM2IWDToizh5GNhMzi3cuI0bpYNJVwxFwnK3DWd+UIBCYJSHeKJz
TWyo2Bg+2sI8owKDIQW+vVRAY74CSEa/kGVu2IP4uccx47hqYhPAE8gKxQ4UmedM
as/3L5nJnRzUnhIzpPhex5gPx0BwvJdiNjpc3GtmpmhfpPZOpxnC9oEpcKgGJKpC
qf62lhposr0FCKIyqBeUVDwr+6pIJvcJD7ZTQYnwH5pcy2sLTY+g2rlz9FeJ5h6Q
hcyw/DsWeIAV7koYVjekQXVMW/qFXyMJ1JThL5L3bs26cYypjCgSNpZObZf7OgUq
Wa47TS1az436goy8N6U7ap6V49WpOwbWnXdDy4VDKaK2zrbTegJ0RfrKW1PT9zuc
CBc1u4yMbeb45RzkL8mVBeZ+gwAIGkMhpkKkdwPuNPVVoSIkBDtpoZ3qS1jksW8/
O6uAr5OEavdn3nA6CVIaBxa4h53waamINXzWUrltnzkEqHKBaARu8fEf3c112h2j
X513Rq67iT1ecwgwTaqZxEJEHY5XNGkz4A+FE0Ux0MCRxeMCfFoRhCWTbEdverBq
a7+WDL1lrwkBJHAbuQzNlAjVvfLTkAiW8OUHWupxkix5OIJakBFIuLRy1Lmq6FKU
YuxA9zeFygbp58hsNZOsWEJxf5eIaALjjnhubSnZo0MGoSooGFC7Q4cLS605lFtD
7ENhLgyc+vMiFR3sZTeiPns7SUjVvaGZEUl1PQLXp30Z4O47Z1mpNytlDYkOj+G2
tDX98IEeDE3IpHzRPS+YgjneaO0Qod93svGU1pI93jeoVHItn3perspPNlbXPDWS
eZO+7AIfGjRuj3clVpnqNmJSn8RssTXMptezUiTFUPePXGudz73AHVSAqsTWqdSl
xosc0h6RHNSwGoWoS1ZKknn+SbZqtm1BKBUZE1ooVsmo2eenq+9ilM3TNP16kyGm
m1HEIH+E4jnz0ze1St9p9t5aYW/7Fzsnn0UdkWbQN/A7AIv7qdYwok3lUY+pUMpv
VSOSLn4FHpH0wm+CAHbPl2TIa6uFd1BmUPVgHmcX9A5kExnmQiQUZ+wJVmZiN5gk
6Auasc2HtrT3UdOsKDkuZ+7rGvgTDg1mx1NKYl4+wSPrA/dIbym9aEqQpQcRlnQr
deKLk/1hq5bpRg5Zpos5IIPCAx1mh/ss19AWipcMPfKRhKnO6cU0/cXGjMAlgUQL
6RnzuMkFwPUJwNgJe+aBuqDrPSGzTUCqV7JmVAcoQeMaLGcSNOO6ZU3R+xExgsPd
gVTd4chG7PHcyydEHqiQ/6CCiLPdcGQcraPhbDqx537ArOmSrz00xMVRT5dAuHBh
QwHGRHs7zeebKi8tN4QPmE8UrmzJrmthZt9apxrUAsdNoim+MEZ67plHzC5plhYN
Qf4YjcT88xKOjU8cwkHBHBT7erVU5woUZ+DgvEPl4oDmb0MSWI50TPHPsbAnDEtF
0AzBcBBPbMP1MMGINTXhki77Bu5zy8cEZTeiPi1FMN6DO7G7ACEqY7CNfue7pPAu
Pu4ZNFb3GWL4W9gPInkaN9FnhH2MlOH34rvjjKNMe/LowzvW7NcDDWkkZZtH43AU
euCuL1BtX0PwcuOdmv2frSCQuAZZccTEbLySdxbpJebepVXH49V6TeB7OEID/KWA
GUk1PIu0r4NiH3WGjvmMtfb4NavEs8SDgA+X6axvo0RrGtQzM+kX1OW68sOpVJ0T
1vhqxh2ugp4yPSlEvR3qaHt2lbHtEAw6f1xBjnrdP+FdAzc2XYaJ37NTLNkCCqUd
w1coorxJ/pn7RyuuxEhuLBmvTZvCshsePqFRzCFPBiHg3y8I4g40ECb1jLEgw+qB
aoYQ3y+9KYzsuphrokX6Hn89QvTyTD+EaCSKqSyZ4dCojHwa6wM5UgN71TxG9Pqj
Osu2DmoQjlLNkalrvPStTwcE5ox3cds1+mAbv2LiPDAqlKc9qLWEM7FHY5DjgZLl
nAfa0R1n/qrpAQ6nyiYxiOugNJtv3fOB0r+vjihmXifTa9Pi9MLP6DVZyb63AupJ
zhv3e6GEfHXowVAcd9VuEEtAG63+EOCgG5antUwDYTZlvx79QqP0NmJGeqWThLSj
eUF5Z5NWdzCKgZwWyBDVZOtAs+aDNKRJDOE+7DuUfXhVMrvP9xUVeDRUC9HDhUsl
mZGj9SIklVQb80Uo1s8LkwSG1NXlFwoVfnY3l8XRZ+Fk8/6ceevb+oF7O5zeR6pP
VTZEVXUVFCzMY7C/9yhNv66wfez1XlJU8MLAvmDBTrJIZJ5sXKWrFr+dsYBbUpV6
3wLfI2Vh906+ExUGjbYBm3Wpi6MX02zmoRZeserbMjPqBK4Qtzm9tGTZCTeQUDwO
pTqY9auWO05TXRik8jl1YYvr9IX5zgqVWbwRulyFaCTJ6txIOGsdd2AficrCYg6S
fsXysov29/iPuXLzM5jyqdam1OV7Lw0giwQ2zSugnJiG73nZ+cEV420tYdVMs1Sl
CwCj/JzANFjoW9RZ8ofATzWBKrHwQK2ulBT6/KCkDAG2M6R4WRe6joi2pLkoXg1N
CgB7pkxf6ctKosOiDsUkJyK39p3tzmqdlfcTx/Roddx1Dy5khrrhxysIzzaYLKhc
ANdo1IB1DCkgjRqvpxxJbQEmYQEpROdwaWRRsCJj+1NKT/0ZIrvFg39H1mUO6j+w
W0SXZ9QKDpnQ6T+SJIjsxPaGThnf1lyzRHusD8Zv0ZkNYbCCIsWCmoF4bsBSdgYZ
a4v75oMkeMPXkQPYyCtq+nOACBv3tJKLbHvCfFR7cE+vHYLfPSzpGXCJjDTMRyld
THguypw/diS4mvaWE7jiqTEQ4L1hXL86FHZ8WU88OET8d/OhK6AuY2Yhn/M0LKw6
8wvE4yPce0unWbZMfNegD6PkqlvQDkTsaHlp3069vahd5jVsdMLlpVa8jYAbeWMq
HM1CNU18u1JeOBBtOWczikD0iA2QfDgruHD0VAI980WiQPKnHmF7wLJsVsHXMH42
5lZ9kFPXHtvZkiFt1FoRpv0vZZOHVOBUl/HbkhTWoJ85U9uVmHflhkN/M+hmR3r7
DPrk7IDFHrI+Tp8ipty1pilzDOBScMxKZlFB6RbXgxTCMEG6g6XCA9XvlI8VdYP/
2sti8BOpn1VoRudik7Z9CHwi3dyLiE4YIj8FP7aWEqayhJamKW66Xhy78UODV4Kz
bm+3yKNTJsB0frrPPlextI0TdnI5DUucV2tEVXNFofpNh4Tbkatd70nCTLAQcimr
0z4b9/j5yzJU/RPBw4lAx6Qz2EvMmAgT8749FTO0kwViL/4h1pb/cF3oG2ojpz+X
CWv9AADTRxx+uD0CMu3Owz2W6E4H1xZ8VGQtvNL7CpKjrNDaCncUFIYZZ0oH3QYr
6cu1VziO2T+9cJWn7fENACOHy+3eyytQeqvjtZTyThBsR7jxHQO/As7VDKMY3WqQ
IeulcWte6g9vjZrtk1tUZ86+oy1T2rauTHGC1+dIXOHvB64rEpPwiJgb6Duo28aQ
ZTbcM5+oS9KN4pKEInuKD0zzVq+Y2PayZ1H0ngK02PgSs0r0WUlhIAnDjIwqImQ3
focUSCtZvUnGGAjfUV0zLdWrdOIwc8lrL0Ra6/sMz5xoOBER5Ozvtbc9SN1V8w4k
RC0V91qGDjAT5UEO9Ke7b6DXs6gHiKTg0vWY4P1fgyt8yh3aOUZCr5aytpCXRs33
n/Yt1XDYhyjQx5MjGTIcVM6SmEwjxm/261BuiNSqU6V8k359L+O1Iivq1WHe1pnu
2E1rMBOxMbCZSAneOnsjb3pIIz4jlMRrtdq4hNOZlHbNk6lcodHHwXPuA+eTXoEO
jZK7KsDVWxPkivv86KZS8oSmZ8Uc9bXmdNUvPmbWYT/g7nE+oq4a6rzIWtnSwVgh
x92WKAMweT7af+si9rb67RJTbht2d+vZRY/0ESa0LXEvs12tvkWegXEpmwbpPYkP
dJ3KBOa5PJ/GCsdZHl3cTFpOiPEMGlaA9PhiaWPEifuP1mu/x0/3C4uL+EiWtLjC
BOpX5skCP3qd0j7ejM0FcpSFzG5pp7VjNvtjBbpfsbdcrpyZ3AyTv4fbLFeXQN9k
f7Pb/QbksNzb/El+SFufrNo13Xv1HvOdeijwaqD6gCLSVhdYMohim79YYiazGUok
JES+NibiU9AjzZ3rMmFpsTGkDPqWipZDsAhnK8j9DagGbpB4/i0/UBHGOgAuFpm3
LTitdID+LluzAkpNCnqHufmu1B8VLdJovCDo53ZMfCjfoQnliQ0d7Ge4L1br+VMz
ysoK9xkj8VhyPNF7corZi6Za3rmmdL0x1p4xi4U8mObaD1m+TwwKjjvuGzWlZVrU
ZIQC+wLJ669KBU4OebPqJj7x8r/5fsuSvExFgOiOmTjHWufMTwTexovXGEt30gvI
cZnJaaNvWgwMcnbjXGOUTBXJ6cY6IB8CkL5H0UP3ObmjYxeAFvbMnVhCGb0/Q7WC
UQ1NB5iysMB+25H/wYFv6lYQj4/AkRJbtI3b5XKti/Nr9GOCNA71/t8KNVT9U1WS
0bJUeW5/+YQslAzXIezS8Cflq7r7ByIv8iN430/VT1b4MrHUHshCAu/buQqJCyso
YN4+KoPcvnCRjHQVlOiLOtWl1QVJL8lZyVnyF7169J7+O+BxUCwG7yF3z9WXIkwe
vihgsBAy5BNED0v31A+9HpnOvTY/GpESgnNs7ccbD1NCTm0dBzGN3iVLk/OC3qKc
OX1HZarhilbX69YXyquMHSzeJenYONJIqZaAKXWuOgaLU5yLCXg7+DSSsT1a/yYt
EcnyDcMrLZUj1fTa5WyEkATO8fN7nlmSdM0proxLtiza+3thust6TWCgC+CvzJxE
+NxmYpwZO2RrqwVYfr6F8HVSzdi51nPF2smQpFmaj6MnGXJjmIy2MQiTVJNvOQ3X
ldZ9ddyL/+zVeGl9XB4giyAMkRtwpAF/d7dGWgB+NcRfmfQfqeeAMi2tpDMmcHB+
Sww75aoJode+Qpr4/Ma2w1Dsv4C3cMCPx2wALdg2RRAAMb/ufsY4e0Rvt5Q32ayq
YrYM8vdQAzEk6c6kHzr4KimGIVHP4/H3s7E2A3EvwWbEYvwzkR1PthY/JGqXg6hZ
dUp3QpDLeSPloawgDBm7SOSQVN5s0tXsdjALmtk4jWaoI8sLWa1/OKBCXQ7iRpZL
IIi5A+y3ZJwBT0xodcPVct2e+POPiptUpZEosN/rFurCttKK3Zb6auUJjROOF64S
Ii3XlcrGt5vaXc/+87FYobScIdu0uKjMXK4z5zAm1xYoDLnEXzSmhC1dwtTqTPzv
YuMQLvX9v9aguv7M2ulGiodw3JrbZ9NUHl8mFyALwXj/Epa/U8KQGuwzlc++z5dp
0IWZL/P9Hz9PEk0y89YDRUgW0OCZvnI+ebvVdJV5UAiu4LKcMQJAoSI8kM9OOg7t
O/Q3xjknApRee5Km5KAwknvwckGQMVhQTkfPelnGigxegbeZXVk1BzQoEWWnOU+X
Y4+1aLYVkEaKOG0J2L96lZK72rCOC9SkRxK5HnaJ5BPCSzVyN7Sh9chlwtpDPLKm
KN3BubG5VlK9WNR5hq2T8y/GXe9gD39rwlVM/TkCAbr6pSlRdylfbpPiHvdWoDxJ
CuqG+AEbsmHcaTOyktxLSlp9cWOh+FczIyCilCnHVwIv8tzlm4Rbd+Vm/XBy8IY8
Nn9yFpsXM5nngMETzvo3wLQct5NjpTiBKXjlvSJYsabu9ReHnhBFLKsqFaBli4At
PdnbYSMTm6icE8RPUFTHAlc8FQaD3IoT5bpMGipUZ888ycOmajQvikuHS/TirAbI
ar3U7sfeMwKtxRdbfMvoBUtt81D3qMhUX4xE7tM4eZntaDMnOqjUsWK5lcbtQwNq
iWUygcuIXnWhHJeRQAiEAssn2ssuTc7KSTJbtB9jETiif05wmtVltgZ/HxPknwDO
ec1eXPkuNlJZqU3hfJgvB1AoI2tvusKzFWBfhCyIirBJ2ariyPjQqGY4KtGRtdQ+
a1x0o+tdQKXXEg3Ttp9pY+TJx2FgQZCQAo/uWvkR+19Skvpts14x+4uTnUXESxeP
K52s4dOKA9n5DnfXbRYKy656W5zSp6+JphIBu5rYKATugwsoGu0RNIqMsEGC6eGS
/Sd327r3SfAI3COYmpCXY9qBD3u9QxlQ1Cc6Of46gGb0F0uanLbP1IPbOHQEOgSz
RtsScntCWoBXqahqkB+Wh1UF/TgY9HPTB2QEqFhw0kdXF5BiwJos9XOcFF0kdFVs
dnuYqaETTm5uK1fx097DB1rdx96zmLxOZJGSFmhR8eAcLmIeygWDY1TfGLyb3KT6
6vq+ZWPqkdmbGn7fHO8FHfC4ec48ZpZwJH1SBezjnOMngYyBf53a0Oos3W8DeGUo
6DyAqfm16Gd4tVt0q2eU99vLri9+Ht5RwtWKek8uXK9piPTPFB+0rJ2xwvXnS7Uf
m+S/bEt09A7sKzCL1VL/7UO6kAo3SYi0yUuRdhlNsYlmEZgh9ZItnbc5Oj5Nw9cU
Cz5oLTeiD0BXP7Uy/pn4Bki9Gyl5j0ZyacVQd8Usc8ythmni3JXQ3g2QY6qWi8ot
/7zmTYWn9WRV+1a1PzT6hyVOfMb5+B0h6FhS9xpAA+v57kVRQvJt0gAN4SyIxTyH
Zi0YNTkelnICpAggg/KcnZXaqGXohOUF0uR+QtiJDrjoj0F4p5sNIjn40VHB0XLo
O3scm2N5Mgjy5VQcEfHHSPzroJZEQBR5FmiuefsU7FRCBlSI5qC3oSPu5cIxdrz9
Wws0sIl5wxI/LtHjawX6SJzF3EDvaVsXcpKvmtQSpnGoUBDtIkV6KHbmj8F0QMoo
+HP396o+8aCQQp9ZgEB0BKQYdNE4eqxdIm4zzRkoggqgTbjmYtJTpgBvI633DSPb
+85it/fSvlf3cH/j5gbEUkDN86n+9ZnLfUp8ALvpDeTIZ3QksZohOQnHgs20fSLJ
4p60xOeDhjYe1p+CfMDaOCzVMwevIhQdwLj5SZ4nnUMUw6cfqQ5qm9h2zfZ1Y2bo
pePoz1js1vSz8tes84YCoJ5rVQqVfbF0v81EDJhzP8D4eBtx4PMFO0Y3+cCA0lOl
ipRweA86zIZhU6vJPePumI1T35kncVfbxtclOeah8OCZmWdFCjjEj+Fz5Vnivxm3
Qiv+V2HJWRaVA9i5FZX07yKMUTbkl2Ii+YH3jrcZtZNWAlb/uL7Ef761FvyF53n4
pw2zW9j7Fv9qgpj95pgbHuTla1qPuCto8NKb7SfbWncBYCWeEVUth0IHHT+Pb6d9
XJRZr+pf1C/b09YffXVSw//iBfTC0xZXqDL7f3s1fFSqWTb9HmbNMC3E+X2FUPUx
Rv7bYBIBFZoem3ZE8oj4yVos3svLCV9nZLlYCX1Q3Q8PlZtmwK+Ov18k6has1iGo
MlTlNz6NFW6nkiFNTpHhJz1q5RwsevkFtxL+yMMbp6wuJTt0vN4cqcFsY52I7FiV
YbeKo1k9rU1Hkf+dyBal0yLaMW9ohCntbZuAiCavt1I9FjdyywWYQ4H2FSCZxF5U
lMnMhrjcek5gi1LR/FpXdkp0v34L3iBXHKtNlf0cSLtkQw7Ws0zC2Elq18kN7qKv
plKXq5t7wmynbjy9dzSERdw0EwSafrq6NulOiMyAflnY6HsccLK7gdv6TbU1ofAp
JFMtOYPbuDUdj05bYu68962vcZrghmkCADtI5kz/p1UnmcoW+sv9Cptuu3CNmr5m
KzhxDjEe6uA6KPBL9Dgdvyl+WqqcWAJT2qUqzDC2qk3qWhr0rKPyDYmirkK4WLgP
xnI+la5mYKp8wxrh/pu47p4yyVy+4cRkSzdmJwmxbuXEwOBLDvgtKg1cukX1MLS9
H0qNcatdyYSfEyy+wlxkj8NXbWvl7wxNMDSCOBQpr0nMifOdYtwlUpDOnL8XVGN4
qGQFwVZmT2ZV8KIDDRnuHgvK6bhCcUUm/nU8kWrNo2Rba6HY/uthbRjC+KvN4h4b
Z3rdX0ILukcl3PwjqurqLYDjQB5t+ogLVu/MQYjy0d9VzpQG09lNRoljADBrVgej
37q/79aBaEaXwLOSuibAwP1YIpEJbe/rIvjQO7WPgh+8A+f9vKjArGJNcxM5bqSj
Zc7W2YJQlKpGR9Hj6I7bD4nlLv3wdd1eo9md/mjX2kTu36K2aMTOIzS3RGjQdgj3
kDgm1MMVTg86rv3Wj35yiR4STWpgzScWzlWNgXWCzOjN7xqJ461s4yuO69lQK7Y1
hwQsJbJpbdkrsDQyxctgor6lDRggMphGwQKsK4vWefuLrZr4dpS/TGOCG8klYtWX
E0TzHFkLmNQ0rICUQ2zgvsQDdbeCgqYoTen92FQDuDZhiSVUoow3DPxP0f9k+3J4
B0W86QVWkZXjT4zoSWrVtpB+nnoxewfk722Tk52Luo7/AGcmm3ICbtzlpjJNMyzH
ytPP/tsQfpKEOhTCkHxZIFDVfdB1168gMWJdco3vWVu90ZChkLRhQdNh6dY36Jai
5XiWDyNfdVZye9MxTCFFYJPMRZ70fdxzYweWvLcL0/p6J01jiHwgpepXmoSONNV0
YnWBYtve6M+W8Va2r2iTu0Ma7s/Ndyq+X20ASSe0w2u/23IJGoU+OwJsLvNGgYY6
2S4GPpm7i5O3LLcFQsYz7OZyZd89F3P/IsBBcI9dgSb87h2Yz5LJypkENlJdpuxR
H/e9SgAE7NQIvYmp+J/t7CM8rm+SxHHqSY1pTW98GoyEvh5QjzPqFj5aVzaagZQS
kXvOXlsBCC97DtvMpmlPb+Y9Jj3cNP8LaTLwCSUl17h432H6z3S8/Q+VMcsW8uct
OREXO1HCaty+5g/HV3rRguMLVn236W+nEUgtSGcYmuH9VTKKi7+2EyOYn8HuBDeT
kSoOCN/7w+k2vRuAvO6sxCONJ9pOoEnNQ9TjLZDosTtMLneLkbndtjQHgtgkMzyd
AIOoNA1G8XPNlKaD5IXJGyHhBq1JqKMY/GgDFn8aADcFM/+K5imQB5aV/SOjIlrS
DaUP9EMbxjclOi3R96WWCeF+cvLMxCODonU+wdxoMlXYb3DJ7o1+pPblVhT+lHOA
av1RjhZyodLI4Akr8kmOxNVfEXvmkAVxH0zBalweV/aKDNs5WC7/K1YuCXQJlE/e
Q3tinrYJ9y/rDg0OgOYC9Sl/DO2KN5CFF+0R8b/hkY2m04mXQypfJFyV779qNYJC
JcVMIAKxYMV2QLBaywNwo9DOxvYAJr1hFmR2Lv8o7ttEr2WoFff8um8fPdvJV8Hu
SnR5Un0I1ruYYxANvWdq9chS1XuuhcFik5PjVV5Pyz4HzhgZ7dW9lW/xVlqQYAKA
tjnbaqd7EPcFvsImUV7faw0WGbgaXWYloMWN0OjES1Zen7iHbgbGAKqOKaAWm6ud
H225CfWInxl3m214hEFSPSRHgRBTngmMLdA0hjFUuu5g839lgjAWAUOijSdPPIGZ
B9OohukYwhAg0vX4Eld0RognnpTrSiJhSeYvz6U7x4dMt24PBAHP81APeFcVhFEg
lAQoJTkYS1x+/o0+/T1ff2oD5HQ5/s31GqZCPfEbMOBQUTDGMf9qXy9gxUZzh/d7
rP4CxPmyCiVjc6cAxjiAU5o/UpYAgUp+b6prHuGTjaqlmJcZTvyR9QAMoQ9MdNid
XptAj12tu33Yi9MyFI9sp0MJ3zWkEFHSJs+j09qXlR/G87cEwChG2ecf3WsUqEWX
ACJagyApl9s7lV+cCVmlYo4M4cTGKe+klHkz5DPPtmYPbB8SQPUrlG/1ZFbX1HEi
FeEuoShehUehHvdID165RyZCUsuXGERCjBCSIkHA9I/JcnDIt8eINtUCgOlyRSSP
sGLloiCN5lq/lgdzIyrtsNe/AZBqY674ghVdLKj1JT0ZpBzzvzNFX4mrJwdxIohN
V7aquumFhISM+x30Htq/ZLKxiqDqfO7FZvN8iEIy9CAVSugeLyt+rl2QySL1hvkx
4fxFmgGv1fxSCxQFSzcjJyFlkrVMJ6t6Bw2JapfEOBQFtfMZKxgOErL3OgbBJ3NP
hqJ/maGSJZwwNI5giZAtJYRx9PgJ+eBB38NPHUchdr1zeiIN0OWfftNnZ6XqdN0x
uKue2bV9lmMWvo8Smsq4SLZmzpgX3ebwlM6kBsj2grCikKMhrccHqsh+Rj1V+6iI
Z3BSNVDqPTfEI2VNWvRbos6MGNkPnPkTTS+ppsi6oESzTO+WRNiDiwXAZqb2DXSA
EBBECxPoI3pM5lirW0mR7RSlDNjr1SNY3T1hAqv6vEJRxKuq2n0JhH99DcnRlPjK
Skk1C5XyhQJI5syYXu/FBY7J8M9LF+rxkPKBFpaXhEqw5daBRaMNILpmXp9hfNVy
FkwmuTCxYgzoEwMHdJ1MmUp62sUeFF+iKLbumrUJEnJrwMBZ42S+LEZIf3qtwbt2
4gTwZXgITpJryMfHsvK/EFUuqbAs0IojZGl+Zrf77hpxHZ/xBVRCzd1dNBDQRN3s
58lYtMADk3V1XzZlkRXR89LizUIAFR+Smm75Pp3s+kA+O34Mk+Y+pu4HvJ9N6Ld1
7tqbaFjvxY4kaVtfJtFjOLku3DltcdhCZj0a7+NO/N60S2sr2mfH7VeKFeieOxXn
NMkziw/HGrib8Zy888ywZovwBL1D0KUycDA5+RAfJKzNo94qqgnSQRL+/Lmr4Y81
RudfjcRAgZV0ezeIIDLCYi/frDwloZsyI8qBeyAhtVxZ2UDE3sg2wIE7HokmiKC0
pbmSTlhyDMZVxrmLL9vPs75I1rTNTtqoll2Fv8Dp8/0OvGUjtFkNaciRh9x8kmNq
HHLyDGBBPzXlwVT2hZsfVp9dufnszsEr1Mn/ZLnsKV15Njtl/KgK2y2iz55yWAyx
UpbsgJOVzILJyLMt6wqw2hiZUDt5O2ZE0sfwEJl1dJVYlwDmFZt2yfiOq6FcrIfR
hEcYf7SvPb9i26osg6WlrJGVMQ/MNVpPtHVt+B17oE0FuTZZjcZdQC8fSJxX8chJ
pTzgreaqgzkE4SrTe2iWyx8D4xftzEyyK0vXPiQScdmD9FKNaKRYHatUH+pVzIwV
SrXDCI2MHlNAzODSQNhWEw/oiVGsFXuOlXqrOix1MVE9Zx0jbp4TKKuSvmsGyBjX
Fgv1+cu7vrV5Irw+s8NrOg98r6T9xeIqRpVm1CNVlZk8rs837JA6HbpXQ+alkbZT
Xk745EuNlcUDs3TwtaLU45Ne6QS/l3gxPSRi1m2bmx+bUqPMyVPMiqgXzKr2NCQG
22iiSdA7rIFiMazCLhqh3OUwwJCI0J6xBvn72IW+4XbtEobaVzA9TQ3XtGviGeCw
FhhxtXoAEe8UPl/rLQJcgac5zL39iF/ZJFKKy0Fu6AcMEgSYTg8eilDt+ghsNvPM
5T1FKZ5WgH53/7BDDoWshW4aPkn0RijY62bczUD++2jVmY074nMjkBlncughO41o
SUPBDJOrSILmQFrKtVcEUiT6qhfPZGvrRCrPNIaZOrTEJ4B5+WM1YsgXcAdDc008
Lq3a7FKP9DNDpeENjL3W1SiM+xQr2q4hdRhgIggw+UB9r9NQLpm/Mb9FpleFBW6/
cwO6OvSblIWNctV5nI6NnIxAAZUOStAqvDYq6TRiGs1hOexPBdu1+QdMM6fJNPHQ
749NMeK0zijs3XLMJf1UHATWzSBYyAuRbn5ZQKY4+4e0Ysy163GVbcj2PuLUuudb
zoWP2599E0d/IH7/Q3x6mCwT0OFuQDNVSWizA019XjQTsuejRfcje5RPrKULuoK8
+aBek3W/w7roAfnWi6R8OAzae4PCHHtaRcNgqDyXN9ln5dOJRnM90Up0qL8sAh/T
dkNzDGH3gsVKNvh50Zp7jP+YmXwtO68mrJdGLJDBXu4Gu2t6KwaHw7Wh5Di//4fz
t7JweAcQn4QnbRRDau4RB3fz4XpUDm+xwavpyIHywFOTib3UhE1t9Ec9a8ltMG1/
tZO7W/0CcOKNMup5lNBEBRSSQBBG6YFJ9QG+dOxaykv7cKmr1Yd8p+ofH6kI74p9
3KPqtImucAFFoxDMzmE8n5/TKE95G8M43dzUZbjXFEC2Hf7sZDqNoAgG+YP2k2Uk
2QEbiOb8j6zuFqe3FauQMn9KfEVYNN6OuyyxJaSLE8Mi5c4HS+7mQLPMkyc82dkI
my09pHQqlWxf7wzZ3TziXaQ4Nv1lEcauBRIi+6f2o/+uEdsTkJ1/ZikEROMeqKwN
yx17jk++CVd7GbgH3AgefH1mB3zdYoAppqVg7441vYn+8TXhB0Sls6m2YzIsLWoH
njG5dEGkuIgZb2bk4yteB2SKDoqw/1m0FDZvCYbmc6MOq/Q3XUfJrfo4VQ/1nTRU
b9+FJBkifa8DXDmbY8G5+0tkl6hTP9moHo/1BD5+/LPVEKBXP0c1XQTL/spoJgGa
QDBVKmRWits835d1LQ727Y3JnAibynWX+eW/5XRX0NWAAiJhX9JO0BKQu54e4U3g
hsaL/dUFYThH976jNK1fi8iJVDwlIA/SiC3MgLrsSAD3BmPmvhAIE7tCjWIWZEPe
1oddFA2+6wCON+BSLDWSt06ta2TxjtrSj2kwZqJhaeTZAAVt5uhlGVgfR9f3sNdj
14CoxYMP9f13jyIyKbhSrB29I/EYvgWwhc12MGNJ+GEQfF7KWXNVMgbQzgmtpnqg
jQAwAIELqNPPfl6dPjlUkDKyDV0bCe69Pu5/HYocXXvmZCVL4E+Pot5nH9hRIyrs
Tnxu8WkPGNMKWVXhr+OWh0B3eaH7xZbaoY/xp0GjAmWW95cJj2xYfXgKh9TAlw2Q
X9P1Bw/pBZHsCJDPR4gCb2lFIlPz5H62+/3qneNChIx2W9CX3B4I7uA4erasG/t4
bsxH0ZtIoyz984i+BODCy/H+1Gnv8HVgr6ylpcxy+4FZ/8V44vzFhImkBemOR6YZ
hPwF6W8T8XdHIZZGVUYnmXNRKjteYxKxkGFzm2T333tZbo0HlXfAvUkAr7ErYSGt
u0jKZBxcrIpKHdIfp7rq18zNn+DNHePWqF5HuFRSRMLJCQ6eu2O/d0fOdPVN8bdm
gcgTudJydZ+VhfyvkbRixNI1m/l++7inRmnS+8opIWrJ2hD/TZxGR5V0OmXwHlAR
7ZySm/wdlB7lX8KAyCEOZeQ7aLv1eblc/Ul23toIBBS/BeoMJRqHzD8EoacV4DUg
8bpfUoAzY9is8w4T5+owFJVLAFvAKA1kp30MReMES+wSyFlMIX8H2kr0iVV9C1ZN
mDSXOGs4n+0Zl4TDpv7Z4cEsd6XMb//SyZ3iFARZHvuuYIyd3qodn5C1npHT95Uc
KX56acjqa3J8R27ppeHdQPUrrVc5eVmJyo9uAHQEeQ/QoKOg+UEmDjGPFSanA8bL
0YJa3McDICvKQaWWS+uP6VmHE2uObeCdhGzgJ1TnaUQLzTcesr9yOCGieXmkqdHt
gFg63NlS4M/dkfsKdyiWb00VLEqX/5Gp7e2hTm6u0VQhLEVa1NMIJmctYmvSrAkH
V486xW9o9d/lJGrvte6VHpVaq/UF/bkf3O714vmOg0c1Z2UasoeI0p7WIaDjxMjj
rchHBIzhEP2CtKojbt41azdTXqhlrhMOlrUjXTq0S9vRr4RAxckjwLZHC7NNshZ4
P+JNDuPOXkq+0FgYimo2Z0A3x88Qtptwj294igMcQm53Ds6RxhMTVOfWct/0naKL
hjOooP+Cv7Sxyq9iOlhUwCYRk8OONrKKLMtilvUqg8SSskY14/dqUTkdO2qif1CC
twcNbS1fDRuLW+1ubOllyu/+5LLYvx8saRGUE+Em9ySxoiqkjSqALZlargMNwP+x
pgZ4kOOgAI7xwqI6528VBAG/fDPX6zFBfcTKwL/CHvPxDua1V498lRkoL45su7UX
7PP9MWMSDPk0Y5+aF6sVk18PnniWdhsqjx04fCTjEn0ddnmU2oMHyhMwwNjpRfjD
2pV7wariXIYw/MoXSwXvZawwnvSNS0TuSu9Ocnh4afKeaZd/Sf2q8GQCFOaCxE2Z
In5nOo5keVeqZAQj3J+M2OgAC/HS03Ip0EjfciXIh7fpsqQrnSRDFjyOxNeGKE1o
EFowtf9rlMsxVEeiqFJ9vu3/PoBNvgnDDZ+c/qY1Tpd0pYbD+qsTBUTpmGjNhCI1
ws4f3Fjr1SEQkS0c+7gmKjSg6Fl/VPe38dBKiXz3sC4gCYQjYZ/MTvge1haoxZEH
ZYLx6OrehqbVwrtTVk4pbRABVxHlETWf2v0S+u+lmIO99tnUSw03jsohD+WdiDz6
Tm8YV4Y4srXFBmZ9ZrvcYNHHBAqwXm73Hg0+Q/niNaVQcMCmE66aGD0Fs5JyN2dg
AB3u/6WwYN2j1g2MnuTYnniG4f7/NlakveFet9dbSXWYoqwAywDq3z+Nhne6B5aF
HQPzxpCxTjJoIQkc30a36BIYwm5bB+B12SE19btP6CPLc81XnYKU8Kr7JDgkR7Im
1IKkW2uA8UFD1VscTJEMM6Xvj2oeNivatsBYGkNJquBBE1az+5CLxeEvi2PZBOJw
/xAKnSNg2Hn32yPq1Gq+4OA4SDPbDC9HtBFpfgXofPul2+neukrSVpgawz4VP1gc
6iYHtpuOgDU2+EMiirH25FDsUMVS22VG6qv95Pr/A/aJQSgbs1iUx55FpI9mlt/N
p/gI1y/102tZ66BKhjjLagufTJxANo7VtBZBAItXAjR9s6EPljsIotEIl/G0/bL1
qb1xRgHlrcvImkGBhXQdPOp+MXX+uGatqMTCmHPGd9+rRChERywN4bTfuPQ22z+Q
K89UwSs0KQrNpQBPrE18xy0MtVo2HM+L32FUdADIblGOFacquO/uIT9Y58ojMbRz
blDfOmGXHzz8W11NOgeNvZZiSODRkgBwqL4v8M1tu7LAcCYXstiQtP8mLjse+JOh
GuAjVR9VNPGkb9xrZMlg7NK/omAm0EO9FGrIy14+rEEQ2NREhCZDJ5gu1eKTkffv
cXPwV21dgrX/D03fowBmHmtO79nrqw6tNeLMeifXxgTTU9P1VeTqnoouZsrePL2I
HXLGil1rIqhtdp1bVQkvd1ekRM0/Ci5yYjWrpsH1JsMDvNxoDG+/NTEliHpXagYz
mJq8Pz79ABy8LoO+xrznimQJuTguo3v1U1bvZlDM3ZYZcpb45n/73ws+LVrvUfCl
yBJ9qZlAkafvncBNZF0RSH0E3uwMbvuRt8/USMWGZEkJBvKrrPunmS9YEiES6ipE
F8QSzBo1SO4NrAW/cxnMpVsXQfBmkUVaE6QhRsV16ZTlBYDUl1kSjEHMi7gohroA
XV0SQhHg5VSTz3xqSV5tUzV9uFM0yo3F+cMj1dAYxezriiWWZ7gzDr0Zl/xAE6Uj
85H+ku0ZVezQE1OeG5oKvQdrIFDbdBVdFpNK403OKiiGWD2/E1m1El3gvXIA9T31
BVsCwC8yDDX83IFhrnRoibauXv+6WF28nI5wT1eZaFYstmbuARRQzLj5GGsmt6qE
im+Q6djkEBjTr3/JO9axyBtw+7wPpxdEmwSrqVgKjf2sCTAI7gpgRoDYMHOqxSIq
exW9Zxbo9iq1ZwjcmUlTR3hwgQVGU+gcVhhJQVo3yF6g1ZSD7HpGmTeqsXLYpbr3
rSe09JcEVZEdFsjuAw+RY/wa9VVZ5Kc9IKv76QyE6lSUoDSsKBK8VEo64kaj9jyG
s7R6sf/Vgxq28Jl9jU0XnN1GpQylO3HelhzERqxd/Iu/Qscruoktfl7JvbvgAr+l
c/QhAJhJS+OLtJTp9bGh77Kq0EW9EIzS7qrpJ6w8iFDd1jRFf2hegPZpEIL2yNAQ
a0SfMjwPJ5Br8RnuciFdepgircxmSGQPe0WDeVwSh0Vx64UoK+sBOjVNtOV/bMB/
1FAZnzLgqjamPdjbxzahjNpO2fyEN/V5AreANaEUV+w3fwRJw+QfRaGhTOdvR11x
zIQxLzZydM+k5fCoNqeMZLm0FRREij2jl8jvt7BPhaggtbuXy5jNtwnyq77JGRja
yD4KFwTRh5hPj5/JTe9QR0jBn5tQDULu7gs/X5eUF5MVhWfB3deqc160fvsZrVI/
DU72D/we7acdwp2u+cEUD0LCz6UutDdshTVHwnNrN0q8VSPMCoO+Dl53/+ho5t7O
6vU8Mf6t892IaEJbIIgr6QbRt6OiTXRS12Lxi2GByDuimG67x5xD5jtf6nUECHfw
6B5YxoDP7sIYQ3y6bBSm3n+NQtStZDmrsRm5IbIEfEsyVJz5Rg/r6nZfaQiN5RrW
ItGwhd7EMi8cdogJ+LvwAYi9SEoHllTqwhlIG2gP1yR9MWns+ZBl0hIJVmqvaqd/
AFaJzjzrhP4ZquXoltfvJLIZFv5d8nN3stEQX9hqyyGiagDo2zyCTtVUIvL/8amd
lxWXgUxFIekP3mxbnm5QebamMRxyNyrj5JYINuqcQyWh5yphU8H/8a+IMRuOwBU7
wP+fgEyN3i9zvPkl88//PsdZZagNagbFlsAECNxaVWmTk6gIS8PpXU8WLG72QKQ2
VC1vP5FYuuFNofW2BKYomHwT0F668tIGyQxWUJCizrHDzzkG+YsK+JWBRZYbNZdW
RsC54Op2CO7IlmlLJLNPts+2Z56aEMf/jvEbVf2eqNXCMqSj19ALl2x4wA1MJpgW
ZJPHMZdL0Fb/cDEnzW28ISVIPFWrDxDAmTQJOuIqv5urJB4ZP2iexL0bH06awRu1
m4wrYup9YYdoXikfajViuKxWWI6DFZl3I1crqaQXOBwK2plRfYoK1iJitOxK4wqK
LQdp4D59a6w4HK+qv7wKanb8ZEDcotxWG6V9QEiwntVAZxlWwEZSja8dxYXEnd61
/7+li80hIuvZ9uxSsY9kXb11t6WSEsAqzZjdY5TNN9TFoCb3EX35vjPp/oItVXvk
ZBgYhXlwpYREo/SlsKKCR3H8IN6uwAalrF46fWVlhxSL3dSOxZtHT3deN6ajAhKa
vb0gL4Z2epQdH8H9mYl0ciVWSZY7rInsl7ThG5oqA7hh0heYz5DQKetjqgcZrSDF
avSHXvcFYOmXi947FiNSrUlUxkgXVO1DXq//2jGHOrigUj6HmhkQQNc4Il1QhDeb
B7nQC07tG3mRu0oXio7jmIbQnZQ1U44cVxKcXFnpdPGzqlrLqdz81xXGQdaIIjJy
tAZSel4N4OQTv8/FEpTHS9M6rQqXa+bP42qv4dGxvj5+ChAYvC5qpVA8/BQLvqYl
qr0ZqoUpLEsp3R1FFsc9s8z5tV8D81sZoPD5eQfBBsZnG/ujdVgNQBWgFvqYmoki
WjC02Nx7JLmFJ1ie4BWJ2bNhzuBG6cScYO7631DAjal+NZkJ+PaEM2q0myBI1zCa
62guu8KnzIk0FHl5q7Tp41bCa+Xgf6Ab5yBUW5TcFmPLiLMGWeWxzstC66E925tQ
CCvBJau9co5MKmTf7kkbMPasU36TcvrorHl51cJS6/j3fsP9cjRMggqd+F4YDhkZ
hAzcG6vLyMnsgArmZ7trKMBoXCfGHnVd6d44ecnQ+kaVc0QR6aDU9wDkTumZm/Ei
dJnyKDce+CTq9SUAokIZeLRJMUz5JaJhfVKtm8Gfi/qN0AZe+p4hgTozW9uWgiFu
r8ubXznsqsgU0T+uixOZdUiqJvogIIBtPcyMcVIRIIvfdZyHHJu0hP0xLfgc/xX4
xpEGHikqxffnQZ3OlHrGeKH4df1tTom/sbutayHFdQaVF0mls3xo+8LF1ofaHzAA
c4JW/9SCFuvSrPeBGan/W0pvzldvyGpEeRKMtfNkNNMfNzuNkx2QR7+PRWSz208C
ggtHpKzfnwoipitIP5/nnU3cRKm4H4JGGSCmRrLw5SeBfajk12sUDKcMEmYerw4z
D9QHw8qLpuuWoRR3MfUPjI6z8vTUiNkbFY+XK+eqZqNdt8lzgU72OoQvGSqDjCnx
SNFqLQyehpBvkW1zlW2Zswx/qGXxfMmWfFGcJkfqWaZD4vkJBaumUn97fsQMKkX+
XKu8uMaYS4f7MIzlPmoLv2hP8lIOr3jGbNytByHoqkKyyrEAat/4kUPfespLXZB9
rCE6iQnisH31zAGDV+6I6KmkstJxYgCYKLFjUnOkRUr1Yao1YXze4KfSN0+7oWrT
RJZuTt2Oy24nSnC8bSiK5hCJMJji88uA+jL5fcom98TwJThkCwSDhTw3fDGmA/xp
PNK7upb9uxkW4JGF1EYVtQB3p1poj/YqocV4GUyPvhZwM5C6HkFeBVpt8639q0i/
lZFYArpmCMn2powNE5Dr0PlS7GSBHV7qNKsdv2u3aCVE5FLyJCTcRKxvD3L2oscM
Ch6MgDFpSAe/XOOpzpyydfLlaivba2+BgK5AOc6AWIvMEVcXzP5MzOvTD6zHcuxb
P+6WTGoyXWXgrnmYzzm20xYFgJiJOttKLgse0GZDnw6m/RoupS8qnSOY2FN55Xz4
0ke7UpL9rMg/3322zZ2cjXpAlFdKplPBCDtiZxdWY7NpQnmVGYkxr646WV823FKl
Kzx8/q+KyKq6R44KQtoONr/I2NESUiV1vIXgOhz19vNZu58qY2rjaZy6+5jIx3F3
JoXZIta6AHsdQqS6rrXX0V+CqnEqk89TmmHaAAeGKAr91yiUhhBJtwELC3BRTPHB
uRxznYRzRLDoUyVaG+x2CqOYJfFLl79iLjXh4k7oTi+okco5RDMod/5SRLQ4BqQb
I7PRcMA79N2a6RMpDG7ZeaJHfg7qJ/uWyN7vAS//FhnD0WfpMdjl7krPvUfV26v7
KZ/BJqubZWZ04gdmch7kLqns1tFVRJh4JgVskw64BsSwgouvqp1JhtnDJrwEV/n1
tOulh1fS25G3RHaGoWpzmQ+kO/8mnlJkNeuzlbp915IdhxrFaLpNn3fGtQOGRe76
g2mrBlRERJUCdjUXvJ3A9bQpfISEdsovshVNDXQ5zM6yhahW5TTAGidyTuIP6Pfo
elZuDbxDTHKfvgHV13CHLkoo4UE5Rn2Ksda95S4+bxuDV8WRL7KIK3zAqcfwmYPt
/lCnAJ8L1paLdfKlVu6vhCHyOCg0ENu9VTEEXLYKBXBDQX6WpwpLKAj7z4a4o7Hx
3XWX0JlWwYDQGN7YWesvYoSipnSmt9V+nkcB3lhyB85pvfvuAsoo+QWy0WsTu6Uv
Tw2PEMZcQjzWVa178xVTy/TPJkZtWkQZKzUzdso7mbzpCq43lAug+taQLUwkg4A8
G9FLycAAoMEX4sNLpJNoiPlja1V0R1uO/D0LkIMpd6IyJgQ2vcC4PUY6JbHXyHd5
ppKwYnBDLU7CahsuBR2We3jG7Qxx65hxVt4GbVo42lHM/TlR3J8AF96JHw/OT8YG
E4ZWDjnDak1DTqoBosnFqblfw56eSBxCX88GWJF8iMFFSgj/nvNDbChTmAGnAinV
yRIsd2Q+dzZgITfGZf+4VVPW77OBlCINJ1AvlTD5i0bAvk+bs6tOmrFshAQbedIc
xTdqxz0FXyf0SmPsLafZE8zbVUufhUYu+0JjoKdySuIOiuHd8nE0ypcR2C969hMr
j/urG9kWj+ofrLlOy3bsY+2wsLPT4qY2xEqdePfcmFx05Rp5ou5+2MJV9pOzQNMK
B8IvzYE5ihP+S7MezzDMX1lKHY7tm6vIAeVHGhqF/kRgAnAzJSawM9BLAbVwtrku
jV1TOLpQh+BE9KDxnVKa3DoBQo3era9+evheJ2nrVwH3gXsciWTTw5osoWQTLVFM
6/UmGCvMjfOJomN/2ubVaL5cNBW7OsOI17Qz5lh/D6kpWqFU52VBSOImP0tsv69L
VYGbM58dgRVt0Jh5uBePUCQEX2HLVTwqoSYe8UOaUqIVtbRANrB5jrzgb8/qd4Tl
3ajezPQPlMSVVE4mKg9nA8RKssBgdWTcbPs+jNqtFAXa0xU3aR4Pp+ErkabQDxj0
68haP12zZQmop9oLaQbTchKmD+9J4WzheGPx67akGzgHZcBaooqMFm4y67aAjmxj
Qx7usTCoZMpgtDRidZ3XeoWppQIceNsP9KlVnk4b5npMIz5Hqcv5iV6rQR3pYtiS
VAkaBbmlVDLI6y4vynedGn15O9reW9J8b9bJgKTBqFQdxHxTsHC3ksa7acATBi+H
cdbRU5fH0ShU4JW+pik5DjP7dTztd0EkxZQFTfSWNIydstY29TUdAwIO/cqgLVST
kjJFvE2yxbPszrxzn05VjUUpSmetlMNemUrS81GBTtpox3BQGp1pokhxCesJsVbP
+csSkO2j5KMSV3t+CYUY4zmVfNvaGHJrIDInOfjO422uBpQBeoHfaWzWZN3UGZzY
E3oJ1CoTf5zhtR7ZxwFzgD3Z3Al4pugOfTMAcddvLIqgTUa79r25XGCNmtCXVvO6
7323RQ9JhUZTtpndCQQRaP5s+o6bEzO3cl/6YfHIPz/0cDsO+373bkx8hZcaLHaN
2kUBKgSPJPSDUKxzu9cpX16+rgRdDoFx8VLM10OAeCvCqLxDFDNgQqNlLCqOi/n2
N+8Yi5hIgZixQwHqfD2HkJLbI5Plz+nmJyWpuwwKwwYAje2ZO3jyO4NAE+udbV6w
e8EZR08OjODic/Fekc4HQqv+zzbvG6PpNITUBDjpfYNluBgR8aV7qb0a+K8Yyyil
S7lhTsnN/Hb09mS7PN0LVeqcd3c4xrVF7Lv/LuDkFdo+gNB+CuqkzIRRpXGIV0On
ATJpU0UrzpjFn1WVYLmW+Hz6Mx6E4JIR3erjvJ+H0JxvhcEYuFrAp9srMzyeJWn+
1FE8oX28p5oKoGjVFdruI0hr7mUG811NnPmtBgssW4gXsRO2Or/hr+DivoJlpHB8
IHxDRvFtsedLJPrsrJ2H0rOSHh9Fko8os4S0mXDK6pGOQ6W4GlRtZOnvJZswjv9x
YxhJFXjSVcP/yqK5gFWgh4g8EOweMXqc6eszXS8VACap8FldALSPpN6GuEuSw2Ar
3UaOI3l0kTky+DnlnkzNGrqjXJATWk4Gud+HEitU6bzZ2x0FC2AElUTEQNA7VJmr
LHV8M8SmChlbOyVhJ4C/X1vKv6xXAmotwEuNUgIIPWF5jgxNi2qktaZR/gA/EXbb
ens2igFnxPXDVusxsgs7kV++SIexiNobduSphJ+1AeyvPOBBSo9LVslQ8yA7JAmM
NcRjgEQmZ2oMzMFr4BrIsDPwdda0qqhz+xl2z/5KttI/ZdgFLnzQ4K4nmYo1caqT
106nTL4SjuSN5CiVmKH8ZA/x6+zvCtBIpkUoIn5NVmcxgICQKifnUtGz2EOtwcHE
XueVGEQLzg5xGmnKhe6fhcvx65nDruwHuMn/9/n7lTz0df3rHMulXKfzl7xQhmI1
28I1EuuS77J73INU/MVF4Jp8G/3E/MHbJvPlNDOmG8fs8SiitV+ZgrQdOTcXpPIW
dTzpxDpCK3ajIxrTR4OkheS/RuhVw73CsU3f6WFSfBcmBHVDJkmP+IsAc0H91LyN
wNnAX5vUlFnSRXwcLu4aRXTQB/gUju4b3Py4rjsBH2Qoixg1lCjUehtFiczGVfLm
UzRG42e6LKjyojaUcfCnJv1S/F5pKBwOlc2/FrU7EOnq++lWIbeW2yN0C3noqOZv
ixqoJRT2sxrYAtVtR7sZ3+kX++eAbVYmtfGnf2imp9TaqmAg6fPHhCce/+ulEN+7
s7rej+bswHkAsgFFMoZE/fWE+LCUg/XEXRLOfnNSiFFQP5gRp3BwCq5xOIWiipqi
7qJSlVK5T7i6oq8luAuLmnDdOGw51quHJDcBlV8O9B+Fv/P9CQ9L6PM5Gwu4z1G7
DzAuKa71Omlj7910lmNjM9GPBq2pLb0VnSPnYg4AzcYuC+4BJgNQSfH9f+9D7xxt
Nj20ipcbc6a1fo0md9qobYCciuBHshDIv70nuEb8qZxyLoTUffjT/QOvc03xujk4
efosxIAQVWIyWZvZDm57HfeeQKK1rTA+WkXcbq7y94iRV0hCO7ypmLze8dcKrw6d
k4TFE6hZ5NrN4yGBKgACXJxGgfdDYPMZLlLnqmgep6Lfpq2EG1KIFHugx4dHtKjv
/KuV9R5mPG/3peivLuugOTV9UAfqzO9JGlT6pWCxJahXdATbi1FiU3gfGUCs3b25
aVPmDDrO0dZD+fC4RAwUx1YPits9Fvo0Z4Yd6/YeFjYxzPEx25AYTkxgcRSxURbr
BTygdqADoywGS9fCFrZlUfx4GUSA59OYFIpElFA3Gel4+XtjnqUz1OoppvEjzulE
74sfoMADgRzZayNeBDG0JUZQB6nV4p9zrL6XvQoxN0DPoEWa/27B4Q4mkQU4a2mZ
hEUlYEedtV51TTbh2R+qrBB2VoRGpgnVUgfoQrA21Nx8STVmQpfn090e3yF9GAZY
/5mLCiVJwapW8zFtky4+iR60KXKLYrxc41BgrpXJpP9cL9kZxmVL5sXuoRwXSGVX
aG+TfSK+1dR7IrQrqbmN9JGTzGawr8IPwpwLf5QRYg1ncfPDP3pVkn9x+lbA3TeZ
piEXGFJQxpPFcXlnuwJKNDC0fBFtQAgfGTZ3UHXtI1kTJmZ6pgejcIZ6Wb5FUs/1
sAga9EDAWgrcL90QLeJJH2qvr/ruC4U57eK/+mACV6ixSte3/XcBVCze1EXoh+gx
ZhtCbvONcLsKjELXkMe/Yw5ql8OZimcqB/ruB8Mm3MatGu2gM2fbGQ/Pg8O8Jlb0
s52qjV+3TInuih00dRCjUsxJyySUP9tmyGnb83DYsCTAyHgMjWkyJbRb+sqZsGpu
KFbSoa5tvzkoIZ2zZexIOILHS73AGfyWCRtwcB5iCNDeKbPBBXQfbbegSY0J8Bl6
tteFYgMA2m5jULGm0RyPsNBE0cdj8mzsj0Wdy4DDhjaH37NYxosh/8YIgpzcQfub
7NvAyS7zt80iP8piHX/LcV1bEmqTLgU16LAfPNN9R4Be1Lxa3CxSI9b5HRmJmpMX
4ef3r5Y8F/wuDBjMyNVoarV0zq9RMFnWFxRqVIDsCTkYxHbdefgSglZIH3VOLOne
dGEWBWg01OncxFee7n2pupDEu22F3+MySL7WpTLfhIwck4s34rK+hHRTCe9wUeYF
3+HgzDksTLrhCxehb1s4GXBMY7LBXugzKs8fqZNVgz/FGrSHSGu7ALFcb8kX85oS
Hh+0E4HARCyjlabwo5u7nh7yJWc4jcEifvOoRg1INkOtVepJJmeRSacPb5Vl60OK
mud75nDEZh6sTIIQFjO/csyU4HOMxqprAFBnFlNsF4B3BNlesoYCaHq0ZulA/zHI
IJB/0VfeKhWtGA/VRPkbm/qfDqtYLt8ES+gplXilZj9daJzxUgRkj1L62gHFfW2B
Fb6sfZKO42296TfursIGCSVTkPT3+LuYvnEoetUfW4aD5cLDFpvl1EmVZL0J7v/N
eHJVeXxYTyyAdzv0cwN0N936Fxfwdw5BIffkw+6SNl+gIInwVnJqlrxQIEX+B3Va
g8fShKJJZct+pSZEDrhnyW5cSgxUC82Uw5kXvQ74cuaP+naR2ax1NkIUrcTOPA3v
U2yqpfsNJeoCp/+1aiwe2gcmGdT1rCihH1iekCj2Sj95JsueP3FtHFeGgq/oM+1Z
lL4C82YxjT7JWpU7wBQlrHq79B1E8dOYzF31LwyJiR9J4FvyKhOOdvHZM2jADApB
VfgkdYouIOR9LUQKMRpz1ZxVtaPhzJQVY6uP1mKv4M4BnF23qigMO35xCTt8e/v1
c9e4Vyd5Eoq46/eBGZXTVJdt0RW0z/l6NKZU3iQey28FwS6OHNO+v9oeMaKtXOR1
SyCuD7Rnvuhe8r/Ak1MXdJ1CKV/H/fJkXHYCWmY9t/4LXYUm0dlvPxnM2cyub2+B
dYDnUqMNptU/rfyZ4XQ6J5q8XPzG8ut4YDjh2FD+2YxXJFGbtJJXS97vrqr0oT4E
MujbID/ECa8/a3tQo4Y7Qa0DGjaNSg9d+vqY6KyA9XpYqvIlMkRRK+I0ZUhHAX7b
0HNmS1RLwwTDhBnahi/APQNB1OtRDg0QM6DC9JC5AaXaQzmGtuncuUhg2p0MNrBi
CMUR8ojbZVtq6hGO8pr+2uS60eFoiYqU8bq/mc3p6WLw/9B9wSWrzbXcvL55nqlC
Ug5LHruneLZI4FYwr3NCKh9MaYURQs4C8D7I7uw8lHjnyp1KfHa5i4LDrOLvUYrB
f/qk6b6yXbw1eoQl2/iVXerDSJfuZZrGjXolFHo4s4IFdAaHTrvaMq7eV+Z4uKEW
6z6b7aqCtfah7b/smFhzU2qFYSqR+hhJMMeniLB+KKcy9sWlUkYjn5C/fqIprb9h
iqkUXi2uroC1CihzCtfGDhGjdHyRw8xhROeWkO3qzQTMZQHz0oGABBrB532jdo1i
omUop12eiPJqeJbNRVi16fFpjKHf3KmowqDjaYFNv0+qxlvK+p5jKH98+JEOaHd1
HxAVpnPkiwE5SK2OQKtaEzPtU/Slz6OtqwNBwgiX+tA1yuPFxyJh51v9UELOqiRb
5GtDR2VaIHXubpgkbyM6e648sR9KsdBmsO6gFsdlstEBSf+iuYSjLrSg1O05EXtf
nAT9O9XrrxTEI8RLu3HbNcJ2jfrxNSkRh0PQgH6uabsdDuT9aNVyFhTAtEEJO9Y3
xHlG8seZrc4vrp4jY8g7VbnFZeTvIVbChnL3Kiab/z5BpmpC59XvWx/jYPO9eik4
7+Z+293Mq9gluuqXyfGflWPnJSyfpqDK40tKR3eW+7Cz5uwd5CgcLDrLV+4B9D1o
d2ZWmo/NJmVE/o3mEYDOVrJu3Qh+rEUPkqxSaf+RjnvLoGuAXHi4WBtnM5cz+xT6
mNtlpqO80X/09HM5IPZM8iFjF8vgYABhBQ6rUpAxBz3X8miyADUKxMNx5/tiSxPW
K8cYJEe7ZNUs+wEcx1WhQ9VwyE7ruX9JiuyldnRoK4+28NJ+TLyR6R92sohEJN5R
rLXBkHax9Fu7xQ5XH0ACnM04f7qUouu6JxrxDIP5PE923AUSJ0bUd/B35sWLilMe
qW0+1JmVqbncM7JGzno4LbxZfy6Fml3pkAjqsmP9gydIFAWN+VMhwAv0wpOaAXJf
EjxHIb/hai0mZR954LnpWbE9sagVQtqwfvKMKw1isD0tOQxld8qbo2jxGFPZ3swq
X54IxJeTQYN5LrAOF0JGTlv01+Vfg9bzRhTkfP8riU5NjBadcRqVLXm2c/DVMrbm
Y/oMUfiinHaEbeiXiKtlUdLv/VkioBOZD3oaBK4V1PI6CmnyhKRKt78mxBLPbRUN
zAz9eNi60UZUOHPT/2rRhLg0n5/fD+dyNP6PMUhPlXwqxUTMvufd4wSojbjBOmMO
nUYt15eyEdL9s8dHHLsltW3nQlL9i50PZWSNBTEzadh/I5J9gyeQfbpfBRzqUSev
3dnKIQFF5k0/zW7GoW7zjgcUwMZwNmmyXjDdgQ+SGD+qXi6YNZIvLKbkyBh4nbMS
dqq4/I5UDfF3Ixq3ltQEZQ8Wb4QWzxLh1kx/7GxyH/GXSJr9QCfu0TJABUiByk1g
yCxWABRhQkdnpLLFs+AMnENV/TIPMCJN0x2/rGx/vumuRpbsaq0WnuA7bWLsDr3O
sK3UBA4NG/9CcfyUTwRhfWgNe/37t6ZQAXth0zKI7pIozVRfd9v7A4f7wGszp5hI
ZYgMVwAnQgWxcBQMw3vgnx2g2Uz6bRfTi+UiJbvlsv4/oXW8U3Rwo+a3OrBnigfy
skeEc1dSad1bGtioX4XXQ0Pc9BJVHXbsa7p9r8weB3A+WYV6CtOIvu6rJ673PMyj
kFrLAHM3GgI1C7pncijI7dUz2dqXDayR11JicvMBuALUfyIWP4CiQPMu2q6L/qt3
fRHuP1+CGgY1EHZ11Ezj4jxSwVfyg75VI45wZTZR3MfU5rX2Md8b1Op4SHfBQqw9
UGM3gTZiZJta/FvSWr2U3Wf7mFph72JC59tz907BANnIFwZ257SCkhYP+CNO747G
PYaP8LVs6V5ZwrYg7hsMN6KjTFBquAQtq1UEMFCRQCwL/Dcrkfg3dkFkDf2+yOhJ
JlYfG1WkG7gh5kL486syUiQ66+vgc/yu7S+8A+b3PwkjUCNTWj+nug08W6TT5Lci
ScEsm9ugBYefjUkhj8+lcCRrl3/p3Zk7iL3xBgZD7as3XoXHIAFihQVYpmhU9D2r
nWjWzL7h93G9AHJqlscjY3QBrQihEAuHK2AYCo4Gxp31a9TTZ/0Ksia7Dzq0APLs
Kd62Nh/12cf1oc/yUq96AuEUoryPYvK6oxXd6E39JVMNFz+qAoaGus8C66u5De/P
/xY9zVySC1ELKnlp4NWcfloSP9KcvCGp1u59RE9i91Cn88nzIv1qZN/DmVgX4H5N
VmwuvPYR25iDKsF1ETy+2Z23nVZW+SfxhatA/mhNz9bvykDE+Jg6weoNhXAwHF65
ptu1AsIpkOtQ+XWkEGG4ld77dX7NPezhsP8hZtk3CYiVdBKuIJwGJ7csgdtgHlgu
Dog9OB9CI4oi8fwR+TEYrulOjCFqQV7kYzt8mQT/a8xIwwekpasG1K6RDhJyedjN
3T+tYwHl3Gex7vifiFhx2KBZ0QGwl2okLKX4sA/TbQsIE+eb/nAUF/k2vXNqunWW
fHguewJParky6mS6kWgwbwAAVJoHA6VJQNBtwmEVJiZc1wKkvj9kwRejIX9Ybj6b
jxMfEwuce8719oBfPwT+tIU6v8B6eOBRFFAls5yGqGU/2S8L1Cl62zShXTYiMIgA
PeBR0Lo6fvNJSk9TO86Kb3lyWx0jCfelvQYq0K6KO+JImh17jNgzMYskud3mfPrA
dGsr8BZWP4bIhN1NNwDKbPSixr7V0HBx7QnEEZ+jn3vWsdu0IgrnvXV70KnEJC9w
AwNM36VQnLirGsm6xU8PBNm5HuA++xAqsFyBtI6mUy8XUKTms50S0HixYiqmv8vI
drvJriCcKGu+b++PSFX/m5yzs2PRAkmgLlUL6GgZ2VcuoMFlkwygFJ4nVcAjsQBq
433DJRtzYmyN7sdrjUAR1PVfD58qh5Y/8W3B7Qrtat4tIcxLnOvKrFySP+ioUaMh
nh6aymLIqb38pMweUoPyUxqMufbtD3UtPBgX893k6pZKqL4cS8pKmXEM0XCEhOHC
yQpcdIakp9IRkv4s+Ni5cmbWbNx6YUp7YOUy1mpFWWKfF5ucQk+DROQneUB2DxXh
FT6ema+JOywCrc2jU62+KC+3P7Mts8pzJtBVx+wXL73+dNoy9c2bfXAshwspbkZF
aGqtUqdIm63vElM4gZH4ofUUqaGqYE+IyQj0iSjaNXZKlRNMY/j2/bIPvSPvz8uS
2kRZWGCpm3/5NdhnSQPP8piGEwuC8aSd+mXyWRZRqimMEhOOxPiaiopLxvw4fywG
cOfrU1i3JKbcZi2aQgQsQlnXUH8uR3bR/+DWH2/6pjdo0EaC8MRyR+s9qwqhXNu4
YCRJzVb5ATEGCU2Lr7NaoEAdaHj/9G4AM0O8/MEmVm9lgEAPWSxey+127J6Lkl8M
B8PDS1ysXrWeor7vTdf2z9lUIR/Sc5Gh1DZE4bKDu43phoUxy+O/Gvj4hiJ7bvRN
AReFY1sRlcb9JivoEgHdA/dwIVsX1Pxfdu5eg1gvb8AV2fmXGjeGFnVfR3xiXlwW
YXwwZuT/0yXM8LabOaErRg+KLFTSokwjazrwD3JcGPHB0Ob3jEHQYJjA2zN9v9Fw
XraEJRVg65DyAnzSjzjzrUhvUdBfmss5qXae9WKh5yzfIj56fBqCkv7WOQHxDXdI
ph1ezjNVp/Ui+jDRLo/Ucm6LLC+uiGcxYw4Kj1vBVhrXRAwY9EJNVw5jVeErWgX4
cC5ndNghFjhry3mWC3wpT2h9SUV8lKk5nrJXZNYhyisWNOpooQ/w/SXOv6IH6XNZ
YhQjP3ZjjyXD4SkqhkwARXRyetoyLUfMPqo/dRLCTTJKgaZITIU97D/OSFF6nw6r
/zyrYJ/f9/a48Yz9MMsAFQZ8MRxvcKpuZoO37nuRkrfjaooEcRW/prF3rZZNP193
pDMvjF8wwWG+RXQQqjar0gibmpScjXVsZ0xNIgeIwM7mAP6w4yjUxXVhSLh4a0Xw
O6NyyxVIGVT46FwVgB+gwmICp6CCzTfIc/uanjgEEaJlUvIMRd02VEBt8d9GrPse
Kr7pLwbaqDjddIY0xhAB24e6cZRRor1SIIhg1velj6+3wW7BYpKBjjbNwIBUfvsQ
8cUa7R10JIz7VUsj3C2hl3aPSD3voKta2w/HxAMkfHA6sx49JGAErl0WtrYSW5Hk
Ln8hNlK8ujSHaU0YN6tugx8UZ44wqOcAwjSgfbIMi4BJegMRPf1+4uvAXrdiYqB4
hOewY/fxWFJ9PpzKUfvEaBrVxel4Zvjja1IPwdvf4KezeTf/cPfbx2eednxxVppM
FrPbreEZC92OPr6de90YMjLYBX0h9m98EiSauj4O0+3oXHYSwDuBVHhnujeqErvP
giWvOs+kxxUv3+E4scy6TMLYK18LuQuhQf+rfl1QLCVIgJ/kVhx+QZENPSbZM5ie
tyaDA4Q2/bWOfz95UbaG+jeAaRgVolo/R6PELuEdLrz5wCrJL6TeENqqpFBc9HuS
fqeWnRRe0Zn01qvsSvCfATfO0iQQlzk6H9oJaZoqYvchtdI7bIZThjyuzloXW8KU
EX3kw+qI6UtApdrBej9VSrc3C+T2pKNjBl7JQbnAbqkQ92LS1pFgb1T+bm8Fj7sB
5zESsEXO1Y/+t/lfYmGIs8rOOCTK03lNmDPIDqXqSA3cBcwodPhqLhIhtwmWz6pu
BgG+JFZ1PDt7N/0kJn0Xu+JkhE846xAH4E2VKAt+dnIusastuqz1NPOsKoFxOL6k
SpZucsTOtF+8yHmoxtdxbLSkBhh8xOxciyQcb7aMjCXgUj4tvIuvpxARqwum0AJJ
2SKgcaqOfezUG6gIJnXnp4souZI1QPX4KE7fNV0Pu1cukSSodIssFDVJIO34DLDT
/xM+QyzpvcFQobWIqTggBfFZY1p3kaS9uQDAWbBLuZvbCoolG3JafLtj96PF1ne7
clGMva58ouJzAYe2zeslfwKwV6y6tVcxWTLXaoYc6+0hd7DdgrofTCYlTBGPEEjB
hvZplt8UNAinRf8vWFQ/a300cTM0hocgWuKh5XQ34Vl3TLNtLMhePY++hbs6TcoJ
NSwgOEcmBfYqjjsQRCs68XzryfJQxLDbNo2sBO4poXTl+SX/IF5jWNRMdy7FVQ3s
tARJ/Ckbg1LiKfEmMQ9BusziG1c7u1McAdvnq/uteT/i6PJeOUtK+gUvpXqWDqsn
USj51TXvS/OTgUIb/f1gUkezYjDpbTJ85uYn3ELNVG2cwhuVzTmMgTKlSMtuYQGm
8ag0hhp8H+E+IDzVpmzqieybyLzR9qceLlz7Sl8tQw3ZUiyxKaeQqm9hOtDm/cAy
d/N6+2fi75Dk6W/IOUPsTWy0QpsoXBWEyxtpAjzzNgj8Fu7xs8O3XRPpYBAm/l+d
T8RlIk0J16UlxoLRICePtZrCB9D8aKrQP/joFk5mQMCAli72sXzC+AsLDkqFja1C
pQWeS6NptshBjqRw/80xQ8J8C/L5W9W5y9qMEcz2Hpdd3GL/5EnzvC2xtB9F5tum
J+ImBnvI68cF/dt2TBXZoj48A/dT77jFP/sxYBpi1GGF0JdOxF7efFMu7A9U45nf
wZ7Cgvqy6rVAUjD2cSyq8CV1CTmXzGnja8N7b/dd+kOY1Yez2VFMQ9q1u5m9ahDT
WHD/c8iELUaTTXgLxf677UVxuf6EayOUxkIZS62mJ62qk+iQstOk+eBacIASXa+b
8tBJuCjaHj5MSvrMhzJK4KUs00LWSCFziIvWIJnSao7jHGIVpl8hEUfa5U2bNnrr
WBoCUjxcanhAEOPHWYLhxYX6Wn0CyAt4jmDCQRqw9C0SsBcWPnzFe4qjWkFsp6Uw
asRcSTJ1RZE3jUaoAw3zkZkwK6iEzMxx8mHdvtyCPxfPXTYFXl5YiTQIngMmrF7s
Y1t/B/twuaFdmghUD5rAmIvLaWD2eEbV5N3meF3yRvwW7A+qB0kl2jF1YbiiSHTF
6c2DiMu+uzEaM475tz+hWPUH2lRgCNyJHmHasZirbCPfU/pLAdvBniq3EsxgG7xM
2xjouhuQLggU2/S8WIqwhAstM9i2KSYT0bS0T0gfDnysuUWhbGOWxxKAuvTygyj+
PaSwiI7SQSPp1xVFqWVm2Zeh++tIhkaoQC2blHJKf3oP81hNj8KamLoXHI2lJ/Di
hJNEoENVqjLQP3GEjiO63MKXfAd8ly0Oee7Cj5bJ7IH7v2mqdOqRN3G8ynXZ8Gh4
yj1CtsZKGA29pOQmF/qaIHirjGv6wNF5G6Wpy/QLo8VY2mq5e2uH7VqcYgwOQ7H/
w6wpcPv6pbC4OQjRR7vKQXPy2TrOgBGAPMPJ957bXNCpe9n6XNrjB8OjdcKLBTXS
XKuddr+ZlZ5mbcU7jQAtxfDu0sdm03dAo2hSVTxZXGcbgZyESnqR/ZULg/kZ1qAU
OyiVJlHoOLhr0dCwtxfzkFzKPACgc3a7jqQekTtFoQlKznS5AfnT5DwDB5KvxS0u
rHaSFdhuAW+KiSCxkU+mzm4ql3zppqENXGXK/V0tdmlA81isERExqgtiLCA4dJ/2
yeyBzhWODkSJtq0c9swHUMsXdUwUDJOuLyso09114Qk2fLKQMPmc15CUkGn9CitS
elyl0dKTld2PVOUS90+vJfF9582rD9vgYVLl2QN6tXmg6USebyFe1Qz6xvzPu0cL
YMq3ZhVKsZxcvrAMTfERysycJS3UgKH0KKtYhgq4WMU5C0pGqzU6YY5xJ+oMDc3F
1O9vyklSOAjWDsSXzKrQeZTIiiVeGx8MqGB7SIuXDqP8cMAi+YKLaQZR1Nn73iUG
ze3w+XQR2UrruKxRi2yKVTs5dERzKUi4RfoHI8/Nbfm7rP0hrETh3j7kL5dxigE8
kHwaBdNiNLDl0IuNEt1aHinGpD6eUTjDeF2eFECEcHnA8jgHmSZYdYsRcQ/YE31e
yUQQ9AwF5+J4spCKISwOoaWXU39RRO4duLv5NjKzaaAkgPQOr0egDCSjy1uH4ufA
lmpA8HgAwVsvcH8z23ST3O/SRhhjPGcteNCvc30wAuZDnGV9P8gcRrX8DafgSpmx
8GyRm9bp7y5zyBk6/rkwO7YVhTdBidm/NeW4FpGsbNOkwzk1Daz+qqqiL8zEz4G4
9xxWqwmQ6mNL6Fj9M/PdcZgqFEJ1w7pbhRH4oOeLmisSYax4P5MLWdvqJGMe2ce2
ha7LqMoXYnGf6+2WK+EBZb5fD1/vo74nAyCSNehPAg2JJgIU0IXsA1ktwWNCOfFz
kjLCBj1dE+CpRM7RPztXCmzstmeki1gaD1OXLA04NcNbEmrurJl2+lXi7coEE+HP
dSMBd9PK2mNDeFIYsHBblRD0lMVmprmOcwJ0eeyDGy69Kr90+gHB1b52987wGzei
ovctzWj8NnqWcP7bHAib8PCGW/JNdtRZWeaIv/IhIc1As3ErCyP5lEBGeuk1fGfQ
RELGD5MeNu5Mb6atucffoseAGtgeSJ22GplAoV29waT3+vk5HKg/pcGC0byS3rWm
ha/MAY2rt4yDM5OOLTNurl3DCfbVtw54s6jNaEZ64gp18euHkvOXC0hK+UUJlxbK
nyV3y4X/ezxB7g7yb8qVOxd0iurgQbhyt4sofKuOfk9UlCoIHlbAVZ8+9bOmQ82q
xe98OKVLmnlw36XSER7/kZz13i+sMfentqjvPQ67XyEtZJRKYeHc2lr11t3a7waK
Ea9BX2pHBFc485X/hgVDEWa9PfJHb2sEgOhgM9fsOCicJzHxrVpd48FFB6kvXuSI
ow1jK4Gd4bezOryrRoBrkCNFCWCBw9Y96Wb+3K4DP9XNPuJtfWS3LTHmR3N6o933
bOqOO3/ZsLPQE+G3tQX6LrLq5l8cBP6m20T+tQD6KGCEHmqUsLOdhQMUoxv0Z3IF
tRlpOBr1lN+5Ak+Ate/4Qe7Yp9HoJLJ3RvsOuUsaWnS4c4UH2gyXRIvMXFEEv+va
9A15UZcbybKQqH3tUkvu4k5Q4jHQBSgFCPQwvV4zZDWK8LwXIJCdtYJSmYTHBnyB
qg39vfB68gMKq+eNBvkKXgMce++Jstz95MGUfw6KWaKh4mrB+CrVdMD+O9JYPanm
FlF/5j5EN0Wk+iWwJ1IwJ6nBMRMInjQ5yZEvBAzIC49V3d90bMn7w7X7OJ7FueNe
TP42+eBKfVREw7R5dOMKeQvZWHkhSxeS4G45U3R4G0NQ6TN6iGsU6hfCZ971RWFl
jpfHfsJDVGT0WGFhITWbXYlpdb+G4MisOizTo6A8jaHqYRqm2xMZisaACKDaoHFl
FyUs5+koOVkPhOp+HuXPcnygJsx0RBzcDnnJwP6HEbCGR5f/6v508aZoC6RvNWDe
bq2ejcDvarKWJGkUuClFlz3nUHBVWm40O0912xQ8PFmt3LLwKYt+umkg0olMVmCa
J6WvnX7HqyA3nWQTpL5dqnJKMg337cChsFlNE91yJPWJWwEDxMz43LlQJ6l7nn/u
IW2h/S+FNIqckCY3P+WV/ZZuxwp1weRGxt9yPSXo8hne4aMkJRsrP/5qIm9z9MC3
0XAeSPPY5FqSdVzRR19qJ9B73cPB9tqdKiYP2mi10KR/7iyXjdxGP0iZHCYIiBPy
dcA1YUNtqys9ENzplU5c6YxkISKr9OUO5AH531SqRHQHDreotlQiV/a+Gb4Kn7Lz
J6UghpWszo56W9cPFgBccXWW0VxaeXNz8zWglW244+35Ji5k0eiLnOjdJeYNiWtb
d1HlA3+SxFVTWE3Oheq/tQw56roVyX5UY0fJEzj+V+CGfQ+HRmRBXBI0gu2QW7SP
TrFeWuHac0MLqS3QIIkFJiir4vvjhvHKHAN5lJvOrhYB3inZma69yYUQoYCZ2spL
Zs3JN4RadgrD9tv9hDLf0M6xQwE6Rh5ILtFGgaDtFpsaoqamEV7vB+i+BTt8GYB7
JSatodKWb+ss8+s6FtPeSQCm8JLBe/aSqpfhb5lttsW6mKjnh6TwXKwz4Zd+qCQR
Fni4pD4pTVJkRkgdZPJSyLerEjoU+9bL6gRh/ft2vxQ1Xpusj+IgC2Vu10N896Ku
4af+C4AZJupohUEHGucuip3Vkubcmt3HbGq/nh1c7xQ2bhexX5byXUUGK6IacBIZ
4AkPHerDD0S4RQa1mzkcTZMUw6OUuMAgPlcgJuQRmi+1f6u7IsSttAGwLL8gDO9y
PG8c7Sa/8BLLuurjxZv8tIBlsBzPVSCrstpHXAf9lKJigGhF92iwWo497sqRyflJ
3RLouKRO/SMM+SFcS77APebxVxBSBgTCdk2a7/yVIQFDEfsjNTvbKe2NELUIDfBV
og32m09vu0h3E5CCGFiU3smCV2Yo3jzmzB1tXPjbvU1LJ7+sDyNphX3/XPK/S0x8
f1zJ7SHTlJQfM4JBc+o59uRAnQHcL90lxdZJSLm2mGEDLAKL4KR712FsoOedrk69
Q2alFvQ+NIfVMMCZGbgY+phmr7MDUz2/a3iwVP0b99Il3+Z/v37kkM2ACH78umHX
bIcaSDVvINNs/6bbm8oE098cAv9iq52w6nSTzsTZZFkcXH/V21/FnhhE6dOfokeU
NxX6slqts5ijzr436l0eVCXR+rqqkZbZx+LONTe0xHSp5xGODEwhmRej09/lN511
xciw57HC3jGUrvZISMhecK8m13AUZ32VrWrTOWt9J9zH1cvCOtgf7kiy/rUZQuNF
jZGfZ9b+OC1rrG2hG3t21DSmK/rCz5WvL7fl8efc1oUOmVbd1EkPwIV6hprIv4y4
6D3E70cXjpYLyhe5FnmljiFXFbuuwG8V6K9UKeQipSXTKNuFcEvOHPy8XNtedJ1c
4GG6UJmi2FgdQFUpb6Y3cGVQEKZ0Ro0YXYjak2laRzznDoCJ99p2YFWemfQemMHS
2SwfFefJ1eR6pXYkZ5EAWFfmXDGqVNE2GBB6ZPpUvTCLDetkgWNs5CjsRa0wQUKm
YS00zevr7uAq+zxQt1G9xtWjf+1PUIkuDOqsnMtm9uXffMCgXWuRG+iwF4ENe66T
1UBM1GInjT0aVisjRYkDYOV9Cvgf1RKmDcYCDxzPVo4NrEId9YiZmGPeW4EfgN92
d1mm2zVQpGQGSix/bddKb1m1IkapEPESsi2ZLqVcTqRHboQsYvg3U4+1DRKXEzvl
yJJyNoseh1oq+n0dXTREuggWX5o/yTXz2931+kvdJR16spNQMPmKIzTyAjS8gvFY
6/Xr11CYO6Fid9h6DInp8n42tIqWUEMNEMUvOkulCLJKTNSdNtj1k/aHVT+JGWUP
MCQZpD+bSwGIDqnprRkhkzotEDouwX17ahtVPanaNgVY2lUW/NspGww+sBy/zA/n
hy2cztceSS9zXkTuirvmfK/Xb3vL2K4NRY17BOvgQVjyOxcx8RMlSZOqnAIEF0IJ
bz0GSMsO75lVmlcdHiKrnSxXeWIP3BLsJ7H2Mg3dWIm7o/DymrN+fv985uSD/dsb
2Df+2cM/8jzNE1HkBmjuyzwnIm3/NEfYCh5OsE+sygC4kglmQ5bgv+RJ+7rlQREl
Sboo8jTd9F/bdnsfykifGjJbbTgVwxyB1KG6LM9+u0f+LW1c3lKEN3ytmkO1o7cV
tQFjrx0DdzFgSFQOUq/Ipie6XiwUgGSWOdKRCiT+zZ1egkzc1Eyb/upfrEroNiQ8
zdq2lZXebXr4WBoImJnUwRfjUj2CtL4kzXrY1fLIW41nBXzRTnU31kaNlDI1nBvz
54rZnHLkLc0WCBnXEMgTfOPux1NLB8NIijJwtJU43P11/HvGMYqzHi+52vBmwbt3
KndHZ6mWBZr5jKRh60fXWdYL7y7ZGdr/Or+LdQFE6xQ7/pqSF9mHEPl4ZD582S5X
xxnwbMqTFPGPwq5M0xiYj5XcUhzc2/P+F3sj7rxRdfzb5ifRcTXGNW6UQBjeaDfJ
FPhqB2wGWNUf3HbvVRU+INKBRRt0x4HWlzCP7LRRIjITykMsQs/r9RE39PMVL3w3
+jryV3tHdBMFMo0VXSE1wa4yA2secVeoUsW39trSXTSaWjvMESrbinsd+GMk5YdT
dSBJsgyjqf3eXp2nCHarFl+ZDd1tssj0daGTJmKrmZVRBFrRqxgJEU93/YUhA7bl
H3X7Iiq/e5w0Nwx+ysjv058I1q6MwJ/fGd3acBf4lScotJTKBe6jSLmNn9nMLygr
0ouVmFuNQiNKmAlsRUFqf7nDHH74KylOyhEwYc4UTzfIO1GOEKiAYddvG+5cMu2c
0lbhz/jSVNqsATlsv7Wl3uZfKBI5jr8MoDYSIeAkFyzjKXTXkicJs3kA5QZl5mPE
P1xF3KFTe8itUa/UIuNblQB301u9AX6qv8LBTTpQ7CY34trMfZK1JkJRGjWsvrFA
/uvqHrtKD71XIvHO5hrpx5HL9zsjmwV27kFBgaNu0VjEY8DyrAusKIrfpcSxZWYR
1rdhfT8GRz/NAIFOujY3BDANZYCIqPAR3v2+QezymiJG46hyrxb7SW//yIei4YGi
pXSEWc/Cx5TsA3aL1AzkH0tYSpO34ehclXcaaM+V62rqybWR2CJFjhexaKDRWOJJ
IxEvB1V6sMhFDrt70hx9BQfOOr/iZS0on7yNEG1rd8jdvUqsh0U3JGg5uhqaTN/A
v6nqouP+Z1Ffc088FxRYXGjFao6g/F6n+ST6oGA2juYPWRnCaP7WICq6ulk19FZy
0SNOF2QFzR//oXm64Vffh2qM4BzL3ZtDwhe6B25gJRBQ8p+CcHeCKZo3XhNBJwmM
j90DTt5ygZNoKzkuLw8c1exdyEAM/h6K1jE1cp52T8QEiqbE6lHKkN8x6Lex4Rtb
rMrg0SY76bxcNzmAqABn4fy7QDABjCfhRF6yss4cmTnv0G6QLtfj6SBR9ezu5rm+
XjkrJ1+4IesaHCDt7FRxeprpJVlRy4PGcRuiIwQ+RBr6whaNZdGoOCU2t0D3IdNY
c5FrSKa+66uqDbSGa/i8AxVd+G2laov9qKRHClAiADSwXslsFmXbaLRTagH7yYf9
GKv2byKK6NtkSiigXPA3+H0IAtDEou7P/Zur7I5fh1FruK8/4eMVcbr9oiQIMnMH
JtFt49HDG58sygEdQ+6NpFD4kZNYS/AxmBrfm7dykdo6GcorBOq+WTvNRwz/GFwM
vIIFKoxACodrY9d1sRLlK8OYxXeYuTWJCXDkHFjaQf1oXewP1EzY0Kx4ypFGE/0c
1G8x2win6NT2XAZF+/QVBJvlzTJ1BE4R8t8WQzSVHnQfOHF4RZ7JeSlP/BiuLcEj
NPJEjMfUxODmDV0zTxvZmL50VjRRcggNrEb3eJYO7DxcouL7Mvnl8ljUtabSx+yL
u/wB2vcBAUMTamMcfty4b+mqshf6TQYI+zKEsbmfQcELqu5rT5HLHtMoI1mbJjOz
0ZfeybuOHBZ8uHV+1uFXBQtwAWGQSV1Nu3MRX1ykt2nnI+Osh72QeQeSmfkZKBln
zrGmanz03m2G16ClW8CN/d6PduhDW0QQS2xD1kdeIgbtM9oduiKIroAM5B9Lwas8
3L/YnzXvkDj6osb/a/++B1czJtQwNiDF0YwlQTPZfc7muPyecV82EzVCrP15xbab
XhUOyLUBdILIACBqlGncGxexh5BkTidrDGiCanCjPzMr8WdRV1VTG3Hbisc2IzVU
UV3zC75Kl4ptnARpRAi+nRQvYhdhUoOhpYztHgUG4xbsulSh5tQ2R2kAkFrGm1gt
o11vqDBvuyvhjvZl+nhU+ls99Y6rP+Rc5+/qjWdgHHo6OOoGFZSNvT52i93Rktiz
3C6gha3defN+CdH5e/wT38tro9Qo47TGbT6fTnEKWTcEjpfXq9w6EkfpX+wIQxQg
kEBzTo4gHPQsP8YZa1p572vsaKmL8HEEGPEt9lQ71nkzJYOU3Vop7EjEDDWWDzH8
z3+dEa4+budHaU2fteG8oGg6Epz9guLkhFHcz2i3Z7lEgxtABU0a4FkzWHDMXE5p
rmfkNRIiJ0o0mhfiH7VoXKO7BIhsK3KeX2kikKuJDKMquFZZpG/bmsc2Yy7+JEKW
IbofbES4ccBuWw0MVeBL5wUpnHdmUlJMYZGAEzaxmk7YYV2IiiHcHosedOqWRLDG
9FRyVzco58YG69MnpdOxaqkT8wwWMv5SUl0mpZGea7IEaIPk4xMf80bn4G6YAe+C
b7nWLDcBIZao8NeB+RTTaDQSHIghup+R/S1HKshDjwJ7QacF7OzqDrtIsQnVsW1a
g01nwzH1aTrFKtmmKAIDrPjqOeVTit35fL4r/c1dY+mGvKjv/X077HgblzbPpEqy
ftxwcAm0XtRvMEMywuY3WZ9VYNGnhZ2u00IUANu1tBDwLp/jjPMSx1MDHRbXyMeJ
UYtn0Db/Xj/3k02ORYwhUEZYDjQPkHOaNgSIwuea7H0GVOVpvQn+iI1v6dJey8QF
Qc0ZspDzng5qTKLxqQGKDjPOV6yPYJoY54FCBBiKxnLL+Lwqyhr2GQuiS2askimh
yPKcaUeZR4LlWP9CvyBj7Zn+qvX2iIg4VFZ+ieOQmwmzPSIXV2NYaJx0xbSZdrcg
TAPANJpplWvAMQjP1IqbSWlcPml6AFcEbzJaITRLriYgoFwAf4JRpi/8Cl4AUlHD
7QVMohKvvJacXMBhXRna3Ao5m1RR43GOfM/DDDh/691sVvDBpyDjol3GyJxDywbk
qoy9Snv0yQMnU0VsaTsMoR/vlJC4GrnhOk0Kn9/EjAZszy6mwvveJuX4gjCeK7Gd
1n9xvzLKCb1BIPbWQfRMVj9G3xT83G34XJ2pq+IPOWR6Mj/GjIH6016txaMPqi8x
uAlZGlhzknN7Q4RbkGrsfk72DDkxHggoSdMaIvv09EInln36wETYgKiNWMcWwpqR
tzwmdGdMa33BJpNivaF1rpIiMpib1WdDa5Pkxa5/S74tnUoCGjt30My9UG0dNl1k
wB6U+aDtICrXAIVlOMDu7ACNKR/4nRLXXdFPerfqAyEX1BITvrNEE/nt2p2ej+eW
xHHLq8tb21LIu+y5PoGK6D8FeyID2nUBvuzYZljYabQzGhM1NU0EH8ijf0063Mbm
SdbN47+gxvHEF5U3kfIC5uSsm4lTltws/encuoQqPKItF/SI7TkGmi+39bEh2xS3
G0K71AE4eKeJy5M6PVDbalVAIgTnNY3mbS3baFdRzH3CM2r6pqS+VOQkuGbU9AE2
kIWzELBqSeaW5t3SnipUIXAZkJt4Ozlbl9Cq/8Jcf2RrZTxUotWwa5LJNOy71ohF
XsSoE8W8E8umXOQ6/Qu+FX8rI99HrX5xvbrorS9435mRdXz4vIPGJABPHHyNnwuz
rCapdd4WjnsUTdhuH/O4zwBRPzf4xmRgipaT88IGIMyjq2pP4jh69wJ+Ke08faIX
ZiLBSpMVfTEajLzEJTE+cx1pFu+5aaiv7ILyI9i1Yt3o29xD3mOx1/JItTEO+44I
JZ2hVn+989OltirimOWBDKBpGTR3ADWH/jHkcojOKGwbMxow9n91rMUvn/oGAWZk
FWG7jxILjBa/kwdsS6+NGsc9AoX1WotyScb72FjOjOTpRuk/mzWlGjL3z2VSiaNV
qINmRGk9vV9WBOp3TTGPebl56Ho+2N/MyVJjdQap5zzRvtV3yJte54BYGE/KrpNn
m5nOkY9c/HTfQ6wbDD89wHyLKzqAW449xfS1nJn/IscdefKJYyCe6eYnrI4TVCA3
m38Jo1ykO66a4cHqNH1Esj5UQbpQ0qEoF2rJxqhT23qw8gBnSkavlhaa4xAAqxxx
cFDPAjLudz5b4UsTPN0bGCEkEh1buZSUZgYCs86BbkxE7zVJivhq7xDCZxoGfWwR
Y+U0lLEUDhNzzOwHVQCayhCFVL5LrR4HZEiORG2fwa0FpvwFLhp3/zYKcS6s4nsn
cS1UfSxW9VUrZr2OJFUIYEauw+Tmzkr43hPcbUIu2OHu21xlQyGZ72SQ2JsTh2bE
2zxS7KJJZXeMAiuIuwHvMbh8EbFOkArVOsI7+YDPHgbIp+diEllTPkkWxqbkdrlx
5LUokVkagdDqXfcaotXX8VgjN+c6qSUF8mWnV9Pd5zrWOp0PckwM2jQz/oJOXaEO
Vff1JIIazu5PyM/MP7fCc6hscEV9ejo93YY2Nqjj3e3L8F4YVazUAeOjgoLRzrPk
XcpsZveIIG7eXyTy0xPmjcL35GnrbAtb7Zp4N8GoWJPzilpWYETuUzkcsyo+d1eR
nxo5kK78Lp/qAAZ/IKG63fZCKBMceVuruvenrAQm252DFd3gE/lQTPQEa39LSv4O
XNwXuQJboUXEkGvD+I8b12Hnk7bZlHsZC89XsTHnzGVeSKUljOOOw8pIBQ9okFPM
MyJJTZtr9/312K7Q3/o5VnTYWQrtWTPIdFp3u1yHQVdz2CHobFr6Yirv9ZM92bCK
3hRjYBV+PpYBNe3qCTrpCEd0cmbvaPhuX8jMyUMG9hyMFBikqfL+bNewHqFCeqyI
8kcFVsQgkKFdNt5acQo2YlqkUtJ/is0W5TOaw7A+0glmdElZ9qjsiYjjxR/vQBp4
FJ5rvqjMxcEr1tRuEi4Hz74hXWKE3Xn3KXsRaL3048adEftDVwmt+uHxJbaYnwZL
AAvJvpEOISUvHMz2PD2BkCWh5ysA2umSJ3kuOv4LZDLLTyUrnJA0So9grE/ygNG9
vzk6w7VfxM+mxtfzYEDDuOdvCWcyCjbWnYpjcCKKTXqm1PZKsUaOayqE3K78iJev
XsVjnJ2HpIi/7XU1vKO921oquN8jIUtigUJxFh0IkCFkrbaVYzrX0fBK+egvYj+a
uloe7kztJzkaslbyMLHpJSlxncK5kber0YvqFnVsIlg/lBEu95bgrM/Mqo1owNbQ
aAjMPHwmnGQIGyztypFg0uEv25IaeXU1olUQeVgKkP2mw7iUokImGCmpLF8Bhn2M
04Vh/F/GPU6FDXq1LQQZ+MF+ZAEvKd813zd/ehL9hY00GBwVacCGqPiip/eA94Iz
7RoHKFIlWQ4/MJ6Q0d7UqdTo9Gd+UGtEqrv8/OSyAR5P8q4q0w1SfGBTmE121MEi
feFMXi0P+REIs1FSg3GsaVffMtdzPHlhw9SuOwdmNyYq/VjixTrSmMmkZoCFJ5Su
vyG2G3NmC3XFG6uvszCMUVL8assce4cW1zY0QgFIzwVoaujZAjEUlgrPjAs3l96I
4r93F4ZxIf4D+XNrVyC4RqY/X11OGMiPnfndTkdYGjFezq5VPozq5ISJJJyPn4Qb
5HpxW2bVNEQ73zIIVxZqJXxONbiFtH/6tcGEcb68xuro34ELHA6lytDx//1TF8ul
l5ef3RoNJDoWgNy4cTGhac4SIfkFEXVpwHg/JkF/nM8etstQ2GOqnyXIKDnxUEPY
WSz+ZDxFW8Xghdl5u8dpGooONpsLDpmY17aO2UXAVaFhQMekVrMY46wPqLXTHelD
MYtbszgiytLDsBJjKqwHjeoKSnBrLm1KMh4bOR+aadE4tEhuOkWGTZ8Wiq5YNwgd
fgPpgYHHwy2/WDWVuLMBWqli4nL+mLIecNCVgHn9mz+jR/NaWxZ+mTMhVtnL0LFZ
GET8mm8Q+D3g76EP49rRSvBii7xcyv9Dh/yjd89VE4MIYpMQ29dy8MELKevMbhVE
FjzWolKu7pcS2T//EGkET8olxysymjyeWtt4oCXOtsj9G5MxL01Ux9nD52cBGkBl
Ws33ok08piKw2a+SUKerTOSNydXc3iGWxlLu0hjLRZ+Z8q8zEcYVG5LaY0zhtPP8
dDRO+CfU8bmcsfq8ZfeLkEQZNcIaS6qUiWEhLixCJTDlYLNlk+B2FuA6ujRl16kc
etkYNkM87amoMIrRs5ld5XVZWENs2aQcSQYDaRQ0PF7E8YLNZAlgazbSkP+722X2
hUxfF8YZHdM7aFkw1SWJMPD03ZSxANtTQXXIeNSL8RXmSiAC1QDiB0itqd7wEHVy
hdLjzR5QaB5+RBrx7uonRKx0Fwfxc6UZF5u4Qy/e8DXPEeMopSXzma3cvpnWQaSo
DIdoDfCQdGc0uVre1iCsgtoB7DlzbCxyCiJijvxTQijGqgwVTGf5OAw9io8srdW1
fgZQt8LX5AFTxr3aeF+lzFFmZw44DCafHJMLqtvHIgIWr00IjeNwkDN9haXWDu/V
H5pPg6dVmMjFdqR4ZtsVD1EP6VBENQLN3W8Awd7rDtb1wgEKmf0tQvQpsZXWKgef
iJCxkAUBrz8iDBTmfwc9COxF+uXcdr8VWKGKkEhp9ZKKXd5QoIhlB3oYvyTUXoUJ
ABr7Fb4nPMcoR6R7DU71JtSC+w3g4dwKB+jcLRkvMghd64E5IzJW0QblVz3EI+Xx
m1AV4oAcil8vZXcIhj+0r2oaqfl8pXm5h5ZOQLMoDA7jJkE9irhGG5t9ZEzNqwTI
GktisDnvZ7BiHh8Hjd1ywP2za8E5RVi8/rY1gMHCMnJIdfSbSClWaUa8UUoFw6o7
vLvyv7D/LDYF7epb3W9u/tssFi4QLObl5wI+k2C3s4/XuLbkAndV/EjHQvPF7gjk
0WrU5quotqh5oRrahOn95quQXkaTJrGn0SI7H5wWgm4olZGeekjfrfwGeeJcK5PX
7qWQ4jqWRb8Rs45OiGdqfdbejGwugwsi/gRIzWnKOq5MAhPSDAj8s5TN/qGWYYQN
+YBsXE5fpL86ZB+iSINXf/Ny2DPWv6iEFrrmMkHou1Ck3422tOEGTMg5EyOGKUeJ
Mfwm/RtXA8h/juvsTdVEWRDjaOJAUGb2ztzIWHXEKIbFGoID3gGqqapFJF4ElWIc
u3jNYC/UhRYszDjOSZS+8ByrSNAwYCq+dGRJPLG4+MZ2+6mn1xWCohwghXiwUnw0
PxJIwu5+fUih2rJYyvmcHpKZKbTDt4egVn/PdmeQ+EBU1aCJD8TFLfW5sw3885gp
NSsuUjq4RgRs3r8JKSzqjZ72yPGKr3kcwo/9U0oMb9abnIOLI3xyrUl0vwJuUTzk
JO9w6Iumr7RQ57r2BNh6heXBf4qKardh90H35eZcTC11Yk2dz+zTQJz0A9MMoQCq
JlybBjlpgMtbGwWOJJ1E+beLGmSXH28MX+SqtEpLiv6UePp9re8kBf2ahkFuacs2
jrg7G1uSRBd2kPLBP7BHXa/QOCug+FSqSNQFNEh2xu2g1oAGU9HfrLsZUxM9JDUP
lHie9SZq8JcX7dkxuP3FICY8rdi5N/nsAy6AIUMdsxcLItJtPmKas2vWm40wPH6D
uNlTKeW7b1aSblSHPEinrrch4dMTkeGznfekiD7BzJhYh6+RfZOH69Teq6xOH8I+
ZZ8qQgZ+P2s0ICjr3GTHxDiyudC3qIQ6HUTU7lsOyZKm0NXWsr+JVsjUWEY+Dv+e
OkxiOqlviVUjKEw+kMmZc5/opAoq0xj1/V8Hbl5tnbWXEpqPQf4XkJBtophC943L
DFlWK+tJ6DV0gq7bamnKy6MAH7Ky69xCzyRqo0zKNSY0gFia2atwxMkV0asr/PIZ
oY69c98x7GBL32ySIPESFeSiQC1IWxrzlE09C1ovGxqmcJ5EqHK4OPPhtIlg8TjB
gWzaJB279Uzee1LJb+MwEYyeNAZDIoR0QtFH7aD0xHawKD+cPkQWXq9TLbd8BFg3
KUR5vTygjzWFAkjdRnwAkSwwHm7RDhK1YwuoYFFlsOq8r3gG/rGv4f13fnUF6f9V
JjbGubKRBdUHLdVANRdVpedUFVi0Bhh9/QF1p1Yf/+Cl425IQQthWOYQVmXFJJDQ
VgClLUZyz49D2YwkfsAxP0jRCnhfEaHWXfZbfbllJx2suGWish5poskedtKoy1nd
LnVDH8KknTrRjHSKZkQl+nBmT6ottggpG7ZY5z2/AepVpsA4qCDWeh2abvgJ9Is4
FlX97p/igJSVj+hcrsXsSAV0HRoc8MOnCHtrHDnlXyKagHi9EHcQx9l5cl7xp36R
UZvk2KiHMtRWe2NdJ0YU5aIa2oF3gU4F6N3eiRW7BONnpQLFK4Cc+S4bfEhiXTOg
bIZACgSBnyLEhzO/UkklcPpnexE8i2FUeCQKBQWrrk+n5QRpYip0Gje8zcWfIBNQ
jSo0GZ5FS3cM3LhV49ekY3uI8aWAmVdpcPxwcLuBdeUFSyLq9fne8orusnUGtdbL
WBbeGp/CMzwoOUUOZAsOKi0nIzGAATbmpyNYtZFNQnmy0Pr/X9ZnauHgHRUe6F7Z
CXKViktTK3LJDqr9/wE4UKYMASOP3dDNTccVKRjqXz3ksSlgdzlOFtpNll+zgwgK
aW3FHs8aEppGP73UCAH+reGscRheFqdNRNlyvkgOqGWvboAR1OhptFQAmlhSzBGy
S2kUQmCMk67xVl/bW30wEwlwFI4yY3zAWP0amLK2Dl2roDYmdV5eCCOv06G5Xlvc
tjxWGeaQr1OCuIGmGipEoXSsqXg8MuclfY7EU87ksQl8kor2QbA18p+yapo6gOuN
vr4KXsptH4pKpMg+CTrU7y7h/81T3TD4loUy68gioeXsIkZWrQUXtcB/luCZBRsJ
hhJqQaqmXoYLC2N+sMSQ2bfoOZYeMYS5Xc1p7Y5N3/0EH293qcpm0VIEIA0Ts/WK
VJb75U3ZJ4WoXuse/V6wvfMIaw9KdDe8KJjb+TjZEyMb+Orz43VeMj9eAC+YqTty
darR4M8Nc5T8Hou3zaRBvtNlARGtInZ1h8JYypxqduJ2TLR24/9EwBBTrTTSGgY8
Ve5n0AYomH4n73zA99HL9MrOfMHikCzuJUOtpRv1rh5uU0vsqKsMqHcwoXjovF6T
eLQYbE0yZCKNUez93ezW/Lm+8SrNvy6H9p9LE1EbRMGWHBOa0qU9UNTlWR3B+cvs
3D1YGdOAu6QjI4gHM9YFqE6Bh6yQX+uh5EVnJuNqRXYxCZja6QM7ZdiBGb7MtDLM
QeVDvk4u7U7c+3p1H0uwziReo4phFqNpyLt5NYU53pdq34AozY5KREQJvrOKDiaT
99KtfCfKtXm8VRQN2g+dlE4hEOJAyDenbP7RLuenl2tZq3h1CnLTEis6NvgvqISN
UTWqmeNnkca0i/xpygaDFQORQCmoFE+olldU1Ds9AfksL4DBI9u9TvuLrTAeeN2t
JOH08ypymZNq7BBGKdiv+r2fafyV8zPPxxDgaoJEzQU/jvZyoPWRhZ/dhN0cjJQc
TITkDhi6k16tkRFD4Kzq+pchHFJ5igC26Y7YHVU2cKpX4nc3aIfFRyRgk3FdNUh7
VR6Jsgd5YsbZG1nucLEItTJPNbRX6eeADMylvpAix1zlEgnm0FjMgQOVePvHIFXo
joz2ELhVMEgwTVjYkY41xz3ftOENxo8NX5hWBeVUSeyUVy/r4np2Ls7qr1YTcRpN
3jwmgA/XQn6V3o1S8FSkrWLFn5/fXjwqFNHIlBAcYJSjXwQliDuT+G54FCMWcBrV
XLGUbKg9swRFO25bVQP4wDrsqwIONKVBiiWb/VcNW2Rf5hpItAsq+GgzHCC5P+Cq
wIlNifC82LQC3X25uY3TKvLdBsBy5ECvunhfQt/Sc4mKcPksKM8FG2spHpB41ZNw
IMqTCYF/U98oh9LBthfffdHF/1phC1n0xFDHbjG2POwi17aFeEl2u/ooCDMcZvSq
PF/q/jSJwhzpnI3BWsSXt+fjJ7K6aUK8L0fig8KVU2tM1YOW+1X4KqK2inmyZxrV
3oVofGdLH2VCcTG/nK3IjTBADn8Eb6+V6wCJSA24kIUYoTAM1uzPJfB+57VlK8T9
b59OEMDy+d7v9kg1UkuRvG4e1aCokiWBvxghUXZ2+pNzuko0c5HGhti7T2LZuqcu
dgn0GoumWwujK/+tJ5pqZJ86JG/1r4sRnPWh9l+33v4Swigl4TLGnMGjPMsT/BU1
lECHC8+p4vPFnnUc7x22ZevOYxaGyx2Aoc7LSDgXu5iac290Mn37Oq3JSLALSj+m
TTbsN9+tIhWSDzLY/9xa5YtsYDxi8Ce3syB1yRKZlMuybSPZOAFvvNdaSflaWaQk
IucAD5L9ipDD089eW9x3OBNIob6isQsN04sYbOgcy9lhDAeU+IpL7movTSVTdku+
h+cFyZ3A0AbHvHCEHAUh1+bPASNwDMKoK9IfDBFRLt4Qe+HO155RNcVhIFm0PHJW
3nfjvBc9siWGWCnn/lsXHPuzcexVREY5eFofoyi9mIOHpgK8Xe7hnpRv6Q+/3DWx
0Pl/Q9LY+3zQvhve8i8oxZww5BZQBp2tnm+ZHMpSFRrm0tBkAGsjlwovdrl4luzu
WWHJFZAizfPRGtNyhuBehhOrta76RP4M9jo0zOXuGSS3fVOgQtsyn2WRg2fwe1PK
SEkxH2hcERKAgxtDGiIwAOD8b7BBUWWrM1viEOUUrUey7to/9AlMBhM2F5K8u37t
BVP+J94DOeSMdepmKfM1hfSD2JFaAwSRerEQTYvTLwFHAU0EplC+aIvq0wLyXmmU
HzcBC/Jtv0mP3XZTUjsIP0fLRaF2cPqQgychcprt1rHkml3le1FEAkLvkWTdxkAc
RWFHDW1i3B2DVSpRwB2m1jYqf2eMQQNE7D7O4Thr9ijOMNl2ZCTDguoe4YMIEAiP
eNrzEObhJVq+2D01xNgKM2gdHIG8O4+lwGFGlo/XzBhH+POc5T8lrS/1SIehq7T3
GK0+i85BbReo9ue82kpVE4aRHZ72e+S6rLYzcLJ1EWJa1IMTzEH2bTHwznXwmQlA
wzry97t9MuHsKOth6gRrU3TaABz4Ko3j+CZQRzI0O4EPj/ZyPWOdIcBrJICRZPJZ
/Ui6MjtAKbx2moNSZfDWkrYIbOtE+PrWgGCrUDvnoVjc+s1255tnphqRXoSNZshG
w0Mr4ETkiFlCvTutxAAV5zdsw8SZXUUWHVieoS404cjIRUAfn1Z0rBymcB2Uhikx
L+DzzFWAKymLaeIx4BMn9m8NDuyqfxj/bpek4S1vMikqE0S+tA9E1tNZsVdxchF3
f7o49ybKyE5jsLMUN53W0wINNRfccBKADd9Mk7li1j7caSk6FpU8p+ROf7fljhFn
NN9x52RRcVDVY5WXEYDyJ0qF9I8tLc5c0ruesT+qwHj2kJfShn5TIGUkMKsOU3cA
7tzEhku1Fbib9ShifaOahfCjkCrAZPsNbd749U92lNMP1uAuHyfyt5Q9Dr2GVY3T
mTOVnh8FqvT4PTQLYcm7rg5kKILDEoxSdWXRuZI0sOZkf+YXn0EVX2c+UcQH4CJX
7oOcTUhlccXhSrLiCDAiFkTZInlrJZEVDRKjgkfSdikA7AbgIxdyS39eyHErppZF
d87AY7+hj7iynJJcrN9r2XG/trENH9dtBzDAVPugsRsKFcGWaxbwiGLINTPhAWdV
2fWaIh7KErTK8kWNta+NYixGW2toQePZ/B1vB2aMl1JUZRH1uleBijc1mCJXDyw+
onb1c9BTlYG5bIUVjiPW6dPOkO2OD4tyigqr5VO/bpKsZe4JY5T/7Fc1lD1IHZO5
pe+OQGc71PKXmdgrymMP71hR1AAu7cUujqjVsegu0VypbcxgOzTPn1V/kj2cDFm5
8qLMECslpgy3PzkfB6bwp8NCxmlfhKjumV1XymWHp+iIRJTHuCud0vNPcv/U0EVF
M8gPr1im6jS27cLLWdLuAFVMZ+1V+U0M2iWAkr21wKDOD3CbpXdyS7DKZpFhGET9
pzYh2TyDFGDaNQ447dwkLPA6dmj88YlV7a7b7APnJRafwaMogd+Mz3Q8WfJrm/bl
b3jMoDezqvzt7AokFAmAB7VgUUuYdiZa41KUJQzHZfxxEXpz5KHVj7ns3UKUIiyE
lTLdeOXM463bJwZbwYQrTknvw2LhzEVeC4qn+LuZVo0JI7JRD0zZzeYtjlryNaLW
GPmlQ0bbhOx9kSeMMuEXskQsTIP3DIP8zTeckKm/o/Y/eeSpq3lCCWRjdkRSircN
dQ4qbN1sRO515JKQzGCg86c7ECIW38P7YmzheninV/E+Y6tbZFmJv0leZAcFNHTl
XTDqbG+1iz4g/Us7DcKOK3PzrpVngWoHZXVj9BfOyE0Sc1lZftzZraxi8rRT/MK0
VEbjbTBWJyFl8HC0zXlMZpTn1c/uq8VpJlXcLWLUZyzdo+EMH99aoar/2LWAZyqN
EEWkd1sSUNUu+Q/mQBV64g58QsL2PEeLT7jdRQ14iNg67NkQe3Al85RFMspEFRYG
k5W6P1QdxbJk0pAWEvtluOeW8YkSpPnr3fH3dY5HWIXMwT93SmeNashg0Z1iu1mL
Fuy/pmA8gAP04FuajsQq7yU7Dc5d+p2UqtCr0Pst/koAEqAeFfWdngdBTM+hU732
KAM5nFbP7mQUp4Zl4osMbf/Ogb0an7JV9VrqSigPn7P0XaOmlFrAuzaeZAOHU+rA
vogtsuxV3IJ98tVY471JH3zjkPP+F9W2L15cDj9SypmPK+69zYcBNI29Fv0xqyTc
XPUxMpgOktaEVfFpd9oOIL2G/SfiVOOk2vhC1ZkqDfI0oPNSn9iQu1jNqeF5K4Lf
rH2T1dcRtQu4L/Qe/+VyYM8o053Q+ivdPNznaefccFWjuAxMBTNu1WhKraCWVk5w
NwxRYo6OMivSTTxiLeJ8JXe4vl1y2E80yUmiJ3BF1m8xekgIVmETuboORb/hhl6D
rcrJK5cjeZhGx8S1mWGpVuvy/ykx2Qd5g4j/ONX2JnWwbED3ypCOhA1qr9CGstNS
RhaXKeAOoBJyLO9b+INcCEuTV3LdcvyRDC/qTvrWLXwiBbiY3XzARG90p7WAXjcu
ELt9QhzWXRKdMqpgXsu3gDbzN2OpqyvVvrFrH04PFlxJDOD15XmG1/UcVbwurVt0
kSWt2TNpfawG3PrCiX+9VYkCkndwgH38Nv4AKtmB9Ayw7064rSaDC+IsMzcj9t1/
cWI7cYctrjT2mp0SPU3khM75R+6MR+FfgG8dVq4Gm40vQobiYTWez5/Cns0J3yCO
AhNLdYzRkNl1jXEd+sAIbLqFhakHhr6hlBcD+vID4ojqXhjuCuWRUkQD3tz6SsOI
hStVK1g4SKr2N9oW2YUTcMfdkzA34n4Z8wKjclsG8u3qx0wVWD/UUJHC1ga7wVcN
kp1z2FyVg2M+4p+ORe9eIQWcFnNHltTFIespbc57Ph5V9vTAj2K0vrGKTjxPCO4q
2bgxXtvJ65XWdAqlEdB54Y27MG24p/aDLjR0/E8rtr7ZJQa7rW98i/1YgbmR1yLC
hhTV2Y1oc8hFR5qzUJdfFtpUY/Ys0F8wN6cFbaOgFx+oHMlwNPeclQuKRTJSSkAb
vicl9s6DgZuge5cm+vDGgNLW9k7nDMDDbbv4k4joHtq/5QBcU1nAjxws4WLQTOGI
Y4WOV0mHGA14h4XjRvFOVFdQ8WWKxvr7xdWaOFjlOorJ7NacDbk9FgIO2KmudMpE
wm9oq8VMCeIhy+1KSLyhjbkd5A9vd6HD+HiYHc6XvJ1TSw+XDHGMhJv9qPUq/2Vc
DtYh/fQf8Xdx9Gsn9FxOIUd+LrJSclI6n7hiyk1DSU08UNyfB+Dv3jTpGk2VTzmJ
Gg5CU88uHERdAZNyReJgUPZJinDjw4fVw6Bx0nn5fbTmMEQWBd3tS5f41A1p3d6A
vdk/cWzcaWa6ZB+LLSLg+IJoC/ivGCibESrSn8H8zX/LurhASZHo1xdjTH9KCRqH
Zw6g+MzW/UcPOuchS1E73Hp/NZsTD1QCWSDdeqAoferT5w11F+CcQ3ZAJ2gqBAEA
/s83VL4sH4QIeQLeQP9GwhkudHy8n9tl4FES3aivDOPYqmbW+UfT2Df6SnfVvUov
rGafE8mSQSfwPF7Xf+0JizEW71dZL6pqJRvjCyVgO/GHLZ3LEnTvIBUlmDHTDaCl
toXmgmw0BQDLE3XsPcGbQJPmH+4ysNxXB/ko0kcdcwOYDW/UuJMTI6UqQ67ASbCw
ptfl3dZR5qm0z1772nYQ20QjLfxqgfPmZ6FB6AU8OcBaUADEyCIRQ3InXoprYUAj
6l7z/BZJMCRFfixIDXXkAKT/OomOHHdqBDoLjToqgHhDdVFJ/XE5f7GHUPQBXqY2
9Q2IZVlrBQeixvbTIvhEmqd2eLxO81cr8wtCJK17BWMLAaD1j3J05LxS/g0lNQv3
rRi7Ff8CbANUWN6eLjMKFxOCHsCp3k2EXjbwbXAETipRWoAjvNIYNprKJorbSCk7
1hI7MQANkhKpOuXMvB3t9VKs8vpEEfQ0ahinJ8Jim11NeejH2sL5WfXdWT6RaMPL
TbDu/0p/WQj2G1lk98Z86PWs4Zw/dV3u4hVDmtIdymDik2kqUmUl8lu8q9APhVOc
QBpLV7Lg86fxxU52SPBvhNyyoGHLwByMcFvqkziGPGgE0Ukcqrh93qu8L5h8zcJ3
3WmqveA1tBp0M3rZGYSv4SfH08wLgNnLMKhwDPchVM3O9Ce6cyZIzkPGZi9OpUjr
GCgAHaS72z01XPGvhlp4lVSdhv2H6oJcnMJQO/s/xyTQ29od0sO2151ABfha+DVa
IFOzA4fdOaksBrYXVswj0/C85O0GABWO7lJ1JYC0is4iMlzuqlANuBP0U5AFkvpZ
lmk3COFlAeGU2k6cBFEy+SXP4sfIv86d8tprjrkSiJDgWsDzo4qadT7txdn0SP5u
L+7vyFrYjj4ufQVTnrczLhE4RuD7tUgl2PQqWu+bjKXY60x7/ytFhlK8xGDEH5jh
TD+ijHO1wB5gOiMLaWSb6oQVyy1h7wwV+rzcAWrHb4jBUMUb7KMr+H1G6ZasJOY8
tsQg30APu6GvSVcLPP+tN+vJJVY2SCs/hknBDjL3LTP096z/ZkgJFJauMYEP7m/o
DAv8elRUQg6eLEUO3w8GvwrOxKBZtFAVJBsRN8Pe8DkQjbp8f2NOquIfXDgJgi7A
yDrSMQr0as8/dYFgbp/V25cpAp6B/WnVcRPcUV2kF+srIWguUqw1USMs3vNvETSJ
sStayOZfNHZihoueI4rDv8KQuAo7HNTaxXZl2L0i30jG/dLHnrmUb7Rm85LNiPQi
iiFVVWBEsnEVlhU7eDpSJZAsysddp4xWW8lWGAZ9Yvo7KqazkfiI0Yfd/L20Yg+b
QBsgwOaRxop8X7LCcfGMjG3hckCQtp+l2gqQSBsOeFMKrpQ0bo+mcipuQGdtzC5d
1QySl7rn6P85ZNcsvmlLHLfIJO4XVSk6M0yE09geXTUtYVq/R5+5tNKZMcBqMc+h
slpDBk9xA2y3lzV/ejmhhJiAdHqgGzSXBnMS7IDgrHbcUSNFgtIKXHxdDwplwK1k
dx/M0Mma0AazcGREtGE9oOjwOyRUeRuWAtnfCZnkYMpiMQ0VAXB4dpunoqja/+ew
8XSphdRhOanwEMfRsbC3wJxVjC8YFCIFJkcwssY1tru9QD2rb+CGs9UuIUs0ol8j
PSbLqy9U2CADTxJxZmYnW0diaHjOnNJRYjuTye08Jz/h93Ao1z1+4BWZ5v2unmO7
2Bo4q7eUFAPnR7fZ2fMZ5K4YN63cHW+WkQapknVEBqDdkIrN6tCDG0DRx7WVUr0D
OS+x8ledR0JsYfOdeptJa9hRIGShOgdOiClJAANQz8MTCCKbRSxDv8B+F4Qa7g2l
ZXdXYn1sHoPTGdum+f/pcNQkM8KjsvC7BRnMDaAL1BeLz4Xux0MGhOp+ATtR+zVm
N8J6wZQ+9RWXcsZavR7mp/jAxoq0KkHPOzGOLvBzeWs31ODLh8WxjXuh3OYjdDqz
Ex8RJaO3rUXPrvPsTrQLkhEslR3Aaz9HjFfH/Nd8YGgYE/a59b/eUZy4AYuEwAfq
C+J32KlpRuhpGFu6Dy9nizF3XQJbVSGH11soLiEM1RzRjXZ8cDC1cf/bHvro8gkb
tfaqwnG6vNaYybsrJU4dAZdlV+tCAIbt5ULPGSuGKK3fVuX6on3WY8jAJcIjch0p
wUHyZMLQuglUADMuhTgMFuLjrBd5DOBQzgInL5C482TwoZWpauWfu9fhxT7cRMUD
XSx6aXkgnqQroQN9mgRHg1qiah8LRWjashmEW/gK9Wab1raxGQR5/D+Ksu7Bc7Cg
SM59nG8y5UGXbBhvwBEfVKPlrac1mCABezHBJ+qlSqWrVicIfFkkhpyAG/KH87PB
vKOuOfxC5Evjj8lXAkqisc/4gu16JFbhoaO5hc3nM9LpAPTlGhXWN1YR7fIKVKOf
7dQIA9KsTMrQU+5X41KIgWYA+ESsnX5x+bNn/MP2CHMVCXiua2RnbpKoL5AHeIGy
rjyBanOrVbuc6zlHsy/Nq3Pon2wGVi234Mst9itiKSkv8UKIVMvqLAtcFpchrQEu
i+xzXFyyxYtuEXemFI3xyXjv06qkVJYm9A2/mdEctfzV2Nq6YZ+8szQvtKmccC4a
ZwgrO2XI6w+HzskrBQxeIHdIzb/m+S5lzELWyYN2CgCHFiHfCHgEmGw/B1TIX58W
PRutp0AM6HZANlJcMP3xltoiM2X610pU4QapBJhQzjH8Sg5qfGh40+hWA6HKvkRL
7eibfy+IF3CLOVglypMWVJrK44mUFJ5fbbOaNrW5oD3dzdZhxOg1vc71MhhOR/69
BRfZYPiT+fcTB7oeX8AqIWfBw5X5mwvBllNUZtlXhhL81sjtFV7ScOhdHgOY21fP
gFsOsBBkVgtY5Qw+egBbi+2vSA/RcSSlYaMrAVvUIN/qpRqsOX7vTBYdlIeT2itu
Sm2jXeKFt5E0fDB5+U5LcwpEQONv5kqU68ZW39RDL2rz29258QLLJ1uOZvypq1t7
8k5QjBoVIeLy7Mj+SfKSNZC1G6PK438I7LBibzbWbmgmmZkqp49KMABFOROdaxpG
+60kuVjE4C1CiPSsKshTu2E1dUPXV9SviD1Fobrx0hqruLFtKKvEt3iWcMK0g/D1
C4YLl0fDtHKApCyC4VBsbfjKPgpfFNfXA2GrlpgWVLwF78rVHW0crzeuy+PBhun5
zl4hdQy1F+xJ7UdHYrDWlHF/6kiSxOrFL8YiDrv8PtO5P2P++flNS2q+9tpRkc/M
+vaO7ZT3qLmKoXbZTsSQzFx69h/d1FKc6nZz+B+7wNndyBDDvakSXtctfPjwhpNG
UhXAgItMfT+43T47Cm01Il3hT6fIWQZzqztzJzfjam7e4Wr+Qorhz3XerjWxb8ek
oe1Oe8OodyPrb2b+ksYf3WVhHZoJ9Emvfn3Ac39ByNhkgYQOINXP6jSvuet2lG+P
harPDBi2GfThUQP5Xg1pbdonvJ/v6a97t1JDFCNSnN0wAXfQKn7vBgxvwIFCOcfx
NyVAuV4qYAQU8wTGK2xlcPRPeshJnGWvEn+yebkcLYa35ITAJitVF+xOM9rC5Tqf
rtQNwtKn+QeUxvHVfZwdC54w13/0wWKXmC3buchto7wTLGvHLjP5Ih4PFH0E9AdG
eGvvdgE0wf8GIG07hLAzqWoTgJm8gsUWybjU5P206YvFM7SD5Sx3C3LR4lg1dFzF
2HNqobGxF9FHDSNmolqdF1RO24xCohVcWxS3HaevVZH3xo9jXhTJulEjyeKwZhZP
+tC6nAgCdB/f5VzGNi4HQTtUiGWPrsvB9PBKBNSp3NNJD/BQNRFihixG8vBJbeUh
Scy7ABMjXT9GoA5Q2YdGVcu3GTRkn1nhIft7SfjSV0OmCtSHUK0HQLJPb302nj4Q
9EaMouXwGqMaiJxm+C2vGyan39Mpz24gW7c055LMOTpbhHOj5bA1GMF1B+B9pygS
EmyuiXleEx8THLezoK6Sq/M2P2ZdU3No3l67V7gF9CAAo6ghnLq1kWa0W9oPY3yO
N3BrElZs5vn7ArhZ20HXsLs46xUA9XzXp6riKAD1VWHuTy+UdvnZNK9kUXt9bCyI
wHJnB9sWXm/dxy57kSORKmQwFjV8LJ9YR4ckIDZOxIWfyRcuk9mfkkJ74JXnthhw
/D8C00YKe9rcM9tpU1BfSH9ThnkM2bcmCau6pdUNHC3F0KOJuBvVA53iADMXs656
Ecr13bXu1R0mMzIROkRUx6weXsRqIGUWxnoKQts/GLRQ5BKCt8PmaIpQKYcMO7Yy
LUxm3Mm9fio6CCWgniLQe2gpJ5yWGtC9i4XRpFvvGidT1fG+uhWXZj72J2n+kL0h
kOjHuNoOC+gG47zaxAd77ocvCjL1kOJgUCNZg19mPNDusCo+2pc2gBFyEPzdw0Qe
OBs76RYeaoEYmdXP7vRopT4HHs+BaMb8s1Oa+Ed2zgcphzwm8zjQ9YRKvQPNT97Q
eRKwBlae1pskS2FqqIYd0HWYL87jT06QA1pS1oHe/YUaSvCc2d3VETw9jHK7Qz/V
s+Xta1O8rhQTgsQ2CnrhADU8p4JWOGnryU8rIbmMSKw7b3PdGiET9sgRMjjg7Cb8
W6br66xscX8VNCVjuTaw73xsokGRBYXt0kty0Aa65qPQCJ2RJMWTTXeUUDkbjFep
7xfvBGTU33rVA+sPJk1NSaS29F4//Dv1FDe7EFTLc3h3a+WLtniAA0wJoQs7gP3/
HGjp6fmHzwaF2C91ZG0NKhFs3dV709x9iWhQ3ASr4RlN6m3FSq6/61hKTv34kAEt
Xddb1D4P4+/AVPMc+p0JS1XiJqMcX+VFwXzyPBD/KhJq3+Om7lUznXkW2drKVcM1
OVE1YI/EUaERFzIaZlBmHk8v5XaHzQT8w2S2BkE54M9pUeJjWrCs98nHFNgUfHVG
Ifc+Rkfk/qKC2N6LFBJECS932DEwhpmCA6Hl0S/eWQvCe+dI3woUzw/ZUChDQP6b
uGELRBnCZo1Nx43YhCXCglfjXpLZ7CxvyZOqHzFzxyehwEXZ98sU9n5tlx7WbRfo
mfiIRYjBN/DLN0aBwrSl9k8jRcMrVrAWgnVFOSY8zWOtCpT2z0+CcG77Wp6HbPmG
r2SlwkhX0Hx5Xzbb+Wu2PibGXo0Igr6BErVrcEPHqONMmtYMfzO+sAveZtwBSasJ
w9xVAd4ka7JDgp5COjsaQhNjZ31tFdgWGtmtEeA1/M6hcQdNKnLWUuMWVn+4cQfb
o6LTu1mSjLqNkzekqR0m3LSKlOFEC4Ja1fRyUoDQIu+2xG1wByJFbn+miRpiEFh5
Hp4MFPsWAlxgcgyOyP6KMTpRKIn6i7K4PAQIRQjmGxpRL4teEZKuvyGeQ32hJyA5
viWI3sT9QQFvzV0zAis+JLlHQnSc8KRr4FSBxbT0qD3ZXw2QB3cjmOkzHK62UASc
lkiY7fhQpbGTba4Pz7E3jQXh3lo28ozQZi6LCjikT8vuC4nlQaI4cbm24eZ0FGue
aF8nFalFwVl3iBW3aexI4WWcy81qwOKiOOl+goERZk97uQ8EISB4Agae6mQ9YBv9
CZvDI/gT70MSS+BSrQy22Flb45PxwXKmWB5LSjnxQCb9jSc0vDEBXCb/FOxKhYgh
OpWrzh3OjEpDkHj2bEQuyhSpnu3yYAGUKEekRFtKVXua1UQpkRTmxLImNPKdy6zE
43dXIhOUTZ29P6TcbD3pQXa+TFN5cHSoe1WfxAT5IlCXDcFhkWEQZrRU/g3gqHLS
/NdQHXMoH46wG0pMLbP0nRqYTMdDL3x5aWzpeEDsVsAimVt0ASi0LJf3f1c25YZK
URmcGcdIq+mV7LH0xbAjoJp2gk3JcAK1Dg5fYhMrK8q1RiQECx8WEkE+VCD+mD0g
ejebYvkFMdqu4XJ8hUwTiMJ28+SIRX6ashmgIC3ctvqqy0WQp3sLzdNG1gTU14gV
GADIi+47dtNC8unrD6tJll5BzBIcRf285OIut9lprbVmZw/5qBz/3K5A6XzvhwBI
DgE99Hh0sbwCMuQq9d0rx95HsqsSnozfYC4vRRVqxIqMEu0c6WfV1GvejB53xevS
zI8MFsiW0goKzrkLj15iBNTCwYLpCzZl4etpSdz32/m82ZPpoc2OMgUpMqVJDC3D
aMMJ7Usgq887NxmYEtFmRD9noDS8LCnCUCvv9+uG8v5fI9Xbn9+yX5x71RpGUI/k
VMkS2gCaad2iSkHsG0n7qO3hkjSBeiwNfg7PvpHbBQ30FFQLrKlA6239ja83d2Ir
RFd+hB/OzwCIXK9Nb+CDT9Ai+KlUKhNmNPIe0yWo2/AEP02eyBQlFy+xb3T8LYp3
SnMUNJPhsWDxIAwzLWkW9ArvhRdKYJx3YjfJyH93JD66mCuYU7OJjO7TuywvgWzQ
7xtx1sj2M9exoXX//VbHWfdZMLYCeaC9OYZ+8l/p/HmvY0ZnrwLuwVYfWEF73pey
azEB5b0wQeFsXaRBWlMhcmtVZF+wrz4rNba5+qnw8xCzdYwvN89WxRxvKzPjqMV0
5+OJzC+J1oolOKCkR/blbyrjFe6xRLxb1EY0CpOlrOoRDBHWz8/aMRskqAmbywLg
Uqr4LGwpcFQr/0gqQWOkiXx7TSJmrEzQRFz4O1iC/A66uGX/lFRGImgd4h/rzmvF
igjVCuUIeHUtyipnObyK0yQBXFr81AgmjCsbp7dPqDm6Zs83eW87Oip+HuOapIXv
bOu761jwVNar8QM5uDKLkPHPkFUuGgmfuthTmhqiGNrfz/MBwM5bZJobWFJJ8S3V
vgCxUk7CCTkBHxSnilyxxZ+GNma7LArIpFA/75TDaJ4+vLx8XFNs35fmC9uD4zj4
DGgcYXQwM8j66UHoeGsPAjNnGx56FnWeNbjZdk1BYJ8ZhxsHIKiaYMw5C6IYdLY4
Nb74zcT/fPI4gAm0KD3/uie+2UgLYuv7mT7KHOMQ/nE3XEDmQNQgHAcQhgtSphiT
xj6RK+AzescVbYexrXwI7goJkhNRHkMlswOyG06bwUX4mYQ5aoyqZ/NduqrBV0Mt
QAXSOblPtUJjPLQx/CB3yYsAk1ZPAhodaG9lC4sYF8qqh/7Wrgoalf9+8q99wEnQ
Alw2IOiwaiPDsWfKqgjugW39szBSrQnSyJIN7nMBlm4EJZIK5poaKhxVymSWv0MJ
6U8JnyIDDx+0lQLJP375Wc0iQ64RqSk9/BamwQuDH86NgRrgVBECkKwYyd2rfKRL
hnupxvPuHuZ3+C6zXBJUVEZGM7sUaKahRABH+lP7QOdTAhCuRkrgYgq9uS0m2it0
ydiwOldtnANSrh3TDMMPc1uFEase1rn5Buk5bERaQqjw6tFSV7BIVTj0d4l3UNli
YZ0nLzHKFJAWvqsNVuUo3TdH9AI+bSEWVnt+fq4dbiq9oRsqWkXYqROemXYf8KwB
MQjVHwL4FFUACLEDDgowlo2FEbvpW2vNwKRZvJl2ZAVITGtIts2MiV5WERg5vL/s
W+NGhYfVJHwpoqMc0hj8Fkj6I5s03X0KB4lKA9UHA6rkm/JuPs/16JktRETxUfdj
Ze1m2hJf4wpL50B4PBvxN+Q3JdQZLKND3s0PHvEWvam1fhnE+eLEEDZ+ptiR3OZ8
fFjclEjE4uUf9hdyUDfnXy+J0A+/R5FpGzueVMR54bHPP/yVIm5efbieGOZfkTas
kNJgE0MPCQAu0j6R/Jj8h1NHGIBNrmsRnYtGPcHf0RFfECfs5mvl8tBlkJusuCib
6Uh/cSg360st+k17CDl2/8B+1Hda4q7cE3JNOGj9NmR5TEpW21vaQRxkfBrKqTlD
v7NfJSSwXtY8f7U5kLxmmaJPxTxqwCahKGLPfPvvIGt8M8kqrc9LI26iN9iDc30v
GuhUvhnt6pRkZ10gDNdMprekpH1Mh1dN60Klo3GIUa0Hvg4yWY2W+forqwTSmb4n
ddAwojJxfqrvgMXGG7J23cX+ZeMeW5GhBuKTVw46N37T18YXevJgT1/dCcGHb95s
oHAOhrH+oFtu9+TXi/75+XPu7Y/z+pcVreAxeN3PQEqnpHcGUwpj7pMb8/YSaO4k
1HMVz7wTvkFSYPId7k3xMwMVdVRJOOODILf6Y6VmhtEZR61K/qh6BsXFLR66dfqC
KwXhL7tnow723MUDmza+pK4uH83mzYYZFynR4gktqTuEmrrkk43VdhsOmW2LpYcP
J5lobu2HS3Y0eRxf/SvVyoFI6Qx8TQEe6kwl+bM29yjtPKcL00PvOaq3hT1bZUSE
AmUIxtoZg1xYPE3oeziczKHu8WJKXT9O+eBGw59TVi5LSDywRVfRGELlvylxJD7w
iTRI2ALojzdgk6Vxoz4/lMbFPGK9DmZpNCiOCxsznZnE6heOBGJW8WhxFaEu4HW6
Cc3YXXMvXSpSnWW1hSDFysNLiAJTjAyfGFFadrH38Ra+1VEVXBq9b+AnrxGEHkiK
gL2eTEcN1EKtQcBay+TMocJn/zcnLWs9EFWFMgS3Py6LNjGbn/cdwo8Pmsb2zm9K
DAJeog9dPk/zJLxROoQC1H42Y/Hu6/ZgWiAh3QKbZtloZtDgz9bBkpnggzM9+LcJ
NaGw7QL4th0Uz3+defNlYHYKs1gj3x+svtV7yHPvj9f8UHLfMo+NMorjOd7aJsrS
I1g8bB2J6Y8v85Rh03H+aKlAtBWW4wbdFuaUmbAvbu7h1/XAZVJnPK9JDTgf2wlL
6EpPJ07SsmuyzytOZ2n4dDF6tcEjU5c+tDMSEzjbLvsZd9HdYuZqf3mh3qhHPzzo
Y11rSw1jdw0AT/ej9YmPCEZuu0d+V7EPZ0bO69vnTLxgZBxO+kdDKgMB5awuXcxK
+sy0MMkz2NgH1xgQ1iNGm9Gsp/zJ+kKbE1PEUnDYVmNxaEJQTVzwyhUnSAv/xMWF
P6ggc2S8r4SwMJWLTTamxIM17jsWK9aEGTXjhwVZ0UuNaIN+xPPUyrcMxw4Q850B
5MWLObcIno16mqklqcFsNhigiuGuxmWrrPyuHTP74ls89hPsJOgQr+IzrNicNcUa
569KlZ6X+QORBe70QwBXZ+yiUKouJdAfFIOE3q9a1gnsQ3usTyjjKwxhFoWhoLez
5odHPJlJEPl/bZsEU9YuWHGe3FmEKAcQiSxG20EcfL+D2SurbBKj+kWFFLzhcvFY
q3liWuUqwo4i+F5qsorZaySwuQ3j+aPoLvrwaVyxHRlDU9p3l3JI7b9CmZvGYuYr
uDQQuoLamp2IJQOS5oqNti58oDN6QwA6nu4C9wacl5BBg3cdZJFvbKPOL1b5K0Nx
2q8Xhg2B9sbDXh5XLhmEAo4iXTMwaVQk4kweegCJBCT2E+AOLtUKI2Q81xPNX+4p
HeQp/334xeEoXOf999LmM1c0WtVS6tQ+5llHm13ERkCxfLpbkYByN612y3WRFQz3
akm+eH/K3znQIDLCOIttXv4dbwB/nZKv5Fyblt3MC6KpzTlNVU8m3nVJ4Xb+mb3s
5i4IG45SblwatYKHMuXs7i+w8gPpfICyKQijHrV6Wha2fNM8BKbnnam57rqnbtyQ
GDhPndp3qH79fj21RHDhvwYgcS4aArBqBgwRhe1LeooAXk+AM3Lsd6uOkePf+GJa
H/azXpr3AVWSLjbICctNQQDLI47iCqzAlppWnh6zEZS3zHiaJcggWP8K+n7vIjXO
NHYf86ohno49Hh4UPSGAegTNL43Ij/x6oGVHdSaK2rNVFdYAB0GaCbs46Afo1x21
1b6+V4KDDLjU+/Zh9LGXprwELTXTLp9vl8MSOIrUqdQYke9B4Hfy7MkFhYCjtx11
R27iokbHkolmCy/h00F114IEjVhZp1RhDteIqgML3qd2aiNKXIfOt5A30A5TqFSo
kHllvFd9DNTYsN6LAMlgRb05dr36Xb4qPzlMEc8t0BcoEJNHcCgeIisFudNo10Zd
Xiig1PYgfYizKsZLpG9wQWjqazla5T0LKJjnfXi+hWf4VeMsiQKcSrKAGDOr6OW2
Gh/gw4+Uc2XxSpB6u6WiQOI1N/etDZ32kDPot4jgBzraRl83yMSC4R6A01xO/8d4
Sp2sGI11fSVn3wCsmPXmR2MK+Xk39pburBuuKXWMUbJ9Kf6J4yxJPYKa7D4euPRt
prNdLmLUVMAHW8nMDz91qTZ0S/RSi1IvQ+scOhOPEGIrhtBxFD6MnPlI1JIaC5eI
kESU3CQ6bQGiWQ/e80Ak9muItG8s8PRW2CZ4EEoiF5IKWVYft9KVJHhXlYhrS2pz
22qjQuzlNXGbYmfuvNY+X8JvXwCJ3DS2KSeD9u3oLIH90Mx4i6mRsX8AltgCF33c
sP2S4LU58xlbaYbpdNY1HvxUHOx2WYRo9Jr0YmLWbh5vTUQal4q/3QARB62vDK2n
I9bcw1ucNUY92mscja2OW/nltpgMdTRVX5LjUKKY2kzF0LSMYdDHlHGj4qKRdJRq
NWwXbdAW0Gze77xKdweaVyAqoWDoHyk8S798SjpqW71xPRV6ZM75HHggnwsmgQKJ
WMZdMMuKUpvw8EA1Qp7BOeKfANlbW5xqxduwcmqUY0Xb4U8C+TYiBjSHXBTJvg6k
Llt4rfXpJbtnPDnSbt3nB70wXuhPRNq6WO9TszFQbFsJ7NPJ8+8EF/IM++vlmc6N
qsxbwOCK2+/sl1kNgycy5cKMzVKLZesPb5rSSz7jMn9+2tojluzd9Vyue9arX103
OA3BO9idZ2VLvo47znkV96Fd04z7EQuibv4u/+HHatNsae/xTbG0Cq3QvohXERyO
DLg8MkFuVE33xmQc/y/8+8U1Qv9OaDSudY2ttrvcjmh2X8FCeb3tZwCwF/bkUeeo
9t5HXbbowT7xkFRWURuAe3SjPh1V9nGxEuy4RG3eXqpsOUo8hwkC+cxiwGhLszhd
pJJxVINVya1FjBUP3Q/xTcjbqBluUq360FoALtsrxBkhfaKDPAsTGsSxRAFXQJRR
gTRuVyc6n4qC3MOV2hQ2luQvY/xfpqNIsDqhFcd8o8FcV3CiYx6gRCdmQU6VoYEk
JedvdNcvLviRetKaVTyumkdHYpZyMGMo7L5OR5IMQYVcqq5QfJipUjGmPdoLBq3R
XHi/M+WeFRbz0BLSg3bD9bqCxDaSMMNnaMOaUIlocJiRdw9sB6jXbSO0fhjyYXn0
79Fbmg9JwKqw2Jj9jFqSEPHcTojCEMm6GHcM+Uy659+5ELPbR3oa2zomPe2S/kQB
5vA0oHI6ZzggJp2e8P6KTwcKkgUuExyO73zKsZOPS39+kAQUg+Dn+CPAYPZj9M/1
FFwcWmNRO9j9kRpWSTmg891V2+Y8nopk+e6aZQYwubwVb+SYa61Zle6pSrJHfTtx
OkbnzwjVZG3UMBSjxshkqxuObzyFlTgmmAfbp2380pw5odo6UjEiA3ggi5E4gGDj
wgvMWqeiJrYXtnKjyzzzFWbEaSTiXjkiNVMBZTsnMVZG+avY1ni/hAQOVOKCkpne
hYLYyvcI6AJEFmv4n0UdhDaZD5wMYit+JrQpYkmtrfj+TYinYwGx/e2TE8CNz95P
mP/264omwlVHC3TY3QTcAmJlLYE6xq5hqTwcIQYCiXX56XKPAcoY6BkgODtE5H/C
1MmXpFfgs/ZHPQnRKMTV9hW/Yp2hQi8LrJtRbfi6QFfhYgUkICX1R+rQCcxqUhxH
hrCgDN6InGCaeyrO2zJ8CI1WIX/JdKSQycmwo7VOOH6IG1XKBAzjRKv1NSS6vaXc
UWYjfRTCcor8NIjLX91QzxajMz6oK7pgUFgLeMGjWapMfDrSC72fza/JEiYdemBV
szhpf2BPXWBsE36GO1wPGtXWESkFiQ9S+C5N17qtUll7Bpy/XU3W/mQeUvBQNavW
SDtWKosAvAIUKEFjkqumPBAa1OnlA0Rboe0GTnkKIe/5kyt5O5bzRs9ZiF0rBmGw
L5LheSTs8D5GR/CtHws03ITjI0BK/Z0qB7grhnJxjm6YAZVWdCcvy9ZSYb7XVCvU
u8rF+S/kxUcxPWVHuWvsNewt6I2QqccPIpI3tTlz92Con0Zcdioi8rvBwPq3L3qZ
wdoMaix5NFW4u8X12KPZxOiNemngRpCcg15brZg+jXcw/MdA/DApzkqvQVyPxoaZ
CuLOqxjRgGcTxcnvhEGhL5oE9IFhHzrhXbeWhJdxS1OlU2l/bxJtR7jjXM14VQSs
R03GpO8HQQI+AWTX3oHEj/zUtPpR2eYF1GDnfwXbCzuVT4vlTn1pvfHl49QbE3Oz
+TvsexDkYyZAaD89WwRpF4or0MbF5q4xhzMFgUAGLTKftTjRERLCkLqxbhlp4o3/
tjwbyJ6pfIVlSQbKygGPWD7IZQjZ7dN3n/A+mmm5rgwFOUYmk2pEb2sodz8aB4UL
VMVrvWrAH8NOgCOZR00az/sh0cRv4kTXeVSSCJ4nNaSWy72Nmwg6wWyAqm+3jRS8
sigh3LDIQUdsxDL8XJWvAz0aOkCCeh6LzdaPiuvR8wy8mVY/9AzYBsiAHeoiFRFV
Bv6TCGyxDYY9eZdtBD3huBXnzpjpWGk3b3/eFZnh+TEmHCkt5Vv0x5mHTEB8Bptx
HgfYIR80h6nieQvMGkNexJqWhzeSa35iWdhgY57QzE+WtznM2wNsORDlL2uQS5f/
5wFIuQyH+T7kCO0idO6sLGOwxW7nSxwi811t3+c59E59fhWzBYtn9TfTuYqQE4Tb
v2vf71ZwtxiKE+MQuMpAgpNxlIA0awvnxP0omvWoe+/rlshjEwMBzd2APQCwZNKT
OMoxRZWh6+f0cOEBRXQCfS4gXoLBauKOh4dnpVfXnQu1PE7mSiEpDi5hlzedgCd5
CX99jGj/pEfKfbpIxwOERNTRH3kbdPWA/rGYhW6Wz+oX4ykz9vPsPVmmcmjX/RQ6
RHqsXLE9infU2X4Ow5+qejKhDQ17MKdyFHEeM+mWvc4swJRJRCWCVwaC3GNZV52f
EhOfm4+vK0Q72EPZ3+EOhkgdfqO7OdyE8u7GQ8geZKW9xKdRK9s61kw7STwEp/8h
+CULZIIgc/ZfaHVdGP8RMbPerST8gVFKuQPx5tobiSgFM4D05p4KwwG+Y8Kg5aBg
ZXbkuIrERK7vJnQdtmFGwkJ+Ocap8FsyvROLg6INJffCtLAejaZXcRN1SBEE0nl3
/C1OF6SrPPmeLg+hDMq01jXpq90jm47Vv+KniDqvAjaJVAJkf70zlVeZQIZdoTFt
fmxHCAr7/YKrzDCrFG7BUuV0yRFmjw90W65PggyS+HIkQyaUcUPLYdfvhdUdBaNp
cH2QUWA+QzMksPUC51+8ylErOJuoggbo3L+Oflx3CHT/xIzB5BN10dARVCNQoHQQ
YGKzzJf3uerncqpdjGdADkE2vQo/txKRD77VNKnALGnaNmkTY/8SijbwXsEeny02
JbV5qkqULXHvcVbWj5pI8AdDwsO1+orclMBnBvKwOUVEYH5LhFOsHCvt/v3uKCsj
XEkw+dWZ3amH1R4+kyuX1JfTahTdj5Ogs7dl8EVvmZHJZ2pyK8axorPdH89pziJh
SNQYVurC4O28lfIO7cKHq4pWq4l6hTy+sAsJEE83SPzt+y9aD/RAWcHrlUoxgCmQ
3wojukyCGGGfgIcuAmdg1MJb5bOSgDFJm51gdNBchOW57vS1+uQWQEIiR6FbZD9t
e6ZmD9MM2csD8TX/R+FJlEwSjoukrGPWFVoHYhJlUMblytZDsnA370YHWl5I3e9E
yaDuxm+IhNZ5sTDeqLQohuFfDGSA+RS4FzQdiMoZGQa8up72zLoNOX89scVyZaMJ
Bv1vl7JPN+vGAgCe1nGL+vIsebG+LfdL++F3chbOAq+dfICHvI4NihCdm0PeDt37
BRymTGnS/bQVtqDq7/QwfLD7yyLUeZcgrhL8tReTQ1D0oLOFuMWp/84t1ZXNVmo/
DmSQ8DFQW9iHTwafHIMqsIRU6dU+dkvtkBLVoTHv59lvze7BqV9M6crYUo168vxT
8+kouFtFBSvnzYgTJyK1uCUJSzGOLf0oCfYuyU2orHAayPfBGZXq6fcinmju7lDE
6xuJDerzmonvk0qu4/i5efpmoTcQbNvBQibjzfkA0u8gXW4DM5mPl8qO8k8dKI9W
Nr8DrAH0CLhfe+xvq1eq2EM5ddh8Hm7vNjh0/b0Zh4/BghtXg8oI53urTtDIs8VI
LxQwCk1b9BhjlP+7E3ObCxRyz4E2ld6v+qJPuE2k5lhCoHwH5AcHlzM9qq5rua/z
zwCoWqLlDyN1FWfikWXhasNlwJ8kSREySDjN1lUC4wUd6RdaUOhFjDGAIBIEU4Df
BE8QvFUlMQHXKTF6DBEmS9Oykl1kU9aNNvi4VWIW1O+M7N3bwakCaBjkw5gQmLTA
u7IHTdV2+mWyRmNvuqcJKh+uCVXQGNwOQ9iK0Lr2DiANk/sBAyXuZX1Tmzu88cUe
zDieRd5BYwmeuJYS5qAyC0HmGZpdrPfGQL8YzCtdulKcrK8iDquqCW1hIpF8ivvI
F765kJe2Q8uxoSjf/RDC3vXT1x1Vx9qMeS1rzstnSvlyVB4YlUxbitfnXnTLT3Oh
VRfLyx3qXZ5maSxw42VnR14C2N80/YKtf6qTbPJYM1qXYbF8ub1yhstPdGmmKdUe
Np9I1KVbDYADJj2Vxf748UEQaE/qAY45NC20ETNGAAvNvHbZhB011mT44GSj5pP4
083xAtRknuuNmxsngHT+bHD8dTrvaoZtiOI+E/UWpaL/vlwudAtQ9KPW501rouZh
eQ4aTSw7dK1h7jrtGuCyPVLqm3RJPpcyAbk4rdRBuksBUC9cR1kei7kXNNFjMM32
yDi2cGd7PK+EI23C0ectDwlzFfVka7LvJTnH7LiJ43kai3n6s4OMMZI02HIs3Ioa
i/WdXuAFEvTtJvXrWIDUQDUVD8GuXH23YqtbsvwumMAQflmLieSu43BaGFEVkXUT
GxE08E/fKM4gbwP0872oPLQnMW48u4tKMwFb15/8F2/eboL5xbVcBQEIOxgko4Pj
z6/1Flj6mAVDhnJNNMC+9ZcNVVIiergaY0ojiiprHhPtnmdyG5ShmApe4MK2dDx8
u0lqCahCRiZKqhJKyTCECAvoFp2jsPlAJHCOQ8GqZGgzLvEHotgK5RWhuskA3A9N
Pv6F6ntPz/FHyIHlJW6r5CckrN31GF59aXjKoHxwG8FWaIxcv9MY6iDcJQUpOryi
lm2WLzOgPjCJhud33JafZKVxvjJNHQmsYTIVoMLDo+mckNVvjdOfbK+tCUhgK70w
FamFu8GqhepkhdBtc3ZEfLF+Cz/IBZo7C4cK8vfpG0+SpIlq7u1vicmMr1q7zxxs
aIQNrdrEm/fl57yq+AGRhJhyyPg8fi1dRV6bZdoDkVprzPIh7ofapk932IHFHoGq
thnv/BHkNTlhHI7arBP+AztVzZn+pL5W13c4fwQV/dyLw9Euils3CwAeThGFcM/N
9VJaPibi7wR+yqhqbao1TzX47qDWrKaEga9O/LbQe36FGxCOad3XMaXCPhh/d/r+
h6+TyFwQt5E7hFEppd+o7XpIrgBUCKReqU7tHtl6b+VJK7hN1LR9iW9b4urYmnkT
xrPe1xhyL3TMHl2Uy4L8jKypIF7fgviZecoYcAfjSAwEH2rS0L5mgwpyaenSZN18
RyWowt89Ttp/eWuxDCr/PxrsDYxcPDpiH+qBlY3u+MVwUpxFO08W5kn51IdHD1la
wfRg6go/OIAMPjOa9P4BU/ZLfsBDKBsChyDtMiAucZcuQPkDJUlXOuh7r15DuQiQ
PdAAOTmDq6PXC6IlzfKpMMNRCNKOa8EbdONpyDftEcwsUeKh5Z12mRDnujB7/TbO
xhpdEKfKkpioUyrVy0LUjahrTidD4OfLX3eBXBKY9z6iQ9LsPVptW4jCy4xXUcQb
gUqyKsemoCh5JMy5/rDte5dcXyft0x1/qQEhzMYTUQYunqs19k1At9GQUPAQGP+v
06WI59hqPlD+lNzsOT6MRqbniTJmmeZT3Nv9UQAsrobD3ry/j8C2bgdZnA/g8i5v
J8BGkFpWS7BZw6aGnLacOyKxi8gQFetXsE69QMwCYMpyOgb//QKDtGcKBpw461Py
Txj6CHLrLqiLZtqNZUaMjKBtKixgkzldH1mKvAt0lSg8PH85bf20C1HGuy60f7AW
xAoanLDqk17LJz4s1GZpScyVZF0Bo2UpR4dLinlprIIO1OGb9z2bzQsUiOMwqN6c
q9VxNKC7aOf+TwUY9sRmYO+Q8CL1CM2KjGDAa5Y9gRr5RGKon4/j+5E9UR9fzd6K
PydZiTS179JFa5oFQBpdKaimkRnGJFhxLfHNYGk+PpcHDiAyQ8KzkXVkzsl8J4hP
t3wajLvca/wmyPF2D/ht4eXvQgR7vn7wXivTxCUWfuRiBg7nCWspeevwrn0hz0kT
lxItgWHghjKLYwigokfUgdtuUeDWZVdOW+fVnJqfLCVUpumAaUVkRNf01DX5FFR1
DIascuhze3WZDehdJ+376LFqUQJy0JZng9R3zIOEzgQ0TYTMmlJA4fJ0Ynk4VBBi
A7xuOYUSWmcVZJeOTeWuRjzLz/cBSCy5IAmmwr2/RvSXgO6gUrflquI3+i6Gt6tq
xDcp7A9KfjOnB/kiKaGm+bN9q44Qi7O/rkRd9I2bW7UnVT7PY+E8kzR7B+x8y0pU
68UEKxWdlZuDUGE9zPuMGSesDfEMti1xlz+HbT4fDWI4Pzmgaue2inzhiP/RfIOX
uIS2CRZk8NtCk44Mn2UAMJv0yhxO2LfRfepg/8EjDV6q3VlVTJAlhd/HbrI8bEhk
+HhW+sGvE4BI6Q04FMoPx2wuqzPG0nZvRr7wvxJ891IpJ/bOb4MNulswmrnH7cZf
Gq48I+kgPqKjjnY9U8sf9iZvLW7Ur3O2nF99YPUu+hgOKVmzzjon+5cTSjZJ2MFR
eATX3ecF5AEJd6o29L1VkcU4eVkkKcgtjOZVdT8w210qzQ9BUsJkpIqfGUh1M/xf
bbRoL0T0MDRxGAgEKlwR4g9/SIvKv/2/9yT/Ai3FHf4q58waFVPInJzw9vQNz/J3
spOMmJgqhgTL1Dm3NY2pcY7O5PdIyCZMIjQIHNQsxrzkhNFh0f/5SQmnOWEeuhvY
Z05RnDYTQhw5scm40bX1btVwJ/JNkfS+qPw2M0ceNUQKcTM/xoBkm6oWAvcAg16L
jfNq+ubwfpSfvgtNk57kXyGaXEDqmCMRujpWhDHpmVuZYYb0q6AwStXDA7KhJiaI
l7zPzR5sfeaD7R88+27D16j7zstzluTmel5ok1vqnbgfdUF3jbfP+UQuCgrnYnEi
C2STVic6CCnA3MnS7EHz9cphc0yNkhS3PgWjX4fDUbySB4wf/faf9Kv9IByeHWR0
7KBHOPs48vA6+PjX5gIGO7sT8ojTMhK+BgpW6qUjDPNjxOsEsm3osKLR7AXGLcQk
VfctZ806ORngKDCP0rg+blqxN5DRd0iU2s14Ce3rkwhYj1BQP7nyyhE4yYxG13ca
niw5uI09vlTodgZuL00UXpsjIrc14SouRlDJEjX47q8LXEDeiRfPXtgNk3Apadxc
grNnvxJ6XZzVPVtvh73/yR5RKQRn0GtSlrXwwyGcBqRXWIbzR45PqnNZ5WIxjkBl
mLsJGcnijO8GfxUCnu09jOURvI+j+h0IPB/k7j7IzshsZOtg/tWebwZldWG4cIDe
1MyJDFfV+H6Txs6SzzSgV4r6zEm5M0OCo7FPhu1p23EuGfwJqAiOWCuY/+ehdIAZ
am+sSyRqRySeLUFM+HO3rX0swqxqjZGO+51U9rlzicXM0j5Rbb/tDOPELO1vVGY8
o8k8vsO6c5wvL2sqwb9/kX876Use+4e2XB7TLEw3X4Ianxh1AyOtWE47VXOINnMm
a1fA7b7CkGfPw2BcfmE4sil3Pq94z+lBPAPYuBq29+QOCL0pov3xT4VzGMw40QWq
nhx766tOETPXg7rsvoLIBg0uIwJqemyfv8YF5E5m5OrDOXNzNsGeEaK5vMc6GVSp
doainGZe6pJR8/pLT6qKUI+hgI1Tf/paRP7XP+l5+ybxSyFIy7vvgHTXkC2FlaTc
LII1ANYRPvsVHBowFZ2/XvkJ+upHZG1jPf5FTeVIEBuCdvKrj4BY+acflgGMASAD
NapaN9bMsI4Zv9MhTbS8NC9civd+uowQFs44I2pj8Q+o4qbF0unaW8hrd01yRTZp
U/n8r6T5chAr1SXdO6anLdD8MQDdG0RE3itMcgQfzOxGNqHFLhxR+w8LZN/6uMI6
MobYvHKcAT3sI/JmiJrhlMLIOTZxbQDJ4f5GDuOENgyJWKXhT6hiTMb6qgKFPNU/
+XNdDcG+bM354LJfRFVsJNtmYSi4A4Lz8/mK4JEYVqVe5V87pDF6jDr/UNsFALtB
MpFJ+OG4gl0Xv2mf++9GX7HhktPYBYERTzA2o7QmZqgsVuYXe5j1LWAn2XOdYjpl
mIcKBaZjiBDeXj54GNE0NFfzzUiDQ7G3u2D1BTjCdDSkQccThGCzHdYcovtomYY2
8x0nRBNQCR4ZZYn/PJ64M2MBSlAnn7DxO7xwtWLXcMtQ6dJzT32WnJI6Vu8T7VJy
yzwHp43nT+ik9Lt529u4zBZV1oQADoluFOfJ2EVrys8TMopSOIcdPA6uZ1s8DQ1w
kBuG8uClKsqqE/eMKTADPw7mkRyjE9NGKCnOJB0AsK5gxWLvBOLhaZsx7b8WxpNn
l2N2NFwRl/pB8TXNfaixWEEm63dpXB9js2RJnkTJQvU3YRtrfkbsidp1h+B7u9Qc
XKKPipVAObksB3OoOJRayKdkT5EMDATzlzsengqOBLOSpHsWkXJM+ccAfoei7VkS
qPh/jzUB+rKyJZ9inBYuGOWhV/TRSj8KHr9HsenqvzLn/w0iLSE1nX267vyVyfZ2
hM+MtIZ/52fd9+1kdNpq1NwtKCH6STI8rYcfaSQHpl6gjPgMoyd4VipknLXuFr/h
1QbS9aefBt3Tf9FUMG3NS6GgPBtVcfKWyE8J3r9SI4q/1AdhGGFIaP1EhvGf/y94
ks+ssrlUqPDmDg+tsMyQxngNSM5BskhKZ7AUmPwppP+gN9X408zxSPwfbZNm2/h/
JAQtUuxcadPj991y4P7Wid/Ak3uIuyqlCIWUCLBPff5AIHS7326+wRBV7fLYK6Gw
s8zZaQ8FK2QNnphMvpum0IJgQ9LOoMvr+WJEdnRkTr5G+aUn1a9kG5DAjn/0P0x8
IzNCJT7/c2Njakk8JHz5Lx9tY9+qxAYNE8Wb2vzaG0iBG+VkgbX7fDZklwHj2mk5
AbGY8qZ+pHqiKunFyf+9GybFvctJoRg0dgr4adiE5dxqpqgkrl3MTvqZpvdS37Tz
aQABBa22EZy50W4D9gEZtDL3bkyF4AATixQAa7f2CGLplguBYH+fYg7V2RN6oFyC
57cjilvFompeLhn+o/ATZ69VT1xDXDVGqKYpS9CZQRmvaNU3sodnY3XK9Oro3s7Y
SEj4v4sC5CFVcL/VCyRgwppdB8NQwQrWNqgTBPepMvZUxYWqdCQ1rbhAeRBWGhjf
ZqmGN8iatRRka46ZmVwcCNeS1ZgW5mx1mfObkELLkXiqRKfNqkHtJ64OvUcRFrpJ
auOhbam7MzAZbms7c/RYGs0XofZaFCelyMR4LKkTHPTqnFaZPA9zORLKGNVZcrvv
20QSiyLV3ENSg/dI3HqZsnPn9W6S+cFzKygSHX4AQe0bs7QJZ4Fzhas8bGOsf6/8
wDjFYVSHW59AD4K8UqsBCp4J6wZstM91rJC/vc9J79fOElVCS9F3Tg/wGGayi/Rs
bLrlXHFEan385VF+LgdRub9+ykzdQJndtSX+z+GkVkT7VUrMVd07EAQZ2FO702G5
5Yjt9KgDlLmlPE0HPJd2ZnV/8qvf+7KQ+cPnjlk5FISflzwrrLqelhZsBzaVMaBZ
YRP6IAGuGYi06dMix7WGvJ2VybQq/qlLVAQyavtvIdnXXgUnB6Z5ykCGSAO4Kecu
bwmCDIx9fw8OLMPbYAziesdEiDMfISoZgqnp4/1WkSTdo422CpfQpB9773ht6gQg
VAOEEW/iXJjpJWPqIhrbVA5fe7eO+7JZ0DMK7hJJQ/FC0rU+Iq0GCitFnKjWNAKD
plgf7FHgjovm2QCrzNWDHxioMV54LsEo0Xa4JuQTZ1n6HqRBv1EA03IIyVSDXRI5
l6SIguH3clEApJaNscJrLIvtEUbrL7wLlZjPw0g2DAksbwyp+AX78VGMrbTYN7pY
5GXt4yz+O8kjo6U0lqxECGD5j0gX5/PmhFlI4ePAZjVAgS4Zdga9f9g8twTeam/E
kS+V1j6G2hr+zXUSqd/vWr01RGLu+TGRjRTu/2Ca3p4EzUcLKTj3YtR8cH87FJfH
X8sXons2Pint1Vj2j5or3VkFa5D8AT/Ht4lfqFaEJE9b5sSV4JE47QBpr9CjGX+f
3X4Y2VMiKF+bBjm/3MWI0B8SUuQ7v7mf8crqdBQwQ3eCOFGJqikId3ByImlVCkUi
Wj2n829MIWHAHNmbemPwUenw/cY4JfmmEVsM3XJSkBpksjoEN0Kb9Ms6x4wsVnmT
+/2ac6AA0y1yXcjMlJ5HmxyHwAp6RUV6icjcS1O+3y39T9rgcuKE9ImKt4q5pNHV
uTWB39Bj8/OJmaj8WR3x11U26V1c2joni5Y6SVlJh0ODLbXwy2phs1MKkkwxwZPb
P+8K4xneNHnPI731De9E+FQcjaoYxWavpbQ2Wvg/zBsxU1pH3M9cLLPgL6+yRFRI
ViZGZ0GqAvoLsfyQzA8YtIuHr34VLfXYJVJCVY9tBUpfo12Y6LtWFwigA4VR5ZjT
+6Aoc/EGaCx9RI0rQuYJCx+McddED0JaNtDBRLQAw4KYMg+WBIhgixfJGr6GSfuK
8GNWGkeoTVUmMdpqNNNMDeePI6zZP13rcUe/8yLb0fKGjs5inLoBiFzQhEMDRvOu
wu0zBcAlN3RkmoYaEPHtF524kHZNQ2iCqAhJKM6r2ciXenk8KQNJTBYjj/04lqSD
i2auNUIy4xKhxQET+e6Xd7Ep4UzkPsNZFRICoLpjBKIpA484uVXD5Z2Zg188Ei69
DZM2wzOvhh6T23FNvG4c8zpmWzkALllsPBRxRbrNfF10IMBuZ/NwoEIayJyCHT6Q
fPXk636olKGJRr1cZuwz5SQwXJIBeO/26qs6AqSdubp6B/1MQD41sMbnMo5NFe4X
bgi9c37fFcVtROBK9d8a3q1SyseQeCxjGiGAlVeBTEZSq9fepLIQ2MYE0qkqmb4W
zlgyintdzsdWTA4G5P+SMTt1YbNbKWnS4ls+CxotysxYU+vBHH6i7CyP4bEhnV07
2LY/WAN5kr0oe5g8kk5i0OpeTG9sGKCkthyfxUgM3+BAHvH4HrqWgFR0SDBgcEr3
gykeNxj1Fey8gfj5Mk4tmSzb7SHGoDqNN1hH1NDBesQWNkA7PmuqI2KJnmv4FLi4
BTA8FgTHPBX7o4Gd4uApO/8XTR76fTFDNMzTe5PjbDm8OLeha74vEofO4WxrcZDx
AXz9qSG/2DH+f1MpAs7TPh99SAQgXUUFv8ir6oMz25XK3X1QS9R53N14Tyy/xUk0
XMCtDxsyv5MQiwrXOB3LLLOg7HxGxfz98WxGWoQRiE4vcWyWtFHdPujcyi6CaRgc
4trIRuEkiNeUoOJR68l9yPZH/l6lmuQzo/6NzGLQnafIEuq9h7TW9mQS+UcflCKJ
fsk7Xb5EVg/r3in7ltRn8kOnl75tzgemNARjSVjGDn3KUqP0Uk3WOhaMnogyj1bq
3pC4G+E8ib3AqE2ygB7JRu0ORCoxrkZyLwGFnQLcOdHe1ZB1pl4Q9f/6f5d6FR3k
7+C0fULWysD9DsDm8cNx8utFVt19iquU1hUiLo4j8j2dHQO6adXMCxcrw/+Fx5ET
fEWwGu2KCFFMN9X/Inzb9ti+8yg+6lH4byGZB/QpmDMzv6PFhASP2oZvR0dDv2rd
MXgky5rRDC/C2HNZriezENGsp14FUJlch9w5UEF/Ecj7QZxfz2cSWo1gzA9Kcukl
4R388yKEfN/iN4611z8txG+tXvKe3FKBT0d2f9oqGIPfMYwDadmIL57iEENF/6iN
F38ms62b146oGY5CnklLQFcBJwgtST+l5wFqrS3+QUELf8XncyzfMvb+k3eD9EmN
nWW434Cu0C0LjE5F/T6A6MCO8tr9lE4yEaJG234FqrDjrr/HzNNfIBlrvgjmH8eb
vLbVme22HvOav372hNpRU9GD7vXDl7tLe1jJ+5uLlhdIDhAUuSG8hmSTgPeYvpGi
RNbUnNzzFCFpkq+upUJL5wNJM+J3ScKRAmvrOPNN21EkYBJfjlg/yLZV0LvA3OIM
hStVO6GWi2USLgFH4wwwG4iQu+oV7FTXtOJGp6nYcmnKPDtKRW4D2BqYIGUQ3ghQ
AwyiJ1c3q6CLZ4d1oGvbsj7ETCzSgM7uSaQrnyEzFDdObjDUzwY1xwz2Po9cSTtS
JRogPcqvd3z1jyLKjG+nRubBPk34qkgAoVOFDJtDYr9O9ZsZG6XGTGx6ZpqfFvYC
3P0SfGH8GyPu/kx/OLJOTwuKA2UxRdM6rFBnnfj6ktWNbvpumTMx35zOTw36yTY+
Aka6hfYehDW0mT9FERwcoHK0Du1laN0ggN5v80/OQj7vZbMoEj4X0WpivDO9DTmS
H2NpFVOJverwH1Q/LPGoHD3n8LYiwYDNF3YOF9sC9q9D3AlB7rTPmzdn7bTwN59X
ndUKfei9xx6scpAxTBHrQVKQ2K1c8sVLgBXhfNxumNIogI5Ki1th5k6rfnwJ/qOT
0lIFteV3kTWjvyJ3ZAbzN/zs001PI/8e1PepslYAMBWj3wvF/wGc2sNTzPTh0rtm
ArkXZhiI8KBOH0sy2aeBv5ZH6AqJXMN8fj2q+zejomjsVTTT09aSLdEHiBR2SjjJ
TRfpc9hPtuLA8d2rsrjXIzbbUiPXTyYfD88DHGYzSed+64dNynrQHedybA7PJ7n9
H2GUF/y7M01LpcrgGnwFI82+EBf7sY66c9Ae87h2dNPOaFJ3Qe1wjiAoQ+l0Odxg
COUcKLitmOO2Yr26dOzTDIaY1LoM5MiN7vsNA1vVRaOGHyHsSIfPh56wBgACb0tX
2T8eCareEqSy1dYFhxmnqzJ2yNOsAh9+jFUM5wmCisu98Wf/9sF20OpDNKDRtYyw
idZxB8tyVE8BDe8FiCZz1IT/OHaA8obQTafLxpWvINjbZAG4ETFifS1QlJxNYAlH
Oi2iy7F+k6xz+MP0D1H1s31N0zbepKRPMlfd1E+oQUVGSx9P8y4aLDchHdBvDCQL
Nj1tKStpKnDUTPocb5rF5nRkTk5D0FmutfK8qPzAimLlq54grIt6lWIL7kKwshv0
gJ1xIdSkN8yaTMSCvfhTmLR+ed/bdSpFge09fVx55vQvRskgrWTHsXqYzNeOeA8M
PP/n+MjgAWIc7KkiZfHlNz8Smc0z202lg+LpAHATk8Mv28nNJ5m0Jez5jxRjEVqY
jEChq6EixF78tCTIs5t2oVRzqENsjcPm6cSLeryEQT88Al/9DocTwbkzp/81ZHr4
RvFy046PQVz+YHOdUarfVsAcV9q9VLUg10TfYxkt5NgslNS6n8Sj4BFfLP9o8kKE
9QLIT/D3CcxmwSPCID2JoF38g7rPoQrpYEYjGYdwgREO9cvqSF0vG/t90NYBB1I7
c0KezBTVcVYJjIgT6oq7lARYYNEbuRNkyfZqkPVZ+7ogEQ7uR3Kil9f2wFD+TNBr
tWoBJr3eB1g4PCphYXUsPxE/GQw7KgqKr/T7696WvC5b+YcwuvnSUuxOgZZhkmul
alOEI1g4aAJgybfR2cNh9Zm1M/IG3rvmgdGzh1DgwBNlukZAn2ByJzV1rfWE0AKQ
HuF5VhWhRqbtESJbLPD4UGUIupxlogvvNJXfUDg8Jrl4O0qzqzWZSiaNbasGip2s
tmRcCXat8KZF4DjTK5D42XIEB13ISPs1O1l9NWXDK+kaT8JbyRs/YY78fRSGuUDd
bCbdbSyFRA2F4Pv5XUCiy+1r9SrPx5uNcgyDoj5xyPuCKUiapMlsnkLFZCg08Zf+
nljH8PfokSp8av5zD3gI5sioo0FQrX92XGSDnyWdVqwa/eD/pdDWH8J8Bzb8i1d5
5mEKzMrR4X+PsTHZey8wWLvhEpe51sQ00zRcRJZIuPf2r6nuo3hee/I33IsVAIQO
Q1sh2ClvCofhxaoJhSgX8b69M7U8FXPsDaFJLyk4PaihYMoNMeOC4FSxGMFkLFtQ
om42ENFpSunBmLxVi/x/2qUMCKfQbNclwWw3OGQaTiEFC28P5R/o6nhH2pR3FggE
CLK0lvKA8GlVy5uV8pAWUbwNgDVtp+56UgFChfRLQm41w5feEvcaN4bll+J3ArZc
lgLzGVM5s6Xgdqy/wcuiT1mz9pD5viNuFpG6TXkUxJlGQqfJlFyzOyFO53fzn7gw
gRVL0LSBtTVuS0Jcagjo/vTyHjERvVlXUUInJRQ6nQPWojmYM6I0pi7sQwtRgdlV
YDDtmixx3AyAmF4k9qDrUJCZcI1iNkOXqhi81ganynLj5/m4lRhsn+MKYyb1FBIE
L69qOr0NMZKJrzYrOxTiOv7x3WcLMCNx9cjmcjpNlc4Fv56IMwyNnmseGcx/yf3c
rVC0t1z7707K8jthXlrloVmUkGm9ApLgPwbQU79T2sr6iucs+EuWwoOHp5onNBAZ
1C0g5MXB6WpcMxRnRnfFjdHzUALhxDqbdFpw1sG1WG5C9eCp4Edw7yMTf2N+bK8e
WhTye4Ym0DMGFbCfuXwAp2tiXZwHy73X0ZD1nNJWvkQJUTrKgFM7hnAklDAlSD7X
vNkBMWp2Yc7F9OieW15Sw40y9paddI1xHabKNdcwtIuuaQ9UfIlUz8zMWyY8OCgb
6J8W1Ghby/vU/MaoAdOMsZ4HLIbYE2InMgVd3UZkpnCT9vNM1SluSxdwu0IeMdcE
xBqzkvblTYhuIASgFZkTd+OCH5uD0MMqdkb8XpiYV52MzO99NR1flyQN2isGOmOO
/c9rgDEK6p/Ptru+R9rvPxxNOAky/O4xqeck6hiJZGxUEqXzVhMAHv9ZUQOoiP5K
zoA5p0Ac+OB2XoMbB+0NGbDRUCt1O3H13Zkb2NrW1LPBtYg/Krh8QErE8AxrYYd8
M0V0dSKCIJEYpuQnVCzJdzWmZAe7u1Blq65stZRSKZ4qymAVoLAWIXDurfo7kUq5
W5eLSzOCBrnlaR6l5DQka6L5iG0eX5KKlN/WOoGBSCzmobt/m7QtHohg+LJmvN9O
NdDIJycPkH37lwXuel5ZRu9lB7wB8nbTgZvAtZ3FiWgZQ4d4+jUbkIk2wO5Uxd3u
BQS/g+Sq4BnBzvrbwvZIS06CWonJ3AfNCwAFCeJsBGe/61q6rDanfSA9z3sZnZ7l
r+gh9+E9ljHAYdP1g1tJLUUrOdFO0ZXvYiJeiVuMB8i/OGkpFuyySoEwIkvjmvmf
7R0GeEL0hPZhZFVZUCYb8i1u8ga46X0svQBrZyxIf86M5b4FzOxvUnzwo9wy/xTk
uOwQxf3zdAstZfsPh1sxyF3vrIFUR/stV+mpFCu7SPIRHyQc0QA8zv2z71u7OIaA
5YU6ZfJipgLmdWQvB3OYz4qbLhK1nOjHIW7Kv57h2fXlRsxNZfWzgi4pDOyRgvRg
W40eiunBSH0Mek8e/mwJfW9n1QB6bHEMGpSkRASGunisIEs5g/mj4991l9lhMX2t
EXI/qzDhMzIWEFNoTchoGJVbXIB4GFsMQMNdRH36QGdWtL3aGREhlPIFB7BSvHW/
b/7yjMumLShiM6xvkG0pf/tCTCoZSKGM1xfGzGVElZZianog1b44NC07NAoKy0Cr
X6cbx7F+oV8+Ch+nESsUVyLuEiFLaejm9VrglRYwCQTmvfTVcvadAO7rn19QOypa
LfxmjQlZnnoM2p4Y2fTa4AYrqLp4IOyd+Vw3TtdyD2vmJ4TI70D3hdhbwrbn82rz
twQSPCklb95g9Jtc0Jk33clHOKy9q81YzXuOyWiUt0SplJuKNlY8ndjhAJaHXIdU
aKmdMtOEke+OfCIhT7R1lKFm9KyYNVdvGBDEpxlo1eaxu2SVOtsa6X/J1niFuqq0
2u7aNAfHQ47xMBmpga2HK4qIvTKBWkx0oX4lwTdzBgNo1DodM8qc23DRylRGI8Mf
EieSV1LbAfiUOSRJnRJLQ/I3SOFF+mxuhoPV3PeHUwIeLhXmJczvKaarTJgWj9hG
GudMZDFhpspwyD0g3rAEFZprttzsHA+Z9Qi7r111Uu6TYnzB4hMR/DGPUaPCIFXP
eIYfVo331UtXoW2d/hwDzxBbQxzsY/YgqqFJ0DbS7kq0DC2zt4yn7cycYgYn/b9G
LDsEMMgQosoL0gqrbLiIVywVYgROGV11KFhCK2EUotbcFTwRvrVhaHuksHAYJVQU
hZ9HUaS1MWrDSvWv0FYEOKARCWXFVvutY+NpcY5/FCVE68vrc9xUg/YZeWQL0I/W
klPM1nQebLodYorh5+i4yv44+B0sC9yyfLA4kcWymiDEo6ce9yT1oZCvdFtJkDd1
l3Z0Kr9nRHa1UsALK8MNq38rGUT1B8VnvQ/juHgPLzESY07YowQfIULNVJI1JbVz
P0nqEHcE9tB/7o2ZORQpx04UpHBZr0hm6YlDWeWy3O2/lc062YjOFrR1IWLKldf8
4WHcp7+Hr2i53S8PO+TXtvb4ZGQfN3fW5kcNEkFhJhJEhyz+n3URZZhRb1l7ue5a
tvdkQIRUvQk9IpZQlC334n48GqHLr5mC0vf8GJT93IDmfrL/HzwDtG4KjnzcbdGP
8yAs+il1acSCIxYEXEdEZsNeHLjPljNiF3n0A2mcdgjbDaGoe1YS3dWG8bTyg9IJ
OkehQRSIeEcg9eGqxxprtUQKlTCrG6xsqogPdVS69Ey4MRMLaMJfGDJrb2WsXvf/
gzJlQWsyeWPo2qayazxBz2BP8Zrl2LIx/wFjlvevJK9T4h0Ek4TpsF6W64rsg/6D
OZfpIpIeBY7rA4ITqR9ncPvMidDtXisQ5dRR+oCEfGqPkkvF379alEVKSPNYEMl/
DCWWoC6eSJN0o0xXLMJxymTsg9QBe22dVcJ6ILDo53ha8q42rPPaY9CSurK3hUGy
h/KVH9d1OpUi4QuNfQYTHqVzwU+uQkqAGPA+WbGpJ/H6rtKRGniDnmw3KaWCUld3
xy+Vq2qMpQ7j79ii3rIbwjVhWW7xl3KfvqgiZnMm4zqs+NMAQ2ZlGEmuAmHLoqlk
/U0vwOYjEEBxgZ81oHg8CRQ6PLllvdaUsnXvDwG29DnK/EEsN13NH741kLzHCW6R
qVj+pRpM7YmeFvt6DR38VHNe+1V1URy3cgKHFqHemmByvmYXeJ64iFtgvgkDaiz7
fUFmGEj6+F5P/xrNHdOcK+dXMOICT/Zomnjs0LA4sUO5bM+0kZxnPO817LrNuvp9
wTCuihLildHd6wqq+uQRFqbagEIV1uFB8Inel3T/NOBryY1L7MfqGBCm3G9bvJwV
S2WUiTFatiLmElib4eXHhEDrNjjFPNwcjchIlOMfTLuI5s0HMzg6BBuFomr/p365
vp5Akc2kUwAE+MrLigF7yepIeUfJwRgfIqBo6RM1nre5VFeYV/mDot0DZwvdR74P
++R5CspmiyvTtOriKm2/Wscz2qeVdDHTjYR8fYBONRPlHVwHlIA+Qyt41QYPIlol
zY7yIV5kkrQEz2mwm97YNpi6o5C0C7SIJl9UZ46c/IJMVsr0wZtnhZR5lcTdoYPO
2uNa6wISUCfLaUuNA0OslBMrWB3dwSKqLbh/ZmOvSOJxzIaXoMkIlFo7FrjnONZW
dvWjSQz1gjxbLOC7g0HxXYRY5wWq1tAiBiXxjMoNH8irc5UTmoNzp9vP/6+2L149
KL8Wm4fNNa0cHI9NLdx751mT+Go+XfNJAFYyFtxQPG+PSS6AE1ROJzspUgD7bZqW
T09zeKYHkiasYuGdM33smlvLtXPc3tHdcrfjohybJMjJWW7DSY3kiWpprBi1NA3F
x/rkp6K1TMu8WsRHeCeR2njtZg4jkLrXaQ01w7zLcTIYECQTaY16VkqzF7Usm5oI
XhvpjZPzOTSzUy0G6j91+cP8wV+cohkJOPbtxiqZ4PybyDhF1ZcKsGAv+XT6+zUi
acTZibQ6YVhe1odeUSaUpnZnb8T0SYf4+qASQE3bE6fcyiUOmUpnTCIhaRC8yMSc
J/YHkZ7UkA4zihdWwpPCXNFfoVw1nXl0mKFtkIMMlUKjI819FHwAf2EL026xdd95
i/Jg0S6AkHVTkbms+vIt8+O3C3SDoyg5oQZrR0q41PeFjdAOMY70gSTYCJsBTSqR
vtpSaRkBjYXaM33mhfvIem+St7BeojW54gyaXsuRBA/N4jaG6gM9Nnrst/zJM1O+
3+hr2gBFkK5+YW1eOe7xs1oZ8tqwBTRiRToHYg71HxCJOe/AMjqnsdAw9ldqW3KW
rz6fYkRaaEoOg4AUx1khzjny89dykj6B18QH9XJUSUpInaTR+jb1vkVUp9XdctXp
IJ2DzJ5WlQt/JLewuLkMLUXn/6bYI+awS02t+ClV6lFekyjqIVWQouDkAky9M220
1q11djaMF/8bHvCjDk7EC3I9d8HRsDgi0mHOUV/acHkxMRobhZG0Ecx88JaLVMq0
rNsqluNWKZAjjT1nEcWBQjd5BLgn0289y6sVV5cJZiPI8IUqOXqyI2fwrXxCR5Qx
4br0Jtc2JealwOfpx5X3WU0iCFZK+PAeL5OEkJMxNAakJuprzJe87vDVCfshGj4H
K2eF5+WrpNmNLZL7fLVHOF7sUvGl62LfjzvxWne1ayabeSSEZb6pQYHidmFX3BHu
H53Cc/mnUM3LS72lcp4H+8B+ZN8Evtv5lev5Te/gSdQEdihtlxs/7l6vtzMuwu8s
WF9r0Z/vNY2qLGJ76BKzx3Pgd5HSeUELKw4Nsm0w94iguLwf8upY3ufVXqp8pqAH
87hOf3jOyjTXNbG+OzUrUSNJlAki1Os3hJvql/HjCmxlVCjHyIRyxq1IR3+Bgwjk
F2phCNQJ6binLFvu0Zkd53neAjYD81jrxrnA1DwYEONMg538RHUgrm6oCn5lqmU1
v4k/1pUsbXdrxjETETXnrR1DJQAvll5rhhAYQseNUrZ3K45T8xqs0dKkCUeFd3RL
zgRtvMVXnZ3Aq3hfG/1W20hCKop2Qmg7sbUgFIGebeUNaTYhDJw2v93DzqveRvZM
0slgm+iH4iZmV6g6XuOY9cb+wSroylREtexhXINMGAQXznfTPboc4307b5csqSZM
rDnll29Db+4hWtN5yJvPoBwCwbWgZXcN4nSswGNQnkmYv89uHcAlGoRuyiLcqeRU
u7iMuQYcOhrMtAbxrJpHQiSq/QBeOtzBuWZ7bkO7qIugwtwxNABpL825Lw+9pMmn
09xL9v5MhGqkwcbN+aYdVr3rZGuYSPepnc8U6x/jBC60sYvAMSjYVLuYng1FHh8W
CqUdqH9Sa763yto+ogfoQAiFnBwplJNELEDlRRpSdz36aadyySDJoVLdvR6hB+kU
MKR+jYAwM1kPBEnMF7+wg6m/K2gS09mnYsK7zO3EICsshdb4ganv0zgiZGiHuxpJ
ipfgZK5WfQ4CdDHnALHuOyzyLEewwf5Nfu3brcADQ7tUsC1fv2WPb0r4hcee6eTJ
VJHCUVuPZCzWvLftpAeDEIhjjm0vwWA6Bny+Wi7i0fJQ92kFyQoElocOrrUNTFm0
/m7GAjzhR8eAp/Z2BVWCw/ALjGcy8U/uoOuI5XLeTNKYqy/CwVE44ZndnEUMYLN6
tiCVnRIX902bh6s0X210JbK5vQE/Y0Sz/rqJ9XJjUEvhedZYFlNrxX9LuZIxvgEk
F+Nqk2piJsIAGG/u8J/QJP294kaL8W2sYz0yqvySwRj/V68NgkVPzZP6Bst8Z/hw
reRm+Jtqyraq5pC+c8/H/kHNl+mlpQVbRHjVPMmBjA8B2QWrmawFV86LQWvvoweU
MsEfWJDATI0nTOblJs7fqQnSwKKV5FTqqk3nbAht5UZNnMJa3/1m+N/8s7claNeh
6x5TcbaWS61XynKb1SU6CKOKaR+ci/JlUW6bli2Lts23PvYae548l1LuSUQm9OrV
RJ50by34BJOMJgnPh+o/mzfdLpEXzTNXbauWGJ0EuPKrQYS+BUviXFpYLk0YFbZW
TiwYMqJxWwx1KV/CGtp+55ieGwToXy78m8gpQWcHPeYHv7t+AJGROCgpz5FZtjbb
GsK3Jd2v3JVi/z+fqd7qKxIf4ml1CRUjk+5yNfNvVk/U7O5fUUY76SaMmvF1i+4L
ksJeKg3BCRCXOaoOWu74vaBoU3U94q+rjHfcwWRRmRPOj8HpIxil1jg3zwBR0mnq
LaPM9EZ1RYaRf2gT0RUql6N8fNoydAPaXu+buu0HdDJxU3TIa51TZfd0pL9alVZm
7EiSHLa6oRJgJYxr0AhDiO7+50ZDghiDWeE0Wbkz0/xROXigXpcFxtJ29BXqHA7X
wHILXNnlO3WjhH7GHci0mICEZjphMQ5Xf44zmalz3xZvKkBSp+8tL8KnSKWy6Qvk
GpVjC5RvQR+rgbhyhlqo/14lb9HC6D1kRGDIQANU4hWLGsxqMHy9Kj6SXB8fEmDF
SPoQ4T2MWvJjlO3UBoXPVK7LyZ8HYTtINBQKRzkubm+FMl2IciFOOaBVF3rsf1vm
GYK6CCI8ldeo+Yt222GJY6JtGmBPHKx60g0MOJuJt+rMpOawyDPwOBg61phYVvOn
6P1o72lSvkqnifB9Yke+UC0fH0vAMA5z86phd9PvohcPJjO1gluMROoMGcuFZL7s
dVX0lhUluBAhTuFrb1MOI9djY/L/Z9aUi/fAGBHnWcmHpKZnla6Ms/3yWx4Ib9G2
8jNeP5ts8SX6MXptVaD+WRnEW3RhPcYCHOsFKClvDQRXMaJCCtRTSs1i8uzvNZfF
aukQYhHs+1Eb10ZAb9m1egTv2xaKK7LyuZ2qSmKZyidjZH/dfzj5/pJTjAt5gRIg
XJ7LAjU4o9X4l0f4Cxyjwnddgjc32k7D0Ke+FqP15/P2p3lyswpQz1AcDImyhwOx
pHb3pjpC+0vH9fZpEZ28+R2bC6gV/Mc2lC4Al2fWEr3UvkhSwT+6xpttyLCgAoKV
dg9Y8Gg8ZxCKMA7vwUvC3ymU/V613UPJTAgnuyuzFEwEc5N2VtbeqMTBUgj1XHCQ
mCEIePJUFmcgQ6ieSfvAxCx6DoMLrPMZP5zXu3J/7ND0yRpZNpfx2O2V4bnIcHoa
aD8pqYwa1Yj8+kjI4Vs/RFS3sXzpyjARtGkyuMxDi6WQ5i7/gRaNgiKLLCJjDQg+
h8DALZ5BmBMS78b57r1kWeNK7kZ5JbDqk5rvcZzDv6Ik1xmFfp0WynDm1lkE3Ieb
wnRs6PVXRYOuFNo4FmOec+2xcLcL63LeBPsACrmGOM2mysk5xrNdzPxGEawL0Kpx
85VT1NBjbXdQLlsxUL4I6APUzTLmK8t5uU5YQ7kuK3mgDOWoHh5UtTEQ3cqg0Hms
mF9u90Fv53A45HNAgjJkq4cO71TtRwYhpmNAEl8S0om+zYc53yV25T/wuz+Ivo+W
z4UYu51LSqHJbG3E1vp/S+jgXhkdEYyBVuTGm7MuZlyvmOOhUKLaf/ez4xNAFGKP
Mie4xhEHvgUllQx2TqDu8s6fmEMHgDKZtIcIHN/HnkudKCTCG/bpw1CWLM3pVzcN
8+9WbtPknLcrjhZnvK3SoqWYQu2wv+IYSp/Iq+pm7rsH90QqLhiAuiccu3n63pt8
1+HiXCXNxpILNMxZQiHjUU+PXrZoE21hhluUV4NofuqDCr4cbpku3W9yVQ+FvVKV
/HLpEV84zIQNX1r7FNPbUiEXzpyAc22naIHTfaQSchvF5nRTAEvvdPDOaoFpdRMg
ieXY0/juxO0MvjoKqbfvl6ZsLksUnJ7EeTRGVTZ5a25ngYO6dcfUDdU9vv086j4k
qkY/zCw1pu0BX8nV/OFODUsGlCEgRbZ4zI96+wB81eBUdJgVj2MEgB92ziPXI358
NUboQm8gjG2PIPPjgiGrMkhAc31Mc8QW1iycc3oQwlwvWYhrcp9vKQXty8ffiPwb
xLNJdr40ES4g6iAYqvCRAKd8ZR6p5nkGS+z5Isjlw2iC0sfhfOTwbr9ZcW6hzrJv
EWjxvdfh64IjuPKv7YFoNmOZSseIoFSxdBhZ79CTQHzcIKkiZtBFxSaFiSCo8/Q6
mX94wO9pvRgsWx8MAIwnrO1YEdHUj8C0R+Vww4HPtimvTwdqbeLz8gNI7p0Qvqwr
rnSEc0OkKFAiBhGCGmPrVOZTUMpaGKU43lYd7VrgBuNTPrUCJ+oY9LL26AygN0dh
4Sgp+83t1Ov4fM65C2EXXHSR0t+xXxXlB6KgXuFGLJ9NEh3VYxKgP9pRmZXBVXEf
ymbK4AlCnE/QcUqSBxspR/YZZTW5ORr90qMJ/ByWMr8pKn/axeSVeC7brmNs/Oum
zdc5db9y0Y4H4jHAL2pyiFyArP7oVwcd9q310rflchcJzh1CnkRnekqsp6byJ4ri
rUlERpDTsIwkZXLldgWRbxvY3htMHJ4DxVez3rGkh9S16SEyNBGn5huSG3J4/2wj
eu6M2PHsthflQjQt47pTq9qA1fV5zn2gSDtQ4ZP52cMDlwYu/zrm+KJxc0JgaWv7
Xx9YjVisu1FVbvndyS/vygxfkanSTYbIonDbZZpPd+3+tq+1RM4WOI6v0ufVa+ed
YN8g1huvsXWjaFWfhSu1dpL2UDk/nkeheddTJ4S7UOW5j1ezEZaW+Q0zpYqhZDtu
7mxOx+39GzwJQuZJgPTP3OHuvDs4tuwSxSbPLAHiCuXhCk5CJKnpLLrCCGOTurl2
mZDvTYwG+0UE3J84V+7QlYyNJb8QkhFJfcODfhK2MTsCuiMeGcG8nnBiFmCoPxbu
s29hxkZyyharU9W63z8Mv4ggKSnIqUvhc9+vIPDJuWys3qui/7YF80aRtBD/P0LX
rve/SSia1187RIRS7rxU1XUi1CqBkx8/J4iRash8llmS6Gof9mDmdKi5xxT9hqJ+
qbMZXpRH4pEFxll32bJGwLnE7wudx9c9xyglHa//M0VkB0g6PJpktCEVXOq6A13C
h99y4lQlBmvZu7Oh9buxxPSxU0xH72D0ITRrdT3ac1R4VJrWcGtoIvYgjs/ntfhQ
oMMqFQ8Z7V3TOlsdCXOeU9OAylIu+FONHR8bCyvl+Ensiyn3YVQacs2LnlgvCVrw
yX+KQyjXc5IYbTT9CmOkoQ1s8frHjlPMyh2zmBobcoXKWnb7yMVZklAv3FZ/moGP
up6gnHry1BfqNLtW5Az2Yo/Isqfw2KgRoa5GLjIAaQBxnpYTmwhdT1JeBNJR03ng
KjHNEunnOJIbMp7mVCGpvwfnbFTKU52TAqg74zpbOxtYrATWGHzmM1NhoYPcC+xh
YUNBanxc9PiWDkHPCrXOA+1kZPv74PclZEHge7ZDqYZ+h3g2/hOUhRJqoXLlAl6v
gXsihfWvH9+sqToorOgkezyndUhB96Mc1J7G+nhgWzFivhyqL6IKdp1hojYf0ugS
IlikCN6nkFHwFH9gW+j67cLRoC9bWMzPfmF7Iu1afprLD1uEch18tn98xpG1YpQZ
3H8UbU0Nj+JqpdnG08PLXxbz1ydCXPVL9CDoUYuYsia2uegkqsVAmwYW19ZPB7xe
qS2Yeul45RYKcQqWBhn5mPTWbgeku2WdNBehDBI4wDE0UpSK4ZraqJL3AJavwVyc
+m8AFLKrck3sMuasIccj28Wmp5/zo3oeNQdtCvruesXT1BVXH0MtfCI0243+Ntwl
vI2VpLd2DZI7BfKxisqfMPiw4Uj26wsqexwhdHlO3FuYFunSPsCxXFVZzcb74bB5
3jMSEZlYQMuQHlNax4om9OJnCD8xpFJLsdXaPgl5dUJBfkktUCDOg68lpS88ap0i
ztfcUinI+nEG18jlgUyC5ubX3JRCzWnLEQnjQ19NEDgTw/fY8uiB1YGpIa5BdkyN
W7do4uiEQAXeb3gBiHJXs23Q+R22co4uHWlECSTRxBYZpO4HxKF1NZOygQJGgwGx
252msDxi1LC0NN6Ny3nInX0GAPjDBn3TNy3tGGvZeoAqle1/GW0qXKSw2JhbdDuC
CbXRex/1KK8p9uPPBw8J9XssIrjUmIM8q1dqTC2LVx6qjyklb4o/9C2zBX/wR3uS
szhJ4nwG1q6taFlwvm8fIQTgJRL5e3w7N5Qi8ZOd9YAISHaovBGM88Ufw9vx9jFq
ZIR9X5lZJ6T2jdSUxUkiGr4uNn05LZJUj64l7QXqbQv4RwIuGutl08VCEu20bsHv
NdaX24cWoVM8ovpTzMUoWVaxOTueX/PjiNK4jA9nYJwsJeL27rfYA7FOzFHMeP8v
eC1q1JXcIxpLemV2R99aIMgJI1vycPIcVqCdIVzejC3NgP41GcFs3UCkJ0FWZ94F
FjugTHCuk8Ajlvae+PPjDCTH4YDPCkrsfEH1Hksao+B4fBDQL3/F/+GxH3zAKLF7
sBOHCe0A2HNwreBqdW/79bUbRPg+5zBeKWvT0U3aWtoYVC2Vp2dwnMbkhhV2FzoG
qEyYpMTYiH4CMW5Arf7wx1ZB8GPNXFcsR23/IJkRSgeAI4/Xo4B2JesQneDxRjDa
hKNGhTnLvh0XYgPLi8CJjgHbicWDNnkmKNXVssDSmI3lA8+4vpXRo7oUSjpbSFEg
eZrJn2SWESvRAP8/BMLm6OyeWPioVR+dTDhNvNvwOit/7n/44wqeE93+c1S7lKRG
1LGDfZWzlTtMRmdzxVkkCfU5n08FZcfbnNZhUMX50AiicFPFhkqoWIWG5LPDWgm4
3xpEc68MW3ppqS/j6UivL5SPm7ZeFYDQS6lj/xNLzqPBEFui85GeJ9Cq0viTTDzh
qlQ1nBlJVE19nyXeylOfLW5Bp/neE/VUENl8hHPR3cBfMNWliQhJOuwsrqgpHLy0
mnP4PvkqBca+Zlm/G2bbCXHuE9X2fi20HVMS1AXktvKyxgwDaIoQTAiI/+PIS+Ln
Sc0jxUzoiXkF1Va1rtxzE7PQdZI3AqJBTLdN9XZJXpTtePWmN8M/XomjUsQksTbW
kOLA1AsLh5avFpwdwtVE/7n0eMjRiOfaevtE7r8zw/kKSC8AaiyYlX4h2wYvhwcT
e9JWOr+ScSX4pLzJLT0W4sldSyOozlof4rHgjwUAT+E3l+9uocjAoTuJtmoNyq5Z
p/qJPamYMQFMkMN5O+EYflpLmKO+uxhrUHfV1pXBzBhFq2/5pgcSleEGd8CvfvaZ
Hn9zYNTNx69ZsO2GnY0DEAf2kX9uRmeAx+xN8jJQNfLUP784aUrPrEO5iCj7VRWy
Uoj2sgHi5tknrb9VsuQUHvvClZWPmJ62oE9/n9o4VjbinUAKdmjg8ufoEARQZvzs
PIbNIAIbfab8YFbuMbIe8MNUg0vBzw1XislxUW4JwJWL6no9b6Z9sJ2CcArG9YGE
b2sZmm6TtKrVVy+ojFr2Z0I/P+b8yVRKrTJnAcCAxwNHjtRNfNXgea3xG8w2rP2o
hRagdumgpydpkZo0dE4XSYYSR5lC2nwsKS3b6xmVYIOnJXZ2YX7K/FRL7XIrAnyR
r6k41xN9ctQhmEVi8f01RreTCL0VN90fzodD1wqW5/OAZu8fM520RoMofqstW1G2
NJb9CmYrQPVOXz1eAwZZkwvqtRag+IfPgR1GNJFJlymUYtK/FxGIMsyV/AhnSquv
XsWh7segtntU6+CP92D+JIjTW5cPFIfW/cxFytNqfabcCsm7+peVR5KMrPhnYPxA
3P11yUkZz2Z1dW3qGG09NB66Kcw4/sCbDPzhk6VJcArn39GRET+qqsB/sYiL8VPV
nW4vPe3pPSh2+W0r4txhFOuAUl3RL2v8pYFouTLjU1MbRLN5TJb95eQdrcHlN2SG
/4XMeSIf4Y2NEjJ7Ici/FtyKv4e8vzWq3I9djRdwSqGUU/56V4pPVdrXH41BrCn3
SasS9Rv2D1uB+qHU9KI9OqGITnRnHpkv/pXmj+t8nqCiybER/w2PCdlHBpEtYgsr
ruxTEO6jRJsb5zgny7GAwwTf9+wOUI5LzQ/qxjveM214EI399jnlY1NBDbe8tUVT
cAtE635WqBrf2RXxKn2x2+pmN2k7bu6szmb8JwX3K+ZRJ8wTapIJ5QrvQ8RRODsq
EXemRU16q49Y0eoar0rByZzEWI5U/NlARcPUxdctD38UwNgHlkbcFvNDg25wgHvK
wsIoSz4yjCqJjIMEQ5kX2rL5M5V3ku57uT/TRC8Z4OaFG0Gz1K1ytsX6Orc59arx
0NvwN7VdLh+2XIDlrhq05E5awHsimDulRzZqpFf7r+Y6fFZpshnMEyxMNRaGTL7W
SdcBetuADnBhKH2WRs+GH5/JcHrsiCiU5fwwIs2Pa5o7GVq3EOw9sfTD0pLalCXl
rlxAXEwBSH8QprfP43ix95HQLQTKo8L5br037FHauzZNU4STEfZ8/iAtkkm9WG7V
uHibiADzS4hjYgCUuPQybC4M4joiBAce8pNJ7APna3Fqun68iVuyj1Q8ouYhIl68
fQ+X0G5gxTPppk/m1UXaMqbXqn51NCtqKakqM9Dxtv68ad6tA71aw4mnDvWb1ruQ
/qJ8nihCS9OM/Lpzml4b9rvndw31r6h7wcDwQvDbKAJOlNxfXQc+VpOM1Q1GmZkh
y24sK0JumtknY3W3ufzqwBy+mHvizaZ4G/+nMLDaCtkwQe7KSb0OfPME56YHH/ZV
ouKRDGeofSKsDVeniOUyQe+VK7Df30BZnKmkUIfm/x3cwrskFYokSyJqAJogFOHs
FlZGH7wHkg9QUCExNfhNwWO3LHwmGfYbGh+EwTSVCQ+ibPV5WVTw8yk+AWqWpljR
egU44/y5+rP5yHNOYlpaQUFgUlq3uQgsWfExDdyMml7ArQZNqP8GsV+U+hHKx7X4
x74HZgI2YZ60qh9Foz9FoGwxJs8Y6INN8odPHwQXu+p3pKM1VKgJokfjkKkGWpj5
FAFJQqPeKug/HCDlhBySwWPSBu1Tf5mjdM2MZL6EQXKgp6q6KTODSqYS0xUSV5Y1
O357tMlJqxtOVU3pV7qM37c7c00nnL4EyhtM1ZUnPdjaAX2tFT7oJWmx9rdmvjVD
HN/mc1EXzXXWl3a71bwMB2zZbx3PvFFutkooYpM4shqlSjBqgZfH17TUWS0TpvJp
f5/QzTah9F4CU8J9krHazKzC7rMJpg/kLfPwpYUIolzW6ZAeuQAes/sf9bKVg8Nk
YHkUUJEgFaD0JFfl6Ppb3ErrahonkVOVqwyGLIB2/ikUS3q5wGBRvXMXQY25qTtb
IM5TRUD358e95yEeJrHRuiWcFVS2xDGWAR0yoOPuO2HMM/M17HlXHkRMc9RnO308
Q/0KknQEJz0CBBF5+tVzIC8+DYanBvktrrjVATpIUXpjC+PF94k66GBRPS0fjHw6
dwyKzFbD7RwYSuh11oI8A5oooxVTBjyM3lDZ76d7E4vTB+u9nGTnZbCF03L1PHTi
oHc+Ea8yf0+OYlVX5SyZxJNIsm8TqTqCYao2jzsMoAtLCzghTWmpcJOhbgqns4KZ
tK/nvj4B6e1BaWvdQhyGXebLEEC67DzNYsYWYzis+NrO1opAv0Pb+bbj5dVY/tVz
YKgf7JEqT3MgkUxcWfEa7C4cvFEv4ue1tvkhgwtybL7cFGecn4QajJ6FNtZW/Uej
Wgvq2vqjYoqBYEBkqUdOgDYRJP0ZtfgkfOcg49soljg+wsvGCMkSrKX2cNuzgszE
PDX1xOVZwHHuSbkVtNmztCxX1+2BJ+uEGwAJSzT+a/ocijJH/jkm04MtvDWaa8h1
snSNLmXrVGCqhHSxeQLDeP7GJ7kuDyJrfKaXkKrOZ/BpLU6q450dUaCpFOgUnkuK
m1GAYOkMwXlviQa4Z4WZeLjwsL/49ZJ5XaihgmvQ5tcpbGcLOdCnZX97HusEvoYY
cZnG9AQyWrWGLn5xHCKWdKYG1Rca/cDjdTI+nz2WyvKkiNQwpIxx0wJF8SbV8WE4
mF6IZtzIxjda84PAoWAm51ekVEArgs2sCAWdIf5aJY+yCs05Amjj1nQK78pKz/ju
9l237RlrFEKyo9AU6h0jQ5VZ0dG1Slun5CcvbMUNWEeKicHYjAdOjSzv4uUo6Cw2
8G8Gq6OUNuPFOCWppb5FPrihWp/OmZ0NmzEHVoLtrj3PZ9zWn9w4gZ5QRR6zXaxz
nu/lBR6gs3Ud58VSEmbtyWtkv4b379642XfhhBlBuuYdHW5dbrUTGW+ieUtMkQHW
WFxdp22M1iO+aKwOEbx9mB6XlwVj7hZ4gM3QTbR2JrL7meNVD38e6BKnecWwR7x0
16vD1OKVIZPuF5ovFGd61Q+44D4o3SoX7DoDGWiTbUrNQ15UUCZICZCbpxCyBj0w
ys9fzdR6TI2d2hX22ABSAPt0+d/HStTBIK84f/XYQ+LN+DDfQL/gLl+9duCeOy8/
ladLKXNL4ACYRWpoVkZf0qgfUrusbgtb9RSPof8B5nmh5J2Ho/7oV2ZdZ1GHGpIV
Xy0sfCOphSEbljBJLKgiTT6pEh360kRswhtb/c1fHr38xX2sahFFk4SbplI1Uo7w
7ImMlPzcv6PoKnReY8QVo8YgQkkyhF7+C2IllfRTdqKkEneR4782QNc3Fq1domXP
BuOharmPLmfa04ZY9s9Ul+DZmARG2WcP2LOV4o8vWfOj2yvN8xckJ6ZUpdIjz01q
p8J6qTPBwKOt09kN6WIKQ3BryNJFOeZF2sv/qnjM/RfhEWiB7DPN27hPouYKn1WZ
99LMNeOv1iDXlL+4nT3zXKFQfBWNuQrhaYdEf4t9tBwIrMj1qVlOPEnvRbHCzMjI
wGg7BA1haTMpGkdGTVE/V2SkBkg7mMWongu7zfPFlIRglHbVDbMlV7YvGpCY+mtL
UZt0ilqHMGURQg8qJ+dlf2s92peulz/L1wK4aJDZWi8cpMPTs2QaAymBqt31PASd
sV1R7GhrMtgtvd5UppBl71HBnpWNwTE99yQgB3e6xxHlRIkRz8qSaM0W9blHpOa9
FAgqE7CqvaKPjVrGgHtmqilQuUlWA8MMuIU3PceqmdemcyERsgor8FrsoTrWxZCC
iMX3ZsyuownXrjNqFNAYhk5ze9AeB3nELRWVHPQpjcwSRGTlj1lsK+RJ80xNr5So
QjuVLNR73SOigzErsJFwC5T8Sbzsp+lr2Iw+bZ5Av9Zn0uW2tUVAXFDRNDsggr8+
veld24qVw8Zlwz8e7GzKh4KSp6D8yY11yedsVNwLOtHRuDxT3hsl9JCNx3J7bWeF
7JQpPDomDLSyFwLqU7FUaTeTrqZnzBmvaDg1n7Nx1GTbr6hnFDzufweD6Y9v4H+o
o8YAY3vHVJT62+l1D7CYysJZnr0MFuHp6efOEdYLD1SGWS5xqUUOmz2GAu6VBbaN
nAYKHMPuO2rKLDtrHA/76DN+guHTE1gV+VR3H0hxEh06RH5QdoOHRhnQyTG2cPFB
J5y/sHM++eiIxbTYp7LtkgSHI9/T8gvC30XslhsZdHGWyJeawrbB38w31rO+5diw
nEWdlibyd76lCoaQjwvq8x8hFU87K3Vd6XNHn1X6s4d+7bGOMZbFrknEV4oaUHW0
kmEMo7jWK4fu7ufGp3I3iYNxxHRSWQ+WPAeYZ8+aAKdz2xiT+4VtN9N/5RAIQnc+
iCXDQ/DDB6Eo8NKh8skCsOCnjopiFBcW82P+jFkp7qxSPlTArTkU3AV9Vbr+Qbij
ArKaIhYYy1KSXupReHQuI28/xPDtlV0ndRFSMh933ycsgS0BSKTy2zpSp/ugIvNZ
itFzNqbPzvM61zDZB+kJaz8bgubM3H5Ar9A9QzK2r2+/XCLmqo/PKQONQ8Erc45F
eRkTzVlivh/uPDfTFlXLLNkn7S6zATKpI5JiuqZLZtipI3bX8as/EmsbIzqC3fOF
1rjoFNEI/K+JTH02vl9TPNsKzx/tmVZpKfCebXiVO4aPQv1qhcIL4yivekORrSmE
2JEcMf37tzxRbtg9jYio2QXs4xF/E5PfGDsAfOEI25RAEWI/9SsDicu2AFJVCmf0
tB+EtnmCyvW3IKgmVZbymHVoqT962MhYHNmt6DO5k0hYEJZa5stt9f3RpPtPYITx
j9AYCmQ0vt/8T5Yonca8YZTfeg+ixOkzB8Pdd9yLCSGwGCum9d1995tcWKHeypQc
q2huAGPd9uhcwH7aYShMbNlZlsW0Qs+u93iIAn1ru5Kipo7gKTbBA69jJu2sFwnK
zfhu9hywt24m0O+rGW2yxmnsZiOgtMZBaWVFdtgycRyKlyDSCgNTf+242iCLmigb
sOAmPwhTVDQ/j+ZD2kY4NCCU3G1ur+3EUybwqZPAcN8lLZHHfiU7ZoNX5PEzAlpk
FcPBNbdRzdkCT8Ku07kuieRuUnUd4t6Ps9zVAH074+7TQ9wVm6mxuuYAkDX1mfqk
uI5Ws/XcEcXf4TYKypk3WoePb/lHp6REtPqyoGJ57U4f1WCwdJLzFALKg4gPmiZU
cAr/e+SCeN+zI/SEBSK3Avbpfp6EHdsJktUDYJXOK4sjrzwawgCEEw8kX8PygHfT
DnTbGROB3gO37eUDD2pEULUS6n5nBTnzVxvtgDGpPClAtgx8fe28FTbpTYq0TfiM
3xOtOHby0IRmBjc4ACOzfjtKchQvaAlYT1TeGC+JvnE1/k+HZWJutBN6CUey5fNp
9lYIF68Avv04mU68sgZlJ4SbfqE3SnMTMyX38UZMhoqyDhj6CIDRDyrouRyKcgFf
NIUfRTEwgqsd+6l5rbryreW5M0SY9cH9JDYKDmTau7A+pgvA/4z9JQmoz3vxA7LR
IO5URwe+WUPfpaplx/wFEcyhHRKalg/xVYtSMNCZPEkwQbcd3HJQwYCyuFY5rRW/
fB15j0d+J4qmiZGLrIT2i77V//L9rEX7I2XJ4MXx9sz3Idid6R88vdC5f2oZlU0G
zjT2B6MFYihMFnGR+ZdqNz3g9v//XARa3XFm1JwdJzUS2MN2aezEU1MNuq35fFrm
f4wwrDpKxyIbYm8j+NwgdJ8+/6XlA2qq8nBptHyy94VyiM4YhwkL4yl6N86mYiSL
hgYbQya29dcKWDzVFai4Z1D97e7PhpI+LAKPDCaORnM3i5SZsEfIJlOwXAKjiyC7
EA0ap1TU14SoNHV2aoYq8hykaLFcKnQXfDN1pNFqLxEHl6AUhl+eKZ1cuPoJec3c
lt8kdMy33R8ZP+J7u+CO8D25bLH5x4mJgbaTjzTpu3LxKZdv6uxNFPX2kUU8LTn+
Ge8+ggQxisOjy+hBWqJTDkkFM+3e7GtbcuPTGpPHfAZGsRFWBUnQgzHjmQs0XpnJ
PdoqUGZ5evVHHWwjpGS5O7QRq6N+taH1Rr2nMTyxxB2y2oSImfXMi84i5eCBt8nd
7ytWX4Tsl1wBo8FYDUjRllz0Yq58sE81vRLmr6SeohofaAlqVWFrUo4TuGiSvYGC
GozPyHfkHaGghW0q/QD0dOuWkxyRn0ay0aRGEUBX6aDZ3plpT8O2X8dWFfnu+jcj
WAzX/gyM9gIzXRssw/HlwQtHJiwhjNWmLkVf72rZxVo1Ti1yaWOyU7tJdsJMgjyY
EODMZe+tV75VfLTte3Ex6nCpTfFCi/JeJ9Z6UeGWUbHsUEYduFfHso6MV7/LVjaW
iMOapcG7fOoVm6pkLGYXfWd2lD1xzK+ze7tl4mVUpksDzPXkRtRlA3E46otC3yOw
mhKQAkAMwdlEAi/ZXd3xtGeR2G4ZXW1hLElW8Ah39Q045vxDC0gGOlB6YvpUs9cN
2STLXiArJRRuSic7YHqOqeuPLHcLJja4Ad58QyQUVTBzFLmxVbBLk1xvMAtf4yfx
2H0XpqUntwBPuMTs9OAZe3gALQg+AvYNtqzKuBESaW/XdTX4wXS+E2Ipl0UDeUtX
4lr0hrzyMf7lcaBpfYfnIHw+BultBzO+1s1sEmGZihDyv/GZGD84ZQPwRO30b15R
uVLBIpe3Pqk21wvhvakarMJR95bWDbFjr1wCBlCfJkYFQouC7jtmOwAxErl+25tt
HUCtKbt8KbqSBLW9XG9I2+xx24SOzxmE7JusyBWNeRr9ZIcwSecnbNyPaB1vIMnE
BM4M08bN5FlIcoGc4KPrdCrntdV2DDejE0n7DFVH2fqB/fLftMVAMDSa1qQYYd7z
snqHeaXv6sT6P8MDbtxpOYKMAlkJwmxphgtS32ODtOWRP1nooI3jtlOVGd+KTOfY
+M+4Yz086qStko+Z0TQPN2jJf0nXczZ7VDyNVVuNjpiPNkTXCn3gfTX9l6DlOjFQ
+lwVyj+P0XaDOyQ35a9fi0eg6VHcBL7Z2cQSXx847IsJZw/DFIGmiwnrp73Up2N9
yjn/FAWL05Wv+9R+RQZU7yfenDUDkO556iT7lUx3TUXMv/mjJeVtSwQIpjq5Jsl/
OAZobD8Qfs2HWocNyVQQWlzlxgxAbk8+TC/XkYU6bk6OLNMuOBDLUOhrVL3Gccba
YveXXxfN67zOpfUh6noP2rBJxJThz703DxktDxdNdpFfV/Mph3+iMCPP5rhQEY9n
eIRUc7kZKBQFkX+iHu2tmA9X768AxAgOztRgLeGL/dkURkVTfegf9/hA5Zyp2ijF
r0lrztrulCQum/cHQBces2hNBBXKBet9Jn5DxCuWOW5mpCkxRr9EyNUM2HC8BGsC
1JNENfJv/v2oElNqh0AhVhmp8I2omLuYH45uOZSRcFX4mo2xCU0lPQSgsHAZz5Ko
J7i+E34pgqH9eC70tgHL3oBdWzWrbnYb94fqK8qogD0zzCmoFt/bNGkFh+a1l533
DTMduWyk8CVMfCvcixlgiUQF5Z8w6jY4r9KxUqvWTnsd/uxW/C64tCv4V2Xl8XjJ
E5mcHuiADPTo2brY6BJlaIdq6xA+osXsQUBQcoPHw+reRaF8Dn5wM+oqDi28REbh
nYDgzWfkrI1nUWrhsxyNNKfIfl8HzkIneVx5yXO4IBMCxM7hcaKBo9McWHVDNR6P
UrT90hoz34iqA37CrYo1afdJU5vsA+gtb3RBJXuXM+2ldXvEIfmQIJ2AP2qN0anx
Ex8bLySUP5wv5rbZeott/M4+c8Hzl7z/xZdjOxvErFGukz57kkqen1rMsSHOP7/1
U3egpNJyIRsDQZHdsNgfGf0QxTuDPh1er5YPvRdNBhgNmPnOh0d8TN5ODpy1VMIA
Jj7Qn+WQCBxLDrPEUud1kFSG9DsrSZbPY1uA+lppTeOKfgeUdhL/8m/UqmKYElJN
vEKDJew9qtVFoN1K/97fekpUaq8lL7MOr+78/2+RmPyZEAeQ7UIFSb1cjwACLOb1
1ifCW1yi8XpDSvxCXEPw4VOGdbSO0HYJU7zT8eLaQEj1KyrU+O95z4Td6QzL7G/j
p6+sI25lbgF715/77Ptaar/gRef6hQXM7sJTpArM+haw5S23WRKuINdcXiXXvgr0
EWXVOZ0yuKpZDw+sE40VKE1cE1smPAcNYHx0jnAfOcvJULBRYZ6WjdaSeQ2C8Sxv
I/iApnsHX+rWjUfsh76BVydYUoHY3EEjIOKv7sndIiYSREyR3NTh5pXS8ZHh45PQ
Ud6oIYte2XXfPNqHI2J6EOzW0oTuGM6p4gUX6k5/tP42LehDWWTEOrIhfgwnQF9s
MPzZLLDsHa2LlfQ4R+oidjlzVqvju+rQyF/ZvqKt9DG5ax2z6mkAknpiCPLLHiTt
0eDuBRw4XM5cc+nC7AcHyViYjg8q2EXFu8lrX6fAzoJuVN8/PQ7xWQ3agKcapNAs
0TDDiwFKNpJAIim3AwLZy1Wc1ymGUlGve5Jz1AaStCWCOFMAYayPIS3yW1TbHzqq
9+5wD4bAHz6yzup45uKOhBsIBsNReD9mu6a9nDaiZFL5QVJ+0lU30f2Tw3T2qNsS
SCqsMPj69ItQye0gSZq4gBCMDor3bzmv15Ojijd0JiSXuLAaKQOayEXOXaDkLRaV
LAiLGdR4K9B5n/YU6aT7Jp2D2xE5NBELlZLfzajhQedR0VRVsSehtHazjvmwR0Lk
PCz8146qLf7jNQVEHp1XkqUYc4YxrqG8MlgF5VcADXdzuiw7nysGJBbl3KxC0X3k
zzvqqT7kXYwAgXkeJqRIr8jiX/K3SF6DILWGNXEyHggCZ+md5lWMW05m7FuhuM2v
qjaV+6JfjA5s5BzbxHKyFRe1QWg9W5IANYnrrJkcAszmXIlrR5qcAXX0id98pWVR
g1r5NCBO0ZokL7S/zQncQylvJ8xneoatThd+l6LWhPYqIQOxZ1GDZn0lHd0YMbcJ
/fl3N42XyeEu7N0T5J+wNJhLqNeCsg4odUmeRvB/nDyN6uvoVAnJcK/ghsGaRPNm
mSnwybZ9BNV3DRxyXAi4mSqXdayjxWgmyEyqUThcVktLp9yTn+k3dehCwRW1tZCT
TBEI9IxNrGY7lHcvvE7+fGsbRObnzangL+Eur5xs+fk/q58c5+OG7TGFZbc0g7aE
9pAOxFns2H0U4QdML9mOg/spZ/gnyvDLVXPvde1GifXOplncE3MecCLE7X4PCfSF
NiRh39w9f9VMWR5wsrPz2LZJXwLrwn85MR/Oh4Iq09/SDXYR/sXQWqpKzRuy56r7
ZaWsPYJdBgYBkjCade2bLy+j47r+K9Z2QEvA71VlY/J20ofU6e2KbBeUb8Xs7jHF
zU3GI231PQ6H0yjDyXcGN2Stv4ECGPfbbnPJii8TYMX8WxV6VV0OlN6syEffDTqr
A9mXduJHYbbwTG+u8q8dMDS9uMXdnB9zJ8EopJsOU2szlKsQeGvty2DN8aVoNHQ9
IHdMC4xBFylNuSMr8rQyqcykRt+36uFS5KLvK2qoyjheuGs28cYqTxN7kGqiFfa7
rTjV2W57ptZ6dooJ01U+ByswHLlYLLpYaIkiIahFT5ACG1UcfUwcMQzdB8xu0kDq
0MYvYQeRjFHc1mmrBCgcgaHj/npWPxIGood4No9fgB3DpKvJRzUBKcnHD6SGKzzo
k9uZTJzU4lKhxPFFS2vHFTXiNRF9F+1ld9givAls6EohdOIb2syh5crydDsjyhnv
sieUWRAfS/MfpzQoHonlVP/oqcASnZJDAH2+kAAbYAT+x8elKFwz3VKtIuNC2WHC
BOIzdd4YQwmZQM9C9uRmj1Y9tBR9Qt/UY3Zr+xkhHuIM15cEeyj87iKJjyxIVql2
07Tcjfzmg8lGPz6XudyHjvLBC2BHd/9Vs69A6z4oRdciKKBu3KMj7oDUeGj0gBij
uSCWe0a6/4YfI/ARfzDGVlOwlzDCeyJ6tMfSJ9dkDvz5Mwrpv0W0FNaN8QGk09Ip
P+GumUTtmPsyNLwr289oxMh5GSLNPfQHj030ZquZMSqG/7S+++GqmZMfymUhTRLM
w+WI4R0F/4moADi3syWnZK6ZzOQhRdiDAzQeLuG1sH5ovHwAf8VYwwnZZzxR3Rdj
bpa1D2U90q9ebAhcwDi+LgQgh6lSPwBxbOW7EvAEnaCFxsHyjz0f5vFGBjgj3+Sn
ApEdA0Lpj5bTCnXj7T+TH6avN3iKqf2V925SdttNObdZA03MK6B4teiaHbdR64T1
vKYKbvOrfmh7QxA2r60GWa/MCoQtSywf3Z/nMJt7Oa9Gk1bVAtKoHd88Ouug3Ck0
IoVclpggJzoKfa36MhTsaYZaIWKJW+q3a7nhQ+4JeQYJBweKeKIuX7yZuaJ0JDC3
DUJLUfL78z+l6LG0jSC5cdZfRQ7DRnnPhpBsP/snp45GE2DZIfVzTjcG7QHJXft/
FpODMN/n4C9UOhql9vbE3ZGGkH7HFw3ywjoGFpY9SsS72VdYIWduocxs2ib3VWut
/QcIeIlmejUAA09Bg5OOce81Awf+RyiCo4O9TafZFhqo9aWr4kgljcwsv09xzfq3
PdpC3qXpu5/yvdLtPs7lkz8pYJAij6220vmeymNubinBE49mlv0tJ1OsSBwfvsQt
wsd+CyVLjN4Pzaai9f560ZkEh8/z4Cm75I8NIQS5CP5zd277IegPAoZQ+u3BIo5T
IT/N4Df1yDZ4gUB80EsIBNWlzV9JVneGkEG6oDUS9PuP9KfuzallUb+vBuLrJGxC
umfHi2w9Ucw0C1QbzEyz0qPya9hbMS+DvXuNVJOZ96hZjL6grxrciANXi+yGf/hB
eNc6cArcvHmtfeQf77CLaNCPBe2AIsK5vzk8lDfa1snnyHMmxQF//emrBLpufcQ9
B2Owh9niUAK/PaBVzyEYTV0AqXdZW7ftvY9rE9UAGx+3f1rzGW6atEOropP8H9PM
y0f30gxkqDgVke8DVANaox6PpnmQsgh6XEH2z5l2q6EX1tICaPzy8jsqfrIBxT3T
qwAK69RZ/BhzAgAQmWSw2Q+Ex60lf6IIX4aU5x4sRku+ASDtd/Lx7MY6k6qcBdD2
TEpiHUOPwqRLzZSzDSGn0KMbT9yk4PprU0HIkGqSLzhQoKmWKZRNBlbH7Y2eUexU
SLcUivXItKY2G7AtuIXRPU+1iO9U3YadRPspbfLDbJa0BiFhw48+39pf3siwhRS1
RDkaJJ9G9G9+QexEkCDa9fK38dsDmStaIjgF5xf4JSMwGBAybeU2lJt8td8I+1T3
84/eh3CgvU0XiNrAVGyffi2rt/BqqEw92vy/jWPe9RVxPdhCSZ79HQndFOSlRAYX
2kcL+CVH/cTujHvyP+rxQXPmq7Z6gIEmvdEBnjjvKWRHUYBs5vvAtr84j2AC1SqC
lgkxSzSv65wWqs444PyPeyWYLyGSd04e9sPmQRLOt+cBzQuqDaX8SKB23gt0gVWu
ZMhCJ5d5SpWWwfstl0lTEFKje6Jx3bHvKhpQ6WE9SvxVxlNnr0NfY4rNjUyW3QH8
QmwdVS53rqXuLF2p/+nzLWQLTetnWAei2g8RalLUdT1HeZEfHnRCdFDYHDMY7qF3
dC+A7Pj7kHz2TVY9jb6kFKHMDhhZ3fGEmS1u0Ge7PzjQ9/jHP3V0idsqCkE7gNzY
L/Xq7s4ORvNjY7kxNLtMPNtkYhNAMRbFRp75Z9LxzUjYIrxoPlLt8xL29njqsPjM
NP31ATI+pyArbyyUbQUp0ZDF9cb+V3e+ICH77GJTozV1xPjw5sW1QPzR3Mp1YgHK
XFuMSNRwIGmJzQd6PAFFDPfvMIgesI/8qkdLBNferwjpWknAuuLUeTSj04V9fS+B
P9bImqtJHwvnuFsH2DEI5fiaOVnUVfeqR2xRM2GfHZa4WNHV6nRcekPd7/2TSRLU
dMKDz+hJStqeQoyqJ9VWrrnYHtEMmPGtYB/n2CA91IFhxxB4DjTH2RPTP1ROybXN
rg93pXCgYSjvD/h+09LdSA/TqTkyHFY7xuS9awVF2XEaSoFRb77AY5sF2Ed49sYU
Mg7ITj/A55qFpMmg4dfo2/FXM/mJBVaaM3qaEjqlcjxfiKFm/jvwUMO2DhPHMjXF
V1/91Po6MqiRxOKga2jEnnVcwXZH/aSwxVjwJxfCEqBKqn8KMoHUuHv83Sv+IEII
uEzCKD0c958mNQGtghO/UmiC1mHLALrLuRxvfT9UWsW+PpaVP7sUwfIdYpWFnME4
gDT27nQexXMYST8cWRi8TAiZxTHST1uULYrLyhOs083gmYwf9acxLl560TauwAJA
0SwsgdJDPSyiEUFPmokMwKDOKbnyM2eiNVXhjE+aKfR0znoncxPp34ypZyUGXPyw
hJ5ZPIAu34SUrAxL2RGQydy/G8w/HKf90C9PUyGPaUR/r+XUvpy9YH1O/mYVUV5M
PUXOu5Jy10TjguY9tsrJw9T1A/3x9qXb4wl7z6XzGt+an8DhasOzyqxzbY5dYVSz
NuVhvJcvWvi61F31ox+PZ6XXO62SRlu8rgZLSI/le0YNSlQMrvSu3ri4qSuEjamX
L3O5IltiXEeUzd4L+x16PgmDWM7vxqdjsokxkvCXNyp0j+IH1BZE1X+EtYqvbwf1
u9N+Ndu2Mk0JzQwqDzRQji80/jO9H1SucGIUybix6Cemtj1d/R9H6+g+tRMW5G19
kEqE4sOoG+l3JWfe2esoi7qm8P4hR5iAGLTBCkjG0dJKl3k2pwx/H5pSO5qqZi30
8dBZlKM7IidKULZogfzOoT8ALlJ8iqsVRWdEPafPE1zjhkbDlR+AytaQCOs7rQrG
dJ0TZLGcB4bBQbYc6qMa1DRroWeZ7uMEx9sY2F73mdaYZ6Y2FLmEBkpzMTkvSAz4
uyBu4HcMI3hMCq+zOZXm7n8h9VBCfiA5CgMP33n6CY7dzsxx0Zr8DNYTt1Vc2jop
UXOK7HoksRCzxzasKefWbyBtyWp3A5b0Cl2YOBctxsNS0J8/KOIsfk2/uNzSzv9B
rTpHP+H4tG9hgjdhR5Za2OW7IjASIBJ4HPWdZfCRkSGs23/sKZvV0CZAEXJJb5Hm
b43q/QQClsCYMmKioo6UxobruBeUA+qpgafhtlRfL/upmln0A/TripimUotLSbOV
QsTA/57Y0Io5gbtLx+B6H1jZXErqXY+ZoaBsbt/zCPw2rC+6zweXFfnnLYU+BUvd
+ZvXF0+DJtse5rLtenmxaXKHn0ltacseHgRjJOOANVNBYmt02meq25FhrboQDAYl
5/Gw4zojxbLn0vMMc+HkFJZu386SaZu8MNh1MIOSk0ZrK/lPFxR1VRhOYWnX0tD+
dPult/0mPL3OJx/KE08ktBUCEfZ7v9BHXAnhtFpEq/LEfE8XesPl+8bFfelq7vO6
aW9h9kuy20ly4ARoU+aS11i9gjnUiOtx21VMuSiMjHwHc1RqptJ+o0W6q7SclalZ
Dz5XZC5UK80UWAbCAAn7Djq+noTIfyJiSX91ArU4lHrTLD5pqQkdVZrJ2Yz6eSFY
OgfV3iaIa4USQgHkTQAkvQ6OXoG/94G5NT0X3ZfvRx9ph+pFcJuHgr3myKDEFUY3
7KowO+BNYhBOxBwR7gFFGpKhlBxJLGODXcYlroZ0Rmzl1rQmLZqTV3RKDty/exy1
HanpZbabkx0K+EieEjKzK5d7P2zPzYuiX/HIROTkHK0pV9ebcUu7FrWBLSdFd5fM
BNc+k9RVpI0qW/AU31uXWvU5XfEpF6iX812pdjpxR7fsj8u/9MHbnNItrzLHOhA1
DbFAH9Hy7GKPhvvMvBrG00jtMUaDIzFdZfADWBGbGuucP4uzAPMyuhTF2s74Ii5L
ewgN4WbR32jBKuWhGZqLC+ZTP+MFuS/NUwGewpqCdFKedkDM/bOwSNxj4+intzxd
QCDpNWrMla2EL+stWqvf0YODZwsM3XiZezqmo03zL6/xuChldpdPTI8VIRVHQ8jx
7SJ0QK9aFF6xVZucDoLWRetZOJVA9bm66F01c8vEmVXkfXwejeSOG9Gn+YeJElk5
6/TLO8Qsl12xRpHhnGmxiBUAl11sqislKVNJFv5RS7TPzxis8TmJ9ZZq/hJTsssr
0YJVqBsujkI1XfmEUEKYKFLs1eC4N8pEpBZbDfM5c/rqLXN9gl15gcxgs24x/4F4
YlhoTMe0cO0G+X0dOlNvu2RxKRTfKKBF9nWCfjW/8RnD68nylgMAH7xB/YIINEmJ
SvA4pfjujvJL+pBNRkwEd+czc16HyZcACkBM3Zquwk4pxe8JDpGVUqpha6bxOMXc
qOof9CeAAI2lPLGGldv7BvQ49UT+I9ozXt63Qoi3fy0U+wvX3suTb/hD1DWw57kx
owwi5j48zfiKP6QCDSJcARx6XMXLPIGqpaYzCQPNFivxl9j+t/JJ5oyLtdKTn/m2
y3y7C8IzFbPArgssA619eHNAgXSGkAlJiUo+QJ6fMLDzMMRDwYg+grjrNu0fIytD
2+d3dT1NMO0HTLQ4t9ELwP1ZXKNYtZ8dau/cjBzn26BAvdVCUa+OggkvCDUbn5nO
Bft+oxbrQXkaeEeU8LzkPDCaGWuyFai2IysOPZPq+AQAwyeUCz3AF2ugAuHO+crx
WOArwfgRePwENU5PpDyj6qsRqcJYXHjF82xp20Svd+krtz3boPi8rjaZPW5HjF72
xn0r87upfpGBwvu7HsYlYqpGnWCWEwrawFI0Kj3gpy1LkhF1dyaEm5naiG1FQjvR
vWdiE7JqkDW9pc3pvSiAZ3t+0kX4I3vBDyOYxdvLGMoNTgPt+JZJdqKgjoSjNayS
OHBTIanFMuKt13qCpSr8/4HsLhjI/3U9mGoiT7xxTDFTqQ1J4huDYMrhKqxFva9K
YSJrj67RnZ8MSmUgxQeRW/IxTtOAxZVEkwn7SFdsSvH1ERQGirCEnVZkBUupXDst
9YjG6In+QMxU3NfTlg2xescEifmMbFncUjDZEcQo1VpRd/KIid+B4Rl3lTOr/eQm
FWok2M6XdzaqCInQMhDf6G/1NWLAuDJ38lI0GzLkpiY2SEoS3Uq0T2RL6XkS1zsq
8xLWh9hlj9rus4qkRhqmm6jLhEVhS6iX+ZSOhI7PSf5TpoFpNLLRFjNjYBbH36ey
YGvEYtSlAFMMVdKbA0mJpIBespATXnBv5DWjgm6kdi3g8XlVNS66xxPHz9zT1P1I
Rwe/AtVNjfhWlv/Py3i8wBoEx10Mt7DCY9xPRmGL012oyQJB+r2TXXd5i1XJMWmK
msEIVXuxW2qpR7ihnlDmF6FN34yXI3lZwXsLMpZt0r12iiglPK87wddzHung4JH2
l2C3ztHHXWs/zUpLL4ftq+aICViUxBkx74SGG0IeY6VPUjcz/uaB9C/LShIyRAo+
aZxZFuptIHsjzgC7p3f4/HtbseBjXaS4hmKHQ1THXVC6jKFrykKyWSHDHD25MbxP
1EKD1qWKg1oiPB3ieVxAqfVqCRhXhWe+dgYmF45ofP8m0ePP3VyyJkn6ann/Hj3G
vLDoNZsklX4OGdIAzHP/dn6z/u48I55iE8Wfb2grFlpd1DJ0JHRjE3GSq6vxgiOP
nk3lpxKaK5845MlzvSRozq14PSK0eCg6QKo2+CD72SVwm0+2E+JP+2huS6eS6oEu
W3R2P5cmx3vtR7hUzIyohI3SXGbl9gPoDVcOx6Nb0IzZbp3BZIb61mzhiVr1JAlV
0r87+5n1huylf0UV8+snhHLvACs6Ty1Y2+RlltUZ00shcN2wLsbPQG3AgxNKlodS
JO52fi1qSiWWN9oazb+rN4WxEWEwOPCYwYlKE9wlo10rl3bN4l08olY7YPHczYom
tdSRy0ssIAlwa2EvWK3C9PGb2t3GAM50YliJPdCcbEY3nFQi/OWpZLsL14MHsON/
GwDGLLwwvxaCGiw6zZnE3RVbo3CTedJmQ3Gk9mWjs6Mug4snPVwb3vN9W9TWOaAS
FJUmAg+e2Dnac9QImZ3bwDUeXSy+jCd/L3Cw+6T+8Ep9ZyH1rynSjtvNRY/4/tFv
FV+/+8eY3B6cIV0dpL1eMdIa0Kvi6ss6Vze7glb+mB5Dcrg5YWaJPEgdkaqctUoe
Zo1uyr6i6vkGSs3vmdf7+N8cqfjqVmd/BObaXAddtuw738AtF2MdPwm8FIyVW69J
SHWzwRW6NtmDX8sZ+Z71hSaq9sug4+w3un6FirWXsJP+wK3kNhSAG5bIooCAGuW4
qid+rkmyJ5VcufcnA8b7sQ8kgriMSH3nsDlPkbX/Inf45YrnBIO7P+scaJgHKegc
R+YR4QTvPuju87JM/G+IMrqwMwHdUam4tQNMnME7ylcg7Tsx9w7C4g+UgwAqbn4Q
MspIjeUSs41CYokJfO430kgbz2oDJO0rLpqJRfCTCXMz2Kq8vrDU0C5uzJhuaVqz
M2+p89v/4jXL6k/rsZkTuvBeppBQcyAiUPsQSTKiVSpXhnCUtVGV9eHAh5GbGm4M
wouwSszX5DUu5MT44peBHl//wbLus9COQHutn3fzz24rzSZVB+IEY5frAQQWRklJ
nL/NUibvv/mADwbKBlapOxuWcRsj62oGfziahRYPhmf6/YfRmR6fRlRzZsW1QB/4
l0H1rLC+hq46xDLnW4ju3H7TKoEA8F6SHCBx0+VPyY5E7zW6jHTIU6K9EB75Rtcj
gqfAcQnN1A5dScd/nfjM0jjxCZnW8yTqbrCxtEFG/rAPOmRURUuUZjr96ajOKpoa
wLaz8koZtY8VxUce1zFn5syvwUK5xT3zeVX3d7flTTJQUkdSPPb4PgufJ5hzHaBo
GZo9SNpZGfgf7QHhyiueM4wcS62ggCGd0rxfBa4pCuCc7bToalsYLpIf946BXLR8
NcLLoyX3gk1KKWgdCicenz9N4bLSN6pc5ZuWUPf2SxM8WAjZwSPEW9dNUSEl2qzt
f93SXURsazkiY+YBRqaFwesmXz2rHDm7ksf4JTZJBprEdHUmZlSKFkfWymJzkHtJ
6d9rKj0XlxnSSHQ6nSoaRvTtM/AcZy1Jzxze4AXVqK5GcO1iETZxsHypzHDGDCZm
dp+ZH1IO18leJGAVo6yr2wBnLUeX4aRwLSfSx0csrgmEInxQohTJDuS5FEbvi6y4
l1KrySMH2oiLQ/3rh9awLQ34r+oIpSXbe6d8GW7gtu4fiqqP2H6N9H23/TnZKyX6
wl/SmrR4Wp2GjyjtP+A6Rt8pZFRheDR4Ud7mp7MxDMsoc+770g/gulq6ueU9w7Mq
KQipbTVE7n8IC6WWaoGlm2w4iwWrPtHYvMRAchz89u/fUlsiDDLTm7ntOVD+YhFT
7icVCqk6HGiRjfu0PYp1skXooNVKWzLU+3Je522nwo3LhBvPcjPsiIbQ9yLTulvu
W1Ag27KyzLkF1GkHGZ8O7kU8peP7qWRHS2PTTnu8hAfQcAcU2P0HUzESG+olfuyd
fiLL9Mid6meu68Zk3MD8SWnHxL4S4cDIJq8wZ1Kn8Uz1WySc+17fLZodUDXqfurP
R/QCSc33tG2g76cHlOxKN5GEkqTqiW0NU07g8Xvo0QT8x41HVEhL0G85ziU5kGkQ
hpU0ehoea9tIkwpb8mxV2+2FwP7FA6sQkQ8YbvnDsyy1A6teF0OUqToAWrnr1WTU
z/lD/CSi4JU2SGMIhSjDrhE132Sklaspu3OxwonWdHXJ8TwZTHS/kGHUM1x8BDsV
octKreMAJxxWoDnD35yDTLpET5D89+dW7rZ5BU43UNoGYAVk84rK/hCailkUpMPe
eYQH38cOMnm7r2u4dwM/CP05vSDJSPHNPv5ZccZJG4pXF2pCN0Wab3KfFqrHG1st
DKIGmKNK+Jtuncby6YLosJ6USZvfCEdYmdCwSWw/e+W02sfRt7gjeShtwZTrsgkQ
VJt8IgwjgpM+ivRkRL02U3Leted0vzeWAUCe6ZpkTcrVs9+wjHkIuVKpPzHPeu7M
MmvV1qWI4aJGRV/VfHjyCDs0G7WjUjYy7r7+Gs42nvnZgEJ7h25CnL9bE68GRtSB
kp+vfsJTJkIWf5A7owc88TapfQFjLCupNRom3x2zS8F4OKoOTBA+achgUK3RU8ia
JAxx7CKcl+cjcRwIhC2ps0jpDH7zEq+lhNnk2QDrrUPPuau7/qhcdJs3oW3B1xXp
6lg42oTQq6CqKoT4Fr68yyf2NQrrUD2l6dm61js1DOOncSFq0PLKLtSw79iGXkJm
/xUdnw/bzt8dEZ4Tc+tFv+gTCcdvoQF+Pq6DxB7QQ3cq60hn/Q6bunfhNyH47/Tg
FjbgF4mfQ2UOaY3SO88uKIYeggNRFL3whKDUa8dG1M+FLWgQ0FdC0ZgmHKVxZGPl
zAQPNSyUEHNTAvgp8bjdI9gYRvmrNVomeAYsyKPd9o/Fh3E392UJzT/RO2xaN4J4
TmJ8ceC7Rq0TTqmddtv8V7Yxw8VUSAvdZEGHmEVmIjX8ujgdgx9VhrPgHH3VunDq
YUpf/mMGxEN//PCyc7EcLByoT2k4yZSR5Pq+QuomWRrDESOqW2Rv+G+uE/CUH9Q/
xahmpGp41kR6cvgrP3nZ/qhS56X8TUicE2PMlvuKmW/9JUfZDzwzFL/O0GMB5A/o
qZVNgA9HcZx254bpjMou1J83GvFu7ct8RRcgfT8QZ5bNrCZPm7UAOMxSN5coea1v
pr/qjvzmSFqx5nmBfpfoW+GagmyOU5qtYIaUTtqe2yJZBRH4ExnlRuSsWUARcPGV
tbXMWs9KGVwdNPL4eF+szbIxC568YojDwyRoZFocLT9ImVNWpg+cr2lWNatWppZj
TM75YionX3T9AYaKWTzi6TbgmlFqYVHoCFduVbS4+is4wiPQ4Dd0en9rMw+gHDKb
XSGRK0hVNFLvzbq6B9iCuHoKvrBpYjO5L4HjPQdiX+NZZHmOhJc8QM0piD8NTFHM
KHLRpWeLN5SfRI1T+YRKovaKAE2f9w1l9Ya9z7+Boo44N9y51EmJbQzXJsCilIJV
mRDhjaQYT8yXTqu9KS39FPnQ9vHiNJ+i0YFNnaklHmBwFeJ1Ty/QQx2k3YEZHxoQ
KU0W+MHGzXuHqs/bklBBVgkJYngki5GKotVUBemCm38gii69R7yQ99441yICPB3V
ulfZWCnlvwet5hy5sSJQOcahi35HSh1xes2RLOzWfWqHWeFyuCyPkgqZpF5FUFo8
pEAhC/9as/Mm878lZNWNA1y4v8tNePC+pNFbJi605nezR5hJUepE1HkIpsRSI3No
eKE7t+YJzqVshNcWQWIF7s+cYytXwLT+EmvsbPUwaz/6IcMYqn0bqj0fwMgAb45R
M3AA/nPkjrij/5XxJZU2U/7wE4IUhS/EM6hGOUeUxfGQqcj8MYiC4VnGdb07z+wQ
BKEj/6ZQyxbulA8Zxrdp7B0GhljoqsOTOVwj8L3ZV6hLzHNZlld2ZehZsp09vEch
qC2iDVEzWtS0ZAD/gFXt/8dAQFmR+97YolKqEwDpPDcXJJkgI4SszBBe7OrShUvU
VhInXCtxTbCtZAnyyASYSO3CtIsgmF7/e/5n78jNSHYyw8svlovAZ6Xs7dVIc6SN
hmZs4Avjv+Rz801aBvOpGLu5R8V6UCR/1WYXUPcFiJUd8nVScedSBKpmgTlg6bzJ
Z+6NIk5E2atPu/83kECO3EHClJpjdY0Rt7NHjHM7ZV97ENUPYdJU7rKj5OZmeFSt
G2sy5QuT4n2Xq3tIle3spe3tN2q4sL0cKZmN/9jheTmCSqmVX3lddGHmGXD4qQt2
8cZd40I/B8iYu+mBYYBkbMmBlo53+pH7Oez3D9nNOFr7/xyG70yOQeWjh++XJE1T
fRydgzQlSHPv8114t9iUj+z2g981iHZtB5qsDvR8kMu5SwKdh4oiSoV8AahzNGRJ
UgrBc6Q+4U6k40Uws9hl7faiUPGyABqFWJfLJw+eShxRcCwGoVqF53kdyrdWxSow
SDJuGPjaE98BWzxVLQnYEJuTmTrUMKMTKe+Cgr4dnnPfX40NZ+YQ5oQV0+euk99z
YJ9oVTUsQJOJKCQzDX45iRnvaIqN3p3YpKqHTq0Ak4C9Q3GVFZ4nuWPyJoBKA5NO
jP6vRKDFsCseYLKg/iwIsoMDcwC2EK2hcd0ON0qbWSiTQftBckx3HHFz6wde6VFJ
WcK9MpQcq7WTEPKXJa2hcHktLHjTYHM5+0WxKXhzH5bWZIajkBqL/3/4PlFAf7Em
GBiZaj50Crf2HejTKfhTHC2avbMfph0qG59nVmN3T4yoTUOx76SIAviiQ/90LoTG
gvylRfp4hOqUJZGV940Rlx28wOTZyGFWbI7gsxKV77ewqgI7iD3hEA5234c0c/IY
pjCwKVnyPcrBOk+hB3rwfz5NQ14y3hCR4+gHadGVgElDEEXMjy2cgHexkMF6UcAo
oyJhAjioEY+SwcDtpKUtx7nxiAdjCwLXC3JKkOgUora8DloKCao2p759nxjQV/4n
FU2IfPLwg2D/5AcIuoU4UJoj2V83iMWhZFhWBR/f4VvaFMasfkUbXfjGUvWLwxS7
ETjVqNpXk+Tl/Nkfvz1EjymtPm5pSscZ6lMDeo06xaFw/Oj89ZR6n7Pauedg470G
SYXPzDiKa9tbC0nbg9jfZtO2kn1hTcSeBVShqaj1b58Yu7WtH/BG0oRr84y9cKZm
a0mKOh560QxM8SY/15TdW+mpAfphhor9UV7L3vSB5hNUb0SVgjlchChs2pMS8j2L
FMzJSst8R6gwaOOMIEd718sDmCkAweaLkeJbllndUV3L8YKlkVUGuVwwwdrXyytu
bg7botWdLLNBxp0MNQkFq0GYTn6uDn4gMustBthbz5Cp0Okqyk8NQF4qDOyt9CWC
Mf9uZjerof3nSmil0J2eER/X3q6BYyANhkqqObsCNkUTu4sWmfAMly14cpS2EjdW
bbHXWKSFcstzqYQecOj9Ar10RbPilf2IEdz0yHVXtLTGejVGp4IpGAVCFAKxfJQx
T8+/uwc3N3rAroAkA0APuaoME6BBwklG6fym85fKUe8kKKXuyyfaK3j54HqPLQny
RMl1ySDUzk3EtnE34bFGdsQ6Jq9DxtMFhe3k/q3lDax7UU4ErtW3QW5k1BZR7WEw
Vei3Zo7+ZTfNxshzuCaAqAc59Ah0FZv8/+nfE2ohJwSqJKdZFyv65Oj+3jPE/Rk/
a+BdCZO8M8zqaNl3X0lNKOtTJJj1zBxJM4M1Rah7485GnC9gqYx4AHZFKsAm0XeZ
n40/GyTMFR7WD9W/8n0RkRfdIVjjiItiyNMZw+5SSoja9VJKD1pCGHcIHZYYPMzB
N9RxucRK/umiLLm41HVzR4CUVpOuiktaMnSNvRJDMkq1oWUANQFNgZ9yadGt90TP
03yLGWYZnxb6ttqxfh7LpX0FzxR///r86CWM+iwy6R6/FnNDCYZwJsLrhkS3anZx
QBKbr6jl5fWSYxj/QBzlmhDeohIEDYTbdpN0wNHTuv+D3AGK1/ZkQIQIiTaIM6GH
WtrfvHgfj+6OpxRG//gYNAhQsKIVt4vrkReuI/MSW0agjlKDfY7HsR83ig1VpXpq
EVtN8ZRZseg6tQrrAtrQnpwocY6d0GXyf2cVU3Y91RgyEuS/h8TJLquMoKz1Zt5I
LAXu2q5xCryQpwx579V0wsL87dsaQ3HcrCy9T1YEA+tY8zKqbgeLphfPsSmkPwQC
t/BHkFCPhpcPLW1kqwlBGyBItfShhj0BR6XYRF2mQJdqphglJm9fp/4UcppRqTMf
UP0TKHUMAx48qpYcqYMUBDLLhwVY4nzIXcd5yk6CQHbi0XM929I8v9AqOCrVUljS
3w3lH7F1fAuHsrElshDb6kIkwkh543BXIDfBwTDMiaFSZeb+mcq8bNoWNwGSwpwI
N9ITnWdi9Mrb2NrdbC78Tipl1pbl1XimF0mpqLtxV5H2japDMeujI/7xIN1NaQiu
aryI78af6SZ+/rc9nfhl8SX1yzhovZsL8jJrU5YX3i74rDMVeBDn21Zu4QArRH3m
pAuGeQjV+h/Sx8SM6sbaMuVKPGW/basnj5QJq9kPvk92Fs0cFxuGvP1ueBGVlmYx
mDHMn4nj9zinmtw8orXmc/eYVzkE9/qTAcf7WpaoKhn10Tqw/sYU7B599kwNCYR6
96+f54ZzcLWnORafxGC+/+ih179bAn2gvcpLLeEd9HR9oIVqoNnU2q0zPOzBu2lx
0GPu5s6NWOogT0E1qlle16NuuRQCJI+/3tBfKs70Ri5KlM+w9KceAXxE69jO5QSb
pVFatoF/u2RQaImDHQJkwKsjCiRZZ/Yp0T+216QWtlhsY6EyOfoqm1mUIrh3tl6k
gUAwVKOohbWhq9orELjsK+PAGQMOO6hlVFOKeDPoujNrXtdhq0jZPu184MTcxzW7
+jqDqOTkublcOk4eS9ineewVLXG8Wj7/Fs6JoAVceahg8gJ90jfKNmnTGjK5czhM
yAPyiHVnpzZWrCI/c6tGgoCEa9GJmnWUIVTZW3ZWD6jzMI4wefhEg1NDJNlQzJ7h
LDkVc2Z+x++Perke944vNWmNGpkLa9b3rUpjTm+0YQJzsyodw9IDs9/K3Y7kRnek
TBQa6QxzG+BQ7eDe/cz3ooCO6PqFoY2H074VVmC9S+aOpdWLNoMc4fROdeOdBDHv
k76h05CwLMjrJUr1mSxz8Bzzc59JtvJC6iOHqLJ5Rfc0bfFDmJ7BvuOrJ2YFLokT
v+Z1hD22EBu9ZsuLfEaTGvEYxPo0ql8rOP+tjXXpTZCukIC4tHDqoCmyMvRrGDH0
G/3wvHfAs0fQCLTiKeozNgJQpfFwcf+qqV4qiUSB/SGXOK9hYedAOBCPwlG6sXFQ
2b9AGNh8pKh2RvSZM64Nh/ldFWfLt+8GOhxZQlu/fUR32S9rx2VjazQ17FEGUSx1
5/OIfya6T2tEczyT/UlJgGt9XYdSte3NK0DzsZ0mYrIWe+sppGlB+qbxRGYo1S03
2C5qQEODNDHtmhAPZrwI90M5Oi+yqH2K+8/fcoiQdxfjKQbVphyyl5DaXwAq+5Ud
7NVbfDp8yHQJudjBUDEFugsbgG+UdjW/M51LI3U/Myf/b0vnwnf+JuVhMTRW+faQ
1fTPaLy0ErQYqQJdBEVbglMjWGwOiyqaGNWXkjOiPlqPWcy6c4tBT8cnFETnN8+F
xSNfx92DmfG2ohJZkCqUnkOGXCaUldXV3y5QDdWLC+DTLx3I2gTRkMw++qF4lZJS
fIcmVPPH7IjGRkQ8Yi2zWo/ydLGcNPhh51jzjYs2Fb10dUqb/5/q0PbCTfC0AUnB
6rDZ+TUBSrEQQsGLbmBdLOZC3IlXWuKjM51YtaLbRug92J/W2BXuPIJ7kNob+UhN
xF+IN714+SYHK6/zBP3wdkRFQhWv8VeaSWUWkDy4Gd57ieek2GHrELWZltzrluE0
XrXgmCTqkkl9Bz2T/GtVHDE6kHF4zc2HoLYszVeUKC7j5bOOLSAVM+0MSa6YhOqa
QFn57IlWeoXMsbdNapHEqyBlu1ukkHYEjqKJYupbnVAxJY4XhCT75Z3JiDuZ7+0z
KzP/ztfIjjcZWYFqpowVVGRChv5vn0GeA8MzxRqVPTL96h6/9Rzasd+qFA7YiJHn
dBSOloCM7heeWcrFVJbpV6m6C8vKI3Bj6Q7Q9F7zRFLLFJAaxC+Cro5tWqQoQbDW
C1X4rvqUx+SHkyJM9bFS1d7Pjlr8o0gHaU3DHhOop7wDQ5E3H6fFsHDybLi5NEED
pbc1dppIQA+EQ+xIwRuY2VX0/wxINWlTs86u7J+uVIhuPdwrsm5EhHy/2jXPBd0V
kz/JYdmDC3fTGVrm6NaFeOPkk/ULIoUTe38D2vzrXF20I/DE5qHSMAVQnfds33Le
9J8v5NI4ma4hqbU2iXAD8oHJQj3PHTCWe2pM488C5SAuB+7mH0wo0Mb4ksQYmB9W
mlMc5G9PvNSoB+Vv7wGqBGvc8Nx8bMThx7LWoctRZsl4FR7GbxBnCg5hJ7RZuf0L
N89niqiUs/oLW35SgIeB07bpXXBqEY2EtujnK6ZZQAAETXR+gwIdKCdnGY5Jq1hr
eBqfZj0zzoijsiW9QtXc2k3J0soIDEiAdZScZXmPspMQCRosvMzOdK8ecR9R3EB1
gI9gJG4NVKVcsnv2Aq14NfprNCfbpobyxdlokuwzlIyxlbW2ppG/doFUlWBrlr3n
Ww7kXG/4DqZEYG1pIpfiVeyC6wqtlkqVy2Pld8NW2iYwYBvVBaf2taaUaLxopIU+
kiF2+OwUKNpB49mXMzN8+TDoB0Xpl+l1liyk8yCyeIZvp2lb7AiHL2o1Ct447+hI
uxeXMkgKQ/pXJuMX64fnvOg0TyIKx00KKsfXV0ZOfc0aGenRZUII5bPq5jBxih/m
GvVbqS+TJ5dXYa6e1pX5wNG2yeJYdM2C2Jt3dFrTSXJQNG7kxneOLDsURJOQFmJl
+SDF6eHSabB1IMNpGqeTRmuHtkXUZc9bUAq+y3aujQwMV8zgskJPylmD6mqvu2M6
IYoodNT6YYa/RdY64/jRaPiIpAd2BFOumuzkejzATo/+xWtLsggXIe9Rk3Q72nau
pngJsf5FhjrpiF9hvR9OjDGXSz2kA9muPzFq0JwCDnAymwSqWmDBLQbxAY01RW5A
GFcGIGfAdDyF5V0kvlZN3dOnavM1bdnvpxxmF6xAsIjHOb46TTbgZnDic8zV+dOD
yo89hrGPuHCXGEp1JAFdRiGBWjfmPbamAKvAu6BhT5NAF42AoLES07emcNr4/KNo
AVBhCZyt9RFaFjD2zmTazdGPcQ52VkR36HPY9hErk6WwfDTiXFV+MUbGXmgKyCBl
ZoIhm8S34gxr16kGMOXLMBg/nxYAhP7NgrIClm70rie/+miP1o31bPw/XBwD+Cvl
fBmYImdvP7/KttIB0qu2B/PhnQC+tD2wUdW1Se+9w2W95hIo/7BOSnqSikJTSO64
I/4V4HDEzSM9BmjEZr4akomKOLUowKt6ZNbNSvkTRj/nx5+XoVeysLaLKfO/y7vO
YhqW7INeohVOSOjZxAj5mcTsiG5j04z2XioTKqZXIqntobz0HRvyuOe7Zwyu03eR
Pzl18BzHq4tS/L9K8vkm5tZTdcsODVWshzLZ0U3HUlHumSG4N8BeaDqhExx7W0Gj
EDpykVOm0ipKl/7LNIAIN7WVZJ/j/x0lH0/Wgi0l0ya0EXRGgcZQhfEjIQn6RbBY
NnlQwVJ4i3cRFCSlMyX57a2ynijDo1ynYiSFE8hYoM6dArRHakbHQJgobSWn/N/y
HAIRcYyLi/qRuVz3LXflyIAdHEvKEa8mV4bUrMW7HQmPkhwD2HhMIFZoQlnfMX4j
NFlGfyC52J0kUQVMxiBfe48wO7SyOcYDXfo/iUfaDzeFglAauItrrYb0u261P6np
pigLEuJ5xRSXbeZoIHojnfjHGA5NH6elCZsIy4J2wgUGyicquraDV9XfVh8SghkB
qkjc785BwRNzCtojOqEPmXyFSWjAiHPi836fZA2QKY3NJPMmE63nCxwY9K8a2wdC
FhDTIgacm4/QJiwwGb4OqYLgH6PEfIaXld+LLSPuRdJHlWqvppsk59OKWclrYbkT
RR8YklOIy3gAm6vT4ctpkpEGRqDyQZKhp5E8+EOyQApzlonOxf3UsDYI/wNwX1Et
5Nk6yFsITfvBhmrMnEUOp4UP/znGMtuV3xEHyZBOMQhxh13G9NJBii2zSGQrdd/B
JGekPkmG8OW/4O0/yN0Ks7ETvKgG8pfj2BxogPRoi3rvi9tjnvNCqcFiQHAVvmSs
JUYpiEJ6u+t8qqv854T1nwEeu5QJxuLDfjvM38JURwWRF96ofrWwDRpXhX5z3HWz
RssxVr73pKN4OPeb+m1PBxXA6zNdsyhJ6HD4n+upATuWWcvw+3xl74pwxNNprshl
uovuktKr43jBolUvM7cpfDL2pjAJ8FwKfSJt6AigoKUBRkJWkAtzdZXydV8aTifd
KBmWkmU/rusCIqudxbMGapL4abAczOuDqo6sIsBuqBlrqZUvhAbQ43PJjW5RNhkW
9hsIfWGqUpeScsyL6VaXwIbD1pedvDZnAlsCcz6GdTOd13qTfLab7cqypw1vNzg0
kRslIYkhL28SA5MjbMG/sOFvn1a46fBms367mcBc62JNohfr6XWTm+fBXKJX31Ol
uZWXxwptUWqirINzFTSWgTvyqTFP1z46rxLMFYhJ1rEi90lnNHYFLbor7ecw+acV
A/X0VomKBIUKiPrfWFyC3Yy+43lvin03sQjki6SHHmKEigocoIkr8g/rgXFvN0yk
Vi9KNvFhR5ODxxmuJV0i46TWCi9CvCouLG/1cOY/7FYbzqnmYZsATzuKPjpdC3l/
2Jq7+MIFtG2sSZ0zEBLw3z48qIv/sI2d9+dFNzoWGEeZ/JQPIfd8452CTFEFvASm
mVQGwIobIxbrLizlvTFMKw72Vwwh2vytm/blaT+x1uHLTaE0nG5tlDqOAXUfpK0z
Gx8bkj0iewRPeZb/pTxhd8lRHyAWLj8pgla/ertADIqHLUgwxhZrw0gLbpboL95A
qA8xeRB7lQ80NxPRwjJ9Mkwu9H6sZgk8dWWz6/6uuAkbeckxKOtTEjR5OprXk/9M
BR8hjP27Z4xtHI2GaUTKl6s9FomaCtvNVFuZ7JdoyOYEqoa062+AUIgvBPmAoE55
NJZjN5X4VKCJbgCB3wwKOtDclxu7NIDpTkK+iFbl4QYAScOPvyD0sWVP9YIAfyLL
YEKiQrmke61ecDDMeiB2cgDYsCouaAN9ggnXpqk6LfnExRR6jeNucHKt9CYevPgn
KO5xWKspKVwlMuu2Q1v2OzsF8PDpO0PHQr6IlldAffZlqqK62hil/QO5OpIbIggp
yIjczGPVEB7df3nuBeWgcT7NCtHSVwrVG4Y2qm/QRf5+R+beHJCBmEfNhAYVa+Bt
JPAyLLTz02+JCtdzf5B0Mx0dfr7YjsqjN0vTBAVXwN/pqeZqqsPLF+1LwUk8L9e1
HMgxWDe0mNPVtyivqQ4LbiOhobf8xlaXtpVX5uBtRdeP8fIpv4fMo8rclJimUMe/
NwBTCrcc1aGn2HIlazPnFo+VBdkagzD4emNtIm+hRM3gLpcywQ/Yr6W/4/LOftkH
aG1a/i3X25kCPrrVtZ6jiYBLhDYsFr89HP1z0trOF4JLcR07nQl2U7OdUP8/xjEO
N80TZATzAvk2UOfHsbxl9IKm1H4kWNbvBCb89cvYzTvFKFte0JMdlsg4gBJpMJum
xA6bp4c5+ailCDB2L+NWU0akPBjpjDRe32CR/e0CAEnr5gZwbWlpfnFsfCsYc/wr
i/VCklyWwwEhTnwWMk4+3BQ7RvxlhbzmuhR86E5xQC1SM0ZURCPicZEUdHgkF7Er
q+zeTz5AjGmbzzfiUbfulu/YYTnFbixSgngq6+wX0hCVU9Xhh6ouNRkoK0dgrrSV
h+E2SoUN6dKhPpMd5XxRAtx94guKWAf7KC+ANvB3S2WtBHwtTdL1giPCw2Iplsih
TnOd6p+aGMEIkSKZc/GNp3TGhsc8uc3TFqrZaGkaX3cSV7aV2TPWDzdEqFOCcdEe
DQ/biGl8o7jj26CUJ44aIqAp+DrrVPrUPD55S+DxKR3qgpOLUXXBVUar667eQQOJ
h9RP2+fjS/X/gNGJlnh17E4fNIY7kyCbIHPBlTFyYBUgMvChJuUHIJmmVoo/Ehu9
T+jZ1g7zpA1bZZb2vFtBHeNQf18VAQVBi15PS97q4PoPjTlqG4sZMgKj95NffRod
MDkQO38opEMzJaiOohoHR0dxwZ4e37TR2lkSJkWgQSe3R7Z0T2eDK7lFuYnnoF8B
VAjpEn5tOD+1QkgaMOY/pahJAsmu0r6xI5romN4kYk60D3zGXnR3t56+8NIG0J0y
/qRJTxNOoa8MZHekjsMxTzEp1v2bsHuNHYLIfdRAI/706y8PvDnv7jHcm8FB2pHe
O1s0qloemfBdCvT8khwXpgGfNQ1U77AoK5W54wtwvJJKRGastifPeA7fEcNUqzwD
QspA2nxW87FPh0yLkrQMU9x54LopveHIIeKrasYYbqV3XMw9SRV8Wd6wFQpiJji5
O1ZuLOvl8L9EkMal25blgs8shwERFr4gJreJ4TJMhpV+CIvHIOmhEL1S2cWQhRNj
Juy3OCmmgFBeLUk17iGf+OiRb54p+NKvInEfWu7hPOWn92lu926D2xveWuJXto1w
x7mMXPMiJcV6w0gOwDyfs5CgbdekaOQ/EzPrwYcXtM87Z20eBBd24caHXdJVC0RQ
2QEYPnvgcHgwz8xODQa8Z0n3rPETpnrku+7AKYE/QzSUdVdcyfdA4pJbGw5A6Dr4
Ql17znO9TjGGgoCpECt3hOJF+/yro70OJ297oUUo1HEUi9rCdfw1geaHoQNjlbjL
Cy3v56VWlA2q3RkfbToacf0fBoQXNUueg4Zk+YKVWY2BOYDWIfNSYD7sO1FiXzfA
PtolVbKs9kTQVjdHe+gMPmfTtxllYw5oe8OlyXWGkxjYcTx9txfwg8xSTOeOrrIy
RZx8StCrKuJkBD888lIm4e3adF426Ki71yqdedqO0Oar/1HZ4KkdNbCHUA9WK8b/
ckJn6YyIkuQNdA3gC7qT4gwnmtAfayQzSG3ZOxAtaKwZAb5ui16yqZWz2XKLOSZQ
zCfK62ngWTBDzguimJzkaD/vcOB4CqZFtPejGNVpVv53qqEwrJ5kRun39YVxzLc1
T8YqEQNK/lwSz4QZhYe0ln15iff9Ek50m/brE9Z7AXs9XlutUSAy5mjK1Tqp2jdL
7we8qGF0W/vUtMDxKx427rLWoSelX8llR6S5eparnfk4MmqDqLcAbNswSOdtzjTq
XQpjaDo1jc2WsjA0yggD17in8fvzDtMU4xeSI1XEKhSHDaGXNZiF0F7zJSwJWV31
RCbxokOsfHm2YWxFhDaSoT2jdMAEmj1GimjUy0Ek6pHmhp/NT1I7RYZS7PiOeyYk
irr+PDUXn0AxBiBzoEDM/zN/7zgg+CzygtNVeLWnFQlCFckujCJlgTtkJ8TmZI7h
hxFxlzZ1R0JcUl5hmXzzLJD2lUOnn9lXS4DSSrKF/2bXPh1AGGqHL42ms5Qw1fr/
GTM3W+gJN/NM1Wa4NBYUNPnimiiPP4/Amkmc5St3oj9L9LMZ9JnwXgz+sRwh6+D/
nPu33kKsaZSE4a3V9Q6JppuLiGQHqH3JgpByY0TJS6/pvx+bR0fXlCi56Xrfvhyg
NTA8ghIQMmH/Zbbkt45eoYo4siJHPiba+weDi9UIRsUtKXiok7WmKF+vfRCuPIVE
1BiMh1xgnk5GM66oKYFoPQJu15wzDcMkmeVXoJb1TI/1YKGF6ET/TonCTPzTJ3t+
mWtKDzQ6ae0jmSEyaZcwwK7wuXkJqb9o6uZEViFTtt0WT0tBx7HnUtv4Vb+wwdIJ
YreZ9mNBf8qPmKAcbrE0IUVlrrXN4BqvqZu6HnDTUVaoCx3Jabqeq0r3gMu2nZV5
8e43/52t0MyVqbYXXTLNdt+se1c1Z3REsF7E3hae/d24ymRRlknHaACZxP0dYwLY
kpCGMUNUBUWkqXw3y85wGBrISi9yJ89/dJBmcQ1yne4oUQUo20FOVYaupT26tnPp
XZJ1N6PjOpqzN7p3JNJbO8G3mFiPaNkRYL8PgAUvxTbJRldP5CsO6WbCcUkICYw6
XcftYi4Ykh1Hu6juQP4E9Ld1/1EuZ5qXwWdmh6v2h7DVq4m7Fw0oAWyYDm5xwcOj
A3b4I3pMpYmyJ3bdfzbIlBAOZDdzUzMIUNwgagXyuGs1Eo5Ubm+AYSD7bc+CtOtF
HJuN/q9WmqLv9rXmWAxCtOBSDTveOgYgaH0dTnJQ+21t9LTLwTiKp+RcmceHqIPu
2kKfoNEJRvsyiVSM/HJYGM9tBKk307C8/DwaSDxpB3O5ty7Tmh2iTuQuXdBBLNr6
tstXExR27RHgQRXnT0jab4leSS3/yFx8c0dfUe0cZgpDbFIn95IafW2IIIHj8Ffd
X3TdirRkF5Sf5FvN8dbKW1L7rRTvp/dzn2EDtya/WICUGa5xwMMbnrQ5azMq6hz3
pVAo5p67lQf6ls21CoAaWj9vRhFq0C+VjHsVVCjbcbTAcJGq77RYMrZeqyls8JXH
4pbQYAtFXn3f0kkp8gSMbmQSwdwoGAhv5uPAsqiRskmSMXJZMpmnN3YUbIJe27If
6nAldgiTHUVRqrW+XWdznIARVpe7eJD/Uu1tcI+GsuWy1hmJlpsP8U3FL7zuyVix
LPu8NzZC8fhLzjruIqUhQG2YAi2Xc8wxxmVcm9cv57HdSLc7LrMNlQiW1cyVg3cP
9t0V5aRmjgYUC9pmfKaycDRH6XrCfgRJAQuMxeTbEaflSBp+OMtwUXdG7cbHBpD5
8XuYsoGyZM82eyGn4kRAWm8LuBc7612ICGTpDg6FtSLZgugCWIvawfdlAxpRdiwm
+Xm9OinpdFBFo7t7NFxIVu4WuUYR+yuRvsGxCTqeJgFs+mX2B44beE7/gox4eBiv
KOF+eX2kd8SjeQ3c7iUDvKHe72Z7MFpgvHnbIezqY0EQ4CqEGuEdc7IJCooVQug3
v6m2E8YEshg3a5pTbYFQ1tEEHeD6q2Pw2/2qpPToydzVz0FuFii93IanRTKL3vbZ
2vh/DVsBa8aL3HMBYFEKCviEtpaa0q7/QhRkfvZqgERAWEBgV/YTtwUCztURn9yE
VVAjqWQ0CCRl8SV/qUEN5do3a2CrIUCdCHQYmClT/kLuwemj5Hk7nRNxhQ0pO+ql
VYGosaHJzpWDvi3vFzVxVZ1pV2wjSnDubw2ol87FgK7X/+j/A1SLNbEHQKtFeiS1
AzNVzS569s86xl+dAoyCwLBCEi+yiMUm8aRtCaMzaKxn7/KxaD6XywH230UoMGsL
17+o2Pi+rcKauJln1xA5y5GZSu2fkDhAElEo3IzdFePTWDrrkOvh5TJseLExuY9t
UJw275/BEdUgKPI5E9fUADrQb7DNmbYInUXTb+qmw0BgHKWAUnRIWcs75OTI3tX4
nxpxPVIrRU/y+GhPs3x5pqp/XkjWPVmj0ue7HzBourgTFGYCdY8OyuPvNSsf9rIx
nRI6mTcH7S4ys9HzGh/rBe6lLB2ZUNB/6fta4I4sVb1mXp0ZwDcQt8JoeAe2puQG
V5jK3k9dy/is/yf2xAKz4i/R+dsF8cYNDu08rkhyngOvc3AV3c1bHnOpbPk2KqDC
f8cQWXLLS0z2mZIu8gqTra2LBASkJcKEcyZvq5XOmp9GSk3HB3PAaVpI2GepHySD
4Ea1rDYeMzYvfXV5gQoGs90/iqA4RTpwEcEKzozFMTrpPAyL6q7uHkvGgyCrnq6I
c68exm/ySPBw83JJSDjGVoAYeIF/S7BLPvnP4/+fJXNiuRWInA4uKs5RyTTmeSQP
qQmZsmYusQkTWPpKS/w69ikunLliIjndUfkfodQvyNu0xX6a0Gnwl1OprzJTc222
xVp8w5Gweg8Ku/dKJmKJDhfm7Fl/WIc+2KjiCzvQMS/QQufwABS5LaPwCHMTyGmn
7bLYQQkgONiudNdfcbcD2GBAoiDBX5Tt97Aj8ZLvU6JZPauxlLoHXpLDcbrvvTnQ
jnVjCyedWkmhQOV/2yh2tCYKc3K5s/1374o+wkwKI+HrAGhyNy+5qCPrhxUj6FAO
Yib1I/FT+gGaPdisoo7BRrOIj5GoigWje0zubCyo91rhO4Ko3h9utrexOWgvbW68
LhVMW4G8/NlZMmwbVt3ERw14l/2bFeyHkeNSOwZqSFqHcjyoGcNsABsnRMkEFr08
EzyS7H47u28W5GGAs1qPyOoA96IEI2ZCrwytN83AZ/CHG9F2iWe1BRy+61xtqM+H
2dywR60plqhSrgJ1fFDhJybkbH+jg8KJaawdWjzV5PCnab0W+sk2uhKFi6ZMY3dB
Cl9qqhyr8tgW1KuEE1Gq/Dmy6IqCmc+5QdBJrDZHObuQNUKcXA3l/joweBUVAEsQ
W5bglG2DwvfuxxQSAn/aX35uv7gS+jXyEXO8HpSC9Rnb08MrU1HD1dZIuUL5Q/Ld
0XxeC8X6XY5QJkp+WgyN67rpUddrBizQRw+jNLClkGBAmvomAifck23eVEqbmnwW
3aE659fXkmMqCJzdxn4g5Y6LjqsSJeRPLJZq/D/cw2Fe4ue/QbDJNTPfJZxY5kdA
4slnWcJXloiFJK/rUnPKSIhY62fjgeRvcVjgDgEibMD3IiD6hi5U1a+9jADlYY7R
w1XKjGG81QaPtWLLVsTy1OUIO+inlvaPa6rWHwursBoecGLLr2G23QZZse8XyERX
F/TVGKM0nqMrsPdWJflqXeWIBCm/B+1IHuttrG7Q7MnBwPahrRL8uxX+yG50MsV9
kTYMDzAW3ZCUSiROhrSOOVOdTn4RDeONVLpOaCyrwkHDgHoEUgKsxsO4JPZBDAq6
iXhFj7COHNXCwU7Qh2dgytKYA9Aq4RWBvKrJ5mA/KlsY4xmIt8HovADRtRm4OhMJ
9XxUdeR+peOyx0CwiJobopT+Cc14qH9WyGAdnMW20TEJtQUPMVRsF8DYmw5IQn67
DFzp2/60MRH9/ysepJuC8NP3gmHBg4wf8JmRpECjb5ibdYOlvaI/inAI2Ryi1yoa
RSb9UiRrxJ/YjT99SMSI1TTPibh/uSmbqN85dOwgG+nlSA8kscmb7wZ5rFS8dDJt
xQdcsGPXpPpKVn8pd75ZLOLUUEUmmC++AO+OegvyPoPoCirh1CvTqThxT/K3gA4b
+wy2gKOEGJz4vYhFX9wDdQcZcxuJoeDUb8UKxJqOKDxpIB3GzmkMUmcJvHFTY27D
Ilj1Pm1T7fWHPr/ioU1s4rbSSydJTkoS4EptNN+6+DO1kdhRBOfZa5aZz+UyUikT
EgJ7xjp6J9KoEr0BncbOBpI1rZ0H7t+yk9ezVvSvi7m7CkgwL27qnhBMJHyNyhhf
Qccf6tsYey9Fjj7sdfyNQDKpWHpAOGV2HkxSiZ16ycfLzUiCFiBHiENWSwjS34r8
6/dsvjT9UeGvfHzQxiltIDAn1YcZ2VqkYsmHviZDb33t0mFXWchi91bTEfXtVHGo
f4BIVtGuFnc8XG5UM9AkhwohQVbK702PaTkrPpklsGg3SeIW4+Src0j2pnVkEp6Z
hnUK+BCnr3xpgAtBwHNCJO4DFlxSYZimNKgNJ5WCGvz+dkAX0tOQQR3y+umlSm8X
EHmJMC2uazjLIkd+py6ae0aglmRG90yYpZCRf8q7Ss8yHhWvUGBk2TbteEHjzlNO
AbxRM+hq7zOgs6KPR8CRhEy+imocCp4Zd80LA8FLOxmw1SDk1KDLK3Sz7T8rWaQv
RPyZdSOnisXGdS+fon4kyO7Qa38YF9HSOMkFONDiRP9HXPBvGVW1a7u65asLGB9H
4Nzt2TShlbFSuZbmil8fyiP4caeOIHo+l+rvPd03MC+X81lDn/7+5H18JkYfusj1
Xv465Gp7YcCo+jg3g892qnvlEQpG9imogQA9vuqC5C/Nlo6nz7rk7TNYHjeUI24n
X5+sRKx5P/v7fnWCQKtXRG8ZsXpMMyEaQvok1YB52/Dv2pUEzsm5qSLXjDBxdhhx
HN2E/Uz61fMojff6961ghgzyF93Yz/gbfi8R0DF0sWmK54PiHZcqL5RW3zJERkiV
C42hadhcvspJkDw72lzsL1560ArIONB/xaD8aPAxX9P59qSHBGK+O3NceOOQ+NxI
QwDGjfGSED7SLQRxznrKQUo2x53Cg6ejq9n5+sHVuTiDWAS+PtJi73BOWBVN/2Y/
EndPri2kMx60ZuMBBeV8dBzzO3B3Cxw8QyEALn2CfSm8iVvA8BZhImRbskJzR8fF
sFGM2jgdUnLIp+NdwUl08lNRBYmvAyuJGa5GjYNvVhY2Tj7pu+lMSn2rV1Nnf7jr
LL8tN4J59LgpPdXxZtzkhrKqSK+IO0Q1cmHsFT9mn8hSxumaiRYqD3WZI5R/CV6f
imlfo6PMeN8+zCQdIaHAgk9cnPivf9G8FRQ2jp0j/HxiA87vziQnaXGfrRY3MqV/
4Q67sdHEPjz3wTLVyshwE5EkY24e5EBqvnIUSBb2GyEuCrbKRBT0hbAqCfMGTpCy
KH3/igV3niDydGuShVSxJLh7hqlAV197WSjSdgOwqAROsnGAtEhNRuCCW4wq8Itc
l20Xk0XrEGu8bPs77Bp4Rl9KmtAOXnT3aL1UeWjaoVjDtF9qsu9lnwIazs7BUQuj
qSWEeqwFiRfjttKGNUbpMPAkHkkafZLwOEkeeCt/A/mCbrNn7Ng55XPDgcA/6fBu
OBPbSc8E4uCj3bZKENsn9K9NrZe9Lji1o4WTYz7uGGKlMsQHYCWbZ40SaEnPQ1OY
G16tJwz3ktAU46qI3VSvBNF3nDXx2Lgqdo7+6MxE/00v9WgcT+Fu+EOBhZoVPncy
TzNeFQ50o6VaIzwBDLWDXl0XNh7iVh9XaVuULrXFmUyghwl6OygcafHatKAKyse3
Tyyoo2e5BFGY+dBs0nt6edgvlg0j6b5jaWKsmZ9isAoQMgzqjAAYhC5ZspGtPm+7
M2RQj1Ay9SmjNOPGWR4eo6wKjoSWv73Myw5ci0tyUkQEsdwTVnUON9uF/E/ep8r4
iN2YRxNBajMC1rudHby+dWm0NoIOc9X4npeVJ8wVL/mOuQXwjfiOZdVAiY3U/B1S
/FouhMgbz9xjTWBB/zDDAU1Rk7Mkqm9lIHwGSjOzFid9JHCg9iQTYrzv6JDBEe+7
I3FNHAikuHrFwmmV+BhMOV59YNxcyzSchzTQ/M5umcvk/+FIltMN+zkFeJh7YgNc
GLjNSZ4DwowEMi6IuyZbC6um8BX5B8ygIyQh/vOh6tR7dwyJkoUhlgoM5AZWrnz3
G+fg7Zm+bvd1KiFusYkn8qaUJ+6eINDNfQjf/UsTqt63Y1bV/k87fbqKwIOCz7Aw
DWKz5zFCaaT3pLG58IfVNK9Wcq/7IGFyaqLaubm36LHIdzpbfXWP2UjqFVtNBHCa
KkUxLA6X5+/jr7bUp6SFH7y/13PNUKls9ZyZEn3foSX7/FS0Pv11GoJSozDIUXXc
jf2xdtjWS3hCa5dSdpHgkkXOjK1rY+xBXA3ttonpzYlrWTxyTvEn6r8uCd1AmFhq
9ZkABrsr68Wx2x7ltE85hJLIlzwr+Raj4JWzsruFtPttkVvKjg6zg5VYHcheWHZJ
X0PV+U5iUMnU4i0uuum+eDrV5Y0ZtrQwGjbkGESnXB3/4Hqhrs7P19Gdu15VIL59
OwjfEuf3WUfOcRg0sd+bAFNhsFjEeFPo1rykrpv49nZLOCKj5zkYrUA2SKheYLii
0Xm1Oh03Cy5mNYb3opqnTveP//W2bly7NJlHaOxdLhVOg7Y78rT+NlRR+kz3C+IH
ngW3T6K1SOY4RM9qHnA0TQIvUtGdvDrlqhu1+X4N8ecrgT9pQ9Bzifsc13615Thu
4ZwsTtdulSB7Rz20x4IspS6k8we4cjykY/9epua00Gk51C463n51HSLz+TSgMUJL
ir/iVDENqwBPm0aOKJSyMXdtQnNQLLSFzgSCly/whv+VYDd1PHGNcuwXnMRHMh/U
TmmYMkQjuhHeSpNEEgllRh3CTphYHaq+8KSjj364fA4Td4grdjH9XmLPYOYPP7ud
1vkle2lYVFyt7NqWmGJPISQ7mYjD4qA4OPOPcL/lGtvgbxN6EyFK5A4o2I1Wk6Fy
3AB08PUPuhzROsluI9CLSkUgJmBw+EFxEsvol22W9b/I5eEetJb6xTDwtKactudJ
PyO5U4TtAMH5ZWl8ahmHuz9jPfedfdNwGaOuvl+wmHWdCwKRelajjvwnKQ+2++Yf
TRBMDaB0RxZb+Diyyp6e8zUF8VtwyenZ59x0hVBLxYB+U9ZXxuDg1Au1HTB/kaKs
Sx9+T8UNtvEXvkxQ/ZwFTb3uZ+XQIUncK1tNLVBWu6ncNa0+M22/KTB5u03kgOOx
f6vYJlOKZWN9OHRQ7HW0Y1Q28bRGI9KhcWgEvHTOQZD21h4DbT8vOZ/Hm3kv9iod
hVEaTpVIx8WGCHrALLISBZ75gts+nwe4Hxg//zo6J3plg2TdBehHEyQIDsSy8O2P
7xidBjTTYZmr2qqHzSYeycXeGmGfKiVyeMu02/QFWzsDTDe0aV2AmIQrcoABDX9C
66uQyUPhbfB7KhsNxg1qSWIVTP2fWKxT3Q1xXcBTBAJl5RguxjYHPoMMCRXek3vq
z1U3mmJ/22AIZMvWQ/JI7YffePhP+Jb58cbvogrblKbNtZz4tM0HBqaQpdjP9bJx
l05WXMPywHQRtus98Mvi7h84l8Ze2w8JNUHjlNn1txzZPZPKHAMi4oIN/3I7jSyG
EqpslBYIbiLWSGUWHzLoy72+ZdUrf8lcqUa0QHVnQLzo5AseZJnouJhMje2Htx3q
qx+FvyAsc1LkcXNq9tirSAuzWX9IJd+Y6tjSzKRGC6EXdpBH2C+WFsHsSGTAJEEX
AvAwHNXM9qStVqy1U7yPnVmEJXYWyAIKhiE8F2TtO2C5JbsAj8VtEr2ERiKO9j/4
BymG4cStDwkklEqflOC4/9E9aFbysCVNhVdwjwBWaYOtzEvqbj9+iw8o11sIhMCj
CTEUJSmxWUG0kjIhLZXTYcjdttBk9FUHIRbKQjDPmrWGv0L2mTidzpkrcg6NpcXL
GxI9FhaK+aVRdBLkIFwouyEigiQnqdfD4zZrTpSlqDLXxcz6NC4EBPa3F7z6nYys
UPgntfbZj37SvxSnvTTQagH6A5H2uZ0LOb6fGUaVGlWYTXRNGRYEdctTNdHrxqB3
BHYFuPkkiIC1+HzFqocuuWqEBIko9kah+TB29ULCKqtofRqVjaP8pN3bfqdaqGby
Tgmd+YjqT1Q3XW67qE5V/6Pqk7i4PFAdZsZTu9tCmOxatGq6UgifdDUMx4GTh90t
ZXSy8K2qmYczRIc4Lz9MiFCI0/pmCfds2Y128nquGtgJ/fE8a4Ju2bLdgvzcbFz1
uaAl0N36TKcvqZ47yCm2Xw59egoGR6BfnuYpYebFXPCvo4+PnnnHeL0KfTYb2n88
RKFi01pOo/snX++13JV+zJDJunxpjtgl/vHa7+hTunfOpR4UgIniw6L0tzU1Qa46
/0in9nXtFC0rmUPbu6ehPpemAm4UG+x+QQ9s0cJqMPZ4KcokJc+AGQYiV8cteRp2
rHfqprukV9L0IBCRjw8wRhtTm5F1hP5uTt2I4uQYmZ/tIaJtsD2FHvtjSmYOA+Rl
jcyGOydzKx/PdZlM27zPhkXRSaqUrljM1ZMs2WqqEHk5tCaV2qQe3amqDun4PpHQ
IwWDhoGqAoqhAa8SUMlJ5nPSX0Yg0nRmr+P0jb/tOB6OTP3gM8l6bRq57gjC6+Ol
VaHqRn0xM8QSWnvYYv4//EtLq2AsWGwH+V+lp08LDu8Ga1/efQsg9LTWrlskZoBY
2oddx5GklaaCZsytm7VJLMq5TAlEXl2PAIPgSAkPyjlAZk9YYqEHwUNkZqnOycuA
pYuh5ls68yVmHhPXdqQKuJ9dkAzrpUIJMeChRg+yh06haPIqhaN4+fAuiV9sbWYS
Nynrr3zuKipmgEGX5bOVG/4aDFqnfcRaLG2MDyTPirsBG3kiLJGn3Epx3NEbtPaR
p6WdI/7KApSMBgA3Q2WwuFuNvPfFLEqivKHyjczppJERmspNaio/TwxuksmD+HmB
cejStx2bdr3TmpargdmB/T5sX36YTmq+9uvS8raLCiRTTKDXGSytJg09RN9mQhnf
xQdYKoogh7yVIDVEj1DBJA/9KdTGJI3wAT6xpOchF/YKrWh1dhHppNY+SCzSL5CB
Gm+L9QIdKyWESGG2IujgDZp+VmyNPrYgIJo97LBsFQT8L7XkUcWVNaix+8EI5u5y
WFSPMzC0SHl2K0k3Pidk/SVRezz/VGBZuvlQ2sj5ko373TIHNgtToKSpQNNHYwAM
/hzkzsRUuACFfyaQ2sSePqRvAL/UAbNlujeZ2V60jXnTeYJ8oGV6rjHTVYdKK5x+
euXAfYjSzaV8ChssoNnIwx2aFRY8ZtSJbcVCdXFF/PimQardcjbvm1JjI+BmOFbp
UjEMwL0UuoKVK54spJSbNII5RjTYLOMGvm0KuPIa39Jpg2qOLZ0X4RtchtuYrW4Y
95QyKpRu3i0XlgnnSDslCNzos/h/Vw22kDv3+YqBBU59n3urZ2YStyaKWM0Rf642
/JOTvgz9rGmCvKqjnFmQJt6MSTMohv1Ud9iLeVq+26Lbek1chH0jJrHEgEOaF6/K
el8TEh3hd0Gn+svpIxd5q/5ziabK+j8JYdamt9LrcNwhXov6YXUiMmaGXfQbwVMx
p4Y+me8P0gg2Q4fiDtdYXSwxSdiHR8YXM2MtiXOjSw1Waykjn4wOHNF2Mrmz1+gu
hwU9A86bdXRudV7P6SXV+HNd3zvN6oxU2kXnguQB6v0bFz4eESLKnC2dLf9HHKlZ
gtwfkXDninbgBtyzllZUvp6O0mN4NvHutPxYkll1W+rPWOrzGcbDysAJDmA332OP
FwNRzieDFVnTTGpDSd69Z/vpBYlPAMr1yIN42AcE/boZNPeHLasvw9b9T8fZtIpN
kzROEIBacBZwkOQ97b/qP/KNhuO29UV2piiYpeRCZE8xRJs5YJt837d4DpNjzPAt
/XzCWZxnoJ4Lwq8rslspaONXKFKUUuGUAKqiNDU2I/5KcWqStrVsOvy+0OesiYQ8
NlWTzU0HyTj/uW8bmqPIPtieOQ7uZxZthre/zQnsFZ+h7PcujCCW7y9mHcnxbbAh
zslFK5JHjKRHywWHG6T0VScHTMart4rHEtHLK2mNk9Km2qjDi38jOJL4rQwyDcJc
qi5Qx0D8EGcvzJw6pko671juIOOCWdDIKOpOVk1cLKOzva5AXiIy0FFeLRDXh7cX
w5S++zzP73i871kGc4dO1FqVkvuRkDVqY6VtZDubb5g1xQ4syrZcgPKzxCQwzVPh
Om14gcqn1VreFtT6eYsbOd1ppjqpuo64JIZKWhF2YaErkVqttqmG0loZM4+xlOdw
1fZW7PsjWJ0CpKRm2RXEtaYCuocO4kzW7hUMjsrIbExK8za7GfxfkvGSN3//XHdC
qL+FU2/3aQJ+iSf9B6CCxqnt4rjuUR8vM/Ez2DCRQa2YtV7CNn574mKH/8k9+vNT
uKnKZ0EW27ECxwybF3yS5Hh5pzb29pb63lWgaYoiP/5XOnOK6WlbOWi6NZfseZdK
kpwO1yhvov8Quap9fYs+ilt+iE6H2XwFcKLfP58gbWVcc2U+lWY4YSusmT5XY0Nw
4huj4Qh2DPCrwwz495tcvNo2qiAW3Dv6xKBnhsF5c3CXTF4KEDtzqgfarokTRoPQ
ajvR8sk6LShz28Rb+poGZ4ZuHvViAowFr4SiGQpRO4EaCRSe1v0vAgcanXnxcLJg
ndhm7l3o6C2nKQUFmxboYGw39/46Hjv1kcufX/hx/IysS5D+zn3P8fE4ky69zYOz
4XhYEyG70JI1eQqakWUZgVb9JLr+b5Lt3/wtGSv0VfB7JuEJOQZLQ0BiXwfKjuSI
N4xK6wyHPRU0F8E7b64FO+vQfT45Wi5R3a4DoZwKPJ1RzIqoCepttAYUJmQW2T2Z
Chb/WFMqqDC5s0tWnAnlg3AyRvwhnxZP98tiNIDYeOHSjjTCKSgroJ0EOmsTCJel
qJuIEAAk486np1dg3xIIqRSsv6+79V5OXyHjxX55xLs8SCui9XnPB8iUd9IGmhVi
Skkj08BqfT2bDKDCC2rPrFq/Ln469tAgk8QTycq3kIry13DguB3CGlt08SqIi+hb
t7byloYV4rRKWREEYOxD70JG7O1KlG26w9YRFt5klViXJ3zkW+bYlLSUml4qENe4
8/x6Omy73P1YSkUtplNFwgv+rGkCOP+7YlQmN1g96GkQGc3Jp+h7hzQgBKdWep7e
pHHHrNkchqFA6I9mcMDV+jLK9ph21IyvvVIIgzusNwbuBQjc8Yf7AA+Fnb4x8Dc2
48S6TTO8E8IPj0fnebi5+T9d+nwJQwJZ9WNiOA/x7vvSWHGKemqxKg1WpkTPIIuz
XdRRaEPiMR6wlM6Ad8XnIYGViRqyCM6BnopmVpArhsysLiF1tZh10Azis7sfeQGO
RNaTGp4wTT23wiDV0yGNSJVbep3KOhGmzeVUh5yyiClrtfqb6pN8ksa1WD4YWhRL
ScRgOfaoUYuhEP8i3IpZO9bP4V9tkXosAbxGgXLAld4AsBxa4wc91YNXJBQ5BbQA
Qd8uJns/G8GrMZzSYpmROJvGmTz1/XVVnOAXhk5JHqH1kpT5MRv64T/KM31EGJJW
eR1/BIU4PkWjMIXFa7Ta/2uXeiIU/YUKOpjgOj52mMTWJrbEYJe3AptlY/wNaC5E
7tRUBMFBjoWi58uCAAPSxx24DbeM92yAo4Ln2B6s/7RIXNc5ZncfBbDvGmOCTInP
KSYjYQR54WCqL301CCiAK8DfiTKC8WhOfu9vflwxWXY9qwXqp7wTfAJkDL+7vt1E
M4nvaUXl5WRsGUn3lwRNF7G0RgKok0gEfHZzlzggLG7F9KwFzlbanxAkApE2QZrC
EkymDcyRmhlKIx4b/m4r62chFe1SSPHbNZvKmhCObuNqUMBp0kZ0VHiCKesydIR7
nSamO0LddyyRXFoJgPC9W+nj4oqkN0QlVajBJMdPXgbQSkX71P3zTnOfSr5nCxa7
MaRcFC7fD8t2KpC2tidg+935hpQPjKpGJttdt4UEKEitCI07F/M2fAk/Dcx6+4+D
/X0yxJU41zIOlppm1xjxXwSUQ116/VhMzaUAZItgOVuhTWpuy6cIkbyEyNM03hE+
K6HqQOyokfWA6+u9Mit7sE0I1ckB5yeYuxn9GWFddZ1P5AYGFxQHaLkd9VqoCNNJ
2COe/oBICy9Fu89sbLAsiJ9v9ScD6kNhqOR3urszbYWCg1MVxZVRjS30DJNtdgDl
OhNzcvOIQDM2T/9uYHyh9S9Hifw315xJNWAWvHk576rTRWeLwdeqEckwDXMpadz9
i3yF0leCAEcV34U4m3VMzUxhlBjEr8UF80COL9SoLccSqfl4Ubshiw41K++zLfwK
MtfnN+YKZLEVOUrxbOX+KFvpJC9TaNcjcqQu9gyZfC6TcbbTHDZ4elUsIoUOfrkR
pq3KSON3NTnTUfVcqAN4n0EhalWhl18BnpDarEGG3/zTXc7+fsQu+GM3lpLZ1P3C
yfkPp4GuXYcWWusTbH7FzhDgr8/PD9vqBIdx6/ktWtwWyX250LQ8K5UhjhhsfCvW
8cHcvi+Ue9Fskv5GYHzjDaLv8rL/KR36/+iby8gnaLq7ZXbjXmEpV4pcFrggCzFa
zdq0BUDPWU2n/cjfE284c/RHdZs9mLGtVTTV0omx/XaUJ73XCD4x7SyPoTVFUWF0
P69rH1DAzI0DP8Rq1OK9RyeHEBwwVUO+YpE0T5TvtDY9v7vz1RxlnwO0eQSODbRe
XUDBhYRqiCCCyeWMuOmoadgFbiWGnCGZxTg6rgyWRqHfV0VBWFCxfb+ZKLVYHhp+
/UimT1Heemyf1t2OmVISKzAzJbLLd937AOMTuMuEvlcCxrdesIA37OaOq4hcVyxq
wLsxazFM97nPtRYGVPSwzjdKscvCqb4qW04RqJk6hVgwkg5NXrin+WjnV1Vu4R7D
nDoHY1p9U5b+8UoO2MjWn7S0r5DudgL5FVbShBX0VWeXjs+XNtWCy/oAu4SaWDsq
bOnMPNV+lCXSS1ZzK2KXYcz8VHTNlglVGmAUR3v2rOWLqAPoOZSbGTbR01WQtFbF
i+5WrSD7PTYm+0ZQg7vpHkqg1Il7HgXUqodZkF1NMA9L8TALS/uUvkMCzxOmzGix
ZEuggtgSxnRqplRWVhkao/CLHvh3jlloPQErm786NJPKE7IEtvDIxCBzP/WcJfyZ
SB27J6XcxgC5RZgb4PVjXZtxlr73aZvznuKji27ELpSXF++MRrYwT7LYO/bt5usc
9YEYH/Toyw1s9sbD4Ndd6XlXo3Vb7rjwoxlsglq+fhx6AEJlUqt1FT3RPuoJGMEx
R+IY/pGwtyQeXrT2u8B9T4KitDjyZFztiWrPYBZTUJvC8j2D1KcjVB2pcYiT2Qdo
8hJDgSD/ldwdwCo6K8SLTWfPA+Te08dlYk3FtDJfDoILOtMvC7jC4zUK080tkXCS
FWJky3h0tE/rlYMXeqZlLsnfyM12gW6R2wb+VDZTvGuFEBqXG8rFxrpkGWCwfMx8
5UH14wNexEKRTrv3pqMkkllDKW3c7Lz+yc4ooXsIqa/wrnbQIKSZftCyyV26dL9g
vxsbMeJ3pp2fNaF0KiigVPMC62+yt+IMlxhMephZZMbMdSXb9QXk2bmZPRj2v7yy
kuPMKAF2HIXidMqFe20VHYdHD5X5o6NKbphNfE9ZfukkVRFtVp9csyi1zGmVUL9u
D8hsTQQT+zIg/uCRlzQ+LgemlMk9X6j1Ts82SRWQBCKgV8/IBT5SpaC5p39m+qi6
KOwO1shyUQM9X/uNwk3X4qFXnMNjQrbPy2x+8qpN8CDRSMFRgiS4u74SzfV5MUpe
UWllmRlZBwc9tL7LwFd5Mm2w+ssFHETPWRV5Clt6bolQfZCLIPAEivy6i20aMcQ8
pnIkIdtieppWq0VW5zC+NZV7s9Al3REU6qtkWTktvLhgWeQb5EffKzC4nPpnJpdU
XPwSlWA+m2Hxu6JGNJu7/MPPdjheNjDHwDnGWIZyyS1lcVeUQdXaolLGPI9RHi3Y
eRWmuX5MpNFEtT8wgz2ljpAjy/Efn8DBFPNa289qgst5e/bfdKn7Qee4c8DoWbNK
tmmx61p8MLdpUDCwGQcr6y6oCWE4vf9D/YNIJ4aCg34TeccR/tXIZBkHxj66nGDx
I95laLsq328VCODRE+1cIh5WLvoEC0aow4nwzp7bZ/74WiqgyW2/w14fL4hY8DAS
kVBEnDZ63P2VYPDuHSnsSMmgYCpEZLjs2s9pQS5t4iZav6Clsqy8p7xKDTnkiKMi
nkRaGTN0Kl9+qSB4EfcznaIWbxLZAe0y9nMWwLDgWcln3/Ai4pOKw9fbjwFieLfy
TSzuo1GIqiGbSJOs/iu8jj6fTwVsC0YtAYGst0A4JCW7UnXg/U1bUbqBksXzqgxI
e6lTOm1TXHhvn1yOAPxJzZsjeOpDWtWZsOKNkVJyrWvGGcZspnloVK1SSQm+3jpx
x5ZaqqGuXHwpGPBIODbircxjxeHO6URkooyOwwc6H5MtE6crEXtIImyggRFhNg/y
3n+DP9V4SWWXuoYHAvd3eGO2GlLb2guqZhEoMACLVavlXBgVSrw4cGjHk+f0lWnc
9IdkhiQRZ+CRWM6OHW8pqKzTd5MLgXrBZyi980hnfdQN4TbmsALCecDMYX6TMN/d
1LPL0S0tRN6GRk5pnA11cMUIrucU7dFdO0IgSg5VrV7V1irUreCOqQQh8IQmUw5e
Qn93hFLHvdiFd/3jQ7zx/y7zDilfj0SWBWhvm7jn38fMSnuV3q5ROVNeqgXRYZfc
iM/4mzb7TJNUBfETxY0JZneEQfWNU/TQZ+WhGM9V0vtJXM3vahNQLyqFy+0sCRFf
Bc0433KtRujOAHdurZ2nJH7uqTy2HROkHZDvDqbElRZAT32pffhwV889Ju2pR8/i
hph7ZQFcdYVD8RtOkTRnh6GBZku8vPu0xTL5EFW0Kir/WrPaldXmNgl/LAkEIl+5
vj/cgEB1ZGWou+XhcrMG9fD+1vXdhfwIXDR6Qvgi7tD6UeNO4s6sfrwbtA4U4lvc
BgYf6laZ/PZoKi4t60F54FKtWLJbTH1cZfhVuWgvqv8DafmwF6k3ARoQVFOnS1wQ
5/2pXzvAj/DsaXgIBDCKpZXE6stK49RPAtVLrUZhA0RVlskPCVd1liAHVpM9aZ/z
wlCVdvv7w2ANp6GZ10/dzRKJ7vXjkKKHpLReRheY3tfyYTuPMzT78amzBMoOClDF
6rU2j9qcMDlaZugPun8sr6PiwPZSL4KdZ4nfDJgQRl9hMwpfaeU+jLyvRdWAKhaA
i1SezJ2XfU32CPPQKKhP9TY8KV5tToYlydKETt14tRlvIOQEEpY/4F6JrgV/DHsX
wlpPq8V/5fIp50ADbDKthx+xCbxjPjX0+1M/Vi3zcBYiUbRNayGYDgcjET3VDHNn
f+Oq/NFMr6TCmCVaDCzGsATAq4zwS9zxq7QmSykLWH3XQLclAwu2UGO7gRVVSzIU
rfL9tRrIOoOVtD0ygRbANBFLb+hdW1j+PzNMYk/jiDb+g4Un/QGmktY1ZLCJtOAC
4S8AwbXk2qf9T0C2O5gWsPmS/j6aOQYIHuVZ8qUJaeeUPPYjrgxwy83AxWhrC84B
xJBUaBxpjK/S1Zvy7ZwGe5nlR+6DrXSILBDuzLx+bLQ/sFE7nb5+uB+2R3mQuaWA
aea6xpAfce68meRue3JrZqmTvojIKdjPyq6ERUps+1NjbdHoEk2L1jgIlQvRcVk7
oHTokzkvhLa0CXDj0I+KZ9yevGJWBJG60wahG6YeNtPt1jNKhuQFlIpk63lAKMN1
3DWwWACB7Rv6mmEV7taJhKqk+SuAt/gSMM+BCEYXnDfMA88NwVMfgHDPOzG780b9
Whh/BrZ1AyFeG4JHb4lcPXdB1BttrBkTTZv8LCbf5hV7yJZuiac82eU4A2IOB3pY
THF1MV0/5GfM4gnbsJPKl2yZ/xQG1vltPctu1mBm4Yh+3krotEam+AwOpsds33RG
o8VgKiWuZLF29rqqqoZFid70O2hdmx36s6kIlyjI2t2rAMeDHe6pOVBrmIXZj4Rr
6MQM3SmQoRKYsMp0Phtx3l0dP3/rbt71AtFGAM4uTTX0tnD2XTxyugUgnwdfzOfL
fqKAClkxIgkDztf8msjx2l++799eymDO+Bca8VhcValCvIX/4avEP3UuRxoGsnk3
aYkvTM4h1dL5m5hUcU5icOU4rveEj+YqEbJyvvErcLNbv8SjFLZ6OyzQMiLKsFrS
gvAW8Mqb0EnQkacY0P1hlvqwh9WZ/BCAPc2Fm0hso/6hpCzUJRFhkl2rKtAI23jl
FeERG+p0VaJpTimhh521IYxSuwPrNoBh23pg1iZf4NUZuOLDdI9BqB8UaYoKSa59
LsS94tFS3YFZjuuJVtzidn7VnJ5OE3PQ6dQ/qRtg53lzNUoHATHUbzHJ0b5T6x4x
h4gPf0J+nAzBGICcZf7HPKBsoZz/RGtqSWKHG+tBOgMNJTAl3pvI6AK6pztgkmwk
LhNPfKQAs0BqmgKfd9qWrqkCpVDcqKKpIJE4ViidspwJ0w2bvSq4U+YWLN63kaSa
vJY2SZDuRJzitWYepDfydAjj14UBXFWdDfzukM2dxe+TpvChy8u0F85oIaeCJiXT
pqR8EFDfV9UYgix+IVLFJLsor3ULp4ku51axxi5/j4ffQjGduD3bMiGeOPoMMjD+
+YwQCTORooKdLfC1gZIo6YnIzdVSXSFtWwomLOKtQzuY3OCusopkMBJ9vca8yzyl
eoDV5HD99nusLa5XWkEcth4TzS2WjSzw9ptPUibXtW4Kv9QMv2EnqHMjL9dg+24X
E2ToaSO9DZh2ZJ7s1gBAcg/KWe236/X2av8XwwpZD6wTuaFdX0s8fDj4ZEZMoZh0
Bz/wj/MSlRv2ZDQi9Dey3AwBJYXz05ovResUX2uhdIbwmfKrM8zXKAR88Jk6y4I9
zswJn8czpJQIuBV8D9GgLBxH2Li7x9Qq2936d7dSxVAqRTfQGuCjYX69WjUQF9tC
1qpKa+MVu7W2iFiQCKmEnRltRpoDxjVLQr/MptDllq0vaqz2oczvBaMaCx6I41Za
MvWbXmCC6Kg0zDrBrXeH6EFzF8BMn7i5+I6mkjiAbwX/PWehU4bTRMkRh+bzkH2o
+BWkkYnJu4+6KEv5CYNL050o1Zr1bdEOg6qPz5F6FNtQaFazSfMbVHwUYo6UNsy0
64EcXd/WU9BZXA9rzB97KZ+6YRjVg2fI+F+YiuZjEDFKaH1kZRgzfRSpl0tEm5lI
yEybohLzTQlfxDYg+oH9sXoBa6rauqtWR2pqMVvy0WiVNheeMB0nMgd1KpJc8i1+
++koBj+cdudbQhhgxxsoHhK2Fa2qFIqVQjAlVP3NYfftOXvv+QtLo2HP2OYUYQ4Y
e38ufaX2eO+9dkkXg/GjS6LC6Ihvfddpf60ku9s8uwXNDCu9hiFLcyIdtZevs+Bo
y9kRidWdBZAA3bRm63azS5+xSzn4UdS+nndYtPJ4xaq+LY5YjUpIDfCabDYgs4m7
CW3mJ7KOncUWO0wKSeP0Oah/tQVdLq6Yo601s18Q+1btCASHCbDAF5vXrRwy7HvN
LgS1FpMABDN+qcKtxSAJspDvH3q+0F+DlK8Oeh7gFYhABTdhf1+3787PjvLbIJex
aKTNfuEqWKV2zlnEsVSafef9oroaQisV8fjLPrT9AeUS7/sOq0O4L6s0htIw9nt8
cA7HOHNhXu2bqH6ldzHfqRPbXCuK43vYIA23FoWoDta5mns0Gii+mnkuiUlJG5/Z
Tn5S5+3CXCAf/8TAYDrrpcYwPs0P1AFMxfwj4x3Uz+CV3hNVOo3T+afg44j8Tn4j
lJIWuz6E2/z9JNqO2z2IJmNjNOpfSmmtnYdFQvtGEI/TCHBcM7epFbcO7yX9xBQ2
mIWQWdR+K+yepfhSWaLd81OnzpkH/rSc1T0SYFxuBSK1xpEhhmMsF9VPhDyWFQzW
a6A0coDzgPp9GdQXOXxZ9z4IBRJ+9EDqCXEQ1NnLLh/u7NP6LvW3wIfkFhxFGLH/
//mU6OFwjv0jqZl8F1ejXYx4WA8pwMLyZTrNDf8HzOCB11bGn/4Aj7Rk4+IgpZA0
LZb6JVoHdgbM88qoaK00qK3Oy2+z43hCk8PlNlvbfMpyeyTspbBCdvNPeKeNuYJb
qsoq6a9IHdlCEWDUPQv8hocrNXz1XpBRAnO8UrN3a97QzXhm3ohUH+TTWXpBF7q2
YQ8KnfbP2QEQaKlW7R3kJyg94bBcXlzXeWkRmynw3ftGHwauniGptXJdei2TRhQb
NgLxoJmSRFohYgp4DHnorbxR80giD3+TC/RASeAUc8SGSFCze2jDbHxNiRVa8VrW
6VwkZQ2hloFxn1YoXRvRcrfd5s5GunSQj+HayszYH2P7bT6gPXYjdZHDnZ1GseuW
sOXZZ16iVEOlxQC5LE9mw1LgHwmxPp0Sm+uqlTGG1d0UKPQd4TEkEMIzGWP/dRIR
rmeZb10LIqpcwmmEDG2AAJUMrkjWuHf65xndgjKshIm9AL79KV836TZYPQhugjiK
XBugi4GJIAxR+0udbPA6DLaX/Ue0QJbCkCLJrmcnH0Se3vJhXD2fcfFjAMNp/fOq
l+i0P9XTpPeBvb//j1jzOlcXqMHB4lE8yYPXRZipjNyG+VJaLgrWT3VJsp5nJIDh
SZHdGtV6SfJ2oe5Y3vDEfYkgruypUg9TmLu2gTzNQTyfJT1M2QW1S40TvwQcb9da
DNV4E1HqVgPqXIKC1zNJaUjLU1EbyACJWhPyMyQDwLwjo8F04Rly9jM52YH12tbE
gnbqi2nlhdIhaMpk/AuO98ieLvOyQJFzSar4IUVLTyOcF+KJxB+eKx5IqrISX/Oe
qzC/DZwKj5UxeHo35AuaU+JozMzJeXGrMFCRttvvmc9hfrWJKECHJ2JRkw4ZDf18
XgWntGYPuZ8LoiXlENx1HKXHX/qVAH9NbX7OF5xfF/sK2mygi0WMcqzAOwaYlfrn
kK0cPOJK1X2TpupS7fK6hk1KrfrMgtDPtx3n1rEJ+DV7tyYv8T5BRL59YvKH8rlI
LrRidp/+akf2/T1EGp7FCRdGd0lzoUh3S7p0rv4vmaxGrf1x9qi+q9oaAu/YlBqS
veHi9PG+uVv6IDG3RGRCtc65SkyD8YvntiXk9yxFPQXHe0SD/ut8zvB5VTwwvF/A
II4RJIiOxR29DrniSC0vHnS5UrUp/P+l6xXqQijtxmfR6rpMYRkHIcpKLpwNfzXg
nh0cmxGeXkeTayEEXD1LYpqBiX0HYRy8ZguCEapHQkpJ66jMznb81xuMNxytGQOO
VN/1p0ZKW9vyWEds9quB1FRocP1Cysz/BEmQp5Nfr1imNGnVGJINJEglyqx1LpB8
s7hhL5/+tASy/1C6s2OFWHDnMyOehwh25KLsRVPbBr1TCUQjpV9dS5Mm9s2w7lqs
oD+12X/ShynIQzhs7pScC5mZ1RSKk+k+0YsTM0yi3Mj4CAk59XxBf5uaxNwNAdrD
iqbK7DCjorOhtRiDA1xVYTXzH+nt7n7aBaGBqLw05fuxF3Zq7JtICNWJwb2+dlSL
jnFg6++B91EyTGe17SNGxYBCcPLf2xQAw7ARXfbmfWc0Kdbk/dKSr6uQRu065htH
`pragma protect end_protected
