// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QTaG/TGFFVZO9mwQc8GtnP0dlK0yBGpKZyDoHHnpp0fFy4aPYy6IClde8V40bIoH
v3XdOxPqxeotmAz9CoERRlDTOuUfLEUW/FibfMlwUyh6/d6pAnbxgOvYYQTET2mp
11ajIU1sSW5n44d91ZCDX4h7RZ+GzCnE7Yq8gpuaNKg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6208)
RAjTRdNj1tJoib/4MIG5VSmyqLCSS0UxePZd50jcotPPGN/ctEA8lyv5PB4vjXjt
xmlkVKOH+3UOi+Kl9uYghQ3N5VG/C+J47yWneXK4LylyOr2gOhsoDl4gBl0EL+6d
uWdsY6KtpnDiwKdc1jKVzrkhZMapKr1yhxJkfwYyAZt/ghh10RIqvJSnWnL80BQw
Gtjgq5G6gZkpNoy8NPszna0hVpDeXSFvqnE19ZK3mhUTWoxo1lT3K2CmkPz3/JoZ
KBdvqw7SaLy8xYepWYasJy0vc81vKlKoh2g78HfDXIHqW9mV3I/znNejIKm0O32T
a/6KeEtE52w/O1jYqY06cUBDQ1zELFZTclLm+W5uZobBIkU8l+Vv8asewkjqMESk
DqyuJ5XpWvlTnns5fT3mZySYroN4Qn5lt9UxQTnH4vhEHwxp6gVTnyFOJifB5XyW
MjIscY1rbu+NKnP7pNZ2qGUQ9lzCzko1CSk+KT6I+hjlu3s27pWLmWfBgT/8DSrL
mUnbsELhA07fDLzR3jKRtAD6O1DDDyZDdmpR8g4pG3iGV6pLrmAXFaayXMLImeAe
wvIH011lF7mTfZ7n00t5paWYyzdrBBb1HglX77ORw88NVvXyOqaeDJj6UmHsaqXb
AcZUgadJUkFX0NcMwi3DT13xz1fdykQMnvF/GjQy/AOnGr6KwKy9w/uDAuvvYshi
ZYC6m9SGYoOp/9iYFCjZu0r5Cksc62gT/bkvHxFSbJcme/2+uDYIKRl6dTkqy5IC
3FYNZgC33VqiUnDK++oA+Pkgu6QEaszhFsrlu8QJL2jFZh96n2o0mKKZduXQKo7H
YJJv98zwUmMGgAWrifM4X9GCw1YsYZIj5lAyZnNLJ1+b8EH0Vl6154O739BQ+iJ/
lpDSuhP9WaQOB2c6ZBYnYy2GnFezf9/RlV5VneLl0A73SUPWMTkcqwOETmrIiiLS
fYYiqswx818evB8gN+v6hzfLGGkSVQh59o3JJ3FPHqIxt293nq1oa7w8+iu91Wrl
A2SiRl47uR0K6Fz8VjXm/4TmGEJj3gBFVVJR8m3hVifuSXZdQWtA+5CZcp+BV5PP
MpNTEQgJJjFvrkXh5GS/X5XR846vM3a9fhP4wAAuXVo+zY4wZjfuT/AOupSOXA1Z
7FyQlsx+ZVgw3GUkuyWAImMDzPqLPFhc+dJ7S4EgBvb4Mm/jh7rxXRAn7meMPpcj
+7HmmQ8/SHSvlfv9Ql9UC6imv3BWWl3Qti2+FJ5BLpOb6GHDgsRaxuFalUJrvBe1
o37RonOjNSgLhMiR/Vox0tFr48c2k3P4fu3N7QdhuYg+9djWzqj8eQbF7TouyNLj
WlG7XsPfffG1xvITHfKXEtGflXp9CPhaCLOUeKXxs7NM2PjAGR3HziHs5GahbZPy
wosiG8dCtYn1AUii1lsLl5JulwR4TsHcypd2KAaMtrfksQnmGsx1XSnr+6M/fs9S
1ykkKT4ZaWnj/NO1Kzz3nbT8wwH/klNDX6hbZ01BwgkpRrfBTpf9XUU/mV5U8rYq
+Yu3jnclU0VdK/oczy6+Kc6kKZMpc8GLPuCxNMJEEp63WTsugf5ncUJvly5E+JOv
Rt+mMNMC5bMpxDGenz2h6u+ZSnXWOtgAk9pnAgQZv80vSRYRjvuslgJN0ogHAPRc
JSFaBz99JpOR6YCl9Eb1R5jQHQFv5YElaBuw+iwhR+knzUyxkGrhTdMLI97PqGsx
fLIha61s878g6J76KH2IuoZQfrGZSKx1N1doxX+TpLflW6ias1b1dOHvx6Pq6yY5
7pHerDIIcnRx+cyT7jpufzIA/gBOVG0SlcHO+8z/b1WnbjkOGmiPyBhFfG6Rs0EY
0B23rOd8yzcPQ8Fe/v8BSXFkaWSelgr65QXGct+t6XgPI+cOFyGzXiLMFm5W0PZC
HfbDcH7z9wSoBADfRSltU4etmyumCqIvG49tvzSFNjEDFRibofVE/6kxm/bYZXbn
h9RNJDg4tYy7EmKE0Gr7Pk+bXCWtu+YT6NMM5hErd87jEXNmK/eeI6x3d84GLjwO
QDWh747+jC5INf0xgHSA7OzlmEEA40alT37pnGcxdVeCf9UAoTB7txXkHGLlJpNF
c46MPoaBgj3V2eInid8fQjApMBHHLctEQ3s1AeuLGY5eZr7dUiKubhvY/uYXvyQs
eF5yTF+6yu0qF6i7lPvIU35w5og7VNSMCJDc/YGRQjF3yF/kJTew/jM2cBwpkyoN
y8gJDBcQStkdePBh9EqEYGl6B9X/J2pyY2F3uJe3EFCpRQwY3c1TfrgSByaDZhzK
D3JGoaTrH1esgK+tpVDRnmxJNt0Eky/CSCGy7iLkvLz48NAbTg77OorQj0Qx+Ttw
pL0BcZ+EhY/vnAY6g3FmXrI6sN2+CmORwTEmolSlxFCJDiJyLNhyuWcACRzOZxKi
nqxgET1vYsgQyxAoBAcyKhjvWDDBD05PTcovZajYcxXUpz9NTIldNVHWoDcgeb2P
qHoAQV72IicqRt5rGWy8ZMv5UcmM6ey4IQnGC/8pZ+VFYITyBaGaZFYzxKBXdWkb
e+rPDVmDWhTTDweDPnrcVNlHBxSa4fGI+8l0XKMt5RCx9VCISTKcNfzUqOdKZv62
j7sK4VyMOMLqZqSVnpVYHNvrhFUC9TxVcS1qEOgDADZ+FWzD9ZIu6dE96VXNtxRp
R77BRTxRHMYGcupG/hbMGIET7Rs8QtA+YiUNzu88hucYwRX9aoLchGZ0pO/EFZ76
I119aqFE+VgC49mDFlYn9m/I8yZacX6d2cwOxlIZV372uQrRGHxaYuP5aOo/db+M
+ocwdmFv3DZm9Li9Xgib8OENY1VTBJlGZbh6Rw3bh2SwBbZIhWamlJz6QoKbnl+6
pVCFaQIl6i8pclX5zGoKX/oE4+9SjYZZe3pofM1zeTOz2ZKYgki4atN3KJxB4gr2
HQTsPXyBMiarg5n5uVCtoh5HqC/kBgNs+sJ56kaUc7ihTsAjBES2FsWPfpXgr5ce
gp+UoNrlkeOPLG8xX4sCOK5yy6YjInECa7ZcnmEDWfwuWZYrfMF/PPvjij2xEpHK
e3ZjluceLIWsnowoHveoYsPbusoqk+5Q+gkplIrMe/znek9hm+Ukrt8tumYDU810
CSjU9j/CrcHKiByZbVwK5P+3WXEBq8jd2rjXMF1wlSdzX6N3HgopsvgT/gOci5N8
55NXd8i2JvnRgzg9ChrrgL1zx+nFvxgGgg+ikl+WLkKM6e72hNsMhqGWSx4x2wjt
3xrvph0Ctd68eBG9jjOXC/boifomJyjx/ircHuibvfENTFLP2lev3ICKOejDReDC
IvyaEbj+emHwtraRwNS4eS8zUZZAWf74VKKI1UzbVceNf4N2dGVf5G6LXybm4yLr
xcpsOTfeXbZGH6J2nrJaW06bnWXfIm1SP9kYClK/KXnRy5uRAh6+9hq1WQZ9KDMK
Q5c4qRE/t8i7MDBjV0FzfPfVg8/eWyyf77zGl/Z679fadbMkA0gmA3PenxU5NlDn
dbZoogSZUSw55IcY9lAKAQCA7Ks/PdEr9cVTZQMo8ayP1rEIHcrBqskWiqRkKKLp
Oswxuq/X4N2ypuOyuF1F9dpOBFeJ95iZ7OQK9AJcfbNj60iYu4aa94pzk736DQ8c
4ru77waKhMlgoMKXnoY5QxHTrDhX5GiqrllYudkcBKVHjccmi7tSri71NkWDEnT9
pFFHELQMNYc0bReCFCFoMtKk78cEnM5CyKquU+++8uOsGKDyORxKp1CA18mKKErw
ro5A/qHhVUckjYAjXSoUTuxsGFgeFHRgVYBTskBsdqVtQMOq61lBoblysI07oZix
1gekpTsplQpzEQdPSOyFigs8XfykMhFfa/fXyCI7P02a5GT6WSkK/YfPBbBhLZBx
0BOw4Ta2tfo7SV0A0+lF6cjkp6vFJ0lpOrjf39DjnjLGLYzDzDPEU/k7us86OUvw
RoXS+7bip7k/y0cG3ppy08OMDor/JGdN5L+WMPZhh2RuPOasBTPqyhWmG2V9M+Uw
3cQ3QV+yCSaAE078ItxtIC71FjFmwxs2HDt/6eWq9kgtW9ui7/E6q6MxQ/2Fmmcv
oj/M4RUzGM03xrWESsLkoVAzoNvBOIdhLpEFb6CcQ9ua68Te1uVLrMDfg/KFzTiy
dPyI6rNA5wNG8KUJUeG/21kNuGYOFTbjbq+/oahY15RULM931575HsPhvuk6/THu
IscdaGyGS+2AUC88S4j5jfOqCY2+MYOJx3ObeZMcv3XCs40+k2illRgzud4pSg3t
xn9K6yBauUxquFRd6/idKGeFQMBM3OTo3C+xKh/+9H8LluKtFa5M82H9ZjxULJ4S
/5PZUZoO0W5uaTYOg5wq1PxFi2z77pR2puimjl/1njwLYiwo2V+NAVf7Rr7PO/va
ro3AnGWbTkHgc6BwbHpm0q9HuMeEPnaYo97lzZ9hl5S5QW8aKJ4Uf0rsrg7pLqzn
tPD2LrNqhCoaB8TnKgrp3HA6t7eYcrADwmExd1/HnIqD1wKZe1SkhOa4SIqw44HN
8fviXdtccrZ14yH1A3G9N6NsUgeiLKsvSpDod5UgOTly+Dpu2VQy84WresRSDXze
e/sr5t7iSALf6C75sZS7QoABwjU4Y/pLEU462C6uKQL66kLiAGspDcJ9FE1sLNcn
iqBiqfpkZjXM0i/gtIA+p3QaBAJmr1kD6fmG7W0+wthkeVHfQAguQx433ggJMJ+7
VLy0LN/yXdVYvVJmABi3ywXysSazfTYla+wATwZLvSllJ++kT23kDdW3fcKdPLHx
jlKLdFHaIpny4vK/hW31KWBMyXWnLHptkk5wfxQ2LDubXu1hO2s+AYuyESX0l9hu
GHtNHF0opWj7pid2YgXHCkQdj4pbJb24wK9F8ZS7PIOWsY7JFrQMjQDsE99WkHGH
N/DpeeaNFPhAnmlq0mdt0hGp+7xbwmvEAh6GVDhzNIF2T7y4NZHLNdo4X8dHfRLZ
WEI1RRZI1WShLujxxOtZg+4y5L+z0YMJxd4udQHEkHilO/+4hA/7w0+nym6Mt0oI
gzEWIBadUWX+nyHstQADa8dpXoS9lxKD0zxegsgmx0O+tV1qGCgYibeW4JAWk2HV
3U0bPNlpJGrSqjFDCDzU1QMdBHpRUHT6rW6b/+gh24BNiM+4y3i0kClrUaeV9U53
yEpoeZu9Ktzy11jkbCs4aQ7ND9i3gLHUJRjehwKP/bGTDvczlmtwzWgufq8n62rW
VrputAQA59BPATaZJOQW5Wsh7/LBKtY6YpSsXEqpyBujUFTy2FcSOvXG6PqdDH8P
7h5s46y0oZin4/n8rkeVhZdFg/gluCLaoAiz6M2DGJep+SGnFkQv8kRLCFQzbddF
Yzz2UwOnleHoThbB0I17axnURNwBW8d1o1MzU8jhPBeZ94beTB+kPrWcedPOXWyd
wd8JIXEg3/c6bard/8nsvU5F6w8Lpt5fPnzyykPijCTrC6b/LxmMBq5A3G8RX9Dm
uHWAoDsE4hUsoAEXjxNKarJUqnRjDKSd1o1t7i2kwK3jnhe7ffodcCP/rOMB8ASe
GqY3DKcSX2KVLRGONDeuepQg8NgmJHsKeYKqiQyfH9R6I5POkABTCHwBBZ4CDTE7
BWwW7y0i+j+HcPyGj1lIitXCYuCXnO4BW+Pq/tMOi3xoC8W4aO9Q9G29sch/X5+q
XJI60fX5aA7pMuHgcrnzgsYHeF3YVOgOGn+Jrd+ytzma/buRveWaslNLakM864zU
UG85E6NT9bVg9DxjcFV9zYzeOhk7BE8ZOPFPKgKWhUvPLfN8iWtg7IrKHpg3keZL
fH9AZlOTEbXEi15MJ6+k7lvjSqm0gpCkPxno4bQ+SeIWTfCOJQlVI5G1MH8OaXbm
G5/LwYS+fHQBh150JpktfDJbqhS25oHhe7GrO7byFFU4biU0UUVCZlCgHwZ94YhK
4q/ItPEQSQOsBBOJbNZ42Gp6f1We1nYChdBODrPJR7j9YpW84RMZpZSPmNy+sSyP
OoAWJaQLQkZ51lGcyoEFaxsb2aUJiC9V2R6BIPLX4kdzHznxUO21CfqILBpTwRsr
QKJlgsjUXyM3tMphji9k3KNrQZawgShzKv20Wg7kw4ytqyh2MgeCH0UGB+AGu+WJ
qiDX4QM7jMS765/98PzmpOpWdEj5lwJBeekRs3arVCdvA8u+/CBbzK8OZSC4MFvs
lXb/rt5i+QAW6mFRMnsHWtZWUJ1oJL3RJbVQkxOLaznTRR3tvOLYfUQ6c8xpvK9a
OJu6S9QN2DCca0KfSldluBBo7tsP5pSb3nREq4YznoXoeZc8qeMNUPe/I4oLn+0Q
SZRkV8JPX+wN4d8rgHcU3WUOq13Hp8tpnRz/Q3PklMvwe1suamyEiOGFJ2hsAH7g
th03bKov2fUHet1Lld/8yMvYLY3RJSiDQMmYKfLDBpis9of674lTpHzUQq/yJMS3
L7yEWVRW55H5icnCwEpcOd6McEGttnMw1SpsN9pAbSr2CcUvuAjJ3yNF8ARpT+QY
P3dzZ5q6KxtNKNLYdCpV2rxiIItHtyqQC+Z2H3yd4pfbCV5R+4pLM1i8WaUCsTzV
xjNteKaH96ckHfwBlqAhJYbt6INCZiua3aFtsmVz5mb+yPXcmr97i0Hsgf5JdesN
3w23zqHHDLQlhKBiFU9G2Is+joFlkg2qE/bXUpg0TuEzmWt5hJ/AkFlFO49hnzLT
DcWThd8HKFfzj1fUWpbuBAhGFba1Ar0eR5gmyS3IqfDpy0V+8jWghXyCl+fmfGx6
rabywO5D1Nsr/mWrD4O+P25BupjAQGzmLoggQzQMqGH61GZqLPS6rk4e4bkZH/MW
pI6wm/3q8RlNIRvbj9bxNEv/XTPnkcSREFGYRz0dgvYbotgBInd51GufesTw9Do+
nWmCX3VmP7g+SEp0NB0BioMSypd9k2BefDZAp0A5nC9j0t/x5chQFqktgqWnGQTw
dxoYBULQr0QEq3VJkdklIfsxS2oHIo8hKNfSSNqjSEwPeg8cFKReC4W8LBOFEqZh
KjJclNA0CC6kMg323eUl210Ohy1z0xCQgJ91trMM2irznWBmuBMzvAx1ej2b0bbd
SAUTumo6K9a+8/L/1JPEAo61Q5GERbAFmjIGwi7ijSKmOLu53g3MLKiJ189LrulP
cz9Tuw5mEA2loVrSyI+XT1hsZ/NancCWXDHOqCkV7B6Z3Ei/OsgKIAweisTlPfPy
FsqoBKfQsV/KItDR/NInJxVT/zAPBniij1fEcx0l71LXnsJiFpHyjW/dIyHRCocA
8TP0MnwEdRhZfqB7SYQgs9r1Xj8nDPwoq8wa6ysRYUO2fc2K5GWzK1h6i848zKus
X0bxQFWP5pxRVrIHj/QjJwu5Mn7k5jjmWnwb3ng0G09sQYkm3+63g9wUhGKbImWx
ojPajbJKB/BA0d5Pp7KG5RjS6WVuYauOEEJkWAqsfY6m/hYfBryB1hODhwe4seoD
6Owi7/Q35Kg8GRjYPQm6uay3BAJjE3cQEjBlUzB1NNGT36xChdsWCTOb6GonNePe
xV5hfKQ3JO6bGau9EjDGYnGh/I2Y0Oj4EZLLeaYztFMfnPo7ho9Yc8hFeXymR8mv
F5OGQnB26BW772vjDn/5flC66mVUwkD+HZ+Ebtj9Mm59Ev2EFOIKIBCcNw0MjIMM
R7QzTXPwG4/ncMaVC207UOPigtyx7yIvdX/SQyYWcLCTYziOp/uAwcmgup6AGzC1
QNo1zfZMJj16kabb/bqMLQXLGr7XAI2elfvAVauyOOdbaHBqA0dVRDAWNwYS7Co8
OnEHbBHYhI/tTvbuDnHO0E+mmdVM/6d/TbVGrt7BybqdxHZmccwfIgo9boJnyICg
k6qVa7RUx0lS/EOkONlC9TWExUEYx+mF2HTzeIuUosaN3yKawMyzeOmlv5210SZT
WhVOYQfeRZhtA1Y1e/e+LEZgD5hDemT9aVxcZuTknA4NYjilmarSu2/lbh/bXUJE
koT1tuBbENkl4q30YDeWKDUew+GOXMYu8lCRYUm1tL2ILK3x0Y96acT1Ifufxi7/
26JuOaou1zchoc0UOgVeNz0/el1oGiWPvPhBLYDda/uV28uiw4RNoon4jipWa+0q
P5qfmvXm24SFF2qgKf7xvt+zx3uiox2ocKbtWCJwD44CBYhGyIJRPLLe/Uvx/w2O
e/Kf2pGsJQRYetZYGwgjAIoBl1uWqtn8rgK5gVvRY0C13ZePT+453bLgd/TEjuqp
qt1pZ9h3dDzExgCNzCyQZg==
`pragma protect end_protected
