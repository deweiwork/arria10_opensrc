// Copyright (C) 2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std
// ALTERA_TIMESTAMP:Thu Sep 13 01:35:02 PDT 2018
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ncSiYm6T7QbPE8NmaklT013m2sUzDLkLC88pfvlV6In9sjCrJRGTnyVikDEB5zc6
1XSAwHxpzer0wfLa+8heU4LbXG1Jnna+IlQ+AphuT+dijN4/DcA4rbO3PNgC9C0M
Huy3ocNdbzPfTyXzaoYFC+HlP555La2mBlbfIqLRxHg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36304)
PCJFN2X2RzV19rTV1rwT8NEkQ3FQu+J59uJpkN8H2kyqztqYAzII57kPrDNFVnGd
JJvO0aK5bGW6G55iso9/g0vHhb64U6FTPeg7y46F6M0EZwPV/sL3YYSWYPGQrcoM
3lVgvN5Kuu896Hc9ZK7ZfjmOZcMfRuzVMEHTwD0s1qeKwmQ6f5xCu2RTHNveLbX/
QaIoCBTzB792WDlKvjALctqbIqqyQgR18Fkyk6aTUtE+JV2HWZSlxLfIlRhv7NXm
H9djO2E1vw/4R2T7rEP4f8GVaO7nl7qWMoisCMklHWHqbDKAOLi+tH5+1w8UIEkf
yM5W7P7YvxsYN/nTYTLS22m26+vSTbv5TvZ465wp8mW/mB/GAxRIH70iyQAKxToq
WlUc0breJe+msOcp1r8jWy5Ptbl7RlgNa5oi8fvEBsYnIOAzh/fKWWgGZyTMZ5nt
5XSxoYmINWkgrsnuu7xG8+2WdSLDGRSjBuoMautR1eTb4+wLiN1yTQOw8shkmxJH
WXQW6Z0rLXFrLboKQdVXVZiXzTNj2aFg3sYPjsFz2uKhuILbdfp/L0ED+XCG1Y7S
u2ijBsGTGLbt5saMkCVrVybC2lp2SFRMVW5F+9d++GdJ8MviEiRtob0tWhd/ZBcb
5sQnB+Ehajte+Si7Gd2PO1yDNWrmvGVumJq2Olbs+p+oXS1Vhy6uBi293XxiTb/q
bE+CPnuogOmiu0Wq0Rwsgrl4vv4LiFoZ7iM9Z2b1LGs/FMth02dZVX+iULPDTS84
l8CYmW/EyGEGOtTw/NhxPQZ6fXtiGCIo/mx8t6FcRA3FHT9DwLY2hfM3ifJa+qgn
EEqpPOUcfTweeQvQkFjkrgwFL0Vscv1Otb5f+bUHitlgBx2+k5wngwJ8YV9ozv5z
LsIEjwxckUYDB1wuka4+pUeX6EE0O7Zt/vjeOkgZnyeztDSDFQdxZ4wud+bBksrL
HmBXMpvBk3TYw2nvAnbEU1kpOHO4cgeS3FaB7b8vi8/0dGUQlFUu8BMEwf+T6O6v
TlkpawLfyIC2Pz65yTUBlqRD8/6wbbEVwPCQEGAH8uYEwv5eJbTxFPuZ12OUQA5l
rD7y37i4MvjCiOfmPJCUZByp6W4TOBH+jmRtBL19AEmP4f4H+7iK/pnMDiAsgJls
0KoU71sFbsNOL7E1cIXRzQKOuKvlPmSUhgyOTIg6bqkPN7f4D1zZctr6ReX0+s2k
gJHHMT+NgML6RTU1SR5uuYppsiIYbgnmhaqgHQKkJnKBwrND7dGuixIgolpbzpiQ
Hsizx2jOkjqEVSweIF9pzfVqVsoNGASLlW/JYz26dk+Jwlh7SPs6twaUcUzsFNt8
gcwtraF1L2vciDh7m0Gr3Z8AoYDIKCnyxldkmry65Ajz7HCkmpSdNhuJ3BXCveXW
TYtJNCsSUiG7BDzFyLnBq3M/ji7s+5+rTCbHU0GlXMpUorTE2KS+FWrTaVefCbig
Qmz851POKmIPuYTOZFK2O3sHNpWOR3jU9WGOlqPX+EMJTBfpSM+DOnsQwJZqYM82
jkB1oab/J+unvx4m2APtIfMLLG65eMk9V7GeG8yoqiS0YfBoE1WPKfpytJGq957k
Sbm9hGeWz7D6JDmUfSKyXOQkgnKnkiSh0KZ55Fx3IYmp685AulL5CF02ei5lrGAg
9A/+FKpBLRiy5NuDyJ7NnntlsMao2xq4YAbO9uo5K6yFS/Cdk1Hia+akds/Rliui
GKomRL0FgPXmTbS8mVZMDWNGYcsUQknCrOLd791nFNt4hwBSbleqNKR7Kzb3VJxp
iVFTCTxGD48bkMSnM5GZ+Qk2bz3eTaApRiEz9UbU672Uxcf9CJMuse4sbPe+XPDx
nWfqTJ9P2VKczC0IdkHxiDci2dz8C+xYPehusj/DigsHPdywfa2xjI9oQR5G993v
GDrLkyg3Xe4iHKugJhnEp3AwZON7HUr7BZ5aLNt22ocsXWPtFLVZVsFvURfX4xC9
54k1W8INtpdTrrWYVyTkB5FXhjq5yvakXkDEStcgUlMs8cjaLof7vG1IEla0McdU
Cxsu73Mrj/HA6HLmlG0xmLiezJa3jaXg2xjLdtHOVOR23ZSHZslKvjQDFUbgkkh8
/M7QruQvPRumCuPrsmTgbyFaOQ7WEwdt8UiMmvKANkzeNq+CFwMOKvnFx6NMpQvM
9XjAZ964o7PlyvRnU49s8kzWmy8On2+o2KyQIz+VDqy7m76tvDDeNDIgKqxwtpgv
mS2VhfU7sYXmMHxNmrp7T+h25sEreBtso4WHo2V4LT1WjXHNR83tsvzJ7LxoywIS
rpN8Ka4DANr62fjaX6ndRwG35kOcja9/GlBTFw5NhcEJcFv8dizcGeutoMZfmD7t
2gbqHo+xXoMxFWirtOKOsyBdjMRBVOcwdFJQ1OYWX+jRIEwde7RY7c42dSgmLzK/
higztFGNLmkyqyH3nQ/MMeOL4tMrXFMWa72s9irMGtFu5G1AXMUOzyb6t7spMnTE
hO4+Zp0IXjIy8/YYdIsTGHvvWYi1m7TwfmJSXdj9eItkSmJ6iRUY/GlzgKceAcVv
zlSkqX9ams20xtrBznOPMRx85Ak4p2RCueg3Ua/89ekjazcSNho2noFX3mygFFZM
OF6nm29uX/lp1J8WufBrqDv4GM46wpGZaJTBCjxqVDzcrLzmXqD4/Kf0l/fqq22r
jmddwulVgbHDc5ILwrBev07B8u1Cnxmdu6UqHZ1tgfIi9Kw5o0qYssfO+m9Loi0P
91VkCKY40+qkfb4iYhpF5actUvFkmg5J3y4eCo326BwDGdce8CzzXw0gorKJtX/p
xIqgyv1mlJOocjW8IVuQco5ywIKlWPS1wCtKZs7VrOd9sEF/q/pIazvfN/d1iL5o
warVOEDELYJodC2TCvsSsLofPCGQvWuIT0c6caP8//Ae9/nzrJ6+5rcHVCOjvK7n
F8mwS+4CvtnZwp4BMfoxlLmhPUhTiA2A/lvj5Pp3EHoZdQOS1EAt1QrNnHwJ5fT8
WP1Tn3mtHN/bRGl+fcteakNEADxBzNM1WBlfv4Ro6/1vdKBOzdm/SYnVxDVGlH0I
96ijy1G8BCkUxax3NeoIMcYkoAUdVfnrysDslaRcs48OxBrBubrIpCBTGJDYSUI2
wiw5Nw4M9RPp9WwmtEuXifReBiSbm2DS9a5KO/81sphJYvZ5FEA6ciYk4ZG4eTZK
0FFNfL2lStQdq+6b8y4QcyChJn+2imYzDZ4vvZrTnyV3f3RWk2vT51VWlBNncjR+
zwgyxGdfWPhsztOFZuFH43eoNaa+HlZrjEU1HXeB30CUo5p+x95EMD0YZeFLfR/f
1K861AnQL+66y4h9DIX9fMiMaL22yvFpVcAdI3YPPrWoqzws87vF7mgf92UdcxPj
l/zkFemMEXS/Rb2Ikx7yaIBlWODlKUoKsLweOP9xTave37+RCeSiRo7ZM3koH/Hj
WZCBjxsWuaTYZcgY6dLoMxuDk41l01BZvRZlLTZJsoX1/yit194i494NbWmUnmSl
/K+VO6hXWSJzedex6bM6C1DbLoyLh2x4/9LRWZAnnme7nIGJMb86Lh8GCLBxFWRw
lC2Z+z33rIN+auCaNKT0qbV+pFucNTmC+o6NvLjH70RH0OlS8pSqoeMUc87z7/C4
IhguIclWz6gWThD5HhjFYVg+RqcypyLH9WJi2zNfg9nVt3T5fimlko+Pmj4W26wB
d9lhOZRThRuqRCFh5MEYmGF9d6k1r3nh1ZYWnsHJ7ywNzFHmGJAB2sJmTKDeYjfm
ZbBJKOsj4lKHObOxjiOX465A4OXQ1hoR1T1eKKFu6Can4Finc/BaeatHtPZUtwjh
mszDt6ZudWGXT4w0miNDOv9XhjS68uzeJgivwKWUlXVBdk9dbUs2Ilch02wI5dNZ
y24W9HfsBGaNxtxArJWE7RKWagv+EWchokloqI+PkGbvbbIOT4F/oMM8HspKxi2I
CTL+8J+I7EXdtu5ex2XaqqoPNBbeUR9ImxBLTxMmg2l/Jzb4asJwmKIPj1LGWM+K
saqVe285OLViwwf6yuWMhVQiZNLm2FBGNZDOWsilmhrq+ktzwLQoysMvk03XuWva
h1GWW0K8sGaHtC3erzCnk+nT3Zlxt3OHE57wU43GjemLTxNAurHE0nLWnn1LwopC
NI6/tP8bPwOdIdcHjrXF9kpkPRoMih7Zm6RxPwXQ4sK7pVAXFGwKymerWSX2msfO
v7c1U3b7Pr6Cpy978XLueO1WtBHow4N4V/k61uzC7GFLtK8+JfA9G2tm8n9eL2/Z
RfyH089achsw9AFo0mMMkLJtCddbRHGO2k0kuhy+fph9WP9y7vje6BlASNymVKv0
OKjJJqpDvH3ZTcz8vuw3sYo3xgkeush39/rgjhCE5nuKrfDUXxUoABct9fJpVOSs
84baYdnOkI5ZyMAAz8WfqmDNhjiFgfTLhsBwa4mmf6WPBz/gV7LZGFllGH0C0lb+
kl2ZD3k/ZHdUX8J1lyvOXSPLxeBzHT4R6fAfMgw25Prszx4f8KheZP9BuSCBwERU
urfjbnoxfDdnR8Lg7+qMiC/KN+NCrnkgZ1/G14szb3H5xBsWJJNONwAX0BaLdInc
8sdiFp7Q8BtGkfW97yZm9aKfwLWhyBEXwjp2RwZgoAa5gvxQULWwgkYPatYlRWHn
+/NXbNi/sdtiCr/11AdRchLooGgOZ+zXYgldbr9M7XsltjqEBMELzpRUYn4f7jCP
fn8/olKVoiKh38Rohtim2XIQpPMrIpdwSJ80E9kNr5uUclp87FoVRXXEcFi40jXY
E7R9WfJdVfOngwOUz0mV4OTmpVcupcr4U2q/qu+0l4o+Fm9q+SKNdnEw+s5RaIKT
yKFspGvocbDdpVeCWAtOtL4eXG5rH6chyHswi5OHOYVMnZ+bLAY2eLrb0YzeJ2NQ
vxMVco3BQkC36qbjT+SoLmmKuA5R0Vhbu3CyntXeFoSGJ/vZnfJO63jIQFcparcs
pTD5UrY5zF612udpel4I5XnqaMqQRm0drtsL1QskaZbB/jOscCkjUDH1Si/z8Bqb
gd75G6eNfO+Higg+JVzhBQhUroDVqHPYZjwQoHzq6LMGIuDD3iqmoNM4aUgbuuwu
m1waYfs9rnNHCkvH14MNNsNJKCYOL08CYYLj85OEKDeKfdVhrzCRLAbJtP8IquAE
I090PU7185XYUxhSEukt0HpWgo+NUNky6Q3FKaLbS5C6x6Z0lWBCNyFFOvKjWQ7R
HJLi/PiiHn93YlqBGhAGAWBC7fUrXizkCxe7lLMc5rV434JbyctIEAy2cOgMKBAC
gn8sRpj2Omsf8j12qy1nWrllE9HzpRxqxwZDIPBxaY+tIBIJM1dUmLKk88hdVnOW
LL4m1JAFf7GP02Ddekec4z5U2JS/5QtfmomtP9CevYuh3kVwNBlUOsiEuZjA94FD
BA5w4/6ZIehjSbM72AkKZR/AT2/JreNUfGsCXAYRVPduAmO+fKksXCeWh36YEjYd
3wIoZ1fIOMkUKj9oD7MJcM+Fbyr1j+6hf0U+cvKyv2cpF7Mm1g8L4b8tOcnfQZ0d
ctwvBecJt/NvyFcTWlWlT++OH4HkoE0nlFt2jFfSB3z9ScnDQ89yc5xANF34b0PE
a9tx1toelfQ6iZg51K9USfybkw31BX6TO99/lmmK4KlluoM8XjWzXQz5vbmKTvkK
moqXYvezPgREstuXYbpVDskUfTvImiVw/eId+Ozv3/esY2dOCdz2vlgaBsR26ccb
7ihWwHVUeX5+K5Hbd+Ug0rXWd31Ij7VmD8U0wBSMXDdeyPZDABzmqiAsWbjgJpfc
KcLMXlUmUu1GfW+nurUxNYDNaypPngijSu5uzLMf1bQzMDhTmi/ZSzoQQVrMWoAR
A6GH2UNqRnEzNsCu6/pNNjzi9cKHrqsU2WcxHD6IEMNotSJo5Sja6UvzlR27GLgA
8yeRdlVWxJbsPp94rCnAhzOKDVUjfIy/61svUFaZrmCfzEMzSp13Gtqt3u2uSy0N
x/GkFFps4DhqO2GFYWWDhC9I7VJ4SkVKdHcWWy5UUxhw+t0LoUX57ftCPAD1Uce8
6uy2WuOiLRtjQpUGOa1GbvU9EvYv1jJ5MTCJS5PMWXwenDXGJQ93y0bCSNz8WwVF
cpzzk495UW41NF+u9vbMC9pNDnh9eAEx0dUyg6cUUChZyqWqdu+BO0q5XyaO/vTU
vcxNoIpv8EUTE4TG8LwwJzW4bud+dQLabwpPjwBJ9DUgT0pdIcBzNE4bhof6npKW
uuwW5zvD01dVTqtewV6vhoGoY5+oLm5bKbQ7M2auoxusdk82fHv2I5gHGPIZW52/
r+dZVgGkdVm1kjk7VP+MSmBg6tatbILhlVjI4xqgLfTlTqMjEt7GJbaT77uwRdIK
yHK44f/G/7ZW2hu6zKp+sECYwjwaKTGfEn4qW0vKPw7YiEDqdNqNGrfPqTiFiRWq
6FY/zDSrOqAoq/wRh81wFAN5ygemmZU63OKo+OkIiA2aeQacp2yZ0rtfpDnqDD0z
SUyo9jfIsYJ/7pUGUdMgAHCDCtwccCCKGq01QAgYKXw64mNMfUvREGQ9/tLEcesl
qhOxKcr2VD/iREItWWWODVUNvYFb5j+jxPy1jRSCTgeh5Y5XzAXv/auidFEiccuK
NrgWaVxS+IY74xnfLpmuWKHQDgCFeUOh8FkJR+TfbI6RI4WlUF2NqxahBXrmFMe8
SE1p7/fKWC4vVBHKeqaNBqD9y+/wIMGz0XWlLDI6eIUDtrxNXIgGSLUmmKeN0+Eo
b23KbiCrkvpXXTjF52gz6LS6t/9IMEkI5xeiXTtKj8glPK0Gw9gHntWn08M8lGDy
hz9Y/9ih7nfymS/VKJ7ynjdHzKe4KcdzCayqhaOvWTdNHa3j3w2KAUGIyD3LMkxI
5F/uEw4AgIAapikPRzwNDuxNWF5e9HLXh7CPOcikgxW2yjRhclKcWSNZL+G1X+rW
sTt2TXTCA9kcwuxsiUp6nx2ntixpUY/UeVKtSGmvS/8j12IVRj8tGzsfdo5jsDXk
z9tLFcVTQoxiBRXGitk05RYB0/yTIgs71Zn40UcnLYlEli/+/bn6L5DqmeHTa1Om
SAwAUfZqSgFSYTCxwPwyQkV0iL6TrzycyR0WtK1YK0yS3ixpJ5OweCL9OdArJ4A8
va1XgoHbARTOZlL3LeL2vgerPruyklEFqn6kEI+bWj97AR7IrJNWUTo/2QypAlGt
JDiRyvyIrVWb5dGkv0N9vSxP+6Vh+JYbwr5ravlTdsn9InTiDZgYmdwhHh4FC3lR
6fMdmugeToRBe4JNazy2YELadz4N3eqJQd71mq2pxX+fu+fjs4qVcYx+/UwBJePJ
P8RS42o4NV/iohPZd3MflH7QHxTVwzxgC1eTWJdJzWWVmsV3bI3bXjJrOED8/K8O
X9tKqRhljB8r0HP16RanbW7FKfAMi+jSyYqJ88q3O/27nZZVVXvTyYXiA5TJnE29
pYgyyR1v4R4svZxvgHqyyHXE74Vw5kTvVfomEH5fZockbwCedjnoEv7nE96+qJ4L
UxczZWw4Xo/1apkIPkNXgtwsTiSqDbGYKiLKHpnYrpb1OXZEMvHkLiiBWXMsWxGi
dam6RaROQscL7okbos+u/0+Xar2CJeKj49MkuMTbmkBBWCwnZcaBi8QWx9hfCNFT
NpSYRawZ0WW+1PnamiZ8t2jJpSZvzziHqIRqqj/SdRwUfUVClFdX5JFbHc2ZSu1O
UJLfnBh41UthGfUUPHjmxcVlBg3DMoHtwxO8MEC1DK5MroOkW2+4CGB9p1kxJvvk
9WnN0hH6ayRsajOLHcj+xu4z87MvSA8xNvJHCPJNsZ2UAHAsVtOI9h5JGEK+Y31A
QGL5dsCuE6i1QNWMlhNF/TuRJDZpn2CmHGDJXh8kSQignhRSHhsWRFcwCKA5gxFW
cw6cdPhin/to5LP6F6SqOPuCDfEaC7Y2xSGboJg3upQXB/vxW4sgc+QbioOCOc3Z
2KTAE21yj0GCyfDwWaDx8a2AqKSnOHi2M4BC5lQq6NGQAkTEnSt8RTITMWxYID1L
NJ6X6uHbPW1tTmPNTj+PYatWw/ik89K71zd9Az/gVndUHC7+awkUz01id2xXPtZx
AAeVpHACceYr3vgZOgMGHen+1HxhfNowEucdgCw9uPHJZYenaH7ccSVt/KJkm0Th
E3CSVwdfdy4r9oVM9/Syz0iSY/kq19YPVvjQ1Xwbd9i0bY2tksmZEhy3Q1Zux+Dj
3bK0KP40CbXwZHAbOpjnPgua9I+Dcf7YxBgUv6zaFj6fT+vfcQVoUIXP9YoDEecm
MzAem1ndqO6I8xxvXu2vuOPzv3Y5ZggWiQE/J2/BPDkm9hS6PZDjoKWx1S81NyCK
9BhRgTMmmwbBhZBEYfNFcelMuF056kHsc4H4wS0lXqyquvcl06fkewbFID8dVAZ8
X0cjvFuB1Ntp2PXUEJxnydAcRnJ/ypMjGHsczw4xsNwV4WWNzwfRFdWvAz7LO16S
Su81byTPxFgWtv3FKkHodj9Ib/HldTCd5P1jxKIYmA5vAWP/NfiZDBZjLIGRKYK4
qtcxzhvmVnv/b2qvbibM6H3jzrq1Yq9WAuH0HRykoAF3OM20f8Djd/VNIrICbxQl
lObuR8D7uDfzSz1OP4MryzxM9iq40WDvG91QEuFuOAa4w7STpqE/H3J7Eqyu7lpW
zIbFW9MwTn53RnscW1OnKFgnZ3gr7O3z02ZjsVv86wgcHhYEjcdu04+ptGyMpHM/
d7aqz/5TRqh3QrLKK8Tw7m7C+ceBEJZdB4eChnth8fNhPdJjMHG3wx5AyOAGtpCQ
3NmN0sEFuu+wPBEiyHt4l1kWwyKH9DKxAhFTQ+1LDvf9lsDSbswVzhkW+zSfIo1O
7wFi4XSx77qUiGRd4aLbmm6iqeqNB9Wwu4Flra85EzgtR/BuZkwxgXdQh2t/HBxb
yGJ3CvJY4AOiiBMYTL1ExiSvT2LRbeVSX3pbZObM6R/lOoaYgw/kjFKJtgOqnCVT
3m4CKcLOGOtq0blfABvNPUxq5QLYKDiahXkVrVX+VciqLgAh82hZdfjc2zOK9Tn0
4lzcJGUfvWveUMnF9gcnhOH++eYFQWUjOVgsTkEhS2eykcMna08P2aAONlMFy+AM
GAVpQZQerWrFB0ssSh+Ady9/yndxH5GXXMEKLC0L8Gg1XKM+YntrWm+7wuBH0OES
gggthOLpoqMjGeNQZcBZanrr50ScDJEg+I+54qeJrQZwl9PwQOe+I+4IDMsUM1GN
MVQctKNBJj+yTwYJi2EwylUcVff102MA8cJ/pqyTUfXuYLn2KwBUtQNcgDkVA0cd
mU/dCgXDXZnNS5Glw8QYXuiO6jLguKL7yspVAUO8cwv70lHHkuVYFbLe1jmJ2L2T
5SKvdXvJ10AxxGkmilByDdLZ3rpp4/cObG80bGWR5XK6Ky9Dud1/7GBfW20RKtRW
iFpwla7XXBtWdxb7TZM/xDgUjuEzfbTvzQPuLxpCFrp/T4ZjgjLfkNlWr8ju5mT4
e5e6V2eYQ3mNE2sA3IqMVmjNASzovT/p2tjJwZpqJg4Roc8TFa3XYg4CGpQibBc8
414Sd3iir1kqqsp2gIr1WaNF8BjhZ1ZU5Ylq/7ccrKqsPM93fynZUYIVoPJyhL+8
f7DPplukuyX2xUIE2YofclcZTNuQfeOYM6+y5mW6NTYr+KCuJrXK+2QayjGIpxIy
voLRfVr05BOgp8WP6ueIVSdDaPhNB7tvaDip26jg6ETdhoXzlX7iSvJcqu8TKnln
xg2Yw7M3O8zM9NkdxIbB+RYS0MTgcwnB6eua+cO75nLuknMDT1K1mcDQ9CGJAMdo
Z41HbGwQ3Rexu7iLwfnUng1aNRBk4Wmxj2BHdMf2kRHQqO/aE0WX7is3RrhgJzgG
pt2kwz9FaA4kMj0NPI7h16nX4xTUV6IFIlNS2cnEjc66d5JG25HM4MpZsZfJvl2T
yBU2mQavytqH4NqHHTBgPXjxOCgIbKydHSWjlqkBK8H5er+nqYLg+jTLusPxqQaP
8Tq2oxNg+hftmORoOn3FWCHybDc+XdXUeRo7uOkIb9RTzjXnV6DWgDPHW+N0Ircp
GJtvJYBrzwpnghm15AvBVZQNfTXBPQzw0c95lCWH3zi0VpLAohbRXPtN+Z90kkaf
JauQR8+3jPJlI2nkQqJ1mpQUkw3nCoaTT8FRroxSNTOf7A8h4y2xdV+9TxrZjPWc
ibcGC9Reg78G08ev0ZxEipqAIwGg5USY4uXNvAvSekFG3RRVIvZQ3EBabdhiZQ+y
ja+FQyATNqfB9iBZkSONusdclDjzDsdFo2NrqunmPycIATBbzbeKdi3TZkNmWEWA
l5o6MRW4epnTm0/2aUSa/CXvJmXtOsBoiKtD6g5LpeDFB72pE2z4Irr9rr6AV+Qu
Ly2AQL6R/sOa4aADQUOm5xNg6gpnkxHmTB3NpFMg2zYdN+omwDptNo17qBSRP8xq
fbaV2S49lcud42X8mdL4HgsrPFt0BO+mWUPEPyrbFo3g6CfhT3Sc27O1Pqo0CaY4
9Ds3fn4IMmbE+Af1Vcr+nX4S+I1WMgkxCKIOBeBjxfxZwGekXC0Eb4DRLNYKFy86
bqwA0Wd+11cDoZiDehdMEMo9cCS9ZQ3U/6zRaG4QYCSnH8VE12moGWWKdTmnCfmR
+jgBjEQm5P3VbQXFXo0sDBQNM8Bif4tkxfRphNa83M1fO+uf519jWPM/L3eIeDtQ
+RwlicwzeXFp3iCO8zoK2lVQygGj9fRnPyMaa/6X5vsHPNl+iF+uBxTMru8CfkY2
3Qa2qxinmd/GIl3+vpLoWGWrT54t91Au/YRgkSl9ZS/0vY5E8tCqJ8anTwqEnq/j
jAYShAhZKngMtOg5isT5FLVbE0tTt7iTgrZQk7G+ACuHG7tKVjv215lu/51xLXl7
90DfYQKslLKAP8KI6iugywcw+tn904Lp+xoCjqaMm2UcP4pF0mMGZfJEf6n/T8NH
nhmZ9tgNAhxjd65LlVMW2pUIQPYhR2KGGsk25BVy3m5BNFL8fGVx/O/tjLBy+e7P
UILBN5IHxPTBE8O5z/FvB0yaAEr4PKxoPjLrsApOfEjqmgD0te2l1Ahoy5I+eKg/
L0tILd5vFCsPOvPQSTGmP75EubG9oq08ikDl7sAu9fFvWe4bx1hrbmUTeXNjrXwP
/5gqcn5Maiv0tOX5qsZ54dOeB72aD0kPWk4ddZVmpvg/rgFB/ur510YXJwLLEaI9
+nrEC3Ch1FKwr1CB7eccINgIq/RKUHjWcwRrgmJZ3TxRHrADhyNNqImUi+bBiX/2
iQLn71HPXk9PhF8pCsfisay8C5xqDnRV0jbYqkOZfEQpItFGCCdY/HuovPfgNpei
pABaOZ++iPOuiGbguWYz5/SJlPdwIgxQ2B4sv7Qurz7N2oztgZgppZY7OxSMmsjA
NyVN/l97fhMzhyDMukfc2RexWWu3PBBMDiChl7a9S1F+5e4WR/fdyqHKbYaybGlp
2I5cxZ0zhRxLyqQJHy/cHni6iDhjrvvZB6JnaP4yW25A5m3B0YCmra/G4wEZs2RL
EOShR3s9urnXy7nElrGFCMyEv2O1dBelilJ5Uw4LfA7mTC7XUeQnzZ5IOWf6rK+X
JDK/6+CeTmHCMzEO3lrEYwbEL54bhqraHLEGMKIfJEdAwP4MYivn6Uerisn0bauV
ODWo+tVD9vfbou2+MmEFEBNpwKRNS0WfT4yIapl/jrfzbyC1hgM6bRLDWQYNH0rh
i+/cKR5dCMfIFqN8Pz4KnUkxTwBihFr23nYPEX1Fd1b3KW9P+mkUTZme1MEk8xzx
1xu0yq4J9//QxRWnsP1l+oYa1WRX+HNNqEPkiHtD2FnDcS/AJi5Zx1zzUqatXE7g
x3IPePa8RcWt/1q7Dwpf1jnUYcY45yfqDClV/G3kbbdjvgzrkdlPqzcVVv5+GP/a
1eHsbFNg/FdJuLzjMR/gPZabVcyB2e7Y5G7mfFWJeMF4OJcRXWAThp3VcqrDW4+K
pW9vQz2yQRX+6GAlvX/piGNYqMgX9/76WRjjkKIA9KjuwABhppNahvi4eZwPNKpW
QnCgkccR/VkttX3JRNE5MM12+v0jMWa1YacR0S4ks8aAwdk8/hzV2ch/j50LgnKL
DleTpH2sFnG3hdEl8v/jisukYmbIJ7Y30jCPa29NeRqNg8XY191pwJIGo1mp4xfU
vf1m0zQr1X6ggWwg/k07+xFmK2pWFZGsjQcT+FE2GeuOhGHaglrFdviEG3HWYkNJ
fGU3CcWjzO4QvFsX9bfWrgxaFMRm6Q/Q2CEj/YqcnzX8WvBUX/ypYYk8kwnByDK/
13obsQ0rThcaRO0imfpwuNS4KlKAUjIBgWZUe52kHlabs/VH8Cw6u7g9pZSqLt85
B8ko26swiU8aziE4js7fL/ErTFGbPzeALeSTqYy/4ioA9HbQL3fPNDGbopTcTe7Z
w05cSpKW5mVQ746zFpq5qnvPend9jC8frJbn53KGtOH6SQ84Q+HlKyP6kgUs3aq8
R/kRhiN18R1S9EHZtg5VF4/9xAaDN9cvDGgCFdVfZuHmPb7y6/zQJPB8RrZqpYdu
mUN1+0dKefvoLyCsioulgsK2xIMzkB7MKhGIP0brSg4Iir3BcSa32azHN4LgZsLv
+iBQZXWu4c8eoLcTQIrjPDfsknj4+tef0JIwqDZw6LspDmsUTjYUvr0HZsX2RnmA
gKZ+hMXS9c1wUKHm2ssShAG1IdE2aDlFV3cx1S55mzJwBUZOctqR+QJmOmmR5yjJ
jHEFwLUnxktfoPL4pe4Jhdd1mFCtrYZ0FejsDVhfbakSWnAyVxKd22xKhYOKz7su
nRbFlXaCX2yUP8H1EXBs5YLmCH+iGC9zBK7TmubfOolPSZQP2Xl3DoCp5dkSta/e
TcaTQmbFPW+RDg8KeQ4rLRgRRFUwi2KNjaTiddq3sYCmdTEsJozj1GKRoLfVJAOa
fbGdFPGYyy36uEMyfP3ftIlFWrRZjUQpwzcWePcpXgTlshis/7UGFDFq7Ihy8cQb
eSalvL2djaV+mB8qdLxNzOluIDhM33/3s+Dk9J1nMw5kAQHrnvuWKHa/YZxs5Dpe
hWA0vvVl4YzVWKJpu662QVNRvNRlvF79oP06jErpHxeMSAYwiHmuEIZhsZJYSvP6
4zAWsoQGWkn6zKt7Lm5eV87GQS5eoAFRph2hHQg1jW1aRjFgsdwsI0YpqFQu9lni
VuRiZYN6M88L1KcDqGApkjQZSXh14qKXWY1wWvPdttWVwW9nYZHTQl6/timx79ti
4evR1rajqZbD/epIXSn7z/PjPTlEQ1AJ6EOhrDU6zPnzAXCQvTB+yweF1CIGTKKy
HPdWN2NVIIUUi7Qhgpv1tye4mqibfOgE9z402eJqY942avpjLL1zYd6fyXeaI2/0
mrOcJnPkTbjatVpmutLWnHuBnG40xkY1ciU3gtN/kI4ZzeUfujI9p9I5ARLjtBSo
flrrs7pk6J/keUJfXS6VO9wvSHBER2mzpBB2EZotiOqBn8xOPFZkXQaIZZMAMATR
77rryakmFce9OwwDX1PQk4boNoCR2Fi9NgxNUmepbNSngVwLo21X9VwwCAmGAARZ
p51g1pgpFguDq/IkP07/iv3gjzpFGO+ACXhAB3+lF/xse5ZHwbNh1OikYhxxQ5Wx
sTnFV26DMv+oq59NwIHPQFjNwuBmuJG+rZnnN0EuM7tCQww4N6UxvMSwFw2X6DTh
xO88UtEfjXmTHJpAxUDUBZ1kNOfSFoa4zNhNmirWyP9wvoWlGrHBVLSJ/JuogrSH
TOYul/Wp+wavtkdhZ8HlJ+jPMlP6GdRG8NSerdIzTDf51zBIhO0i0GNIhOI80+sN
2FU6EGP0O0iT0goI2HTSZUGpLyzBdHuj8/IxnXPqU3/XjaZsnz2dUROPtPt8/u0s
OQLkgsi1dyylj2MRwT5174tY8RpRH2FfdlkZiioL8b99AWFiqzm9rGqjqqKXrEDO
iFij1ch9Y7MpqA3ti67OlcVSS1l+bBnb51cHb1fOC9mE0LsiLeVOE1HxLzBAHKbK
K/MmYMHDPW0RfLw22xJEYsxwv3N1C/LQmRsNW0+boo1DRq3T9IzmtkWE2D7G7k1s
L83I9w/lp9LyhNq0BFYclj31ia9t2WS0/zOng0WFPc2RiFXYaegP3mpWKA0Cwgr0
62G0RdM8wSSpVF+IamQz3l2E9bgCuzbVg8Tb4HFqH09QAnu1ufu+UYqb2mK6LP7m
ZGcwZNEUs/1AGmn95xxRVZNu9sFXjJJx+wD5lXOOMl4AlHf8nQELaj502Qniizvx
rN73Pp78b2KN2N98fBU7W+TZhyvLrC7ZHKbjSlwcLEjy9Qh+GiRlph1UUAy8/9UP
26bjGkk0l3vX137tPyT1qIe8MOma17HgYEvfuIw30LkBsmOeWYu6+z2zhEfFdbZW
HoSM2LgC310tPLKIkCfCcp0PCUmUg+ck/dz6KI9Yo1r5jNBXYHzH0R0pb/vs3C6i
milfQ016SRFctNSb1nc5YWtafoB0aiukr7NtpZANHXR0WgWFLJ4jLuGhGPRz+51G
LWenJn71WwXPqHJ+SRf2Buw4f3uJ2wkvjtS2mXvPkmspeZPNJlngZKDaUeziw0s6
N/CIbeNnIxzrtozGhv+7s2xdm6rUS0Z4+yiUUbPU2TrnX22xBfoE9plhkmPcd0zx
u8V2nheXcg1QYt5Qb2ojEh749Z+nkReklgfgMcAIpJ2MNKSeqMTO0vOG2UyYO3Np
yvr62Bp3RpVupYIHLdVqah9Oh/Wl/M1rR4LX0IdFNa4X4n+9stZyUjMp8tTtFNK4
7qA5M6I0gOxEbpbuOSOZAFl31zPKftIoo/PQmj9YGlADHPrvMUngnyEt/n6u538H
R+guAwzg8lJN7fpwO4d0/DS1G9gh/zi8TMfv/HZVWLVJjpqqL9Rk1l5laCOAycVY
uT6YndhhiHZXVUJyxVBO/YceU8JqDHc0mdJoUspoUFgwEi8Zog055GGiiHMHoiza
SzNUcWf2ZKRvbKRMxdfcNGRgsHMP1CxnxadTGURGL2WBapO1f57ARstOjJTgn9ns
imagxi8ybHnJ6SJGmDEnBL/GoLiCG1NO9Rg/cl9K2kvvPLAfZYRxwGSIaCUY3bYL
IbcSAO53liYomg9ZOVRz4BArUQEGrNi1n0tfYoEDBmkfyJ5Cstpt6BQbDaPGNkDQ
v5u4wYeJoPITlhVmrhRm7OwKgswAmlfOxuH226Dsu+AnGS9j1FGMe/r/l1vvjHY9
bnSQukNr1MohVjHF2TTQbI9X+crZiwCPm5oQ3cqNiRHTxe9oaisvxBtDFdSgdS2Y
Nu9dyjdNCvHWq/xbwr6wLy8QP20o0AwuOmYZmCJPfu8RK1wQr5VhAcQ9WCMHLmhU
fXRaMa2g389n+N4VUgSzmAfc8KJP3GUJbzKpzy46rfZZ4lf3X4/B4GV1Iz0/+luG
Hb5X++ACCM7IYensvw1127/b7YftseknAzb7mvq+iMnfcTsMvS5zoUsFNgl7GJEp
uHUkhLVvZC4QXnl507RZTYcYatF8bhuDhxoWqatClKfq9pFmH+jyOzt6tnA4GBi2
F/Aj7OOOCNNcw4G1reyzXvIbMMR2izDroLPmviSsybbqMGrq/ZLOS42W8gMg/lp2
f2BlY8PYgUQ3r/TlpCyZCH1R97eUSw8x9iVkWSwmYvEVyS6a8LN2li2ewvnamrWX
rjlsq9Wrd80x0wi0QyWaOWxAtI+F9Ho+9u5QFTCiRVzJxMqFFECyh6+879Yipnt/
0tpjE2l0cgvCfCwrggRpvJS8P6QMxdHprx8eQFmzmWAkVsrUEbeJej/20ZMCY5T4
oJxKJlc/aJJxBtze0E2a9n+aSbBMWyq1aEMSw06gozyN9WHYO221hlx5gqFmxBzH
x76VfBbKq2t5952Svlnc1Ur9+YAiYwzB3mTHN75ySQ1LlBOZK7wJha9WaHCdjPZf
+SA+GVmMlJkuc/h0XFr/RfczSt0O3ACV4hlr5YlyX6dECFKqeMBeHz1Wn/mLYnyz
JlDGTONsCoyUw/0TJ7fiYE3OQEWREpLzpOVHZyPqjGkQ1z9SLMATcH1Y1wF/PUI6
0WKPyY8URsMt4kEJH+i5Zxvk+MB6IkNLRjaVTnTyKOz76dxtBPYGTDlJwJOMo779
GmcDbs6PqiTSby0eE7h5qZG10ucfvMYH3+OHl7vYNkGy9opbwf2E5Rjs8nSS0jN+
jXoy6JUaP5IYbiLCGNBgBEqwscRAmM7dObBC1tqMF0clk+XRHrLKaqeHO8RAgfHI
Y5US5X/X3LYr5OgmL3+/FHCfrynqtabaX5+eQ8xIbT9hI9F1324s+ZSK/Koj6Zs/
hc9fEvE+DkhANxP9p2cr+YwPBn8CJhzdfdXPu/6FJ1vPNxIq8l2QLNYtOsoE1j9z
Bf65GT95DQ9d0WSKAFdzxReFJz/GW937Ld5T5keiJxtSpdGAkfdLmAWekqNXyFGQ
xfhE6jC+EEKAlXXNOtE2sjNagaFI5EelcOwfKPpBkhCtuZTwe4ecYdedPwxIcP5M
9UbZE8Za5NQfiCZx3d0p7Kwus1llwsU0TUnjvKk0SW3AAJGGxI2KmUdNIaPSevvt
uZ3AwkCurbP4hmou5fIolzyfovjXu9lCi2iyEZykwASIgOEEgvho+w12FfOoDBzz
ivnLmFT+V7X0UD/OZ/bQxFvdrABS2DAskOeXeBVdiHkoy9AUXCMDnAoqPlMSdcV0
oqDeu64niOCMRPtsZbD2EFcFcOlqGb0Beb+iH4kfzG+JxSMAzLvfWOmZ01QKRSpr
l9vqq7yrxp1KBPBtkn29T6UYLIiKwVNkh2s645vObQLxjbq58N0RnkFgH9jpgo2P
5VJpz7s2N8XIvtflmtv3/cz//+XBU8rOqE4gJlrk4/Q2Kkejtg0io0QT+XBetbMs
ITJq8rGznps2Ybk9T8k8PItj6TJpZA8BlloMUIu65/kvfXqqSQmFyPWnaOIrXH0G
t/F8NnAHuvIdQw7snXdRcNQ/tLmhdkcZmgVw9/z13agJRbJmUSD3JCQIYv1db5c7
+ovcG3XzV4vu3Z0VIz6Xr8N9h2spx8UyoK1DH/CsAdV+jo7u8Gsg/OuJZJxBPLF1
yXU5wP/KiKaFfW5V/c/64J++RiSXxDrQBvPcth9QPZ4YR4r+DNcmCsxiLBAiFNLI
0ITRS+aerX1H2sO97ZW+yKznPN9ZxDP9Jt2vVPtfObUe+m7e4H1r0Af4Fmnjd+ct
NwDwSj6GbHwvS4aQN/jxYRdO6USRP4WdotuYY/4cz+vHa31JXf8rOcJaEcImS9jl
5YVH+48qbshMrzQ3wxjr6IW/iyE0MkRWB4mSBvbpoEqWB6AW7vvCHb7nhtcPQAIA
k+3UysQgsQc7yexApuxeYMMX45NK4GopPOAK/t5G6AeU03rsUUcCNOqp1VAD4ehY
QLBOfixxc5r50l7obIu3kK23Ia27M/pkydwmQ7i1sPWZVJpjMzQk8eeKsbtvA3Rm
LlKnOcyqnfDqD+K3qBO8Bc0SxohCJd/yg2KKeKqW9VuqqxmtuRFQWo84XbTeVd6u
k84mGuhQAt9ITjZPm79tQIkfbM9OaSFeKN45O2dLWYIZhJFdo87zZqdB3sp25t1o
NZ7NTiPfYNMOfVRPDUjGN1wCWnS/D4jfi7DIYOAu6cjanJBQ753y5GEu3zAJV/Gb
qPaDHlxmX2Nl+gO8mMzW3lKjt0qfftDzd2XAx9AWXm8jnkBBC6IUxaG6Y2W9AXv7
MV9j2hteow5OP16/1PRDpv7AcGcWyD2BvsdDfZitdw+OcC0SgY4ZG7JsrkjcY/fn
wUxH9ZfhTMWh0bSfP5+cLjqmRiK3GpDQmUnPY/Lzic0IUesIRQHWu0djpNjMZy17
i1Pcv3xuZl1V9xqtnTrsuiMyyDbAVTN6/BmyI10KQmr9kR04v68Wo1rS8Ny3PHTD
10FzZXSbgugG0SMIKiRwR8bcxfn4uFtUhknUQlg988KqrPxONzfYK2nGxRqWMkj3
deNms/49lOcUjk895JmDPNAAdcjTmTCCZK7MD0QnfEAFAa+qljAP6x52vgxyO1dt
GMRNHbspkYOdbdNl+NiZKcFRxEYiLQ5FN2uSLbvOPLFuOou28b0aVTnBuBWWIFtU
tB2O4kLnIRJPsNW4KVMg5ZIsY0/vqAAmqHMdlfnbR4wEQL5GOmfOMUOYmpsXvgzA
KOASYN28xPnVb8M3KaTjCQdOHB13Y9oGgOdlSdL63eDpv0Jk1HvAjxbPbVpYSjng
o/ynn0TEsphab7hFjXbS5rJGYShDHMrO8EWYr9ye/KmfQdf/+X/M++2L/njQu96r
jSbkaWc66jtGBjE3euQxHyxCDITz2wSUI5TXOu3286dBeDDrhj210xy4vxfz+ZsG
ikakKbZMahJbvl0J/kcJrpQVysKyKb8eJ1Unmj5qzBaBlvyvUVAwpVxbDMuGtaFo
8ILRON5VIEzWjQ9HeCFmCLUNctCi6wf1XgBLMB7/Ly4s2IiPbk+b126shSGuKVKQ
oN0BlmT/XtqGHzRl30+2js8zn1MQ8pzcVsW752LKcAX7d9wL2A7193D3CsKYEcS+
nChuOtCiopMyga+T3DQd2+I5YuA35U+RWLQlNm7NyQO69oCeGq69yYkC33MrnOvD
J7ZeJu/H6eT74n/rnrAJu3FRXlqmHvqqtas1HvOsVkbwisdGBge3n9UzuSt0SJmg
i3bmA9iJXj4qyQAFoYi5j28OblagRA24S9GWwyKA4N5acofKjdkzeqpiTveFYVCH
rPc/wHBciZrL//rBmObOPIrxC9N+HXxUxnz4QH+5JlqfQI9Kzu+hr4lQQQ8no0O8
tAuvFqmvtg4bBNhOKPnZG+UiCED4ycHcaz/F+wsX5lVyy9nMynvqHlTeIpAXA9KB
X5FdLyQxqPUkf0z4+uaeJ3MXZJJG9l315ij9YFNbOaNN0JZKl9Mo/n4SyD35crl9
uw2VnIjDhOc23SegMvxpZrDyP3FBiENKRlrpZVxEWiqne6mJtmtsHMo/nDT4fNCt
WbpJWfDh+4lCgPxKNWrqIkLeeHbtY+g7+vycGOJ6276RtAjtT1vW7jjxoMyM83tc
K6XYy7jqn+ZiWt/XKXG+PuBPIeFY4mBfHkBNMJUE4UH6XSxK5VWe+uM4pBMMB3rp
5+KYTkdK+4f+22nuo7rqgIZVE7q2wCN/aCyTvR5fHmrtqanhw9E6HZe1E3i9d1xy
ozU+/LRyTGeX/0h7pIBVs4d7gh9/Wz/ovDNMJWlQgHuyBRiOLIIpEY93CTYBuJOe
xXj7ytDJ3E50E/UrIGClSl+UykInNfdFejO+iXeuYmUQrmHfJi0AfHA9ATAKT8Rf
GszfLQ1l6hRzSDiBdemU8Ci9qNNRiOEVlHwMzPkj8IXNY5v9n/gTLt8qq6UwG9lR
rbbNMNV6kEzovjniOlLMJYSbZIzjn+nWvryM2W6T9Tq8G+YGWKL3YTtBf/guDOQE
so191elS6uSm8BC/L7IAGbuz9IHf3qQMbl+Wom853UjivE7rZX1n7Tf8J16VUm4X
PlNVnNx+aLe+7xBzjD4zTSZs6Etxls6+MoKIYtM8nJ8DNqhP3IDGK2Rst7puhv01
nOcyr8dsNR/N9MrHuCkrf44iuJTZJZGwJS2Sv5Qm1JJX/Ye/pejjNH/fqKfFS9Uj
Sug1dVvOaRrFE+2dKOeRkYCS6PQ12zxUsZLCVyLwLCQyvKo76b0Qckp8/4A4uErJ
n7RzgW7DdZMzwr2cJogoAKm9AWEta1BIm3aqLRgBjbdWB8eYSSh2WTmRT4c0DbM8
Ft7TGClfQUBkKwfOauyQU73cAlASgtYqRJ3QQdM/2Ow1yLK9WtMemLPcE090Pcuk
8cW3LyTruJgFR+9Jm/uwidUlmBXPAuk+knw68NBv1mjX/69g2cqTq1ZuG0sF/0DA
n3UtyfXxbYHB1jN+pR7ZWcUZ1i4nrhP4VDy//ef868yz4Y84npz7H2IX1+22jTFU
1gqs0mtQDIJg1eE9aPlPS2qEU1Ec2SMH+60G1U03kx5/jmXbDQUY56a+8VqVpBw/
6pDaQO+FwT/yJfafr/PcvPtjHIZXnJ8z3A3kjIMJB6exXCxkswVbgIqwvgO2eDwC
/P4/kiygF+DOzxhbYR9+BvdS/2tEPgr62PM5HH5kwKhfUjON6GUodJr2ZC2X8k6a
GrttxFYmZeqm2AGLKV0hJf9eVTEoxd5LpP3jWJiy/RjTRnpsvzVu6U9Eq0d01orM
OD3vGqYxhcOa474Jn2NUgaDsZ0SPpisO7JeJu+mhMm+03Z+rcTdJnSCYgIircm3X
DTcHeMAhnsp67g9Sojlgm83Y1vZDSgbvTf+rgl8wlSFbaVbrfz7Zz2l5jU2+0myb
SI6X1SV+i/ioYzDG5VH3giKIWmMBRWgCWkYel51PdZzD5+GtWySkFCkvBnvhm+6S
TNOeB8zy14zcquQ6j5IAaOHEbyLPrVVL7qSv33B5sIrjJBPdDJR8rqGJuWAiel2h
1QG3fnj1wFrJiepOsgRQGDyUEi9hnuz1HSD8U9OaN+NGjAWylbtoGySmpyYcfnqr
qmPDXk2aloXKFTxb3xkQiFp/4jPE+bg5l3MRecTjUo9ExKhpDNkPplByTrrEDDSB
O8/EbC13G5VNn7MlGmN0Pw08GtwrC6pdZ0HI9y/xpW1zPM4fBp9QVhPr6Yf6tWfK
wAAiZxEj04xm37MEVFHiF5RBvhsQAFf4Y5b2YQ9ZApikBPx42P0bcicZ41YAIt+5
yPtBykQeKHNQg8PxDYLksnd3eAZqJlYNm7SUHMkFEEq9LvhPgovPZcu74Z4KgfA9
Tj7U/8/6TovXfCWZfo/cM+F+RsJ0x//qlXeGsfFJjfeo3pVlQ2x/FS2NDcbENZ98
j20vFIXALQ4Fxmk3cQWj7BFT30tK/xUqUXQ9W2nzv01LFROI3tJ7IvjCM1NjVz6S
0X2Ojg4lixf3oWnW6yxeVr8GYM0mi4fR7Bnt1lhbR2sWNI88DQJm+kGSi85ybabc
zBbUhORU1ZvOljikIE0mP54ItjbPMfRpBsUevdZI0b1vJh13vwR2ojJ0uoGN91bL
2P8io5b72OkLsEPA6cNnkgdZvfkiEA6lIjEd2znIYRuoDJlY7eZihJpjXboZmZVA
rAuTNX5rF8MWtVLz0Ctm2wYzyZO8KdtOMaKRLOOo/5Vfdv8JtQQ9iGh0Y2Ejul1s
MUK8l29NdKNKV4WGwiHPzgTb7USwurWqz2h6Gi42p3EFx63IG2iFByx4SPEKBFdp
ePu7Kud4if22wjmNzkG7RfctPGUeDzBmTjvqy5J0qmrfK9avuPt3Nqobk9lDelax
acl1kUNJZTAlF9DFlOL4UEobkK7cQNxvzmaojrjgzJP3N2p7TY30h3EVYKyYdvAs
D1ZgJFNhCTfGBe3sLhzdel9Ov2f6fzRy3Sd/4EP4qnwNUObmvqv76uuyHSbNyycH
ts7pzfZfRCwZ8nBq18muePq1mSZS4d9W3VKxgExiMe/gUuyUYEb2yYZ/bOGr6oJu
cMfN2IwCSdEHQop/SX4q492W6JGO7n2wxhfr6UTrgwLkr+OGg7oUimiwVZ6CdLRp
i7eNV+xjOOhdHTR/uOsY7PjIc2fFXABBB4E/2MJWSPklTYsch7SRL9f67wvrKl8c
S9//7XwqwjezXUB8oRq3rpcJRlo7SXXdnDsyIqVffogrTzp5FypUTQl1qj1t8HSn
PGOC3kY1YjIaoSEe7x4J3BngA/0d3XyQMyey1a6c5EMjMK04qi3IWfBHhWE5VPdF
CwGFp8kqgvKRAAmcrF2ra6V4nutN+luk16U068ex+29yD5AVw3dMBBXiZOkFx11H
aWH5PDdv0gEvwo1CSlWS/mHASivtQcisrGrB8UTwJT7g+ePazkderJ98mdVbnuKG
YfmpCf51FeVDU0p54TfnyTDjq2VgVGhTJ1i/fjT2Koezvsr2aCQ5cyMstGhe+QZp
UrSKm3+O9HBnrZbDMOiqEqQmrkbFh8wMbLXIf7QDkLDLHdAdWQK4CDt0A3wbTGmv
M8c4MOYg1NKOwIm9xnHGUXPVLMaiGqNKBaSPxs3S3w4sRL5G+oQTekB2Ah5EbsbJ
SFFhqwB6AAr1AxYjWzfI0pq5DFfyE9YQ1zBB530DtpDANvUIqs0WE+owXSSVPHnu
dvZnXdzPuh9a9sIi/fb1wGDiEiG6yXMZyL/pReZUGkY+286McO/R+qfPqI+wM1Io
RR8W2MbUL36NuLKaH4Bt5uk0hpvaJGurJ6luqHVpDs4QvCPBkl+HIFLb5CmuVWDT
o6CodzduonAsNMhkqBpzpJg1AeCZyAgFYK0JMkOhsILwvbMzQccKSmjeJSnKY+I/
q4uuYdMGXtmeb8EaF1BI1yC1jCeUzaocpy+T0tZZKJaIb7dVGChexu/ERonsLMtx
VMTCEqUF83QXXehvMy/16dIYxbVntl9rDAFe9E9h/ERh3xRXg/Rk15wwdYpaliwm
nLQpC3DsLPxg/xKwa6IbiFd5bN4rhgWEOu0VBHo4YNyjRsNy3X2nBHvzmaw9dWz5
+F6wDcawpORS+hH5VnrxxnhE8jbjnB4WngTYSPcSLffZv+JdOCg491AQag/i5jca
qw54hCywURZg/cmZDZgxtx83IeEaGvJT03hVpsTjlVsBxqoY2jtdkugYWImhftOA
fgS4L4scYsVqDOvJ8aAFvcCNFThoBwSuPccqLmEkTJhZD2rOPRvgRhRsvsQkeSWK
t3i6x3cenvw/xVEwGXMn95/9HJZD/j2q2dpH572SCUKIQfhv+ZNnfu7uqM1DhiW1
85ogoMI8F0iFumhXGZj9kz4iUQEF0l0XOlukEOcIsMgSOQXSvN2xC0fuQddcL5Qn
9hvor1qMm54gvk6WoeSE/EeRLcWHNZ3k8GcZTcX1E0D7t6a4Z/lpEDtuM5vIq2Xo
tko8PHnxkz07reOktQy5FwWWOjO8HoXOt8vzePwVCtz7PMHbFtOXsnEo70MtiIB1
fNdrInUimPDpeoumXUJxPAwv9muuouqdTKS3eVaLioK1JeRuzWbcu5p/qTEfRqBa
r9h/rj26YhlHsr2ld0lhOG5JtzKPRYVO1dw/v6ES9HTEPUCLvhZi2WUuHOdbnug0
rlqsHAGMW1mK9BBBzOkWo32m5aKqCK/CLzDq/8iBN6xBnBrXmpVe96dqqONGDNah
t+c38oGw2en7afNRbDkJynHKqAtZDPLM8QZuybFkzLSA5np2l198u7Sson3b1ZSL
MZvBsoFd4ZRJT9Q2VWW8SAKx8OiiI2ybGive4Pv5iyWZnS04bWWyOdoB4FlY0g6i
zHYarq5sE5ECv84Y0wzELbPEMDvfyYotnlOdPfc8Dd6Bcz836tuS5LxhBgi5nCmm
hm0o7ZVQyhbUKtTIxfGYtC0Y+PXdOeVteWSk2PXQHHREweKoUY/G0NnC92Dy7dBl
Tl7qA2pfbC9jOd4zMnI6nPRkeJBD1I8cqipI/CfLBCAuye5R2SQwjZ7uJsjId/5l
capBha/GXv0BVbl25q20x8RplHHOEoiZqlVJJcOEdQ4XD/or4rLj41fgeCGec6jG
yV7aKdvn6UPHbYKdIXg3zWA0AMzaQ2ZfUOuVmRNKNnt65zOlaCBHkSJcs2Yo51Q3
8H4IM7eTfS+m34L6gtfd/RfRo76+9r5K3FXWZAhAdihCENwQm45uMSAEh86Z1PFc
wZiKrhL17FQd+IL7jQL/CE2HPr1b29oTPtL8ATUYGHaq4fH91HZLj7cOfrfvQL7V
oFAGuEhiFH9r/JwvM4Ewc4CVhLZrQHvgPeOyRJxG0CmYzsy+bNfZBT+91nE+OlJS
tBkP4qu/FN60x8sOeyKo3H8YdFSHxPpLluBxgQdUAUvlmwM4NvYxsjV/Jm0Ia+pS
cuGkdBGWX/VPAR0pM84UluHGiqoJzVcVVMpIquni9Wb+PP09TqTCUxmCGudBLgJS
WG/++mGuZkqdImnGXy82xMy9bvP1Ffh4XC+ekibHxg2qJtj4ua3mjVZc5uMHw8Kw
C3Nuv78SKjDe0tZ6kn8KMforQMIJXkiel9IgXc4tMCGBNeAs1vn6JtyTP0YDwGN5
x0ktoz9sGwkwAu8IdS0m9xKJQExPZI3F/Do0kOKpT/DFJgYspV8giwR2G1DGyx80
ywwmHIm+qLmnv49JK1/8VRcCQgqGAq4NLcVbZ3IkjYU+znTLKerdkGc7XFUd/5Pw
Iq3ku3bt8WNUlwMcMHylW/KLus7K2Phg8yffGQCeSSEQPOITQF+qqjCYlIUlpwR1
fo7F8OcH0gvmLfY5Py/O2BTydeyyl5gaol57zdJlDp6k9LoYrLQMCT2Ra+pcl7ex
FvAeFUSQrOqtIiKH7w8N2TKjSa5xjadF5wxmGXSmsIwmitdFBvvMGcWg639P4MFJ
BVLT7VR3cg4SZYZ7+pRnzV2+CrHjUId3bim79NbUOWLNe4wN2iJYEONAcjoTzhpe
LiyTXcRZwgFmsUrKSaJrEyvjJQpuX+pMYVhr0dSpzng/SLX5/VGDiZK6DgIu0S/E
BgxT5mefbp4cexI5U6TtIun07+IBaWO/xEi5gj47dz6aaHbM5NV9hd5/u7ZGX04G
pL1F/p1YyxLByxCHhb1A3/2upyU8jdpNmujRliZdFzYFkJwFbNCcIG+PedpyFMCE
KGyzPLRAe82pvFFIz8l07Jml7Ol2IUpSAw8YxXmZM+h3xQ1UTZspue2t2MHMJBMX
t37chGA9p9Yo42yDinuLbpRaqFs20knmuhFdDSM8IuIVSYiTMWLqIXAKtGa/3Rya
rWMA8JT2SCQVBi5tia1HTC8w12SHagA+LFE4ikrhGqTeyDXjDxYs5RrWcudJ8ODq
6RKBENcnO6Pmib3NXKP6oog3SnmrvRfU7Ukqe3ICNSEhjdygEyPEVYCY40/6ONoC
zECtcDWJi+62iNduZ3VOFCyZSGUvgFzoLlHHttUGqCu62O4fMD763j0OTYVq6hea
IT8AJirWv6B3HXf2XUm5t9IR0/+tNnqGxvYv4XRaP0E+lUKh+2NXWTTFEwNSugCP
vZsSBSgiFEYEA29dzcp37yEyniVJr7WLqFpUozbOMsn+L+53zV3Wu5AjlUUTrPQz
9Z4/kQrPJTzMCoCx04/29WkpWFYWUJwTjdEAJlRanxbbqx7qiRPJPSAosyc1aQzC
jr5r2OMRotbiS5yL9XP/Vb0Z4UCwcMGrCqnJIjr/Z6FFyc53LUn/sd3z85k0gWUG
FT+peRGhT57+1At8mqbLk35dTlf8jfjKuGsqLsF7daAw4xG4An7FR0sweBgYIIvx
Ma10VFDWCCxGOddsdUa8zWwiqv6qXBDjrQSZVjt2yQ9Wh4z4rUKIh8jdfyPVRoB0
/Wn6bSaZ3nZlxX5ZgU6310LQIKeiY9bmYPaKSKWGcf2LdWfVuH+DvEj8JMP3eljh
NegNyBpTLK29CPtg4FJ24XHgm7gs/PlCUVFIouQ/8ztHb3cUGkCiYbUIww9rgfk3
hEf460g9fw3A5IhibXZ3Kka42+f1XwZ0XFoTV2QRvLWRNpkydvpyoWreo02w8Hjt
mzeicyK6snaW5lsoGUEkRr+qwFqpbOHF3JgHqbdh94xF7WaD9//nC5IRVKtk1Spg
Ygt8s4wN5fITz1sOsZeGhbePm3pQOGHt6YqCYGGRVrKnk07vQEqJJZ41S2qKwTje
hgcMbj/YJANN77U20b5KIt438ZHOav3dPIbUfip6jnXZwYi0B+wKcupo/rR0L+fo
mt8gkhjQV6SXmFpWLD6otGWwlR/nkaRq34sqVvbplWBuKyCEzSgwDa53uCXdZw2s
EN2mgqkSTKD+bM3CdrXLIHLOe76FOw9iXOFxhLr8b66gPBRnmaoxhiFqx5erMto8
2XzhcKTEIkIutsOfnFocy3zwxAQdZ7xHfMS108LdhXHPpsrqdVanhLCUsJ2a+EVL
ZqXdj27PNIPDJLgTp4kbzyUcCGafSvCWvCgQ2iHE7fWkcfpNS5NyQxe9ZS8yN4iL
vuKd0GM/0OmKSiXexF/aIzyYqW8KjjCNpbMni8CcLanYbmoUAFCClBe4Uq/C/XGN
/MhHZKyZTW6IGSKMT9E3qFC5x063v/m4dDxTFaqO/6G5vGOvmvdcV1WfuYjk5Ahx
gMN08WT+i8LclvIfSwWQ+D40CWULe6iaZqFZYGy6kjsprEunjUYVA1KbLeumNJwX
KBtCC+W2hJN7pqVTC3p3KFN6j3wlgUIZ4PaCk4q6j3RHeYPKi0KOMk2LEYX2bmPC
9DozZEGwrDO7s4vgnD4dNYo4cGFOiuRm5545v6UPYaY3RL0nh6jKpb/bmQKOLWEV
mzWEdUHTwWZZ8/HgQeDfbE3zMXMcQd+uQZxZHZ2YpyfaiT7BSxOWvLMuNr3Q52B+
2+56r8/Bq+L2hpsyQ28R/k5VTSPPuMyByioEQ9/HXJczXu/JMyWCCCS3dDHriqrV
rDzHU7ySOos7V9JFjVz2vS8yI7dWs5cpGEzCEdBi4JndnOGY4XrsSyjsP3zaC0b5
3irbN2P/cO2tbVEliSYauWF9Ui/O7H7qK88pRUfr67anvKAKqPBVhekJnnagGKhN
yPeLNOUrasxXwJDEm/yccFI1nzGg2ug2MTQgA0Z+1Qu2WFznUh+y15kAtkyNBLj+
KrrfUE3jj7qVw5/FcfQvBPT/Knlu7kGuJChteUOHHdc19IK83XEsbOjRXO58jPQs
yq7OdjoyNtgriXQkN5vE76fBeNzScFZIJOiKRryEiZuOVmWB2AkWBPVjxrwhoXQU
dgFHxRYHNlghgE3ctPAK9+ZMGfvFajNkyB54EOZAp6wGb/uShq5Q5+CmR8IZgU6T
fKZj/8OKZ4r/BwesQNixQXUtTSBnHnbCg8FglTeksNajH5NVcEp2ibt/jh8itbbO
AXxB3cei8N6cEFllBKJVyvAukD2Pe2HhKcHSqyh8n+xbDjhv4HgzvHYXBVCePhAF
wltEcmp/trfj0ID4yzkHt209jDaQod6NL9IQVWBCkRlgn0zJbgnIEzsvCaReN1qF
2TWFbF0s0/1u2shf2z4DBXyNNy4LLCIfaKkV7rMBcjygse9ATlL7yc2TBziG0Wok
KC5aid5NbGI/rSuxQBctX//Wd6wLcDplD8MH1l60HNO1EwxJmyk1nGZiioSPQ0gU
PwGQITfknIY5MDvKij3LmdmxV9gJlDiTHGcl+IoFjjhQK77YwVWmSI9iTgA64/+W
scFwSSiWYhW63avz3oT2k/wHNl+8fgUG1LSajtWjh2vhKlf38kcGqYW+5OCvulrU
YgHVUJ8lP8BkITRTiff/S+fxC6lckvYcqlcf2qvg88hn9IO7tNEFmuwMs19PyODo
TviA7Y9jseVteRc07lJFLLJphUT5UY0Bjnx1VhUhnIPaUpCay3Z6TvWPagBfHJro
MjXjvecQ0Cn/uqCyRZom+66vXdMdckkJydZxQjP6icOJs3aqRy6ouwxZmijQnhrB
dd4h0fzHg6IaJiDHEtWf63ArtX2fBEuG9m1lgCjmi8xOIUqnB+bMp2h3Os112L3B
EppbnPWEaB7ptZ/hLOCdKwBCQzxOr2XBY7lVpxWPMowi3b3V5Q7jEEHk6xw7LRUn
A2XKnwovzM+yOna9VsuOd24DRvulsm0own7YKEpkjEHZejF+1tekjJx1QsZKZZBD
4v4Jii5vuPEeZDdB/VSG24OxMS+VEXaEDm4GSDe0BrhtNV7CfjZTyf58UBxxYasZ
ouiNGEBC3OUPONb5LAf02YWoL6gwWt9LTqAP8Jm1qy1DPHPNn1yzgWHyumTVpdxJ
j35P/9nL2uiP/sf+3m7ePiqD3NVoPfNRslEDm8Gu/wDcwxbM/dFZ5+UOoI48YDCH
tbKE5hHbBBea6GTc8X94BWFBGrHgHTjcFGScOv3cO03zqIZgkws4odf6cYX1922x
LJrRiJAkylYRI5nhlWcMvxM4rpsZXADHdS6s87wy9VEbGcAC27/gqW7IWU5PYJ/d
ECS7PlADdROTTKQdcHgNWFFEpcSE8BudA4HYWXJoqf5eby3NyOG7dvAbSnM5EBsj
Q2NAUycen9r1GJm+KGCWVASG/mNEcsnsRaPW3fDZehTlOtTCk7Dv1hGcfs5ZRkhx
fT9df+V2pL69wRLaSM7PT03S1CeGE/w4mYctckV+LtzYfM64BewjvyGP9EFRMZzI
QeYGfs+6xj7acabB7Byskp4fqAC75akpv+Vzq1YNsPMO843kSr+lU2tZJ+KHJy6j
iaRLLSYy2eHxSoHOCEIfrTa6f0JqsqKu8G4ktOQgyKZbkNNN2eODfXazebqEgOqt
smQBGh8cKJkz8O5ZHpqPQJYbGe8F83U5CZ2dVsHzI968NtZg3RIoaGPm0dKXTEDe
rqdhvgpB/GJxUwolhOTQI5y8iGV7/E8ocQg+zcd6Dk3w4tJHF76wCxI7CLpDtBOj
r+zAt8+YOQvEgrOi+mFI912OSGpF83FfU+6O8yHimF/i3nsB2C51tPE5jezH7hBa
RMtEvKVeLuYqqkduKekWzUDZFxGMakgI+NntXQ6B9lqx4jgC2ptHVjbiUCppvGAR
mmYduRvq9W7iQ1yYWVVtXDKDD1IDa1p0tErPaDOmvXl/8EcJOS38jK5JgMgnFQJ4
XeUzf6+nHjtmz406WspAPJqp05qd8UMgPcRHW5fY7C29yOirYpEGz9VHBHfGTxki
JBmauDMULi3wKau5fD+TgsElqcFYA4bnt/yPzQupHkWA3XfTN7IYMKgpUwObiFBJ
9jR62R5UF6MKvlyc9C76uGPTZeKYJANuUEQNcyw7pOV2nPMUvLaMT2n3pTx0AXLC
0/8gLYfBvGW/0fkUpTWSeVuOyN+CykJjatueCacwEDeub+m8TXg898kb9/J2+hmi
sRPRsCUYQ752KINep5EFax6WpfvR77BQXl5LoGFvE0QkYaSgQTXYhUOtNY4JuG/T
QgVb8/M6bO5bWYTfrLNVYkTTQd5Dbnra3cFonnN4KUSUDOID34ritYtM6VarI6MQ
eNicvun8ed8W+0Z13Aus3F6jxjMrnBox9OE/b5OVr1TKtGXskIIuq69Pp5SkBfbZ
HJyeJ3h8TB7nToGeF7WfdDC9bFMNwmiWeF56OYO5BkzvAP8NJnBgM94F9VKxRbX6
MNxeRxVwT2DiNNQMo5uEjJBN8K6sT/RJynGBLGWIs63Ky5JNFk2zXWChFpiler24
a+FNHBZHtaLTrFseUgF5Hsl0o+AijcW30EwyNAMNs4MrYPiXtyAzONSAsURufiHB
8Dj4iFxOyVmixe7tpGdcyVKIVTg1fVhnioTree5bYBbsp3Ohl5lYKSmO6TmifmzF
8JBt3gJRtCZED6al3nwTs7LKLbV6r62oyEWtpReremRfZcVRDFbBOdNXP1oa4ZVq
wo1g8yFxt/CaEsIHVp/8mETC5Rk7XVCteER6T9UmNcLHAh71t4ieH/5MUhWmBL1f
drM2XCLQ9byPqCOVQwRnhfuwF6r44qhjy/kL4BuPOiPQfiqVnKDgE57jSFwcmsg8
ULZrswb2RnVgj0mcHJjkmn4mHvI0mRBpty8783FrvJEgjkDFqdc1SJvQc9/C62CL
UnjYBFvYY8tJ8Z4QmOketv03d4y0TxI9Wj9ScSPEhNm0SLe+ysZ+oMZ+kbuCKVy3
aKs/XH6AMybiL7cs3XJxYv1tYTip7EnpMyGzyAHcsZcrhwq2nfa6nb6KgWtCTGAZ
0ZuLiZMVQbjMdhicW50WpD82fJAP9M7h3nytQPpHKqYKqBxWJHrZWBFGmYs4DHx8
qCOeh4Cm3+JV473uTNqFh5x3dRK/Nfbe1qXMz2tctNxbbekgABIXTzcasKeERQ/V
ct8RTx59el/Y4cGpp/39EnVHiEnd5JnuqmMG86MyHZY90MyFxbhM971/c1HTe84N
UtDZ7T9z4LjOUIdMrpnavqgEY3T3KyLcYstztCA500aYhDWECyL+DpENkvzxSv8f
AzBA5iT2tj4arty6JDkgk8csKzDjYIPVI8aGkDm8QNfYR6yUOxAro75EA0mGXPvC
FQLCkvPUb9rp/4MSsIjMvQsgghz3l9EKuV3nfA4AOkeZusvHboRethXhQtLNLYVr
jbhxIhw4+RRubhlY4a+XrR8ewkWnNktzFnhTsmxv2PND/ATJFQsN3KompTPijhyN
g6XzlOeXFrUYvLyOaLPTqmPaO/Ufy+hc97rZDoughxRCqC9xJiaOgPcg+dg3iVaS
9p4umJvTgbEC09cOTQDgttWjFzY2EkoMR+m6Y5x4uOgStM6IbcU7F/tszChj22Rq
CCxtx+OTg06huxYC/Xdulhjul2gEpexg5cC2hOJiZMUSSiJ4jHbAt0qUMZoTdrpX
kskIVdfWupFN5z7R1tbxnZaF0lqKn8j1AG6fBNYt3H0s7xUzo9Wc6764VEbsPBll
xp0/kvyynhQCrzPxh0qbxOZ5w/IgL/XlFHoV3Tg91agszYYjQMxGKkcOYbAEz/MP
yVqDaFoMCHyTyw8XGNw47TnTaXXg6Mg0IDx3UcASMY81U86BmY0JbUf2EBljQXJQ
2rxvQt8rS/L6B1HibjnSzhsMA1tcPjMMTz/DIe0KiYbBz9O2i0fsTZ/XjOmhsWhc
HFIfqK7n3xEBrBFppMfsS+0TlGIltwpZAurxuAeDbwzPEhBXShBYBNcDqHZ8hje8
emhAQqMayVSlwSHIzZi9Y8hdwQZeVW6U9AQbbbIuDEBEfOH33i0iDSMG2Mpu3CjQ
C8GtqyJ0Xt3cP1uM3UDwdBy8kocAgMLXWIjz1ATL8RJXP7FkN0yPARPUS0sA4srz
kAH63m7OkmRyWbIhxbZQ7+rfJ6dp0hGkKwlqYhFil10bjfWS5NsuAoV084Umjxji
1U35DY/AO6qUxW4NB4Z55ufkvuzrGuuYDS12kFejXFrd/vE3yAmXTZaCrwr/d6Ib
asd8GtSk+vxaKkYhRmQ68wCoJ4Gmt/oZDE4R+YA+mapOhULyymt1zKlclf3De6rH
IcAtJyxHpG7/HnFCC8bBVg2hMBJKYkBddYXIxDCWHv4/Oyrdua6JOcyAH9wiqdA/
7Bcnrrfh6NyHa7fABK0/iEnOBCPY/E1xETkxFfkTX38LBB5qXzO9k+Nib4h6XBII
PwB3uAOSjgnXXAHXsY+cfyWw9qW5XehgfTNJWMnEP4v9ZzZzlz4YPD52iS5AO6RV
/pSsHd2C7JXY3osEjxNcHDFMEQGv6ty1eXrQOq48S7ZDZNaov0Urg+d/pyOLOTOJ
8PX3jRSR9UbsggY4D6pNGT8OSvcde80V82xzD4uKEtoY2iNBzRcKwrMIGWb2RSD/
T+v7eYITFPWB8FuRj/3gbAFVinslsa3VRHSlzLCaK5FigLe0k9D2rxxKbJH/Zjfq
sTt4eLMNxUNN5DHVB5tDGgwT8JAEZFweSfWfHx6sjmfvYw6rrykUdmook684Vbwk
lT6lQ0A2CpiKPoerXB985P+T6DL9dM0kxrnunKuqjRjSDLmv+ufT4cgYBbm8LRet
bV/UAa4LFBaMe69KmM/LIhDAwRqtWtkolLADxWZf3sJ2FSRHngicPCdueqV5WpV6
Iz0cjpc3XhInreDBBeRUvSLhCv6lKz9wIMl7w6W4ktlFk6XqQpgT5YV2X1FEY1Qj
0sGGhC7yng1P1dZ/89ZGuZGhHk+QYMSEHQspyEQ3LhTu2pB34Lg+t3xpE0qUuCTP
C3KrlSStpyTQ+1HOywQWwHOlPNFGul/ezIsi+zaPOHRg7eOk4hoolB0Ja54A51A2
QuTiZvlf/fDzA6Z3655vhubUZECpPrYz99zDs9JZA9YZJHjEiST2wis/wXQB14NN
/Jl0SgHGmGuIkLyq4FiSH1Ki89EJJbyR63fEwfY3ExsnigsSuHs/cgpSVF3ipOUD
2OsEOkhatfeQ+sBfos6WYblEJk+NCET0Rv+RS93BAEiGoPLp632YV1PVpmT7Th6S
zOvzTDByisxAruTQWwToDW7HeEK9P6wTcLk7PvZ+RA7H2RFsI1leeCEuRS4hLTlH
J+ycvIBptkctr4i0HViCDJlI/Xz1bgD3Dn+lH/c6vrYY5FgDEtXvcesE7QB6ziEr
Ft/uG8gZtPvH0UfV5FOoUvuCHKJKl2Dr+Iw5IYly1l7Kn+3ZVRcTT2O9Q+igJxO9
PfF+9k4OJUi6cugqS8FA8ec/og585B0bkuq1Rz3wNEyrUnrwkmg6iD2CdvMLRkDn
y4g8B1ZQfT4x3PU+EsWIaC5kRt0Z512EmraqA0WyRbK7I3RvRTvhAgOpmif+O0od
mAqgDsYdfQZf2pA7+BfEpEX6qc2BSWq6aNjJX10fe+wlmlnPvNz5tREibiAM6Yq3
ETh6L7mY+2y9MNUVPcna1RcPztjVW0knYtTaeKvRksaiOrwTk/jvayAig0hzywEe
tFfXOAkiY3TLCWUlNlI2xBzfBmAyYl3t/Hqc4YfhmxfgXn9dZnNea7Eg8gLnB017
yt62Lxo1likDmY1+V1V6OuqVvlfYsc/6qQbs976fEn+SY8bSBvtvezJvo2E30FVs
0wbQ3y0ILZv5zxSdKFarAZpT+RT9FZ2+EhQPznhXdcsM6Ey7W28N+9g2ymLWqr1B
r4DWduC86w7t4jhfUQbGPybRPmFTDajeP0EAbs9MuEfgMtW3jT3elFMlN7wpYWzu
5sKuAWAfkyR77cWM3MkJ8ANCTqUDibUNE9qdK9vOt7O6TEPx0+ixaShL8VOFeGZe
vkTPvJOOvnCDGEijwi3MPPtuJz2zIl/NawZ2YRvREHYmZowoHHrb2QUfmgfKqEgG
x0sd42hug0Hj7Qzf1B7FHYKwrJJPuAeWCzGU+gdWwVU0pbs+dYsolGVmuLABRyqF
Q0Ul/IlqhZo2YjdFfYleTdO5Z1006NbJfcaytjY7iodTHQ0Bj95sA3Gd0kOkjSbs
Sss88gL9PGGoxzsDavyPv1MPtnqTqmQCgQlU9G4cyIh/ZtpgU3N4FrHmy/q6Y3fk
9jeZeslOgr6MI/IgB5q73zxUtJ9LG7AqxY23giypIfW4NtHH8oQJ1RP5ZWEd75V2
pD93EDHC2GNLUgIamqO8mgeVxpI8ZWJfVesdWp9X/DlDqTfep+AghXzKZYmeqPrh
FOqqZM5jckI9YH03uX754Y76+kXvl65Yxk5BFGxeDl4OU0eFaROkinajC5ihn4Ef
0cr7ibIuMscIuIR3Mt0uecmIen9cVewFrfcevNB4F8Wot9KfPdvSff01pHdDi8jj
3duwspcvZae7i8CYatP8ciHpryGtK/DLZDMc6JW/ykrluH0l6uLmx1W+GkmsozNh
TYtpKRzpV5UoqssB4uN8v6xGpLM/mJzCl3KwE6t/v6arn7Trcn2wvjTlITpkTQmp
g3ck099oR+vXg1q3Tzh4ZP77hf+qxh1rxYxWyI/qiuJNhMrOohpShrvr38HUrjM8
5SlRE3fVDk7Eodxz8XiRAkifwCOISi3VWiVhzjLwlYnfkBY9SSAy2WgmbK1g73zl
r5rW5Kk+vXnvTpvf/76c82jaHiFKaRSrT8OO9aXjq9kwb1/9wOv7/AUbwFnUQUlv
v4QRB2tTSWMvGKZyrM/e0mjc1qjTQk0fT39MWmA3/X52YkihVd90XN5IiUjWpj59
jqOiM9oJCp/X56FHZVsrg34R/NS/ozNQteabP2Ocq8ulP+dHtB5moBEEm3SIgC1q
+DK1Bf1q9SEMO34O2Q/wHsQUsXIimPicrDpqwrHDkDmaf2AArru4GMLK0kqpqKR7
syDKdHhy//iwNbwlJxwFb+Ab68Uq3SLmS9h6a+YDnPdn7ASCPMO5XJxd9XHD3ZPm
o4LhBdXcomoFuZora2YL3KLXEIkWzoNYhmvOb7z20C/M3vapOQTMq1RvmjIYUJAg
WBLW+NjU57cmVlnDr7SswnRNqzf5GFNNC1HelrXNBv6UID5V0VOYeSfW9BLI0PKu
Q/sSoST7kYX2RiIBKsx8jIQrHl6WvZOv6oriJcmvGO6X7uftTZPy6FKAGtY9sTG9
hFB1BAaiOsdx8QO0EKVet7Kntho+i8Ws4SzejQl8crMwoa4VKabThgtJPrn7z+uh
9AQlvl7iSzQH25t+5TAXrGi2xispOASMySXPdDAnPLZMMO0HhLe3Yu6FrnuRQK33
+7u7aW7DTs2emxOZfZtka3iOGlcnKhSbheS6TvNBJ9H9AKhR8Q32LqEu/CbwuC8w
mofgUbUXQLVk0V1sPbEhO/8oWqsEJhEUqiud1H3fXJJhkczh5sb2auxGu56+ptEA
l6VoqyExmaRvnzBYTP+TlyTExHQEghAQRyhjdjYth8mIY2aJe0jpKjPQGiFReHn2
dhOmIwqSDA5k0v138WwYRyzw4AaZSJkTQhF8/WKsiTFV4AORifJUfROGjNC5PdFX
LVVwDW/yoe3f5S9+gIUFYeu+dEDaNiEh2fXjBu++vy7nQ6Vt/8o/S0PgpLbY4WM8
3l+bbghQKY0LUlX1F7vZ2zB2qk6e6ueNMpC37CnohL44qKjX0Vg0JOycloDh/DHd
5s9v26fBupenkHh0B1AKbp4NtsIYGWCaAhNsuGPSERmDXA0djKutPhD96FUdWf7/
PjvmvgsGx8ELXtYe3qEHbuQZ1Oj/Tq10OgY3aqHJxeiEMpyY3g7xLEpEfWw0RW7c
ZV6zRLFd2mno7PntmZqyVxnVMDNty2Z7IquRZxkH7zUKaD+Iq1TqLnl7kESkoY8I
AFihoSGK2BgG37lhtRSc6Glikw3qapjTWfx52Aqc8gJL2XlchcsrQnH6pyYDF6IN
NQ3DgYqGfpkoqxLzhkB8C4T2E0JiQI09SpViPIbjuuzW5ZIEqPGgfkbFhK+/Y4uN
vkCIfHYJaZVTN6ZDXzxLe3GE9VAIvhLQNn3up+NhzrVQsPQUhCmX4KC4QlONR5Jp
5FzYviwrfo1rabuh6ETx44cizeGEOc3jkWYfQmHysXsEU+l4hE91Aux2KkSTdvol
DBOhHTE6hohp30ePbITtwD/NTJ9jRE5Rtc5Tb27BMGvdGrFHUsmedjRucW0xQFLE
IJVI/JIW2OYf8nzD0mLhGiDmnT5bS96fmTLiExrwIi0uxt0W9WnSi823CNLel5oc
65CGHza0ahPOWt14b+Ujj2AGKJLcLdI8w8QZk3U9lBEbVolkCTpfxTZKNuOHM3F/
aqeg9/O4fWQ4X9vjVlVlQ3hC+AQV65bHCAddJQ19UtcrXh2dBOvwmlGJ/tub5UaB
ACORkKu7q7rx5ORBSe2BtmOIOzP1Yaj34wLHCTBF/KAuLgfAhXUpbtRs+AfpS5tR
KsI09o7W462COueMmejzQHI/aenE7YtBLlmolHi9zhRn0acwb2KY08Xpw2X9I5lw
QSYhug8BLVo3sElg0Hb7CDHZvCjG9Kdbf3WN4a6Eksz0GI/XSxGp8PDjqAeOOWVe
PFkUpyosXs7QPLul4DIj9sj7SraxEptAtzsNW/x5y/yL0+3jF43cxCMyipvUKr1Z
LIcBWqdekt7PJfW8gq47TJ/AqxVE+5V5Xg3kDTEHUQdeHHlDAYL22+lY7gF0+QK9
/MgH08Mk5RvMDSnO7pZIClXOGBEGN9ZQrtgQ2uNo6xtu+ht/Dwj+NTDAv0xecntd
aAVRQOZYiM+REVjOK4TBcOb+jZ6vUVbGU45qlR+wycfbHjGdgAawl7ATxQ3szQhk
ikMWflH6ve3r+WfCJeL1VG/7pJhhn6saazty6KxiMr1Y01Wyz5l+KHB7oCmdZYAu
FDluixboWO+lfjm+Qc9SpFQjFhWRjeNB+QHmKJKb2IqnMJeS3QcKp3NySZtb8fqc
WAZHtOlmZp55csvcVAjKi+13eiq2PqYSFmNTG4oIsQKpoeZoRJ1PZNMKu/4QmrtO
EdaEcKMvrwrq7DI2FsUXbue3nFbFO9ON8q0vBeY4q/HKdW/QOObXMeBj2RTVIdNV
DTZVMIl4Fck65V6iHBVZnEmY0qI2W9ltF19GBoGT691ywFLPo0oCT5PYxa1I0yF+
c4TxhF4j9lXyJwlP1yG8WmxsyU+GOWYoa1T+admjsTcUqjmX4SpDYjETaZkFBrN9
kucTgZUwfiQvpvgO3pquC4Zuk/xq3yK7cIMvWNq2sAtrAilVdkqLMBvUx8rdOnNG
uYvI3ImADH0WXZo0kBKuR20DSeCX+WQsM7ut12S24ydhbIToGOnkEyc5MSc5QJaR
ninLbdvWqwyXdux3KqnrhfT4TQ2eC9yvH9DQ5Dl13eEr1Ln4vEIEGKKX8Q5/QatN
lFb4L3el9svqGmMEXmvmXBxOif5Lmwlax1caX6uDzJ1B7Cj4+4oMxHRYcdbLH+e8
Lr3C5refABuS9y4wlOzzNg9VS6vCqBjEd2GHbXSot0u1LBC+w0g1KYES1YrshIFN
gK2f8FGdgTMpX2XjRqHTgtPzuv9H2I5h5ao0vnowZaY3sFiLsRNSRNel69aIX8nh
YypbZ78q9s3XPYk6fodgijpa8ofvseo/84MOn34/Y/BCFbDdR9CiEqdNJJDn83QC
a40Kvz+5UpYgWQj1/ngfvkQdI/bs8wSSqHbA/28BRCAEvMWFuo6r/UwmfD8IOBv/
gvahGrdAMudnm8vVYQNq3V/qBlznA0+ZMD8djk8YEuZf70yMGQkTS13Y7XRX7YeW
+PPeYfcH76GNCVL2V54V7dxfmF3vyJE7w9+snHZkbfF9f9MrUe+WuTQm18Jxuv/+
ZrEWO7l0t6rCIOYZLssAgTe8leC98NBroijPBItycDZQMhHNGwNesS2DUSA//h1c
lavEHtvyD09FyyZz0qkR2bT6wYZ4imgFEYVN/jCZkwsgnUknYvQyhVlDqjdVTO1/
pnAZQQEMIsv1RGLlHs89Vqel7Nj4BpO8wUMGFF3JYITPxE5IDO2qcivbfI8dNAlS
YHlnrYA7m+r2TwcC8c/4/1I8shLFUmhFl5jOi9KE31j6LshVBhjpdMCJ+scPuTSv
2NNgTFUZdpoD8Zo4IjI4OMagoBxBT5cxRWSKAKq4hE0MePL8HaiWsDhlFwL4uyEw
BV7IY+vRzgTicFIwzw5Imw9rH4llMvebhsIh7HC57H91uMBaE8s/yQ97kwhMEIvz
4PrPBBOc8dfAtDPRMt4/1Nc3trcqgOMFRJv1wBjFMFJ0ahebldTAzDw8JPTvgd4Y
WUnYqRtGtuvYUMXQ6jgsmr3WQHc/NGCwwRy22FJsIcW+B6c+rDPlhMWNdreWFqYC
6pL4PhXDOXp76Jc45p7cxJ7nu9lpt5AGTLg5foOEQIruBDs8fYI5D+HmwKIT6LcQ
EecYIDO3ZdPsXuOzuQWfqaVrdkV/zOnr3MYxLzWoYEpUzsZZqg6jwGuVsbxVyVPs
WzivRvSjE6+vzdNqm+iFqrodsNwKxpuVCBq8E9+whubCc5kE2PO6KXASSvAid72B
YzIxjgNUB5OHHExFJ9pQ5IxgqIbwO9hTevtx54LqnFuKNfbS0HEyCBXF8fwAbDS+
YpB48XPmw2s6XtSkw3hh5V3Dopby+DlYwp+BFsnaPmDkoZIhEselwWjq8RxvjKw1
Zn1bLcas5FE9OUXU287fkBcGKz+QAYYGnCrNPdfpgzmIzSnG647h9aYHnMGawn4H
c7ygRDr/Cwle+pA3NdqKPu+BS+U4gmi3r4gTvSGnKQ9Id0/bPQm4YPsjJCo5YxZt
lHXcbc/Y0sHawZSfEGmD/myA5SBUMgSdxXEz4Xe7dd8Vl81kYW/E+KQ/BLydoaMX
/4v8qZ1omhKPTNVD9XeinO671qV9S4LHO12+gcvHN3oYz0jqSGqgT/dUx2NSoGfH
F64BGxdB2MqhEEGelBEbBOMC7+e7cYuPzYSddmu863qW0vndpLkdakvODlcIO2hD
SwSA5BFTNHeydG4N3pE4hbYpec+qC1lXoZYqhMfpdSRsFAMU9wCfmDDdzpKB0GYh
qJWcoxiNT/tF3697b5Nu/Avf0vXeLV3wTgSLaY9xp6R/SqBQtB5KopuxdrpZyk7c
pV0eLivTDt485RA3/QzQXoYcqaHu7c/rW+Bfu421pDqGx3aeVTIUrN+iQjO29Rae
EwOHqODVrKF42XIaOI5ZV58ggWyZck1+w/Q1ijeAtPHGhvBS00ZAmLa9i7Gi3Nt8
BO+qUzcWUHBKynfsdjuLOqQwFhEEIfkYSwf3HstRI416VhEbrjabUmNaJ1b+h7oM
2ecZ4YETDbAxaePmweZiDsdtSPL1tt1nCJkMcY9y2I7Cnp/VqmS6/nXQ4yN8zluK
qK5Z94EtuOU9IxH6B0tT8g/vUfj63kA0kgko+yYfkW0zMcZiqwJUdmJqw1HMvbud
XRcN0QpH1uZp8dPpcBBjM1UriHnFr+VD53ef+FCjpyiY/8g13xYX1FgNmsD6INDR
H6/SvwyG1lL6O+XsDQT86A9koOkMPriaWM4bMplNiWoWTdUsb0ihuuKNsGLfwAIi
NSeES4WAe5/2cP9YjMUhcM+J2KY32i3AFX5RWvFKLaNmwPnTgrKtkN0I7EFQ/Enl
j9F1Z/czPa4of4mWe/64KWH7uNE07oTNEN2R5eoaMAJ9klM7BNfWchMehKncMfov
6XJUYZ3Roi0OuEn7UcRla/RKTcUfR50sbI6/FfKctcehP8VQpckBGEnki1XfUlsK
dH4Anr9HGdgm3owKPw/SCPy/h+hhca/8JgwztGKcvkN5884aEOP8Y7t61sFGGudo
CbWFMAg9znwx0yrgb4bP+wUDD/emmNccLfqAKMP8UR62LNI1yCk3yzIcO/Tin2Nh
7dFSqPNfdf1E/Sqt1JwKlBqVPT53fjce45D8l5ZsTrKkcLv0ZjcDGH9x7965IcFV
tI0h59Zs3HrCuBW1VJBogLzzrd0EAjhO1DFLjIWiDy3MAWQ/7zdtuYfe/9blviXi
b+uxNK22IRD5A8dGuaqH5Iza4q4ntFxCnAWJKPN1EuR8Almc9jlfaAZF6c6xfEpV
qNOc+CiQCeNjrBMBBem28DP1NoyXQBDUL4dpMji1UCmal6GkLoBWL7aT3zI2qA6l
Y2kkmNeiT2v02R4KTXLACpqfH37TpLwEtCBP8yy/oac/ijK+9Uj+AmohwjXSh6zV
ridxUBtIWdJvrsvCac1sNXd4SDquUkDJlYu9L7dWYDaoyabXaQv70j5Ehwil4fvb
ViD1jMxMl0ZVReeGwwbEUGmovLMmlQNg8c+14Cou5EEE+gA1KA2PZRUeD3N08rz4
LtOhkIIpINPJ1jB4hJas5AYSIe/Irx8X9R89kqJtQxIgYgHQnCLgyz3Pbfb/FVRu
sU5UKZ4tfSOi68/wq507Jog62b5lNA68NTx2CI4Mm1NB28pHLbjtgCoJjW05VYFQ
R1HC8iAUbZlNmhGyzfVsLIL4ul+6r047TUKaUJuDS+qeK/SixOoXYB030pkgHh1d
fqu1RSvsV8e8erIDmwi01EiMyqZRxzsQq3Rk4NBw4eBNizYCDx3f1WREujTsGheZ
8Ghwg90ori0km1Y2q35RpeH4No+OueT3ZG+JxgXWBSd97Q2bRThad3Rn+IfyzuMK
21uImuzLrXGLc0Hg9JDmoSeYKRYrqGqghqHksKbbiEnyq8NUYcVoMFjurB/3WLGl
dBBcX25SgGShu/iBLpRqkd43UdPx5CKTOcnlFPHb4j4+SEvRS+vDE5UGSeqB8vO/
S8g1/Dz+zQi0bWu+zEX3y/fyMWZewZD/04kseJLQn1neeDiADBkk5rcCd3LDEMPj
nteOCaQDVKexQO1v8ofaJyBOzAHStF7eDW/pcBAPgZRfsAel22h18SBEcqlBa1Th
riEXT+jlL8d3D4ipzPMpV7bgfiq0cRw1YQnH19OtgqkPeAuNampSWDl+IuDjoFdj
yf5SF6lOgKt17cG2CWjGwIQMoYiebsE/CurSPuHkfDqHJB+uXzTzsdpaQrQP832b
WZzKlHKT7lbG7NrtWxWc99Ja//ZxxznphSXfh8dmuirBTsC0s4wQFcGxSqZAgR2c
AS7PJv2oxd3FNM4q4ciZoXJygCs7GJju+RHoI3sm8qql45W0rHcsRddnh9bzNIvm
GwXuKyrESKHCgdrhLMvYNe+cqJLaMZb5Dp3BqmweRTJjKWMtC0Jhg8aTocTYmhzQ
jbZa0gaJ/nyu1bsQq07ZqRA3m8Eq2Q+0H9DJmLoO6k3H85IiCFouqn/gMcfr7zIf
bKRukwbFxL+bEy6iEwX+7cuvxlodrw6Zp8s5SABfLXTCL8Cha5RapzvEGl7+ge+M
Csfr+QcAW2MlediIu17oROxE55qa8i8e8OKyW1mN2Sde36b3HPHDFgUHLE+pa5tY
qzlpyX6QYTa3VRZjzzqx8d35EO8mma1P25SV8Ay/nsMl6dAH8/fWI6t6QYinj8PE
G6VPPCRSBja8GQ/O4PZrpPLz14A5JBWZ2Sz2bnjS+WGskioDDMlCVD3A0NLyetbu
xRPgkqSa2R4mUpiaaTAmoYrofZxrb+ADA1mG5S7lm/5L+VESiVEn2W+/HMk+K4+T
3MZIhfW4f2hPlbRGG24ArhZNC3McpU36kFioKhSJLXGt0h2oVd9wowtNPbI2X2ML
j3Y+E0qGPj7f2qqI/zBSpu2FwWHr29O4FC9h4JdG/P43UMEnAuB49/L7WPAjarbf
oqVJT8xWmxPTCmiH05qtedFjZZ2PAsQbZzIf3CZr6Ly9hDiJQwQgJhd3tTb316+Z
48/ptF3jdQjqbtB6whQQ1/K+sOxgkab8fg/TpK0LkwdLGhzG1uDhojGpcv4+GNb+
SO2YaRZiYvXqnNWwItJjiLJHKfu2hP0k4e0zvAx7vBOxh/yOv0kAYGAr7/ZOboXa
0bYRV/jS13bWQkMnVRsNPf+FCx2GC2CF0N8KfoliAx4yosI92lE6tkPRBZLtA+0K
1ZLng5uAMboTOKhcWYzRDyHL8IZxctzQviy+qxpMFoh9cIziMsLvC8DPstcHAc16
9NvHSsYYJlFFZuFIvx5Ue+cet2XhQvz2gNSfUZBULm6h1padk1vHtdg9asCiqPLd
9wZH/MVJVA1rXtlhy/RsNY7dqGfMhqZ4q0BqglYy6SGIbgc84LR0kzfXKmBHk0Zg
yP6UOXejEhRp/ZfNXO1z+v5KmUNh6NaM+21M9dGSSvLu0Mv5WMcYeJeKRLCX/8O/
wCftTttXylRcYa0C8V2fXcpOgI0Y/D1j5geCYnYayanrsrkWWzPjIQmQ5szic9rR
p928NIS+JqU7tl+yZt617+1bNKhYFWxyv0QRUV1Z/DsGl8dbLcL8sU7jineF5Ors
MJj8KD8W0L4f9LkGBPWAs28UFNcVA9bQPZs1OhfA/im9keOpPX+rYbU6TjS8aHuv
aXbub1+o8XP0qxUeJ0bApCH99cYeLLF3kbAWJLTuiKtE1cqW7EcmWKKh+bBR9lPB
+V8RR8Usc8Ai6pv50Sbka+Si26fX+whowpnUg6BrnuAymWygNWa7J8BYHmAbveFL
884Ycrm1xL/mnFgUzTNfpQT1E2ViZWYrwateyZ3bWziFshUuZPtlhuAlxjbn+dIt
eMWH3NdOIl+hZJ7bKGLcyJemVFZDEQz/9URHPzRwtj4Zv5Kgp9ucPXDeCtyEAFip
nZZdojYbpsT70GzRycuBNp+cmXBOWoRxmWHSRwlC2XYTYXjjVVkepMHNopLUKKms
H6iDsk/koFINJBMlnLU/S5hlAop7HzUnsRdawCkV/d78ux0zH/PXPf6lCEDUtCzn
t7ZtmcgyiH5NrOGOyYYojW8Ujtk2NgEP1B8A+i+mQ5WGtXwfK9Efo4ekYkdbdFhW
wZD/eegnouNoKRWR3hnWmbV6QJokaVmiLe+YbzqrhugVgoZGrCwXK+CserWvWBIc
DcScD+4SDF2eecqH3DWQ8bfBVbJwYcHwQ36LxlRcqO68UhINFr7yTlEp/pHBBTTm
JVTsuqFtTEHMzTOUAv3kwuXBLEZqxuZsg8VrDJebQYavf69+9C61dbLz+9PGUYaI
MtQNn7n3Ogu41SUdCbo9/7oF1fVG135t46UfF/ZItu7cbRAuo6l1sFj3jMzIUDn3
paz9IxSusKkF7GhwoVmdLtuQowxPP4dDUPW/wLThl7ghl27yZfmzxeQW/DFLfOg9
FjA8sFfbTSgT3kpB+tNvlf4WOAgOhoEPe2ZKGcvAKduzmtqgnphbnjFNPyd7G+VO
zeWqilalkgznAYymVdgcnT/wctNw5spGqziNiQhLm6XSOR2hEcpGtbvRiw+ZmO48
3Fsul14egzEz+TYGfdLcE3bpDNPJidGkbgrK0p9uFKUsFIIOsCj6ZvtM6EyABvTW
J1zfnQ+fEhNn1Zy0ovE1qGP0sk0IJZ1e9ocRJjNWGGcJdoiEyGXVBJF4/bf+477l
KI4IDdof9RgqkEkK1lCuTw0NXfDVqeYWXmVH2ag4SpzFuezsKJKb/7IzOv8Qme4N
umLVcFFuFkQqyGX241MYbTNiVtmOvaiVXBxmRvgLEBH/ugzeAfuOVL1jyAFeOAy4
AkgbuWWuLiP2+Ywso9e5q0jnnwwRbMCw+XJfBhAkz7RaiZV7grFJYa6yz1gA3CIt
V6HAf7lvRfw8P18k+uiDo+pzaSeZs/N9efMF+EaWwPDOeXcHDZkCsm0LwhMbQncn
kXdx2gXyo+D76EQQIL/4fp0NdNakhMsTjQ/V8Ju9zHq1I3Kx6lknEQcxM8CYNbbS
Nbh9EC9tvdPIqk1t6R4ZS+pZY0RQXQZse66GIElKqCSsCsFOw+Z0gsSQFJB6x4IV
kRVL9Wtfn/8uLNdrwfFQEzGbRMQqCyLocUavLqSVRpYj6CDNCmFm9+Ec7aW1fFc4
8XdkWcqkFXbpzzYqgXtQZ51xREHwzYtBhYEwGDrQG7sl5Mg+4wHOKYP4zPoVtc6B
sQP0/zqSPbqfz8ulMeHaaNryyPfvjeXLC3FJ1WA35N3TL3MNvQm8v6qZqob+o6ZC
R+iObqyRUfKTHwYQXO5M5Y9T24yeSS6iNwj5qrHkQTxRtd8ZmWpJmKJf+vVreMh5
UdOSKjvSAUjBu1cva07JIvoC+OPGI6LV8AU/OQRFH76LY2lsxPCT2zDWIz+OUVOb
GmQE+Ex7gtdcyXEsfdL4vfobh9hOF3wSyAzjC2eMF0FDVPdmgVkHxQZpkt2eMcaM
UtsWslTMK6WJgKY86cEcimH+dVyno2O6Cxh0qIk8UM51sakRoulMiYr2s9Omz3fc
iLSYIYDj0/a1RRi1g4CTSa6SafJFTuo+j871EtVXAGHmivluALYkH+KgyiRMZkzA
kgy1rF/kcI/m+/d7RQsMupgBSHCzf/4ag3ud+fIksAUHzWqxawc2Oo/0K2Vq7qFY
ZP25NL0JM8U/gVjHDTDfC/33vVGPEPObzqJFfyqndKNfzwMb9NxXzCqtTf0H8wnk
o8h8Visgcqn9VJSi7226xhTbQz6YHtz5v0o/TEWhjlHRYCaBNxiKJ32r3DNrmHNr
UdbX7Dcs/O2Ww91CxJFux/kHI6xsOx+UzuJysgp89jfOV/NRqEKTdZvAEsNFBgXk
2NUGsAQy5XLmorpEFULYk/ngC3/7KwIyo0GDY2hqTaJ15OtLZz07bt9SqSUdvdSR
D9gzpyjhkWCX3u7+S0OU/B3h7LXE+TAswYTr5+UOFkIIPZmqVxWBr5YdXVRlnrYB
miW1fTOk39CvEV3hq0zYQ58uqs+NwRGQ4CN4g0ikUvT7oRhan40ybygSUvAIIGUw
GZJklqwIYGyZbCChN30GurFZVg60mkqufuv7q5cKYewF42MRJK5NBwkYT43mwNGm
j4Kt7uCT2NB9+nHKDCbBWbYvX8QOaGf8yc/Y+P4iQcx0tTisr0M29QHEHqrXh3nV
y8x7SSNAEgsklpk4VyoJdTVXQ//OnVs/SmC0pvcV13513KTOBQUbOT/Hq8F1e83T
mQUoYGKtwWTICQzclvY3iuwYrVKCnx1QvWVXQWK1YrADGwsgj8mghFIot4s4p9Rb
9Hqy1aga1w34+gLTiKR/E67YDbA2ESeGh0M6W+2qsVSf79vIMrbl4nR0lzoOspmR
bmAnVVFi6P9W4JVPPZr/2f8atb7YivVie8TurPatvbXe2TF+zoTzkaiEg94MKFtw
30zxKDc2Jie5TV556slAQwYfxFOrIZULPpea/iFty1mRi0rwu5QCMRkuHdAwc3Vd
eENahjGvc4C+qiKUWpcK4eVNLkpGBhwxB+ozwOSQDGGtZtZ0cO2e0fLyREUxtj/j
AaraDWPRoi19blr2kd6pC/EqMtdSyHNrFyJwoE4DjdNlvfwvpw7IpdmWnlRF73r9
vec2cs0+Si9bpi0do8xZqW9B5Hd/M8OXe0ATdkinoq/G3ccdhUfmdex4RRaHU2Qr
TQDniIWx75AN4+u3TqD1uNEwuPJbdLDCNp3blqnlanroKVjuddPTmBRm9Es2GBwZ
ZIzwWiBAn/eoICpyQCwd2Roj2RyJjIKAzmimjALzTV8IjFsSnBAi3yP8S8uf8prb
i1HzGAxTAeFX+d8V16pHgGgwgBfTKP5VNLjls5ETbZH9y/yPa5tQDAWPAQcURMqE
YSCC5m3+5xDkpUPN+q5roRIAK8Yy3+Pl/ZMYbTmwPmZwoqytvzqTfaz7GuT6TxWv
Olgh7LyciDBvWtjSZadrh8PS7PvdxeBD1QA67OZz3gDJhnBoYkIe8tTzt4qtJHC8
FuPEftAGlqb3Xi+RYknUjlwN9mgCXXK3ggB5nyCVL1qCHt4VaCtyb1O/ffegZMk4
ho1uXWYHn9Yr0aW3iNRfBm8HLVZD4hR6Dzsig6oLHjGlcQo8WziFGn53fmyVxVuB
gOI6tnDsXzfPO+ixU9KnkDzmsvoKKdWk9TGJOqRBtlxW3Bf+TWY1QXFsrsL2yKhc
Um1/FRcvcxtrn/FFdcOsLOdhjZCff0M4HVUBbGMNaXXP0UaCL3HaPJE+IwQwkR76
pUNEAVY8zMvvK4vjFd2BfPC4ddAB+HV3ah0bqeo99Fc170NR6j6Y29AwUxeoo1Wz
sh5Agfj5g+UpIcArGnUAUFukVRLkIhkoIs+ZrlCeKZl4epc4t1+L6mpGhom2QSAk
OgeQwNWOWjhgOB6Olp99BQHTwz2V955ZCBhw2A+gdnJqsUldeScM2Ylcj+kQk7fH
P1KhG/AsCuiqMkd0M4Z+VLghyfFQgxvCD3Hnxr8tiqtf0sP8sNSEb8v4yOqmZBlG
vlLeqA1pm10zE66BdFGh1RC0I3d3eEmMl2zCY1TcfHPnfW0ATvpEYqSegofsyQHB
QF0nbsxI8gxVAk50bFqvKc6zgGeOoKVlj79CKzAXsCdSDhY6jQ1aa+g5DO+IvfPI
YadgvnCI3HtYi5yXTaPPI+iPdtUNGipXUGIWnDbVHwwN/1ROE2yPxbzRWhQYyDAX
c/2CO7qE3ShQwuukv+4/tcOnEXfnU6LHlOqMPB1H0Oc5mbxtRTAA+klidT1ut4qr
18lP0DAg7CBBrZhnS0/mnkbO9QdCEiG+vQWWtZMdHjX4aPqlrQzoO23KRNCFZIFY
iyKsfNEncWoq2d9chDovNGc1RGlHRPzwyAyUzv6s4HyOrmzm0IySZospOxVm4jID
k+5nJNUGeFTr1I0mFlC8RH+VMhnJEGzwtHKNyC+/wJg4T78FSvxtj7wflzv90XPP
9GUE6r3YcuFe360iJTnOS+VVldnCmdRPdYI16mZOxd4k6iSqSwA/PORQ7mnaiSQB
av+domcqSIs69njAZaRbH/eGKzqswi8MIE28kNjvRqdjlSvJCGevN58Gtzd7lmJU
BMXirkn6lngXV+8Ka8zef5BmYxwjvnziaova4PFBSO/l4iyvryMQUhsaZFBwKl7g
vHI+gE0ddBbc2BpgNseaHnIHe+HTT/LAuiaaO4V1QW/vsCBYtr8/oObwCOgAlCF9
CjtHoTOymIg3g6GYBFk6tZ35iwQ4YYx2lEwwL/TjG1cwfOFC2T0TEatAi6Vi6vg+
TyBuy94anoj0D1u7A3Vw0C8/1BYB8u/CNi59wYfsLYp7j+xmnQwJZvetu9aUeXLY
3qagvFV7xDq9hpIemh/24UZ3P3YZAxqLkJ68Hb/KwGA0ELUSINpOWrmd851zgLsK
RBKGWqcYhzqcRoKvmgVX9XmvHfShhroWhljsNSD+8o1qGOTG2cy4qY23nd2t2lrk
KefhnDPDzcvPKThaeVMQ0ficyvj4RwlqAlcoHRSrMBBRXpb2fOfMD43oeXGNVrBl
7hTEYARDBCeAwLflWAJO/0YQ83bc60IrHRKgaoNsMPI9fSLRD7yNzuoO7B+zE1mr
WeyhslB5Yn5SR+iU+A7CMGdIQiXjipTP0GxSMd+gD2GYdw4A/hnfYTjfXjzuc8QO
WuukQty/wccbcXmZTvXTR7wxpl2k1Q5YNZOAivLFbDCOuKmCIoDPTMrzqWfsBijD
vJ/BGKjjWPrYDEdAC+M5cBC6mx/ce5MCfxczj7NBaq86H95ViEWFlcXsuFJ+L11h
XnhGgVMAnpJ72TAU7nOROzggtX2A+byHyWHMH4pfsJTdwdN53Kxs3qKddlpPOrou
0G1LduAaxK+nnIGzoWEfeqe1jl7rNtwBjQAgtboBNUsouZkOAG2tYDYGH/0Dwnpz
ts/lGZjn4YyY13KH7ZtwKCNXQ3mkb7Japp+PjOpBar4kvdBXdvaCQBQ71KbUrLdG
Ti54XrjUYUYuKjgeWHWuFpEovVSfzlrszJdM5RXRACS6v6kWQUlVHQPtGGFUaTtS
VL9DOzO8AxpFxFs9GcqsgI9JEICaja5cCwOcNr+vmjYY8zsoXU9Zdx+BSNhayaDA
bEcFJbOFMAc2neQ8jGggA8Y2XDO3xWF7KR47vzfytDx+MUtHW38yG/7CXK8NY4DA
tvcpVxnrT4DRIwe3yZvQc3n17yBBDHA4Is3WQ9rQwe65DImu8qQbN+bjVk2n1KQf
Ktk+6i1y5DoF4f0YNxOvxcWRwzmsrIemDDohyisxV73YGLKzaBJz5/OwIcFEewAt
Sdp56VFOOix/QmaoPZf81hTwSNecnIUwaFBPF9g6apdngqS1JoUywGmGy+vmqQ9R
JTDmSVmD0b2835+kTKGQsC5TPuGR8KBiVb1ewlR4hmbH/ypFzfgl0rsEjJN03tRw
Y6oczdzLekeftWPcXm6iM8HTClcF2m83V7QkxoMSpXJvE1Ug7n5pHHviYE/m2RtC
USad/gbky2OK9zXrFoeBQu+rfoatQGL+07hiidAYTA3BOaUYxsBCLqUAl0C/lPih
CQ2TqQTp1FmOMYOlGA+Tm8lBQo+qVsZ/m7x1CAttS3Da6iSN6H2//wF9WoGKkGGq
fktqjnpdyW1K7yKhSiMFU9nqR7ErN6JFyN4hqsMqR8WWJVSTTp82O/47e/l6pO4r
d680GoVNmfjwsl1kuICGPAeTQnjZCjyhgWsPauuflV6bEM8ETNuEYX/o8xcVPdfI
cd1Rfu16WkmCuRA8H68guOdQKWsHuAs5IuLYtJOOpA1kLwBmkxl2C3JuGJML5AzY
qZ931YgYe9PfXiGAYdz2bLpbjOtMitRTGlelt6+CqQi4jIClLZi3f5RfHZ/zCuXK
WmwpaaWbJb8rs+sWguyDKZGC5ArU8WhqB6/4D+WhUlhzsxUirEvGjW7Y7KjI4cwz
VdTFJBjt20r3boB5AbayUNhryYwJGPybwlxe2+3m2f2VnqTjROJnIrqfCNA0nF50
s8TE4p3rac5hh7cDfuloOB5ALWw6XPhIg1x56as7vN5+LPmKAsyogg4yXYbfOoDY
HoKFLam3jzwYPR8AabkeBmUkOy5UsECzAI+UVWKpsaf2SCDe6CcmAZNe4Xxs0TCQ
wkgI7k3TzrNwoOTUD1+Gg2azPGfoCdEa1HyE+ol4ezjR2GSNZ/L4qZDWNt2GiVa8
DhyOUnF0F1qoOTGhkF6odRTzstLSR8VtgpJTkoe/xnAHOxgK6sXtBJC8vOQfIMqb
9hNZUVg1PBzUv9wzeqJB7tHLc41IogWyyo2rQZM6xfHJrnM3X6QvtnrGnct+8wm1
NjFpc+2QBPs40Jj7RhzjsDNoMC99yU8VfFXvN9PVx8mWQzuCgUNRT7rAWLMq0260
9/NLb7G/0xQPKlWVOq1wDYMM6k0IUtvMkXVu/DCPkTf2kBnduP5+YgkMuYq5L4ZH
6gPgZYSIMbab0VTv+JfqV9VFyWh7R2oVckC/lIp6JcRG2YUVLZlp8WfWg5Ycp9uL
iqUyRUZvaFDVgYqF2dc/+ZPrUyIe1G3ulvnrYV+WzB6t4n7j1cV5Y9RY2+kCCy69
dl4QlPqM5nOyi7uhYEJqQIbzppMS46AHKKo0Ex4oA2dU5H2y5fc6ZItr6GShsODh
+/cuTHmpYnstgBVx2C6ZH1aDD9TJBh6XUsjRfJbH1URUPqeJJvx2oFLI2rVKy/1S
SMYsVAvPcUp4zfhHuc60jQ==
`pragma protect end_protected
