-- xcvr_8B10B.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
library xcvr_8B10B_altera_xcvr_atx_pll_a10_181;
library xcvr_8B10B_altera_xcvr_native_a10_181;
library xcvr_8B10B_altera_xcvr_reset_control_181;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity xcvr_8B10B is
	port (
		clk_clk                                                             : in  std_logic                      := '0';             --                                          clk.clk
		reset_reset_n                                                       : in  std_logic                      := '0';             --                                        reset.reset_n
		xcvr_native_a10_0_rx_clkout_ch0_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_rx_clkout_ch0.clk
		xcvr_native_a10_0_rx_clkout_ch1_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_rx_clkout_ch1.clk
		xcvr_native_a10_0_rx_clkout_ch2_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_rx_clkout_ch2.clk
		xcvr_native_a10_0_rx_clkout_ch3_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_rx_clkout_ch3.clk
		xcvr_native_a10_0_rx_coreclkin_ch0_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_rx_coreclkin_ch0.clk
		xcvr_native_a10_0_rx_coreclkin_ch1_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_rx_coreclkin_ch1.clk
		xcvr_native_a10_0_rx_coreclkin_ch2_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_rx_coreclkin_ch2.clk
		xcvr_native_a10_0_rx_coreclkin_ch3_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_rx_coreclkin_ch3.clk
		xcvr_native_a10_0_rx_parallel_data_ch0_rx_parallel_data             : out std_logic_vector(19 downto 0);                     --       xcvr_native_a10_0_rx_parallel_data_ch0.rx_parallel_data
		xcvr_native_a10_0_rx_parallel_data_ch1_rx_parallel_data             : out std_logic_vector(19 downto 0);                     --       xcvr_native_a10_0_rx_parallel_data_ch1.rx_parallel_data
		xcvr_native_a10_0_rx_parallel_data_ch2_rx_parallel_data             : out std_logic_vector(19 downto 0);                     --       xcvr_native_a10_0_rx_parallel_data_ch2.rx_parallel_data
		xcvr_native_a10_0_rx_parallel_data_ch3_rx_parallel_data             : out std_logic_vector(19 downto 0);                     --       xcvr_native_a10_0_rx_parallel_data_ch3.rx_parallel_data
		xcvr_native_a10_0_rx_patterndetect_ch0_rx_patterndetect             : out std_logic_vector(1 downto 0);                      --       xcvr_native_a10_0_rx_patterndetect_ch0.rx_patterndetect
		xcvr_native_a10_0_rx_patterndetect_ch1_rx_patterndetect             : out std_logic_vector(1 downto 0);                      --       xcvr_native_a10_0_rx_patterndetect_ch1.rx_patterndetect
		xcvr_native_a10_0_rx_patterndetect_ch2_rx_patterndetect             : out std_logic_vector(1 downto 0);                      --       xcvr_native_a10_0_rx_patterndetect_ch2.rx_patterndetect
		xcvr_native_a10_0_rx_patterndetect_ch3_rx_patterndetect             : out std_logic_vector(1 downto 0);                      --       xcvr_native_a10_0_rx_patterndetect_ch3.rx_patterndetect
		xcvr_native_a10_0_rx_serial_data_ch0_rx_serial_data                 : in  std_logic                      := '0';             --         xcvr_native_a10_0_rx_serial_data_ch0.rx_serial_data
		xcvr_native_a10_0_rx_serial_data_ch1_rx_serial_data                 : in  std_logic                      := '0';             --         xcvr_native_a10_0_rx_serial_data_ch1.rx_serial_data
		xcvr_native_a10_0_rx_serial_data_ch2_rx_serial_data                 : in  std_logic                      := '0';             --         xcvr_native_a10_0_rx_serial_data_ch2.rx_serial_data
		xcvr_native_a10_0_rx_serial_data_ch3_rx_serial_data                 : in  std_logic                      := '0';             --         xcvr_native_a10_0_rx_serial_data_ch3.rx_serial_data
		xcvr_native_a10_0_rx_seriallpbken_ch0_rx_seriallpbken               : in  std_logic                      := '0';             --        xcvr_native_a10_0_rx_seriallpbken_ch0.rx_seriallpbken
		xcvr_native_a10_0_rx_seriallpbken_ch1_rx_seriallpbken               : in  std_logic                      := '0';             --        xcvr_native_a10_0_rx_seriallpbken_ch1.rx_seriallpbken
		xcvr_native_a10_0_rx_seriallpbken_ch2_rx_seriallpbken               : in  std_logic                      := '0';             --        xcvr_native_a10_0_rx_seriallpbken_ch2.rx_seriallpbken
		xcvr_native_a10_0_rx_seriallpbken_ch3_rx_seriallpbken               : in  std_logic                      := '0';             --        xcvr_native_a10_0_rx_seriallpbken_ch3.rx_seriallpbken
		xcvr_native_a10_0_rx_std_wa_patternalign_ch0_rx_std_wa_patternalign : in  std_logic                      := '0';             -- xcvr_native_a10_0_rx_std_wa_patternalign_ch0.rx_std_wa_patternalign
		xcvr_native_a10_0_rx_std_wa_patternalign_ch1_rx_std_wa_patternalign : in  std_logic                      := '0';             -- xcvr_native_a10_0_rx_std_wa_patternalign_ch1.rx_std_wa_patternalign
		xcvr_native_a10_0_rx_std_wa_patternalign_ch2_rx_std_wa_patternalign : in  std_logic                      := '0';             -- xcvr_native_a10_0_rx_std_wa_patternalign_ch2.rx_std_wa_patternalign
		xcvr_native_a10_0_rx_std_wa_patternalign_ch3_rx_std_wa_patternalign : in  std_logic                      := '0';             -- xcvr_native_a10_0_rx_std_wa_patternalign_ch3.rx_std_wa_patternalign
		xcvr_native_a10_0_rx_syncstatus_ch0_rx_syncstatus                   : out std_logic_vector(1 downto 0);                      --          xcvr_native_a10_0_rx_syncstatus_ch0.rx_syncstatus
		xcvr_native_a10_0_rx_syncstatus_ch1_rx_syncstatus                   : out std_logic_vector(1 downto 0);                      --          xcvr_native_a10_0_rx_syncstatus_ch1.rx_syncstatus
		xcvr_native_a10_0_rx_syncstatus_ch2_rx_syncstatus                   : out std_logic_vector(1 downto 0);                      --          xcvr_native_a10_0_rx_syncstatus_ch2.rx_syncstatus
		xcvr_native_a10_0_rx_syncstatus_ch3_rx_syncstatus                   : out std_logic_vector(1 downto 0);                      --          xcvr_native_a10_0_rx_syncstatus_ch3.rx_syncstatus
		xcvr_native_a10_0_tx_clkout_ch0_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_tx_clkout_ch0.clk
		xcvr_native_a10_0_tx_clkout_ch1_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_tx_clkout_ch1.clk
		xcvr_native_a10_0_tx_clkout_ch2_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_tx_clkout_ch2.clk
		xcvr_native_a10_0_tx_clkout_ch3_clk                                 : out std_logic;                                         --              xcvr_native_a10_0_tx_clkout_ch3.clk
		xcvr_native_a10_0_tx_coreclkin_ch0_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_tx_coreclkin_ch0.clk
		xcvr_native_a10_0_tx_coreclkin_ch1_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_tx_coreclkin_ch1.clk
		xcvr_native_a10_0_tx_coreclkin_ch2_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_tx_coreclkin_ch2.clk
		xcvr_native_a10_0_tx_coreclkin_ch3_clk                              : in  std_logic                      := '0';             --           xcvr_native_a10_0_tx_coreclkin_ch3.clk
		xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data             : in  std_logic_vector(19 downto 0)  := (others => '0'); --       xcvr_native_a10_0_tx_parallel_data_ch0.tx_parallel_data
		xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data             : in  std_logic_vector(19 downto 0)  := (others => '0'); --       xcvr_native_a10_0_tx_parallel_data_ch1.tx_parallel_data
		xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data             : in  std_logic_vector(19 downto 0)  := (others => '0'); --       xcvr_native_a10_0_tx_parallel_data_ch2.tx_parallel_data
		xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data             : in  std_logic_vector(19 downto 0)  := (others => '0'); --       xcvr_native_a10_0_tx_parallel_data_ch3.tx_parallel_data
		xcvr_native_a10_0_tx_serial_data_ch0_tx_serial_data                 : out std_logic;                                         --         xcvr_native_a10_0_tx_serial_data_ch0.tx_serial_data
		xcvr_native_a10_0_tx_serial_data_ch1_tx_serial_data                 : out std_logic;                                         --         xcvr_native_a10_0_tx_serial_data_ch1.tx_serial_data
		xcvr_native_a10_0_tx_serial_data_ch2_tx_serial_data                 : out std_logic;                                         --         xcvr_native_a10_0_tx_serial_data_ch2.tx_serial_data
		xcvr_native_a10_0_tx_serial_data_ch3_tx_serial_data                 : out std_logic;                                         --         xcvr_native_a10_0_tx_serial_data_ch3.tx_serial_data
		xcvr_native_a10_0_unused_rx_parallel_data_unused_rx_parallel_data   : out std_logic_vector(415 downto 0);                    --    xcvr_native_a10_0_unused_rx_parallel_data.unused_rx_parallel_data
		xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data   : in  std_logic_vector(431 downto 0) := (others => '0'); --    xcvr_native_a10_0_unused_tx_parallel_data.unused_tx_parallel_data
		xcvr_reset_control_0_clock_clk                                      : in  std_logic                      := '0';             --                   xcvr_reset_control_0_clock.clk
		xcvr_reset_control_0_pll_select_pll_select                          : in  std_logic_vector(0 downto 0)   := (others => '0'); --              xcvr_reset_control_0_pll_select.pll_select
		xcvr_reset_control_0_reset_reset                                    : in  std_logic                      := '0';             --                   xcvr_reset_control_0_reset.reset
		xcvr_reset_control_0_rx_ready0_rx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_rx_ready0.rx_ready
		xcvr_reset_control_0_rx_ready1_rx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_rx_ready1.rx_ready
		xcvr_reset_control_0_rx_ready2_rx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_rx_ready2.rx_ready
		xcvr_reset_control_0_rx_ready3_rx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_rx_ready3.rx_ready
		xcvr_reset_control_0_tx_ready0_tx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_tx_ready0.tx_ready
		xcvr_reset_control_0_tx_ready1_tx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_tx_ready1.tx_ready
		xcvr_reset_control_0_tx_ready2_tx_ready                             : out std_logic;                                         --               xcvr_reset_control_0_tx_ready2.tx_ready
		xcvr_reset_control_0_tx_ready3_tx_ready                             : out std_logic                                          --               xcvr_reset_control_0_tx_ready3.tx_ready
	);
end entity xcvr_8B10B;

architecture rtl of xcvr_8B10B is
	component xcvr_8B10B_altera_xcvr_atx_pll_a10_181_ubmonnq is
		generic (
			enable_pll_reconfig                                              : integer := 0;
			rcfg_jtag_enable                                                 : integer := 0;
			rcfg_separate_avmm_busy                                          : integer := 0;
			dbg_embedded_debug_enable                                        : integer := 0;
			dbg_capability_reg_enable                                        : integer := 0;
			dbg_user_identifier                                              : integer := 0;
			dbg_stat_soft_logic_enable                                       : integer := 0;
			dbg_ctrl_soft_logic_enable                                       : integer := 0;
			rcfg_emb_strm_enable                                             : integer := 0;
			rcfg_profile_cnt                                                 : integer := 2;
			hssi_pma_lc_refclk_select_mux_powerdown_mode                     : string  := "powerup";
			hssi_pma_lc_refclk_select_mux_refclk_select                      : string  := "ref_iqclk0";
			hssi_pma_lc_refclk_select_mux_silicon_rev                        : string  := "20nm5es";
			hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping : string  := "ref_iqclk0";
			hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping : string  := "ref_iqclk0";
			hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping : string  := "ref_iqclk0";
			hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping : string  := "ref_iqclk0";
			hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping : string  := "ref_iqclk0";
			hssi_refclk_divider_silicon_rev                                  : string  := "20nm5es";
			atx_pll_silicon_rev                                              : string  := "20nm5es";
			atx_pll_is_cascaded_pll                                          : string  := "false";
			atx_pll_cgb_div                                                  : integer := 1;
			atx_pll_pma_width                                                : integer := 8;
			atx_pll_cp_compensation_enable                                   : string  := "true";
			atx_pll_cp_current_setting                                       : string  := "cp_current_setting0";
			atx_pll_cp_testmode                                              : string  := "cp_normal";
			atx_pll_cp_lf_3rd_pole_freq                                      : string  := "lf_3rd_pole_setting0";
			atx_pll_lf_cbig_size                                             : string  := "lf_cbig_setting0";
			atx_pll_cp_lf_order                                              : string  := "lf_2nd_order";
			atx_pll_lf_resistance                                            : string  := "lf_setting0";
			atx_pll_lf_ripplecap                                             : string  := "lf_ripple_cap_0";
			atx_pll_tank_sel                                                 : string  := "lctank0";
			atx_pll_tank_band                                                : string  := "lc_band0";
			atx_pll_tank_voltage_coarse                                      : string  := "vreg_setting_coarse0";
			atx_pll_tank_voltage_fine                                        : string  := "vreg_setting5";
			atx_pll_output_regulator_supply                                  : string  := "vreg1v_setting3";
			atx_pll_overrange_voltage                                        : string  := "over_setting5";
			atx_pll_underrange_voltage                                       : string  := "under_setting4";
			atx_pll_fb_select                                                : string  := "direct_fb";
			atx_pll_d2a_voltage                                              : string  := "d2a_disable";
			atx_pll_dsm_mode                                                 : string  := "dsm_mode_integer";
			atx_pll_dsm_out_sel                                              : string  := "pll_dsm_disable";
			atx_pll_dsm_ecn_bypass                                           : string  := "false";
			atx_pll_dsm_ecn_test_en                                          : string  := "false";
			atx_pll_dsm_fractional_division                                  : string  := "0";
			atx_pll_dsm_fractional_value_ready                               : string  := "pll_k_ready";
			atx_pll_iqclk_mux_sel                                            : string  := "power_down";
			atx_pll_vco_bypass_enable                                        : string  := "false";
			atx_pll_l_counter                                                : integer := 1;
			atx_pll_l_counter_enable                                         : string  := "false";
			atx_pll_cascadeclk_test                                          : string  := "cascadetest_off";
			atx_pll_hclk_divide                                              : integer := 1;
			atx_pll_enable_hclk                                              : string  := "hclk_disabled";
			atx_pll_m_counter                                                : integer := 8;
			atx_pll_ref_clk_div                                              : integer := 1;
			atx_pll_bw_sel                                                   : string  := "low";
			atx_pll_datarate                                                 : string  := "0 bps";
			atx_pll_device_variant                                           : string  := "device1";
			atx_pll_initial_settings                                         : string  := "true";
			atx_pll_lc_mode                                                  : string  := "lccmu_pd";
			atx_pll_output_clock_frequency                                   : string  := "0 hz";
			atx_pll_powerdown_mode                                           : string  := "powerup";
			atx_pll_prot_mode                                                : string  := "basic_tx";
			atx_pll_reference_clock_frequency                                : string  := "0 hz";
			atx_pll_sup_mode                                                 : string  := "user_mode";
			atx_pll_regulator_bypass                                         : string  := "reg_enable";
			atx_pll_vco_freq                                                 : string  := "0 hz";
			atx_pll_is_otn                                                   : string  := "false";
			atx_pll_is_sdi                                                   : string  := "false";
			atx_pll_primary_use                                              : string  := "hssi_x1";
			atx_pll_fpll_refclk_selection                                    : string  := "select_div_by_2";
			atx_pll_lc_to_fpll_l_counter_scratch                             : integer := 1;
			atx_pll_lc_to_fpll_l_counter                                     : string  := "lcounter_setting0";
			atx_pll_pfd_delay_compensation                                   : string  := "normal_delay";
			atx_pll_xcpvco_xchgpmplf_cp_current_boost                        : string  := "normal_setting";
			atx_pll_pfd_pulse_width                                          : string  := "pulse_width_setting0";
			hip_cal_en                                                       : string  := "disable";
			calibration_en                                                   : string  := "enable";
			enable_analog_resets                                             : integer := 0;
			atx_pll_bonding_mode                                             : string  := "";
			enable_mcgb                                                      : integer := 0;
			enable_mcgb_debug_ports_parameters                               : integer := 0;
			hssi_pma_cgb_master_prot_mode                                    : string  := "";
			hssi_pma_cgb_master_silicon_rev                                  : string  := "";
			hssi_pma_cgb_master_x1_div_m_sel                                 : string  := "";
			hssi_pma_cgb_master_cgb_enable_iqtxrxclk                         : string  := "";
			hssi_pma_cgb_master_ser_mode                                     : string  := "";
			hssi_pma_cgb_master_datarate                                     : string  := "";
			hssi_pma_cgb_master_cgb_power_down                               : string  := "normal_cgb";
			hssi_pma_cgb_master_observe_cgb_clocks                           : string  := "observe_nothing";
			hssi_pma_cgb_master_op_mode                                      : string  := "enabled";
			hssi_pma_cgb_master_tx_ucontrol_reset_pcie                       : string  := "pcscorehip_controls_mcgb";
			hssi_pma_cgb_master_vccdreg_output                               : string  := "vccdreg_nominal";
			hssi_pma_cgb_master_input_select                                 : string  := "fpll_top";
			hssi_pma_cgb_master_input_select_gen3                            : string  := "unused"
		);
		port (
			pll_powerdown           : in  std_logic                     := 'X';             -- pll_powerdown
			pll_refclk0             : in  std_logic                     := 'X';             -- clk
			tx_serial_clk           : out std_logic;                                        -- clk
			pll_locked              : out std_logic;                                        -- pll_locked
			pll_cal_busy            : out std_logic;                                        -- pll_cal_busy
			pll_refclk1             : in  std_logic                     := 'X';             -- clk
			pll_refclk2             : in  std_logic                     := 'X';             -- clk
			pll_refclk3             : in  std_logic                     := 'X';             -- clk
			pll_refclk4             : in  std_logic                     := 'X';             -- clk
			tx_serial_clk_gt        : out std_logic;                                        -- clk
			pll_pcie_clk            : out std_logic;                                        -- pll_pcie_clk
			pll_cascade_clk         : out std_logic;                                        -- clk
			atx_to_fpll_cascade_clk : out std_logic;                                        -- clk
			reconfig_clk0           : in  std_logic                     := 'X';             -- clk
			reconfig_reset0         : in  std_logic                     := 'X';             -- reset
			reconfig_write0         : in  std_logic                     := 'X';             -- write
			reconfig_read0          : in  std_logic                     := 'X';             -- read
			reconfig_address0       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			reconfig_writedata0     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_readdata0      : out std_logic_vector(31 downto 0);                    -- readdata
			reconfig_waitrequest0   : out std_logic;                                        -- waitrequest
			avmm_busy0              : out std_logic;                                        -- avmm_busy0
			hip_cal_done            : out std_logic;                                        -- hip_cal_done
			clklow                  : out std_logic;                                        -- clk
			fref                    : out std_logic;                                        -- clk
			overrange               : out std_logic;                                        -- debug
			underrange              : out std_logic;                                        -- debug
			mcgb_rst                : in  std_logic                     := 'X';             -- mcgb_rst
			mcgb_aux_clk0           : in  std_logic                     := 'X';             -- tx_serial_clk
			mcgb_aux_clk1           : in  std_logic                     := 'X';             -- tx_serial_clk
			mcgb_aux_clk2           : in  std_logic                     := 'X';             -- tx_serial_clk
			tx_bonding_clocks       : out std_logic_vector(5 downto 0);                     -- clk
			mcgb_serial_clk         : out std_logic;                                        -- clk
			pcie_sw                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- pcie_sw
			pcie_sw_done            : out std_logic_vector(1 downto 0);                     -- pcie_sw_done
			reconfig_clk1           : in  std_logic                     := 'X';             -- clk
			reconfig_reset1         : in  std_logic                     := 'X';             -- reset
			reconfig_write1         : in  std_logic                     := 'X';             -- write
			reconfig_read1          : in  std_logic                     := 'X';             -- read
			reconfig_address1       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			reconfig_writedata1     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_readdata1      : out std_logic_vector(31 downto 0);                    -- readdata
			reconfig_waitrequest1   : out std_logic;                                        -- waitrequest
			mcgb_cal_busy           : out std_logic;                                        -- mcgb_cal_busy
			mcgb_hip_cal_done       : out std_logic                                         -- hip_cal_done
		);
	end component xcvr_8B10B_altera_xcvr_atx_pll_a10_181_ubmonnq;

	component xcvr_8B10B_altera_xcvr_native_a10_181_b5mzony is
		generic (
			device_revision                                                        : string  := "20nm5es";
			duplex_mode                                                            : string  := "duplex";
			channels                                                               : integer := 1;
			enable_calibration                                                     : integer := 0;
			enable_analog_resets                                                   : integer := 1;
			enable_reset_sequence                                                  : integer := 0;
			bonded_mode                                                            : string  := "not_bonded";
			pcs_bonding_master                                                     : integer := 0;
			plls                                                                   : integer := 1;
			number_physical_bonding_clocks                                         : integer := 1;
			cdr_refclk_cnt                                                         : integer := 1;
			enable_hip                                                             : integer := 0;
			hip_cal_en                                                             : string  := "disable";
			rcfg_enable                                                            : integer := 0;
			rcfg_shared                                                            : integer := 0;
			rcfg_jtag_enable                                                       : integer := 0;
			rcfg_separate_avmm_busy                                                : integer := 0;
			adme_prot_mode                                                         : string  := "basic_tx";
			adme_data_rate                                                         : string  := "5000000000";
			enable_pcie_dfe_ip                                                     : boolean := false;
			sim_reduced_counters                                                   : boolean := false;
			disable_continuous_dfe                                                 : boolean := false;
			dbg_embedded_debug_enable                                              : integer := 0;
			dbg_capability_reg_enable                                              : integer := 0;
			dbg_user_identifier                                                    : integer := 0;
			dbg_stat_soft_logic_enable                                             : integer := 0;
			dbg_ctrl_soft_logic_enable                                             : integer := 0;
			dbg_prbs_soft_logic_enable                                             : integer := 0;
			dbg_odi_soft_logic_enable                                              : integer := 0;
			rcfg_emb_strm_enable                                                   : integer := 0;
			rcfg_profile_cnt                                                       : integer := 2;
			hssi_gen3_rx_pcs_block_sync                                            : string  := "enable_block_sync";
			hssi_gen3_rx_pcs_block_sync_sm                                         : string  := "enable_blk_sync_sm";
			hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                                 : string  := "enable";
			hssi_gen3_rx_pcs_lpbk_force                                            : string  := "lpbk_frce_dis";
			hssi_gen3_rx_pcs_mode                                                  : string  := "gen3_func";
			hssi_gen3_rx_pcs_rate_match_fifo                                       : string  := "enable_rm_fifo_600ppm";
			hssi_gen3_rx_pcs_rate_match_fifo_latency                               : string  := "regular_latency";
			hssi_gen3_rx_pcs_reverse_lpbk                                          : string  := "rev_lpbk_en";
			hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                                      : string  := "b4gb_par_lpbk_dis";
			hssi_gen3_rx_pcs_rx_force_balign                                       : string  := "en_force_balign";
			hssi_gen3_rx_pcs_rx_ins_del_one_skip                                   : string  := "ins_del_one_skip_en";
			hssi_gen3_rx_pcs_rx_num_fixed_pat                                      : integer := 8;
			hssi_gen3_rx_pcs_rx_test_out_sel                                       : string  := "rx_test_out0";
			hssi_gen3_rx_pcs_sup_mode                                              : string  := "user_mode";
			hssi_gen3_tx_pcs_mode                                                  : string  := "gen3_func";
			hssi_gen3_tx_pcs_reverse_lpbk                                          : string  := "rev_lpbk_en";
			hssi_gen3_tx_pcs_sup_mode                                              : string  := "user_mode";
			hssi_gen3_tx_pcs_tx_bitslip                                            : integer := 0;
			hssi_gen3_tx_pcs_tx_gbox_byp                                           : string  := "bypass_gbox";
			hssi_krfec_rx_pcs_blksync_cor_en                                       : string  := "detect";
			hssi_krfec_rx_pcs_bypass_gb                                            : string  := "bypass_dis";
			hssi_krfec_rx_pcs_clr_ctrl                                             : string  := "both_enabled";
			hssi_krfec_rx_pcs_ctrl_bit_reverse                                     : string  := "ctrl_bit_reverse_dis";
			hssi_krfec_rx_pcs_data_bit_reverse                                     : string  := "data_bit_reverse_dis";
			hssi_krfec_rx_pcs_dv_start                                             : string  := "with_blklock";
			hssi_krfec_rx_pcs_err_mark_type                                        : string  := "err_mark_10g";
			hssi_krfec_rx_pcs_error_marking_en                                     : string  := "err_mark_dis";
			hssi_krfec_rx_pcs_low_latency_en                                       : string  := "disable";
			hssi_krfec_rx_pcs_lpbk_mode                                            : string  := "lpbk_dis";
			hssi_krfec_rx_pcs_parity_invalid_enum                                  : integer := 8;
			hssi_krfec_rx_pcs_parity_valid_num                                     : integer := 4;
			hssi_krfec_rx_pcs_pipeln_blksync                                       : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_descrm                                        : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errcorrect                                    : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_ind                                   : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_lfsr                                  : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_loc                                   : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_errtrap_pat                                   : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_gearbox                                       : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_syndrm                                        : string  := "enable";
			hssi_krfec_rx_pcs_pipeln_trans_dec                                     : string  := "enable";
			hssi_krfec_rx_pcs_prot_mode                                            : string  := "disable_mode";
			hssi_krfec_rx_pcs_receive_order                                        : string  := "receive_lsb";
			hssi_krfec_rx_pcs_rx_testbus_sel                                       : string  := "overall";
			hssi_krfec_rx_pcs_signal_ok_en                                         : string  := "sig_ok_dis";
			hssi_krfec_rx_pcs_sup_mode                                             : string  := "user_mode";
			hssi_krfec_tx_pcs_burst_err                                            : string  := "burst_err_dis";
			hssi_krfec_tx_pcs_burst_err_len                                        : string  := "burst_err_len1";
			hssi_krfec_tx_pcs_ctrl_bit_reverse                                     : string  := "ctrl_bit_reverse_dis";
			hssi_krfec_tx_pcs_data_bit_reverse                                     : string  := "data_bit_reverse_dis";
			hssi_krfec_tx_pcs_enc_frame_query                                      : string  := "enc_query_dis";
			hssi_krfec_tx_pcs_low_latency_en                                       : string  := "disable";
			hssi_krfec_tx_pcs_pipeln_encoder                                       : string  := "enable";
			hssi_krfec_tx_pcs_pipeln_scrambler                                     : string  := "enable";
			hssi_krfec_tx_pcs_prot_mode                                            : string  := "disable_mode";
			hssi_krfec_tx_pcs_sup_mode                                             : string  := "user_mode";
			hssi_krfec_tx_pcs_transcode_err                                        : string  := "trans_err_dis";
			hssi_krfec_tx_pcs_transmit_order                                       : string  := "transmit_lsb";
			hssi_krfec_tx_pcs_tx_testbus_sel                                       : string  := "overall";
			hssi_10g_rx_pcs_align_del                                              : string  := "align_del_en";
			hssi_10g_rx_pcs_ber_bit_err_total_cnt                                  : string  := "bit_err_total_cnt_10g";
			hssi_10g_rx_pcs_ber_clken                                              : string  := "ber_clk_dis";
			hssi_10g_rx_pcs_ber_xus_timer_window                                   : integer := 19530;
			hssi_10g_rx_pcs_bitslip_mode                                           : string  := "bitslip_dis";
			hssi_10g_rx_pcs_blksync_bitslip_type                                   : string  := "bitslip_comb";
			hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                               : integer := 1;
			hssi_10g_rx_pcs_blksync_bitslip_wait_type                              : string  := "bitslip_match";
			hssi_10g_rx_pcs_blksync_bypass                                         : string  := "blksync_bypass_dis";
			hssi_10g_rx_pcs_blksync_clken                                          : string  := "blksync_clk_dis";
			hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt                            : string  := "enum_invalid_sh_cnt_10g";
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock                           : string  := "knum_sh_cnt_postlock_10g";
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock                            : string  := "knum_sh_cnt_prelock_10g";
			hssi_10g_rx_pcs_blksync_pipeln                                         : string  := "blksync_pipeln_dis";
			hssi_10g_rx_pcs_clr_errblk_cnt_en                                      : string  := "disable";
			hssi_10g_rx_pcs_control_del                                            : string  := "control_del_all";
			hssi_10g_rx_pcs_crcchk_bypass                                          : string  := "crcchk_bypass_dis";
			hssi_10g_rx_pcs_crcchk_clken                                           : string  := "crcchk_clk_dis";
			hssi_10g_rx_pcs_crcchk_inv                                             : string  := "crcchk_inv_dis";
			hssi_10g_rx_pcs_crcchk_pipeln                                          : string  := "crcchk_pipeln_dis";
			hssi_10g_rx_pcs_crcflag_pipeln                                         : string  := "crcflag_pipeln_dis";
			hssi_10g_rx_pcs_ctrl_bit_reverse                                       : string  := "ctrl_bit_reverse_dis";
			hssi_10g_rx_pcs_data_bit_reverse                                       : string  := "data_bit_reverse_dis";
			hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                                 : string  := "dec_64b66b_rxsm_bypass_dis";
			hssi_10g_rx_pcs_dec64b66b_clken                                        : string  := "dec64b66b_clk_dis";
			hssi_10g_rx_pcs_descrm_bypass                                          : string  := "descrm_bypass_en";
			hssi_10g_rx_pcs_descrm_clken                                           : string  := "descrm_clk_dis";
			hssi_10g_rx_pcs_descrm_mode                                            : string  := "async";
			hssi_10g_rx_pcs_descrm_pipeln                                          : string  := "enable";
			hssi_10g_rx_pcs_dft_clk_out_sel                                        : string  := "rx_master_clk";
			hssi_10g_rx_pcs_dis_signal_ok                                          : string  := "dis_signal_ok_dis";
			hssi_10g_rx_pcs_dispchk_bypass                                         : string  := "dispchk_bypass_dis";
			hssi_10g_rx_pcs_empty_flag_type                                        : string  := "empty_rd_side";
			hssi_10g_rx_pcs_fast_path                                              : string  := "fast_path_dis";
			hssi_10g_rx_pcs_fec_clken                                              : string  := "fec_clk_dis";
			hssi_10g_rx_pcs_fec_enable                                             : string  := "fec_dis";
			hssi_10g_rx_pcs_fifo_double_read                                       : string  := "fifo_double_read_dis";
			hssi_10g_rx_pcs_fifo_stop_rd                                           : string  := "n_rd_empty";
			hssi_10g_rx_pcs_fifo_stop_wr                                           : string  := "n_wr_full";
			hssi_10g_rx_pcs_force_align                                            : string  := "force_align_dis";
			hssi_10g_rx_pcs_frmsync_bypass                                         : string  := "frmsync_bypass_dis";
			hssi_10g_rx_pcs_frmsync_clken                                          : string  := "frmsync_clk_dis";
			hssi_10g_rx_pcs_frmsync_enum_scrm                                      : string  := "enum_scrm_default";
			hssi_10g_rx_pcs_frmsync_enum_sync                                      : string  := "enum_sync_default";
			hssi_10g_rx_pcs_frmsync_flag_type                                      : string  := "all_framing_words";
			hssi_10g_rx_pcs_frmsync_knum_sync                                      : string  := "knum_sync_default";
			hssi_10g_rx_pcs_frmsync_mfrm_length                                    : integer := 2048;
			hssi_10g_rx_pcs_frmsync_pipeln                                         : string  := "frmsync_pipeln_dis";
			hssi_10g_rx_pcs_full_flag_type                                         : string  := "full_wr_side";
			hssi_10g_rx_pcs_gb_rx_idwidth                                          : string  := "width_32";
			hssi_10g_rx_pcs_gb_rx_odwidth                                          : string  := "width_66";
			hssi_10g_rx_pcs_gbexp_clken                                            : string  := "gbexp_clk_dis";
			hssi_10g_rx_pcs_low_latency_en                                         : string  := "enable";
			hssi_10g_rx_pcs_lpbk_mode                                              : string  := "lpbk_dis";
			hssi_10g_rx_pcs_master_clk_sel                                         : string  := "master_rx_pma_clk";
			hssi_10g_rx_pcs_pempty_flag_type                                       : string  := "pempty_rd_side";
			hssi_10g_rx_pcs_pfull_flag_type                                        : string  := "pfull_wr_side";
			hssi_10g_rx_pcs_phcomp_rd_del                                          : string  := "phcomp_rd_del2";
			hssi_10g_rx_pcs_pld_if_type                                            : string  := "fifo";
			hssi_10g_rx_pcs_prot_mode                                              : string  := "disable_mode";
			hssi_10g_rx_pcs_rand_clken                                             : string  := "rand_clk_dis";
			hssi_10g_rx_pcs_rd_clk_sel                                             : string  := "rd_rx_pma_clk";
			hssi_10g_rx_pcs_rdfifo_clken                                           : string  := "rdfifo_clk_dis";
			hssi_10g_rx_pcs_rx_fifo_write_ctrl                                     : string  := "blklock_stops";
			hssi_10g_rx_pcs_rx_scrm_width                                          : string  := "bit64";
			hssi_10g_rx_pcs_rx_sh_location                                         : string  := "lsb";
			hssi_10g_rx_pcs_rx_signal_ok_sel                                       : string  := "synchronized_ver";
			hssi_10g_rx_pcs_rx_sm_bypass                                           : string  := "rx_sm_bypass_dis";
			hssi_10g_rx_pcs_rx_sm_hiber                                            : string  := "rx_sm_hiber_en";
			hssi_10g_rx_pcs_rx_sm_pipeln                                           : string  := "rx_sm_pipeln_dis";
			hssi_10g_rx_pcs_rx_testbus_sel                                         : string  := "rx_fifo_testbus1";
			hssi_10g_rx_pcs_rx_true_b2b                                            : string  := "b2b";
			hssi_10g_rx_pcs_rxfifo_empty                                           : string  := "empty_default";
			hssi_10g_rx_pcs_rxfifo_full                                            : string  := "full_default";
			hssi_10g_rx_pcs_rxfifo_mode                                            : string  := "phase_comp";
			hssi_10g_rx_pcs_rxfifo_pempty                                          : integer := 2;
			hssi_10g_rx_pcs_rxfifo_pfull                                           : integer := 23;
			hssi_10g_rx_pcs_stretch_num_stages                                     : string  := "zero_stage";
			hssi_10g_rx_pcs_sup_mode                                               : string  := "user_mode";
			hssi_10g_rx_pcs_test_mode                                              : string  := "test_off";
			hssi_10g_rx_pcs_wrfifo_clken                                           : string  := "wrfifo_clk_dis";
			hssi_10g_rx_pcs_advanced_user_mode                                     : string  := "disable";
			hssi_10g_tx_pcs_bitslip_en                                             : string  := "bitslip_dis";
			hssi_10g_tx_pcs_bonding_dft_en                                         : string  := "dft_dis";
			hssi_10g_tx_pcs_bonding_dft_val                                        : string  := "dft_0";
			hssi_10g_tx_pcs_crcgen_bypass                                          : string  := "crcgen_bypass_dis";
			hssi_10g_tx_pcs_crcgen_clken                                           : string  := "crcgen_clk_dis";
			hssi_10g_tx_pcs_crcgen_err                                             : string  := "crcgen_err_dis";
			hssi_10g_tx_pcs_crcgen_inv                                             : string  := "crcgen_inv_dis";
			hssi_10g_tx_pcs_ctrl_bit_reverse                                       : string  := "ctrl_bit_reverse_dis";
			hssi_10g_tx_pcs_data_bit_reverse                                       : string  := "data_bit_reverse_dis";
			hssi_10g_tx_pcs_dft_clk_out_sel                                        : string  := "tx_master_clk";
			hssi_10g_tx_pcs_dispgen_bypass                                         : string  := "dispgen_bypass_dis";
			hssi_10g_tx_pcs_dispgen_clken                                          : string  := "dispgen_clk_dis";
			hssi_10g_tx_pcs_dispgen_err                                            : string  := "dispgen_err_dis";
			hssi_10g_tx_pcs_dispgen_pipeln                                         : string  := "dispgen_pipeln_dis";
			hssi_10g_tx_pcs_empty_flag_type                                        : string  := "empty_rd_side";
			hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                                 : string  := "enc_64b66b_txsm_bypass_dis";
			hssi_10g_tx_pcs_enc64b66b_txsm_clken                                   : string  := "enc64b66b_txsm_clk_dis";
			hssi_10g_tx_pcs_fastpath                                               : string  := "fastpath_dis";
			hssi_10g_tx_pcs_fec_clken                                              : string  := "fec_clk_dis";
			hssi_10g_tx_pcs_fec_enable                                             : string  := "fec_dis";
			hssi_10g_tx_pcs_fifo_double_write                                      : string  := "fifo_double_write_dis";
			hssi_10g_tx_pcs_fifo_reg_fast                                          : string  := "fifo_reg_fast_dis";
			hssi_10g_tx_pcs_fifo_stop_rd                                           : string  := "n_rd_empty";
			hssi_10g_tx_pcs_fifo_stop_wr                                           : string  := "n_wr_full";
			hssi_10g_tx_pcs_frmgen_burst                                           : string  := "frmgen_burst_dis";
			hssi_10g_tx_pcs_frmgen_bypass                                          : string  := "frmgen_bypass_dis";
			hssi_10g_tx_pcs_frmgen_clken                                           : string  := "frmgen_clk_dis";
			hssi_10g_tx_pcs_frmgen_mfrm_length                                     : integer := 2048;
			hssi_10g_tx_pcs_frmgen_pipeln                                          : string  := "frmgen_pipeln_dis";
			hssi_10g_tx_pcs_frmgen_pyld_ins                                        : string  := "frmgen_pyld_ins_dis";
			hssi_10g_tx_pcs_frmgen_wordslip                                        : string  := "frmgen_wordslip_dis";
			hssi_10g_tx_pcs_full_flag_type                                         : string  := "full_wr_side";
			hssi_10g_tx_pcs_gb_pipeln_bypass                                       : string  := "disable";
			hssi_10g_tx_pcs_gb_tx_idwidth                                          : string  := "width_50";
			hssi_10g_tx_pcs_gb_tx_odwidth                                          : string  := "width_32";
			hssi_10g_tx_pcs_gbred_clken                                            : string  := "gbred_clk_dis";
			hssi_10g_tx_pcs_low_latency_en                                         : string  := "enable";
			hssi_10g_tx_pcs_master_clk_sel                                         : string  := "master_tx_pma_clk";
			hssi_10g_tx_pcs_pempty_flag_type                                       : string  := "pempty_rd_side";
			hssi_10g_tx_pcs_pfull_flag_type                                        : string  := "pfull_wr_side";
			hssi_10g_tx_pcs_phcomp_rd_del                                          : string  := "phcomp_rd_del2";
			hssi_10g_tx_pcs_pld_if_type                                            : string  := "fifo";
			hssi_10g_tx_pcs_prot_mode                                              : string  := "disable_mode";
			hssi_10g_tx_pcs_pseudo_random                                          : string  := "all_0";
			hssi_10g_tx_pcs_pseudo_seed_a                                          : string  := "288230376151711743";
			hssi_10g_tx_pcs_pseudo_seed_b                                          : string  := "288230376151711743";
			hssi_10g_tx_pcs_random_disp                                            : string  := "disable";
			hssi_10g_tx_pcs_rdfifo_clken                                           : string  := "rdfifo_clk_dis";
			hssi_10g_tx_pcs_scrm_bypass                                            : string  := "scrm_bypass_dis";
			hssi_10g_tx_pcs_scrm_clken                                             : string  := "scrm_clk_dis";
			hssi_10g_tx_pcs_scrm_mode                                              : string  := "async";
			hssi_10g_tx_pcs_scrm_pipeln                                            : string  := "enable";
			hssi_10g_tx_pcs_sh_err                                                 : string  := "sh_err_dis";
			hssi_10g_tx_pcs_sop_mark                                               : string  := "sop_mark_dis";
			hssi_10g_tx_pcs_stretch_num_stages                                     : string  := "zero_stage";
			hssi_10g_tx_pcs_sup_mode                                               : string  := "user_mode";
			hssi_10g_tx_pcs_test_mode                                              : string  := "test_off";
			hssi_10g_tx_pcs_tx_scrm_err                                            : string  := "scrm_err_dis";
			hssi_10g_tx_pcs_tx_scrm_width                                          : string  := "bit64";
			hssi_10g_tx_pcs_tx_sh_location                                         : string  := "lsb";
			hssi_10g_tx_pcs_tx_sm_bypass                                           : string  := "tx_sm_bypass_dis";
			hssi_10g_tx_pcs_tx_sm_pipeln                                           : string  := "tx_sm_pipeln_dis";
			hssi_10g_tx_pcs_tx_testbus_sel                                         : string  := "tx_fifo_testbus1";
			hssi_10g_tx_pcs_txfifo_empty                                           : string  := "empty_default";
			hssi_10g_tx_pcs_txfifo_full                                            : string  := "full_default";
			hssi_10g_tx_pcs_txfifo_mode                                            : string  := "phase_comp";
			hssi_10g_tx_pcs_txfifo_pempty                                          : integer := 2;
			hssi_10g_tx_pcs_txfifo_pfull                                           : integer := 11;
			hssi_10g_tx_pcs_wr_clk_sel                                             : string  := "wr_tx_pma_clk";
			hssi_10g_tx_pcs_wrfifo_clken                                           : string  := "wrfifo_clk_dis";
			hssi_10g_tx_pcs_advanced_user_mode                                     : string  := "disable";
			hssi_8g_rx_pcs_auto_error_replacement                                  : string  := "dis_err_replace";
			hssi_8g_rx_pcs_bit_reversal                                            : string  := "dis_bit_reversal";
			hssi_8g_rx_pcs_bonding_dft_en                                          : string  := "dft_dis";
			hssi_8g_rx_pcs_bonding_dft_val                                         : string  := "dft_0";
			hssi_8g_rx_pcs_bypass_pipeline_reg                                     : string  := "dis_bypass_pipeline";
			hssi_8g_rx_pcs_byte_deserializer                                       : string  := "dis_bds";
			hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                                   : string  := "dis_rxvalid_mask";
			hssi_8g_rx_pcs_clkcmp_pattern_n                                        : integer := 0;
			hssi_8g_rx_pcs_clkcmp_pattern_p                                        : integer := 0;
			hssi_8g_rx_pcs_clock_gate_bds_dec_asn                                  : string  := "dis_bds_dec_asn_clk_gating";
			hssi_8g_rx_pcs_clock_gate_cdr_eidle                                    : string  := "dis_cdr_eidle_clk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                                  : string  := "dis_dw_pc_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_rm_rd                                     : string  := "dis_dw_rm_rdclk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_rm_wr                                     : string  := "dis_dw_rm_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_dw_wa                                        : string  := "dis_dw_wa_clk_gating";
			hssi_8g_rx_pcs_clock_gate_pc_rdclk                                     : string  := "dis_pc_rdclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                                  : string  := "dis_sw_pc_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_rm_rd                                     : string  := "dis_sw_rm_rdclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_rm_wr                                     : string  := "dis_sw_rm_wrclk_gating";
			hssi_8g_rx_pcs_clock_gate_sw_wa                                        : string  := "dis_sw_wa_clk_gating";
			hssi_8g_rx_pcs_clock_observation_in_pld_core                           : string  := "internal_sw_wa_clk";
			hssi_8g_rx_pcs_eidle_entry_eios                                        : string  := "dis_eidle_eios";
			hssi_8g_rx_pcs_eidle_entry_iei                                         : string  := "dis_eidle_iei";
			hssi_8g_rx_pcs_eidle_entry_sd                                          : string  := "dis_eidle_sd";
			hssi_8g_rx_pcs_eightb_tenb_decoder                                     : string  := "dis_8b10b";
			hssi_8g_rx_pcs_err_flags_sel                                           : string  := "err_flags_wa";
			hssi_8g_rx_pcs_fixed_pat_det                                           : string  := "dis_fixed_patdet";
			hssi_8g_rx_pcs_fixed_pat_num                                           : integer := 15;
			hssi_8g_rx_pcs_force_signal_detect                                     : string  := "en_force_signal_detect";
			hssi_8g_rx_pcs_gen3_clk_en                                             : string  := "disable_clk";
			hssi_8g_rx_pcs_gen3_rx_clk_sel                                         : string  := "rcvd_clk";
			hssi_8g_rx_pcs_gen3_tx_clk_sel                                         : string  := "tx_pma_clk";
			hssi_8g_rx_pcs_hip_mode                                                : string  := "dis_hip";
			hssi_8g_rx_pcs_ibm_invalid_code                                        : string  := "dis_ibm_invalid_code";
			hssi_8g_rx_pcs_invalid_code_flag_only                                  : string  := "dis_invalid_code_only";
			hssi_8g_rx_pcs_pad_or_edb_error_replace                                : string  := "replace_edb";
			hssi_8g_rx_pcs_pcs_bypass                                              : string  := "dis_pcs_bypass";
			hssi_8g_rx_pcs_phase_comp_rdptr                                        : string  := "enable_rdptr";
			hssi_8g_rx_pcs_phase_compensation_fifo                                 : string  := "low_latency";
			hssi_8g_rx_pcs_pipe_if_enable                                          : string  := "dis_pipe_rx";
			hssi_8g_rx_pcs_pma_dw                                                  : string  := "eight_bit";
			hssi_8g_rx_pcs_polinv_8b10b_dec                                        : string  := "dis_polinv_8b10b_dec";
			hssi_8g_rx_pcs_prot_mode                                               : string  := "gige";
			hssi_8g_rx_pcs_rate_match                                              : string  := "dis_rm";
			hssi_8g_rx_pcs_rate_match_del_thres                                    : string  := "dis_rm_del_thres";
			hssi_8g_rx_pcs_rate_match_empty_thres                                  : string  := "dis_rm_empty_thres";
			hssi_8g_rx_pcs_rate_match_full_thres                                   : string  := "dis_rm_full_thres";
			hssi_8g_rx_pcs_rate_match_ins_thres                                    : string  := "dis_rm_ins_thres";
			hssi_8g_rx_pcs_rate_match_start_thres                                  : string  := "dis_rm_start_thres";
			hssi_8g_rx_pcs_rx_clk_free_running                                     : string  := "en_rx_clk_free_run";
			hssi_8g_rx_pcs_rx_clk2                                                 : string  := "rcvd_clk_clk2";
			hssi_8g_rx_pcs_rx_pcs_urst                                             : string  := "en_rx_pcs_urst";
			hssi_8g_rx_pcs_rx_rcvd_clk                                             : string  := "rcvd_clk_rcvd_clk";
			hssi_8g_rx_pcs_rx_rd_clk                                               : string  := "pld_rx_clk";
			hssi_8g_rx_pcs_rx_refclk                                               : string  := "dis_refclk_sel";
			hssi_8g_rx_pcs_rx_wr_clk                                               : string  := "rx_clk2_div_1_2_4";
			hssi_8g_rx_pcs_sup_mode                                                : string  := "user_mode";
			hssi_8g_rx_pcs_symbol_swap                                             : string  := "dis_symbol_swap";
			hssi_8g_rx_pcs_sync_sm_idle_eios                                       : string  := "dis_syncsm_idle";
			hssi_8g_rx_pcs_test_bus_sel                                            : string  := "tx_testbus";
			hssi_8g_rx_pcs_tx_rx_parallel_loopback                                 : string  := "dis_plpbk";
			hssi_8g_rx_pcs_wa_boundary_lock_ctrl                                   : string  := "bit_slip";
			hssi_8g_rx_pcs_wa_clk_slip_spacing                                     : integer := 16;
			hssi_8g_rx_pcs_wa_det_latency_sync_status_beh                          : string  := "dont_care_assert_sync";
			hssi_8g_rx_pcs_wa_disp_err_flag                                        : string  := "dis_disp_err_flag";
			hssi_8g_rx_pcs_wa_kchar                                                : string  := "dis_kchar";
			hssi_8g_rx_pcs_wa_pd                                                   : string  := "wa_pd_10";
			hssi_8g_rx_pcs_wa_pd_data                                              : string  := "0";
			hssi_8g_rx_pcs_wa_pd_polarity                                          : string  := "dis_pd_both_pol";
			hssi_8g_rx_pcs_wa_pld_controlled                                       : string  := "dis_pld_ctrl";
			hssi_8g_rx_pcs_wa_renumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_rgnumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_rknumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_rosnumber_data                                       : integer := 0;
			hssi_8g_rx_pcs_wa_rvnumber_data                                        : integer := 0;
			hssi_8g_rx_pcs_wa_sync_sm_ctrl                                         : string  := "gige_sync_sm";
			hssi_8g_rx_pcs_wait_cnt                                                : integer := 0;
			hssi_8g_tx_pcs_bit_reversal                                            : string  := "dis_bit_reversal";
			hssi_8g_tx_pcs_bonding_dft_en                                          : string  := "dft_dis";
			hssi_8g_tx_pcs_bonding_dft_val                                         : string  := "dft_0";
			hssi_8g_tx_pcs_bypass_pipeline_reg                                     : string  := "dis_bypass_pipeline";
			hssi_8g_tx_pcs_byte_serializer                                         : string  := "dis_bs";
			hssi_8g_tx_pcs_clock_gate_bs_enc                                       : string  := "dis_bs_enc_clk_gating";
			hssi_8g_tx_pcs_clock_gate_dw_fifowr                                    : string  := "dis_dw_fifowr_clk_gating";
			hssi_8g_tx_pcs_clock_gate_fiford                                       : string  := "dis_fiford_clk_gating";
			hssi_8g_tx_pcs_clock_gate_sw_fifowr                                    : string  := "dis_sw_fifowr_clk_gating";
			hssi_8g_tx_pcs_clock_observation_in_pld_core                           : string  := "internal_refclk_b";
			hssi_8g_tx_pcs_data_selection_8b10b_encoder_input                      : string  := "normal_data_path";
			hssi_8g_tx_pcs_dynamic_clk_switch                                      : string  := "dis_dyn_clk_switch";
			hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                                   : string  := "dis_disp_ctrl";
			hssi_8g_tx_pcs_eightb_tenb_encoder                                     : string  := "dis_8b10b";
			hssi_8g_tx_pcs_force_echar                                             : string  := "dis_force_echar";
			hssi_8g_tx_pcs_force_kchar                                             : string  := "dis_force_kchar";
			hssi_8g_tx_pcs_gen3_tx_clk_sel                                         : string  := "tx_pma_clk";
			hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                                    : string  := "func_clk";
			hssi_8g_tx_pcs_hip_mode                                                : string  := "dis_hip";
			hssi_8g_tx_pcs_pcs_bypass                                              : string  := "dis_pcs_bypass";
			hssi_8g_tx_pcs_phase_comp_rdptr                                        : string  := "enable_rdptr";
			hssi_8g_tx_pcs_phase_compensation_fifo                                 : string  := "low_latency";
			hssi_8g_tx_pcs_phfifo_write_clk_sel                                    : string  := "pld_tx_clk";
			hssi_8g_tx_pcs_pma_dw                                                  : string  := "eight_bit";
			hssi_8g_tx_pcs_prot_mode                                               : string  := "basic";
			hssi_8g_tx_pcs_refclk_b_clk_sel                                        : string  := "tx_pma_clock";
			hssi_8g_tx_pcs_revloop_back_rm                                         : string  := "dis_rev_loopback_rx_rm";
			hssi_8g_tx_pcs_sup_mode                                                : string  := "user_mode";
			hssi_8g_tx_pcs_symbol_swap                                             : string  := "dis_symbol_swap";
			hssi_8g_tx_pcs_tx_bitslip                                              : string  := "dis_tx_bitslip";
			hssi_8g_tx_pcs_tx_compliance_controlled_disparity                      : string  := "dis_txcompliance";
			hssi_8g_tx_pcs_tx_fast_pld_reg                                         : string  := "dis_tx_fast_pld_reg";
			hssi_8g_tx_pcs_txclk_freerun                                           : string  := "dis_freerun_tx";
			hssi_8g_tx_pcs_txpcs_urst                                              : string  := "en_txpcs_urst";
			hssi_tx_pld_pcs_interface_hd_chnl_hip_en                               : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx                         : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx                : string  := "individual_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx                            : string  := "pma_8b_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx                     : string  := "fifo_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx                 : string  := "single_tx";
			hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx                    : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_func_mode                            : string  := "enable";
			hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en                              : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en                   : string  := "enable";
			hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz                        : integer := 0;
			hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz                        : integer := 0;
			hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz                  : integer := 0;
			hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx                         : string  := "teng_mode_tx";
			hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx                 : string  := "single_tx";
			hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode                : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_10g_lpbk_en                               : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx                 : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx                             : string  := "pma_64b_tx";
			hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx                          : string  := "fifo_tx";
			hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx                          : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx                     : string  := "enable";
			hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx                  : string  := "single_tx";
			hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode                 : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_8g_lpbk_en                                : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx                           : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_8g_hip_mode                               : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx                              : string  := "pma_8b_tx";
			hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx                           : string  := "fifo_tx";
			hssi_tx_pld_pcs_interface_hd_g3_prot_mode                              : string  := "disabled_prot_mode";
			hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en                             : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx                        : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx                   : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en                             : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode                            : string  := "disable";
			hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx                        : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx                           : string  := "pma_8b_tx";
			hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx                        : string  := "disabled_prot_mode_tx";
			hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        : string  := "disable";
			hssi_tx_pld_pcs_interface_pcs_tx_clk_source                            : string  := "teng";
			hssi_tx_pld_pcs_interface_pcs_tx_data_source                           : string  := "hip_disable";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en                         : string  := "delay1_clk_disable";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel                        : string  := "pld_tx_clk";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl                           : string  := "delay1_path0";
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel                       : string  := "one_ff_delay";
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en                         : string  := "delay2_clk_disable";
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl                           : string  := "delay2_path0";
			hssi_tx_pld_pcs_interface_pcs_tx_output_sel                            : string  := "teng_output";
			hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel                           : string  := "teng_clk_out";
			hssi_rx_pld_pcs_interface_hd_chnl_hip_en                               : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx                   : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx                         : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx                : string  := "individual_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx                            : string  := "pma_8b_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx                     : string  := "fifo_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx                 : string  := "single_rx";
			hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx                    : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_func_mode                            : string  := "enable";
			hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en                              : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx                 : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en                   : string  := "enable";
			hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz                        : integer := 0;
			hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz                        : integer := 0;
			hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz                          : integer := 0;
			hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz                        : integer := 0;
			hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode               : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx                         : string  := "teng_mode_rx";
			hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx                 : string  := "single_rx";
			hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode                : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_10g_lpbk_en                               : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx                             : string  := "pma_64b_rx";
			hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx                          : string  := "fifo_rx";
			hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx                          : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx                     : string  := "enable";
			hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx                  : string  := "single_rx";
			hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode                         : string  := "tx";
			hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode                 : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_8g_lpbk_en                                : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx                           : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_8g_hip_mode                               : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx                              : string  := "pma_8b_rx";
			hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx                           : string  := "fifo_rx";
			hssi_rx_pld_pcs_interface_hd_g3_prot_mode                              : string  := "disabled_prot_mode";
			hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en                             : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx                        : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx                   : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode                       : string  := "tx";
			hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en                             : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode              : string  := "tx_rx_pair_enabled";
			hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode                            : string  := "disable";
			hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx                        : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx                           : string  := "pma_8b_rx";
			hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx                        : string  := "disabled_prot_mode_rx";
			hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        : string  := "disable";
			hssi_rx_pld_pcs_interface_pcs_rx_block_sel                             : string  := "pcs_direct";
			hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                               : string  := "pld_rx_clk";
			hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en                            : string  := "hip_rx_enable";
			hssi_rx_pld_pcs_interface_pcs_rx_output_sel                            : string  := "teng_output";
			hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel                           : string  := "teng_clk_out";
			hssi_common_pld_pcs_interface_dft_clk_out_en                           : string  := "dft_clk_out_disable";
			hssi_common_pld_pcs_interface_dft_clk_out_sel                          : string  := "teng_rx_dft_clk";
			hssi_common_pld_pcs_interface_hrdrstctrl_en                            : string  := "hrst_dis";
			hssi_common_pld_pcs_interface_pcs_testbus_block_sel                    : string  := "pma_if";
			hssi_rx_pcs_pma_interface_block_sel                                    : string  := "eight_g_pcs";
			hssi_rx_pcs_pma_interface_channel_operation_mode                       : string  := "tx_rx_pair_enabled";
			hssi_rx_pcs_pma_interface_clkslip_sel                                  : string  := "pld";
			hssi_rx_pcs_pma_interface_lpbk_en                                      : string  := "disable";
			hssi_rx_pcs_pma_interface_master_clk_sel                               : string  := "master_rx_pma_clk";
			hssi_rx_pcs_pma_interface_pldif_datawidth_mode                         : string  := "pldif_data_10bit";
			hssi_rx_pcs_pma_interface_pma_dw_rx                                    : string  := "pma_8b_rx";
			hssi_rx_pcs_pma_interface_pma_if_dft_en                                : string  := "dft_dis";
			hssi_rx_pcs_pma_interface_pma_if_dft_val                               : string  := "dft_0";
			hssi_rx_pcs_pma_interface_prbs_clken                                   : string  := "prbs_clk_dis";
			hssi_rx_pcs_pma_interface_prbs_ver                                     : string  := "prbs_off";
			hssi_rx_pcs_pma_interface_prbs9_dwidth                                 : string  := "prbs9_64b";
			hssi_rx_pcs_pma_interface_prot_mode_rx                                 : string  := "disabled_prot_mode_rx";
			hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion                    : string  := "rx_dyn_polinv_dis";
			hssi_rx_pcs_pma_interface_rx_lpbk_en                                   : string  := "lpbk_dis";
			hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok                      : string  := "unforce_sig_ok";
			hssi_rx_pcs_pma_interface_rx_prbs_mask                                 : string  := "prbsmask128";
			hssi_rx_pcs_pma_interface_rx_prbs_mode                                 : string  := "teng_mode";
			hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel                    : string  := "sel_sig_det";
			hssi_rx_pcs_pma_interface_rx_static_polarity_inversion                 : string  := "rx_stat_polinv_dis";
			hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en                             : string  := "uhsif_lpbk_dis";
			hssi_rx_pcs_pma_interface_sup_mode                                     : string  := "user_mode";
			hssi_tx_pcs_pma_interface_bypass_pma_txelecidle                        : string  := "false";
			hssi_tx_pcs_pma_interface_channel_operation_mode                       : string  := "tx_rx_pair_enabled";
			hssi_tx_pcs_pma_interface_lpbk_en                                      : string  := "disable";
			hssi_tx_pcs_pma_interface_master_clk_sel                               : string  := "master_tx_pma_clk";
			hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx                        : string  := "other_prot_mode";
			hssi_tx_pcs_pma_interface_pldif_datawidth_mode                         : string  := "pldif_data_10bit";
			hssi_tx_pcs_pma_interface_pma_dw_tx                                    : string  := "pma_8b_tx";
			hssi_tx_pcs_pma_interface_pma_if_dft_en                                : string  := "dft_dis";
			hssi_tx_pcs_pma_interface_pmagate_en                                   : string  := "pmagate_dis";
			hssi_tx_pcs_pma_interface_prbs_clken                                   : string  := "prbs_clk_dis";
			hssi_tx_pcs_pma_interface_prbs_gen_pat                                 : string  := "prbs_gen_dis";
			hssi_tx_pcs_pma_interface_prbs9_dwidth                                 : string  := "prbs9_64b";
			hssi_tx_pcs_pma_interface_prot_mode_tx                                 : string  := "disabled_prot_mode_tx";
			hssi_tx_pcs_pma_interface_sq_wave_num                                  : string  := "sq_wave_4";
			hssi_tx_pcs_pma_interface_sqwgen_clken                                 : string  := "sqwgen_clk_dis";
			hssi_tx_pcs_pma_interface_sup_mode                                     : string  := "user_mode";
			hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion                    : string  := "tx_dyn_polinv_dis";
			hssi_tx_pcs_pma_interface_tx_pma_data_sel                              : string  := "pld_dir";
			hssi_tx_pcs_pma_interface_tx_static_polarity_inversion                 : string  := "tx_stat_polinv_dis";
			hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock              : string  := "uhsif_filt_stepsz_b4lock_4";
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value       : integer := 11;
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock            : string  := "uhsif_filt_cntthr_b4lock_16";
			hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period                 : string  := "uhsif_dcn_test_period_4";
			hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable                    : string  := "uhsif_dcn_test_mode_disable";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh                 : string  := "uhsif_dzt_cnt_thr_4";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable             : string  := "uhsif_dzt_enable";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window                 : string  := "uhsif_dzt_obr_win_32";
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size                    : string  := "uhsif_dzt_skipsz_8";
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel                   : string  := "uhsif_index_internal";
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin                      : string  := "uhsif_dcn_margin_4";
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value          : integer := 128;
			hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control                  : string  := "uhsif_dft_dz_det_val_0";
			hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control                    : string  := "uhsif_dft_up_val_0";
			hssi_tx_pcs_pma_interface_uhsif_enable                                 : string  := "uhsif_disable";
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock              : string  := "uhsif_lkd_segsz_aflock_2048";
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock             : string  := "uhsif_lkd_segsz_b4lock_32";
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value   : integer := 8;
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value  : integer := 8;
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value  : integer := 3;
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value : integer := 3;
			hssi_common_pcs_pma_interface_asn_clk_enable                           : string  := "false";
			hssi_common_pcs_pma_interface_asn_enable                               : string  := "dis_asn";
			hssi_common_pcs_pma_interface_block_sel                                : string  := "eight_g_pcs";
			hssi_common_pcs_pma_interface_bypass_early_eios                        : string  := "false";
			hssi_common_pcs_pma_interface_bypass_pcie_switch                       : string  := "false";
			hssi_common_pcs_pma_interface_bypass_pma_ltr                           : string  := "false";
			hssi_common_pcs_pma_interface_bypass_pma_sw_done                       : string  := "false";
			hssi_common_pcs_pma_interface_bypass_ppm_lock                          : string  := "false";
			hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp                   : string  := "false";
			hssi_common_pcs_pma_interface_bypass_txdetectrx                        : string  := "false";
			hssi_common_pcs_pma_interface_cdr_control                              : string  := "en_cdr_ctrl";
			hssi_common_pcs_pma_interface_cid_enable                               : string  := "en_cid_mode";
			hssi_common_pcs_pma_interface_data_mask_count                          : integer := 2500;
			hssi_common_pcs_pma_interface_data_mask_count_multi                    : integer := 1;
			hssi_common_pcs_pma_interface_dft_observation_clock_selection          : string  := "dft_clk_obsrv_tx0";
			hssi_common_pcs_pma_interface_early_eios_counter                       : integer := 50;
			hssi_common_pcs_pma_interface_force_freqdet                            : string  := "force_freqdet_dis";
			hssi_common_pcs_pma_interface_free_run_clk_enable                      : string  := "true";
			hssi_common_pcs_pma_interface_ignore_sigdet_g23                        : string  := "false";
			hssi_common_pcs_pma_interface_pc_en_counter                            : integer := 55;
			hssi_common_pcs_pma_interface_pc_rst_counter                           : integer := 23;
			hssi_common_pcs_pma_interface_pcie_hip_mode                            : string  := "hip_disable";
			hssi_common_pcs_pma_interface_ph_fifo_reg_mode                         : string  := "phfifo_reg_mode_dis";
			hssi_common_pcs_pma_interface_phfifo_flush_wait                        : integer := 36;
			hssi_common_pcs_pma_interface_pipe_if_g3pcs                            : string  := "pipe_if_8gpcs";
			hssi_common_pcs_pma_interface_pma_done_counter                         : integer := 175000;
			hssi_common_pcs_pma_interface_pma_if_dft_en                            : string  := "dft_dis";
			hssi_common_pcs_pma_interface_pma_if_dft_val                           : string  := "dft_0";
			hssi_common_pcs_pma_interface_ppm_cnt_rst                              : string  := "ppm_cnt_rst_dis";
			hssi_common_pcs_pma_interface_ppm_deassert_early                       : string  := "deassert_early_dis";
			hssi_common_pcs_pma_interface_ppm_gen1_2_cnt                           : string  := "cnt_32k";
			hssi_common_pcs_pma_interface_ppm_post_eidle_delay                     : string  := "cnt_200_cycles";
			hssi_common_pcs_pma_interface_ppmsel                                   : string  := "ppmsel_300";
			hssi_common_pcs_pma_interface_prot_mode                                : string  := "disable_prot_mode";
			hssi_common_pcs_pma_interface_rxvalid_mask                             : string  := "rxvalid_mask_en";
			hssi_common_pcs_pma_interface_sigdet_wait_counter                      : integer := 2500;
			hssi_common_pcs_pma_interface_sigdet_wait_counter_multi                : integer := 1;
			hssi_common_pcs_pma_interface_sim_mode                                 : string  := "disable";
			hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en                  : string  := "true";
			hssi_common_pcs_pma_interface_sup_mode                                 : string  := "user_mode";
			hssi_common_pcs_pma_interface_testout_sel                              : string  := "asn_test";
			hssi_common_pcs_pma_interface_wait_clk_on_off_timer                    : integer := 4;
			hssi_common_pcs_pma_interface_wait_pipe_synchronizing                  : integer := 23;
			hssi_common_pcs_pma_interface_wait_send_syncp_fbkp                     : integer := 250;
			hssi_common_pcs_pma_interface_ppm_det_buckets                          : string  := "ppm_100_bucket";
			hssi_fifo_rx_pcs_double_read_mode                                      : string  := "double_read_dis";
			hssi_fifo_rx_pcs_prot_mode                                             : string  := "teng_mode";
			hssi_fifo_tx_pcs_double_write_mode                                     : string  := "double_write_dis";
			hssi_fifo_tx_pcs_prot_mode                                             : string  := "teng_mode";
			hssi_pipe_gen3_bypass_rx_detection_enable                              : string  := "false";
			hssi_pipe_gen3_bypass_rx_preset                                        : integer := 0;
			hssi_pipe_gen3_bypass_rx_preset_enable                                 : string  := "false";
			hssi_pipe_gen3_bypass_tx_coefficent                                    : integer := 0;
			hssi_pipe_gen3_bypass_tx_coefficent_enable                             : string  := "false";
			hssi_pipe_gen3_elecidle_delay_g3                                       : integer := 6;
			hssi_pipe_gen3_ind_error_reporting                                     : string  := "dis_ind_error_reporting";
			hssi_pipe_gen3_mode                                                    : string  := "pipe_g1";
			hssi_pipe_gen3_phy_status_delay_g12                                    : integer := 5;
			hssi_pipe_gen3_phy_status_delay_g3                                     : integer := 5;
			hssi_pipe_gen3_phystatus_rst_toggle_g12                                : string  := "dis_phystatus_rst_toggle";
			hssi_pipe_gen3_phystatus_rst_toggle_g3                                 : string  := "dis_phystatus_rst_toggle_g3";
			hssi_pipe_gen3_rate_match_pad_insertion                                : string  := "dis_rm_fifo_pad_ins";
			hssi_pipe_gen3_sup_mode                                                : string  := "user_mode";
			hssi_pipe_gen3_test_out_sel                                            : string  := "disable_test_out";
			hssi_pipe_gen1_2_elec_idle_delay_val                                   : integer := 0;
			hssi_pipe_gen1_2_error_replace_pad                                     : string  := "replace_edb";
			hssi_pipe_gen1_2_hip_mode                                              : string  := "dis_hip";
			hssi_pipe_gen1_2_ind_error_reporting                                   : string  := "dis_ind_error_reporting";
			hssi_pipe_gen1_2_phystatus_delay_val                                   : integer := 0;
			hssi_pipe_gen1_2_phystatus_rst_toggle                                  : string  := "dis_phystatus_rst_toggle";
			hssi_pipe_gen1_2_pipe_byte_de_serializer_en                            : string  := "dont_care_bds";
			hssi_pipe_gen1_2_prot_mode                                             : string  := "pipe_g1";
			hssi_pipe_gen1_2_rx_pipe_enable                                        : string  := "dis_pipe_rx";
			hssi_pipe_gen1_2_rxdetect_bypass                                       : string  := "dis_rxdetect_bypass";
			hssi_pipe_gen1_2_sup_mode                                              : string  := "user_mode";
			hssi_pipe_gen1_2_tx_pipe_enable                                        : string  := "dis_pipe_tx";
			hssi_pipe_gen1_2_txswing                                               : string  := "dis_txswing";
			pma_adapt_adp_1s_ctle_bypass                                           : string  := "radp_1s_ctle_bypass_0";
			pma_adapt_adp_4s_ctle_bypass                                           : string  := "radp_4s_ctle_bypass_0";
			pma_adapt_adp_ctle_en                                                  : string  := "radp_ctle_disable";
			pma_adapt_adp_dfe_fltap_bypass                                         : string  := "radp_dfe_fltap_bypass_0";
			pma_adapt_adp_dfe_fltap_en                                             : string  := "radp_dfe_fltap_disable";
			pma_adapt_adp_dfe_fxtap_bypass                                         : string  := "radp_dfe_fxtap_bypass_0";
			pma_adapt_adp_dfe_fxtap_en                                             : string  := "radp_dfe_fxtap_disable";
			pma_adapt_adp_dfe_fxtap_hold_en                                        : string  := "radp_dfe_fxtap_not_held";
			pma_adapt_adp_dfe_mode                                                 : string  := "radp_dfe_mode_0";
			pma_adapt_adp_vga_bypass                                               : string  := "radp_vga_bypass_0";
			pma_adapt_adp_vga_en                                                   : string  := "radp_vga_disable";
			pma_adapt_adp_vref_bypass                                              : string  := "radp_vref_bypass_0";
			pma_adapt_adp_vref_en                                                  : string  := "radp_vref_disable";
			pma_adapt_datarate                                                     : string  := "0 bps";
			pma_adapt_prot_mode                                                    : string  := "basic_rx";
			pma_adapt_sup_mode                                                     : string  := "user_mode";
			pma_adapt_adp_ctle_adapt_cycle_window                                  : string  := "radp_ctle_adapt_cycle_window_6";
			pma_adapt_odi_dfe_spec_en                                              : string  := "rodi_dfe_spec_en_0";
			pma_adapt_adapt_mode                                                   : string  := "dfe_vga";
			pma_adapt_adp_onetime_dfe                                              : string  := "radp_onetime_dfe_0";
			pma_adapt_adp_mode                                                     : string  := "radp_mode_0";
			pma_cdr_refclk_powerdown_mode                                          : string  := "powerup";
			pma_cdr_refclk_refclk_select                                           : string  := "ref_iqclk0";
			pma_cgb_bitslip_enable                                                 : string  := "enable_bitslip";
			pma_cgb_bonding_reset_enable                                           : string  := "disallow_bonding_reset";
			pma_cgb_datarate                                                       : string  := "0 bps";
			pma_cgb_pcie_gen3_bitwidth                                             : string  := "pciegen3_wide";
			pma_cgb_prot_mode                                                      : string  := "basic_tx";
			pma_cgb_ser_mode                                                       : string  := "eight_bit";
			pma_cgb_sup_mode                                                       : string  := "user_mode";
			pma_cgb_x1_div_m_sel                                                   : string  := "divbypass";
			pma_cgb_input_select_x1                                                : string  := "fpll_bot";
			pma_cgb_input_select_gen3                                              : string  := "unused";
			pma_cgb_input_select_xn                                                : string  := "unused";
			pma_cgb_tx_ucontrol_en                                                 : string  := "disable";
			pma_rx_dfe_datarate                                                    : string  := "0 bps";
			pma_rx_dfe_dft_en                                                      : string  := "dft_disable";
			pma_rx_dfe_pdb                                                         : string  := "dfe_enable";
			pma_rx_dfe_pdb_fixedtap                                                : string  := "fixtap_dfe_powerdown";
			pma_rx_dfe_pdb_floattap                                                : string  := "floattap_dfe_powerdown";
			pma_rx_dfe_pdb_fxtap4t7                                                : string  := "fxtap4t7_powerdown";
			pma_rx_dfe_sup_mode                                                    : string  := "user_mode";
			pma_rx_dfe_prot_mode                                                   : string  := "basic_rx";
			pma_rx_odi_datarate                                                    : string  := "0 bps";
			pma_rx_odi_sup_mode                                                    : string  := "user_mode";
			pma_rx_odi_step_ctrl_sel                                               : string  := "feedback_mode";
			pma_rx_odi_prot_mode                                                   : string  := "basic_rx";
			pma_rx_buf_bypass_eqz_stages_234                                       : string  := "bypass_off";
			pma_rx_buf_datarate                                                    : string  := "0 bps";
			pma_rx_buf_diag_lp_en                                                  : string  := "dlp_off";
			pma_rx_buf_prot_mode                                                   : string  := "basic_rx";
			pma_rx_buf_qpi_enable                                                  : string  := "non_qpi_mode";
			pma_rx_buf_rx_refclk_divider                                           : string  := "bypass_divider";
			pma_rx_buf_sup_mode                                                    : string  := "user_mode";
			pma_rx_buf_loopback_modes                                              : string  := "lpbk_disable";
			pma_rx_buf_refclk_en                                                   : string  := "enable";
			pma_rx_buf_pm_tx_rx_pcie_gen                                           : string  := "non_pcie";
			pma_rx_buf_pm_tx_rx_pcie_gen_bitwidth                                  : string  := "pcie_gen3_32b";
			pma_rx_buf_pm_tx_rx_cvp_mode                                           : string  := "cvp_off";
			pma_rx_buf_xrx_path_uc_cal_enable                                      : string  := "rx_cal_off";
			pma_rx_buf_xrx_path_sup_mode                                           : string  := "user_mode";
			pma_rx_buf_xrx_path_prot_mode                                          : string  := "unused";
			pma_rx_buf_xrx_path_datarate                                           : string  := "0 bps";
			pma_rx_buf_xrx_path_datawidth                                          : integer := 0;
			pma_rx_buf_xrx_path_pma_rx_divclk_hz                                   : string  := "0";
			pma_rx_sd_prot_mode                                                    : string  := "basic_rx";
			pma_rx_sd_sd_output_off                                                : integer := 1;
			pma_rx_sd_sd_output_on                                                 : integer := 1;
			pma_rx_sd_sd_pdb                                                       : string  := "sd_off";
			pma_rx_sd_sup_mode                                                     : string  := "user_mode";
			pma_tx_ser_ser_clk_divtx_user_sel                                      : string  := "divtx_user_33";
			pma_tx_ser_sup_mode                                                    : string  := "user_mode";
			pma_tx_ser_prot_mode                                                   : string  := "basic_tx";
			pma_tx_buf_datarate                                                    : string  := "0 bps";
			pma_tx_buf_prot_mode                                                   : string  := "basic_tx";
			pma_tx_buf_rx_det                                                      : string  := "mode_0";
			pma_tx_buf_rx_det_output_sel                                           : string  := "rx_det_pcie_out";
			pma_tx_buf_rx_det_pdb                                                  : string  := "rx_det_off";
			pma_tx_buf_sup_mode                                                    : string  := "user_mode";
			pma_tx_buf_user_fir_coeff_ctrl_sel                                     : string  := "ram_ctl";
			pma_tx_buf_xtx_path_prot_mode                                          : string  := "basic_tx";
			pma_tx_buf_xtx_path_datarate                                           : string  := "0 bps";
			pma_tx_buf_xtx_path_datawidth                                          : integer := 0;
			pma_tx_buf_xtx_path_clock_divider_ratio                                : integer := 0;
			pma_tx_buf_xtx_path_pma_tx_divclk_hz                                   : string  := "0";
			pma_tx_buf_xtx_path_tx_pll_clk_hz                                      : string  := "0 hz";
			pma_tx_buf_xtx_path_sup_mode                                           : string  := "user_mode";
			cdr_pll_pma_width                                                      : integer := 8;
			cdr_pll_cgb_div                                                        : integer := 1;
			cdr_pll_is_cascaded_pll                                                : string  := "false";
			cdr_pll_datarate                                                       : string  := "0 bps";
			cdr_pll_lpd_counter                                                    : integer := 1;
			cdr_pll_lpfd_counter                                                   : integer := 1;
			cdr_pll_n_counter_scratch                                              : integer := 1;
			cdr_pll_output_clock_frequency                                         : string  := "0 hz";
			cdr_pll_reference_clock_frequency                                      : string  := "0 hz";
			cdr_pll_set_cdr_vco_speed                                              : integer := 1;
			cdr_pll_set_cdr_vco_speed_fix                                          : integer := 0;
			cdr_pll_vco_freq                                                       : string  := "0 hz";
			cdr_pll_atb_select_control                                             : string  := "atb_off";
			cdr_pll_auto_reset_on                                                  : string  := "auto_reset_on";
			cdr_pll_bbpd_data_pattern_filter_select                                : string  := "bbpd_data_pat_off";
			cdr_pll_bw_sel                                                         : string  := "low";
			cdr_pll_cdr_odi_select                                                 : string  := "sel_cdr";
			cdr_pll_cdr_phaselock_mode                                             : string  := "no_ignore_lock";
			cdr_pll_cdr_powerdown_mode                                             : string  := "power_up";
			cdr_pll_chgpmp_current_pd                                              : string  := "cp_current_pd_setting0";
			cdr_pll_chgpmp_current_pfd                                             : string  := "cp_current_pfd_setting0";
			cdr_pll_chgpmp_replicate                                               : string  := "false";
			cdr_pll_chgpmp_testmode                                                : string  := "cp_test_disable";
			cdr_pll_clklow_mux_select                                              : string  := "clklow_mux_cdr_fbclk";
			cdr_pll_diag_loopback_enable                                           : string  := "false";
			cdr_pll_disable_up_dn                                                  : string  := "true";
			cdr_pll_fref_clklow_div                                                : integer := 1;
			cdr_pll_fref_mux_select                                                : string  := "fref_mux_cdr_refclk";
			cdr_pll_gpon_lck2ref_control                                           : string  := "gpon_lck2ref_off";
			cdr_pll_initial_settings                                               : string  := "true";
			cdr_pll_lck2ref_delay_control                                          : string  := "lck2ref_delay_off";
			cdr_pll_lf_resistor_pd                                                 : string  := "lf_pd_setting0";
			cdr_pll_lf_resistor_pfd                                                : string  := "lf_pfd_setting0";
			cdr_pll_lf_ripple_cap                                                  : string  := "lf_no_ripple";
			cdr_pll_loop_filter_bias_select                                        : string  := "lpflt_bias_off";
			cdr_pll_loopback_mode                                                  : string  := "loopback_disabled";
			cdr_pll_ltd_ltr_micro_controller_select                                : string  := "ltd_ltr_pcs";
			cdr_pll_m_counter                                                      : integer := 1;
			cdr_pll_n_counter                                                      : integer := 1;
			cdr_pll_pd_fastlock_mode                                               : string  := "false";
			cdr_pll_pd_l_counter                                                   : integer := 1;
			cdr_pll_pfd_l_counter                                                  : integer := 1;
			cdr_pll_primary_use                                                    : string  := "cdr";
			cdr_pll_prot_mode                                                      : string  := "unused";
			cdr_pll_reverse_serial_loopback                                        : string  := "no_loopback";
			cdr_pll_set_cdr_v2i_enable                                             : string  := "true";
			cdr_pll_set_cdr_vco_reset                                              : string  := "false";
			cdr_pll_set_cdr_vco_speed_pciegen3                                     : string  := "cdr_vco_max_speedbin_pciegen3";
			cdr_pll_sup_mode                                                       : string  := "user_mode";
			cdr_pll_tx_pll_prot_mode                                               : string  := "txpll_unused";
			cdr_pll_txpll_hclk_driver_enable                                       : string  := "false";
			cdr_pll_vco_overrange_voltage                                          : string  := "vco_overrange_off";
			cdr_pll_vco_underrange_voltage                                         : string  := "vco_underange_off";
			cdr_pll_fb_select                                                      : string  := "direct_fb";
			cdr_pll_uc_ro_cal                                                      : string  := "uc_ro_cal_off";
			cdr_pll_iqclk_mux_sel                                                  : string  := "power_down";
			cdr_pll_pcie_gen                                                       : string  := "non_pcie";
			cdr_pll_set_cdr_input_freq_range                                       : integer := 0;
			cdr_pll_chgpmp_current_dn_trim                                         : string  := "cp_current_trimming_dn_setting0";
			cdr_pll_chgpmp_up_pd_trim_double                                       : string  := "normal_up_trim_current";
			cdr_pll_chgpmp_current_up_pd                                           : string  := "cp_current_pd_up_setting0";
			cdr_pll_chgpmp_current_up_trim                                         : string  := "cp_current_trimming_up_setting0";
			cdr_pll_chgpmp_dn_pd_trim_double                                       : string  := "normal_dn_trim_current";
			cdr_pll_cal_vco_count_length                                           : string  := "sel_8b_count";
			cdr_pll_chgpmp_current_dn_pd                                           : string  := "cp_current_pd_dn_setting0";
			pma_rx_deser_clkdiv_source                                             : string  := "vco_bypass_normal";
			pma_rx_deser_clkdivrx_user_mode                                        : string  := "clkdivrx_user_disabled";
			pma_rx_deser_datarate                                                  : string  := "0 bps";
			pma_rx_deser_deser_factor                                              : integer := 8;
			pma_rx_deser_force_clkdiv_for_testing                                  : string  := "normal_clkdiv";
			pma_rx_deser_sdclk_enable                                              : string  := "false";
			pma_rx_deser_sup_mode                                                  : string  := "user_mode";
			pma_rx_deser_rst_n_adapt_odi                                           : string  := "no_rst_adapt_odi";
			pma_rx_deser_bitslip_bypass                                            : string  := "bs_bypass_no";
			pma_rx_deser_prot_mode                                                 : string  := "basic_rx";
			pma_rx_deser_pcie_gen                                                  : string  := "non_pcie";
			pma_rx_deser_pcie_gen_bitwidth                                         : string  := "pcie_gen3_32b"
		);
		port (
			tx_analogreset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_analogreset
			tx_digitalreset           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_digitalreset
			rx_analogreset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_analogreset
			rx_digitalreset           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_digitalreset
			tx_cal_busy               : out std_logic_vector(3 downto 0);                      -- tx_cal_busy
			rx_cal_busy               : out std_logic_vector(3 downto 0);                      -- rx_cal_busy
			tx_serial_clk0            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			rx_cdr_refclk0            : in  std_logic                      := 'X';             -- clk
			tx_serial_data            : out std_logic_vector(3 downto 0);                      -- tx_serial_data
			rx_serial_data            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_serial_data
			rx_seriallpbken           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_seriallpbken
			rx_is_lockedtodata        : out std_logic_vector(3 downto 0);                      -- rx_is_lockedtodata
			tx_coreclkin              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			rx_coreclkin              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			tx_clkout                 : out std_logic_vector(3 downto 0);                      -- clk
			rx_clkout                 : out std_logic_vector(3 downto 0);                      -- clk
			tx_parallel_data          : in  std_logic_vector(511 downto 0) := (others => 'X'); -- unused_tx_parallel_data
			rx_parallel_data          : out std_logic_vector(511 downto 0);                    -- unused_rx_parallel_data
			rx_std_wa_patternalign    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_wa_patternalign
			tx_analogreset_ack        : out std_logic_vector(3 downto 0);                      -- tx_analogreset_ack
			rx_analogreset_ack        : out std_logic_vector(3 downto 0);                      -- rx_analogreset_ack
			tx_serial_clk1            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			tx_serial_clk2            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			tx_serial_clk3            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			tx_bonding_clocks         : in  std_logic_vector(23 downto 0)  := (others => 'X'); -- clk
			tx_bonding_clocks1        : in  std_logic_vector(23 downto 0)  := (others => 'X'); -- clk
			tx_bonding_clocks2        : in  std_logic_vector(23 downto 0)  := (others => 'X'); -- clk
			tx_bonding_clocks3        : in  std_logic_vector(23 downto 0)  := (others => 'X'); -- clk
			rx_cdr_refclk1            : in  std_logic                      := 'X';             -- clk
			rx_cdr_refclk2            : in  std_logic                      := 'X';             -- clk
			rx_cdr_refclk3            : in  std_logic                      := 'X';             -- clk
			rx_cdr_refclk4            : in  std_logic                      := 'X';             -- clk
			rx_pma_clkslip            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_pma_clkslip
			rx_set_locktodata         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_set_locktodata
			rx_set_locktoref          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_set_locktoref
			rx_is_lockedtoref         : out std_logic_vector(3 downto 0);                      -- rx_is_lockedtoref
			rx_pma_qpipulldn          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_pma_qpipulldn
			tx_pma_qpipulldn          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_pma_qpipulldn
			tx_pma_qpipullup          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_pma_qpipullup
			tx_pma_txdetectrx         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_pma_txdetectrx
			tx_pma_elecidle           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_pma_elecidle
			tx_pma_rxfound            : out std_logic_vector(3 downto 0);                      -- tx_pma_rxfound
			rx_clklow                 : out std_logic_vector(3 downto 0);                      -- rx_clklow
			rx_fref                   : out std_logic_vector(3 downto 0);                      -- rx_fref
			tx_pma_clkout             : out std_logic_vector(3 downto 0);                      -- clk
			tx_pma_div_clkout         : out std_logic_vector(3 downto 0);                      -- clk
			tx_pma_iqtxrx_clkout      : out std_logic_vector(3 downto 0);                      -- clk
			rx_pma_clkout             : out std_logic_vector(3 downto 0);                      -- clk
			rx_pma_div_clkout         : out std_logic_vector(3 downto 0);                      -- clk
			rx_pma_iqtxrx_clkout      : out std_logic_vector(3 downto 0);                      -- clk
			tx_control                : in  std_logic_vector(71 downto 0)  := (others => 'X'); -- tx_control
			rx_control                : out std_logic_vector(79 downto 0);                     -- rx_control
			rx_bitslip                : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_bitslip
			rx_adapt_reset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_adapt_reset
			rx_adapt_start            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_adapt_start
			rx_prbs_err_clr           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_prbs_err_clr
			rx_prbs_done              : out std_logic_vector(3 downto 0);                      -- rx_prbs_done
			rx_prbs_err               : out std_logic_vector(3 downto 0);                      -- rx_prbs_err
			tx_uhsif_clk              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			tx_uhsif_clkout           : out std_logic_vector(3 downto 0);                      -- clk
			tx_uhsif_lock             : out std_logic_vector(3 downto 0);                      -- tx_uhsif_lock
			tx_std_pcfifo_full        : out std_logic_vector(3 downto 0);                      -- tx_std_pcfifo_full
			tx_std_pcfifo_empty       : out std_logic_vector(3 downto 0);                      -- tx_std_pcfifo_empty
			rx_std_pcfifo_full        : out std_logic_vector(3 downto 0);                      -- rx_std_pcfifo_full
			rx_std_pcfifo_empty       : out std_logic_vector(3 downto 0);                      -- rx_std_pcfifo_empty
			rx_std_bitrev_ena         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_bitrev_ena
			rx_std_byterev_ena        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_byterev_ena
			tx_polinv                 : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_polinv
			rx_polinv                 : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_polinv
			tx_std_bitslipboundarysel : in  std_logic_vector(19 downto 0)  := (others => 'X'); -- tx_std_bitslipboundarysel
			rx_std_bitslipboundarysel : out std_logic_vector(19 downto 0);                     -- rx_std_bitslipboundarysel
			rx_std_wa_a1a2size        : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_std_wa_a1a2size
			rx_std_rmfifo_full        : out std_logic_vector(3 downto 0);                      -- rx_std_rmfifo_full
			rx_std_rmfifo_empty       : out std_logic_vector(3 downto 0);                      -- rx_std_rmfifo_empty
			rx_std_signaldetect       : out std_logic_vector(3 downto 0);                      -- rx_std_signaldetect
			tx_enh_data_valid         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_enh_data_valid
			tx_enh_fifo_full          : out std_logic_vector(3 downto 0);                      -- tx_enh_fifo_full
			tx_enh_fifo_pfull         : out std_logic_vector(3 downto 0);                      -- tx_enh_fifo_pfull
			tx_enh_fifo_empty         : out std_logic_vector(3 downto 0);                      -- tx_enh_fifo_empty
			tx_enh_fifo_pempty        : out std_logic_vector(3 downto 0);                      -- tx_enh_fifo_pempty
			tx_enh_fifo_cnt           : out std_logic_vector(15 downto 0);                     -- tx_enh_fifo_cnt
			rx_enh_fifo_rd_en         : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_enh_fifo_rd_en
			rx_enh_data_valid         : out std_logic_vector(3 downto 0);                      -- rx_enh_data_valid
			rx_enh_fifo_full          : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_full
			rx_enh_fifo_pfull         : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_pfull
			rx_enh_fifo_empty         : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_empty
			rx_enh_fifo_pempty        : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_pempty
			rx_enh_fifo_del           : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_del
			rx_enh_fifo_insert        : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_insert
			rx_enh_fifo_cnt           : out std_logic_vector(19 downto 0);                     -- rx_enh_fifo_cnt
			rx_enh_fifo_align_val     : out std_logic_vector(3 downto 0);                      -- rx_enh_fifo_align_val
			rx_enh_fifo_align_clr     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_enh_fifo_align_clr
			tx_enh_frame              : out std_logic_vector(3 downto 0);                      -- tx_enh_frame
			tx_enh_frame_burst_en     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- tx_enh_frame_burst_en
			tx_enh_frame_diag_status  : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- tx_enh_frame_diag_status
			rx_enh_frame              : out std_logic_vector(3 downto 0);                      -- rx_enh_frame
			rx_enh_frame_lock         : out std_logic_vector(3 downto 0);                      -- rx_enh_frame_lock
			rx_enh_frame_diag_status  : out std_logic_vector(7 downto 0);                      -- rx_enh_frame_diag_status
			rx_enh_crc32_err          : out std_logic_vector(3 downto 0);                      -- rx_enh_crc32err
			rx_enh_highber            : out std_logic_vector(3 downto 0);                      -- rx_enh_highber
			rx_enh_highber_clr_cnt    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_enh_highber_clr_cnt
			rx_enh_clr_errblk_count   : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- rx_enh_clr_errblk_count
			rx_enh_blk_lock           : out std_logic_vector(3 downto 0);                      -- rx_enh_blk_lock
			tx_enh_bitslip            : in  std_logic_vector(27 downto 0)  := (others => 'X'); -- tx_enh_bitslip
			tx_hip_data               : in  std_logic_vector(255 downto 0) := (others => 'X'); -- tx_hip_data
			rx_hip_data               : out std_logic_vector(203 downto 0);                    -- rx_hip_data
			hip_pipe_pclk             : out std_logic;                                         -- hip_pipe_pclk
			hip_fixedclk              : out std_logic;                                         -- hip_fixedclk
			hip_frefclk               : out std_logic_vector(3 downto 0);                      -- hip_frefclk
			hip_ctrl                  : out std_logic_vector(31 downto 0);                     -- hip_ctrl
			hip_cal_done              : out std_logic_vector(3 downto 0);                      -- hip_cal_done
			ltssm_detect_quiet        : in  std_logic                      := 'X';             -- ltssm_detect_quiet
			ltssm_detect_active       : in  std_logic                      := 'X';             -- ltssm_detect_active
			ltssm_rcvr_phase_two      : in  std_logic                      := 'X';             -- ltssm_rcvr_phase_two
			hip_reduce_counters       : in  std_logic                      := 'X';             -- hip_reduce_counters
			pcie_rate                 : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- pcie_rate
			pipe_rate                 : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- pipe_rate
			pipe_sw_done              : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- pipe_sw_done
			pipe_sw                   : out std_logic_vector(1 downto 0);                      -- pipe_sw
			pipe_hclk_in              : in  std_logic                      := 'X';             -- clk
			pipe_hclk_out             : out std_logic;                                         -- clk
			pipe_g3_txdeemph          : in  std_logic_vector(71 downto 0)  := (others => 'X'); -- pipe_g3_txdeemph
			pipe_g3_rxpresethint      : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- pipe_g3_rxpresethint
			pipe_rx_eidleinfersel     : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- pipe_rx_eidleinfersel
			pipe_rx_elecidle          : out std_logic_vector(3 downto 0);                      -- pipe_rx_elecidle
			pipe_rx_polarity          : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- pipe_rx_polarity
			reconfig_clk              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- clk
			reconfig_reset            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- reset
			reconfig_write            : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- write
			reconfig_read             : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- read
			reconfig_address          : in  std_logic_vector(39 downto 0)  := (others => 'X'); -- address
			reconfig_writedata        : in  std_logic_vector(127 downto 0) := (others => 'X'); -- writedata
			reconfig_readdata         : out std_logic_vector(127 downto 0);                    -- readdata
			reconfig_waitrequest      : out std_logic_vector(3 downto 0);                      -- waitrequest
			avmm_busy                 : out std_logic_vector(3 downto 0)                       -- avmm_busy
		);
	end component xcvr_8B10B_altera_xcvr_native_a10_181_b5mzony;

	component altera_xcvr_reset_control is
		generic (
			CHANNELS              : integer := 1;
			PLLS                  : integer := 1;
			SYS_CLK_IN_MHZ        : integer := 250;
			SYNCHRONIZE_RESET     : integer := 1;
			REDUCED_SIM_TIME      : integer := 1;
			TX_PLL_ENABLE         : integer := 1;
			T_PLL_POWERDOWN       : integer := 1000;
			SYNCHRONIZE_PLL_RESET : integer := 0;
			TX_ENABLE             : integer := 1;
			TX_PER_CHANNEL        : integer := 0;
			T_TX_ANALOGRESET      : integer := 0;
			T_TX_DIGITALRESET     : integer := 20;
			T_PLL_LOCK_HYST       : integer := 0;
			EN_PLL_CAL_BUSY       : integer := 0;
			RX_ENABLE             : integer := 1;
			RX_PER_CHANNEL        : integer := 0;
			T_RX_ANALOGRESET      : integer := 40;
			T_RX_DIGITALRESET     : integer := 4000
		);
		port (
			clock              : in  std_logic                    := 'X';             -- clk
			reset              : in  std_logic                    := 'X';             -- reset
			pll_powerdown      : out std_logic_vector(0 downto 0);                    -- pll_powerdown
			tx_analogreset     : out std_logic_vector(3 downto 0);                    -- tx_analogreset
			tx_digitalreset    : out std_logic_vector(3 downto 0);                    -- tx_digitalreset
			tx_ready           : out std_logic_vector(3 downto 0);                    -- tx_ready
			pll_locked         : in  std_logic_vector(0 downto 0) := (others => 'X'); -- pll_locked
			pll_select         : in  std_logic_vector(0 downto 0) := (others => 'X'); -- pll_select
			tx_cal_busy        : in  std_logic_vector(3 downto 0) := (others => 'X'); -- tx_cal_busy
			pll_cal_busy       : in  std_logic_vector(0 downto 0) := (others => 'X'); -- pll_cal_busy
			rx_analogreset     : out std_logic_vector(3 downto 0);                    -- rx_analogreset
			rx_digitalreset    : out std_logic_vector(3 downto 0);                    -- rx_digitalreset
			rx_ready           : out std_logic_vector(3 downto 0);                    -- rx_ready
			rx_is_lockedtodata : in  std_logic_vector(3 downto 0) := (others => 'X'); -- rx_is_lockedtodata
			rx_cal_busy        : in  std_logic_vector(3 downto 0) := (others => 'X'); -- rx_cal_busy
			tx_manual          : in  std_logic_vector(3 downto 0) := (others => 'X'); -- tx_reset_mode
			rx_manual          : in  std_logic_vector(3 downto 0) := (others => 'X'); -- rx_reset_mode
			tx_digitalreset_or : in  std_logic_vector(3 downto 0) := (others => 'X'); -- tx_digitalreset_or
			rx_digitalreset_or : in  std_logic_vector(3 downto 0) := (others => 'X')  -- rx_digitalreset_or
		);
	end component altera_xcvr_reset_control;

	signal xcvr_atx_pll_a10_0_pll_cal_busy_pll_cal_busy                : std_logic;                      -- xcvr_atx_pll_a10_0:pll_cal_busy -> xcvr_reset_control_0:pll_cal_busy0
	signal xcvr_atx_pll_a10_0_pll_locked_pll_locked                    : std_logic;                      -- xcvr_atx_pll_a10_0:pll_locked -> xcvr_reset_control_0:pll_locked0
	signal xcvr_reset_control_0_pll_powerdown0_pll_powerdown           : std_logic;                      -- xcvr_reset_control_0:pll_powerdown0 -> xcvr_atx_pll_a10_0:pll_powerdown
	signal xcvr_reset_control_0_rx_analogreset0_rx_analogreset         : std_logic;                      -- xcvr_reset_control_0:rx_analogreset0 -> xcvr_native_a10_0:rx_analogreset_ch0
	signal xcvr_reset_control_0_rx_analogreset1_rx_analogreset         : std_logic;                      -- xcvr_reset_control_0:rx_analogreset1 -> xcvr_native_a10_0:rx_analogreset_ch1
	signal xcvr_reset_control_0_rx_analogreset3_rx_analogreset         : std_logic;                      -- xcvr_reset_control_0:rx_analogreset3 -> xcvr_native_a10_0:rx_analogreset_ch3
	signal xcvr_reset_control_0_rx_analogreset2_rx_analogreset         : std_logic;                      -- xcvr_reset_control_0:rx_analogreset2 -> xcvr_native_a10_0:rx_analogreset_ch2
	signal xcvr_native_a10_0_rx_cal_busy_ch0_rx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:rx_cal_busy_ch0 -> xcvr_reset_control_0:rx_cal_busy0
	signal xcvr_native_a10_0_rx_cal_busy_ch2_rx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:rx_cal_busy_ch2 -> xcvr_reset_control_0:rx_cal_busy2
	signal xcvr_native_a10_0_rx_cal_busy_ch1_rx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:rx_cal_busy_ch1 -> xcvr_reset_control_0:rx_cal_busy1
	signal xcvr_native_a10_0_rx_cal_busy_ch3_rx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:rx_cal_busy_ch3 -> xcvr_reset_control_0:rx_cal_busy3
	signal xcvr_reset_control_0_rx_digitalreset0_rx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:rx_digitalreset0 -> xcvr_native_a10_0:rx_digitalreset_ch0
	signal xcvr_reset_control_0_rx_digitalreset2_rx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:rx_digitalreset2 -> xcvr_native_a10_0:rx_digitalreset_ch2
	signal xcvr_reset_control_0_rx_digitalreset1_rx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:rx_digitalreset1 -> xcvr_native_a10_0:rx_digitalreset_ch1
	signal xcvr_reset_control_0_rx_digitalreset3_rx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:rx_digitalreset3 -> xcvr_native_a10_0:rx_digitalreset_ch3
	signal xcvr_native_a10_0_rx_is_lockedtodata_ch1_rx_is_lockedtodata : std_logic;                      -- xcvr_native_a10_0:rx_is_lockedtodata_ch1 -> xcvr_reset_control_0:rx_is_lockedtodata1
	signal xcvr_native_a10_0_rx_is_lockedtodata_ch3_rx_is_lockedtodata : std_logic;                      -- xcvr_native_a10_0:rx_is_lockedtodata_ch3 -> xcvr_reset_control_0:rx_is_lockedtodata3
	signal xcvr_native_a10_0_rx_is_lockedtodata_ch0_rx_is_lockedtodata : std_logic;                      -- xcvr_native_a10_0:rx_is_lockedtodata_ch0 -> xcvr_reset_control_0:rx_is_lockedtodata0
	signal xcvr_native_a10_0_rx_is_lockedtodata_ch2_rx_is_lockedtodata : std_logic;                      -- xcvr_native_a10_0:rx_is_lockedtodata_ch2 -> xcvr_reset_control_0:rx_is_lockedtodata2
	signal xcvr_reset_control_0_tx_analogreset0_tx_analogreset         : std_logic;                      -- xcvr_reset_control_0:tx_analogreset0 -> xcvr_native_a10_0:tx_analogreset_ch0
	signal xcvr_reset_control_0_tx_analogreset2_tx_analogreset         : std_logic;                      -- xcvr_reset_control_0:tx_analogreset2 -> xcvr_native_a10_0:tx_analogreset_ch2
	signal xcvr_reset_control_0_tx_analogreset1_tx_analogreset         : std_logic;                      -- xcvr_reset_control_0:tx_analogreset1 -> xcvr_native_a10_0:tx_analogreset_ch1
	signal xcvr_reset_control_0_tx_analogreset3_tx_analogreset         : std_logic;                      -- xcvr_reset_control_0:tx_analogreset3 -> xcvr_native_a10_0:tx_analogreset_ch3
	signal xcvr_native_a10_0_tx_cal_busy_ch0_tx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:tx_cal_busy_ch0 -> xcvr_reset_control_0:tx_cal_busy0
	signal xcvr_native_a10_0_tx_cal_busy_ch2_tx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:tx_cal_busy_ch2 -> xcvr_reset_control_0:tx_cal_busy2
	signal xcvr_native_a10_0_tx_cal_busy_ch1_tx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:tx_cal_busy_ch1 -> xcvr_reset_control_0:tx_cal_busy1
	signal xcvr_native_a10_0_tx_cal_busy_ch3_tx_cal_busy               : std_logic;                      -- xcvr_native_a10_0:tx_cal_busy_ch3 -> xcvr_reset_control_0:tx_cal_busy3
	signal xcvr_reset_control_0_tx_digitalreset0_tx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:tx_digitalreset0 -> xcvr_native_a10_0:tx_digitalreset_ch0
	signal xcvr_reset_control_0_tx_digitalreset2_tx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:tx_digitalreset2 -> xcvr_native_a10_0:tx_digitalreset_ch2
	signal xcvr_reset_control_0_tx_digitalreset1_tx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:tx_digitalreset1 -> xcvr_native_a10_0:tx_digitalreset_ch1
	signal xcvr_reset_control_0_tx_digitalreset3_tx_digitalreset       : std_logic;                      -- xcvr_reset_control_0:tx_digitalreset3 -> xcvr_native_a10_0:tx_digitalreset_ch3
	signal xcvr_atx_pll_a10_0_tx_serial_clk_clk                        : std_logic;                      -- xcvr_atx_pll_a10_0:tx_serial_clk -> [xcvr_native_a10_0:tx_serial_clk0_ch0, xcvr_native_a10_0:tx_serial_clk0_ch1, xcvr_native_a10_0:tx_serial_clk0_ch2, xcvr_native_a10_0:tx_serial_clk0_ch3]
	signal xcvr_native_a10_0_tx_clkout                                 : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_native_a10_0_tx_serial_data                            : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_native_a10_0_rx_parallel_data                          : std_logic_vector(511 downto 0); -- port fragment
	signal xcvr_native_a10_0_rx_cal_busy                               : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_native_a10_0_rx_is_lockedtodata                        : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_native_a10_0_tx_cal_busy                               : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_native_a10_0_rx_clkout                                 : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_reset_control_0_pll_powerdown                          : std_logic_vector(0 downto 0);   -- port fragment
	signal xcvr_reset_control_0_rx_digitalreset                        : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_reset_control_0_tx_analogreset                         : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_reset_control_0_rx_ready                               : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_reset_control_0_tx_digitalreset                        : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_reset_control_0_rx_analogreset                         : std_logic_vector(3 downto 0);   -- port fragment
	signal xcvr_reset_control_0_tx_ready                               : std_logic_vector(3 downto 0);   -- port fragment

	for xcvr_atx_pll_a10_0 : xcvr_8B10B_altera_xcvr_atx_pll_a10_181_ubmonnq
		use entity xcvr_8B10B_altera_xcvr_atx_pll_a10_181.xcvr_8B10B_altera_xcvr_atx_pll_a10_181_ubmonnq;
	for xcvr_native_a10_0 : xcvr_8B10B_altera_xcvr_native_a10_181_b5mzony
		use entity xcvr_8B10B_altera_xcvr_native_a10_181.xcvr_8B10B_altera_xcvr_native_a10_181_b5mzony;
	for xcvr_reset_control_0 : altera_xcvr_reset_control
		use entity xcvr_8B10B_altera_xcvr_reset_control_181.altera_xcvr_reset_control;
begin

	xcvr_atx_pll_a10_0 : component xcvr_8B10B_altera_xcvr_atx_pll_a10_181_ubmonnq
		generic map (
			enable_pll_reconfig                                              => 0,
			rcfg_jtag_enable                                                 => 0,
			rcfg_separate_avmm_busy                                          => 0,
			dbg_embedded_debug_enable                                        => 0,
			dbg_capability_reg_enable                                        => 0,
			dbg_user_identifier                                              => 0,
			dbg_stat_soft_logic_enable                                       => 0,
			dbg_ctrl_soft_logic_enable                                       => 0,
			rcfg_emb_strm_enable                                             => 0,
			rcfg_profile_cnt                                                 => 2,
			hssi_pma_lc_refclk_select_mux_powerdown_mode                     => "powerup",
			hssi_pma_lc_refclk_select_mux_refclk_select                      => "ref_iqclk0",
			hssi_pma_lc_refclk_select_mux_silicon_rev                        => "20nm4",
			hssi_pma_lc_refclk_select_mux_inclk0_logical_to_physical_mapping => "ref_iqclk0",
			hssi_pma_lc_refclk_select_mux_inclk1_logical_to_physical_mapping => "power_down",
			hssi_pma_lc_refclk_select_mux_inclk2_logical_to_physical_mapping => "power_down",
			hssi_pma_lc_refclk_select_mux_inclk3_logical_to_physical_mapping => "power_down",
			hssi_pma_lc_refclk_select_mux_inclk4_logical_to_physical_mapping => "power_down",
			hssi_refclk_divider_silicon_rev                                  => "20nm4",
			atx_pll_silicon_rev                                              => "20nm4",
			atx_pll_is_cascaded_pll                                          => "false",
			atx_pll_cgb_div                                                  => 1,
			atx_pll_pma_width                                                => 64,
			atx_pll_cp_compensation_enable                                   => "true",
			atx_pll_cp_current_setting                                       => "cp_current_setting26",
			atx_pll_cp_testmode                                              => "cp_normal",
			atx_pll_cp_lf_3rd_pole_freq                                      => "lf_3rd_pole_setting1",
			atx_pll_lf_cbig_size                                             => "lf_cbig_setting4",
			atx_pll_cp_lf_order                                              => "lf_3rd_order",
			atx_pll_lf_resistance                                            => "lf_setting1",
			atx_pll_lf_ripplecap                                             => "lf_ripple_cap_0",
			atx_pll_tank_sel                                                 => "lctank1",
			atx_pll_tank_band                                                => "lc_band4",
			atx_pll_tank_voltage_coarse                                      => "vreg_setting_coarse0",
			atx_pll_tank_voltage_fine                                        => "vreg_setting5",
			atx_pll_output_regulator_supply                                  => "vreg1v_setting0",
			atx_pll_overrange_voltage                                        => "over_setting0",
			atx_pll_underrange_voltage                                       => "under_setting4",
			atx_pll_fb_select                                                => "direct_fb",
			atx_pll_d2a_voltage                                              => "d2a_setting_4",
			atx_pll_dsm_mode                                                 => "dsm_mode_integer",
			atx_pll_dsm_out_sel                                              => "pll_dsm_disable",
			atx_pll_dsm_ecn_bypass                                           => "false",
			atx_pll_dsm_ecn_test_en                                          => "false",
			atx_pll_dsm_fractional_division                                  => "1",
			atx_pll_dsm_fractional_value_ready                               => "pll_k_ready",
			atx_pll_iqclk_mux_sel                                            => "iqtxrxclk0",
			atx_pll_vco_bypass_enable                                        => "false",
			atx_pll_l_counter                                                => 8,
			atx_pll_l_counter_enable                                         => "true",
			atx_pll_cascadeclk_test                                          => "cascadetest_off",
			atx_pll_hclk_divide                                              => 1,
			atx_pll_enable_hclk                                              => "hclk_disabled",
			atx_pll_m_counter                                                => 40,
			atx_pll_ref_clk_div                                              => 1,
			atx_pll_bw_sel                                                   => "medium",
			atx_pll_datarate                                                 => "2540000000 bps",
			atx_pll_device_variant                                           => "device1",
			atx_pll_initial_settings                                         => "true",
			atx_pll_lc_mode                                                  => "lccmu_normal",
			atx_pll_output_clock_frequency                                   => "1270000000 Hz",
			atx_pll_powerdown_mode                                           => "powerup",
			atx_pll_prot_mode                                                => "basic_tx",
			atx_pll_reference_clock_frequency                                => "127000000 Hz",
			atx_pll_sup_mode                                                 => "user_mode",
			atx_pll_regulator_bypass                                         => "reg_enable",
			atx_pll_vco_freq                                                 => "10160000000 Hz",
			atx_pll_is_otn                                                   => "false",
			atx_pll_is_sdi                                                   => "false",
			atx_pll_primary_use                                              => "hssi_x1",
			atx_pll_fpll_refclk_selection                                    => "select_vco_output",
			atx_pll_lc_to_fpll_l_counter_scratch                             => 1,
			atx_pll_lc_to_fpll_l_counter                                     => "lcounter_setting0",
			atx_pll_pfd_delay_compensation                                   => "normal_delay",
			atx_pll_xcpvco_xchgpmplf_cp_current_boost                        => "normal_setting",
			atx_pll_pfd_pulse_width                                          => "pulse_width_setting0",
			hip_cal_en                                                       => "disable",
			calibration_en                                                   => "enable",
			enable_analog_resets                                             => 0,
			atx_pll_bonding_mode                                             => "cpri_bonding",
			enable_mcgb                                                      => 0,
			enable_mcgb_debug_ports_parameters                               => 0,
			hssi_pma_cgb_master_prot_mode                                    => "basic_tx",
			hssi_pma_cgb_master_silicon_rev                                  => "20nm4",
			hssi_pma_cgb_master_x1_div_m_sel                                 => "divbypass",
			hssi_pma_cgb_master_cgb_enable_iqtxrxclk                         => "disable_iqtxrxclk",
			hssi_pma_cgb_master_ser_mode                                     => "sixty_four_bit",
			hssi_pma_cgb_master_datarate                                     => "2540000000 bps",
			hssi_pma_cgb_master_cgb_power_down                               => "normal_cgb",
			hssi_pma_cgb_master_observe_cgb_clocks                           => "observe_nothing",
			hssi_pma_cgb_master_op_mode                                      => "enabled",
			hssi_pma_cgb_master_tx_ucontrol_reset_pcie                       => "pcscorehip_controls_mcgb",
			hssi_pma_cgb_master_vccdreg_output                               => "vccdreg_nominal",
			hssi_pma_cgb_master_input_select                                 => "lcpll_top",
			hssi_pma_cgb_master_input_select_gen3                            => "unused"
		)
		port map (
			pll_powerdown           => xcvr_reset_control_0_pll_powerdown0_pll_powerdown, -- pll_powerdown.pll_powerdown
			pll_refclk0             => clk_clk,                                           --   pll_refclk0.clk
			tx_serial_clk           => xcvr_atx_pll_a10_0_tx_serial_clk_clk,              -- tx_serial_clk.clk
			pll_locked              => xcvr_atx_pll_a10_0_pll_locked_pll_locked,          --    pll_locked.pll_locked
			pll_cal_busy            => xcvr_atx_pll_a10_0_pll_cal_busy_pll_cal_busy,      --  pll_cal_busy.pll_cal_busy
			pll_refclk1             => '0',                                               --   (terminated)
			pll_refclk2             => '0',                                               --   (terminated)
			pll_refclk3             => '0',                                               --   (terminated)
			pll_refclk4             => '0',                                               --   (terminated)
			tx_serial_clk_gt        => open,                                              --   (terminated)
			pll_pcie_clk            => open,                                              --   (terminated)
			pll_cascade_clk         => open,                                              --   (terminated)
			atx_to_fpll_cascade_clk => open,                                              --   (terminated)
			reconfig_clk0           => '0',                                               --   (terminated)
			reconfig_reset0         => '0',                                               --   (terminated)
			reconfig_write0         => '0',                                               --   (terminated)
			reconfig_read0          => '0',                                               --   (terminated)
			reconfig_address0       => "0000000000",                                      --   (terminated)
			reconfig_writedata0     => "00000000000000000000000000000000",                --   (terminated)
			reconfig_readdata0      => open,                                              --   (terminated)
			reconfig_waitrequest0   => open,                                              --   (terminated)
			avmm_busy0              => open,                                              --   (terminated)
			hip_cal_done            => open,                                              --   (terminated)
			clklow                  => open,                                              --   (terminated)
			fref                    => open,                                              --   (terminated)
			overrange               => open,                                              --   (terminated)
			underrange              => open,                                              --   (terminated)
			mcgb_rst                => '0',                                               --   (terminated)
			mcgb_aux_clk0           => '0',                                               --   (terminated)
			mcgb_aux_clk1           => '0',                                               --   (terminated)
			mcgb_aux_clk2           => '0',                                               --   (terminated)
			tx_bonding_clocks       => open,                                              --   (terminated)
			mcgb_serial_clk         => open,                                              --   (terminated)
			pcie_sw                 => "00",                                              --   (terminated)
			pcie_sw_done            => open,                                              --   (terminated)
			reconfig_clk1           => '0',                                               --   (terminated)
			reconfig_reset1         => '0',                                               --   (terminated)
			reconfig_write1         => '0',                                               --   (terminated)
			reconfig_read1          => '0',                                               --   (terminated)
			reconfig_address1       => "0000000000",                                      --   (terminated)
			reconfig_writedata1     => "00000000000000000000000000000000",                --   (terminated)
			reconfig_readdata1      => open,                                              --   (terminated)
			reconfig_waitrequest1   => open,                                              --   (terminated)
			mcgb_cal_busy           => open,                                              --   (terminated)
			mcgb_hip_cal_done       => open                                               --   (terminated)
		);

	xcvr_native_a10_0 : component xcvr_8B10B_altera_xcvr_native_a10_181_b5mzony
		generic map (
			device_revision                                                        => "20nm4",
			duplex_mode                                                            => "duplex",
			channels                                                               => 4,
			enable_calibration                                                     => 1,
			enable_analog_resets                                                   => 1,
			enable_reset_sequence                                                  => 1,
			bonded_mode                                                            => "not_bonded",
			pcs_bonding_master                                                     => 0,
			plls                                                                   => 1,
			number_physical_bonding_clocks                                         => 1,
			cdr_refclk_cnt                                                         => 1,
			enable_hip                                                             => 0,
			hip_cal_en                                                             => "disable",
			rcfg_enable                                                            => 0,
			rcfg_shared                                                            => 0,
			rcfg_jtag_enable                                                       => 0,
			rcfg_separate_avmm_busy                                                => 0,
			adme_prot_mode                                                         => "basic_std",
			adme_data_rate                                                         => "2540000000",
			enable_pcie_dfe_ip                                                     => false,
			sim_reduced_counters                                                   => false,
			disable_continuous_dfe                                                 => false,
			dbg_embedded_debug_enable                                              => 0,
			dbg_capability_reg_enable                                              => 0,
			dbg_user_identifier                                                    => 0,
			dbg_stat_soft_logic_enable                                             => 0,
			dbg_ctrl_soft_logic_enable                                             => 0,
			dbg_prbs_soft_logic_enable                                             => 0,
			dbg_odi_soft_logic_enable                                              => 0,
			rcfg_emb_strm_enable                                                   => 0,
			rcfg_profile_cnt                                                       => 2,
			hssi_gen3_rx_pcs_block_sync                                            => "bypass_block_sync",
			hssi_gen3_rx_pcs_block_sync_sm                                         => "disable_blk_sync_sm",
			hssi_gen3_rx_pcs_cdr_ctrl_force_unalgn                                 => "disable",
			hssi_gen3_rx_pcs_lpbk_force                                            => "lpbk_frce_dis",
			hssi_gen3_rx_pcs_mode                                                  => "disable_pcs",
			hssi_gen3_rx_pcs_rate_match_fifo                                       => "bypass_rm_fifo",
			hssi_gen3_rx_pcs_rate_match_fifo_latency                               => "low_latency",
			hssi_gen3_rx_pcs_reverse_lpbk                                          => "rev_lpbk_dis",
			hssi_gen3_rx_pcs_rx_b4gb_par_lpbk                                      => "b4gb_par_lpbk_dis",
			hssi_gen3_rx_pcs_rx_force_balign                                       => "dis_force_balign",
			hssi_gen3_rx_pcs_rx_ins_del_one_skip                                   => "ins_del_one_skip_dis",
			hssi_gen3_rx_pcs_rx_num_fixed_pat                                      => 0,
			hssi_gen3_rx_pcs_rx_test_out_sel                                       => "rx_test_out0",
			hssi_gen3_rx_pcs_sup_mode                                              => "user_mode",
			hssi_gen3_tx_pcs_mode                                                  => "disable_pcs",
			hssi_gen3_tx_pcs_reverse_lpbk                                          => "rev_lpbk_dis",
			hssi_gen3_tx_pcs_sup_mode                                              => "user_mode",
			hssi_gen3_tx_pcs_tx_bitslip                                            => 0,
			hssi_gen3_tx_pcs_tx_gbox_byp                                           => "bypass_gbox",
			hssi_krfec_rx_pcs_blksync_cor_en                                       => "detect",
			hssi_krfec_rx_pcs_bypass_gb                                            => "bypass_dis",
			hssi_krfec_rx_pcs_clr_ctrl                                             => "both_enabled",
			hssi_krfec_rx_pcs_ctrl_bit_reverse                                     => "ctrl_bit_reverse_en",
			hssi_krfec_rx_pcs_data_bit_reverse                                     => "data_bit_reverse_dis",
			hssi_krfec_rx_pcs_dv_start                                             => "with_blklock",
			hssi_krfec_rx_pcs_err_mark_type                                        => "err_mark_10g",
			hssi_krfec_rx_pcs_error_marking_en                                     => "err_mark_dis",
			hssi_krfec_rx_pcs_low_latency_en                                       => "disable",
			hssi_krfec_rx_pcs_lpbk_mode                                            => "lpbk_dis",
			hssi_krfec_rx_pcs_parity_invalid_enum                                  => 8,
			hssi_krfec_rx_pcs_parity_valid_num                                     => 4,
			hssi_krfec_rx_pcs_pipeln_blksync                                       => "enable",
			hssi_krfec_rx_pcs_pipeln_descrm                                        => "disable",
			hssi_krfec_rx_pcs_pipeln_errcorrect                                    => "disable",
			hssi_krfec_rx_pcs_pipeln_errtrap_ind                                   => "enable",
			hssi_krfec_rx_pcs_pipeln_errtrap_lfsr                                  => "disable",
			hssi_krfec_rx_pcs_pipeln_errtrap_loc                                   => "disable",
			hssi_krfec_rx_pcs_pipeln_errtrap_pat                                   => "disable",
			hssi_krfec_rx_pcs_pipeln_gearbox                                       => "enable",
			hssi_krfec_rx_pcs_pipeln_syndrm                                        => "enable",
			hssi_krfec_rx_pcs_pipeln_trans_dec                                     => "disable",
			hssi_krfec_rx_pcs_prot_mode                                            => "disable_mode",
			hssi_krfec_rx_pcs_receive_order                                        => "receive_lsb",
			hssi_krfec_rx_pcs_rx_testbus_sel                                       => "overall",
			hssi_krfec_rx_pcs_signal_ok_en                                         => "sig_ok_en",
			hssi_krfec_rx_pcs_sup_mode                                             => "user_mode",
			hssi_krfec_tx_pcs_burst_err                                            => "burst_err_dis",
			hssi_krfec_tx_pcs_burst_err_len                                        => "burst_err_len1",
			hssi_krfec_tx_pcs_ctrl_bit_reverse                                     => "ctrl_bit_reverse_en",
			hssi_krfec_tx_pcs_data_bit_reverse                                     => "data_bit_reverse_dis",
			hssi_krfec_tx_pcs_enc_frame_query                                      => "enc_query_dis",
			hssi_krfec_tx_pcs_low_latency_en                                       => "disable",
			hssi_krfec_tx_pcs_pipeln_encoder                                       => "enable",
			hssi_krfec_tx_pcs_pipeln_scrambler                                     => "enable",
			hssi_krfec_tx_pcs_prot_mode                                            => "disable_mode",
			hssi_krfec_tx_pcs_sup_mode                                             => "user_mode",
			hssi_krfec_tx_pcs_transcode_err                                        => "trans_err_dis",
			hssi_krfec_tx_pcs_transmit_order                                       => "transmit_lsb",
			hssi_krfec_tx_pcs_tx_testbus_sel                                       => "overall",
			hssi_10g_rx_pcs_align_del                                              => "align_del_dis",
			hssi_10g_rx_pcs_ber_bit_err_total_cnt                                  => "bit_err_total_cnt_10g",
			hssi_10g_rx_pcs_ber_clken                                              => "ber_clk_dis",
			hssi_10g_rx_pcs_ber_xus_timer_window                                   => 19530,
			hssi_10g_rx_pcs_bitslip_mode                                           => "bitslip_dis",
			hssi_10g_rx_pcs_blksync_bitslip_type                                   => "bitslip_comb",
			hssi_10g_rx_pcs_blksync_bitslip_wait_cnt                               => 1,
			hssi_10g_rx_pcs_blksync_bitslip_wait_type                              => "bitslip_cnt",
			hssi_10g_rx_pcs_blksync_bypass                                         => "blksync_bypass_en",
			hssi_10g_rx_pcs_blksync_clken                                          => "blksync_clk_dis",
			hssi_10g_rx_pcs_blksync_enum_invalid_sh_cnt                            => "enum_invalid_sh_cnt_10g",
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_postlock                           => "knum_sh_cnt_postlock_10g",
			hssi_10g_rx_pcs_blksync_knum_sh_cnt_prelock                            => "knum_sh_cnt_prelock_10g",
			hssi_10g_rx_pcs_blksync_pipeln                                         => "blksync_pipeln_dis",
			hssi_10g_rx_pcs_clr_errblk_cnt_en                                      => "disable",
			hssi_10g_rx_pcs_control_del                                            => "control_del_none",
			hssi_10g_rx_pcs_crcchk_bypass                                          => "crcchk_bypass_en",
			hssi_10g_rx_pcs_crcchk_clken                                           => "crcchk_clk_dis",
			hssi_10g_rx_pcs_crcchk_inv                                             => "crcchk_inv_en",
			hssi_10g_rx_pcs_crcchk_pipeln                                          => "crcchk_pipeln_en",
			hssi_10g_rx_pcs_crcflag_pipeln                                         => "crcflag_pipeln_en",
			hssi_10g_rx_pcs_ctrl_bit_reverse                                       => "ctrl_bit_reverse_dis",
			hssi_10g_rx_pcs_data_bit_reverse                                       => "data_bit_reverse_dis",
			hssi_10g_rx_pcs_dec_64b66b_rxsm_bypass                                 => "dec_64b66b_rxsm_bypass_en",
			hssi_10g_rx_pcs_dec64b66b_clken                                        => "dec64b66b_clk_dis",
			hssi_10g_rx_pcs_descrm_bypass                                          => "descrm_bypass_en",
			hssi_10g_rx_pcs_descrm_clken                                           => "descrm_clk_dis",
			hssi_10g_rx_pcs_descrm_mode                                            => "async",
			hssi_10g_rx_pcs_descrm_pipeln                                          => "enable",
			hssi_10g_rx_pcs_dft_clk_out_sel                                        => "rx_master_clk",
			hssi_10g_rx_pcs_dis_signal_ok                                          => "dis_signal_ok_en",
			hssi_10g_rx_pcs_dispchk_bypass                                         => "dispchk_bypass_en",
			hssi_10g_rx_pcs_empty_flag_type                                        => "empty_rd_side",
			hssi_10g_rx_pcs_fast_path                                              => "fast_path_en",
			hssi_10g_rx_pcs_fec_clken                                              => "fec_clk_dis",
			hssi_10g_rx_pcs_fec_enable                                             => "fec_dis",
			hssi_10g_rx_pcs_fifo_double_read                                       => "fifo_double_read_dis",
			hssi_10g_rx_pcs_fifo_stop_rd                                           => "n_rd_empty",
			hssi_10g_rx_pcs_fifo_stop_wr                                           => "n_wr_full",
			hssi_10g_rx_pcs_force_align                                            => "force_align_dis",
			hssi_10g_rx_pcs_frmsync_bypass                                         => "frmsync_bypass_en",
			hssi_10g_rx_pcs_frmsync_clken                                          => "frmsync_clk_dis",
			hssi_10g_rx_pcs_frmsync_enum_scrm                                      => "enum_scrm_default",
			hssi_10g_rx_pcs_frmsync_enum_sync                                      => "enum_sync_default",
			hssi_10g_rx_pcs_frmsync_flag_type                                      => "location_only",
			hssi_10g_rx_pcs_frmsync_knum_sync                                      => "knum_sync_default",
			hssi_10g_rx_pcs_frmsync_mfrm_length                                    => 2048,
			hssi_10g_rx_pcs_frmsync_pipeln                                         => "frmsync_pipeln_en",
			hssi_10g_rx_pcs_full_flag_type                                         => "full_wr_side",
			hssi_10g_rx_pcs_gb_rx_idwidth                                          => "width_64",
			hssi_10g_rx_pcs_gb_rx_odwidth                                          => "width_64",
			hssi_10g_rx_pcs_gbexp_clken                                            => "gbexp_clk_dis",
			hssi_10g_rx_pcs_low_latency_en                                         => "disable",
			hssi_10g_rx_pcs_lpbk_mode                                              => "lpbk_dis",
			hssi_10g_rx_pcs_master_clk_sel                                         => "master_rx_pma_clk",
			hssi_10g_rx_pcs_pempty_flag_type                                       => "pempty_rd_side",
			hssi_10g_rx_pcs_pfull_flag_type                                        => "pfull_wr_side",
			hssi_10g_rx_pcs_phcomp_rd_del                                          => "phcomp_rd_del2",
			hssi_10g_rx_pcs_pld_if_type                                            => "fifo",
			hssi_10g_rx_pcs_prot_mode                                              => "disable_mode",
			hssi_10g_rx_pcs_rand_clken                                             => "rand_clk_dis",
			hssi_10g_rx_pcs_rd_clk_sel                                             => "rd_rx_pld_clk",
			hssi_10g_rx_pcs_rdfifo_clken                                           => "rdfifo_clk_dis",
			hssi_10g_rx_pcs_rx_fifo_write_ctrl                                     => "blklock_stops",
			hssi_10g_rx_pcs_rx_scrm_width                                          => "bit64",
			hssi_10g_rx_pcs_rx_sh_location                                         => "msb",
			hssi_10g_rx_pcs_rx_signal_ok_sel                                       => "synchronized_ver",
			hssi_10g_rx_pcs_rx_sm_bypass                                           => "rx_sm_bypass_en",
			hssi_10g_rx_pcs_rx_sm_hiber                                            => "rx_sm_hiber_en",
			hssi_10g_rx_pcs_rx_sm_pipeln                                           => "rx_sm_pipeln_en",
			hssi_10g_rx_pcs_rx_testbus_sel                                         => "rx_fifo_testbus1",
			hssi_10g_rx_pcs_rx_true_b2b                                            => "b2b",
			hssi_10g_rx_pcs_rxfifo_empty                                           => "empty_default",
			hssi_10g_rx_pcs_rxfifo_full                                            => "full_default",
			hssi_10g_rx_pcs_rxfifo_mode                                            => "phase_comp",
			hssi_10g_rx_pcs_rxfifo_pempty                                          => 2,
			hssi_10g_rx_pcs_rxfifo_pfull                                           => 23,
			hssi_10g_rx_pcs_stretch_num_stages                                     => "zero_stage",
			hssi_10g_rx_pcs_sup_mode                                               => "user_mode",
			hssi_10g_rx_pcs_test_mode                                              => "test_off",
			hssi_10g_rx_pcs_wrfifo_clken                                           => "wrfifo_clk_dis",
			hssi_10g_rx_pcs_advanced_user_mode                                     => "disable",
			hssi_10g_tx_pcs_bitslip_en                                             => "bitslip_dis",
			hssi_10g_tx_pcs_bonding_dft_en                                         => "dft_dis",
			hssi_10g_tx_pcs_bonding_dft_val                                        => "dft_0",
			hssi_10g_tx_pcs_crcgen_bypass                                          => "crcgen_bypass_en",
			hssi_10g_tx_pcs_crcgen_clken                                           => "crcgen_clk_dis",
			hssi_10g_tx_pcs_crcgen_err                                             => "crcgen_err_dis",
			hssi_10g_tx_pcs_crcgen_inv                                             => "crcgen_inv_en",
			hssi_10g_tx_pcs_ctrl_bit_reverse                                       => "ctrl_bit_reverse_dis",
			hssi_10g_tx_pcs_data_bit_reverse                                       => "data_bit_reverse_dis",
			hssi_10g_tx_pcs_dft_clk_out_sel                                        => "tx_master_clk",
			hssi_10g_tx_pcs_dispgen_bypass                                         => "dispgen_bypass_en",
			hssi_10g_tx_pcs_dispgen_clken                                          => "dispgen_clk_dis",
			hssi_10g_tx_pcs_dispgen_err                                            => "dispgen_err_dis",
			hssi_10g_tx_pcs_dispgen_pipeln                                         => "dispgen_pipeln_dis",
			hssi_10g_tx_pcs_empty_flag_type                                        => "empty_rd_side",
			hssi_10g_tx_pcs_enc_64b66b_txsm_bypass                                 => "enc_64b66b_txsm_bypass_en",
			hssi_10g_tx_pcs_enc64b66b_txsm_clken                                   => "enc64b66b_txsm_clk_dis",
			hssi_10g_tx_pcs_fastpath                                               => "fastpath_en",
			hssi_10g_tx_pcs_fec_clken                                              => "fec_clk_dis",
			hssi_10g_tx_pcs_fec_enable                                             => "fec_dis",
			hssi_10g_tx_pcs_fifo_double_write                                      => "fifo_double_write_dis",
			hssi_10g_tx_pcs_fifo_reg_fast                                          => "fifo_reg_fast_dis",
			hssi_10g_tx_pcs_fifo_stop_rd                                           => "rd_empty",
			hssi_10g_tx_pcs_fifo_stop_wr                                           => "n_wr_full",
			hssi_10g_tx_pcs_frmgen_burst                                           => "frmgen_burst_dis",
			hssi_10g_tx_pcs_frmgen_bypass                                          => "frmgen_bypass_en",
			hssi_10g_tx_pcs_frmgen_clken                                           => "frmgen_clk_dis",
			hssi_10g_tx_pcs_frmgen_mfrm_length                                     => 2048,
			hssi_10g_tx_pcs_frmgen_pipeln                                          => "frmgen_pipeln_en",
			hssi_10g_tx_pcs_frmgen_pyld_ins                                        => "frmgen_pyld_ins_dis",
			hssi_10g_tx_pcs_frmgen_wordslip                                        => "frmgen_wordslip_dis",
			hssi_10g_tx_pcs_full_flag_type                                         => "full_wr_side",
			hssi_10g_tx_pcs_gb_pipeln_bypass                                       => "disable",
			hssi_10g_tx_pcs_gb_tx_idwidth                                          => "width_64",
			hssi_10g_tx_pcs_gb_tx_odwidth                                          => "width_64",
			hssi_10g_tx_pcs_gbred_clken                                            => "gbred_clk_dis",
			hssi_10g_tx_pcs_low_latency_en                                         => "disable",
			hssi_10g_tx_pcs_master_clk_sel                                         => "master_tx_pma_clk",
			hssi_10g_tx_pcs_pempty_flag_type                                       => "pempty_rd_side",
			hssi_10g_tx_pcs_pfull_flag_type                                        => "pfull_wr_side",
			hssi_10g_tx_pcs_phcomp_rd_del                                          => "phcomp_rd_del2",
			hssi_10g_tx_pcs_pld_if_type                                            => "fifo",
			hssi_10g_tx_pcs_prot_mode                                              => "disable_mode",
			hssi_10g_tx_pcs_pseudo_random                                          => "all_0",
			hssi_10g_tx_pcs_pseudo_seed_a                                          => "288230376151711743",
			hssi_10g_tx_pcs_pseudo_seed_b                                          => "288230376151711743",
			hssi_10g_tx_pcs_random_disp                                            => "disable",
			hssi_10g_tx_pcs_rdfifo_clken                                           => "rdfifo_clk_dis",
			hssi_10g_tx_pcs_scrm_bypass                                            => "scrm_bypass_en",
			hssi_10g_tx_pcs_scrm_clken                                             => "scrm_clk_dis",
			hssi_10g_tx_pcs_scrm_mode                                              => "async",
			hssi_10g_tx_pcs_scrm_pipeln                                            => "enable",
			hssi_10g_tx_pcs_sh_err                                                 => "sh_err_dis",
			hssi_10g_tx_pcs_sop_mark                                               => "sop_mark_dis",
			hssi_10g_tx_pcs_stretch_num_stages                                     => "zero_stage",
			hssi_10g_tx_pcs_sup_mode                                               => "user_mode",
			hssi_10g_tx_pcs_test_mode                                              => "test_off",
			hssi_10g_tx_pcs_tx_scrm_err                                            => "scrm_err_dis",
			hssi_10g_tx_pcs_tx_scrm_width                                          => "bit64",
			hssi_10g_tx_pcs_tx_sh_location                                         => "msb",
			hssi_10g_tx_pcs_tx_sm_bypass                                           => "tx_sm_bypass_en",
			hssi_10g_tx_pcs_tx_sm_pipeln                                           => "tx_sm_pipeln_en",
			hssi_10g_tx_pcs_tx_testbus_sel                                         => "tx_fifo_testbus1",
			hssi_10g_tx_pcs_txfifo_empty                                           => "empty_default",
			hssi_10g_tx_pcs_txfifo_full                                            => "full_default",
			hssi_10g_tx_pcs_txfifo_mode                                            => "phase_comp",
			hssi_10g_tx_pcs_txfifo_pempty                                          => 2,
			hssi_10g_tx_pcs_txfifo_pfull                                           => 11,
			hssi_10g_tx_pcs_wr_clk_sel                                             => "wr_tx_pld_clk",
			hssi_10g_tx_pcs_wrfifo_clken                                           => "wrfifo_clk_dis",
			hssi_10g_tx_pcs_advanced_user_mode                                     => "disable",
			hssi_8g_rx_pcs_auto_error_replacement                                  => "dis_err_replace",
			hssi_8g_rx_pcs_bit_reversal                                            => "dis_bit_reversal",
			hssi_8g_rx_pcs_bonding_dft_en                                          => "dft_dis",
			hssi_8g_rx_pcs_bonding_dft_val                                         => "dft_0",
			hssi_8g_rx_pcs_bypass_pipeline_reg                                     => "dis_bypass_pipeline",
			hssi_8g_rx_pcs_byte_deserializer                                       => "dis_bds",
			hssi_8g_rx_pcs_cdr_ctrl_rxvalid_mask                                   => "dis_rxvalid_mask",
			hssi_8g_rx_pcs_clkcmp_pattern_n                                        => 0,
			hssi_8g_rx_pcs_clkcmp_pattern_p                                        => 0,
			hssi_8g_rx_pcs_clock_gate_bds_dec_asn                                  => "dis_bds_dec_asn_clk_gating",
			hssi_8g_rx_pcs_clock_gate_cdr_eidle                                    => "en_cdr_eidle_clk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_pc_wrclk                                  => "dis_dw_pc_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_rm_rd                                     => "en_dw_rm_rdclk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_rm_wr                                     => "en_dw_rm_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_dw_wa                                        => "dis_dw_wa_clk_gating",
			hssi_8g_rx_pcs_clock_gate_pc_rdclk                                     => "dis_pc_rdclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_pc_wrclk                                  => "dis_sw_pc_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_rm_rd                                     => "en_sw_rm_rdclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_rm_wr                                     => "en_sw_rm_wrclk_gating",
			hssi_8g_rx_pcs_clock_gate_sw_wa                                        => "dis_sw_wa_clk_gating",
			hssi_8g_rx_pcs_clock_observation_in_pld_core                           => "internal_sw_wa_clk",
			hssi_8g_rx_pcs_eidle_entry_eios                                        => "dis_eidle_eios",
			hssi_8g_rx_pcs_eidle_entry_iei                                         => "dis_eidle_iei",
			hssi_8g_rx_pcs_eidle_entry_sd                                          => "dis_eidle_sd",
			hssi_8g_rx_pcs_eightb_tenb_decoder                                     => "dis_8b10b",
			hssi_8g_rx_pcs_err_flags_sel                                           => "err_flags_wa",
			hssi_8g_rx_pcs_fixed_pat_det                                           => "dis_fixed_patdet",
			hssi_8g_rx_pcs_fixed_pat_num                                           => 0,
			hssi_8g_rx_pcs_force_signal_detect                                     => "en_force_signal_detect",
			hssi_8g_rx_pcs_gen3_clk_en                                             => "disable_clk",
			hssi_8g_rx_pcs_gen3_rx_clk_sel                                         => "rcvd_clk",
			hssi_8g_rx_pcs_gen3_tx_clk_sel                                         => "tx_pma_clk",
			hssi_8g_rx_pcs_hip_mode                                                => "dis_hip",
			hssi_8g_rx_pcs_ibm_invalid_code                                        => "dis_ibm_invalid_code",
			hssi_8g_rx_pcs_invalid_code_flag_only                                  => "dis_invalid_code_only",
			hssi_8g_rx_pcs_pad_or_edb_error_replace                                => "replace_edb",
			hssi_8g_rx_pcs_pcs_bypass                                              => "dis_pcs_bypass",
			hssi_8g_rx_pcs_phase_comp_rdptr                                        => "enable_rdptr",
			hssi_8g_rx_pcs_phase_compensation_fifo                                 => "low_latency",
			hssi_8g_rx_pcs_pipe_if_enable                                          => "dis_pipe_rx",
			hssi_8g_rx_pcs_pma_dw                                                  => "twenty_bit",
			hssi_8g_rx_pcs_polinv_8b10b_dec                                        => "dis_polinv_8b10b_dec",
			hssi_8g_rx_pcs_prot_mode                                               => "basic_rm_disable",
			hssi_8g_rx_pcs_rate_match                                              => "dis_rm",
			hssi_8g_rx_pcs_rate_match_del_thres                                    => "dis_rm_del_thres",
			hssi_8g_rx_pcs_rate_match_empty_thres                                  => "dis_rm_empty_thres",
			hssi_8g_rx_pcs_rate_match_full_thres                                   => "dis_rm_full_thres",
			hssi_8g_rx_pcs_rate_match_ins_thres                                    => "dis_rm_ins_thres",
			hssi_8g_rx_pcs_rate_match_start_thres                                  => "dis_rm_start_thres",
			hssi_8g_rx_pcs_rx_clk_free_running                                     => "en_rx_clk_free_run",
			hssi_8g_rx_pcs_rx_clk2                                                 => "rcvd_clk_clk2",
			hssi_8g_rx_pcs_rx_pcs_urst                                             => "en_rx_pcs_urst",
			hssi_8g_rx_pcs_rx_rcvd_clk                                             => "rcvd_clk_rcvd_clk",
			hssi_8g_rx_pcs_rx_rd_clk                                               => "pld_rx_clk",
			hssi_8g_rx_pcs_rx_refclk                                               => "dis_refclk_sel",
			hssi_8g_rx_pcs_rx_wr_clk                                               => "rx_clk2_div_1_2_4",
			hssi_8g_rx_pcs_sup_mode                                                => "user_mode",
			hssi_8g_rx_pcs_symbol_swap                                             => "dis_symbol_swap",
			hssi_8g_rx_pcs_sync_sm_idle_eios                                       => "dis_syncsm_idle",
			hssi_8g_rx_pcs_test_bus_sel                                            => "tx_testbus",
			hssi_8g_rx_pcs_tx_rx_parallel_loopback                                 => "dis_plpbk",
			hssi_8g_rx_pcs_wa_boundary_lock_ctrl                                   => "auto_align_pld_ctrl",
			hssi_8g_rx_pcs_wa_clk_slip_spacing                                     => 16,
			hssi_8g_rx_pcs_wa_det_latency_sync_status_beh                          => "dont_care_assert_sync",
			hssi_8g_rx_pcs_wa_disp_err_flag                                        => "dis_disp_err_flag",
			hssi_8g_rx_pcs_wa_kchar                                                => "dis_kchar",
			hssi_8g_rx_pcs_wa_pd                                                   => "wa_pd_10",
			hssi_8g_rx_pcs_wa_pd_data                                              => "380",
			hssi_8g_rx_pcs_wa_pd_polarity                                          => "en_pd_both_pol",
			hssi_8g_rx_pcs_wa_pld_controlled                                       => "rising_edge_sensitive_dw",
			hssi_8g_rx_pcs_wa_renumber_data                                        => 3,
			hssi_8g_rx_pcs_wa_rgnumber_data                                        => 3,
			hssi_8g_rx_pcs_wa_rknumber_data                                        => 3,
			hssi_8g_rx_pcs_wa_rosnumber_data                                       => 1,
			hssi_8g_rx_pcs_wa_rvnumber_data                                        => 0,
			hssi_8g_rx_pcs_wa_sync_sm_ctrl                                         => "gige_sync_sm",
			hssi_8g_rx_pcs_wait_cnt                                                => 0,
			hssi_8g_tx_pcs_bit_reversal                                            => "dis_bit_reversal",
			hssi_8g_tx_pcs_bonding_dft_en                                          => "dft_dis",
			hssi_8g_tx_pcs_bonding_dft_val                                         => "dft_0",
			hssi_8g_tx_pcs_bypass_pipeline_reg                                     => "dis_bypass_pipeline",
			hssi_8g_tx_pcs_byte_serializer                                         => "dis_bs",
			hssi_8g_tx_pcs_clock_gate_bs_enc                                       => "dis_bs_enc_clk_gating",
			hssi_8g_tx_pcs_clock_gate_dw_fifowr                                    => "dis_dw_fifowr_clk_gating",
			hssi_8g_tx_pcs_clock_gate_fiford                                       => "dis_fiford_clk_gating",
			hssi_8g_tx_pcs_clock_gate_sw_fifowr                                    => "dis_sw_fifowr_clk_gating",
			hssi_8g_tx_pcs_clock_observation_in_pld_core                           => "internal_refclk_b",
			hssi_8g_tx_pcs_data_selection_8b10b_encoder_input                      => "normal_data_path",
			hssi_8g_tx_pcs_dynamic_clk_switch                                      => "dis_dyn_clk_switch",
			hssi_8g_tx_pcs_eightb_tenb_disp_ctrl                                   => "dis_disp_ctrl",
			hssi_8g_tx_pcs_eightb_tenb_encoder                                     => "dis_8b10b",
			hssi_8g_tx_pcs_force_echar                                             => "dis_force_echar",
			hssi_8g_tx_pcs_force_kchar                                             => "dis_force_kchar",
			hssi_8g_tx_pcs_gen3_tx_clk_sel                                         => "dis_tx_clk",
			hssi_8g_tx_pcs_gen3_tx_pipe_clk_sel                                    => "dis_tx_pipe_clk",
			hssi_8g_tx_pcs_hip_mode                                                => "dis_hip",
			hssi_8g_tx_pcs_pcs_bypass                                              => "dis_pcs_bypass",
			hssi_8g_tx_pcs_phase_comp_rdptr                                        => "enable_rdptr",
			hssi_8g_tx_pcs_phase_compensation_fifo                                 => "low_latency",
			hssi_8g_tx_pcs_phfifo_write_clk_sel                                    => "pld_tx_clk",
			hssi_8g_tx_pcs_pma_dw                                                  => "twenty_bit",
			hssi_8g_tx_pcs_prot_mode                                               => "basic",
			hssi_8g_tx_pcs_refclk_b_clk_sel                                        => "tx_pma_clock",
			hssi_8g_tx_pcs_revloop_back_rm                                         => "dis_rev_loopback_rx_rm",
			hssi_8g_tx_pcs_sup_mode                                                => "user_mode",
			hssi_8g_tx_pcs_symbol_swap                                             => "dis_symbol_swap",
			hssi_8g_tx_pcs_tx_bitslip                                              => "dis_tx_bitslip",
			hssi_8g_tx_pcs_tx_compliance_controlled_disparity                      => "dis_txcompliance",
			hssi_8g_tx_pcs_tx_fast_pld_reg                                         => "dis_tx_fast_pld_reg",
			hssi_8g_tx_pcs_txclk_freerun                                           => "en_freerun_tx",
			hssi_8g_tx_pcs_txpcs_urst                                              => "en_txpcs_urst",
			hssi_tx_pld_pcs_interface_hd_chnl_hip_en                               => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_prot_mode_tx                         => "basic_8gpcs_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_tx                => "individual_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_pma_dw_tx                            => "pma_20b_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_pld_fifo_mode_tx                     => "fifo_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_shared_fifo_width_tx                 => "single_tx",
			hssi_tx_pld_pcs_interface_hd_chnl_low_latency_en_tx                    => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_func_mode                            => "enable",
			hssi_tx_pld_pcs_interface_hd_chnl_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_chnl_lpbk_en                              => "disable",
			hssi_tx_pld_pcs_interface_hd_chnl_frequency_rules_en                   => "enable",
			hssi_tx_pld_pcs_interface_hd_chnl_pma_tx_clk_hz                        => 127000000,
			hssi_tx_pld_pcs_interface_hd_chnl_pld_tx_clk_hz                        => 127000000,
			hssi_tx_pld_pcs_interface_hd_chnl_pld_uhsif_tx_clk_hz                  => 0,
			hssi_tx_pld_pcs_interface_hd_fifo_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_fifo_prot_mode_tx                         => "non_teng_mode_tx",
			hssi_tx_pld_pcs_interface_hd_fifo_shared_fifo_width_tx                 => "single_tx",
			hssi_tx_pld_pcs_interface_hd_10g_channel_operation_mode                => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_10g_lpbk_en                               => "disable",
			hssi_tx_pld_pcs_interface_hd_10g_advanced_user_mode_tx                 => "disable",
			hssi_tx_pld_pcs_interface_hd_10g_pma_dw_tx                             => "pma_64b_tx",
			hssi_tx_pld_pcs_interface_hd_10g_fifo_mode_tx                          => "fifo_tx",
			hssi_tx_pld_pcs_interface_hd_10g_prot_mode_tx                          => "disabled_prot_mode_tx",
			hssi_tx_pld_pcs_interface_hd_10g_low_latency_en_tx                     => "disable",
			hssi_tx_pld_pcs_interface_hd_10g_shared_fifo_width_tx                  => "single_tx",
			hssi_tx_pld_pcs_interface_hd_8g_channel_operation_mode                 => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_8g_lpbk_en                                => "disable",
			hssi_tx_pld_pcs_interface_hd_8g_prot_mode_tx                           => "basic_tx",
			hssi_tx_pld_pcs_interface_hd_8g_hip_mode                               => "disable",
			hssi_tx_pld_pcs_interface_hd_8g_pma_dw_tx                              => "pma_20b_tx",
			hssi_tx_pld_pcs_interface_hd_8g_fifo_mode_tx                           => "fifo_tx",
			hssi_tx_pld_pcs_interface_hd_g3_prot_mode                              => "disabled_prot_mode",
			hssi_tx_pld_pcs_interface_hd_krfec_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_krfec_lpbk_en                             => "disable",
			hssi_tx_pld_pcs_interface_hd_krfec_prot_mode_tx                        => "disabled_prot_mode_tx",
			hssi_tx_pld_pcs_interface_hd_krfec_low_latency_en_tx                   => "disable",
			hssi_tx_pld_pcs_interface_hd_pmaif_lpbk_en                             => "disable",
			hssi_tx_pld_pcs_interface_hd_pmaif_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_tx_pld_pcs_interface_hd_pmaif_sim_mode                            => "disable",
			hssi_tx_pld_pcs_interface_hd_pmaif_prot_mode_tx                        => "eightg_basic_mode_tx",
			hssi_tx_pld_pcs_interface_hd_pmaif_pma_dw_tx                           => "pma_20b_tx",
			hssi_tx_pld_pcs_interface_hd_pldif_prot_mode_tx                        => "eightg_and_g3_pld_fifo_mode_tx",
			hssi_tx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        => "disable",
			hssi_tx_pld_pcs_interface_pcs_tx_clk_source                            => "eightg",
			hssi_tx_pld_pcs_interface_pcs_tx_data_source                           => "hip_disable",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_en                         => "delay1_clk_disable",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_clk_sel                        => "pcs_tx_clk",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_ctrl                           => "delay1_path0",
			hssi_tx_pld_pcs_interface_pcs_tx_delay1_data_sel                       => "one_ff_delay",
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_clk_en                         => "delay2_clk_disable",
			hssi_tx_pld_pcs_interface_pcs_tx_delay2_ctrl                           => "delay2_path0",
			hssi_tx_pld_pcs_interface_pcs_tx_output_sel                            => "teng_output",
			hssi_tx_pld_pcs_interface_pcs_tx_clk_out_sel                           => "eightg_clk_out",
			hssi_rx_pld_pcs_interface_hd_chnl_hip_en                               => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_transparent_pcs_rx                   => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_hrdrstctl_en                         => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_prot_mode_rx                         => "basic_8gpcs_rm_disable_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_ctrl_plane_bonding_rx                => "individual_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_pma_dw_rx                            => "pma_20b_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_pld_fifo_mode_rx                     => "fifo_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_shared_fifo_width_rx                 => "single_rx",
			hssi_rx_pld_pcs_interface_hd_chnl_low_latency_en_rx                    => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_func_mode                            => "enable",
			hssi_rx_pld_pcs_interface_hd_chnl_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_chnl_lpbk_en                              => "disable",
			hssi_rx_pld_pcs_interface_hd_10g_advanced_user_mode_rx                 => "disable",
			hssi_rx_pld_pcs_interface_hd_chnl_frequency_rules_en                   => "enable",
			hssi_rx_pld_pcs_interface_hd_chnl_pma_rx_clk_hz                        => 127000000,
			hssi_rx_pld_pcs_interface_hd_chnl_pld_rx_clk_hz                        => 127000000,
			hssi_rx_pld_pcs_interface_hd_chnl_fref_clk_hz                          => 127000000,
			hssi_rx_pld_pcs_interface_hd_chnl_clklow_clk_hz                        => 127000000,
			hssi_rx_pld_pcs_interface_hd_fifo_channel_operation_mode               => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_fifo_prot_mode_rx                         => "non_teng_mode_rx",
			hssi_rx_pld_pcs_interface_hd_fifo_shared_fifo_width_rx                 => "single_rx",
			hssi_rx_pld_pcs_interface_hd_10g_channel_operation_mode                => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_10g_lpbk_en                               => "disable",
			hssi_rx_pld_pcs_interface_hd_10g_pma_dw_rx                             => "pma_64b_rx",
			hssi_rx_pld_pcs_interface_hd_10g_fifo_mode_rx                          => "fifo_rx",
			hssi_rx_pld_pcs_interface_hd_10g_prot_mode_rx                          => "disabled_prot_mode_rx",
			hssi_rx_pld_pcs_interface_hd_10g_low_latency_en_rx                     => "disable",
			hssi_rx_pld_pcs_interface_hd_10g_shared_fifo_width_rx                  => "single_rx",
			hssi_rx_pld_pcs_interface_hd_10g_test_bus_mode                         => "rx",
			hssi_rx_pld_pcs_interface_hd_8g_channel_operation_mode                 => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_8g_lpbk_en                                => "disable",
			hssi_rx_pld_pcs_interface_hd_8g_prot_mode_rx                           => "basic_rm_disable_rx",
			hssi_rx_pld_pcs_interface_hd_8g_hip_mode                               => "disable",
			hssi_rx_pld_pcs_interface_hd_8g_pma_dw_rx                              => "pma_20b_rx",
			hssi_rx_pld_pcs_interface_hd_8g_fifo_mode_rx                           => "fifo_rx",
			hssi_rx_pld_pcs_interface_hd_g3_prot_mode                              => "disabled_prot_mode",
			hssi_rx_pld_pcs_interface_hd_krfec_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_krfec_lpbk_en                             => "disable",
			hssi_rx_pld_pcs_interface_hd_krfec_prot_mode_rx                        => "disabled_prot_mode_rx",
			hssi_rx_pld_pcs_interface_hd_krfec_low_latency_en_rx                   => "disable",
			hssi_rx_pld_pcs_interface_hd_krfec_test_bus_mode                       => "tx",
			hssi_rx_pld_pcs_interface_hd_pmaif_lpbk_en                             => "disable",
			hssi_rx_pld_pcs_interface_hd_pmaif_channel_operation_mode              => "tx_rx_pair_enabled",
			hssi_rx_pld_pcs_interface_hd_pmaif_sim_mode                            => "disable",
			hssi_rx_pld_pcs_interface_hd_pmaif_prot_mode_rx                        => "eightg_basic_mode_rx",
			hssi_rx_pld_pcs_interface_hd_pmaif_pma_dw_rx                           => "pma_20b_rx",
			hssi_rx_pld_pcs_interface_hd_pldif_prot_mode_rx                        => "eightg_and_g3_pld_fifo_mode_rx",
			hssi_rx_pld_pcs_interface_hd_pldif_hrdrstctl_en                        => "disable",
			hssi_rx_pld_pcs_interface_pcs_rx_block_sel                             => "eightg",
			hssi_rx_pld_pcs_interface_pcs_rx_clk_sel                               => "pld_rx_clk",
			hssi_rx_pld_pcs_interface_pcs_rx_hip_clk_en                            => "hip_rx_disable",
			hssi_rx_pld_pcs_interface_pcs_rx_output_sel                            => "teng_output",
			hssi_rx_pld_pcs_interface_pcs_rx_clk_out_sel                           => "eightg_clk_out",
			hssi_common_pld_pcs_interface_dft_clk_out_en                           => "dft_clk_out_disable",
			hssi_common_pld_pcs_interface_dft_clk_out_sel                          => "teng_rx_dft_clk",
			hssi_common_pld_pcs_interface_hrdrstctrl_en                            => "hrst_dis",
			hssi_common_pld_pcs_interface_pcs_testbus_block_sel                    => "pma_if",
			hssi_rx_pcs_pma_interface_block_sel                                    => "eight_g_pcs",
			hssi_rx_pcs_pma_interface_channel_operation_mode                       => "tx_rx_pair_enabled",
			hssi_rx_pcs_pma_interface_clkslip_sel                                  => "pld",
			hssi_rx_pcs_pma_interface_lpbk_en                                      => "disable",
			hssi_rx_pcs_pma_interface_master_clk_sel                               => "master_rx_pma_clk",
			hssi_rx_pcs_pma_interface_pldif_datawidth_mode                         => "pldif_data_10bit",
			hssi_rx_pcs_pma_interface_pma_dw_rx                                    => "pma_20b_rx",
			hssi_rx_pcs_pma_interface_pma_if_dft_en                                => "dft_dis",
			hssi_rx_pcs_pma_interface_pma_if_dft_val                               => "dft_0",
			hssi_rx_pcs_pma_interface_prbs_clken                                   => "prbs_clk_dis",
			hssi_rx_pcs_pma_interface_prbs_ver                                     => "prbs_off",
			hssi_rx_pcs_pma_interface_prbs9_dwidth                                 => "prbs9_64b",
			hssi_rx_pcs_pma_interface_prot_mode_rx                                 => "eightg_basic_mode_rx",
			hssi_rx_pcs_pma_interface_rx_dyn_polarity_inversion                    => "rx_dyn_polinv_dis",
			hssi_rx_pcs_pma_interface_rx_lpbk_en                                   => "lpbk_dis",
			hssi_rx_pcs_pma_interface_rx_prbs_force_signal_ok                      => "force_sig_ok",
			hssi_rx_pcs_pma_interface_rx_prbs_mask                                 => "prbsmask128",
			hssi_rx_pcs_pma_interface_rx_prbs_mode                                 => "teng_mode",
			hssi_rx_pcs_pma_interface_rx_signalok_signaldet_sel                    => "sel_sig_det",
			hssi_rx_pcs_pma_interface_rx_static_polarity_inversion                 => "rx_stat_polinv_dis",
			hssi_rx_pcs_pma_interface_rx_uhsif_lpbk_en                             => "uhsif_lpbk_dis",
			hssi_rx_pcs_pma_interface_sup_mode                                     => "user_mode",
			hssi_tx_pcs_pma_interface_bypass_pma_txelecidle                        => "true",
			hssi_tx_pcs_pma_interface_channel_operation_mode                       => "tx_rx_pair_enabled",
			hssi_tx_pcs_pma_interface_lpbk_en                                      => "disable",
			hssi_tx_pcs_pma_interface_master_clk_sel                               => "master_tx_pma_clk",
			hssi_tx_pcs_pma_interface_pcie_sub_prot_mode_tx                        => "other_prot_mode",
			hssi_tx_pcs_pma_interface_pldif_datawidth_mode                         => "pldif_data_10bit",
			hssi_tx_pcs_pma_interface_pma_dw_tx                                    => "pma_20b_tx",
			hssi_tx_pcs_pma_interface_pma_if_dft_en                                => "dft_dis",
			hssi_tx_pcs_pma_interface_pmagate_en                                   => "pmagate_dis",
			hssi_tx_pcs_pma_interface_prbs_clken                                   => "prbs_clk_dis",
			hssi_tx_pcs_pma_interface_prbs_gen_pat                                 => "prbs_gen_dis",
			hssi_tx_pcs_pma_interface_prbs9_dwidth                                 => "prbs9_64b",
			hssi_tx_pcs_pma_interface_prot_mode_tx                                 => "eightg_basic_mode_tx",
			hssi_tx_pcs_pma_interface_sq_wave_num                                  => "sq_wave_default",
			hssi_tx_pcs_pma_interface_sqwgen_clken                                 => "sqwgen_clk_dis",
			hssi_tx_pcs_pma_interface_sup_mode                                     => "user_mode",
			hssi_tx_pcs_pma_interface_tx_dyn_polarity_inversion                    => "tx_dyn_polinv_dis",
			hssi_tx_pcs_pma_interface_tx_pma_data_sel                              => "eight_g_pcs",
			hssi_tx_pcs_pma_interface_tx_static_polarity_inversion                 => "tx_stat_polinv_dis",
			hssi_tx_pcs_pma_interface_uhsif_cnt_step_filt_before_lock              => "uhsif_filt_stepsz_b4lock_2",
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_after_lock_value       => 0,
			hssi_tx_pcs_pma_interface_uhsif_cnt_thresh_filt_before_lock            => "uhsif_filt_cntthr_b4lock_8",
			hssi_tx_pcs_pma_interface_uhsif_dcn_test_update_period                 => "uhsif_dcn_test_period_4",
			hssi_tx_pcs_pma_interface_uhsif_dcn_testmode_enable                    => "uhsif_dcn_test_mode_disable",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_count_thresh                 => "uhsif_dzt_cnt_thr_2",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_detection_enable             => "uhsif_dzt_disable",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_obser_window                 => "uhsif_dzt_obr_win_16",
			hssi_tx_pcs_pma_interface_uhsif_dead_zone_skip_size                    => "uhsif_dzt_skipsz_4",
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_index_sel                   => "uhsif_index_cram",
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_margin                      => "uhsif_dcn_margin_2",
			hssi_tx_pcs_pma_interface_uhsif_delay_cell_static_index_value          => 0,
			hssi_tx_pcs_pma_interface_uhsif_dft_dead_zone_control                  => "uhsif_dft_dz_det_val_0",
			hssi_tx_pcs_pma_interface_uhsif_dft_up_filt_control                    => "uhsif_dft_up_val_0",
			hssi_tx_pcs_pma_interface_uhsif_enable                                 => "uhsif_disable",
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_after_lock              => "uhsif_lkd_segsz_aflock_512",
			hssi_tx_pcs_pma_interface_uhsif_lock_det_segsz_before_lock             => "uhsif_lkd_segsz_b4lock_16",
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_after_lock_value   => 0,
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_cnt_before_lock_value  => 0,
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_after_lock_value  => 0,
			hssi_tx_pcs_pma_interface_uhsif_lock_det_thresh_diff_before_lock_value => 0,
			hssi_common_pcs_pma_interface_asn_clk_enable                           => "false",
			hssi_common_pcs_pma_interface_asn_enable                               => "dis_asn",
			hssi_common_pcs_pma_interface_block_sel                                => "eight_g_pcs",
			hssi_common_pcs_pma_interface_bypass_early_eios                        => "true",
			hssi_common_pcs_pma_interface_bypass_pcie_switch                       => "true",
			hssi_common_pcs_pma_interface_bypass_pma_ltr                           => "true",
			hssi_common_pcs_pma_interface_bypass_pma_sw_done                       => "true",
			hssi_common_pcs_pma_interface_bypass_ppm_lock                          => "false",
			hssi_common_pcs_pma_interface_bypass_send_syncp_fbkp                   => "true",
			hssi_common_pcs_pma_interface_bypass_txdetectrx                        => "true",
			hssi_common_pcs_pma_interface_cdr_control                              => "dis_cdr_ctrl",
			hssi_common_pcs_pma_interface_cid_enable                               => "dis_cid_mode",
			hssi_common_pcs_pma_interface_data_mask_count                          => 0,
			hssi_common_pcs_pma_interface_data_mask_count_multi                    => 0,
			hssi_common_pcs_pma_interface_dft_observation_clock_selection          => "dft_clk_obsrv_tx0",
			hssi_common_pcs_pma_interface_early_eios_counter                       => 0,
			hssi_common_pcs_pma_interface_force_freqdet                            => "force_freqdet_dis",
			hssi_common_pcs_pma_interface_free_run_clk_enable                      => "false",
			hssi_common_pcs_pma_interface_ignore_sigdet_g23                        => "false",
			hssi_common_pcs_pma_interface_pc_en_counter                            => 0,
			hssi_common_pcs_pma_interface_pc_rst_counter                           => 0,
			hssi_common_pcs_pma_interface_pcie_hip_mode                            => "hip_disable",
			hssi_common_pcs_pma_interface_ph_fifo_reg_mode                         => "phfifo_reg_mode_dis",
			hssi_common_pcs_pma_interface_phfifo_flush_wait                        => 0,
			hssi_common_pcs_pma_interface_pipe_if_g3pcs                            => "pipe_if_8gpcs",
			hssi_common_pcs_pma_interface_pma_done_counter                         => 0,
			hssi_common_pcs_pma_interface_pma_if_dft_en                            => "dft_dis",
			hssi_common_pcs_pma_interface_pma_if_dft_val                           => "dft_0",
			hssi_common_pcs_pma_interface_ppm_cnt_rst                              => "ppm_cnt_rst_dis",
			hssi_common_pcs_pma_interface_ppm_deassert_early                       => "deassert_early_dis",
			hssi_common_pcs_pma_interface_ppm_gen1_2_cnt                           => "cnt_32k",
			hssi_common_pcs_pma_interface_ppm_post_eidle_delay                     => "cnt_200_cycles",
			hssi_common_pcs_pma_interface_ppmsel                                   => "ppmsel_1000",
			hssi_common_pcs_pma_interface_prot_mode                                => "other_protocols",
			hssi_common_pcs_pma_interface_rxvalid_mask                             => "rxvalid_mask_dis",
			hssi_common_pcs_pma_interface_sigdet_wait_counter                      => 0,
			hssi_common_pcs_pma_interface_sigdet_wait_counter_multi                => 0,
			hssi_common_pcs_pma_interface_sim_mode                                 => "disable",
			hssi_common_pcs_pma_interface_spd_chg_rst_wait_cnt_en                  => "false",
			hssi_common_pcs_pma_interface_sup_mode                                 => "user_mode",
			hssi_common_pcs_pma_interface_testout_sel                              => "asn_test",
			hssi_common_pcs_pma_interface_wait_clk_on_off_timer                    => 0,
			hssi_common_pcs_pma_interface_wait_pipe_synchronizing                  => 0,
			hssi_common_pcs_pma_interface_wait_send_syncp_fbkp                     => 0,
			hssi_common_pcs_pma_interface_ppm_det_buckets                          => "ppm_300_100_bucket",
			hssi_fifo_rx_pcs_double_read_mode                                      => "double_read_dis",
			hssi_fifo_rx_pcs_prot_mode                                             => "non_teng_mode",
			hssi_fifo_tx_pcs_double_write_mode                                     => "double_write_dis",
			hssi_fifo_tx_pcs_prot_mode                                             => "non_teng_mode",
			hssi_pipe_gen3_bypass_rx_detection_enable                              => "false",
			hssi_pipe_gen3_bypass_rx_preset                                        => 0,
			hssi_pipe_gen3_bypass_rx_preset_enable                                 => "false",
			hssi_pipe_gen3_bypass_tx_coefficent                                    => 0,
			hssi_pipe_gen3_bypass_tx_coefficent_enable                             => "false",
			hssi_pipe_gen3_elecidle_delay_g3                                       => 0,
			hssi_pipe_gen3_ind_error_reporting                                     => "dis_ind_error_reporting",
			hssi_pipe_gen3_mode                                                    => "disable_pcs",
			hssi_pipe_gen3_phy_status_delay_g12                                    => 0,
			hssi_pipe_gen3_phy_status_delay_g3                                     => 0,
			hssi_pipe_gen3_phystatus_rst_toggle_g12                                => "dis_phystatus_rst_toggle",
			hssi_pipe_gen3_phystatus_rst_toggle_g3                                 => "dis_phystatus_rst_toggle_g3",
			hssi_pipe_gen3_rate_match_pad_insertion                                => "dis_rm_fifo_pad_ins",
			hssi_pipe_gen3_sup_mode                                                => "user_mode",
			hssi_pipe_gen3_test_out_sel                                            => "disable_test_out",
			hssi_pipe_gen1_2_elec_idle_delay_val                                   => 0,
			hssi_pipe_gen1_2_error_replace_pad                                     => "replace_edb",
			hssi_pipe_gen1_2_hip_mode                                              => "dis_hip",
			hssi_pipe_gen1_2_ind_error_reporting                                   => "dis_ind_error_reporting",
			hssi_pipe_gen1_2_phystatus_delay_val                                   => 0,
			hssi_pipe_gen1_2_phystatus_rst_toggle                                  => "dis_phystatus_rst_toggle",
			hssi_pipe_gen1_2_pipe_byte_de_serializer_en                            => "dont_care_bds",
			hssi_pipe_gen1_2_prot_mode                                             => "basic",
			hssi_pipe_gen1_2_rx_pipe_enable                                        => "dis_pipe_rx",
			hssi_pipe_gen1_2_rxdetect_bypass                                       => "dis_rxdetect_bypass",
			hssi_pipe_gen1_2_sup_mode                                              => "user_mode",
			hssi_pipe_gen1_2_tx_pipe_enable                                        => "dis_pipe_tx",
			hssi_pipe_gen1_2_txswing                                               => "dis_txswing",
			pma_adapt_adp_1s_ctle_bypass                                           => "radp_1s_ctle_bypass_1",
			pma_adapt_adp_4s_ctle_bypass                                           => "radp_4s_ctle_bypass_1",
			pma_adapt_adp_ctle_en                                                  => "radp_ctle_disable",
			pma_adapt_adp_dfe_fltap_bypass                                         => "radp_dfe_fltap_bypass_1",
			pma_adapt_adp_dfe_fltap_en                                             => "radp_dfe_fltap_disable",
			pma_adapt_adp_dfe_fxtap_bypass                                         => "radp_dfe_fxtap_bypass_1",
			pma_adapt_adp_dfe_fxtap_en                                             => "radp_dfe_fxtap_disable",
			pma_adapt_adp_dfe_fxtap_hold_en                                        => "radp_dfe_fxtap_not_held",
			pma_adapt_adp_dfe_mode                                                 => "radp_dfe_mode_4",
			pma_adapt_adp_vga_bypass                                               => "radp_vga_bypass_1",
			pma_adapt_adp_vga_en                                                   => "radp_vga_disable",
			pma_adapt_adp_vref_bypass                                              => "radp_vref_bypass_1",
			pma_adapt_adp_vref_en                                                  => "radp_vref_disable",
			pma_adapt_datarate                                                     => "2540000000 bps",
			pma_adapt_prot_mode                                                    => "basic_rx",
			pma_adapt_sup_mode                                                     => "user_mode",
			pma_adapt_adp_ctle_adapt_cycle_window                                  => "radp_ctle_adapt_cycle_window_7",
			pma_adapt_odi_dfe_spec_en                                              => "rodi_dfe_spec_en_0",
			pma_adapt_adapt_mode                                                   => "manual",
			pma_adapt_adp_onetime_dfe                                              => "radp_onetime_dfe_0",
			pma_adapt_adp_mode                                                     => "radp_mode_8",
			pma_cdr_refclk_powerdown_mode                                          => "powerup",
			pma_cdr_refclk_refclk_select                                           => "ref_iqclk0",
			pma_cgb_bitslip_enable                                                 => "disable_bitslip",
			pma_cgb_bonding_reset_enable                                           => "disallow_bonding_reset",
			pma_cgb_datarate                                                       => "2540000000 bps",
			pma_cgb_pcie_gen3_bitwidth                                             => "pciegen3_wide",
			pma_cgb_prot_mode                                                      => "basic_tx",
			pma_cgb_ser_mode                                                       => "twenty_bit",
			pma_cgb_sup_mode                                                       => "user_mode",
			pma_cgb_x1_div_m_sel                                                   => "divbypass",
			pma_cgb_input_select_x1                                                => "fpll_bot",
			pma_cgb_input_select_gen3                                              => "unused",
			pma_cgb_input_select_xn                                                => "unused",
			pma_cgb_tx_ucontrol_en                                                 => "disable",
			pma_rx_dfe_datarate                                                    => "2540000000 bps",
			pma_rx_dfe_dft_en                                                      => "dft_disable",
			pma_rx_dfe_pdb                                                         => "dfe_enable",
			pma_rx_dfe_pdb_fixedtap                                                => "fixtap_dfe_powerdown",
			pma_rx_dfe_pdb_floattap                                                => "floattap_dfe_powerdown",
			pma_rx_dfe_pdb_fxtap4t7                                                => "fxtap4t7_powerdown",
			pma_rx_dfe_sup_mode                                                    => "user_mode",
			pma_rx_dfe_prot_mode                                                   => "basic_rx",
			pma_rx_odi_datarate                                                    => "2540000000 bps",
			pma_rx_odi_sup_mode                                                    => "user_mode",
			pma_rx_odi_step_ctrl_sel                                               => "dprio_mode",
			pma_rx_odi_prot_mode                                                   => "basic_rx",
			pma_rx_buf_bypass_eqz_stages_234                                       => "bypass_off",
			pma_rx_buf_datarate                                                    => "2540000000 bps",
			pma_rx_buf_diag_lp_en                                                  => "dlp_off",
			pma_rx_buf_prot_mode                                                   => "basic_rx",
			pma_rx_buf_qpi_enable                                                  => "non_qpi_mode",
			pma_rx_buf_rx_refclk_divider                                           => "bypass_divider",
			pma_rx_buf_sup_mode                                                    => "user_mode",
			pma_rx_buf_loopback_modes                                              => "lpbk_disable",
			pma_rx_buf_refclk_en                                                   => "disable",
			pma_rx_buf_pm_tx_rx_pcie_gen                                           => "non_pcie",
			pma_rx_buf_pm_tx_rx_pcie_gen_bitwidth                                  => "pcie_gen3_32b",
			pma_rx_buf_pm_tx_rx_cvp_mode                                           => "cvp_off",
			pma_rx_buf_xrx_path_uc_cal_enable                                      => "rx_cal_off",
			pma_rx_buf_xrx_path_sup_mode                                           => "user_mode",
			pma_rx_buf_xrx_path_prot_mode                                          => "basic_rx",
			pma_rx_buf_xrx_path_datarate                                           => "2540000000 bps",
			pma_rx_buf_xrx_path_datawidth                                          => 20,
			pma_rx_buf_xrx_path_pma_rx_divclk_hz                                   => "127000000",
			pma_rx_sd_prot_mode                                                    => "basic_rx",
			pma_rx_sd_sd_output_off                                                => 1,
			pma_rx_sd_sd_output_on                                                 => 15,
			pma_rx_sd_sd_pdb                                                       => "sd_off",
			pma_rx_sd_sup_mode                                                     => "user_mode",
			pma_tx_ser_ser_clk_divtx_user_sel                                      => "divtx_user_off",
			pma_tx_ser_sup_mode                                                    => "user_mode",
			pma_tx_ser_prot_mode                                                   => "basic_tx",
			pma_tx_buf_datarate                                                    => "2540000000 bps",
			pma_tx_buf_prot_mode                                                   => "basic_tx",
			pma_tx_buf_rx_det                                                      => "mode_0",
			pma_tx_buf_rx_det_output_sel                                           => "rx_det_pcie_out",
			pma_tx_buf_rx_det_pdb                                                  => "rx_det_off",
			pma_tx_buf_sup_mode                                                    => "user_mode",
			pma_tx_buf_user_fir_coeff_ctrl_sel                                     => "ram_ctl",
			pma_tx_buf_xtx_path_prot_mode                                          => "basic_tx",
			pma_tx_buf_xtx_path_datarate                                           => "2540000000 bps",
			pma_tx_buf_xtx_path_datawidth                                          => 20,
			pma_tx_buf_xtx_path_clock_divider_ratio                                => 1,
			pma_tx_buf_xtx_path_pma_tx_divclk_hz                                   => "127000000",
			pma_tx_buf_xtx_path_tx_pll_clk_hz                                      => "1270000000",
			pma_tx_buf_xtx_path_sup_mode                                           => "user_mode",
			cdr_pll_pma_width                                                      => 20,
			cdr_pll_cgb_div                                                        => 1,
			cdr_pll_is_cascaded_pll                                                => "false",
			cdr_pll_datarate                                                       => "2540000000 bps",
			cdr_pll_lpd_counter                                                    => 4,
			cdr_pll_lpfd_counter                                                   => 1,
			cdr_pll_n_counter_scratch                                              => 1,
			cdr_pll_output_clock_frequency                                         => "1270000000 Hz",
			cdr_pll_reference_clock_frequency                                      => "127000000 hz",
			cdr_pll_set_cdr_vco_speed                                              => 3,
			cdr_pll_set_cdr_vco_speed_fix                                          => 60,
			cdr_pll_vco_freq                                                       => "5080000000 Hz",
			cdr_pll_atb_select_control                                             => "atb_off",
			cdr_pll_auto_reset_on                                                  => "auto_reset_off",
			cdr_pll_bbpd_data_pattern_filter_select                                => "bbpd_data_pat_off",
			cdr_pll_bw_sel                                                         => "medium",
			cdr_pll_cdr_odi_select                                                 => "sel_cdr",
			cdr_pll_cdr_phaselock_mode                                             => "no_ignore_lock",
			cdr_pll_cdr_powerdown_mode                                             => "power_up",
			cdr_pll_chgpmp_current_pd                                              => "cp_current_pd_setting0",
			cdr_pll_chgpmp_current_pfd                                             => "cp_current_pfd_setting3",
			cdr_pll_chgpmp_replicate                                               => "false",
			cdr_pll_chgpmp_testmode                                                => "cp_test_disable",
			cdr_pll_clklow_mux_select                                              => "clklow_mux_cdr_fbclk",
			cdr_pll_diag_loopback_enable                                           => "false",
			cdr_pll_disable_up_dn                                                  => "true",
			cdr_pll_fref_clklow_div                                                => 1,
			cdr_pll_fref_mux_select                                                => "fref_mux_cdr_refclk",
			cdr_pll_gpon_lck2ref_control                                           => "gpon_lck2ref_off",
			cdr_pll_initial_settings                                               => "true",
			cdr_pll_lck2ref_delay_control                                          => "lck2ref_delay_2",
			cdr_pll_lf_resistor_pd                                                 => "lf_pd_setting3",
			cdr_pll_lf_resistor_pfd                                                => "lf_pfd_setting2",
			cdr_pll_lf_ripple_cap                                                  => "lf_no_ripple",
			cdr_pll_loop_filter_bias_select                                        => "lpflt_bias_7",
			cdr_pll_loopback_mode                                                  => "loopback_disabled",
			cdr_pll_ltd_ltr_micro_controller_select                                => "ltd_ltr_pcs",
			cdr_pll_m_counter                                                      => 40,
			cdr_pll_n_counter                                                      => 1,
			cdr_pll_pd_fastlock_mode                                               => "false",
			cdr_pll_pd_l_counter                                                   => 4,
			cdr_pll_pfd_l_counter                                                  => 1,
			cdr_pll_primary_use                                                    => "cdr",
			cdr_pll_prot_mode                                                      => "basic_rx",
			cdr_pll_reverse_serial_loopback                                        => "no_loopback",
			cdr_pll_set_cdr_v2i_enable                                             => "true",
			cdr_pll_set_cdr_vco_reset                                              => "false",
			cdr_pll_set_cdr_vco_speed_pciegen3                                     => "cdr_vco_max_speedbin_pciegen3",
			cdr_pll_sup_mode                                                       => "user_mode",
			cdr_pll_tx_pll_prot_mode                                               => "txpll_unused",
			cdr_pll_txpll_hclk_driver_enable                                       => "false",
			cdr_pll_vco_overrange_voltage                                          => "vco_overrange_off",
			cdr_pll_vco_underrange_voltage                                         => "vco_underange_off",
			cdr_pll_fb_select                                                      => "direct_fb",
			cdr_pll_uc_ro_cal                                                      => "uc_ro_cal_on",
			cdr_pll_iqclk_mux_sel                                                  => "power_down",
			cdr_pll_pcie_gen                                                       => "non_pcie",
			cdr_pll_set_cdr_input_freq_range                                       => 0,
			cdr_pll_chgpmp_current_dn_trim                                         => "cp_current_trimming_dn_setting0",
			cdr_pll_chgpmp_up_pd_trim_double                                       => "normal_up_trim_current",
			cdr_pll_chgpmp_current_up_pd                                           => "cp_current_pd_up_setting4",
			cdr_pll_chgpmp_current_up_trim                                         => "cp_current_trimming_up_setting0",
			cdr_pll_chgpmp_dn_pd_trim_double                                       => "normal_dn_trim_current",
			cdr_pll_cal_vco_count_length                                           => "sel_8b_count",
			cdr_pll_chgpmp_current_dn_pd                                           => "cp_current_pd_dn_setting4",
			pma_rx_deser_clkdiv_source                                             => "vco_bypass_normal",
			pma_rx_deser_clkdivrx_user_mode                                        => "clkdivrx_user_disabled",
			pma_rx_deser_datarate                                                  => "2540000000 bps",
			pma_rx_deser_deser_factor                                              => 20,
			pma_rx_deser_force_clkdiv_for_testing                                  => "normal_clkdiv",
			pma_rx_deser_sdclk_enable                                              => "false",
			pma_rx_deser_sup_mode                                                  => "user_mode",
			pma_rx_deser_rst_n_adapt_odi                                           => "no_rst_adapt_odi",
			pma_rx_deser_bitslip_bypass                                            => "bs_bypass_yes",
			pma_rx_deser_prot_mode                                                 => "basic_rx",
			pma_rx_deser_pcie_gen                                                  => "non_pcie",
			pma_rx_deser_pcie_gen_bitwidth                                         => "pcie_gen3_32b"
		)
		port map (
			tx_analogreset(0)         => xcvr_reset_control_0_tx_analogreset0_tx_analogreset,                                                                                                                                                                                                                --         tx_analogreset_ch0.tx_analogreset
			tx_analogreset(1)         => xcvr_reset_control_0_tx_analogreset1_tx_analogreset,                                                                                                                                                                                                                --                           .tx_analogreset
			tx_analogreset(2)         => xcvr_reset_control_0_tx_analogreset2_tx_analogreset,                                                                                                                                                                                                                --                           .tx_analogreset
			tx_analogreset(3)         => xcvr_reset_control_0_tx_analogreset3_tx_analogreset,                                                                                                                                                                                                                --                           .tx_analogreset
			tx_digitalreset(0)        => xcvr_reset_control_0_tx_digitalreset0_tx_digitalreset,                                                                                                                                                                                                              --        tx_digitalreset_ch0.tx_digitalreset
			tx_digitalreset(1)        => xcvr_reset_control_0_tx_digitalreset1_tx_digitalreset,                                                                                                                                                                                                              --                           .tx_digitalreset
			tx_digitalreset(2)        => xcvr_reset_control_0_tx_digitalreset2_tx_digitalreset,                                                                                                                                                                                                              --                           .tx_digitalreset
			tx_digitalreset(3)        => xcvr_reset_control_0_tx_digitalreset3_tx_digitalreset,                                                                                                                                                                                                              --                           .tx_digitalreset
			rx_analogreset(0)         => xcvr_reset_control_0_rx_analogreset0_rx_analogreset,                                                                                                                                                                                                                --         rx_analogreset_ch0.rx_analogreset
			rx_analogreset(1)         => xcvr_reset_control_0_rx_analogreset1_rx_analogreset,                                                                                                                                                                                                                --                           .rx_analogreset
			rx_analogreset(2)         => xcvr_reset_control_0_rx_analogreset2_rx_analogreset,                                                                                                                                                                                                                --                           .rx_analogreset
			rx_analogreset(3)         => xcvr_reset_control_0_rx_analogreset3_rx_analogreset,                                                                                                                                                                                                                --                           .rx_analogreset
			rx_digitalreset(0)        => xcvr_reset_control_0_rx_digitalreset0_rx_digitalreset,                                                                                                                                                                                                              --        rx_digitalreset_ch0.rx_digitalreset
			rx_digitalreset(1)        => xcvr_reset_control_0_rx_digitalreset1_rx_digitalreset,                                                                                                                                                                                                              --                           .rx_digitalreset
			rx_digitalreset(2)        => xcvr_reset_control_0_rx_digitalreset2_rx_digitalreset,                                                                                                                                                                                                              --                           .rx_digitalreset
			rx_digitalreset(3)        => xcvr_reset_control_0_rx_digitalreset3_rx_digitalreset,                                                                                                                                                                                                              --                           .rx_digitalreset
			tx_cal_busy(0)            => xcvr_native_a10_0_tx_cal_busy(0),                                                                                                                                                                                                                                   --            tx_cal_busy_ch0.tx_cal_busy
			tx_cal_busy(1)            => xcvr_native_a10_0_tx_cal_busy(1),                                                                                                                                                                                                                                   --                           .tx_cal_busy
			tx_cal_busy(2)            => xcvr_native_a10_0_tx_cal_busy(2),                                                                                                                                                                                                                                   --                           .tx_cal_busy
			tx_cal_busy(3)            => xcvr_native_a10_0_tx_cal_busy(3),                                                                                                                                                                                                                                   --                           .tx_cal_busy
			rx_cal_busy(0)            => xcvr_native_a10_0_rx_cal_busy(0),                                                                                                                                                                                                                                   --            rx_cal_busy_ch0.rx_cal_busy
			rx_cal_busy(1)            => xcvr_native_a10_0_rx_cal_busy(1),                                                                                                                                                                                                                                   --                           .rx_cal_busy
			rx_cal_busy(2)            => xcvr_native_a10_0_rx_cal_busy(2),                                                                                                                                                                                                                                   --                           .rx_cal_busy
			rx_cal_busy(3)            => xcvr_native_a10_0_rx_cal_busy(3),                                                                                                                                                                                                                                   --                           .rx_cal_busy
			tx_serial_clk0(0)         => xcvr_atx_pll_a10_0_tx_serial_clk_clk,                                                                                                                                                                                                                               --         tx_serial_clk0_ch0.clk
			tx_serial_clk0(1)         => xcvr_atx_pll_a10_0_tx_serial_clk_clk,                                                                                                                                                                                                                               --                           .clk
			tx_serial_clk0(2)         => xcvr_atx_pll_a10_0_tx_serial_clk_clk,                                                                                                                                                                                                                               --                           .clk
			tx_serial_clk0(3)         => xcvr_atx_pll_a10_0_tx_serial_clk_clk,                                                                                                                                                                                                                               --                           .clk
			rx_cdr_refclk0            => clk_clk,                                                                                                                                                                                                                                                            --             rx_cdr_refclk0.clk
			tx_serial_data(0)         => xcvr_native_a10_0_tx_serial_data(0),                                                                                                                                                                                                                                --         tx_serial_data_ch0.tx_serial_data
			tx_serial_data(1)         => xcvr_native_a10_0_tx_serial_data(1),                                                                                                                                                                                                                                --                           .tx_serial_data
			tx_serial_data(2)         => xcvr_native_a10_0_tx_serial_data(2),                                                                                                                                                                                                                                --                           .tx_serial_data
			tx_serial_data(3)         => xcvr_native_a10_0_tx_serial_data(3),                                                                                                                                                                                                                                --                           .tx_serial_data
			rx_serial_data(0)         => xcvr_native_a10_0_rx_serial_data_ch0_rx_serial_data,                                                                                                                                                                                                                --         rx_serial_data_ch0.rx_serial_data
			rx_serial_data(1)         => xcvr_native_a10_0_rx_serial_data_ch1_rx_serial_data,                                                                                                                                                                                                                --                           .rx_serial_data
			rx_serial_data(2)         => xcvr_native_a10_0_rx_serial_data_ch2_rx_serial_data,                                                                                                                                                                                                                --                           .rx_serial_data
			rx_serial_data(3)         => xcvr_native_a10_0_rx_serial_data_ch3_rx_serial_data,                                                                                                                                                                                                                --                           .rx_serial_data
			rx_seriallpbken(0)        => xcvr_native_a10_0_rx_seriallpbken_ch0_rx_seriallpbken,                                                                                                                                                                                                              --        rx_seriallpbken_ch0.rx_seriallpbken
			rx_seriallpbken(1)        => xcvr_native_a10_0_rx_seriallpbken_ch1_rx_seriallpbken,                                                                                                                                                                                                              --                           .rx_seriallpbken
			rx_seriallpbken(2)        => xcvr_native_a10_0_rx_seriallpbken_ch2_rx_seriallpbken,                                                                                                                                                                                                              --                           .rx_seriallpbken
			rx_seriallpbken(3)        => xcvr_native_a10_0_rx_seriallpbken_ch3_rx_seriallpbken,                                                                                                                                                                                                              --                           .rx_seriallpbken
			rx_is_lockedtodata(0)     => xcvr_native_a10_0_rx_is_lockedtodata(0),                                                                                                                                                                                                                            --     rx_is_lockedtodata_ch0.rx_is_lockedtodata
			rx_is_lockedtodata(1)     => xcvr_native_a10_0_rx_is_lockedtodata(1),                                                                                                                                                                                                                            --                           .rx_is_lockedtodata
			rx_is_lockedtodata(2)     => xcvr_native_a10_0_rx_is_lockedtodata(2),                                                                                                                                                                                                                            --                           .rx_is_lockedtodata
			rx_is_lockedtodata(3)     => xcvr_native_a10_0_rx_is_lockedtodata(3),                                                                                                                                                                                                                            --                           .rx_is_lockedtodata
			tx_coreclkin(0)           => xcvr_native_a10_0_tx_coreclkin_ch0_clk,                                                                                                                                                                                                                             --           tx_coreclkin_ch0.clk
			tx_coreclkin(1)           => xcvr_native_a10_0_tx_coreclkin_ch1_clk,                                                                                                                                                                                                                             --                           .clk
			tx_coreclkin(2)           => xcvr_native_a10_0_tx_coreclkin_ch2_clk,                                                                                                                                                                                                                             --                           .clk
			tx_coreclkin(3)           => xcvr_native_a10_0_tx_coreclkin_ch3_clk,                                                                                                                                                                                                                             --                           .clk
			rx_coreclkin(0)           => xcvr_native_a10_0_rx_coreclkin_ch0_clk,                                                                                                                                                                                                                             --           rx_coreclkin_ch0.clk
			rx_coreclkin(1)           => xcvr_native_a10_0_rx_coreclkin_ch1_clk,                                                                                                                                                                                                                             --                           .clk
			rx_coreclkin(2)           => xcvr_native_a10_0_rx_coreclkin_ch2_clk,                                                                                                                                                                                                                             --                           .clk
			rx_coreclkin(3)           => xcvr_native_a10_0_rx_coreclkin_ch3_clk,                                                                                                                                                                                                                             --                           .clk
			tx_clkout(0)              => xcvr_native_a10_0_tx_clkout(0),                                                                                                                                                                                                                                     --              tx_clkout_ch0.clk
			tx_clkout(1)              => xcvr_native_a10_0_tx_clkout(1),                                                                                                                                                                                                                                     --                           .clk
			tx_clkout(2)              => xcvr_native_a10_0_tx_clkout(2),                                                                                                                                                                                                                                     --                           .clk
			tx_clkout(3)              => xcvr_native_a10_0_tx_clkout(3),                                                                                                                                                                                                                                     --                           .clk
			rx_clkout(0)              => xcvr_native_a10_0_rx_clkout(0),                                                                                                                                                                                                                                     --              rx_clkout_ch0.clk
			rx_clkout(1)              => xcvr_native_a10_0_rx_clkout(1),                                                                                                                                                                                                                                     --                           .clk
			rx_clkout(2)              => xcvr_native_a10_0_rx_clkout(2),                                                                                                                                                                                                                                     --                           .clk
			rx_clkout(3)              => xcvr_native_a10_0_rx_clkout(3),                                                                                                                                                                                                                                     --                           .clk
			tx_parallel_data(0)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(0),                                                                                                                                                                                                         --       tx_parallel_data_ch0.tx_parallel_data
			tx_parallel_data(1)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(1),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(2)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(2),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(3)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(3),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(4)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(4),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(5)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(5),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(6)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(6),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(7)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(7),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(8)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(8),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(9)       => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(9),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(10)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(0),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(11)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(10),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(12)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(11),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(13)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(12),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(14)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(13),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(15)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(14),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(16)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(15),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(17)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(16),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(18)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(17),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(19)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(18),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(20)      => xcvr_native_a10_0_tx_parallel_data_ch0_tx_parallel_data(19),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(21)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(1),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(22)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(2),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(23)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(3),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(24)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(4),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(25)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(5),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(26)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(6),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(27)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(7),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(28)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(8),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(29)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(9),                                                                                                                                                                                               --                           .tx_parallel_data
			tx_parallel_data(30)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(10),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(31)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(11),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(32)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(12),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(33)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(13),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(34)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(14),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(35)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(15),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(36)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(16),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(37)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(17),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(38)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(18),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(39)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(19),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(40)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(20),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(41)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(21),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(42)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(22),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(43)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(23),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(44)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(24),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(45)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(25),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(46)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(26),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(47)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(27),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(48)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(28),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(49)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(29),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(50)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(30),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(51)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(31),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(52)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(32),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(53)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(33),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(54)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(34),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(55)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(35),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(56)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(36),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(57)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(37),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(58)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(38),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(59)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(39),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(60)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(40),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(61)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(41),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(62)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(42),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(63)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(43),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(64)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(44),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(65)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(45),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(66)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(46),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(67)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(47),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(68)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(48),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(69)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(49),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(70)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(50),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(71)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(51),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(72)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(52),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(73)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(53),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(74)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(54),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(75)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(55),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(76)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(56),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(77)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(57),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(78)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(58),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(79)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(59),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(80)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(60),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(81)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(61),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(82)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(62),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(83)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(63),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(84)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(64),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(85)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(65),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(86)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(66),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(87)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(67),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(88)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(68),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(89)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(69),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(90)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(70),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(91)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(71),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(92)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(72),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(93)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(73),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(94)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(74),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(95)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(75),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(96)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(76),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(97)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(77),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(98)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(78),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(99)      => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(79),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(100)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(80),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(101)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(81),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(102)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(82),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(103)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(83),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(104)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(84),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(105)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(85),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(106)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(86),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(107)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(87),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(108)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(88),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(109)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(89),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(110)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(90),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(111)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(91),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(112)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(92),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(113)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(93),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(114)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(94),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(115)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(95),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(116)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(96),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(117)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(97),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(118)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(98),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(119)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(99),                                                                                                                                                                                              --                           .tx_parallel_data
			tx_parallel_data(120)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(100),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(121)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(101),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(122)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(102),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(123)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(103),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(124)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(104),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(125)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(105),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(126)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(106),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(127)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(107),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(128)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(0),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(129)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(1),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(130)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(2),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(131)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(3),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(132)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(4),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(133)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(5),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(134)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(6),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(135)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(7),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(136)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(8),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(137)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(9),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(138)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(108),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(139)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(10),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(140)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(11),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(141)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(12),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(142)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(13),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(143)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(14),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(144)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(15),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(145)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(16),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(146)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(17),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(147)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(18),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(148)     => xcvr_native_a10_0_tx_parallel_data_ch1_tx_parallel_data(19),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(149)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(109),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(150)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(110),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(151)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(111),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(152)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(112),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(153)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(113),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(154)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(114),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(155)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(115),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(156)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(116),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(157)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(117),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(158)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(118),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(159)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(119),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(160)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(120),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(161)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(121),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(162)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(122),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(163)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(123),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(164)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(124),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(165)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(125),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(166)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(126),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(167)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(127),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(168)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(128),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(169)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(129),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(170)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(130),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(171)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(131),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(172)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(132),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(173)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(133),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(174)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(134),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(175)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(135),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(176)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(136),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(177)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(137),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(178)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(138),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(179)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(139),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(180)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(140),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(181)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(141),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(182)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(142),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(183)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(143),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(184)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(144),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(185)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(145),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(186)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(146),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(187)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(147),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(188)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(148),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(189)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(149),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(190)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(150),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(191)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(151),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(192)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(152),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(193)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(153),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(194)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(154),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(195)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(155),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(196)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(156),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(197)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(157),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(198)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(158),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(199)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(159),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(200)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(160),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(201)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(161),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(202)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(162),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(203)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(163),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(204)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(164),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(205)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(165),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(206)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(166),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(207)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(167),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(208)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(168),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(209)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(169),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(210)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(170),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(211)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(171),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(212)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(172),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(213)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(173),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(214)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(174),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(215)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(175),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(216)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(176),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(217)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(177),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(218)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(178),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(219)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(179),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(220)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(180),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(221)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(181),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(222)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(182),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(223)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(183),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(224)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(184),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(225)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(185),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(226)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(186),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(227)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(187),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(228)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(188),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(229)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(189),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(230)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(190),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(231)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(191),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(232)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(192),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(233)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(193),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(234)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(194),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(235)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(195),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(236)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(196),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(237)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(197),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(238)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(198),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(239)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(199),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(240)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(200),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(241)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(201),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(242)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(202),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(243)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(203),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(244)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(204),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(245)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(205),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(246)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(206),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(247)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(207),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(248)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(208),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(249)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(209),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(250)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(210),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(251)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(211),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(252)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(212),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(253)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(213),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(254)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(214),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(255)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(215),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(256)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(0),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(257)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(1),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(258)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(2),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(259)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(3),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(260)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(4),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(261)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(5),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(262)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(6),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(263)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(7),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(264)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(8),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(265)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(9),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(266)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(216),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(267)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(10),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(268)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(11),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(269)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(12),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(270)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(13),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(271)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(14),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(272)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(15),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(273)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(16),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(274)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(17),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(275)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(18),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(276)     => xcvr_native_a10_0_tx_parallel_data_ch2_tx_parallel_data(19),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(277)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(217),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(278)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(218),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(279)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(219),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(280)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(220),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(281)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(221),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(282)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(222),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(283)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(223),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(284)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(224),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(285)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(225),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(286)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(226),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(287)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(227),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(288)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(228),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(289)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(229),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(290)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(230),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(291)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(231),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(292)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(232),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(293)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(233),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(294)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(234),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(295)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(235),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(296)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(236),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(297)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(237),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(298)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(238),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(299)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(239),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(300)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(240),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(301)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(241),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(302)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(242),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(303)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(243),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(304)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(244),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(305)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(245),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(306)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(246),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(307)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(247),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(308)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(248),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(309)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(249),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(310)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(250),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(311)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(251),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(312)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(252),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(313)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(253),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(314)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(254),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(315)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(255),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(316)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(256),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(317)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(257),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(318)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(258),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(319)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(259),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(320)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(260),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(321)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(261),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(322)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(262),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(323)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(263),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(324)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(264),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(325)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(265),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(326)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(266),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(327)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(267),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(328)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(268),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(329)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(269),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(330)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(270),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(331)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(271),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(332)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(272),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(333)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(273),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(334)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(274),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(335)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(275),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(336)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(276),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(337)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(277),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(338)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(278),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(339)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(279),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(340)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(280),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(341)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(281),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(342)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(282),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(343)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(283),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(344)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(284),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(345)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(285),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(346)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(286),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(347)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(287),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(348)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(288),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(349)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(289),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(350)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(290),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(351)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(291),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(352)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(292),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(353)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(293),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(354)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(294),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(355)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(295),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(356)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(296),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(357)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(297),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(358)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(298),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(359)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(299),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(360)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(300),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(361)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(301),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(362)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(302),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(363)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(303),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(364)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(304),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(365)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(305),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(366)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(306),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(367)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(307),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(368)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(308),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(369)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(309),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(370)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(310),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(371)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(311),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(372)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(312),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(373)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(313),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(374)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(314),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(375)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(315),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(376)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(316),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(377)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(317),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(378)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(318),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(379)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(319),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(380)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(320),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(381)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(321),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(382)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(322),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(383)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(323),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(384)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(0),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(385)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(1),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(386)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(2),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(387)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(3),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(388)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(4),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(389)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(5),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(390)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(6),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(391)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(7),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(392)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(8),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(393)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(9),                                                                                                                                                                                                         --                           .tx_parallel_data
			tx_parallel_data(394)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(324),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(395)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(10),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(396)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(11),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(397)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(12),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(398)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(13),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(399)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(14),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(400)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(15),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(401)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(16),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(402)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(17),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(403)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(18),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(404)     => xcvr_native_a10_0_tx_parallel_data_ch3_tx_parallel_data(19),                                                                                                                                                                                                        --                           .tx_parallel_data
			tx_parallel_data(405)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(325),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(406)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(326),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(407)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(327),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(408)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(328),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(409)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(329),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(410)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(330),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(411)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(331),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(412)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(332),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(413)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(333),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(414)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(334),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(415)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(335),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(416)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(336),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(417)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(337),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(418)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(338),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(419)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(339),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(420)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(340),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(421)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(341),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(422)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(342),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(423)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(343),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(424)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(344),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(425)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(345),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(426)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(346),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(427)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(347),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(428)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(348),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(429)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(349),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(430)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(350),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(431)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(351),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(432)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(352),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(433)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(353),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(434)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(354),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(435)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(355),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(436)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(356),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(437)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(357),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(438)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(358),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(439)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(359),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(440)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(360),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(441)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(361),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(442)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(362),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(443)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(363),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(444)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(364),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(445)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(365),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(446)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(366),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(447)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(367),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(448)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(368),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(449)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(369),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(450)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(370),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(451)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(371),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(452)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(372),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(453)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(373),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(454)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(374),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(455)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(375),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(456)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(376),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(457)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(377),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(458)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(378),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(459)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(379),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(460)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(380),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(461)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(381),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(462)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(382),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(463)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(383),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(464)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(384),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(465)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(385),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(466)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(386),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(467)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(387),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(468)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(388),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(469)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(389),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(470)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(390),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(471)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(391),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(472)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(392),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(473)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(393),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(474)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(394),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(475)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(395),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(476)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(396),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(477)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(397),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(478)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(398),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(479)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(399),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(480)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(400),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(481)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(401),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(482)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(402),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(483)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(403),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(484)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(404),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(485)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(405),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(486)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(406),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(487)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(407),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(488)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(408),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(489)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(409),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(490)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(410),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(491)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(411),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(492)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(412),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(493)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(413),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(494)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(414),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(495)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(415),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(496)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(416),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(497)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(417),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(498)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(418),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(499)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(419),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(500)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(420),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(501)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(421),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(502)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(422),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(503)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(423),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(504)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(424),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(505)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(425),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(506)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(426),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(507)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(427),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(508)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(428),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(509)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(429),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(510)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(430),                                                                                                                                                                                             --                           .tx_parallel_data
			tx_parallel_data(511)     => xcvr_native_a10_0_unused_tx_parallel_data_unused_tx_parallel_data(431),                                                                                                                                                                                             --                           .tx_parallel_data
			rx_parallel_data(0)       => xcvr_native_a10_0_rx_parallel_data(0),                                                                                                                                                                                                                              --       rx_parallel_data_ch0.rx_parallel_data
			rx_parallel_data(1)       => xcvr_native_a10_0_rx_parallel_data(1),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(2)       => xcvr_native_a10_0_rx_parallel_data(2),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(3)       => xcvr_native_a10_0_rx_parallel_data(3),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(4)       => xcvr_native_a10_0_rx_parallel_data(4),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(5)       => xcvr_native_a10_0_rx_parallel_data(5),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(6)       => xcvr_native_a10_0_rx_parallel_data(6),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(7)       => xcvr_native_a10_0_rx_parallel_data(7),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(8)       => xcvr_native_a10_0_rx_parallel_data(8),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(9)       => xcvr_native_a10_0_rx_parallel_data(9),                                                                                                                                                                                                                              --                           .rx_parallel_data
			rx_parallel_data(10)      => xcvr_native_a10_0_rx_parallel_data(10),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(11)      => xcvr_native_a10_0_rx_parallel_data(11),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(12)      => xcvr_native_a10_0_rx_parallel_data(12),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(13)      => xcvr_native_a10_0_rx_parallel_data(13),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(14)      => xcvr_native_a10_0_rx_parallel_data(14),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(15)      => xcvr_native_a10_0_rx_parallel_data(15),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(16)      => xcvr_native_a10_0_rx_parallel_data(16),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(17)      => xcvr_native_a10_0_rx_parallel_data(17),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(18)      => xcvr_native_a10_0_rx_parallel_data(18),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(19)      => xcvr_native_a10_0_rx_parallel_data(19),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(20)      => xcvr_native_a10_0_rx_parallel_data(20),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(21)      => xcvr_native_a10_0_rx_parallel_data(21),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(22)      => xcvr_native_a10_0_rx_parallel_data(22),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(23)      => xcvr_native_a10_0_rx_parallel_data(23),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(24)      => xcvr_native_a10_0_rx_parallel_data(24),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(25)      => xcvr_native_a10_0_rx_parallel_data(25),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(26)      => xcvr_native_a10_0_rx_parallel_data(26),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(27)      => xcvr_native_a10_0_rx_parallel_data(27),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(28)      => xcvr_native_a10_0_rx_parallel_data(28),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(29)      => xcvr_native_a10_0_rx_parallel_data(29),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(30)      => xcvr_native_a10_0_rx_parallel_data(30),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(31)      => xcvr_native_a10_0_rx_parallel_data(31),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(32)      => xcvr_native_a10_0_rx_parallel_data(32),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(33)      => xcvr_native_a10_0_rx_parallel_data(33),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(34)      => xcvr_native_a10_0_rx_parallel_data(34),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(35)      => xcvr_native_a10_0_rx_parallel_data(35),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(36)      => xcvr_native_a10_0_rx_parallel_data(36),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(37)      => xcvr_native_a10_0_rx_parallel_data(37),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(38)      => xcvr_native_a10_0_rx_parallel_data(38),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(39)      => xcvr_native_a10_0_rx_parallel_data(39),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(40)      => xcvr_native_a10_0_rx_parallel_data(40),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(41)      => xcvr_native_a10_0_rx_parallel_data(41),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(42)      => xcvr_native_a10_0_rx_parallel_data(42),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(43)      => xcvr_native_a10_0_rx_parallel_data(43),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(44)      => xcvr_native_a10_0_rx_parallel_data(44),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(45)      => xcvr_native_a10_0_rx_parallel_data(45),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(46)      => xcvr_native_a10_0_rx_parallel_data(46),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(47)      => xcvr_native_a10_0_rx_parallel_data(47),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(48)      => xcvr_native_a10_0_rx_parallel_data(48),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(49)      => xcvr_native_a10_0_rx_parallel_data(49),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(50)      => xcvr_native_a10_0_rx_parallel_data(50),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(51)      => xcvr_native_a10_0_rx_parallel_data(51),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(52)      => xcvr_native_a10_0_rx_parallel_data(52),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(53)      => xcvr_native_a10_0_rx_parallel_data(53),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(54)      => xcvr_native_a10_0_rx_parallel_data(54),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(55)      => xcvr_native_a10_0_rx_parallel_data(55),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(56)      => xcvr_native_a10_0_rx_parallel_data(56),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(57)      => xcvr_native_a10_0_rx_parallel_data(57),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(58)      => xcvr_native_a10_0_rx_parallel_data(58),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(59)      => xcvr_native_a10_0_rx_parallel_data(59),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(60)      => xcvr_native_a10_0_rx_parallel_data(60),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(61)      => xcvr_native_a10_0_rx_parallel_data(61),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(62)      => xcvr_native_a10_0_rx_parallel_data(62),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(63)      => xcvr_native_a10_0_rx_parallel_data(63),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(64)      => xcvr_native_a10_0_rx_parallel_data(64),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(65)      => xcvr_native_a10_0_rx_parallel_data(65),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(66)      => xcvr_native_a10_0_rx_parallel_data(66),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(67)      => xcvr_native_a10_0_rx_parallel_data(67),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(68)      => xcvr_native_a10_0_rx_parallel_data(68),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(69)      => xcvr_native_a10_0_rx_parallel_data(69),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(70)      => xcvr_native_a10_0_rx_parallel_data(70),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(71)      => xcvr_native_a10_0_rx_parallel_data(71),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(72)      => xcvr_native_a10_0_rx_parallel_data(72),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(73)      => xcvr_native_a10_0_rx_parallel_data(73),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(74)      => xcvr_native_a10_0_rx_parallel_data(74),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(75)      => xcvr_native_a10_0_rx_parallel_data(75),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(76)      => xcvr_native_a10_0_rx_parallel_data(76),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(77)      => xcvr_native_a10_0_rx_parallel_data(77),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(78)      => xcvr_native_a10_0_rx_parallel_data(78),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(79)      => xcvr_native_a10_0_rx_parallel_data(79),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(80)      => xcvr_native_a10_0_rx_parallel_data(80),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(81)      => xcvr_native_a10_0_rx_parallel_data(81),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(82)      => xcvr_native_a10_0_rx_parallel_data(82),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(83)      => xcvr_native_a10_0_rx_parallel_data(83),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(84)      => xcvr_native_a10_0_rx_parallel_data(84),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(85)      => xcvr_native_a10_0_rx_parallel_data(85),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(86)      => xcvr_native_a10_0_rx_parallel_data(86),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(87)      => xcvr_native_a10_0_rx_parallel_data(87),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(88)      => xcvr_native_a10_0_rx_parallel_data(88),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(89)      => xcvr_native_a10_0_rx_parallel_data(89),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(90)      => xcvr_native_a10_0_rx_parallel_data(90),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(91)      => xcvr_native_a10_0_rx_parallel_data(91),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(92)      => xcvr_native_a10_0_rx_parallel_data(92),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(93)      => xcvr_native_a10_0_rx_parallel_data(93),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(94)      => xcvr_native_a10_0_rx_parallel_data(94),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(95)      => xcvr_native_a10_0_rx_parallel_data(95),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(96)      => xcvr_native_a10_0_rx_parallel_data(96),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(97)      => xcvr_native_a10_0_rx_parallel_data(97),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(98)      => xcvr_native_a10_0_rx_parallel_data(98),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(99)      => xcvr_native_a10_0_rx_parallel_data(99),                                                                                                                                                                                                                             --                           .rx_parallel_data
			rx_parallel_data(100)     => xcvr_native_a10_0_rx_parallel_data(100),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(101)     => xcvr_native_a10_0_rx_parallel_data(101),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(102)     => xcvr_native_a10_0_rx_parallel_data(102),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(103)     => xcvr_native_a10_0_rx_parallel_data(103),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(104)     => xcvr_native_a10_0_rx_parallel_data(104),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(105)     => xcvr_native_a10_0_rx_parallel_data(105),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(106)     => xcvr_native_a10_0_rx_parallel_data(106),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(107)     => xcvr_native_a10_0_rx_parallel_data(107),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(108)     => xcvr_native_a10_0_rx_parallel_data(108),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(109)     => xcvr_native_a10_0_rx_parallel_data(109),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(110)     => xcvr_native_a10_0_rx_parallel_data(110),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(111)     => xcvr_native_a10_0_rx_parallel_data(111),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(112)     => xcvr_native_a10_0_rx_parallel_data(112),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(113)     => xcvr_native_a10_0_rx_parallel_data(113),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(114)     => xcvr_native_a10_0_rx_parallel_data(114),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(115)     => xcvr_native_a10_0_rx_parallel_data(115),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(116)     => xcvr_native_a10_0_rx_parallel_data(116),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(117)     => xcvr_native_a10_0_rx_parallel_data(117),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(118)     => xcvr_native_a10_0_rx_parallel_data(118),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(119)     => xcvr_native_a10_0_rx_parallel_data(119),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(120)     => xcvr_native_a10_0_rx_parallel_data(120),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(121)     => xcvr_native_a10_0_rx_parallel_data(121),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(122)     => xcvr_native_a10_0_rx_parallel_data(122),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(123)     => xcvr_native_a10_0_rx_parallel_data(123),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(124)     => xcvr_native_a10_0_rx_parallel_data(124),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(125)     => xcvr_native_a10_0_rx_parallel_data(125),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(126)     => xcvr_native_a10_0_rx_parallel_data(126),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(127)     => xcvr_native_a10_0_rx_parallel_data(127),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(128)     => xcvr_native_a10_0_rx_parallel_data(128),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(129)     => xcvr_native_a10_0_rx_parallel_data(129),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(130)     => xcvr_native_a10_0_rx_parallel_data(130),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(131)     => xcvr_native_a10_0_rx_parallel_data(131),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(132)     => xcvr_native_a10_0_rx_parallel_data(132),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(133)     => xcvr_native_a10_0_rx_parallel_data(133),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(134)     => xcvr_native_a10_0_rx_parallel_data(134),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(135)     => xcvr_native_a10_0_rx_parallel_data(135),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(136)     => xcvr_native_a10_0_rx_parallel_data(136),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(137)     => xcvr_native_a10_0_rx_parallel_data(137),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(138)     => xcvr_native_a10_0_rx_parallel_data(138),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(139)     => xcvr_native_a10_0_rx_parallel_data(139),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(140)     => xcvr_native_a10_0_rx_parallel_data(140),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(141)     => xcvr_native_a10_0_rx_parallel_data(141),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(142)     => xcvr_native_a10_0_rx_parallel_data(142),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(143)     => xcvr_native_a10_0_rx_parallel_data(143),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(144)     => xcvr_native_a10_0_rx_parallel_data(144),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(145)     => xcvr_native_a10_0_rx_parallel_data(145),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(146)     => xcvr_native_a10_0_rx_parallel_data(146),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(147)     => xcvr_native_a10_0_rx_parallel_data(147),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(148)     => xcvr_native_a10_0_rx_parallel_data(148),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(149)     => xcvr_native_a10_0_rx_parallel_data(149),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(150)     => xcvr_native_a10_0_rx_parallel_data(150),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(151)     => xcvr_native_a10_0_rx_parallel_data(151),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(152)     => xcvr_native_a10_0_rx_parallel_data(152),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(153)     => xcvr_native_a10_0_rx_parallel_data(153),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(154)     => xcvr_native_a10_0_rx_parallel_data(154),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(155)     => xcvr_native_a10_0_rx_parallel_data(155),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(156)     => xcvr_native_a10_0_rx_parallel_data(156),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(157)     => xcvr_native_a10_0_rx_parallel_data(157),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(158)     => xcvr_native_a10_0_rx_parallel_data(158),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(159)     => xcvr_native_a10_0_rx_parallel_data(159),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(160)     => xcvr_native_a10_0_rx_parallel_data(160),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(161)     => xcvr_native_a10_0_rx_parallel_data(161),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(162)     => xcvr_native_a10_0_rx_parallel_data(162),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(163)     => xcvr_native_a10_0_rx_parallel_data(163),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(164)     => xcvr_native_a10_0_rx_parallel_data(164),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(165)     => xcvr_native_a10_0_rx_parallel_data(165),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(166)     => xcvr_native_a10_0_rx_parallel_data(166),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(167)     => xcvr_native_a10_0_rx_parallel_data(167),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(168)     => xcvr_native_a10_0_rx_parallel_data(168),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(169)     => xcvr_native_a10_0_rx_parallel_data(169),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(170)     => xcvr_native_a10_0_rx_parallel_data(170),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(171)     => xcvr_native_a10_0_rx_parallel_data(171),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(172)     => xcvr_native_a10_0_rx_parallel_data(172),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(173)     => xcvr_native_a10_0_rx_parallel_data(173),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(174)     => xcvr_native_a10_0_rx_parallel_data(174),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(175)     => xcvr_native_a10_0_rx_parallel_data(175),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(176)     => xcvr_native_a10_0_rx_parallel_data(176),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(177)     => xcvr_native_a10_0_rx_parallel_data(177),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(178)     => xcvr_native_a10_0_rx_parallel_data(178),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(179)     => xcvr_native_a10_0_rx_parallel_data(179),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(180)     => xcvr_native_a10_0_rx_parallel_data(180),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(181)     => xcvr_native_a10_0_rx_parallel_data(181),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(182)     => xcvr_native_a10_0_rx_parallel_data(182),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(183)     => xcvr_native_a10_0_rx_parallel_data(183),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(184)     => xcvr_native_a10_0_rx_parallel_data(184),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(185)     => xcvr_native_a10_0_rx_parallel_data(185),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(186)     => xcvr_native_a10_0_rx_parallel_data(186),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(187)     => xcvr_native_a10_0_rx_parallel_data(187),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(188)     => xcvr_native_a10_0_rx_parallel_data(188),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(189)     => xcvr_native_a10_0_rx_parallel_data(189),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(190)     => xcvr_native_a10_0_rx_parallel_data(190),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(191)     => xcvr_native_a10_0_rx_parallel_data(191),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(192)     => xcvr_native_a10_0_rx_parallel_data(192),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(193)     => xcvr_native_a10_0_rx_parallel_data(193),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(194)     => xcvr_native_a10_0_rx_parallel_data(194),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(195)     => xcvr_native_a10_0_rx_parallel_data(195),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(196)     => xcvr_native_a10_0_rx_parallel_data(196),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(197)     => xcvr_native_a10_0_rx_parallel_data(197),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(198)     => xcvr_native_a10_0_rx_parallel_data(198),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(199)     => xcvr_native_a10_0_rx_parallel_data(199),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(200)     => xcvr_native_a10_0_rx_parallel_data(200),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(201)     => xcvr_native_a10_0_rx_parallel_data(201),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(202)     => xcvr_native_a10_0_rx_parallel_data(202),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(203)     => xcvr_native_a10_0_rx_parallel_data(203),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(204)     => xcvr_native_a10_0_rx_parallel_data(204),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(205)     => xcvr_native_a10_0_rx_parallel_data(205),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(206)     => xcvr_native_a10_0_rx_parallel_data(206),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(207)     => xcvr_native_a10_0_rx_parallel_data(207),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(208)     => xcvr_native_a10_0_rx_parallel_data(208),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(209)     => xcvr_native_a10_0_rx_parallel_data(209),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(210)     => xcvr_native_a10_0_rx_parallel_data(210),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(211)     => xcvr_native_a10_0_rx_parallel_data(211),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(212)     => xcvr_native_a10_0_rx_parallel_data(212),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(213)     => xcvr_native_a10_0_rx_parallel_data(213),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(214)     => xcvr_native_a10_0_rx_parallel_data(214),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(215)     => xcvr_native_a10_0_rx_parallel_data(215),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(216)     => xcvr_native_a10_0_rx_parallel_data(216),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(217)     => xcvr_native_a10_0_rx_parallel_data(217),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(218)     => xcvr_native_a10_0_rx_parallel_data(218),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(219)     => xcvr_native_a10_0_rx_parallel_data(219),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(220)     => xcvr_native_a10_0_rx_parallel_data(220),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(221)     => xcvr_native_a10_0_rx_parallel_data(221),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(222)     => xcvr_native_a10_0_rx_parallel_data(222),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(223)     => xcvr_native_a10_0_rx_parallel_data(223),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(224)     => xcvr_native_a10_0_rx_parallel_data(224),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(225)     => xcvr_native_a10_0_rx_parallel_data(225),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(226)     => xcvr_native_a10_0_rx_parallel_data(226),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(227)     => xcvr_native_a10_0_rx_parallel_data(227),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(228)     => xcvr_native_a10_0_rx_parallel_data(228),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(229)     => xcvr_native_a10_0_rx_parallel_data(229),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(230)     => xcvr_native_a10_0_rx_parallel_data(230),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(231)     => xcvr_native_a10_0_rx_parallel_data(231),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(232)     => xcvr_native_a10_0_rx_parallel_data(232),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(233)     => xcvr_native_a10_0_rx_parallel_data(233),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(234)     => xcvr_native_a10_0_rx_parallel_data(234),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(235)     => xcvr_native_a10_0_rx_parallel_data(235),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(236)     => xcvr_native_a10_0_rx_parallel_data(236),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(237)     => xcvr_native_a10_0_rx_parallel_data(237),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(238)     => xcvr_native_a10_0_rx_parallel_data(238),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(239)     => xcvr_native_a10_0_rx_parallel_data(239),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(240)     => xcvr_native_a10_0_rx_parallel_data(240),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(241)     => xcvr_native_a10_0_rx_parallel_data(241),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(242)     => xcvr_native_a10_0_rx_parallel_data(242),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(243)     => xcvr_native_a10_0_rx_parallel_data(243),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(244)     => xcvr_native_a10_0_rx_parallel_data(244),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(245)     => xcvr_native_a10_0_rx_parallel_data(245),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(246)     => xcvr_native_a10_0_rx_parallel_data(246),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(247)     => xcvr_native_a10_0_rx_parallel_data(247),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(248)     => xcvr_native_a10_0_rx_parallel_data(248),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(249)     => xcvr_native_a10_0_rx_parallel_data(249),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(250)     => xcvr_native_a10_0_rx_parallel_data(250),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(251)     => xcvr_native_a10_0_rx_parallel_data(251),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(252)     => xcvr_native_a10_0_rx_parallel_data(252),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(253)     => xcvr_native_a10_0_rx_parallel_data(253),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(254)     => xcvr_native_a10_0_rx_parallel_data(254),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(255)     => xcvr_native_a10_0_rx_parallel_data(255),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(256)     => xcvr_native_a10_0_rx_parallel_data(256),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(257)     => xcvr_native_a10_0_rx_parallel_data(257),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(258)     => xcvr_native_a10_0_rx_parallel_data(258),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(259)     => xcvr_native_a10_0_rx_parallel_data(259),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(260)     => xcvr_native_a10_0_rx_parallel_data(260),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(261)     => xcvr_native_a10_0_rx_parallel_data(261),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(262)     => xcvr_native_a10_0_rx_parallel_data(262),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(263)     => xcvr_native_a10_0_rx_parallel_data(263),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(264)     => xcvr_native_a10_0_rx_parallel_data(264),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(265)     => xcvr_native_a10_0_rx_parallel_data(265),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(266)     => xcvr_native_a10_0_rx_parallel_data(266),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(267)     => xcvr_native_a10_0_rx_parallel_data(267),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(268)     => xcvr_native_a10_0_rx_parallel_data(268),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(269)     => xcvr_native_a10_0_rx_parallel_data(269),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(270)     => xcvr_native_a10_0_rx_parallel_data(270),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(271)     => xcvr_native_a10_0_rx_parallel_data(271),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(272)     => xcvr_native_a10_0_rx_parallel_data(272),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(273)     => xcvr_native_a10_0_rx_parallel_data(273),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(274)     => xcvr_native_a10_0_rx_parallel_data(274),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(275)     => xcvr_native_a10_0_rx_parallel_data(275),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(276)     => xcvr_native_a10_0_rx_parallel_data(276),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(277)     => xcvr_native_a10_0_rx_parallel_data(277),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(278)     => xcvr_native_a10_0_rx_parallel_data(278),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(279)     => xcvr_native_a10_0_rx_parallel_data(279),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(280)     => xcvr_native_a10_0_rx_parallel_data(280),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(281)     => xcvr_native_a10_0_rx_parallel_data(281),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(282)     => xcvr_native_a10_0_rx_parallel_data(282),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(283)     => xcvr_native_a10_0_rx_parallel_data(283),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(284)     => xcvr_native_a10_0_rx_parallel_data(284),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(285)     => xcvr_native_a10_0_rx_parallel_data(285),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(286)     => xcvr_native_a10_0_rx_parallel_data(286),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(287)     => xcvr_native_a10_0_rx_parallel_data(287),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(288)     => xcvr_native_a10_0_rx_parallel_data(288),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(289)     => xcvr_native_a10_0_rx_parallel_data(289),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(290)     => xcvr_native_a10_0_rx_parallel_data(290),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(291)     => xcvr_native_a10_0_rx_parallel_data(291),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(292)     => xcvr_native_a10_0_rx_parallel_data(292),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(293)     => xcvr_native_a10_0_rx_parallel_data(293),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(294)     => xcvr_native_a10_0_rx_parallel_data(294),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(295)     => xcvr_native_a10_0_rx_parallel_data(295),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(296)     => xcvr_native_a10_0_rx_parallel_data(296),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(297)     => xcvr_native_a10_0_rx_parallel_data(297),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(298)     => xcvr_native_a10_0_rx_parallel_data(298),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(299)     => xcvr_native_a10_0_rx_parallel_data(299),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(300)     => xcvr_native_a10_0_rx_parallel_data(300),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(301)     => xcvr_native_a10_0_rx_parallel_data(301),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(302)     => xcvr_native_a10_0_rx_parallel_data(302),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(303)     => xcvr_native_a10_0_rx_parallel_data(303),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(304)     => xcvr_native_a10_0_rx_parallel_data(304),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(305)     => xcvr_native_a10_0_rx_parallel_data(305),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(306)     => xcvr_native_a10_0_rx_parallel_data(306),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(307)     => xcvr_native_a10_0_rx_parallel_data(307),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(308)     => xcvr_native_a10_0_rx_parallel_data(308),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(309)     => xcvr_native_a10_0_rx_parallel_data(309),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(310)     => xcvr_native_a10_0_rx_parallel_data(310),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(311)     => xcvr_native_a10_0_rx_parallel_data(311),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(312)     => xcvr_native_a10_0_rx_parallel_data(312),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(313)     => xcvr_native_a10_0_rx_parallel_data(313),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(314)     => xcvr_native_a10_0_rx_parallel_data(314),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(315)     => xcvr_native_a10_0_rx_parallel_data(315),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(316)     => xcvr_native_a10_0_rx_parallel_data(316),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(317)     => xcvr_native_a10_0_rx_parallel_data(317),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(318)     => xcvr_native_a10_0_rx_parallel_data(318),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(319)     => xcvr_native_a10_0_rx_parallel_data(319),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(320)     => xcvr_native_a10_0_rx_parallel_data(320),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(321)     => xcvr_native_a10_0_rx_parallel_data(321),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(322)     => xcvr_native_a10_0_rx_parallel_data(322),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(323)     => xcvr_native_a10_0_rx_parallel_data(323),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(324)     => xcvr_native_a10_0_rx_parallel_data(324),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(325)     => xcvr_native_a10_0_rx_parallel_data(325),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(326)     => xcvr_native_a10_0_rx_parallel_data(326),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(327)     => xcvr_native_a10_0_rx_parallel_data(327),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(328)     => xcvr_native_a10_0_rx_parallel_data(328),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(329)     => xcvr_native_a10_0_rx_parallel_data(329),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(330)     => xcvr_native_a10_0_rx_parallel_data(330),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(331)     => xcvr_native_a10_0_rx_parallel_data(331),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(332)     => xcvr_native_a10_0_rx_parallel_data(332),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(333)     => xcvr_native_a10_0_rx_parallel_data(333),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(334)     => xcvr_native_a10_0_rx_parallel_data(334),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(335)     => xcvr_native_a10_0_rx_parallel_data(335),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(336)     => xcvr_native_a10_0_rx_parallel_data(336),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(337)     => xcvr_native_a10_0_rx_parallel_data(337),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(338)     => xcvr_native_a10_0_rx_parallel_data(338),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(339)     => xcvr_native_a10_0_rx_parallel_data(339),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(340)     => xcvr_native_a10_0_rx_parallel_data(340),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(341)     => xcvr_native_a10_0_rx_parallel_data(341),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(342)     => xcvr_native_a10_0_rx_parallel_data(342),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(343)     => xcvr_native_a10_0_rx_parallel_data(343),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(344)     => xcvr_native_a10_0_rx_parallel_data(344),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(345)     => xcvr_native_a10_0_rx_parallel_data(345),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(346)     => xcvr_native_a10_0_rx_parallel_data(346),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(347)     => xcvr_native_a10_0_rx_parallel_data(347),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(348)     => xcvr_native_a10_0_rx_parallel_data(348),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(349)     => xcvr_native_a10_0_rx_parallel_data(349),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(350)     => xcvr_native_a10_0_rx_parallel_data(350),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(351)     => xcvr_native_a10_0_rx_parallel_data(351),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(352)     => xcvr_native_a10_0_rx_parallel_data(352),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(353)     => xcvr_native_a10_0_rx_parallel_data(353),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(354)     => xcvr_native_a10_0_rx_parallel_data(354),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(355)     => xcvr_native_a10_0_rx_parallel_data(355),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(356)     => xcvr_native_a10_0_rx_parallel_data(356),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(357)     => xcvr_native_a10_0_rx_parallel_data(357),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(358)     => xcvr_native_a10_0_rx_parallel_data(358),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(359)     => xcvr_native_a10_0_rx_parallel_data(359),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(360)     => xcvr_native_a10_0_rx_parallel_data(360),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(361)     => xcvr_native_a10_0_rx_parallel_data(361),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(362)     => xcvr_native_a10_0_rx_parallel_data(362),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(363)     => xcvr_native_a10_0_rx_parallel_data(363),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(364)     => xcvr_native_a10_0_rx_parallel_data(364),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(365)     => xcvr_native_a10_0_rx_parallel_data(365),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(366)     => xcvr_native_a10_0_rx_parallel_data(366),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(367)     => xcvr_native_a10_0_rx_parallel_data(367),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(368)     => xcvr_native_a10_0_rx_parallel_data(368),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(369)     => xcvr_native_a10_0_rx_parallel_data(369),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(370)     => xcvr_native_a10_0_rx_parallel_data(370),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(371)     => xcvr_native_a10_0_rx_parallel_data(371),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(372)     => xcvr_native_a10_0_rx_parallel_data(372),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(373)     => xcvr_native_a10_0_rx_parallel_data(373),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(374)     => xcvr_native_a10_0_rx_parallel_data(374),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(375)     => xcvr_native_a10_0_rx_parallel_data(375),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(376)     => xcvr_native_a10_0_rx_parallel_data(376),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(377)     => xcvr_native_a10_0_rx_parallel_data(377),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(378)     => xcvr_native_a10_0_rx_parallel_data(378),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(379)     => xcvr_native_a10_0_rx_parallel_data(379),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(380)     => xcvr_native_a10_0_rx_parallel_data(380),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(381)     => xcvr_native_a10_0_rx_parallel_data(381),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(382)     => xcvr_native_a10_0_rx_parallel_data(382),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(383)     => xcvr_native_a10_0_rx_parallel_data(383),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(384)     => xcvr_native_a10_0_rx_parallel_data(384),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(385)     => xcvr_native_a10_0_rx_parallel_data(385),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(386)     => xcvr_native_a10_0_rx_parallel_data(386),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(387)     => xcvr_native_a10_0_rx_parallel_data(387),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(388)     => xcvr_native_a10_0_rx_parallel_data(388),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(389)     => xcvr_native_a10_0_rx_parallel_data(389),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(390)     => xcvr_native_a10_0_rx_parallel_data(390),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(391)     => xcvr_native_a10_0_rx_parallel_data(391),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(392)     => xcvr_native_a10_0_rx_parallel_data(392),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(393)     => xcvr_native_a10_0_rx_parallel_data(393),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(394)     => xcvr_native_a10_0_rx_parallel_data(394),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(395)     => xcvr_native_a10_0_rx_parallel_data(395),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(396)     => xcvr_native_a10_0_rx_parallel_data(396),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(397)     => xcvr_native_a10_0_rx_parallel_data(397),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(398)     => xcvr_native_a10_0_rx_parallel_data(398),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(399)     => xcvr_native_a10_0_rx_parallel_data(399),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(400)     => xcvr_native_a10_0_rx_parallel_data(400),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(401)     => xcvr_native_a10_0_rx_parallel_data(401),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(402)     => xcvr_native_a10_0_rx_parallel_data(402),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(403)     => xcvr_native_a10_0_rx_parallel_data(403),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(404)     => xcvr_native_a10_0_rx_parallel_data(404),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(405)     => xcvr_native_a10_0_rx_parallel_data(405),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(406)     => xcvr_native_a10_0_rx_parallel_data(406),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(407)     => xcvr_native_a10_0_rx_parallel_data(407),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(408)     => xcvr_native_a10_0_rx_parallel_data(408),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(409)     => xcvr_native_a10_0_rx_parallel_data(409),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(410)     => xcvr_native_a10_0_rx_parallel_data(410),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(411)     => xcvr_native_a10_0_rx_parallel_data(411),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(412)     => xcvr_native_a10_0_rx_parallel_data(412),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(413)     => xcvr_native_a10_0_rx_parallel_data(413),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(414)     => xcvr_native_a10_0_rx_parallel_data(414),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(415)     => xcvr_native_a10_0_rx_parallel_data(415),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(416)     => xcvr_native_a10_0_rx_parallel_data(416),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(417)     => xcvr_native_a10_0_rx_parallel_data(417),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(418)     => xcvr_native_a10_0_rx_parallel_data(418),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(419)     => xcvr_native_a10_0_rx_parallel_data(419),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(420)     => xcvr_native_a10_0_rx_parallel_data(420),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(421)     => xcvr_native_a10_0_rx_parallel_data(421),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(422)     => xcvr_native_a10_0_rx_parallel_data(422),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(423)     => xcvr_native_a10_0_rx_parallel_data(423),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(424)     => xcvr_native_a10_0_rx_parallel_data(424),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(425)     => xcvr_native_a10_0_rx_parallel_data(425),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(426)     => xcvr_native_a10_0_rx_parallel_data(426),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(427)     => xcvr_native_a10_0_rx_parallel_data(427),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(428)     => xcvr_native_a10_0_rx_parallel_data(428),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(429)     => xcvr_native_a10_0_rx_parallel_data(429),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(430)     => xcvr_native_a10_0_rx_parallel_data(430),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(431)     => xcvr_native_a10_0_rx_parallel_data(431),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(432)     => xcvr_native_a10_0_rx_parallel_data(432),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(433)     => xcvr_native_a10_0_rx_parallel_data(433),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(434)     => xcvr_native_a10_0_rx_parallel_data(434),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(435)     => xcvr_native_a10_0_rx_parallel_data(435),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(436)     => xcvr_native_a10_0_rx_parallel_data(436),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(437)     => xcvr_native_a10_0_rx_parallel_data(437),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(438)     => xcvr_native_a10_0_rx_parallel_data(438),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(439)     => xcvr_native_a10_0_rx_parallel_data(439),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(440)     => xcvr_native_a10_0_rx_parallel_data(440),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(441)     => xcvr_native_a10_0_rx_parallel_data(441),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(442)     => xcvr_native_a10_0_rx_parallel_data(442),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(443)     => xcvr_native_a10_0_rx_parallel_data(443),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(444)     => xcvr_native_a10_0_rx_parallel_data(444),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(445)     => xcvr_native_a10_0_rx_parallel_data(445),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(446)     => xcvr_native_a10_0_rx_parallel_data(446),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(447)     => xcvr_native_a10_0_rx_parallel_data(447),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(448)     => xcvr_native_a10_0_rx_parallel_data(448),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(449)     => xcvr_native_a10_0_rx_parallel_data(449),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(450)     => xcvr_native_a10_0_rx_parallel_data(450),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(451)     => xcvr_native_a10_0_rx_parallel_data(451),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(452)     => xcvr_native_a10_0_rx_parallel_data(452),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(453)     => xcvr_native_a10_0_rx_parallel_data(453),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(454)     => xcvr_native_a10_0_rx_parallel_data(454),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(455)     => xcvr_native_a10_0_rx_parallel_data(455),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(456)     => xcvr_native_a10_0_rx_parallel_data(456),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(457)     => xcvr_native_a10_0_rx_parallel_data(457),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(458)     => xcvr_native_a10_0_rx_parallel_data(458),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(459)     => xcvr_native_a10_0_rx_parallel_data(459),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(460)     => xcvr_native_a10_0_rx_parallel_data(460),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(461)     => xcvr_native_a10_0_rx_parallel_data(461),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(462)     => xcvr_native_a10_0_rx_parallel_data(462),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(463)     => xcvr_native_a10_0_rx_parallel_data(463),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(464)     => xcvr_native_a10_0_rx_parallel_data(464),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(465)     => xcvr_native_a10_0_rx_parallel_data(465),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(466)     => xcvr_native_a10_0_rx_parallel_data(466),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(467)     => xcvr_native_a10_0_rx_parallel_data(467),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(468)     => xcvr_native_a10_0_rx_parallel_data(468),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(469)     => xcvr_native_a10_0_rx_parallel_data(469),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(470)     => xcvr_native_a10_0_rx_parallel_data(470),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(471)     => xcvr_native_a10_0_rx_parallel_data(471),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(472)     => xcvr_native_a10_0_rx_parallel_data(472),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(473)     => xcvr_native_a10_0_rx_parallel_data(473),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(474)     => xcvr_native_a10_0_rx_parallel_data(474),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(475)     => xcvr_native_a10_0_rx_parallel_data(475),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(476)     => xcvr_native_a10_0_rx_parallel_data(476),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(477)     => xcvr_native_a10_0_rx_parallel_data(477),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(478)     => xcvr_native_a10_0_rx_parallel_data(478),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(479)     => xcvr_native_a10_0_rx_parallel_data(479),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(480)     => xcvr_native_a10_0_rx_parallel_data(480),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(481)     => xcvr_native_a10_0_rx_parallel_data(481),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(482)     => xcvr_native_a10_0_rx_parallel_data(482),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(483)     => xcvr_native_a10_0_rx_parallel_data(483),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(484)     => xcvr_native_a10_0_rx_parallel_data(484),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(485)     => xcvr_native_a10_0_rx_parallel_data(485),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(486)     => xcvr_native_a10_0_rx_parallel_data(486),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(487)     => xcvr_native_a10_0_rx_parallel_data(487),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(488)     => xcvr_native_a10_0_rx_parallel_data(488),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(489)     => xcvr_native_a10_0_rx_parallel_data(489),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(490)     => xcvr_native_a10_0_rx_parallel_data(490),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(491)     => xcvr_native_a10_0_rx_parallel_data(491),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(492)     => xcvr_native_a10_0_rx_parallel_data(492),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(493)     => xcvr_native_a10_0_rx_parallel_data(493),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(494)     => xcvr_native_a10_0_rx_parallel_data(494),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(495)     => xcvr_native_a10_0_rx_parallel_data(495),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(496)     => xcvr_native_a10_0_rx_parallel_data(496),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(497)     => xcvr_native_a10_0_rx_parallel_data(497),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(498)     => xcvr_native_a10_0_rx_parallel_data(498),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(499)     => xcvr_native_a10_0_rx_parallel_data(499),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(500)     => xcvr_native_a10_0_rx_parallel_data(500),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(501)     => xcvr_native_a10_0_rx_parallel_data(501),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(502)     => xcvr_native_a10_0_rx_parallel_data(502),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(503)     => xcvr_native_a10_0_rx_parallel_data(503),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(504)     => xcvr_native_a10_0_rx_parallel_data(504),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(505)     => xcvr_native_a10_0_rx_parallel_data(505),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(506)     => xcvr_native_a10_0_rx_parallel_data(506),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(507)     => xcvr_native_a10_0_rx_parallel_data(507),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(508)     => xcvr_native_a10_0_rx_parallel_data(508),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(509)     => xcvr_native_a10_0_rx_parallel_data(509),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(510)     => xcvr_native_a10_0_rx_parallel_data(510),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_parallel_data(511)     => xcvr_native_a10_0_rx_parallel_data(511),                                                                                                                                                                                                                            --                           .rx_parallel_data
			rx_std_wa_patternalign(0) => xcvr_native_a10_0_rx_std_wa_patternalign_ch0_rx_std_wa_patternalign,                                                                                                                                                                                                -- rx_std_wa_patternalign_ch0.rx_std_wa_patternalign
			rx_std_wa_patternalign(1) => xcvr_native_a10_0_rx_std_wa_patternalign_ch1_rx_std_wa_patternalign,                                                                                                                                                                                                --                           .rx_std_wa_patternalign
			rx_std_wa_patternalign(2) => xcvr_native_a10_0_rx_std_wa_patternalign_ch2_rx_std_wa_patternalign,                                                                                                                                                                                                --                           .rx_std_wa_patternalign
			rx_std_wa_patternalign(3) => xcvr_native_a10_0_rx_std_wa_patternalign_ch3_rx_std_wa_patternalign,                                                                                                                                                                                                --                           .rx_std_wa_patternalign
			tx_analogreset_ack        => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_analogreset_ack        => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_serial_clk1            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_serial_clk2            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_serial_clk3            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_bonding_clocks         => "000000000000000000000000",                                                                                                                                                                                                                                         --                (terminated)
			tx_bonding_clocks1        => "000000000000000000000000",                                                                                                                                                                                                                                         --                (terminated)
			tx_bonding_clocks2        => "000000000000000000000000",                                                                                                                                                                                                                                         --                (terminated)
			tx_bonding_clocks3        => "000000000000000000000000",                                                                                                                                                                                                                                         --                (terminated)
			rx_cdr_refclk1            => '0',                                                                                                                                                                                                                                                                --                (terminated)
			rx_cdr_refclk2            => '0',                                                                                                                                                                                                                                                                --                (terminated)
			rx_cdr_refclk3            => '0',                                                                                                                                                                                                                                                                --                (terminated)
			rx_cdr_refclk4            => '0',                                                                                                                                                                                                                                                                --                (terminated)
			rx_pma_clkslip            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_set_locktodata         => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_set_locktoref          => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_is_lockedtoref         => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_pma_qpipulldn          => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_pma_qpipulldn          => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_pma_qpipullup          => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_pma_txdetectrx         => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_pma_elecidle           => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_pma_rxfound            => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_clklow                 => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_fref                   => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_pma_clkout             => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_pma_div_clkout         => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_pma_iqtxrx_clkout      => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_pma_clkout             => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_pma_div_clkout         => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_pma_iqtxrx_clkout      => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_control                => "000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                                                         --                (terminated)
			rx_control                => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_bitslip                => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_adapt_reset            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_adapt_start            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_prbs_err_clr           => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_prbs_done              => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_prbs_err               => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_uhsif_clk              => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_uhsif_clkout           => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_uhsif_lock             => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_std_pcfifo_full        => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_std_pcfifo_empty       => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_std_bitrev_ena         => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_std_byterev_ena        => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_polinv                 => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_polinv                 => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_std_bitslipboundarysel => "00000000000000000000",                                                                                                                                                                                                                                             --                (terminated)
			rx_std_bitslipboundarysel => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_std_wa_a1a2size        => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_std_rmfifo_full        => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_std_rmfifo_empty       => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_std_signaldetect       => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_data_valid         => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_enh_fifo_full          => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_fifo_pfull         => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_fifo_empty         => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_fifo_pempty        => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_fifo_cnt           => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_rd_en         => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_enh_data_valid         => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_full          => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_pfull         => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_empty         => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_pempty        => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_del           => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_insert        => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_cnt           => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_align_val     => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_fifo_align_clr     => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_enh_frame              => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_frame_burst_en     => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			tx_enh_frame_diag_status  => "00000000",                                                                                                                                                                                                                                                         --                (terminated)
			rx_enh_frame              => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_frame_lock         => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_frame_diag_status  => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_crc32_err          => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_highber            => open,                                                                                                                                                                                                                                                               --                (terminated)
			rx_enh_highber_clr_cnt    => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_enh_clr_errblk_count   => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			rx_enh_blk_lock           => open,                                                                                                                                                                                                                                                               --                (terminated)
			tx_enh_bitslip            => "0000000000000000000000000000",                                                                                                                                                                                                                                     --                (terminated)
			tx_hip_data               => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", --                (terminated)
			rx_hip_data               => open,                                                                                                                                                                                                                                                               --                (terminated)
			hip_pipe_pclk             => open,                                                                                                                                                                                                                                                               --                (terminated)
			hip_fixedclk              => open,                                                                                                                                                                                                                                                               --                (terminated)
			hip_frefclk               => open,                                                                                                                                                                                                                                                               --                (terminated)
			hip_ctrl                  => open,                                                                                                                                                                                                                                                               --                (terminated)
			hip_cal_done              => open,                                                                                                                                                                                                                                                               --                (terminated)
			ltssm_detect_quiet        => '0',                                                                                                                                                                                                                                                                --                (terminated)
			ltssm_detect_active       => '0',                                                                                                                                                                                                                                                                --                (terminated)
			ltssm_rcvr_phase_two      => '0',                                                                                                                                                                                                                                                                --                (terminated)
			hip_reduce_counters       => '0',                                                                                                                                                                                                                                                                --                (terminated)
			pcie_rate                 => "00",                                                                                                                                                                                                                                                               --                (terminated)
			pipe_rate                 => "00",                                                                                                                                                                                                                                                               --                (terminated)
			pipe_sw_done              => "00",                                                                                                                                                                                                                                                               --                (terminated)
			pipe_sw                   => open,                                                                                                                                                                                                                                                               --                (terminated)
			pipe_hclk_in              => '0',                                                                                                                                                                                                                                                                --                (terminated)
			pipe_hclk_out             => open,                                                                                                                                                                                                                                                               --                (terminated)
			pipe_g3_txdeemph          => "000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                                                                         --                (terminated)
			pipe_g3_rxpresethint      => "000000000000",                                                                                                                                                                                                                                                     --                (terminated)
			pipe_rx_eidleinfersel     => "000000000000",                                                                                                                                                                                                                                                     --                (terminated)
			pipe_rx_elecidle          => open,                                                                                                                                                                                                                                                               --                (terminated)
			pipe_rx_polarity          => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			reconfig_clk              => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			reconfig_reset            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			reconfig_write            => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			reconfig_read             => "0000",                                                                                                                                                                                                                                                             --                (terminated)
			reconfig_address          => "0000000000000000000000000000000000000000",                                                                                                                                                                                                                         --                (terminated)
			reconfig_writedata        => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",                                                                                                                                 --                (terminated)
			reconfig_readdata         => open,                                                                                                                                                                                                                                                               --                (terminated)
			reconfig_waitrequest      => open,                                                                                                                                                                                                                                                               --                (terminated)
			avmm_busy                 => open                                                                                                                                                                                                                                                                --                (terminated)
		);

	xcvr_reset_control_0 : component altera_xcvr_reset_control
		generic map (
			CHANNELS              => 4,
			PLLS                  => 1,
			SYS_CLK_IN_MHZ        => 127,
			SYNCHRONIZE_RESET     => 1,
			REDUCED_SIM_TIME      => 1,
			TX_PLL_ENABLE         => 1,
			T_PLL_POWERDOWN       => 1000,
			SYNCHRONIZE_PLL_RESET => 0,
			TX_ENABLE             => 1,
			TX_PER_CHANNEL        => 0,
			T_TX_ANALOGRESET      => 70000,
			T_TX_DIGITALRESET     => 70000,
			T_PLL_LOCK_HYST       => 0,
			EN_PLL_CAL_BUSY       => 1,
			RX_ENABLE             => 1,
			RX_PER_CHANNEL        => 0,
			T_RX_ANALOGRESET      => 70000,
			T_RX_DIGITALRESET     => 4000
		)
		port map (
			clock                 => xcvr_reset_control_0_clock_clk,                              --               clock.clk
			reset                 => xcvr_reset_control_0_reset_reset,                            --               reset.reset
			pll_powerdown(0)      => xcvr_reset_control_0_pll_powerdown(0),                       --      pll_powerdown0.pll_powerdown
			tx_analogreset(0)     => xcvr_reset_control_0_tx_analogreset(0),                      --     tx_analogreset0.tx_analogreset
			tx_analogreset(1)     => xcvr_reset_control_0_tx_analogreset(1),                      --                    .tx_analogreset
			tx_analogreset(2)     => xcvr_reset_control_0_tx_analogreset(2),                      --                    .tx_analogreset
			tx_analogreset(3)     => xcvr_reset_control_0_tx_analogreset(3),                      --                    .tx_analogreset
			tx_digitalreset(0)    => xcvr_reset_control_0_tx_digitalreset(0),                     --    tx_digitalreset0.tx_digitalreset
			tx_digitalreset(1)    => xcvr_reset_control_0_tx_digitalreset(1),                     --                    .tx_digitalreset
			tx_digitalreset(2)    => xcvr_reset_control_0_tx_digitalreset(2),                     --                    .tx_digitalreset
			tx_digitalreset(3)    => xcvr_reset_control_0_tx_digitalreset(3),                     --                    .tx_digitalreset
			tx_ready(0)           => xcvr_reset_control_0_tx_ready(0),                            --           tx_ready0.tx_ready
			tx_ready(1)           => xcvr_reset_control_0_tx_ready(1),                            --                    .tx_ready
			tx_ready(2)           => xcvr_reset_control_0_tx_ready(2),                            --                    .tx_ready
			tx_ready(3)           => xcvr_reset_control_0_tx_ready(3),                            --                    .tx_ready
			pll_locked(0)         => xcvr_atx_pll_a10_0_pll_locked_pll_locked,                    --         pll_locked0.pll_locked
			pll_select            => xcvr_reset_control_0_pll_select_pll_select,                  --          pll_select.pll_select
			tx_cal_busy(0)        => xcvr_native_a10_0_tx_cal_busy_ch0_tx_cal_busy,               --        tx_cal_busy0.tx_cal_busy
			tx_cal_busy(1)        => xcvr_native_a10_0_tx_cal_busy_ch1_tx_cal_busy,               --                    .tx_cal_busy
			tx_cal_busy(2)        => xcvr_native_a10_0_tx_cal_busy_ch2_tx_cal_busy,               --                    .tx_cal_busy
			tx_cal_busy(3)        => xcvr_native_a10_0_tx_cal_busy_ch3_tx_cal_busy,               --                    .tx_cal_busy
			pll_cal_busy(0)       => xcvr_atx_pll_a10_0_pll_cal_busy_pll_cal_busy,                --       pll_cal_busy0.pll_cal_busy
			rx_analogreset(0)     => xcvr_reset_control_0_rx_analogreset(0),                      --     rx_analogreset0.rx_analogreset
			rx_analogreset(1)     => xcvr_reset_control_0_rx_analogreset(1),                      --                    .rx_analogreset
			rx_analogreset(2)     => xcvr_reset_control_0_rx_analogreset(2),                      --                    .rx_analogreset
			rx_analogreset(3)     => xcvr_reset_control_0_rx_analogreset(3),                      --                    .rx_analogreset
			rx_digitalreset(0)    => xcvr_reset_control_0_rx_digitalreset(0),                     --    rx_digitalreset0.rx_digitalreset
			rx_digitalreset(1)    => xcvr_reset_control_0_rx_digitalreset(1),                     --                    .rx_digitalreset
			rx_digitalreset(2)    => xcvr_reset_control_0_rx_digitalreset(2),                     --                    .rx_digitalreset
			rx_digitalreset(3)    => xcvr_reset_control_0_rx_digitalreset(3),                     --                    .rx_digitalreset
			rx_ready(0)           => xcvr_reset_control_0_rx_ready(0),                            --           rx_ready0.rx_ready
			rx_ready(1)           => xcvr_reset_control_0_rx_ready(1),                            --                    .rx_ready
			rx_ready(2)           => xcvr_reset_control_0_rx_ready(2),                            --                    .rx_ready
			rx_ready(3)           => xcvr_reset_control_0_rx_ready(3),                            --                    .rx_ready
			rx_is_lockedtodata(0) => xcvr_native_a10_0_rx_is_lockedtodata_ch0_rx_is_lockedtodata, -- rx_is_lockedtodata0.rx_is_lockedtodata
			rx_is_lockedtodata(1) => xcvr_native_a10_0_rx_is_lockedtodata_ch1_rx_is_lockedtodata, --                    .rx_is_lockedtodata
			rx_is_lockedtodata(2) => xcvr_native_a10_0_rx_is_lockedtodata_ch2_rx_is_lockedtodata, --                    .rx_is_lockedtodata
			rx_is_lockedtodata(3) => xcvr_native_a10_0_rx_is_lockedtodata_ch3_rx_is_lockedtodata, --                    .rx_is_lockedtodata
			rx_cal_busy(0)        => xcvr_native_a10_0_rx_cal_busy_ch0_rx_cal_busy,               --        rx_cal_busy0.rx_cal_busy
			rx_cal_busy(1)        => xcvr_native_a10_0_rx_cal_busy_ch1_rx_cal_busy,               --                    .rx_cal_busy
			rx_cal_busy(2)        => xcvr_native_a10_0_rx_cal_busy_ch2_rx_cal_busy,               --                    .rx_cal_busy
			rx_cal_busy(3)        => xcvr_native_a10_0_rx_cal_busy_ch3_rx_cal_busy,               --                    .rx_cal_busy
			tx_manual             => "0000",                                                      --         (terminated)
			rx_manual             => "0000",                                                      --         (terminated)
			tx_digitalreset_or    => "0000",                                                      --         (terminated)
			rx_digitalreset_or    => "0000"                                                       --         (terminated)
		);

	xcvr_native_a10_0_rx_clkout_ch0_clk <= xcvr_native_a10_0_rx_clkout(0);

	xcvr_native_a10_0_rx_clkout_ch1_clk <= xcvr_native_a10_0_rx_clkout(1);

	xcvr_native_a10_0_rx_clkout_ch2_clk <= xcvr_native_a10_0_rx_clkout(2);

	xcvr_native_a10_0_rx_clkout_ch3_clk <= xcvr_native_a10_0_rx_clkout(3);

	xcvr_native_a10_0_rx_parallel_data_ch0_rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(25) & xcvr_native_a10_0_rx_parallel_data(24) & xcvr_native_a10_0_rx_parallel_data(23) & xcvr_native_a10_0_rx_parallel_data(22) & xcvr_native_a10_0_rx_parallel_data(21) & xcvr_native_a10_0_rx_parallel_data(20) & xcvr_native_a10_0_rx_parallel_data(19) & xcvr_native_a10_0_rx_parallel_data(18) & xcvr_native_a10_0_rx_parallel_data(17) & xcvr_native_a10_0_rx_parallel_data(16) & xcvr_native_a10_0_rx_parallel_data(9) & xcvr_native_a10_0_rx_parallel_data(8) & xcvr_native_a10_0_rx_parallel_data(7) & xcvr_native_a10_0_rx_parallel_data(6) & xcvr_native_a10_0_rx_parallel_data(5) & xcvr_native_a10_0_rx_parallel_data(4) & xcvr_native_a10_0_rx_parallel_data(3) & xcvr_native_a10_0_rx_parallel_data(2) & xcvr_native_a10_0_rx_parallel_data(1) & xcvr_native_a10_0_rx_parallel_data(0);

	xcvr_native_a10_0_rx_parallel_data_ch1_rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(153) & xcvr_native_a10_0_rx_parallel_data(152) & xcvr_native_a10_0_rx_parallel_data(151) & xcvr_native_a10_0_rx_parallel_data(150) & xcvr_native_a10_0_rx_parallel_data(149) & xcvr_native_a10_0_rx_parallel_data(148) & xcvr_native_a10_0_rx_parallel_data(147) & xcvr_native_a10_0_rx_parallel_data(146) & xcvr_native_a10_0_rx_parallel_data(145) & xcvr_native_a10_0_rx_parallel_data(144) & xcvr_native_a10_0_rx_parallel_data(137) & xcvr_native_a10_0_rx_parallel_data(136) & xcvr_native_a10_0_rx_parallel_data(135) & xcvr_native_a10_0_rx_parallel_data(134) & xcvr_native_a10_0_rx_parallel_data(133) & xcvr_native_a10_0_rx_parallel_data(132) & xcvr_native_a10_0_rx_parallel_data(131) & xcvr_native_a10_0_rx_parallel_data(130) & xcvr_native_a10_0_rx_parallel_data(129) & xcvr_native_a10_0_rx_parallel_data(128);

	xcvr_native_a10_0_rx_parallel_data_ch2_rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(281) & xcvr_native_a10_0_rx_parallel_data(280) & xcvr_native_a10_0_rx_parallel_data(279) & xcvr_native_a10_0_rx_parallel_data(278) & xcvr_native_a10_0_rx_parallel_data(277) & xcvr_native_a10_0_rx_parallel_data(276) & xcvr_native_a10_0_rx_parallel_data(275) & xcvr_native_a10_0_rx_parallel_data(274) & xcvr_native_a10_0_rx_parallel_data(273) & xcvr_native_a10_0_rx_parallel_data(272) & xcvr_native_a10_0_rx_parallel_data(265) & xcvr_native_a10_0_rx_parallel_data(264) & xcvr_native_a10_0_rx_parallel_data(263) & xcvr_native_a10_0_rx_parallel_data(262) & xcvr_native_a10_0_rx_parallel_data(261) & xcvr_native_a10_0_rx_parallel_data(260) & xcvr_native_a10_0_rx_parallel_data(259) & xcvr_native_a10_0_rx_parallel_data(258) & xcvr_native_a10_0_rx_parallel_data(257) & xcvr_native_a10_0_rx_parallel_data(256);

	xcvr_native_a10_0_rx_parallel_data_ch3_rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(409) & xcvr_native_a10_0_rx_parallel_data(408) & xcvr_native_a10_0_rx_parallel_data(407) & xcvr_native_a10_0_rx_parallel_data(406) & xcvr_native_a10_0_rx_parallel_data(405) & xcvr_native_a10_0_rx_parallel_data(404) & xcvr_native_a10_0_rx_parallel_data(403) & xcvr_native_a10_0_rx_parallel_data(402) & xcvr_native_a10_0_rx_parallel_data(401) & xcvr_native_a10_0_rx_parallel_data(400) & xcvr_native_a10_0_rx_parallel_data(393) & xcvr_native_a10_0_rx_parallel_data(392) & xcvr_native_a10_0_rx_parallel_data(391) & xcvr_native_a10_0_rx_parallel_data(390) & xcvr_native_a10_0_rx_parallel_data(389) & xcvr_native_a10_0_rx_parallel_data(388) & xcvr_native_a10_0_rx_parallel_data(387) & xcvr_native_a10_0_rx_parallel_data(386) & xcvr_native_a10_0_rx_parallel_data(385) & xcvr_native_a10_0_rx_parallel_data(384);

	xcvr_native_a10_0_rx_patterndetect_ch0_rx_patterndetect <= xcvr_native_a10_0_rx_parallel_data(28) & xcvr_native_a10_0_rx_parallel_data(12);

	xcvr_native_a10_0_rx_patterndetect_ch1_rx_patterndetect <= xcvr_native_a10_0_rx_parallel_data(156) & xcvr_native_a10_0_rx_parallel_data(140);

	xcvr_native_a10_0_rx_patterndetect_ch2_rx_patterndetect <= xcvr_native_a10_0_rx_parallel_data(284) & xcvr_native_a10_0_rx_parallel_data(268);

	xcvr_native_a10_0_rx_patterndetect_ch3_rx_patterndetect <= xcvr_native_a10_0_rx_parallel_data(412) & xcvr_native_a10_0_rx_parallel_data(396);

	xcvr_native_a10_0_rx_syncstatus_ch0_rx_syncstatus <= xcvr_native_a10_0_rx_parallel_data(26) & xcvr_native_a10_0_rx_parallel_data(10);

	xcvr_native_a10_0_rx_syncstatus_ch1_rx_syncstatus <= xcvr_native_a10_0_rx_parallel_data(154) & xcvr_native_a10_0_rx_parallel_data(138);

	xcvr_native_a10_0_rx_syncstatus_ch2_rx_syncstatus <= xcvr_native_a10_0_rx_parallel_data(282) & xcvr_native_a10_0_rx_parallel_data(266);

	xcvr_native_a10_0_rx_syncstatus_ch3_rx_syncstatus <= xcvr_native_a10_0_rx_parallel_data(410) & xcvr_native_a10_0_rx_parallel_data(394);

	xcvr_native_a10_0_tx_clkout_ch0_clk <= xcvr_native_a10_0_tx_clkout(0);

	xcvr_native_a10_0_tx_clkout_ch1_clk <= xcvr_native_a10_0_tx_clkout(1);

	xcvr_native_a10_0_tx_clkout_ch2_clk <= xcvr_native_a10_0_tx_clkout(2);

	xcvr_native_a10_0_tx_clkout_ch3_clk <= xcvr_native_a10_0_tx_clkout(3);

	xcvr_native_a10_0_tx_serial_data_ch0_tx_serial_data <= xcvr_native_a10_0_tx_serial_data(0);

	xcvr_native_a10_0_tx_serial_data_ch1_tx_serial_data <= xcvr_native_a10_0_tx_serial_data(1);

	xcvr_native_a10_0_tx_serial_data_ch2_tx_serial_data <= xcvr_native_a10_0_tx_serial_data(2);

	xcvr_native_a10_0_tx_serial_data_ch3_tx_serial_data <= xcvr_native_a10_0_tx_serial_data(3);

	xcvr_native_a10_0_unused_rx_parallel_data_unused_rx_parallel_data <= xcvr_native_a10_0_rx_parallel_data(511) & xcvr_native_a10_0_rx_parallel_data(510) & xcvr_native_a10_0_rx_parallel_data(509) & xcvr_native_a10_0_rx_parallel_data(508) & xcvr_native_a10_0_rx_parallel_data(507) & xcvr_native_a10_0_rx_parallel_data(506) & xcvr_native_a10_0_rx_parallel_data(505) & xcvr_native_a10_0_rx_parallel_data(504) & xcvr_native_a10_0_rx_parallel_data(503) & xcvr_native_a10_0_rx_parallel_data(502) & xcvr_native_a10_0_rx_parallel_data(501) & xcvr_native_a10_0_rx_parallel_data(500) & xcvr_native_a10_0_rx_parallel_data(499) & xcvr_native_a10_0_rx_parallel_data(498) & xcvr_native_a10_0_rx_parallel_data(497) & xcvr_native_a10_0_rx_parallel_data(496) & xcvr_native_a10_0_rx_parallel_data(495) & xcvr_native_a10_0_rx_parallel_data(494) & xcvr_native_a10_0_rx_parallel_data(493) & xcvr_native_a10_0_rx_parallel_data(492) & xcvr_native_a10_0_rx_parallel_data(491) & xcvr_native_a10_0_rx_parallel_data(490) & xcvr_native_a10_0_rx_parallel_data(489) & xcvr_native_a10_0_rx_parallel_data(488) & xcvr_native_a10_0_rx_parallel_data(487) & xcvr_native_a10_0_rx_parallel_data(486) & xcvr_native_a10_0_rx_parallel_data(485) & xcvr_native_a10_0_rx_parallel_data(484) & xcvr_native_a10_0_rx_parallel_data(483) & xcvr_native_a10_0_rx_parallel_data(482) & xcvr_native_a10_0_rx_parallel_data(481) & xcvr_native_a10_0_rx_parallel_data(480) & xcvr_native_a10_0_rx_parallel_data(479) & xcvr_native_a10_0_rx_parallel_data(478) & xcvr_native_a10_0_rx_parallel_data(477) & xcvr_native_a10_0_rx_parallel_data(476) & xcvr_native_a10_0_rx_parallel_data(475) & xcvr_native_a10_0_rx_parallel_data(474) & xcvr_native_a10_0_rx_parallel_data(473) & xcvr_native_a10_0_rx_parallel_data(472) & xcvr_native_a10_0_rx_parallel_data(471) & xcvr_native_a10_0_rx_parallel_data(470) & xcvr_native_a10_0_rx_parallel_data(469) & xcvr_native_a10_0_rx_parallel_data(468) & xcvr_native_a10_0_rx_parallel_data(467) & xcvr_native_a10_0_rx_parallel_data(466) & xcvr_native_a10_0_rx_parallel_data(465) & xcvr_native_a10_0_rx_parallel_data(464) & xcvr_native_a10_0_rx_parallel_data(463) & xcvr_native_a10_0_rx_parallel_data(462) & xcvr_native_a10_0_rx_parallel_data(461) & xcvr_native_a10_0_rx_parallel_data(460) & xcvr_native_a10_0_rx_parallel_data(459) & xcvr_native_a10_0_rx_parallel_data(458) & xcvr_native_a10_0_rx_parallel_data(457) & xcvr_native_a10_0_rx_parallel_data(456) & xcvr_native_a10_0_rx_parallel_data(455) & xcvr_native_a10_0_rx_parallel_data(454) & xcvr_native_a10_0_rx_parallel_data(453) & xcvr_native_a10_0_rx_parallel_data(452) & xcvr_native_a10_0_rx_parallel_data(451) & xcvr_native_a10_0_rx_parallel_data(450) & xcvr_native_a10_0_rx_parallel_data(449) & xcvr_native_a10_0_rx_parallel_data(448) & xcvr_native_a10_0_rx_parallel_data(447) & xcvr_native_a10_0_rx_parallel_data(446) & xcvr_native_a10_0_rx_parallel_data(445) & xcvr_native_a10_0_rx_parallel_data(444) & xcvr_native_a10_0_rx_parallel_data(443) & xcvr_native_a10_0_rx_parallel_data(442) & xcvr_native_a10_0_rx_parallel_data(441) & xcvr_native_a10_0_rx_parallel_data(440) & xcvr_native_a10_0_rx_parallel_data(439) & xcvr_native_a10_0_rx_parallel_data(438) & xcvr_native_a10_0_rx_parallel_data(437) & xcvr_native_a10_0_rx_parallel_data(436) & xcvr_native_a10_0_rx_parallel_data(435) & xcvr_native_a10_0_rx_parallel_data(434) & xcvr_native_a10_0_rx_parallel_data(433) & xcvr_native_a10_0_rx_parallel_data(432) & xcvr_native_a10_0_rx_parallel_data(431) & xcvr_native_a10_0_rx_parallel_data(430) & xcvr_native_a10_0_rx_parallel_data(429) & xcvr_native_a10_0_rx_parallel_data(428) & xcvr_native_a10_0_rx_parallel_data(427) & xcvr_native_a10_0_rx_parallel_data(426) & xcvr_native_a10_0_rx_parallel_data(425) & xcvr_native_a10_0_rx_parallel_data(424) & xcvr_native_a10_0_rx_parallel_data(423) & xcvr_native_a10_0_rx_parallel_data(422) & xcvr_native_a10_0_rx_parallel_data(421) & xcvr_native_a10_0_rx_parallel_data(420) & xcvr_native_a10_0_rx_parallel_data(419) & xcvr_native_a10_0_rx_parallel_data(418) & xcvr_native_a10_0_rx_parallel_data(417) & xcvr_native_a10_0_rx_parallel_data(416) & xcvr_native_a10_0_rx_parallel_data(415) & xcvr_native_a10_0_rx_parallel_data(414) & xcvr_native_a10_0_rx_parallel_data(413) & xcvr_native_a10_0_rx_parallel_data(411) & xcvr_native_a10_0_rx_parallel_data(399) & xcvr_native_a10_0_rx_parallel_data(398) & xcvr_native_a10_0_rx_parallel_data(397) & xcvr_native_a10_0_rx_parallel_data(395) & xcvr_native_a10_0_rx_parallel_data(383) & xcvr_native_a10_0_rx_parallel_data(382) & xcvr_native_a10_0_rx_parallel_data(381) & xcvr_native_a10_0_rx_parallel_data(380) & xcvr_native_a10_0_rx_parallel_data(379) & xcvr_native_a10_0_rx_parallel_data(378) & xcvr_native_a10_0_rx_parallel_data(377) & xcvr_native_a10_0_rx_parallel_data(376) & xcvr_native_a10_0_rx_parallel_data(375) & xcvr_native_a10_0_rx_parallel_data(374) & xcvr_native_a10_0_rx_parallel_data(373) & xcvr_native_a10_0_rx_parallel_data(372) & xcvr_native_a10_0_rx_parallel_data(371) & xcvr_native_a10_0_rx_parallel_data(370) & xcvr_native_a10_0_rx_parallel_data(369) & xcvr_native_a10_0_rx_parallel_data(368) & xcvr_native_a10_0_rx_parallel_data(367) & xcvr_native_a10_0_rx_parallel_data(366) & xcvr_native_a10_0_rx_parallel_data(365) & xcvr_native_a10_0_rx_parallel_data(364) & xcvr_native_a10_0_rx_parallel_data(363) & xcvr_native_a10_0_rx_parallel_data(362) & xcvr_native_a10_0_rx_parallel_data(361) & xcvr_native_a10_0_rx_parallel_data(360) & xcvr_native_a10_0_rx_parallel_data(359) & xcvr_native_a10_0_rx_parallel_data(358) & xcvr_native_a10_0_rx_parallel_data(357) & xcvr_native_a10_0_rx_parallel_data(356) & xcvr_native_a10_0_rx_parallel_data(355) & xcvr_native_a10_0_rx_parallel_data(354) & xcvr_native_a10_0_rx_parallel_data(353) & xcvr_native_a10_0_rx_parallel_data(352) & xcvr_native_a10_0_rx_parallel_data(351) & xcvr_native_a10_0_rx_parallel_data(350) & xcvr_native_a10_0_rx_parallel_data(349) & xcvr_native_a10_0_rx_parallel_data(348) & xcvr_native_a10_0_rx_parallel_data(347) & xcvr_native_a10_0_rx_parallel_data(346) & xcvr_native_a10_0_rx_parallel_data(345) & xcvr_native_a10_0_rx_parallel_data(344) & xcvr_native_a10_0_rx_parallel_data(343) & xcvr_native_a10_0_rx_parallel_data(342) & xcvr_native_a10_0_rx_parallel_data(341) & xcvr_native_a10_0_rx_parallel_data(340) & xcvr_native_a10_0_rx_parallel_data(339) & xcvr_native_a10_0_rx_parallel_data(338) & xcvr_native_a10_0_rx_parallel_data(337) & xcvr_native_a10_0_rx_parallel_data(336) & xcvr_native_a10_0_rx_parallel_data(335) & xcvr_native_a10_0_rx_parallel_data(334) & xcvr_native_a10_0_rx_parallel_data(333) & xcvr_native_a10_0_rx_parallel_data(332) & xcvr_native_a10_0_rx_parallel_data(331) & xcvr_native_a10_0_rx_parallel_data(330) & xcvr_native_a10_0_rx_parallel_data(329) & xcvr_native_a10_0_rx_parallel_data(328) & xcvr_native_a10_0_rx_parallel_data(327) & xcvr_native_a10_0_rx_parallel_data(326) & xcvr_native_a10_0_rx_parallel_data(325) & xcvr_native_a10_0_rx_parallel_data(324) & xcvr_native_a10_0_rx_parallel_data(323) & xcvr_native_a10_0_rx_parallel_data(322) & xcvr_native_a10_0_rx_parallel_data(321) & xcvr_native_a10_0_rx_parallel_data(320) & xcvr_native_a10_0_rx_parallel_data(319) & xcvr_native_a10_0_rx_parallel_data(318) & xcvr_native_a10_0_rx_parallel_data(317) & xcvr_native_a10_0_rx_parallel_data(316) & xcvr_native_a10_0_rx_parallel_data(315) & xcvr_native_a10_0_rx_parallel_data(314) & xcvr_native_a10_0_rx_parallel_data(313) & xcvr_native_a10_0_rx_parallel_data(312) & xcvr_native_a10_0_rx_parallel_data(311) & xcvr_native_a10_0_rx_parallel_data(310) & xcvr_native_a10_0_rx_parallel_data(309) & xcvr_native_a10_0_rx_parallel_data(308) & xcvr_native_a10_0_rx_parallel_data(307) & xcvr_native_a10_0_rx_parallel_data(306) & xcvr_native_a10_0_rx_parallel_data(305) & xcvr_native_a10_0_rx_parallel_data(304) & xcvr_native_a10_0_rx_parallel_data(303) & xcvr_native_a10_0_rx_parallel_data(302) & xcvr_native_a10_0_rx_parallel_data(301) & xcvr_native_a10_0_rx_parallel_data(300) & xcvr_native_a10_0_rx_parallel_data(299) & xcvr_native_a10_0_rx_parallel_data(298) & xcvr_native_a10_0_rx_parallel_data(297) & xcvr_native_a10_0_rx_parallel_data(296) & xcvr_native_a10_0_rx_parallel_data(295) & xcvr_native_a10_0_rx_parallel_data(294) & xcvr_native_a10_0_rx_parallel_data(293) & xcvr_native_a10_0_rx_parallel_data(292) & xcvr_native_a10_0_rx_parallel_data(291) & xcvr_native_a10_0_rx_parallel_data(290) & xcvr_native_a10_0_rx_parallel_data(289) & xcvr_native_a10_0_rx_parallel_data(288) & xcvr_native_a10_0_rx_parallel_data(287) & xcvr_native_a10_0_rx_parallel_data(286) & xcvr_native_a10_0_rx_parallel_data(285) & xcvr_native_a10_0_rx_parallel_data(283) & xcvr_native_a10_0_rx_parallel_data(271) & xcvr_native_a10_0_rx_parallel_data(270) & xcvr_native_a10_0_rx_parallel_data(269) & xcvr_native_a10_0_rx_parallel_data(267) & xcvr_native_a10_0_rx_parallel_data(255) & xcvr_native_a10_0_rx_parallel_data(254) & xcvr_native_a10_0_rx_parallel_data(253) & xcvr_native_a10_0_rx_parallel_data(252) & xcvr_native_a10_0_rx_parallel_data(251) & xcvr_native_a10_0_rx_parallel_data(250) & xcvr_native_a10_0_rx_parallel_data(249) & xcvr_native_a10_0_rx_parallel_data(248) & xcvr_native_a10_0_rx_parallel_data(247) & xcvr_native_a10_0_rx_parallel_data(246) & xcvr_native_a10_0_rx_parallel_data(245) & xcvr_native_a10_0_rx_parallel_data(244) & xcvr_native_a10_0_rx_parallel_data(243) & xcvr_native_a10_0_rx_parallel_data(242) & xcvr_native_a10_0_rx_parallel_data(241) & xcvr_native_a10_0_rx_parallel_data(240) & xcvr_native_a10_0_rx_parallel_data(239) & xcvr_native_a10_0_rx_parallel_data(238) & xcvr_native_a10_0_rx_parallel_data(237) & xcvr_native_a10_0_rx_parallel_data(236) & xcvr_native_a10_0_rx_parallel_data(235) & xcvr_native_a10_0_rx_parallel_data(234) & xcvr_native_a10_0_rx_parallel_data(233) & xcvr_native_a10_0_rx_parallel_data(232) & xcvr_native_a10_0_rx_parallel_data(231) & xcvr_native_a10_0_rx_parallel_data(230) & xcvr_native_a10_0_rx_parallel_data(229) & xcvr_native_a10_0_rx_parallel_data(228) & xcvr_native_a10_0_rx_parallel_data(227) & xcvr_native_a10_0_rx_parallel_data(226) & xcvr_native_a10_0_rx_parallel_data(225) & xcvr_native_a10_0_rx_parallel_data(224) & xcvr_native_a10_0_rx_parallel_data(223) & xcvr_native_a10_0_rx_parallel_data(222) & xcvr_native_a10_0_rx_parallel_data(221) & xcvr_native_a10_0_rx_parallel_data(220) & xcvr_native_a10_0_rx_parallel_data(219) & xcvr_native_a10_0_rx_parallel_data(218) & xcvr_native_a10_0_rx_parallel_data(217) & xcvr_native_a10_0_rx_parallel_data(216) & xcvr_native_a10_0_rx_parallel_data(215) & xcvr_native_a10_0_rx_parallel_data(214) & xcvr_native_a10_0_rx_parallel_data(213) & xcvr_native_a10_0_rx_parallel_data(212) & xcvr_native_a10_0_rx_parallel_data(211) & xcvr_native_a10_0_rx_parallel_data(210) & xcvr_native_a10_0_rx_parallel_data(209) & xcvr_native_a10_0_rx_parallel_data(208) & xcvr_native_a10_0_rx_parallel_data(207) & xcvr_native_a10_0_rx_parallel_data(206) & xcvr_native_a10_0_rx_parallel_data(205) & xcvr_native_a10_0_rx_parallel_data(204) & xcvr_native_a10_0_rx_parallel_data(203) & xcvr_native_a10_0_rx_parallel_data(202) & xcvr_native_a10_0_rx_parallel_data(201) & xcvr_native_a10_0_rx_parallel_data(200) & xcvr_native_a10_0_rx_parallel_data(199) & xcvr_native_a10_0_rx_parallel_data(198) & xcvr_native_a10_0_rx_parallel_data(197) & xcvr_native_a10_0_rx_parallel_data(196) & xcvr_native_a10_0_rx_parallel_data(195) & xcvr_native_a10_0_rx_parallel_data(194) & xcvr_native_a10_0_rx_parallel_data(193) & xcvr_native_a10_0_rx_parallel_data(192) & xcvr_native_a10_0_rx_parallel_data(191) & xcvr_native_a10_0_rx_parallel_data(190) & xcvr_native_a10_0_rx_parallel_data(189) & xcvr_native_a10_0_rx_parallel_data(188) & xcvr_native_a10_0_rx_parallel_data(187) & xcvr_native_a10_0_rx_parallel_data(186) & xcvr_native_a10_0_rx_parallel_data(185) & xcvr_native_a10_0_rx_parallel_data(184) & xcvr_native_a10_0_rx_parallel_data(183) & xcvr_native_a10_0_rx_parallel_data(182) & xcvr_native_a10_0_rx_parallel_data(181) & xcvr_native_a10_0_rx_parallel_data(180) & xcvr_native_a10_0_rx_parallel_data(179) & xcvr_native_a10_0_rx_parallel_data(178) & xcvr_native_a10_0_rx_parallel_data(177) & xcvr_native_a10_0_rx_parallel_data(176) & xcvr_native_a10_0_rx_parallel_data(175) & xcvr_native_a10_0_rx_parallel_data(174) & xcvr_native_a10_0_rx_parallel_data(173) & xcvr_native_a10_0_rx_parallel_data(172) & xcvr_native_a10_0_rx_parallel_data(171) & xcvr_native_a10_0_rx_parallel_data(170) & xcvr_native_a10_0_rx_parallel_data(169) & xcvr_native_a10_0_rx_parallel_data(168) & xcvr_native_a10_0_rx_parallel_data(167) & xcvr_native_a10_0_rx_parallel_data(166) & xcvr_native_a10_0_rx_parallel_data(165) & xcvr_native_a10_0_rx_parallel_data(164) & xcvr_native_a10_0_rx_parallel_data(163) & xcvr_native_a10_0_rx_parallel_data(162) & xcvr_native_a10_0_rx_parallel_data(161) & xcvr_native_a10_0_rx_parallel_data(160) & xcvr_native_a10_0_rx_parallel_data(159) & xcvr_native_a10_0_rx_parallel_data(158) & xcvr_native_a10_0_rx_parallel_data(157) & xcvr_native_a10_0_rx_parallel_data(155) & xcvr_native_a10_0_rx_parallel_data(143) & xcvr_native_a10_0_rx_parallel_data(142) & xcvr_native_a10_0_rx_parallel_data(141) & xcvr_native_a10_0_rx_parallel_data(139) & xcvr_native_a10_0_rx_parallel_data(127) & xcvr_native_a10_0_rx_parallel_data(126) & xcvr_native_a10_0_rx_parallel_data(125) & xcvr_native_a10_0_rx_parallel_data(124) & xcvr_native_a10_0_rx_parallel_data(123) & xcvr_native_a10_0_rx_parallel_data(122) & xcvr_native_a10_0_rx_parallel_data(121) & xcvr_native_a10_0_rx_parallel_data(120) & xcvr_native_a10_0_rx_parallel_data(119) & xcvr_native_a10_0_rx_parallel_data(118) & xcvr_native_a10_0_rx_parallel_data(117) & xcvr_native_a10_0_rx_parallel_data(116) & xcvr_native_a10_0_rx_parallel_data(115) & xcvr_native_a10_0_rx_parallel_data(114) & xcvr_native_a10_0_rx_parallel_data(113) & xcvr_native_a10_0_rx_parallel_data(112) & xcvr_native_a10_0_rx_parallel_data(111) & xcvr_native_a10_0_rx_parallel_data(110) & xcvr_native_a10_0_rx_parallel_data(109) & xcvr_native_a10_0_rx_parallel_data(108) & xcvr_native_a10_0_rx_parallel_data(107) & xcvr_native_a10_0_rx_parallel_data(106) & xcvr_native_a10_0_rx_parallel_data(105) & xcvr_native_a10_0_rx_parallel_data(104) & xcvr_native_a10_0_rx_parallel_data(103) & xcvr_native_a10_0_rx_parallel_data(102) & xcvr_native_a10_0_rx_parallel_data(101) & xcvr_native_a10_0_rx_parallel_data(100) & xcvr_native_a10_0_rx_parallel_data(99) & xcvr_native_a10_0_rx_parallel_data(98) & xcvr_native_a10_0_rx_parallel_data(97) & xcvr_native_a10_0_rx_parallel_data(96) & xcvr_native_a10_0_rx_parallel_data(95) & xcvr_native_a10_0_rx_parallel_data(94) & xcvr_native_a10_0_rx_parallel_data(93) & xcvr_native_a10_0_rx_parallel_data(92) & xcvr_native_a10_0_rx_parallel_data(91) & xcvr_native_a10_0_rx_parallel_data(90) & xcvr_native_a10_0_rx_parallel_data(89) & xcvr_native_a10_0_rx_parallel_data(88) & xcvr_native_a10_0_rx_parallel_data(87) & xcvr_native_a10_0_rx_parallel_data(86) & xcvr_native_a10_0_rx_parallel_data(85) & xcvr_native_a10_0_rx_parallel_data(84) & xcvr_native_a10_0_rx_parallel_data(83) & xcvr_native_a10_0_rx_parallel_data(82) & xcvr_native_a10_0_rx_parallel_data(81) & xcvr_native_a10_0_rx_parallel_data(80) & xcvr_native_a10_0_rx_parallel_data(79) & xcvr_native_a10_0_rx_parallel_data(78) & xcvr_native_a10_0_rx_parallel_data(77) & xcvr_native_a10_0_rx_parallel_data(76) & xcvr_native_a10_0_rx_parallel_data(75) & xcvr_native_a10_0_rx_parallel_data(74) & xcvr_native_a10_0_rx_parallel_data(73) & xcvr_native_a10_0_rx_parallel_data(72) & xcvr_native_a10_0_rx_parallel_data(71) & xcvr_native_a10_0_rx_parallel_data(70) & xcvr_native_a10_0_rx_parallel_data(69) & xcvr_native_a10_0_rx_parallel_data(68) & xcvr_native_a10_0_rx_parallel_data(67) & xcvr_native_a10_0_rx_parallel_data(66) & xcvr_native_a10_0_rx_parallel_data(65) & xcvr_native_a10_0_rx_parallel_data(64) & xcvr_native_a10_0_rx_parallel_data(63) & xcvr_native_a10_0_rx_parallel_data(62) & xcvr_native_a10_0_rx_parallel_data(61) & xcvr_native_a10_0_rx_parallel_data(60) & xcvr_native_a10_0_rx_parallel_data(59) & xcvr_native_a10_0_rx_parallel_data(58) & xcvr_native_a10_0_rx_parallel_data(57) & xcvr_native_a10_0_rx_parallel_data(56) & xcvr_native_a10_0_rx_parallel_data(55) & xcvr_native_a10_0_rx_parallel_data(54) & xcvr_native_a10_0_rx_parallel_data(53) & xcvr_native_a10_0_rx_parallel_data(52) & xcvr_native_a10_0_rx_parallel_data(51) & xcvr_native_a10_0_rx_parallel_data(50) & xcvr_native_a10_0_rx_parallel_data(49) & xcvr_native_a10_0_rx_parallel_data(48) & xcvr_native_a10_0_rx_parallel_data(47) & xcvr_native_a10_0_rx_parallel_data(46) & xcvr_native_a10_0_rx_parallel_data(45) & xcvr_native_a10_0_rx_parallel_data(44) & xcvr_native_a10_0_rx_parallel_data(43) & xcvr_native_a10_0_rx_parallel_data(42) & xcvr_native_a10_0_rx_parallel_data(41) & xcvr_native_a10_0_rx_parallel_data(40) & xcvr_native_a10_0_rx_parallel_data(39) & xcvr_native_a10_0_rx_parallel_data(38) & xcvr_native_a10_0_rx_parallel_data(37) & xcvr_native_a10_0_rx_parallel_data(36) & xcvr_native_a10_0_rx_parallel_data(35) & xcvr_native_a10_0_rx_parallel_data(34) & xcvr_native_a10_0_rx_parallel_data(33) & xcvr_native_a10_0_rx_parallel_data(32) & xcvr_native_a10_0_rx_parallel_data(31) & xcvr_native_a10_0_rx_parallel_data(30) & xcvr_native_a10_0_rx_parallel_data(29) & xcvr_native_a10_0_rx_parallel_data(27) & xcvr_native_a10_0_rx_parallel_data(15) & xcvr_native_a10_0_rx_parallel_data(14) & xcvr_native_a10_0_rx_parallel_data(13) & xcvr_native_a10_0_rx_parallel_data(11);

	xcvr_reset_control_0_rx_ready0_rx_ready <= xcvr_reset_control_0_rx_ready(0);

	xcvr_reset_control_0_rx_ready1_rx_ready <= xcvr_reset_control_0_rx_ready(1);

	xcvr_reset_control_0_rx_ready2_rx_ready <= xcvr_reset_control_0_rx_ready(2);

	xcvr_reset_control_0_rx_ready3_rx_ready <= xcvr_reset_control_0_rx_ready(3);

	xcvr_reset_control_0_tx_ready0_tx_ready <= xcvr_reset_control_0_tx_ready(0);

	xcvr_reset_control_0_tx_ready1_tx_ready <= xcvr_reset_control_0_tx_ready(1);

	xcvr_reset_control_0_tx_ready2_tx_ready <= xcvr_reset_control_0_tx_ready(2);

	xcvr_reset_control_0_tx_ready3_tx_ready <= xcvr_reset_control_0_tx_ready(3);

	xcvr_reset_control_0_pll_powerdown0_pll_powerdown <= xcvr_reset_control_0_pll_powerdown(0);

	xcvr_reset_control_0_rx_analogreset0_rx_analogreset <= xcvr_reset_control_0_rx_analogreset(0);

	xcvr_reset_control_0_rx_analogreset1_rx_analogreset <= xcvr_reset_control_0_rx_analogreset(1);

	xcvr_reset_control_0_rx_analogreset3_rx_analogreset <= xcvr_reset_control_0_rx_analogreset(3);

	xcvr_reset_control_0_rx_analogreset2_rx_analogreset <= xcvr_reset_control_0_rx_analogreset(2);

	xcvr_native_a10_0_rx_cal_busy_ch0_rx_cal_busy <= xcvr_native_a10_0_rx_cal_busy(0);

	xcvr_native_a10_0_rx_cal_busy_ch2_rx_cal_busy <= xcvr_native_a10_0_rx_cal_busy(2);

	xcvr_native_a10_0_rx_cal_busy_ch1_rx_cal_busy <= xcvr_native_a10_0_rx_cal_busy(1);

	xcvr_native_a10_0_rx_cal_busy_ch3_rx_cal_busy <= xcvr_native_a10_0_rx_cal_busy(3);

	xcvr_reset_control_0_rx_digitalreset0_rx_digitalreset <= xcvr_reset_control_0_rx_digitalreset(0);

	xcvr_reset_control_0_rx_digitalreset2_rx_digitalreset <= xcvr_reset_control_0_rx_digitalreset(2);

	xcvr_reset_control_0_rx_digitalreset1_rx_digitalreset <= xcvr_reset_control_0_rx_digitalreset(1);

	xcvr_reset_control_0_rx_digitalreset3_rx_digitalreset <= xcvr_reset_control_0_rx_digitalreset(3);

	xcvr_native_a10_0_rx_is_lockedtodata_ch1_rx_is_lockedtodata <= xcvr_native_a10_0_rx_is_lockedtodata(1);

	xcvr_native_a10_0_rx_is_lockedtodata_ch3_rx_is_lockedtodata <= xcvr_native_a10_0_rx_is_lockedtodata(3);

	xcvr_native_a10_0_rx_is_lockedtodata_ch0_rx_is_lockedtodata <= xcvr_native_a10_0_rx_is_lockedtodata(0);

	xcvr_native_a10_0_rx_is_lockedtodata_ch2_rx_is_lockedtodata <= xcvr_native_a10_0_rx_is_lockedtodata(2);

	xcvr_reset_control_0_tx_analogreset0_tx_analogreset <= xcvr_reset_control_0_tx_analogreset(0);

	xcvr_reset_control_0_tx_analogreset2_tx_analogreset <= xcvr_reset_control_0_tx_analogreset(2);

	xcvr_reset_control_0_tx_analogreset1_tx_analogreset <= xcvr_reset_control_0_tx_analogreset(1);

	xcvr_reset_control_0_tx_analogreset3_tx_analogreset <= xcvr_reset_control_0_tx_analogreset(3);

	xcvr_native_a10_0_tx_cal_busy_ch0_tx_cal_busy <= xcvr_native_a10_0_tx_cal_busy(0);

	xcvr_native_a10_0_tx_cal_busy_ch2_tx_cal_busy <= xcvr_native_a10_0_tx_cal_busy(2);

	xcvr_native_a10_0_tx_cal_busy_ch1_tx_cal_busy <= xcvr_native_a10_0_tx_cal_busy(1);

	xcvr_native_a10_0_tx_cal_busy_ch3_tx_cal_busy <= xcvr_native_a10_0_tx_cal_busy(3);

	xcvr_reset_control_0_tx_digitalreset0_tx_digitalreset <= xcvr_reset_control_0_tx_digitalreset(0);

	xcvr_reset_control_0_tx_digitalreset2_tx_digitalreset <= xcvr_reset_control_0_tx_digitalreset(2);

	xcvr_reset_control_0_tx_digitalreset1_tx_digitalreset <= xcvr_reset_control_0_tx_digitalreset(1);

	xcvr_reset_control_0_tx_digitalreset3_tx_digitalreset <= xcvr_reset_control_0_tx_digitalreset(3);

end architecture rtl; -- of xcvr_8B10B
